VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r1
  CLASS BLOCK ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.725 BY 12.455 ;
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 18.465 8.225 18.635 9.495 ;
        RECT 29.690 8.230 29.860 9.500 ;
        RECT 29.690 2.960 29.860 4.230 ;
      LAYER met1 ;
        RECT 18.380 8.400 18.720 8.450 ;
        RECT 18.380 8.395 18.725 8.400 ;
        RECT 18.380 8.365 18.865 8.395 ;
        RECT 20.690 8.365 21.030 8.455 ;
        RECT 18.380 8.190 21.030 8.365 ;
        RECT 18.380 8.170 18.720 8.190 ;
        RECT 20.690 8.175 21.030 8.190 ;
        RECT 29.620 8.400 29.945 8.475 ;
        RECT 29.620 8.230 30.090 8.400 ;
        RECT 29.620 8.150 29.945 8.230 ;
        RECT 29.615 4.930 29.940 5.255 ;
        RECT 29.690 4.260 29.870 4.930 ;
        RECT 29.630 4.230 29.920 4.260 ;
        RECT 29.630 4.060 30.090 4.230 ;
        RECT 29.630 4.030 29.920 4.060 ;
      LAYER met2 ;
        RECT 20.775 9.315 29.860 9.485 ;
        RECT 18.410 8.125 18.690 8.495 ;
        RECT 20.775 8.485 20.945 9.315 ;
        RECT 20.720 8.145 21.000 8.485 ;
        RECT 29.685 8.475 29.860 9.315 ;
        RECT 29.620 8.150 29.945 8.475 ;
        RECT 29.685 5.255 29.860 8.150 ;
        RECT 29.615 4.930 29.940 5.255 ;
      LAYER met3 ;
        RECT 18.380 8.125 18.720 12.455 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 35.050 8.225 35.220 9.495 ;
        RECT 46.275 8.230 46.445 9.500 ;
        RECT 46.275 2.960 46.445 4.230 ;
      LAYER met1 ;
        RECT 34.965 8.400 35.305 8.450 ;
        RECT 34.965 8.395 35.310 8.400 ;
        RECT 34.965 8.365 35.450 8.395 ;
        RECT 37.275 8.365 37.615 8.455 ;
        RECT 34.965 8.190 37.615 8.365 ;
        RECT 34.965 8.170 35.305 8.190 ;
        RECT 37.275 8.175 37.615 8.190 ;
        RECT 46.205 8.400 46.530 8.475 ;
        RECT 46.205 8.230 46.675 8.400 ;
        RECT 46.205 8.150 46.530 8.230 ;
        RECT 46.200 4.930 46.525 5.255 ;
        RECT 46.275 4.260 46.455 4.930 ;
        RECT 46.215 4.230 46.505 4.260 ;
        RECT 46.215 4.060 46.675 4.230 ;
        RECT 46.215 4.030 46.505 4.060 ;
      LAYER met2 ;
        RECT 37.360 9.315 46.445 9.485 ;
        RECT 34.995 8.125 35.275 8.495 ;
        RECT 37.360 8.485 37.530 9.315 ;
        RECT 37.305 8.145 37.585 8.485 ;
        RECT 46.270 8.475 46.445 9.315 ;
        RECT 46.205 8.150 46.530 8.475 ;
        RECT 46.270 5.255 46.445 8.150 ;
        RECT 46.200 4.930 46.525 5.255 ;
      LAYER met3 ;
        RECT 34.965 8.125 35.305 12.455 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 51.635 8.225 51.805 9.495 ;
        RECT 62.860 8.230 63.030 9.500 ;
        RECT 62.860 2.960 63.030 4.230 ;
      LAYER met1 ;
        RECT 51.550 8.400 51.890 8.450 ;
        RECT 51.550 8.395 51.895 8.400 ;
        RECT 51.550 8.365 52.035 8.395 ;
        RECT 53.860 8.365 54.200 8.455 ;
        RECT 51.550 8.190 54.200 8.365 ;
        RECT 51.550 8.170 51.890 8.190 ;
        RECT 53.860 8.175 54.200 8.190 ;
        RECT 62.790 8.400 63.115 8.475 ;
        RECT 62.790 8.230 63.260 8.400 ;
        RECT 62.790 8.150 63.115 8.230 ;
        RECT 62.785 4.930 63.110 5.255 ;
        RECT 62.860 4.260 63.040 4.930 ;
        RECT 62.800 4.230 63.090 4.260 ;
        RECT 62.800 4.060 63.260 4.230 ;
        RECT 62.800 4.030 63.090 4.060 ;
      LAYER met2 ;
        RECT 53.945 9.315 63.030 9.485 ;
        RECT 51.580 8.125 51.860 8.495 ;
        RECT 53.945 8.485 54.115 9.315 ;
        RECT 53.890 8.145 54.170 8.485 ;
        RECT 62.855 8.475 63.030 9.315 ;
        RECT 62.790 8.150 63.115 8.475 ;
        RECT 62.855 5.255 63.030 8.150 ;
        RECT 62.785 4.930 63.110 5.255 ;
      LAYER met3 ;
        RECT 51.550 8.125 51.890 12.455 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 68.220 8.225 68.390 9.495 ;
        RECT 79.445 8.230 79.615 9.500 ;
        RECT 79.445 2.960 79.615 4.230 ;
      LAYER met1 ;
        RECT 68.135 8.400 68.475 8.450 ;
        RECT 68.135 8.395 68.480 8.400 ;
        RECT 68.135 8.365 68.620 8.395 ;
        RECT 70.445 8.365 70.785 8.455 ;
        RECT 68.135 8.190 70.785 8.365 ;
        RECT 68.135 8.170 68.475 8.190 ;
        RECT 70.445 8.175 70.785 8.190 ;
        RECT 79.375 8.400 79.700 8.475 ;
        RECT 79.375 8.230 79.845 8.400 ;
        RECT 79.375 8.150 79.700 8.230 ;
        RECT 79.370 4.930 79.695 5.255 ;
        RECT 79.445 4.260 79.625 4.930 ;
        RECT 79.385 4.230 79.675 4.260 ;
        RECT 79.385 4.060 79.845 4.230 ;
        RECT 79.385 4.030 79.675 4.060 ;
      LAYER met2 ;
        RECT 70.530 9.315 79.615 9.485 ;
        RECT 68.165 8.125 68.445 8.495 ;
        RECT 70.530 8.485 70.700 9.315 ;
        RECT 70.475 8.145 70.755 8.485 ;
        RECT 79.440 8.475 79.615 9.315 ;
        RECT 79.375 8.150 79.700 8.475 ;
        RECT 79.440 5.255 79.615 8.150 ;
        RECT 79.370 4.930 79.695 5.255 ;
      LAYER met3 ;
        RECT 68.135 8.125 68.475 12.455 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 84.800 8.225 84.970 9.495 ;
        RECT 96.025 8.230 96.195 9.500 ;
        RECT 96.025 2.960 96.195 4.230 ;
      LAYER met1 ;
        RECT 84.715 8.400 85.055 8.450 ;
        RECT 84.715 8.395 85.060 8.400 ;
        RECT 84.715 8.365 85.200 8.395 ;
        RECT 87.025 8.365 87.365 8.455 ;
        RECT 84.715 8.190 87.365 8.365 ;
        RECT 84.715 8.170 85.055 8.190 ;
        RECT 87.025 8.175 87.365 8.190 ;
        RECT 95.955 8.400 96.280 8.475 ;
        RECT 95.955 8.230 96.425 8.400 ;
        RECT 95.955 8.150 96.280 8.230 ;
        RECT 95.950 4.930 96.275 5.255 ;
        RECT 96.025 4.260 96.205 4.930 ;
        RECT 95.965 4.230 96.255 4.260 ;
        RECT 95.965 4.060 96.425 4.230 ;
        RECT 95.965 4.030 96.255 4.060 ;
      LAYER met2 ;
        RECT 87.110 9.315 96.195 9.485 ;
        RECT 84.745 8.125 85.025 8.495 ;
        RECT 87.110 8.485 87.280 9.315 ;
        RECT 87.055 8.145 87.335 8.485 ;
        RECT 96.020 8.475 96.195 9.315 ;
        RECT 95.955 8.150 96.280 8.475 ;
        RECT 96.020 5.255 96.195 8.150 ;
        RECT 95.950 4.930 96.275 5.255 ;
      LAYER met3 ;
        RECT 84.715 8.125 85.055 12.455 ;
    END
  END s5
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 100.180 4.015 100.355 5.160 ;
        RECT 100.180 3.580 100.350 4.015 ;
        RECT 100.185 1.870 100.355 2.380 ;
      LAYER met1 ;
        RECT 100.120 3.545 100.410 3.780 ;
        RECT 100.120 3.540 100.350 3.545 ;
        RECT 100.180 2.440 100.350 3.540 ;
        RECT 100.120 2.180 100.415 2.440 ;
    END
  END X5_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 83.600 4.015 83.775 5.160 ;
        RECT 83.600 3.580 83.770 4.015 ;
        RECT 83.605 1.870 83.775 2.380 ;
      LAYER met1 ;
        RECT 83.540 3.545 83.830 3.780 ;
        RECT 83.540 3.540 83.770 3.545 ;
        RECT 83.600 2.440 83.770 3.540 ;
        RECT 83.540 2.180 83.835 2.440 ;
    END
  END X4_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 67.015 4.015 67.190 5.160 ;
        RECT 67.015 3.580 67.185 4.015 ;
        RECT 67.020 1.870 67.190 2.380 ;
      LAYER met1 ;
        RECT 66.955 3.545 67.245 3.780 ;
        RECT 66.955 3.540 67.185 3.545 ;
        RECT 67.015 2.440 67.185 3.540 ;
        RECT 66.955 2.180 67.250 2.440 ;
    END
  END X3_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 50.430 4.015 50.605 5.160 ;
        RECT 50.430 3.580 50.600 4.015 ;
        RECT 50.435 1.870 50.605 2.380 ;
      LAYER met1 ;
        RECT 50.370 3.545 50.660 3.780 ;
        RECT 50.370 3.540 50.600 3.545 ;
        RECT 50.430 2.440 50.600 3.540 ;
        RECT 50.370 2.180 50.665 2.440 ;
    END
  END X2_Y1
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 33.845 4.015 34.020 5.160 ;
        RECT 33.845 3.580 34.015 4.015 ;
        RECT 33.850 1.870 34.020 2.380 ;
      LAYER met1 ;
        RECT 33.785 3.545 34.075 3.780 ;
        RECT 33.785 3.540 34.015 3.545 ;
        RECT 33.845 2.440 34.015 3.540 ;
        RECT 33.785 2.180 34.080 2.440 ;
    END
  END X1_Y1
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 15.235 8.225 15.405 9.495 ;
      LAYER met1 ;
        RECT 15.175 8.395 15.470 8.425 ;
        RECT 15.175 8.225 15.635 8.395 ;
        RECT 15.175 8.195 15.470 8.225 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 17.765 8.735 21.310 8.740 ;
        RECT 14.985 8.130 21.310 8.735 ;
        RECT 28.535 8.130 37.895 8.740 ;
        RECT 45.120 8.130 54.480 8.740 ;
        RECT 61.705 8.130 71.065 8.740 ;
        RECT 78.290 8.130 87.645 8.740 ;
        RECT 14.985 7.620 21.330 8.130 ;
        RECT 14.995 7.135 21.330 7.620 ;
        RECT 28.535 7.135 37.915 8.130 ;
        RECT 45.120 7.135 54.500 8.130 ;
        RECT 61.705 7.135 71.085 8.130 ;
        RECT 78.290 7.135 87.665 8.130 ;
        RECT 94.870 7.135 100.725 8.740 ;
        RECT 14.995 5.425 100.725 7.135 ;
        RECT 14.985 4.305 100.725 5.425 ;
        RECT 14.985 3.715 21.005 4.305 ;
        RECT 28.695 3.720 37.590 4.305 ;
        RECT 45.280 3.720 54.175 4.305 ;
        RECT 61.865 3.720 70.760 4.305 ;
        RECT 78.450 3.720 87.340 4.305 ;
        RECT 95.030 3.720 100.725 4.305 ;
        RECT 34.240 3.715 37.590 3.720 ;
        RECT 50.810 3.715 54.175 3.720 ;
        RECT 67.405 3.715 70.760 3.720 ;
        RECT 83.960 3.715 87.340 3.720 ;
        RECT 17.800 3.710 20.775 3.715 ;
        RECT 34.385 3.710 37.360 3.715 ;
        RECT 50.810 3.710 53.945 3.715 ;
        RECT 67.405 3.710 70.530 3.715 ;
        RECT 83.960 3.710 87.110 3.715 ;
      LAYER li1 ;
        RECT 17.040 10.035 17.215 10.585 ;
        RECT 17.040 8.435 17.210 10.035 ;
        RECT 15.225 7.025 15.395 7.755 ;
        RECT 17.040 7.295 17.215 8.435 ;
        RECT 17.040 7.025 17.210 7.295 ;
        RECT 18.455 7.025 18.625 7.755 ;
        RECT 29.680 7.030 29.850 7.760 ;
        RECT 32.425 7.030 32.595 7.760 ;
        RECT 33.415 7.030 33.585 7.760 ;
        RECT 35.040 7.030 35.210 7.755 ;
        RECT 46.265 7.030 46.435 7.760 ;
        RECT 49.010 7.030 49.180 7.760 ;
        RECT 50.000 7.030 50.170 7.760 ;
        RECT 51.625 7.030 51.795 7.755 ;
        RECT 62.850 7.030 63.020 7.760 ;
        RECT 65.595 7.030 65.765 7.760 ;
        RECT 66.585 7.030 66.755 7.760 ;
        RECT 68.210 7.030 68.380 7.755 ;
        RECT 79.435 7.030 79.605 7.760 ;
        RECT 82.180 7.030 82.350 7.760 ;
        RECT 83.170 7.030 83.340 7.760 ;
        RECT 84.790 7.030 84.960 7.755 ;
        RECT 96.015 7.030 96.185 7.760 ;
        RECT 98.760 7.030 98.930 7.760 ;
        RECT 99.750 7.030 99.920 7.760 ;
        RECT 0.000 5.805 21.620 7.025 ;
        RECT 22.710 5.805 23.040 6.525 ;
        RECT 23.725 5.805 24.005 6.265 ;
        RECT 24.870 5.805 25.140 6.585 ;
        RECT 25.690 5.805 26.060 6.185 ;
        RECT 28.450 5.965 38.205 7.030 ;
        RECT 28.320 5.805 38.205 5.965 ;
        RECT 39.295 5.805 39.625 6.525 ;
        RECT 40.310 5.805 40.590 6.265 ;
        RECT 41.455 5.805 41.725 6.585 ;
        RECT 42.275 5.805 42.645 6.185 ;
        RECT 45.035 5.965 54.790 7.030 ;
        RECT 44.905 5.805 54.790 5.965 ;
        RECT 55.880 5.805 56.210 6.525 ;
        RECT 56.895 5.805 57.175 6.265 ;
        RECT 58.040 5.805 58.310 6.585 ;
        RECT 58.860 5.805 59.230 6.185 ;
        RECT 61.620 5.965 71.375 7.030 ;
        RECT 61.490 5.805 71.375 5.965 ;
        RECT 72.465 5.805 72.795 6.525 ;
        RECT 73.480 5.805 73.760 6.265 ;
        RECT 74.625 5.805 74.895 6.585 ;
        RECT 75.445 5.805 75.815 6.185 ;
        RECT 78.205 5.965 87.960 7.030 ;
        RECT 78.075 5.805 87.960 5.965 ;
        RECT 89.045 5.805 89.375 6.525 ;
        RECT 90.060 5.805 90.340 6.265 ;
        RECT 91.205 5.805 91.475 6.585 ;
        RECT 92.025 5.805 92.395 6.185 ;
        RECT 94.785 5.965 100.725 7.030 ;
        RECT 94.655 5.805 100.725 5.965 ;
        RECT 0.000 5.635 100.725 5.805 ;
        RECT 0.000 5.425 21.620 5.635 ;
        RECT 21.295 5.125 21.555 5.425 ;
        RECT 22.520 5.135 23.140 5.635 ;
        RECT 22.940 4.955 23.140 5.135 ;
        RECT 23.950 5.095 24.170 5.635 ;
        RECT 24.820 4.985 25.430 5.635 ;
        RECT 26.250 5.095 26.510 5.635 ;
        RECT 27.990 5.430 38.205 5.635 ;
        RECT 25.250 4.955 25.440 4.985 ;
        RECT 22.940 4.765 23.270 4.955 ;
        RECT 25.250 4.715 25.580 4.955 ;
        RECT 27.990 4.495 28.320 5.430 ;
        RECT 29.680 4.700 29.850 5.430 ;
        RECT 32.425 4.700 32.595 5.430 ;
        RECT 33.415 4.700 33.585 5.430 ;
        RECT 34.225 5.425 38.205 5.430 ;
        RECT 37.880 5.125 38.140 5.425 ;
        RECT 39.105 5.135 39.725 5.635 ;
        RECT 39.525 4.955 39.725 5.135 ;
        RECT 40.535 5.095 40.755 5.635 ;
        RECT 41.405 4.985 42.015 5.635 ;
        RECT 42.835 5.095 43.095 5.635 ;
        RECT 44.575 5.430 54.790 5.635 ;
        RECT 41.835 4.955 42.025 4.985 ;
        RECT 39.525 4.765 39.855 4.955 ;
        RECT 41.835 4.715 42.165 4.955 ;
        RECT 44.575 4.495 44.905 5.430 ;
        RECT 46.265 4.700 46.435 5.430 ;
        RECT 49.010 4.700 49.180 5.430 ;
        RECT 50.000 4.700 50.170 5.430 ;
        RECT 50.805 5.425 54.790 5.430 ;
        RECT 54.465 5.125 54.725 5.425 ;
        RECT 55.690 5.135 56.310 5.635 ;
        RECT 56.110 4.955 56.310 5.135 ;
        RECT 57.120 5.095 57.340 5.635 ;
        RECT 57.990 4.985 58.600 5.635 ;
        RECT 59.420 5.095 59.680 5.635 ;
        RECT 61.160 5.430 71.375 5.635 ;
        RECT 58.420 4.955 58.610 4.985 ;
        RECT 56.110 4.765 56.440 4.955 ;
        RECT 58.420 4.715 58.750 4.955 ;
        RECT 61.160 4.495 61.490 5.430 ;
        RECT 62.850 4.700 63.020 5.430 ;
        RECT 65.595 4.700 65.765 5.430 ;
        RECT 66.585 4.700 66.755 5.430 ;
        RECT 67.385 5.425 71.375 5.430 ;
        RECT 71.050 5.125 71.310 5.425 ;
        RECT 72.275 5.135 72.895 5.635 ;
        RECT 72.695 4.955 72.895 5.135 ;
        RECT 73.705 5.095 73.925 5.635 ;
        RECT 74.575 4.985 75.185 5.635 ;
        RECT 76.005 5.095 76.265 5.635 ;
        RECT 77.745 5.430 87.960 5.635 ;
        RECT 75.005 4.955 75.195 4.985 ;
        RECT 72.695 4.765 73.025 4.955 ;
        RECT 75.005 4.715 75.335 4.955 ;
        RECT 77.745 4.495 78.075 5.430 ;
        RECT 79.435 4.700 79.605 5.430 ;
        RECT 82.180 4.700 82.350 5.430 ;
        RECT 83.170 4.700 83.340 5.430 ;
        RECT 83.965 5.425 87.955 5.430 ;
        RECT 87.630 5.125 87.890 5.425 ;
        RECT 88.855 5.135 89.475 5.635 ;
        RECT 89.275 4.955 89.475 5.135 ;
        RECT 90.285 5.095 90.505 5.635 ;
        RECT 91.155 4.985 91.765 5.635 ;
        RECT 92.585 5.095 92.845 5.635 ;
        RECT 94.325 5.430 100.725 5.635 ;
        RECT 91.585 4.955 91.775 4.985 ;
        RECT 89.275 4.765 89.605 4.955 ;
        RECT 91.585 4.715 91.915 4.955 ;
        RECT 94.325 4.495 94.655 5.430 ;
        RECT 96.015 4.700 96.185 5.430 ;
        RECT 98.760 4.700 98.930 5.430 ;
        RECT 99.750 4.700 99.920 5.430 ;
      LAYER met1 ;
        RECT 16.980 9.135 17.270 9.165 ;
        RECT 16.810 8.965 17.270 9.135 ;
        RECT 16.980 8.935 17.270 8.965 ;
        RECT 0.000 5.965 21.620 7.025 ;
        RECT 23.130 5.965 23.280 5.970 ;
        RECT 28.450 5.965 38.205 7.030 ;
        RECT 39.715 5.965 39.865 5.970 ;
        RECT 45.035 5.965 54.790 7.030 ;
        RECT 56.300 5.965 56.450 5.970 ;
        RECT 61.620 5.965 71.375 7.030 ;
        RECT 72.885 5.965 73.035 5.970 ;
        RECT 78.205 5.965 87.960 7.030 ;
        RECT 89.465 5.965 89.615 5.970 ;
        RECT 94.785 5.965 100.725 7.030 ;
        RECT 0.000 5.485 100.725 5.965 ;
        RECT 0.000 5.425 21.620 5.485 ;
        RECT 28.320 5.430 38.205 5.485 ;
        RECT 44.905 5.430 54.790 5.485 ;
        RECT 61.490 5.430 71.375 5.485 ;
        RECT 78.075 5.430 87.960 5.485 ;
        RECT 94.655 5.430 100.725 5.485 ;
        RECT 34.225 5.425 38.205 5.430 ;
        RECT 50.805 5.425 54.790 5.430 ;
        RECT 67.385 5.425 71.375 5.430 ;
        RECT 83.965 5.425 87.955 5.430 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.055 10.855 100.725 12.455 ;
        RECT 15.225 10.225 15.395 10.855 ;
        RECT 18.455 10.225 18.625 10.855 ;
        RECT 19.410 10.305 19.580 10.585 ;
        RECT 19.410 10.135 19.640 10.305 ;
        RECT 19.470 8.525 19.640 10.135 ;
        RECT 21.515 8.525 21.765 10.855 ;
        RECT 22.040 8.525 22.315 10.855 ;
        RECT 22.590 8.525 22.865 10.855 ;
        RECT 23.140 8.525 23.415 10.855 ;
        RECT 23.690 8.525 23.965 10.855 ;
        RECT 24.240 8.525 24.515 10.855 ;
        RECT 24.790 8.525 25.065 10.855 ;
        RECT 25.340 8.525 25.615 10.855 ;
        RECT 25.890 8.525 26.165 10.855 ;
        RECT 26.440 8.525 26.715 10.855 ;
        RECT 26.990 8.525 27.265 10.855 ;
        RECT 27.540 8.525 27.815 10.855 ;
        RECT 28.090 8.525 28.435 10.855 ;
        RECT 29.680 10.230 29.850 10.855 ;
        RECT 32.425 10.230 32.595 10.855 ;
        RECT 33.415 10.230 33.585 10.855 ;
        RECT 35.040 10.225 35.210 10.855 ;
        RECT 35.995 10.305 36.165 10.585 ;
        RECT 35.995 10.135 36.225 10.305 ;
        RECT 36.055 8.525 36.225 10.135 ;
        RECT 38.100 8.525 38.350 10.855 ;
        RECT 38.625 8.525 38.900 10.855 ;
        RECT 39.175 8.525 39.450 10.855 ;
        RECT 39.725 8.525 40.000 10.855 ;
        RECT 40.275 8.525 40.550 10.855 ;
        RECT 40.825 8.525 41.100 10.855 ;
        RECT 41.375 8.525 41.650 10.855 ;
        RECT 41.925 8.525 42.200 10.855 ;
        RECT 42.475 8.525 42.750 10.855 ;
        RECT 43.025 8.525 43.300 10.855 ;
        RECT 43.575 8.525 43.850 10.855 ;
        RECT 44.125 8.525 44.400 10.855 ;
        RECT 44.675 8.525 45.020 10.855 ;
        RECT 46.265 10.230 46.435 10.855 ;
        RECT 49.010 10.230 49.180 10.855 ;
        RECT 50.000 10.230 50.170 10.855 ;
        RECT 51.625 10.225 51.795 10.855 ;
        RECT 52.580 10.305 52.750 10.585 ;
        RECT 52.580 10.135 52.810 10.305 ;
        RECT 52.640 8.525 52.810 10.135 ;
        RECT 54.685 8.525 54.935 10.855 ;
        RECT 55.210 8.525 55.485 10.855 ;
        RECT 55.760 8.525 56.035 10.855 ;
        RECT 56.310 8.525 56.585 10.855 ;
        RECT 56.860 8.525 57.135 10.855 ;
        RECT 57.410 8.525 57.685 10.855 ;
        RECT 57.960 8.525 58.235 10.855 ;
        RECT 58.510 8.525 58.785 10.855 ;
        RECT 59.060 8.525 59.335 10.855 ;
        RECT 59.610 8.525 59.885 10.855 ;
        RECT 60.160 8.525 60.435 10.855 ;
        RECT 60.710 8.525 60.985 10.855 ;
        RECT 61.260 8.525 61.605 10.855 ;
        RECT 62.850 10.230 63.020 10.855 ;
        RECT 65.595 10.230 65.765 10.855 ;
        RECT 66.585 10.230 66.755 10.855 ;
        RECT 68.210 10.225 68.380 10.855 ;
        RECT 69.165 10.305 69.335 10.585 ;
        RECT 69.165 10.135 69.395 10.305 ;
        RECT 69.225 8.525 69.395 10.135 ;
        RECT 71.270 8.525 71.520 10.855 ;
        RECT 71.795 8.525 72.070 10.855 ;
        RECT 72.345 8.525 72.620 10.855 ;
        RECT 72.895 8.525 73.170 10.855 ;
        RECT 73.445 8.525 73.720 10.855 ;
        RECT 73.995 8.525 74.270 10.855 ;
        RECT 74.545 8.525 74.820 10.855 ;
        RECT 75.095 8.525 75.370 10.855 ;
        RECT 75.645 8.525 75.920 10.855 ;
        RECT 76.195 8.525 76.470 10.855 ;
        RECT 76.745 8.525 77.020 10.855 ;
        RECT 77.295 8.525 77.570 10.855 ;
        RECT 77.845 8.525 78.190 10.855 ;
        RECT 79.435 10.230 79.605 10.855 ;
        RECT 82.180 10.230 82.350 10.855 ;
        RECT 83.170 10.230 83.340 10.855 ;
        RECT 84.790 10.225 84.960 10.855 ;
        RECT 85.745 10.305 85.915 10.585 ;
        RECT 85.745 10.135 85.975 10.305 ;
        RECT 85.805 8.525 85.975 10.135 ;
        RECT 87.850 8.525 88.100 10.855 ;
        RECT 88.375 8.525 88.650 10.855 ;
        RECT 88.925 8.525 89.200 10.855 ;
        RECT 89.475 8.525 89.750 10.855 ;
        RECT 90.025 8.525 90.300 10.855 ;
        RECT 90.575 8.525 90.850 10.855 ;
        RECT 91.125 8.525 91.400 10.855 ;
        RECT 91.675 8.525 91.950 10.855 ;
        RECT 92.225 8.525 92.500 10.855 ;
        RECT 92.775 8.525 93.050 10.855 ;
        RECT 93.325 8.525 93.600 10.855 ;
        RECT 93.875 8.525 94.150 10.855 ;
        RECT 94.425 8.525 94.770 10.855 ;
        RECT 96.015 10.230 96.185 10.855 ;
        RECT 98.760 10.230 98.930 10.855 ;
        RECT 99.750 10.230 99.920 10.855 ;
        RECT 19.410 8.355 19.640 8.525 ;
        RECT 21.380 8.355 28.435 8.525 ;
        RECT 35.995 8.355 36.225 8.525 ;
        RECT 37.965 8.355 45.020 8.525 ;
        RECT 52.580 8.355 52.810 8.525 ;
        RECT 54.550 8.355 61.605 8.525 ;
        RECT 69.165 8.355 69.395 8.525 ;
        RECT 71.135 8.355 78.190 8.525 ;
        RECT 85.745 8.355 85.975 8.525 ;
        RECT 87.715 8.355 94.770 8.525 ;
        RECT 19.410 7.295 19.580 8.355 ;
        RECT 22.790 7.895 23.040 8.355 ;
        RECT 24.860 7.955 25.190 8.355 ;
        RECT 26.950 7.845 27.400 8.355 ;
        RECT 22.940 7.115 23.280 7.365 ;
        RECT 25.160 7.115 25.490 7.445 ;
        RECT 35.995 7.295 36.165 8.355 ;
        RECT 39.375 7.895 39.625 8.355 ;
        RECT 41.445 7.955 41.775 8.355 ;
        RECT 43.535 7.845 43.985 8.355 ;
        RECT 39.525 7.115 39.865 7.365 ;
        RECT 41.745 7.115 42.075 7.445 ;
        RECT 52.580 7.295 52.750 8.355 ;
        RECT 55.960 7.895 56.210 8.355 ;
        RECT 58.030 7.955 58.360 8.355 ;
        RECT 60.120 7.845 60.570 8.355 ;
        RECT 56.110 7.115 56.450 7.365 ;
        RECT 58.330 7.115 58.660 7.445 ;
        RECT 69.165 7.295 69.335 8.355 ;
        RECT 72.545 7.895 72.795 8.355 ;
        RECT 74.615 7.955 74.945 8.355 ;
        RECT 76.705 7.845 77.155 8.355 ;
        RECT 72.695 7.115 73.035 7.365 ;
        RECT 74.915 7.115 75.245 7.445 ;
        RECT 85.745 7.295 85.915 8.355 ;
        RECT 89.125 7.895 89.375 8.355 ;
        RECT 91.195 7.955 91.525 8.355 ;
        RECT 93.285 7.845 93.735 8.355 ;
        RECT 89.275 7.115 89.615 7.365 ;
        RECT 91.495 7.115 91.825 7.445 ;
      LAYER met1 ;
        RECT 0.055 10.855 100.725 12.455 ;
        RECT 19.245 8.805 19.415 10.855 ;
        RECT 19.245 8.775 19.700 8.805 ;
        RECT 19.235 8.605 19.700 8.775 ;
        RECT 21.515 8.685 21.765 10.855 ;
        RECT 22.040 8.685 22.315 10.855 ;
        RECT 22.590 8.685 22.865 10.855 ;
        RECT 23.140 8.685 23.415 10.855 ;
        RECT 23.690 8.685 23.965 10.855 ;
        RECT 24.240 8.685 24.515 10.855 ;
        RECT 24.790 8.685 25.065 10.855 ;
        RECT 25.340 8.685 25.615 10.855 ;
        RECT 25.890 8.685 26.165 10.855 ;
        RECT 26.440 8.685 26.715 10.855 ;
        RECT 26.990 8.685 27.265 10.855 ;
        RECT 27.540 8.685 27.815 10.855 ;
        RECT 28.090 8.685 28.435 10.855 ;
        RECT 35.830 8.805 36.000 10.855 ;
        RECT 35.830 8.775 36.285 8.805 ;
        RECT 19.245 8.600 19.700 8.605 ;
        RECT 19.410 8.575 19.700 8.600 ;
        RECT 21.380 8.325 28.435 8.685 ;
        RECT 35.820 8.605 36.285 8.775 ;
        RECT 38.100 8.685 38.350 10.855 ;
        RECT 38.625 8.685 38.900 10.855 ;
        RECT 39.175 8.685 39.450 10.855 ;
        RECT 39.725 8.685 40.000 10.855 ;
        RECT 40.275 8.685 40.550 10.855 ;
        RECT 40.825 8.685 41.100 10.855 ;
        RECT 41.375 8.685 41.650 10.855 ;
        RECT 41.925 8.685 42.200 10.855 ;
        RECT 42.475 8.685 42.750 10.855 ;
        RECT 43.025 8.685 43.300 10.855 ;
        RECT 43.575 8.685 43.850 10.855 ;
        RECT 44.125 8.685 44.400 10.855 ;
        RECT 44.675 8.685 45.020 10.855 ;
        RECT 52.415 8.805 52.585 10.855 ;
        RECT 52.415 8.775 52.870 8.805 ;
        RECT 35.830 8.600 36.285 8.605 ;
        RECT 35.995 8.575 36.285 8.600 ;
        RECT 37.965 8.325 45.020 8.685 ;
        RECT 52.405 8.605 52.870 8.775 ;
        RECT 54.685 8.685 54.935 10.855 ;
        RECT 55.210 8.685 55.485 10.855 ;
        RECT 55.760 8.685 56.035 10.855 ;
        RECT 56.310 8.685 56.585 10.855 ;
        RECT 56.860 8.685 57.135 10.855 ;
        RECT 57.410 8.685 57.685 10.855 ;
        RECT 57.960 8.685 58.235 10.855 ;
        RECT 58.510 8.685 58.785 10.855 ;
        RECT 59.060 8.685 59.335 10.855 ;
        RECT 59.610 8.685 59.885 10.855 ;
        RECT 60.160 8.685 60.435 10.855 ;
        RECT 60.710 8.685 60.985 10.855 ;
        RECT 61.260 8.685 61.605 10.855 ;
        RECT 69.000 8.805 69.170 10.855 ;
        RECT 69.000 8.775 69.455 8.805 ;
        RECT 52.415 8.600 52.870 8.605 ;
        RECT 52.580 8.575 52.870 8.600 ;
        RECT 54.550 8.325 61.605 8.685 ;
        RECT 68.990 8.605 69.455 8.775 ;
        RECT 71.270 8.685 71.520 10.855 ;
        RECT 71.795 8.685 72.070 10.855 ;
        RECT 72.345 8.685 72.620 10.855 ;
        RECT 72.895 8.685 73.170 10.855 ;
        RECT 73.445 8.685 73.720 10.855 ;
        RECT 73.995 8.685 74.270 10.855 ;
        RECT 74.545 8.685 74.820 10.855 ;
        RECT 75.095 8.685 75.370 10.855 ;
        RECT 75.645 8.685 75.920 10.855 ;
        RECT 76.195 8.685 76.470 10.855 ;
        RECT 76.745 8.685 77.020 10.855 ;
        RECT 77.295 8.685 77.570 10.855 ;
        RECT 77.845 8.685 78.190 10.855 ;
        RECT 85.580 8.805 85.750 10.855 ;
        RECT 85.580 8.775 86.035 8.805 ;
        RECT 69.000 8.600 69.455 8.605 ;
        RECT 69.165 8.575 69.455 8.600 ;
        RECT 71.135 8.325 78.190 8.685 ;
        RECT 85.570 8.605 86.035 8.775 ;
        RECT 87.850 8.685 88.100 10.855 ;
        RECT 88.375 8.685 88.650 10.855 ;
        RECT 88.925 8.685 89.200 10.855 ;
        RECT 89.475 8.685 89.750 10.855 ;
        RECT 90.025 8.685 90.300 10.855 ;
        RECT 90.575 8.685 90.850 10.855 ;
        RECT 91.125 8.685 91.400 10.855 ;
        RECT 91.675 8.685 91.950 10.855 ;
        RECT 92.225 8.685 92.500 10.855 ;
        RECT 92.775 8.685 93.050 10.855 ;
        RECT 93.325 8.685 93.600 10.855 ;
        RECT 93.875 8.685 94.150 10.855 ;
        RECT 94.425 8.685 94.770 10.855 ;
        RECT 85.580 8.600 86.035 8.605 ;
        RECT 85.745 8.575 86.035 8.600 ;
        RECT 87.715 8.325 94.770 8.685 ;
        RECT 22.980 7.945 23.120 8.325 ;
        RECT 23.910 7.945 24.340 8.045 ;
        RECT 39.565 7.945 39.705 8.325 ;
        RECT 40.495 7.945 40.925 8.045 ;
        RECT 56.150 7.945 56.290 8.325 ;
        RECT 57.080 7.945 57.510 8.045 ;
        RECT 72.735 7.945 72.875 8.325 ;
        RECT 73.665 7.945 74.095 8.045 ;
        RECT 89.315 7.945 89.455 8.325 ;
        RECT 90.245 7.945 90.675 8.045 ;
        RECT 22.980 7.805 25.330 7.945 ;
        RECT 22.980 7.365 23.120 7.805 ;
        RECT 23.920 7.775 24.200 7.805 ;
        RECT 23.940 7.745 24.200 7.775 ;
        RECT 25.190 7.365 25.330 7.805 ;
        RECT 39.565 7.805 41.915 7.945 ;
        RECT 39.565 7.365 39.705 7.805 ;
        RECT 40.505 7.775 40.785 7.805 ;
        RECT 40.525 7.745 40.785 7.775 ;
        RECT 41.775 7.365 41.915 7.805 ;
        RECT 56.150 7.805 58.500 7.945 ;
        RECT 56.150 7.365 56.290 7.805 ;
        RECT 57.090 7.775 57.370 7.805 ;
        RECT 57.110 7.745 57.370 7.775 ;
        RECT 58.360 7.365 58.500 7.805 ;
        RECT 72.735 7.805 75.085 7.945 ;
        RECT 72.735 7.365 72.875 7.805 ;
        RECT 73.675 7.775 73.955 7.805 ;
        RECT 73.695 7.745 73.955 7.775 ;
        RECT 74.945 7.365 75.085 7.805 ;
        RECT 89.315 7.805 91.665 7.945 ;
        RECT 89.315 7.365 89.455 7.805 ;
        RECT 90.255 7.775 90.535 7.805 ;
        RECT 90.275 7.745 90.535 7.775 ;
        RECT 91.525 7.365 91.665 7.805 ;
        RECT 22.900 7.135 23.190 7.365 ;
        RECT 25.110 7.135 25.400 7.365 ;
        RECT 39.485 7.135 39.775 7.365 ;
        RECT 41.695 7.135 41.985 7.365 ;
        RECT 56.070 7.135 56.360 7.365 ;
        RECT 58.280 7.135 58.570 7.365 ;
        RECT 72.655 7.135 72.945 7.365 ;
        RECT 74.865 7.135 75.155 7.365 ;
        RECT 89.235 7.135 89.525 7.365 ;
        RECT 91.445 7.135 91.735 7.365 ;
      LAYER met2 ;
        RECT 23.920 7.715 24.200 8.095 ;
        RECT 40.505 7.715 40.785 8.095 ;
        RECT 57.090 7.715 57.370 8.095 ;
        RECT 73.675 7.715 73.955 8.095 ;
        RECT 90.255 7.715 90.535 8.095 ;
      LAYER met3 ;
        RECT 23.860 8.095 24.200 8.195 ;
        RECT 40.445 8.095 40.785 8.195 ;
        RECT 57.030 8.095 57.370 8.195 ;
        RECT 73.615 8.095 73.955 8.195 ;
        RECT 90.195 8.095 90.535 8.195 ;
        RECT 23.860 8.085 24.220 8.095 ;
        RECT 40.445 8.085 40.805 8.095 ;
        RECT 57.030 8.085 57.390 8.095 ;
        RECT 73.615 8.085 73.975 8.095 ;
        RECT 90.195 8.085 90.555 8.095 ;
        RECT 23.420 8.065 24.220 8.085 ;
        RECT 40.005 8.065 40.805 8.085 ;
        RECT 56.590 8.065 57.390 8.085 ;
        RECT 73.175 8.065 73.975 8.085 ;
        RECT 89.755 8.065 90.555 8.085 ;
        RECT 23.420 7.785 24.225 8.065 ;
        RECT 40.005 7.785 40.810 8.065 ;
        RECT 56.590 7.785 57.395 8.065 ;
        RECT 73.175 7.785 73.980 8.065 ;
        RECT 89.755 7.785 90.560 8.065 ;
        RECT 23.880 7.755 24.225 7.785 ;
        RECT 40.465 7.755 40.810 7.785 ;
        RECT 57.050 7.755 57.395 7.785 ;
        RECT 73.635 7.755 73.980 7.785 ;
        RECT 90.215 7.755 90.560 7.785 ;
        RECT 23.890 7.725 24.225 7.755 ;
        RECT 40.475 7.725 40.810 7.755 ;
        RECT 57.060 7.725 57.395 7.755 ;
        RECT 73.645 7.725 73.980 7.755 ;
        RECT 90.225 7.725 90.560 7.755 ;
    END
    PORT
      LAYER li1 ;
        RECT 21.300 3.355 21.555 3.905 ;
        RECT 21.300 3.095 21.560 3.355 ;
        RECT 23.890 3.095 24.220 3.545 ;
        RECT 26.270 3.095 26.520 3.625 ;
        RECT 27.140 3.095 27.380 3.895 ;
        RECT 28.050 3.095 28.320 3.895 ;
        RECT 37.885 3.355 38.140 3.905 ;
        RECT 37.885 3.095 38.145 3.355 ;
        RECT 40.475 3.095 40.805 3.545 ;
        RECT 42.855 3.095 43.105 3.625 ;
        RECT 43.725 3.095 43.965 3.895 ;
        RECT 44.635 3.095 44.905 3.895 ;
        RECT 54.470 3.355 54.725 3.905 ;
        RECT 54.470 3.095 54.730 3.355 ;
        RECT 57.060 3.095 57.390 3.545 ;
        RECT 59.440 3.095 59.690 3.625 ;
        RECT 60.310 3.095 60.550 3.895 ;
        RECT 61.220 3.095 61.490 3.895 ;
        RECT 71.055 3.355 71.310 3.905 ;
        RECT 71.055 3.095 71.315 3.355 ;
        RECT 73.645 3.095 73.975 3.545 ;
        RECT 76.025 3.095 76.275 3.625 ;
        RECT 76.895 3.095 77.135 3.895 ;
        RECT 77.805 3.095 78.075 3.895 ;
        RECT 87.635 3.355 87.890 3.905 ;
        RECT 87.635 3.095 87.895 3.355 ;
        RECT 90.225 3.095 90.555 3.545 ;
        RECT 92.605 3.095 92.855 3.625 ;
        RECT 93.475 3.095 93.715 3.895 ;
        RECT 94.385 3.095 94.655 3.895 ;
        RECT 21.220 2.925 28.610 3.095 ;
        RECT 37.805 2.925 45.195 3.095 ;
        RECT 54.390 2.925 61.780 3.095 ;
        RECT 70.975 2.925 78.365 3.095 ;
        RECT 87.555 2.925 94.945 3.095 ;
        RECT 21.265 1.600 21.525 2.925 ;
        RECT 21.815 1.600 22.075 2.925 ;
        RECT 22.355 1.600 22.615 2.925 ;
        RECT 22.895 1.600 23.135 2.925 ;
        RECT 23.435 1.600 23.675 2.925 ;
        RECT 23.955 1.600 24.195 2.925 ;
        RECT 24.475 1.600 24.715 2.925 ;
        RECT 24.995 1.600 25.235 2.925 ;
        RECT 25.515 1.600 25.755 2.925 ;
        RECT 25.995 1.600 26.235 2.925 ;
        RECT 26.475 1.600 26.715 2.925 ;
        RECT 26.955 1.600 27.195 2.925 ;
        RECT 27.435 1.600 27.675 2.925 ;
        RECT 27.915 1.600 28.155 2.925 ;
        RECT 28.395 1.600 28.610 2.925 ;
        RECT 29.680 1.600 29.850 2.230 ;
        RECT 32.425 1.600 32.595 2.230 ;
        RECT 33.415 1.600 33.585 2.230 ;
        RECT 37.850 1.600 38.110 2.925 ;
        RECT 38.400 1.600 38.660 2.925 ;
        RECT 38.940 1.600 39.200 2.925 ;
        RECT 39.480 1.600 39.720 2.925 ;
        RECT 40.020 1.600 40.260 2.925 ;
        RECT 40.540 1.600 40.780 2.925 ;
        RECT 41.060 1.600 41.300 2.925 ;
        RECT 41.580 1.600 41.820 2.925 ;
        RECT 42.100 1.600 42.340 2.925 ;
        RECT 42.580 1.600 42.820 2.925 ;
        RECT 43.060 1.600 43.300 2.925 ;
        RECT 43.540 1.600 43.780 2.925 ;
        RECT 44.020 1.600 44.260 2.925 ;
        RECT 44.500 1.600 44.740 2.925 ;
        RECT 44.980 1.600 45.195 2.925 ;
        RECT 46.265 1.600 46.435 2.230 ;
        RECT 49.010 1.600 49.180 2.230 ;
        RECT 50.000 1.600 50.170 2.230 ;
        RECT 54.435 1.600 54.695 2.925 ;
        RECT 54.985 1.600 55.245 2.925 ;
        RECT 55.525 1.600 55.785 2.925 ;
        RECT 56.065 1.600 56.305 2.925 ;
        RECT 56.605 1.600 56.845 2.925 ;
        RECT 57.125 1.600 57.365 2.925 ;
        RECT 57.645 1.600 57.885 2.925 ;
        RECT 58.165 1.600 58.405 2.925 ;
        RECT 58.685 1.600 58.925 2.925 ;
        RECT 59.165 1.600 59.405 2.925 ;
        RECT 59.645 1.600 59.885 2.925 ;
        RECT 60.125 1.600 60.365 2.925 ;
        RECT 60.605 1.600 60.845 2.925 ;
        RECT 61.085 1.600 61.325 2.925 ;
        RECT 61.565 1.600 61.780 2.925 ;
        RECT 62.850 1.600 63.020 2.230 ;
        RECT 65.595 1.600 65.765 2.230 ;
        RECT 66.585 1.600 66.755 2.230 ;
        RECT 71.020 1.600 71.280 2.925 ;
        RECT 71.570 1.600 71.830 2.925 ;
        RECT 72.110 1.600 72.370 2.925 ;
        RECT 72.650 1.600 72.890 2.925 ;
        RECT 73.190 1.600 73.430 2.925 ;
        RECT 73.710 1.600 73.950 2.925 ;
        RECT 74.230 1.600 74.470 2.925 ;
        RECT 74.750 1.600 74.990 2.925 ;
        RECT 75.270 1.600 75.510 2.925 ;
        RECT 75.750 1.600 75.990 2.925 ;
        RECT 76.230 1.600 76.470 2.925 ;
        RECT 76.710 1.600 76.950 2.925 ;
        RECT 77.190 1.600 77.430 2.925 ;
        RECT 77.670 1.600 77.910 2.925 ;
        RECT 78.150 1.600 78.365 2.925 ;
        RECT 79.435 1.600 79.605 2.230 ;
        RECT 82.180 1.600 82.350 2.230 ;
        RECT 83.170 1.600 83.340 2.230 ;
        RECT 87.600 1.600 87.860 2.925 ;
        RECT 88.150 1.600 88.410 2.925 ;
        RECT 88.690 1.600 88.950 2.925 ;
        RECT 89.230 1.600 89.470 2.925 ;
        RECT 89.770 1.600 90.010 2.925 ;
        RECT 90.290 1.600 90.530 2.925 ;
        RECT 90.810 1.600 91.050 2.925 ;
        RECT 91.330 1.600 91.570 2.925 ;
        RECT 91.850 1.600 92.090 2.925 ;
        RECT 92.330 1.600 92.570 2.925 ;
        RECT 92.810 1.600 93.050 2.925 ;
        RECT 93.290 1.600 93.530 2.925 ;
        RECT 93.770 1.600 94.010 2.925 ;
        RECT 94.250 1.600 94.490 2.925 ;
        RECT 94.730 1.600 94.945 2.925 ;
        RECT 96.015 1.600 96.185 2.230 ;
        RECT 98.760 1.600 98.930 2.230 ;
        RECT 99.750 1.600 99.920 2.230 ;
        RECT 0.000 0.000 100.725 1.600 ;
      LAYER met1 ;
        RECT 21.220 2.765 28.610 3.125 ;
        RECT 37.805 2.765 45.195 3.125 ;
        RECT 54.390 2.765 61.780 3.125 ;
        RECT 70.975 2.765 78.365 3.125 ;
        RECT 87.555 2.765 94.945 3.125 ;
        RECT 21.265 1.600 21.525 2.765 ;
        RECT 21.815 1.600 22.075 2.765 ;
        RECT 22.355 1.600 22.615 2.765 ;
        RECT 22.895 1.600 23.135 2.765 ;
        RECT 23.435 1.600 23.675 2.765 ;
        RECT 23.955 1.600 24.195 2.765 ;
        RECT 24.475 1.600 24.715 2.765 ;
        RECT 24.995 1.600 25.235 2.765 ;
        RECT 25.515 1.600 25.755 2.765 ;
        RECT 25.995 1.600 26.235 2.765 ;
        RECT 26.475 1.600 26.715 2.765 ;
        RECT 26.955 1.600 27.195 2.765 ;
        RECT 27.435 1.600 27.675 2.765 ;
        RECT 27.915 1.600 28.155 2.765 ;
        RECT 28.395 1.600 28.610 2.765 ;
        RECT 37.850 1.600 38.110 2.765 ;
        RECT 38.400 1.600 38.660 2.765 ;
        RECT 38.940 1.600 39.200 2.765 ;
        RECT 39.480 1.600 39.720 2.765 ;
        RECT 40.020 1.600 40.260 2.765 ;
        RECT 40.540 1.600 40.780 2.765 ;
        RECT 41.060 1.600 41.300 2.765 ;
        RECT 41.580 1.600 41.820 2.765 ;
        RECT 42.100 1.600 42.340 2.765 ;
        RECT 42.580 1.600 42.820 2.765 ;
        RECT 43.060 1.600 43.300 2.765 ;
        RECT 43.540 1.600 43.780 2.765 ;
        RECT 44.020 1.600 44.260 2.765 ;
        RECT 44.500 1.600 44.740 2.765 ;
        RECT 44.980 1.600 45.195 2.765 ;
        RECT 54.435 1.600 54.695 2.765 ;
        RECT 54.985 1.600 55.245 2.765 ;
        RECT 55.525 1.600 55.785 2.765 ;
        RECT 56.065 1.600 56.305 2.765 ;
        RECT 56.605 1.600 56.845 2.765 ;
        RECT 57.125 1.600 57.365 2.765 ;
        RECT 57.645 1.600 57.885 2.765 ;
        RECT 58.165 1.600 58.405 2.765 ;
        RECT 58.685 1.600 58.925 2.765 ;
        RECT 59.165 1.600 59.405 2.765 ;
        RECT 59.645 1.600 59.885 2.765 ;
        RECT 60.125 1.600 60.365 2.765 ;
        RECT 60.605 1.600 60.845 2.765 ;
        RECT 61.085 1.600 61.325 2.765 ;
        RECT 61.565 1.600 61.780 2.765 ;
        RECT 71.020 1.600 71.280 2.765 ;
        RECT 71.570 1.600 71.830 2.765 ;
        RECT 72.110 1.600 72.370 2.765 ;
        RECT 72.650 1.600 72.890 2.765 ;
        RECT 73.190 1.600 73.430 2.765 ;
        RECT 73.710 1.600 73.950 2.765 ;
        RECT 74.230 1.600 74.470 2.765 ;
        RECT 74.750 1.600 74.990 2.765 ;
        RECT 75.270 1.600 75.510 2.765 ;
        RECT 75.750 1.600 75.990 2.765 ;
        RECT 76.230 1.600 76.470 2.765 ;
        RECT 76.710 1.600 76.950 2.765 ;
        RECT 77.190 1.600 77.430 2.765 ;
        RECT 77.670 1.600 77.910 2.765 ;
        RECT 78.150 1.600 78.365 2.765 ;
        RECT 87.600 1.600 87.860 2.765 ;
        RECT 88.150 1.600 88.410 2.765 ;
        RECT 88.690 1.600 88.950 2.765 ;
        RECT 89.230 1.600 89.470 2.765 ;
        RECT 89.770 1.600 90.010 2.765 ;
        RECT 90.290 1.600 90.530 2.765 ;
        RECT 90.810 1.600 91.050 2.765 ;
        RECT 91.330 1.600 91.570 2.765 ;
        RECT 91.850 1.600 92.090 2.765 ;
        RECT 92.330 1.600 92.570 2.765 ;
        RECT 92.810 1.600 93.050 2.765 ;
        RECT 93.290 1.600 93.530 2.765 ;
        RECT 93.770 1.600 94.010 2.765 ;
        RECT 94.250 1.600 94.490 2.765 ;
        RECT 94.730 1.600 94.945 2.765 ;
        RECT 0.000 0.000 100.725 1.600 ;
    END
  END vssd1
  OBS
      LAYER pwell ;
        RECT 21.320 8.335 22.050 8.745 ;
        RECT 23.960 8.495 24.130 8.525 ;
        RECT 27.180 8.495 27.350 8.525 ;
        RECT 23.960 8.335 24.540 8.495 ;
        RECT 27.180 8.385 27.810 8.495 ;
        RECT 27.180 8.335 27.490 8.385 ;
        RECT 21.320 8.145 27.490 8.335 ;
        RECT 37.905 8.335 38.635 8.745 ;
        RECT 40.545 8.495 40.715 8.525 ;
        RECT 43.765 8.495 43.935 8.525 ;
        RECT 40.545 8.335 41.125 8.495 ;
        RECT 43.765 8.385 44.395 8.495 ;
        RECT 43.765 8.335 44.075 8.385 ;
        RECT 37.905 8.145 44.075 8.335 ;
        RECT 54.490 8.335 55.220 8.745 ;
        RECT 57.130 8.495 57.300 8.525 ;
        RECT 60.350 8.495 60.520 8.525 ;
        RECT 57.130 8.335 57.710 8.495 ;
        RECT 60.350 8.385 60.980 8.495 ;
        RECT 60.350 8.335 60.660 8.385 ;
        RECT 54.490 8.145 60.660 8.335 ;
        RECT 71.075 8.335 71.805 8.745 ;
        RECT 73.715 8.495 73.885 8.525 ;
        RECT 76.935 8.495 77.105 8.525 ;
        RECT 73.715 8.335 74.295 8.495 ;
        RECT 76.935 8.385 77.565 8.495 ;
        RECT 76.935 8.335 77.245 8.385 ;
        RECT 71.075 8.145 77.245 8.335 ;
        RECT 87.655 8.335 88.385 8.745 ;
        RECT 90.295 8.495 90.465 8.525 ;
        RECT 93.515 8.495 93.685 8.525 ;
        RECT 90.295 8.335 90.875 8.495 ;
        RECT 93.515 8.385 94.145 8.495 ;
        RECT 93.515 8.335 93.825 8.385 ;
        RECT 87.655 8.145 93.825 8.335 ;
        RECT 22.180 7.515 27.490 8.145 ;
        RECT 22.180 7.425 23.130 7.515 ;
        RECT 24.740 7.425 27.490 7.515 ;
        RECT 38.765 7.515 44.075 8.145 ;
        RECT 38.765 7.425 39.715 7.515 ;
        RECT 41.325 7.425 44.075 7.515 ;
        RECT 55.350 7.515 60.660 8.145 ;
        RECT 55.350 7.425 56.300 7.515 ;
        RECT 57.910 7.425 60.660 7.515 ;
        RECT 71.935 7.515 77.245 8.145 ;
        RECT 71.935 7.425 72.885 7.515 ;
        RECT 74.495 7.425 77.245 7.515 ;
        RECT 88.515 7.515 93.825 8.145 ;
        RECT 88.515 7.425 89.465 7.515 ;
        RECT 91.075 7.425 93.825 7.515 ;
        RECT 21.220 3.815 22.450 4.015 ;
        RECT 23.780 3.815 24.730 4.015 ;
        RECT 21.220 3.790 24.730 3.815 ;
        RECT 26.110 3.790 28.390 4.015 ;
        RECT 21.220 3.305 28.390 3.790 ;
        RECT 37.805 3.815 39.035 4.015 ;
        RECT 40.365 3.815 41.315 4.015 ;
        RECT 37.805 3.790 41.315 3.815 ;
        RECT 42.695 3.790 44.975 4.015 ;
        RECT 37.805 3.305 44.975 3.790 ;
        RECT 54.390 3.815 55.620 4.015 ;
        RECT 56.950 3.815 57.900 4.015 ;
        RECT 54.390 3.790 57.900 3.815 ;
        RECT 59.280 3.790 61.560 4.015 ;
        RECT 54.390 3.305 61.560 3.790 ;
        RECT 70.975 3.815 72.205 4.015 ;
        RECT 73.535 3.815 74.485 4.015 ;
        RECT 70.975 3.790 74.485 3.815 ;
        RECT 75.865 3.790 78.145 4.015 ;
        RECT 70.975 3.305 78.145 3.790 ;
        RECT 87.555 3.815 88.785 4.015 ;
        RECT 90.115 3.815 91.065 4.015 ;
        RECT 87.555 3.790 91.065 3.815 ;
        RECT 92.445 3.790 94.725 4.015 ;
        RECT 87.555 3.305 94.725 3.790 ;
        RECT 21.160 3.135 28.390 3.305 ;
        RECT 21.160 2.705 21.750 3.135 ;
        RECT 23.800 3.110 28.390 3.135 ;
        RECT 37.745 3.135 44.975 3.305 ;
        RECT 24.880 2.925 25.050 3.105 ;
        RECT 27.190 3.095 27.360 3.105 ;
        RECT 27.180 3.085 27.360 3.095 ;
        RECT 27.190 2.925 27.360 3.085 ;
        RECT 37.745 2.705 38.335 3.135 ;
        RECT 40.385 3.110 44.975 3.135 ;
        RECT 54.330 3.135 61.560 3.305 ;
        RECT 41.465 2.925 41.635 3.105 ;
        RECT 43.775 3.095 43.945 3.105 ;
        RECT 43.765 3.085 43.945 3.095 ;
        RECT 43.775 2.925 43.945 3.085 ;
        RECT 54.330 2.705 54.920 3.135 ;
        RECT 56.970 3.110 61.560 3.135 ;
        RECT 70.915 3.135 78.145 3.305 ;
        RECT 58.050 2.925 58.220 3.105 ;
        RECT 60.360 3.095 60.530 3.105 ;
        RECT 60.350 3.085 60.530 3.095 ;
        RECT 60.360 2.925 60.530 3.085 ;
        RECT 70.915 2.705 71.505 3.135 ;
        RECT 73.555 3.110 78.145 3.135 ;
        RECT 87.495 3.135 94.725 3.305 ;
        RECT 74.635 2.925 74.805 3.105 ;
        RECT 76.945 3.095 77.115 3.105 ;
        RECT 76.935 3.085 77.115 3.095 ;
        RECT 76.945 2.925 77.115 3.085 ;
        RECT 87.495 2.705 88.085 3.135 ;
        RECT 90.135 3.110 94.725 3.135 ;
        RECT 91.215 2.925 91.385 3.105 ;
        RECT 93.525 3.095 93.695 3.105 ;
        RECT 93.515 3.085 93.695 3.095 ;
        RECT 93.525 2.925 93.695 3.085 ;
      LAYER li1 ;
        RECT 15.655 10.095 15.830 10.585 ;
        RECT 16.180 10.305 16.350 10.585 ;
        RECT 16.180 10.135 16.410 10.305 ;
        RECT 15.655 9.925 15.825 10.095 ;
        RECT 15.655 9.595 16.065 9.925 ;
        RECT 15.655 9.085 15.825 9.595 ;
        RECT 15.655 8.755 16.065 9.085 ;
        RECT 15.655 8.555 15.825 8.755 ;
        RECT 15.655 7.295 15.830 8.555 ;
        RECT 16.240 8.525 16.410 10.135 ;
        RECT 16.610 10.075 16.785 10.585 ;
        RECT 18.885 10.095 19.060 10.585 ;
        RECT 18.885 9.925 19.055 10.095 ;
        RECT 19.840 10.075 20.015 10.585 ;
        RECT 20.270 10.035 20.445 10.585 ;
        RECT 30.110 10.100 30.285 10.590 ;
        RECT 30.635 10.310 30.805 10.590 ;
        RECT 30.635 10.140 30.865 10.310 ;
        RECT 18.885 9.595 19.295 9.925 ;
        RECT 16.180 8.355 16.410 8.525 ;
        RECT 16.610 8.555 16.780 9.505 ;
        RECT 18.885 9.085 19.055 9.595 ;
        RECT 18.885 8.755 19.295 9.085 ;
        RECT 18.885 8.555 19.055 8.755 ;
        RECT 19.840 8.555 20.010 9.505 ;
        RECT 16.180 7.295 16.350 8.355 ;
        RECT 16.610 7.295 16.785 8.555 ;
        RECT 18.885 7.295 19.060 8.555 ;
        RECT 19.840 7.295 20.015 8.555 ;
        RECT 20.270 8.435 20.440 10.035 ;
        RECT 30.110 9.930 30.280 10.100 ;
        RECT 30.110 9.600 30.520 9.930 ;
        RECT 30.110 9.090 30.280 9.600 ;
        RECT 30.110 8.760 30.520 9.090 ;
        RECT 30.110 8.560 30.280 8.760 ;
        RECT 20.270 7.295 20.445 8.435 ;
        RECT 22.060 7.895 22.620 8.185 ;
        RECT 23.660 8.055 23.920 8.085 ;
        RECT 22.060 6.525 22.310 7.895 ;
        RECT 23.660 7.725 23.990 8.055 ;
        RECT 25.370 7.935 26.680 8.185 ;
        RECT 25.370 7.785 25.550 7.935 ;
        RECT 22.600 7.535 23.990 7.725 ;
        RECT 24.820 7.615 25.550 7.785 ;
        RECT 22.600 7.445 22.770 7.535 ;
        RECT 22.480 7.115 22.770 7.445 ;
        RECT 23.500 7.115 24.180 7.365 ;
        RECT 22.600 6.865 22.770 7.115 ;
        RECT 22.600 6.695 23.545 6.865 ;
        RECT 23.910 6.755 24.180 7.115 ;
        RECT 24.820 6.945 24.990 7.615 ;
        RECT 25.800 7.365 26.010 7.765 ;
        RECT 25.660 7.165 26.010 7.365 ;
        RECT 26.260 7.365 26.510 7.765 ;
        RECT 26.260 7.165 26.730 7.365 ;
        RECT 26.920 7.165 27.370 7.675 ;
        RECT 30.110 7.300 30.285 8.560 ;
        RECT 30.695 8.530 30.865 10.140 ;
        RECT 31.065 10.080 31.240 10.590 ;
        RECT 31.495 10.040 31.670 10.590 ;
        RECT 32.860 10.080 33.030 10.590 ;
        RECT 33.850 10.080 34.020 10.590 ;
        RECT 35.470 10.095 35.645 10.585 ;
        RECT 30.635 8.360 30.865 8.530 ;
        RECT 31.065 8.560 31.235 9.510 ;
        RECT 30.635 7.300 30.805 8.360 ;
        RECT 31.065 7.300 31.240 8.560 ;
        RECT 31.495 8.440 31.665 10.040 ;
        RECT 35.470 9.925 35.640 10.095 ;
        RECT 36.425 10.075 36.600 10.585 ;
        RECT 36.855 10.035 37.030 10.585 ;
        RECT 46.695 10.100 46.870 10.590 ;
        RECT 47.220 10.310 47.390 10.590 ;
        RECT 47.220 10.140 47.450 10.310 ;
        RECT 35.470 9.595 35.880 9.925 ;
        RECT 32.035 9.475 32.265 9.570 ;
        RECT 32.035 9.420 32.655 9.475 ;
        RECT 32.035 9.305 32.955 9.420 ;
        RECT 32.485 9.250 32.955 9.305 ;
        RECT 33.475 9.250 33.945 9.420 ;
        RECT 32.485 8.560 32.655 9.250 ;
        RECT 32.855 8.770 33.025 8.880 ;
        RECT 33.475 8.770 33.645 9.250 ;
        RECT 35.470 9.085 35.640 9.595 ;
        RECT 32.855 8.600 33.645 8.770 ;
        RECT 31.495 7.300 31.670 8.440 ;
        RECT 32.855 7.300 33.030 8.600 ;
        RECT 33.475 8.560 33.645 8.600 ;
        RECT 33.845 8.445 34.015 8.880 ;
        RECT 35.470 8.755 35.880 9.085 ;
        RECT 35.470 8.555 35.640 8.755 ;
        RECT 36.425 8.555 36.595 9.505 ;
        RECT 33.845 7.300 34.020 8.445 ;
        RECT 35.470 7.295 35.645 8.555 ;
        RECT 36.425 7.295 36.600 8.555 ;
        RECT 36.855 8.435 37.025 10.035 ;
        RECT 46.695 9.930 46.865 10.100 ;
        RECT 46.695 9.600 47.105 9.930 ;
        RECT 46.695 9.090 46.865 9.600 ;
        RECT 46.695 8.760 47.105 9.090 ;
        RECT 46.695 8.560 46.865 8.760 ;
        RECT 36.855 7.295 37.030 8.435 ;
        RECT 38.645 7.895 39.205 8.185 ;
        RECT 40.245 8.055 40.505 8.085 ;
        RECT 25.660 6.945 27.400 6.995 ;
        RECT 24.820 6.815 27.400 6.945 ;
        RECT 24.820 6.775 25.880 6.815 ;
        RECT 22.060 5.975 22.520 6.525 ;
        RECT 23.240 5.975 23.545 6.695 ;
        RECT 26.020 6.605 26.900 6.645 ;
        RECT 25.370 6.405 26.900 6.605 ;
        RECT 25.370 6.275 25.540 6.405 ;
        RECT 26.290 6.355 26.900 6.405 ;
        RECT 26.670 6.315 26.900 6.355 ;
        RECT 27.070 6.315 27.400 6.815 ;
        RECT 38.645 6.525 38.895 7.895 ;
        RECT 40.245 7.725 40.575 8.055 ;
        RECT 41.955 7.935 43.265 8.185 ;
        RECT 41.955 7.785 42.135 7.935 ;
        RECT 39.185 7.535 40.575 7.725 ;
        RECT 41.405 7.615 42.135 7.785 ;
        RECT 39.185 7.445 39.355 7.535 ;
        RECT 39.065 7.115 39.355 7.445 ;
        RECT 40.085 7.115 40.765 7.365 ;
        RECT 39.185 6.865 39.355 7.115 ;
        RECT 39.185 6.695 40.130 6.865 ;
        RECT 40.495 6.755 40.765 7.115 ;
        RECT 41.405 6.945 41.575 7.615 ;
        RECT 42.385 7.365 42.595 7.765 ;
        RECT 42.245 7.165 42.595 7.365 ;
        RECT 42.845 7.365 43.095 7.765 ;
        RECT 42.845 7.165 43.315 7.365 ;
        RECT 43.505 7.165 43.955 7.675 ;
        RECT 46.695 7.300 46.870 8.560 ;
        RECT 47.280 8.530 47.450 10.140 ;
        RECT 47.650 10.080 47.825 10.590 ;
        RECT 48.080 10.040 48.255 10.590 ;
        RECT 49.445 10.080 49.615 10.590 ;
        RECT 50.435 10.080 50.605 10.590 ;
        RECT 52.055 10.095 52.230 10.585 ;
        RECT 47.220 8.360 47.450 8.530 ;
        RECT 47.650 8.560 47.820 9.510 ;
        RECT 47.220 7.300 47.390 8.360 ;
        RECT 47.650 7.300 47.825 8.560 ;
        RECT 48.080 8.440 48.250 10.040 ;
        RECT 52.055 9.925 52.225 10.095 ;
        RECT 53.010 10.075 53.185 10.585 ;
        RECT 53.440 10.035 53.615 10.585 ;
        RECT 63.280 10.100 63.455 10.590 ;
        RECT 63.805 10.310 63.975 10.590 ;
        RECT 63.805 10.140 64.035 10.310 ;
        RECT 52.055 9.595 52.465 9.925 ;
        RECT 48.620 9.475 48.850 9.570 ;
        RECT 48.620 9.420 49.240 9.475 ;
        RECT 48.620 9.305 49.540 9.420 ;
        RECT 49.070 9.250 49.540 9.305 ;
        RECT 50.060 9.250 50.530 9.420 ;
        RECT 49.070 8.560 49.240 9.250 ;
        RECT 49.440 8.770 49.610 8.880 ;
        RECT 50.060 8.770 50.230 9.250 ;
        RECT 52.055 9.085 52.225 9.595 ;
        RECT 49.440 8.600 50.230 8.770 ;
        RECT 48.080 7.300 48.255 8.440 ;
        RECT 49.440 7.300 49.615 8.600 ;
        RECT 50.060 8.560 50.230 8.600 ;
        RECT 50.430 8.445 50.600 8.880 ;
        RECT 52.055 8.755 52.465 9.085 ;
        RECT 52.055 8.555 52.225 8.755 ;
        RECT 53.010 8.555 53.180 9.505 ;
        RECT 50.430 7.300 50.605 8.445 ;
        RECT 52.055 7.295 52.230 8.555 ;
        RECT 53.010 7.295 53.185 8.555 ;
        RECT 53.440 8.435 53.610 10.035 ;
        RECT 63.280 9.930 63.450 10.100 ;
        RECT 63.280 9.600 63.690 9.930 ;
        RECT 63.280 9.090 63.450 9.600 ;
        RECT 63.280 8.760 63.690 9.090 ;
        RECT 63.280 8.560 63.450 8.760 ;
        RECT 53.440 7.295 53.615 8.435 ;
        RECT 55.230 7.895 55.790 8.185 ;
        RECT 56.830 8.055 57.090 8.085 ;
        RECT 42.245 6.945 43.985 6.995 ;
        RECT 41.405 6.815 43.985 6.945 ;
        RECT 41.405 6.775 42.465 6.815 ;
        RECT 26.230 6.145 26.560 6.185 ;
        RECT 27.070 6.145 27.890 6.315 ;
        RECT 26.230 5.975 27.400 6.145 ;
        RECT 38.645 5.975 39.105 6.525 ;
        RECT 39.825 5.975 40.130 6.695 ;
        RECT 42.605 6.605 43.485 6.645 ;
        RECT 41.955 6.405 43.485 6.605 ;
        RECT 41.955 6.275 42.125 6.405 ;
        RECT 42.875 6.355 43.485 6.405 ;
        RECT 43.255 6.315 43.485 6.355 ;
        RECT 43.655 6.315 43.985 6.815 ;
        RECT 55.230 6.525 55.480 7.895 ;
        RECT 56.830 7.725 57.160 8.055 ;
        RECT 58.540 7.935 59.850 8.185 ;
        RECT 58.540 7.785 58.720 7.935 ;
        RECT 55.770 7.535 57.160 7.725 ;
        RECT 57.990 7.615 58.720 7.785 ;
        RECT 55.770 7.445 55.940 7.535 ;
        RECT 55.650 7.115 55.940 7.445 ;
        RECT 56.670 7.115 57.350 7.365 ;
        RECT 55.770 6.865 55.940 7.115 ;
        RECT 55.770 6.695 56.715 6.865 ;
        RECT 57.080 6.755 57.350 7.115 ;
        RECT 57.990 6.945 58.160 7.615 ;
        RECT 58.970 7.365 59.180 7.765 ;
        RECT 58.830 7.165 59.180 7.365 ;
        RECT 59.430 7.365 59.680 7.765 ;
        RECT 59.430 7.165 59.900 7.365 ;
        RECT 60.090 7.165 60.540 7.675 ;
        RECT 63.280 7.300 63.455 8.560 ;
        RECT 63.865 8.530 64.035 10.140 ;
        RECT 64.235 10.080 64.410 10.590 ;
        RECT 64.665 10.040 64.840 10.590 ;
        RECT 66.030 10.080 66.200 10.590 ;
        RECT 67.020 10.080 67.190 10.590 ;
        RECT 68.640 10.095 68.815 10.585 ;
        RECT 63.805 8.360 64.035 8.530 ;
        RECT 64.235 8.560 64.405 9.510 ;
        RECT 63.805 7.300 63.975 8.360 ;
        RECT 64.235 7.300 64.410 8.560 ;
        RECT 64.665 8.440 64.835 10.040 ;
        RECT 68.640 9.925 68.810 10.095 ;
        RECT 69.595 10.075 69.770 10.585 ;
        RECT 70.025 10.035 70.200 10.585 ;
        RECT 79.865 10.100 80.040 10.590 ;
        RECT 80.390 10.310 80.560 10.590 ;
        RECT 80.390 10.140 80.620 10.310 ;
        RECT 68.640 9.595 69.050 9.925 ;
        RECT 65.205 9.475 65.435 9.570 ;
        RECT 65.205 9.420 65.825 9.475 ;
        RECT 65.205 9.305 66.125 9.420 ;
        RECT 65.655 9.250 66.125 9.305 ;
        RECT 66.645 9.250 67.115 9.420 ;
        RECT 65.655 8.560 65.825 9.250 ;
        RECT 66.025 8.770 66.195 8.880 ;
        RECT 66.645 8.770 66.815 9.250 ;
        RECT 68.640 9.085 68.810 9.595 ;
        RECT 66.025 8.600 66.815 8.770 ;
        RECT 64.665 7.300 64.840 8.440 ;
        RECT 66.025 7.300 66.200 8.600 ;
        RECT 66.645 8.560 66.815 8.600 ;
        RECT 67.015 8.445 67.185 8.880 ;
        RECT 68.640 8.755 69.050 9.085 ;
        RECT 68.640 8.555 68.810 8.755 ;
        RECT 69.595 8.555 69.765 9.505 ;
        RECT 67.015 7.300 67.190 8.445 ;
        RECT 68.640 7.295 68.815 8.555 ;
        RECT 69.595 7.295 69.770 8.555 ;
        RECT 70.025 8.435 70.195 10.035 ;
        RECT 79.865 9.930 80.035 10.100 ;
        RECT 79.865 9.600 80.275 9.930 ;
        RECT 79.865 9.090 80.035 9.600 ;
        RECT 79.865 8.760 80.275 9.090 ;
        RECT 79.865 8.560 80.035 8.760 ;
        RECT 70.025 7.295 70.200 8.435 ;
        RECT 71.815 7.895 72.375 8.185 ;
        RECT 73.415 8.055 73.675 8.085 ;
        RECT 58.830 6.945 60.570 6.995 ;
        RECT 57.990 6.815 60.570 6.945 ;
        RECT 57.990 6.775 59.050 6.815 ;
        RECT 42.815 6.145 43.145 6.185 ;
        RECT 43.655 6.145 44.475 6.315 ;
        RECT 42.815 5.975 43.985 6.145 ;
        RECT 55.230 5.975 55.690 6.525 ;
        RECT 56.410 5.975 56.715 6.695 ;
        RECT 59.190 6.605 60.070 6.645 ;
        RECT 58.540 6.405 60.070 6.605 ;
        RECT 58.540 6.275 58.710 6.405 ;
        RECT 59.460 6.355 60.070 6.405 ;
        RECT 59.840 6.315 60.070 6.355 ;
        RECT 60.240 6.315 60.570 6.815 ;
        RECT 71.815 6.525 72.065 7.895 ;
        RECT 73.415 7.725 73.745 8.055 ;
        RECT 75.125 7.935 76.435 8.185 ;
        RECT 75.125 7.785 75.305 7.935 ;
        RECT 72.355 7.535 73.745 7.725 ;
        RECT 74.575 7.615 75.305 7.785 ;
        RECT 72.355 7.445 72.525 7.535 ;
        RECT 72.235 7.115 72.525 7.445 ;
        RECT 73.255 7.115 73.935 7.365 ;
        RECT 72.355 6.865 72.525 7.115 ;
        RECT 72.355 6.695 73.300 6.865 ;
        RECT 73.665 6.755 73.935 7.115 ;
        RECT 74.575 6.945 74.745 7.615 ;
        RECT 75.555 7.365 75.765 7.765 ;
        RECT 75.415 7.165 75.765 7.365 ;
        RECT 76.015 7.365 76.265 7.765 ;
        RECT 76.015 7.165 76.485 7.365 ;
        RECT 76.675 7.165 77.125 7.675 ;
        RECT 79.865 7.300 80.040 8.560 ;
        RECT 80.450 8.530 80.620 10.140 ;
        RECT 80.820 10.080 80.995 10.590 ;
        RECT 81.250 10.040 81.425 10.590 ;
        RECT 82.615 10.080 82.785 10.590 ;
        RECT 83.605 10.080 83.775 10.590 ;
        RECT 85.220 10.095 85.395 10.585 ;
        RECT 80.390 8.360 80.620 8.530 ;
        RECT 80.820 8.560 80.990 9.510 ;
        RECT 80.390 7.300 80.560 8.360 ;
        RECT 80.820 7.300 80.995 8.560 ;
        RECT 81.250 8.440 81.420 10.040 ;
        RECT 85.220 9.925 85.390 10.095 ;
        RECT 86.175 10.075 86.350 10.585 ;
        RECT 86.605 10.035 86.780 10.585 ;
        RECT 96.445 10.100 96.620 10.590 ;
        RECT 96.970 10.310 97.140 10.590 ;
        RECT 96.970 10.140 97.200 10.310 ;
        RECT 85.220 9.595 85.630 9.925 ;
        RECT 81.790 9.475 82.020 9.570 ;
        RECT 81.790 9.420 82.410 9.475 ;
        RECT 81.790 9.305 82.710 9.420 ;
        RECT 82.240 9.250 82.710 9.305 ;
        RECT 83.230 9.250 83.700 9.420 ;
        RECT 82.240 8.560 82.410 9.250 ;
        RECT 82.610 8.770 82.780 8.880 ;
        RECT 83.230 8.770 83.400 9.250 ;
        RECT 85.220 9.085 85.390 9.595 ;
        RECT 82.610 8.600 83.400 8.770 ;
        RECT 81.250 7.300 81.425 8.440 ;
        RECT 82.610 7.300 82.785 8.600 ;
        RECT 83.230 8.560 83.400 8.600 ;
        RECT 83.600 8.445 83.770 8.880 ;
        RECT 85.220 8.755 85.630 9.085 ;
        RECT 85.220 8.555 85.390 8.755 ;
        RECT 86.175 8.555 86.345 9.505 ;
        RECT 83.600 7.300 83.775 8.445 ;
        RECT 85.220 7.295 85.395 8.555 ;
        RECT 86.175 7.295 86.350 8.555 ;
        RECT 86.605 8.435 86.775 10.035 ;
        RECT 96.445 9.930 96.615 10.100 ;
        RECT 96.445 9.600 96.855 9.930 ;
        RECT 96.445 9.090 96.615 9.600 ;
        RECT 96.445 8.760 96.855 9.090 ;
        RECT 96.445 8.560 96.615 8.760 ;
        RECT 86.605 7.295 86.780 8.435 ;
        RECT 88.395 7.895 88.955 8.185 ;
        RECT 89.995 8.055 90.255 8.085 ;
        RECT 75.415 6.945 77.155 6.995 ;
        RECT 74.575 6.815 77.155 6.945 ;
        RECT 74.575 6.775 75.635 6.815 ;
        RECT 59.400 6.145 59.730 6.185 ;
        RECT 60.240 6.145 61.060 6.315 ;
        RECT 59.400 5.975 60.570 6.145 ;
        RECT 71.815 5.975 72.275 6.525 ;
        RECT 72.995 5.975 73.300 6.695 ;
        RECT 75.775 6.605 76.655 6.645 ;
        RECT 75.125 6.405 76.655 6.605 ;
        RECT 75.125 6.275 75.295 6.405 ;
        RECT 76.045 6.355 76.655 6.405 ;
        RECT 76.425 6.315 76.655 6.355 ;
        RECT 76.825 6.315 77.155 6.815 ;
        RECT 88.395 6.525 88.645 7.895 ;
        RECT 89.995 7.725 90.325 8.055 ;
        RECT 91.705 7.935 93.015 8.185 ;
        RECT 91.705 7.785 91.885 7.935 ;
        RECT 88.935 7.535 90.325 7.725 ;
        RECT 91.155 7.615 91.885 7.785 ;
        RECT 88.935 7.445 89.105 7.535 ;
        RECT 88.815 7.115 89.105 7.445 ;
        RECT 89.835 7.115 90.515 7.365 ;
        RECT 88.935 6.865 89.105 7.115 ;
        RECT 88.935 6.695 89.880 6.865 ;
        RECT 90.245 6.755 90.515 7.115 ;
        RECT 91.155 6.945 91.325 7.615 ;
        RECT 92.135 7.365 92.345 7.765 ;
        RECT 91.995 7.165 92.345 7.365 ;
        RECT 92.595 7.365 92.845 7.765 ;
        RECT 92.595 7.165 93.065 7.365 ;
        RECT 93.255 7.165 93.705 7.675 ;
        RECT 96.445 7.300 96.620 8.560 ;
        RECT 97.030 8.530 97.200 10.140 ;
        RECT 97.400 10.080 97.575 10.590 ;
        RECT 97.830 10.040 98.005 10.590 ;
        RECT 99.195 10.080 99.365 10.590 ;
        RECT 100.185 10.080 100.355 10.590 ;
        RECT 96.970 8.360 97.200 8.530 ;
        RECT 97.400 8.560 97.570 9.510 ;
        RECT 96.970 7.300 97.140 8.360 ;
        RECT 97.400 7.300 97.575 8.560 ;
        RECT 97.830 8.440 98.000 10.040 ;
        RECT 98.370 9.475 98.600 9.570 ;
        RECT 98.370 9.420 98.990 9.475 ;
        RECT 98.370 9.305 99.290 9.420 ;
        RECT 98.820 9.250 99.290 9.305 ;
        RECT 99.810 9.250 100.280 9.420 ;
        RECT 98.820 8.560 98.990 9.250 ;
        RECT 99.190 8.770 99.360 8.880 ;
        RECT 99.810 8.770 99.980 9.250 ;
        RECT 99.190 8.600 99.980 8.770 ;
        RECT 97.830 7.300 98.005 8.440 ;
        RECT 99.190 7.300 99.365 8.600 ;
        RECT 99.810 8.560 99.980 8.600 ;
        RECT 100.180 8.445 100.350 8.880 ;
        RECT 100.180 7.300 100.355 8.445 ;
        RECT 91.995 6.945 93.735 6.995 ;
        RECT 91.155 6.815 93.735 6.945 ;
        RECT 91.155 6.775 92.215 6.815 ;
        RECT 75.985 6.145 76.315 6.185 ;
        RECT 76.825 6.145 77.645 6.315 ;
        RECT 75.985 5.975 77.155 6.145 ;
        RECT 88.395 5.975 88.855 6.525 ;
        RECT 89.575 5.975 89.880 6.695 ;
        RECT 92.355 6.605 93.235 6.645 ;
        RECT 91.705 6.405 93.235 6.605 ;
        RECT 91.705 6.275 91.875 6.405 ;
        RECT 92.625 6.355 93.235 6.405 ;
        RECT 93.005 6.315 93.235 6.355 ;
        RECT 93.405 6.315 93.735 6.815 ;
        RECT 92.565 6.145 92.895 6.185 ;
        RECT 93.405 6.145 94.225 6.315 ;
        RECT 92.565 5.975 93.735 6.145 ;
        RECT 21.815 5.125 21.985 5.465 ;
        RECT 23.310 5.125 23.780 5.465 ;
        RECT 21.810 5.065 21.985 5.125 ;
        RECT 21.300 4.075 21.640 4.955 ;
        RECT 21.810 4.245 21.980 5.065 ;
        RECT 22.520 4.595 22.770 4.965 ;
        RECT 23.490 4.595 24.210 4.895 ;
        RECT 24.380 4.765 24.650 5.465 ;
        RECT 25.600 5.125 26.080 5.465 ;
        RECT 22.520 4.425 24.310 4.595 ;
        RECT 21.810 3.995 22.910 4.245 ;
        RECT 21.810 3.905 22.060 3.995 ;
        RECT 21.760 3.485 22.060 3.905 ;
        RECT 23.080 3.575 23.330 4.425 ;
        RECT 22.540 3.305 23.330 3.575 ;
        RECT 23.500 3.725 23.910 4.245 ;
        RECT 24.080 3.995 24.310 4.425 ;
        RECT 24.480 3.735 24.650 4.765 ;
        RECT 24.820 4.365 25.080 4.815 ;
        RECT 25.750 4.635 26.510 4.885 ;
        RECT 26.680 4.765 26.950 5.465 ;
        RECT 25.740 4.605 26.510 4.635 ;
        RECT 25.720 4.595 26.510 4.605 ;
        RECT 25.720 4.575 26.610 4.595 ;
        RECT 25.700 4.565 26.610 4.575 ;
        RECT 25.680 4.555 26.610 4.565 ;
        RECT 25.650 4.545 26.610 4.555 ;
        RECT 25.580 4.515 26.610 4.545 ;
        RECT 25.560 4.485 26.610 4.515 ;
        RECT 25.540 4.455 26.610 4.485 ;
        RECT 25.510 4.425 26.610 4.455 ;
        RECT 25.480 4.395 26.610 4.425 ;
        RECT 25.450 4.385 26.610 4.395 ;
        RECT 25.450 4.375 25.810 4.385 ;
        RECT 25.450 4.365 25.800 4.375 ;
        RECT 24.820 4.355 25.780 4.365 ;
        RECT 24.820 4.345 25.770 4.355 ;
        RECT 24.820 4.325 25.750 4.345 ;
        RECT 24.820 4.315 25.740 4.325 ;
        RECT 24.820 4.195 25.710 4.315 ;
        RECT 23.500 3.305 23.700 3.725 ;
        RECT 24.390 3.265 24.650 3.735 ;
        RECT 24.820 3.635 25.370 4.025 ;
        RECT 25.540 3.465 25.710 4.195 ;
        RECT 24.820 3.295 25.710 3.465 ;
        RECT 25.880 3.795 26.210 4.215 ;
        RECT 26.380 3.995 26.610 4.385 ;
        RECT 26.780 4.275 26.950 4.765 ;
        RECT 27.130 4.665 27.460 5.455 ;
        RECT 27.130 4.495 27.810 4.665 ;
        RECT 27.120 4.275 27.470 4.325 ;
        RECT 26.780 4.105 27.470 4.275 ;
        RECT 25.880 3.305 26.100 3.795 ;
        RECT 26.780 3.735 26.950 4.105 ;
        RECT 27.120 4.075 27.470 4.105 ;
        RECT 27.640 3.895 27.810 4.495 ;
        RECT 27.980 4.075 28.330 4.325 ;
        RECT 30.110 3.900 30.285 5.160 ;
        RECT 30.635 4.100 30.805 5.160 ;
        RECT 30.635 3.930 30.865 4.100 ;
        RECT 26.690 3.265 26.950 3.735 ;
        RECT 27.550 3.265 27.880 3.895 ;
        RECT 30.110 3.700 30.280 3.900 ;
        RECT 30.110 3.370 30.520 3.700 ;
        RECT 30.110 2.860 30.280 3.370 ;
        RECT 30.110 2.530 30.520 2.860 ;
        RECT 30.110 2.360 30.280 2.530 ;
        RECT 30.110 1.870 30.285 2.360 ;
        RECT 30.695 2.320 30.865 3.930 ;
        RECT 31.065 3.900 31.240 5.160 ;
        RECT 31.495 4.020 31.670 5.160 ;
        RECT 31.065 2.950 31.235 3.900 ;
        RECT 31.495 2.420 31.665 4.020 ;
        RECT 32.855 4.015 33.030 5.160 ;
        RECT 38.400 5.125 38.570 5.465 ;
        RECT 39.895 5.125 40.365 5.465 ;
        RECT 38.395 5.065 38.570 5.125 ;
        RECT 37.885 4.075 38.225 4.955 ;
        RECT 38.395 4.245 38.565 5.065 ;
        RECT 39.105 4.595 39.355 4.965 ;
        RECT 40.075 4.595 40.795 4.895 ;
        RECT 40.965 4.765 41.235 5.465 ;
        RECT 42.185 5.125 42.665 5.465 ;
        RECT 39.105 4.425 40.895 4.595 ;
        RECT 32.485 3.210 32.655 3.900 ;
        RECT 32.855 3.750 33.025 4.015 ;
        RECT 38.395 3.995 39.495 4.245 ;
        RECT 38.395 3.905 38.645 3.995 ;
        RECT 33.475 3.750 33.645 3.900 ;
        RECT 32.855 3.580 33.645 3.750 ;
        RECT 33.475 3.210 33.645 3.580 ;
        RECT 38.345 3.485 38.645 3.905 ;
        RECT 39.665 3.575 39.915 4.425 ;
        RECT 39.125 3.305 39.915 3.575 ;
        RECT 40.085 3.725 40.495 4.245 ;
        RECT 40.665 3.995 40.895 4.425 ;
        RECT 41.065 3.735 41.235 4.765 ;
        RECT 41.405 4.365 41.665 4.815 ;
        RECT 42.335 4.635 43.095 4.885 ;
        RECT 43.265 4.765 43.535 5.465 ;
        RECT 42.325 4.605 43.095 4.635 ;
        RECT 42.305 4.595 43.095 4.605 ;
        RECT 42.305 4.575 43.195 4.595 ;
        RECT 42.285 4.565 43.195 4.575 ;
        RECT 42.265 4.555 43.195 4.565 ;
        RECT 42.235 4.545 43.195 4.555 ;
        RECT 42.165 4.515 43.195 4.545 ;
        RECT 42.145 4.485 43.195 4.515 ;
        RECT 42.125 4.455 43.195 4.485 ;
        RECT 42.095 4.425 43.195 4.455 ;
        RECT 42.065 4.395 43.195 4.425 ;
        RECT 42.035 4.385 43.195 4.395 ;
        RECT 42.035 4.375 42.395 4.385 ;
        RECT 42.035 4.365 42.385 4.375 ;
        RECT 41.405 4.355 42.365 4.365 ;
        RECT 41.405 4.345 42.355 4.355 ;
        RECT 41.405 4.325 42.335 4.345 ;
        RECT 41.405 4.315 42.325 4.325 ;
        RECT 41.405 4.195 42.295 4.315 ;
        RECT 40.085 3.305 40.285 3.725 ;
        RECT 40.975 3.265 41.235 3.735 ;
        RECT 41.405 3.635 41.955 4.025 ;
        RECT 42.125 3.465 42.295 4.195 ;
        RECT 41.405 3.295 42.295 3.465 ;
        RECT 42.465 3.795 42.795 4.215 ;
        RECT 42.965 3.995 43.195 4.385 ;
        RECT 43.365 4.275 43.535 4.765 ;
        RECT 43.715 4.665 44.045 5.455 ;
        RECT 43.715 4.495 44.395 4.665 ;
        RECT 43.705 4.275 44.055 4.325 ;
        RECT 43.365 4.105 44.055 4.275 ;
        RECT 42.465 3.305 42.685 3.795 ;
        RECT 43.365 3.735 43.535 4.105 ;
        RECT 43.705 4.075 44.055 4.105 ;
        RECT 44.225 3.895 44.395 4.495 ;
        RECT 44.565 4.075 44.915 4.325 ;
        RECT 46.695 3.900 46.870 5.160 ;
        RECT 47.220 4.100 47.390 5.160 ;
        RECT 47.220 3.930 47.450 4.100 ;
        RECT 43.275 3.265 43.535 3.735 ;
        RECT 44.135 3.265 44.465 3.895 ;
        RECT 46.695 3.700 46.865 3.900 ;
        RECT 46.695 3.370 47.105 3.700 ;
        RECT 32.035 3.040 32.955 3.210 ;
        RECT 33.475 3.040 33.945 3.210 ;
        RECT 32.035 2.890 32.265 3.040 ;
        RECT 46.695 2.860 46.865 3.370 ;
        RECT 46.695 2.530 47.105 2.860 ;
        RECT 30.635 2.150 30.865 2.320 ;
        RECT 30.635 1.870 30.805 2.150 ;
        RECT 31.065 1.870 31.240 2.380 ;
        RECT 31.495 1.870 31.670 2.420 ;
        RECT 32.860 1.870 33.030 2.380 ;
        RECT 46.695 2.360 46.865 2.530 ;
        RECT 46.695 1.870 46.870 2.360 ;
        RECT 47.280 2.320 47.450 3.930 ;
        RECT 47.650 3.900 47.825 5.160 ;
        RECT 48.080 4.020 48.255 5.160 ;
        RECT 47.650 2.950 47.820 3.900 ;
        RECT 48.080 2.420 48.250 4.020 ;
        RECT 49.440 4.015 49.615 5.160 ;
        RECT 54.985 5.125 55.155 5.465 ;
        RECT 56.480 5.125 56.950 5.465 ;
        RECT 54.980 5.065 55.155 5.125 ;
        RECT 54.470 4.075 54.810 4.955 ;
        RECT 54.980 4.245 55.150 5.065 ;
        RECT 55.690 4.595 55.940 4.965 ;
        RECT 56.660 4.595 57.380 4.895 ;
        RECT 57.550 4.765 57.820 5.465 ;
        RECT 58.770 5.125 59.250 5.465 ;
        RECT 55.690 4.425 57.480 4.595 ;
        RECT 49.070 3.210 49.240 3.900 ;
        RECT 49.440 3.750 49.610 4.015 ;
        RECT 54.980 3.995 56.080 4.245 ;
        RECT 54.980 3.905 55.230 3.995 ;
        RECT 50.060 3.750 50.230 3.900 ;
        RECT 49.440 3.580 50.230 3.750 ;
        RECT 50.060 3.210 50.230 3.580 ;
        RECT 54.930 3.485 55.230 3.905 ;
        RECT 56.250 3.575 56.500 4.425 ;
        RECT 55.710 3.305 56.500 3.575 ;
        RECT 56.670 3.725 57.080 4.245 ;
        RECT 57.250 3.995 57.480 4.425 ;
        RECT 57.650 3.735 57.820 4.765 ;
        RECT 57.990 4.365 58.250 4.815 ;
        RECT 58.920 4.635 59.680 4.885 ;
        RECT 59.850 4.765 60.120 5.465 ;
        RECT 58.910 4.605 59.680 4.635 ;
        RECT 58.890 4.595 59.680 4.605 ;
        RECT 58.890 4.575 59.780 4.595 ;
        RECT 58.870 4.565 59.780 4.575 ;
        RECT 58.850 4.555 59.780 4.565 ;
        RECT 58.820 4.545 59.780 4.555 ;
        RECT 58.750 4.515 59.780 4.545 ;
        RECT 58.730 4.485 59.780 4.515 ;
        RECT 58.710 4.455 59.780 4.485 ;
        RECT 58.680 4.425 59.780 4.455 ;
        RECT 58.650 4.395 59.780 4.425 ;
        RECT 58.620 4.385 59.780 4.395 ;
        RECT 58.620 4.375 58.980 4.385 ;
        RECT 58.620 4.365 58.970 4.375 ;
        RECT 57.990 4.355 58.950 4.365 ;
        RECT 57.990 4.345 58.940 4.355 ;
        RECT 57.990 4.325 58.920 4.345 ;
        RECT 57.990 4.315 58.910 4.325 ;
        RECT 57.990 4.195 58.880 4.315 ;
        RECT 56.670 3.305 56.870 3.725 ;
        RECT 57.560 3.265 57.820 3.735 ;
        RECT 57.990 3.635 58.540 4.025 ;
        RECT 58.710 3.465 58.880 4.195 ;
        RECT 57.990 3.295 58.880 3.465 ;
        RECT 59.050 3.795 59.380 4.215 ;
        RECT 59.550 3.995 59.780 4.385 ;
        RECT 59.950 4.275 60.120 4.765 ;
        RECT 60.300 4.665 60.630 5.455 ;
        RECT 60.300 4.495 60.980 4.665 ;
        RECT 60.290 4.275 60.640 4.325 ;
        RECT 59.950 4.105 60.640 4.275 ;
        RECT 59.050 3.305 59.270 3.795 ;
        RECT 59.950 3.735 60.120 4.105 ;
        RECT 60.290 4.075 60.640 4.105 ;
        RECT 60.810 3.895 60.980 4.495 ;
        RECT 61.150 4.075 61.500 4.325 ;
        RECT 63.280 3.900 63.455 5.160 ;
        RECT 63.805 4.100 63.975 5.160 ;
        RECT 63.805 3.930 64.035 4.100 ;
        RECT 59.860 3.265 60.120 3.735 ;
        RECT 60.720 3.265 61.050 3.895 ;
        RECT 63.280 3.700 63.450 3.900 ;
        RECT 63.280 3.370 63.690 3.700 ;
        RECT 48.620 3.040 49.540 3.210 ;
        RECT 50.060 3.040 50.530 3.210 ;
        RECT 48.620 2.890 48.850 3.040 ;
        RECT 63.280 2.860 63.450 3.370 ;
        RECT 63.280 2.530 63.690 2.860 ;
        RECT 47.220 2.150 47.450 2.320 ;
        RECT 47.220 1.870 47.390 2.150 ;
        RECT 47.650 1.870 47.825 2.380 ;
        RECT 48.080 1.870 48.255 2.420 ;
        RECT 49.445 1.870 49.615 2.380 ;
        RECT 63.280 2.360 63.450 2.530 ;
        RECT 63.280 1.870 63.455 2.360 ;
        RECT 63.865 2.320 64.035 3.930 ;
        RECT 64.235 3.900 64.410 5.160 ;
        RECT 64.665 4.020 64.840 5.160 ;
        RECT 64.235 2.950 64.405 3.900 ;
        RECT 64.665 2.420 64.835 4.020 ;
        RECT 66.025 4.015 66.200 5.160 ;
        RECT 71.570 5.125 71.740 5.465 ;
        RECT 73.065 5.125 73.535 5.465 ;
        RECT 71.565 5.065 71.740 5.125 ;
        RECT 71.055 4.075 71.395 4.955 ;
        RECT 71.565 4.245 71.735 5.065 ;
        RECT 72.275 4.595 72.525 4.965 ;
        RECT 73.245 4.595 73.965 4.895 ;
        RECT 74.135 4.765 74.405 5.465 ;
        RECT 75.355 5.125 75.835 5.465 ;
        RECT 72.275 4.425 74.065 4.595 ;
        RECT 65.655 3.210 65.825 3.900 ;
        RECT 66.025 3.750 66.195 4.015 ;
        RECT 71.565 3.995 72.665 4.245 ;
        RECT 71.565 3.905 71.815 3.995 ;
        RECT 66.645 3.750 66.815 3.900 ;
        RECT 66.025 3.580 66.815 3.750 ;
        RECT 66.645 3.210 66.815 3.580 ;
        RECT 71.515 3.485 71.815 3.905 ;
        RECT 72.835 3.575 73.085 4.425 ;
        RECT 72.295 3.305 73.085 3.575 ;
        RECT 73.255 3.725 73.665 4.245 ;
        RECT 73.835 3.995 74.065 4.425 ;
        RECT 74.235 3.735 74.405 4.765 ;
        RECT 74.575 4.365 74.835 4.815 ;
        RECT 75.505 4.635 76.265 4.885 ;
        RECT 76.435 4.765 76.705 5.465 ;
        RECT 75.495 4.605 76.265 4.635 ;
        RECT 75.475 4.595 76.265 4.605 ;
        RECT 75.475 4.575 76.365 4.595 ;
        RECT 75.455 4.565 76.365 4.575 ;
        RECT 75.435 4.555 76.365 4.565 ;
        RECT 75.405 4.545 76.365 4.555 ;
        RECT 75.335 4.515 76.365 4.545 ;
        RECT 75.315 4.485 76.365 4.515 ;
        RECT 75.295 4.455 76.365 4.485 ;
        RECT 75.265 4.425 76.365 4.455 ;
        RECT 75.235 4.395 76.365 4.425 ;
        RECT 75.205 4.385 76.365 4.395 ;
        RECT 75.205 4.375 75.565 4.385 ;
        RECT 75.205 4.365 75.555 4.375 ;
        RECT 74.575 4.355 75.535 4.365 ;
        RECT 74.575 4.345 75.525 4.355 ;
        RECT 74.575 4.325 75.505 4.345 ;
        RECT 74.575 4.315 75.495 4.325 ;
        RECT 74.575 4.195 75.465 4.315 ;
        RECT 73.255 3.305 73.455 3.725 ;
        RECT 74.145 3.265 74.405 3.735 ;
        RECT 74.575 3.635 75.125 4.025 ;
        RECT 75.295 3.465 75.465 4.195 ;
        RECT 74.575 3.295 75.465 3.465 ;
        RECT 75.635 3.795 75.965 4.215 ;
        RECT 76.135 3.995 76.365 4.385 ;
        RECT 76.535 4.275 76.705 4.765 ;
        RECT 76.885 4.665 77.215 5.455 ;
        RECT 76.885 4.495 77.565 4.665 ;
        RECT 76.875 4.275 77.225 4.325 ;
        RECT 76.535 4.105 77.225 4.275 ;
        RECT 75.635 3.305 75.855 3.795 ;
        RECT 76.535 3.735 76.705 4.105 ;
        RECT 76.875 4.075 77.225 4.105 ;
        RECT 77.395 3.895 77.565 4.495 ;
        RECT 77.735 4.075 78.085 4.325 ;
        RECT 79.865 3.900 80.040 5.160 ;
        RECT 80.390 4.100 80.560 5.160 ;
        RECT 80.390 3.930 80.620 4.100 ;
        RECT 76.445 3.265 76.705 3.735 ;
        RECT 77.305 3.265 77.635 3.895 ;
        RECT 79.865 3.700 80.035 3.900 ;
        RECT 79.865 3.370 80.275 3.700 ;
        RECT 65.205 3.040 66.125 3.210 ;
        RECT 66.645 3.040 67.115 3.210 ;
        RECT 65.205 2.890 65.435 3.040 ;
        RECT 79.865 2.860 80.035 3.370 ;
        RECT 79.865 2.530 80.275 2.860 ;
        RECT 63.805 2.150 64.035 2.320 ;
        RECT 63.805 1.870 63.975 2.150 ;
        RECT 64.235 1.870 64.410 2.380 ;
        RECT 64.665 1.870 64.840 2.420 ;
        RECT 66.030 1.870 66.200 2.380 ;
        RECT 79.865 2.360 80.035 2.530 ;
        RECT 79.865 1.870 80.040 2.360 ;
        RECT 80.450 2.320 80.620 3.930 ;
        RECT 80.820 3.900 80.995 5.160 ;
        RECT 81.250 4.020 81.425 5.160 ;
        RECT 80.820 2.950 80.990 3.900 ;
        RECT 81.250 2.420 81.420 4.020 ;
        RECT 82.610 4.015 82.785 5.160 ;
        RECT 88.150 5.125 88.320 5.465 ;
        RECT 89.645 5.125 90.115 5.465 ;
        RECT 88.145 5.065 88.320 5.125 ;
        RECT 87.635 4.075 87.975 4.955 ;
        RECT 88.145 4.245 88.315 5.065 ;
        RECT 88.855 4.595 89.105 4.965 ;
        RECT 89.825 4.595 90.545 4.895 ;
        RECT 90.715 4.765 90.985 5.465 ;
        RECT 91.935 5.125 92.415 5.465 ;
        RECT 88.855 4.425 90.645 4.595 ;
        RECT 82.240 3.210 82.410 3.900 ;
        RECT 82.610 3.750 82.780 4.015 ;
        RECT 88.145 3.995 89.245 4.245 ;
        RECT 88.145 3.905 88.395 3.995 ;
        RECT 83.230 3.750 83.400 3.900 ;
        RECT 82.610 3.580 83.400 3.750 ;
        RECT 83.230 3.210 83.400 3.580 ;
        RECT 88.095 3.485 88.395 3.905 ;
        RECT 89.415 3.575 89.665 4.425 ;
        RECT 88.875 3.305 89.665 3.575 ;
        RECT 89.835 3.725 90.245 4.245 ;
        RECT 90.415 3.995 90.645 4.425 ;
        RECT 90.815 3.735 90.985 4.765 ;
        RECT 91.155 4.365 91.415 4.815 ;
        RECT 92.085 4.635 92.845 4.885 ;
        RECT 93.015 4.765 93.285 5.465 ;
        RECT 92.075 4.605 92.845 4.635 ;
        RECT 92.055 4.595 92.845 4.605 ;
        RECT 92.055 4.575 92.945 4.595 ;
        RECT 92.035 4.565 92.945 4.575 ;
        RECT 92.015 4.555 92.945 4.565 ;
        RECT 91.985 4.545 92.945 4.555 ;
        RECT 91.915 4.515 92.945 4.545 ;
        RECT 91.895 4.485 92.945 4.515 ;
        RECT 91.875 4.455 92.945 4.485 ;
        RECT 91.845 4.425 92.945 4.455 ;
        RECT 91.815 4.395 92.945 4.425 ;
        RECT 91.785 4.385 92.945 4.395 ;
        RECT 91.785 4.375 92.145 4.385 ;
        RECT 91.785 4.365 92.135 4.375 ;
        RECT 91.155 4.355 92.115 4.365 ;
        RECT 91.155 4.345 92.105 4.355 ;
        RECT 91.155 4.325 92.085 4.345 ;
        RECT 91.155 4.315 92.075 4.325 ;
        RECT 91.155 4.195 92.045 4.315 ;
        RECT 89.835 3.305 90.035 3.725 ;
        RECT 90.725 3.265 90.985 3.735 ;
        RECT 91.155 3.635 91.705 4.025 ;
        RECT 91.875 3.465 92.045 4.195 ;
        RECT 91.155 3.295 92.045 3.465 ;
        RECT 92.215 3.795 92.545 4.215 ;
        RECT 92.715 3.995 92.945 4.385 ;
        RECT 93.115 4.275 93.285 4.765 ;
        RECT 93.465 4.665 93.795 5.455 ;
        RECT 93.465 4.495 94.145 4.665 ;
        RECT 93.455 4.275 93.805 4.325 ;
        RECT 93.115 4.105 93.805 4.275 ;
        RECT 92.215 3.305 92.435 3.795 ;
        RECT 93.115 3.735 93.285 4.105 ;
        RECT 93.455 4.075 93.805 4.105 ;
        RECT 93.975 3.895 94.145 4.495 ;
        RECT 94.315 4.075 94.665 4.325 ;
        RECT 96.445 3.900 96.620 5.160 ;
        RECT 96.970 4.100 97.140 5.160 ;
        RECT 96.970 3.930 97.200 4.100 ;
        RECT 93.025 3.265 93.285 3.735 ;
        RECT 93.885 3.265 94.215 3.895 ;
        RECT 96.445 3.700 96.615 3.900 ;
        RECT 96.445 3.370 96.855 3.700 ;
        RECT 81.790 3.040 82.710 3.210 ;
        RECT 83.230 3.040 83.700 3.210 ;
        RECT 81.790 2.890 82.020 3.040 ;
        RECT 96.445 2.860 96.615 3.370 ;
        RECT 96.445 2.530 96.855 2.860 ;
        RECT 80.390 2.150 80.620 2.320 ;
        RECT 80.390 1.870 80.560 2.150 ;
        RECT 80.820 1.870 80.995 2.380 ;
        RECT 81.250 1.870 81.425 2.420 ;
        RECT 82.615 1.870 82.785 2.380 ;
        RECT 96.445 2.360 96.615 2.530 ;
        RECT 96.445 1.870 96.620 2.360 ;
        RECT 97.030 2.320 97.200 3.930 ;
        RECT 97.400 3.900 97.575 5.160 ;
        RECT 97.830 4.020 98.005 5.160 ;
        RECT 97.400 2.950 97.570 3.900 ;
        RECT 97.830 2.420 98.000 4.020 ;
        RECT 99.190 4.015 99.365 5.160 ;
        RECT 98.820 3.210 98.990 3.900 ;
        RECT 99.190 3.750 99.360 4.015 ;
        RECT 99.810 3.750 99.980 3.900 ;
        RECT 99.190 3.580 99.980 3.750 ;
        RECT 99.810 3.210 99.980 3.580 ;
        RECT 98.370 3.040 99.290 3.210 ;
        RECT 99.810 3.040 100.280 3.210 ;
        RECT 98.370 2.890 98.600 3.040 ;
        RECT 96.970 2.150 97.200 2.320 ;
        RECT 96.970 1.870 97.140 2.150 ;
        RECT 97.400 1.870 97.575 2.380 ;
        RECT 97.830 1.870 98.005 2.420 ;
        RECT 99.195 1.870 99.365 2.380 ;
      LAYER met1 ;
        RECT 16.550 10.045 16.840 10.275 ;
        RECT 19.780 10.045 20.070 10.275 ;
        RECT 31.005 10.050 31.295 10.280 ;
        RECT 16.610 9.585 16.780 10.045 ;
        RECT 19.840 9.675 20.010 10.045 ;
        RECT 16.520 9.305 16.860 9.585 ;
        RECT 19.740 9.305 20.110 9.675 ;
        RECT 31.065 9.575 31.235 10.050 ;
        RECT 32.795 10.020 33.090 10.280 ;
        RECT 33.785 10.020 34.080 10.280 ;
        RECT 36.365 10.045 36.655 10.275 ;
        RECT 47.590 10.050 47.880 10.280 ;
        RECT 31.975 9.575 32.325 9.600 ;
        RECT 31.065 9.540 32.325 9.575 ;
        RECT 31.005 9.405 32.325 9.540 ;
        RECT 31.005 9.310 31.295 9.405 ;
        RECT 31.975 9.310 32.325 9.405 ;
        RECT 20.240 9.165 20.580 9.195 ;
        RECT 31.460 9.170 31.785 9.265 ;
        RECT 20.210 9.135 20.580 9.165 ;
        RECT 31.435 9.140 31.785 9.170 ;
        RECT 20.040 8.965 20.580 9.135 ;
        RECT 31.265 8.970 31.785 9.140 ;
        RECT 20.210 8.935 20.580 8.965 ;
        RECT 31.435 8.940 31.785 8.970 ;
        RECT 20.240 8.915 20.580 8.935 ;
        RECT 32.855 8.920 33.025 10.020 ;
        RECT 33.845 9.270 34.015 10.020 ;
        RECT 36.425 9.675 36.595 10.045 ;
        RECT 36.325 9.305 36.695 9.675 ;
        RECT 47.650 9.575 47.820 10.050 ;
        RECT 49.380 10.020 49.675 10.280 ;
        RECT 50.370 10.020 50.665 10.280 ;
        RECT 52.950 10.045 53.240 10.275 ;
        RECT 64.175 10.050 64.465 10.280 ;
        RECT 48.560 9.575 48.910 9.600 ;
        RECT 47.650 9.540 48.910 9.575 ;
        RECT 47.590 9.405 48.910 9.540 ;
        RECT 47.590 9.310 47.880 9.405 ;
        RECT 48.560 9.310 48.910 9.405 ;
        RECT 33.845 8.945 34.175 9.270 ;
        RECT 36.825 9.165 37.165 9.195 ;
        RECT 48.045 9.170 48.370 9.265 ;
        RECT 36.795 9.135 37.165 9.165 ;
        RECT 48.020 9.140 48.370 9.170 ;
        RECT 36.625 8.965 37.165 9.135 ;
        RECT 47.850 8.970 48.370 9.140 ;
        RECT 33.845 8.920 34.135 8.945 ;
        RECT 36.795 8.935 37.165 8.965 ;
        RECT 48.020 8.940 48.370 8.970 ;
        RECT 32.795 8.915 33.025 8.920 ;
        RECT 16.145 8.775 16.485 8.845 ;
        RECT 30.660 8.810 30.980 8.890 ;
        RECT 30.635 8.780 30.980 8.810 ;
        RECT 16.005 8.605 16.485 8.775 ;
        RECT 30.460 8.610 30.980 8.780 ;
        RECT 32.795 8.680 33.085 8.915 ;
        RECT 33.785 8.795 34.135 8.920 ;
        RECT 36.825 8.915 37.165 8.935 ;
        RECT 49.440 8.920 49.610 10.020 ;
        RECT 50.430 9.270 50.600 10.020 ;
        RECT 53.010 9.675 53.180 10.045 ;
        RECT 52.910 9.305 53.280 9.675 ;
        RECT 64.235 9.575 64.405 10.050 ;
        RECT 65.965 10.020 66.260 10.280 ;
        RECT 66.955 10.020 67.250 10.280 ;
        RECT 69.535 10.045 69.825 10.275 ;
        RECT 80.760 10.050 81.050 10.280 ;
        RECT 65.145 9.575 65.495 9.600 ;
        RECT 64.235 9.540 65.495 9.575 ;
        RECT 64.175 9.405 65.495 9.540 ;
        RECT 64.175 9.310 64.465 9.405 ;
        RECT 65.145 9.310 65.495 9.405 ;
        RECT 50.430 8.945 50.760 9.270 ;
        RECT 53.410 9.165 53.750 9.195 ;
        RECT 64.630 9.170 64.955 9.265 ;
        RECT 53.380 9.135 53.750 9.165 ;
        RECT 64.605 9.140 64.955 9.170 ;
        RECT 53.210 8.965 53.750 9.135 ;
        RECT 64.435 8.970 64.955 9.140 ;
        RECT 50.430 8.920 50.720 8.945 ;
        RECT 53.380 8.935 53.750 8.965 ;
        RECT 64.605 8.940 64.955 8.970 ;
        RECT 49.380 8.915 49.610 8.920 ;
        RECT 47.245 8.810 47.565 8.890 ;
        RECT 33.785 8.680 34.075 8.795 ;
        RECT 47.220 8.780 47.565 8.810 ;
        RECT 47.045 8.610 47.565 8.780 ;
        RECT 49.380 8.680 49.670 8.915 ;
        RECT 50.370 8.805 50.720 8.920 ;
        RECT 53.410 8.915 53.750 8.935 ;
        RECT 66.025 8.920 66.195 10.020 ;
        RECT 67.015 9.270 67.185 10.020 ;
        RECT 69.595 9.675 69.765 10.045 ;
        RECT 69.495 9.305 69.865 9.675 ;
        RECT 80.820 9.575 80.990 10.050 ;
        RECT 82.550 10.020 82.845 10.280 ;
        RECT 83.540 10.020 83.835 10.280 ;
        RECT 86.115 10.045 86.405 10.275 ;
        RECT 97.340 10.050 97.630 10.280 ;
        RECT 81.730 9.575 82.080 9.600 ;
        RECT 80.820 9.540 82.080 9.575 ;
        RECT 80.760 9.405 82.080 9.540 ;
        RECT 80.760 9.310 81.050 9.405 ;
        RECT 81.730 9.310 82.080 9.405 ;
        RECT 67.015 8.945 67.345 9.270 ;
        RECT 69.995 9.165 70.335 9.195 ;
        RECT 81.215 9.170 81.540 9.265 ;
        RECT 69.965 9.135 70.335 9.165 ;
        RECT 81.190 9.140 81.540 9.170 ;
        RECT 69.795 8.965 70.335 9.135 ;
        RECT 81.020 8.970 81.540 9.140 ;
        RECT 67.015 8.920 67.305 8.945 ;
        RECT 69.965 8.935 70.335 8.965 ;
        RECT 81.190 8.940 81.540 8.970 ;
        RECT 65.965 8.915 66.195 8.920 ;
        RECT 63.830 8.810 64.150 8.890 ;
        RECT 50.370 8.680 50.660 8.805 ;
        RECT 63.805 8.780 64.150 8.810 ;
        RECT 63.630 8.610 64.150 8.780 ;
        RECT 65.965 8.680 66.255 8.915 ;
        RECT 66.955 8.805 67.305 8.920 ;
        RECT 69.995 8.915 70.335 8.935 ;
        RECT 82.610 8.920 82.780 10.020 ;
        RECT 83.600 9.270 83.770 10.020 ;
        RECT 86.175 9.675 86.345 10.045 ;
        RECT 86.075 9.305 86.445 9.675 ;
        RECT 97.400 9.575 97.570 10.050 ;
        RECT 99.130 10.020 99.425 10.280 ;
        RECT 100.120 10.020 100.415 10.280 ;
        RECT 98.310 9.575 98.660 9.600 ;
        RECT 97.400 9.540 98.660 9.575 ;
        RECT 97.340 9.405 98.660 9.540 ;
        RECT 97.340 9.310 97.630 9.405 ;
        RECT 98.310 9.310 98.660 9.405 ;
        RECT 83.600 8.945 83.930 9.270 ;
        RECT 86.575 9.165 86.915 9.195 ;
        RECT 97.795 9.170 98.120 9.265 ;
        RECT 86.545 9.135 86.915 9.165 ;
        RECT 97.770 9.140 98.120 9.170 ;
        RECT 86.375 8.965 86.915 9.135 ;
        RECT 97.600 8.970 98.120 9.140 ;
        RECT 83.600 8.920 83.890 8.945 ;
        RECT 86.545 8.935 86.915 8.965 ;
        RECT 97.770 8.940 98.120 8.970 ;
        RECT 82.550 8.915 82.780 8.920 ;
        RECT 80.415 8.810 80.735 8.890 ;
        RECT 66.955 8.680 67.245 8.805 ;
        RECT 80.390 8.780 80.735 8.810 ;
        RECT 80.215 8.610 80.735 8.780 ;
        RECT 82.550 8.680 82.840 8.915 ;
        RECT 83.540 8.805 83.890 8.920 ;
        RECT 86.575 8.915 86.915 8.935 ;
        RECT 99.190 8.920 99.360 10.020 ;
        RECT 100.150 9.985 100.415 10.020 ;
        RECT 100.150 9.585 100.475 9.985 ;
        RECT 100.180 8.920 100.350 9.585 ;
        RECT 99.130 8.915 99.360 8.920 ;
        RECT 100.120 8.915 100.350 8.920 ;
        RECT 96.995 8.810 97.315 8.890 ;
        RECT 83.540 8.680 83.830 8.805 ;
        RECT 96.970 8.780 97.315 8.810 ;
        RECT 96.795 8.610 97.315 8.780 ;
        RECT 99.130 8.680 99.420 8.915 ;
        RECT 100.120 8.680 100.410 8.915 ;
        RECT 16.145 8.565 16.485 8.605 ;
        RECT 30.635 8.580 30.980 8.610 ;
        RECT 47.220 8.580 47.565 8.610 ;
        RECT 63.805 8.580 64.150 8.610 ;
        RECT 80.390 8.580 80.735 8.610 ;
        RECT 96.970 8.580 97.315 8.610 ;
        RECT 30.660 8.565 30.980 8.580 ;
        RECT 47.245 8.565 47.565 8.580 ;
        RECT 63.830 8.565 64.150 8.580 ;
        RECT 80.415 8.565 80.735 8.580 ;
        RECT 96.995 8.565 97.315 8.580 ;
        RECT 23.920 7.325 24.210 7.365 ;
        RECT 24.590 7.325 24.910 7.385 ;
        RECT 23.920 7.185 24.910 7.325 ;
        RECT 23.920 7.135 24.210 7.185 ;
        RECT 24.590 7.125 24.910 7.185 ;
        RECT 25.610 7.125 25.930 7.385 ;
        RECT 26.300 7.135 26.590 7.365 ;
        RECT 26.970 7.325 27.290 7.385 ;
        RECT 40.505 7.325 40.795 7.365 ;
        RECT 41.175 7.325 41.495 7.385 ;
        RECT 26.970 7.185 27.560 7.325 ;
        RECT 40.505 7.185 41.495 7.325 ;
        RECT 24.680 6.985 24.820 7.125 ;
        RECT 26.380 6.985 26.520 7.135 ;
        RECT 26.970 7.125 27.290 7.185 ;
        RECT 40.505 7.135 40.795 7.185 ;
        RECT 41.175 7.125 41.495 7.185 ;
        RECT 42.195 7.125 42.515 7.385 ;
        RECT 42.885 7.135 43.175 7.365 ;
        RECT 43.555 7.325 43.875 7.385 ;
        RECT 57.090 7.325 57.380 7.365 ;
        RECT 57.760 7.325 58.080 7.385 ;
        RECT 43.555 7.185 44.145 7.325 ;
        RECT 57.090 7.185 58.080 7.325 ;
        RECT 24.680 6.845 26.520 6.985 ;
        RECT 41.265 6.985 41.405 7.125 ;
        RECT 42.965 6.985 43.105 7.135 ;
        RECT 43.555 7.125 43.875 7.185 ;
        RECT 57.090 7.135 57.380 7.185 ;
        RECT 57.760 7.125 58.080 7.185 ;
        RECT 58.780 7.125 59.100 7.385 ;
        RECT 59.470 7.135 59.760 7.365 ;
        RECT 60.140 7.325 60.460 7.385 ;
        RECT 73.675 7.325 73.965 7.365 ;
        RECT 74.345 7.325 74.665 7.385 ;
        RECT 60.140 7.185 60.730 7.325 ;
        RECT 73.675 7.185 74.665 7.325 ;
        RECT 41.265 6.845 43.105 6.985 ;
        RECT 57.850 6.985 57.990 7.125 ;
        RECT 59.550 6.985 59.690 7.135 ;
        RECT 60.140 7.125 60.460 7.185 ;
        RECT 73.675 7.135 73.965 7.185 ;
        RECT 74.345 7.125 74.665 7.185 ;
        RECT 75.365 7.125 75.685 7.385 ;
        RECT 76.055 7.135 76.345 7.365 ;
        RECT 76.725 7.325 77.045 7.385 ;
        RECT 90.255 7.325 90.545 7.365 ;
        RECT 90.925 7.325 91.245 7.385 ;
        RECT 76.725 7.185 77.315 7.325 ;
        RECT 90.255 7.185 91.245 7.325 ;
        RECT 57.850 6.845 59.690 6.985 ;
        RECT 74.435 6.985 74.575 7.125 ;
        RECT 76.135 6.985 76.275 7.135 ;
        RECT 76.725 7.125 77.045 7.185 ;
        RECT 90.255 7.135 90.545 7.185 ;
        RECT 90.925 7.125 91.245 7.185 ;
        RECT 91.945 7.125 92.265 7.385 ;
        RECT 92.635 7.135 92.925 7.365 ;
        RECT 93.305 7.325 93.625 7.385 ;
        RECT 93.305 7.185 93.895 7.325 ;
        RECT 74.435 6.845 76.275 6.985 ;
        RECT 91.015 6.985 91.155 7.125 ;
        RECT 92.715 6.985 92.855 7.135 ;
        RECT 93.305 7.125 93.625 7.185 ;
        RECT 91.015 6.845 92.855 6.985 ;
        RECT 22.220 6.305 22.510 6.345 ;
        RECT 24.930 6.305 25.250 6.365 ;
        RECT 22.220 6.165 25.250 6.305 ;
        RECT 22.220 6.115 22.510 6.165 ;
        RECT 24.930 6.105 25.250 6.165 ;
        RECT 27.660 6.105 28.310 6.365 ;
        RECT 38.805 6.305 39.095 6.345 ;
        RECT 41.515 6.305 41.835 6.365 ;
        RECT 38.805 6.165 41.835 6.305 ;
        RECT 38.805 6.115 39.095 6.165 ;
        RECT 41.515 6.105 41.835 6.165 ;
        RECT 44.245 6.105 44.895 6.365 ;
        RECT 55.390 6.305 55.680 6.345 ;
        RECT 58.100 6.305 58.420 6.365 ;
        RECT 55.390 6.165 58.420 6.305 ;
        RECT 55.390 6.115 55.680 6.165 ;
        RECT 58.100 6.105 58.420 6.165 ;
        RECT 60.830 6.105 61.480 6.365 ;
        RECT 71.975 6.305 72.265 6.345 ;
        RECT 74.685 6.305 75.005 6.365 ;
        RECT 71.975 6.165 75.005 6.305 ;
        RECT 71.975 6.115 72.265 6.165 ;
        RECT 74.685 6.105 75.005 6.165 ;
        RECT 77.415 6.105 78.065 6.365 ;
        RECT 88.555 6.305 88.845 6.345 ;
        RECT 91.265 6.305 91.585 6.365 ;
        RECT 88.555 6.165 91.585 6.305 ;
        RECT 88.555 6.115 88.845 6.165 ;
        RECT 91.265 6.105 91.585 6.165 ;
        RECT 93.995 6.105 94.645 6.365 ;
        RECT 23.410 5.285 23.700 5.325 ;
        RECT 25.620 5.285 25.910 5.325 ;
        RECT 26.290 5.285 26.610 5.345 ;
        RECT 23.410 5.145 26.610 5.285 ;
        RECT 23.410 5.095 23.700 5.145 ;
        RECT 25.620 5.095 25.910 5.145 ;
        RECT 26.290 5.085 26.610 5.145 ;
        RECT 39.995 5.285 40.285 5.325 ;
        RECT 42.205 5.285 42.495 5.325 ;
        RECT 42.875 5.285 43.195 5.345 ;
        RECT 39.995 5.145 43.195 5.285 ;
        RECT 39.995 5.095 40.285 5.145 ;
        RECT 42.205 5.095 42.495 5.145 ;
        RECT 42.875 5.085 43.195 5.145 ;
        RECT 56.580 5.285 56.870 5.325 ;
        RECT 58.790 5.285 59.080 5.325 ;
        RECT 59.460 5.285 59.780 5.345 ;
        RECT 56.580 5.145 59.780 5.285 ;
        RECT 56.580 5.095 56.870 5.145 ;
        RECT 58.790 5.095 59.080 5.145 ;
        RECT 59.460 5.085 59.780 5.145 ;
        RECT 73.165 5.285 73.455 5.325 ;
        RECT 75.375 5.285 75.665 5.325 ;
        RECT 76.045 5.285 76.365 5.345 ;
        RECT 73.165 5.145 76.365 5.285 ;
        RECT 73.165 5.095 73.455 5.145 ;
        RECT 75.375 5.095 75.665 5.145 ;
        RECT 76.045 5.085 76.365 5.145 ;
        RECT 89.745 5.285 90.035 5.325 ;
        RECT 91.955 5.285 92.245 5.325 ;
        RECT 92.625 5.285 92.945 5.345 ;
        RECT 89.745 5.145 92.945 5.285 ;
        RECT 89.745 5.095 90.035 5.145 ;
        RECT 91.955 5.095 92.245 5.145 ;
        RECT 92.625 5.085 92.945 5.145 ;
        RECT 25.610 4.605 25.930 4.665 ;
        RECT 27.580 4.605 27.870 4.645 ;
        RECT 28.405 4.620 28.730 4.805 ;
        RECT 28.305 4.605 28.730 4.620 ;
        RECT 25.610 4.480 28.730 4.605 ;
        RECT 42.195 4.605 42.515 4.665 ;
        RECT 44.165 4.605 44.455 4.645 ;
        RECT 44.990 4.620 45.315 4.805 ;
        RECT 44.890 4.605 45.315 4.620 ;
        RECT 42.195 4.480 45.315 4.605 ;
        RECT 58.780 4.605 59.100 4.665 ;
        RECT 60.750 4.605 61.040 4.645 ;
        RECT 61.575 4.620 61.900 4.805 ;
        RECT 61.475 4.605 61.900 4.620 ;
        RECT 58.780 4.480 61.900 4.605 ;
        RECT 75.365 4.605 75.685 4.665 ;
        RECT 77.335 4.605 77.625 4.645 ;
        RECT 78.160 4.620 78.485 4.805 ;
        RECT 78.060 4.605 78.485 4.620 ;
        RECT 75.365 4.480 78.485 4.605 ;
        RECT 91.945 4.605 92.265 4.665 ;
        RECT 93.915 4.605 94.205 4.645 ;
        RECT 94.740 4.620 95.065 4.805 ;
        RECT 94.640 4.605 95.065 4.620 ;
        RECT 91.945 4.480 95.065 4.605 ;
        RECT 25.610 4.465 28.445 4.480 ;
        RECT 42.195 4.465 45.030 4.480 ;
        RECT 58.780 4.465 61.615 4.480 ;
        RECT 75.365 4.465 78.200 4.480 ;
        RECT 91.945 4.465 94.780 4.480 ;
        RECT 25.610 4.405 25.930 4.465 ;
        RECT 27.580 4.415 27.870 4.465 ;
        RECT 42.195 4.405 42.515 4.465 ;
        RECT 44.165 4.415 44.455 4.465 ;
        RECT 58.780 4.405 59.100 4.465 ;
        RECT 60.750 4.415 61.040 4.465 ;
        RECT 75.365 4.405 75.685 4.465 ;
        RECT 77.335 4.415 77.625 4.465 ;
        RECT 91.945 4.405 92.265 4.465 ;
        RECT 93.915 4.415 94.205 4.465 ;
        RECT 21.250 4.265 21.540 4.305 ;
        RECT 23.985 4.265 24.855 4.295 ;
        RECT 26.290 4.265 26.610 4.325 ;
        RECT 27.990 4.265 28.310 4.325 ;
        RECT 21.250 4.155 26.610 4.265 ;
        RECT 21.250 4.125 24.125 4.155 ;
        RECT 24.715 4.125 26.610 4.155 ;
        RECT 27.710 4.125 28.310 4.265 ;
        RECT 21.250 4.075 21.540 4.125 ;
        RECT 26.290 4.065 26.610 4.125 ;
        RECT 27.990 4.065 28.310 4.125 ;
        RECT 37.835 4.265 38.125 4.305 ;
        RECT 40.570 4.265 41.440 4.295 ;
        RECT 42.875 4.265 43.195 4.325 ;
        RECT 44.575 4.265 44.895 4.325 ;
        RECT 37.835 4.155 43.195 4.265 ;
        RECT 37.835 4.125 40.710 4.155 ;
        RECT 41.300 4.125 43.195 4.155 ;
        RECT 44.295 4.125 44.895 4.265 ;
        RECT 37.835 4.075 38.125 4.125 ;
        RECT 42.875 4.065 43.195 4.125 ;
        RECT 44.575 4.065 44.895 4.125 ;
        RECT 54.420 4.265 54.710 4.305 ;
        RECT 57.155 4.265 58.025 4.295 ;
        RECT 59.460 4.265 59.780 4.325 ;
        RECT 61.160 4.265 61.480 4.325 ;
        RECT 54.420 4.155 59.780 4.265 ;
        RECT 54.420 4.125 57.295 4.155 ;
        RECT 57.885 4.125 59.780 4.155 ;
        RECT 60.880 4.125 61.480 4.265 ;
        RECT 54.420 4.075 54.710 4.125 ;
        RECT 59.460 4.065 59.780 4.125 ;
        RECT 61.160 4.065 61.480 4.125 ;
        RECT 71.005 4.265 71.295 4.305 ;
        RECT 73.740 4.265 74.610 4.295 ;
        RECT 76.045 4.265 76.365 4.325 ;
        RECT 77.745 4.265 78.065 4.325 ;
        RECT 71.005 4.155 76.365 4.265 ;
        RECT 71.005 4.125 73.880 4.155 ;
        RECT 74.470 4.125 76.365 4.155 ;
        RECT 77.465 4.125 78.065 4.265 ;
        RECT 71.005 4.075 71.295 4.125 ;
        RECT 76.045 4.065 76.365 4.125 ;
        RECT 77.745 4.065 78.065 4.125 ;
        RECT 87.585 4.265 87.875 4.305 ;
        RECT 90.320 4.265 91.190 4.295 ;
        RECT 92.625 4.265 92.945 4.325 ;
        RECT 94.325 4.265 94.645 4.325 ;
        RECT 87.585 4.155 92.945 4.265 ;
        RECT 87.585 4.125 90.460 4.155 ;
        RECT 91.050 4.125 92.945 4.155 ;
        RECT 94.045 4.125 94.645 4.265 ;
        RECT 87.585 4.075 87.875 4.125 ;
        RECT 92.625 4.065 92.945 4.125 ;
        RECT 94.325 4.065 94.645 4.125 ;
        RECT 24.250 3.965 24.570 3.975 ;
        RECT 23.580 3.735 23.870 3.965 ;
        RECT 24.250 3.925 24.710 3.965 ;
        RECT 24.930 3.925 25.250 3.985 ;
        RECT 26.380 3.925 26.520 4.065 ;
        RECT 24.250 3.785 24.730 3.925 ;
        RECT 24.930 3.785 25.520 3.925 ;
        RECT 26.380 3.785 26.860 3.925 ;
        RECT 30.660 3.880 30.980 3.980 ;
        RECT 40.835 3.965 41.155 3.975 ;
        RECT 30.635 3.860 30.980 3.880 ;
        RECT 24.250 3.735 24.710 3.785 ;
        RECT 23.660 3.535 23.800 3.735 ;
        RECT 24.250 3.715 24.570 3.735 ;
        RECT 24.930 3.725 25.250 3.785 ;
        RECT 25.980 3.665 26.240 3.695 ;
        RECT 25.950 3.645 26.270 3.665 ;
        RECT 26.720 3.645 26.860 3.785 ;
        RECT 30.345 3.690 30.980 3.860 ;
        RECT 30.460 3.680 30.980 3.690 ;
        RECT 30.635 3.660 30.980 3.680 ;
        RECT 30.635 3.650 30.925 3.660 ;
        RECT 25.850 3.535 26.270 3.645 ;
        RECT 23.660 3.405 26.270 3.535 ;
        RECT 26.640 3.415 26.930 3.645 ;
        RECT 28.990 3.490 29.315 3.615 ;
        RECT 31.435 3.490 31.785 3.610 ;
        RECT 32.795 3.545 33.085 3.780 ;
        RECT 40.165 3.735 40.455 3.965 ;
        RECT 40.835 3.925 41.295 3.965 ;
        RECT 41.515 3.925 41.835 3.985 ;
        RECT 42.965 3.925 43.105 4.065 ;
        RECT 40.835 3.785 41.315 3.925 ;
        RECT 41.515 3.785 42.105 3.925 ;
        RECT 42.965 3.785 43.445 3.925 ;
        RECT 47.245 3.880 47.565 3.980 ;
        RECT 57.420 3.965 57.740 3.975 ;
        RECT 47.220 3.860 47.565 3.880 ;
        RECT 40.835 3.735 41.295 3.785 ;
        RECT 32.795 3.540 33.025 3.545 ;
        RECT 23.660 3.395 25.910 3.405 ;
        RECT 28.990 3.320 31.785 3.490 ;
        RECT 28.990 3.290 29.315 3.320 ;
        RECT 31.435 3.260 31.785 3.320 ;
        RECT 31.005 3.120 31.295 3.150 ;
        RECT 31.975 3.120 32.325 3.150 ;
        RECT 31.005 2.950 32.325 3.120 ;
        RECT 31.005 2.920 31.295 2.950 ;
        RECT 31.065 2.410 31.235 2.920 ;
        RECT 31.975 2.860 32.325 2.950 ;
        RECT 32.855 2.440 33.025 3.540 ;
        RECT 40.245 3.535 40.385 3.735 ;
        RECT 40.835 3.715 41.155 3.735 ;
        RECT 41.515 3.725 41.835 3.785 ;
        RECT 42.565 3.665 42.825 3.695 ;
        RECT 42.535 3.645 42.855 3.665 ;
        RECT 43.305 3.645 43.445 3.785 ;
        RECT 46.930 3.690 47.565 3.860 ;
        RECT 47.045 3.680 47.565 3.690 ;
        RECT 47.220 3.660 47.565 3.680 ;
        RECT 47.220 3.650 47.510 3.660 ;
        RECT 42.435 3.535 42.855 3.645 ;
        RECT 40.245 3.405 42.855 3.535 ;
        RECT 43.225 3.415 43.515 3.645 ;
        RECT 45.575 3.490 45.900 3.615 ;
        RECT 48.020 3.490 48.370 3.610 ;
        RECT 49.380 3.545 49.670 3.780 ;
        RECT 56.750 3.735 57.040 3.965 ;
        RECT 57.420 3.925 57.880 3.965 ;
        RECT 58.100 3.925 58.420 3.985 ;
        RECT 59.550 3.925 59.690 4.065 ;
        RECT 57.420 3.785 57.900 3.925 ;
        RECT 58.100 3.785 58.690 3.925 ;
        RECT 59.550 3.785 60.030 3.925 ;
        RECT 63.830 3.880 64.150 3.980 ;
        RECT 74.005 3.965 74.325 3.975 ;
        RECT 63.805 3.860 64.150 3.880 ;
        RECT 57.420 3.735 57.880 3.785 ;
        RECT 49.380 3.540 49.610 3.545 ;
        RECT 40.245 3.395 42.495 3.405 ;
        RECT 45.575 3.320 48.370 3.490 ;
        RECT 45.575 3.290 45.900 3.320 ;
        RECT 48.020 3.260 48.370 3.320 ;
        RECT 47.590 3.120 47.880 3.150 ;
        RECT 48.560 3.120 48.910 3.150 ;
        RECT 47.590 2.950 48.910 3.120 ;
        RECT 47.590 2.920 47.880 2.950 ;
        RECT 31.005 2.180 31.295 2.410 ;
        RECT 32.795 2.180 33.090 2.440 ;
        RECT 47.650 2.410 47.820 2.920 ;
        RECT 48.560 2.860 48.910 2.950 ;
        RECT 49.440 2.440 49.610 3.540 ;
        RECT 56.830 3.535 56.970 3.735 ;
        RECT 57.420 3.715 57.740 3.735 ;
        RECT 58.100 3.725 58.420 3.785 ;
        RECT 59.150 3.665 59.410 3.695 ;
        RECT 59.120 3.645 59.440 3.665 ;
        RECT 59.890 3.645 60.030 3.785 ;
        RECT 63.515 3.690 64.150 3.860 ;
        RECT 63.630 3.680 64.150 3.690 ;
        RECT 63.805 3.660 64.150 3.680 ;
        RECT 63.805 3.650 64.095 3.660 ;
        RECT 59.020 3.535 59.440 3.645 ;
        RECT 56.830 3.405 59.440 3.535 ;
        RECT 59.810 3.415 60.100 3.645 ;
        RECT 62.160 3.490 62.485 3.615 ;
        RECT 64.605 3.490 64.955 3.610 ;
        RECT 65.965 3.545 66.255 3.780 ;
        RECT 73.335 3.735 73.625 3.965 ;
        RECT 74.005 3.925 74.465 3.965 ;
        RECT 74.685 3.925 75.005 3.985 ;
        RECT 76.135 3.925 76.275 4.065 ;
        RECT 74.005 3.785 74.485 3.925 ;
        RECT 74.685 3.785 75.275 3.925 ;
        RECT 76.135 3.785 76.615 3.925 ;
        RECT 80.415 3.880 80.735 3.980 ;
        RECT 90.585 3.965 90.905 3.975 ;
        RECT 80.390 3.860 80.735 3.880 ;
        RECT 74.005 3.735 74.465 3.785 ;
        RECT 65.965 3.540 66.195 3.545 ;
        RECT 56.830 3.395 59.080 3.405 ;
        RECT 62.160 3.320 64.955 3.490 ;
        RECT 62.160 3.290 62.485 3.320 ;
        RECT 64.605 3.260 64.955 3.320 ;
        RECT 64.175 3.120 64.465 3.150 ;
        RECT 65.145 3.120 65.495 3.150 ;
        RECT 64.175 2.950 65.495 3.120 ;
        RECT 64.175 2.920 64.465 2.950 ;
        RECT 47.590 2.180 47.880 2.410 ;
        RECT 49.380 2.180 49.675 2.440 ;
        RECT 64.235 2.410 64.405 2.920 ;
        RECT 65.145 2.860 65.495 2.950 ;
        RECT 66.025 2.440 66.195 3.540 ;
        RECT 73.415 3.535 73.555 3.735 ;
        RECT 74.005 3.715 74.325 3.735 ;
        RECT 74.685 3.725 75.005 3.785 ;
        RECT 75.735 3.665 75.995 3.695 ;
        RECT 75.705 3.645 76.025 3.665 ;
        RECT 76.475 3.645 76.615 3.785 ;
        RECT 80.100 3.690 80.735 3.860 ;
        RECT 80.215 3.680 80.735 3.690 ;
        RECT 80.390 3.660 80.735 3.680 ;
        RECT 80.390 3.650 80.680 3.660 ;
        RECT 75.605 3.535 76.025 3.645 ;
        RECT 73.415 3.405 76.025 3.535 ;
        RECT 76.395 3.415 76.685 3.645 ;
        RECT 78.745 3.490 79.070 3.615 ;
        RECT 81.190 3.490 81.540 3.610 ;
        RECT 82.550 3.545 82.840 3.780 ;
        RECT 89.915 3.735 90.205 3.965 ;
        RECT 90.585 3.925 91.045 3.965 ;
        RECT 91.265 3.925 91.585 3.985 ;
        RECT 92.715 3.925 92.855 4.065 ;
        RECT 90.585 3.785 91.065 3.925 ;
        RECT 91.265 3.785 91.855 3.925 ;
        RECT 92.715 3.785 93.195 3.925 ;
        RECT 96.995 3.880 97.315 3.980 ;
        RECT 96.970 3.860 97.315 3.880 ;
        RECT 90.585 3.735 91.045 3.785 ;
        RECT 82.550 3.540 82.780 3.545 ;
        RECT 73.415 3.395 75.665 3.405 ;
        RECT 78.745 3.320 81.540 3.490 ;
        RECT 78.745 3.290 79.070 3.320 ;
        RECT 81.190 3.260 81.540 3.320 ;
        RECT 80.760 3.120 81.050 3.150 ;
        RECT 81.730 3.120 82.080 3.150 ;
        RECT 80.760 2.950 82.080 3.120 ;
        RECT 80.760 2.920 81.050 2.950 ;
        RECT 64.175 2.180 64.465 2.410 ;
        RECT 65.965 2.180 66.260 2.440 ;
        RECT 80.820 2.410 80.990 2.920 ;
        RECT 81.730 2.860 82.080 2.950 ;
        RECT 82.610 2.440 82.780 3.540 ;
        RECT 89.995 3.535 90.135 3.735 ;
        RECT 90.585 3.715 90.905 3.735 ;
        RECT 91.265 3.725 91.585 3.785 ;
        RECT 92.315 3.665 92.575 3.695 ;
        RECT 92.285 3.645 92.605 3.665 ;
        RECT 93.055 3.645 93.195 3.785 ;
        RECT 96.680 3.690 97.315 3.860 ;
        RECT 96.795 3.680 97.315 3.690 ;
        RECT 96.970 3.660 97.315 3.680 ;
        RECT 96.970 3.650 97.260 3.660 ;
        RECT 92.185 3.535 92.605 3.645 ;
        RECT 89.995 3.405 92.605 3.535 ;
        RECT 92.975 3.415 93.265 3.645 ;
        RECT 95.325 3.490 95.650 3.615 ;
        RECT 97.770 3.490 98.120 3.610 ;
        RECT 99.130 3.545 99.420 3.780 ;
        RECT 99.130 3.540 99.360 3.545 ;
        RECT 89.995 3.395 92.245 3.405 ;
        RECT 95.325 3.320 98.120 3.490 ;
        RECT 95.325 3.290 95.650 3.320 ;
        RECT 97.770 3.260 98.120 3.320 ;
        RECT 97.340 3.120 97.630 3.150 ;
        RECT 98.310 3.120 98.660 3.150 ;
        RECT 97.340 2.950 98.660 3.120 ;
        RECT 97.340 2.920 97.630 2.950 ;
        RECT 80.760 2.180 81.050 2.410 ;
        RECT 82.550 2.180 82.845 2.440 ;
        RECT 97.400 2.410 97.570 2.920 ;
        RECT 98.310 2.860 98.660 2.950 ;
        RECT 99.190 2.440 99.360 3.540 ;
        RECT 97.340 2.180 97.630 2.410 ;
        RECT 99.130 2.180 99.425 2.440 ;
      LAYER met2 ;
        RECT 17.765 10.285 100.355 10.290 ;
        RECT 16.230 10.120 100.355 10.285 ;
        RECT 16.230 10.115 17.765 10.120 ;
        RECT 16.230 8.875 16.400 10.115 ;
        RECT 100.185 9.910 100.355 10.120 ;
        RECT 20.325 9.720 30.505 9.890 ;
        RECT 16.550 9.510 16.830 9.615 ;
        RECT 16.550 9.340 17.715 9.510 ;
        RECT 16.550 9.275 16.830 9.340 ;
        RECT 17.545 9.145 17.715 9.340 ;
        RECT 19.740 9.305 20.110 9.675 ;
        RECT 20.325 9.225 20.495 9.720 ;
        RECT 17.545 9.140 17.865 9.145 ;
        RECT 20.270 9.140 20.550 9.225 ;
        RECT 17.545 8.970 20.550 9.140 ;
        RECT 20.270 8.885 20.550 8.970 ;
        RECT 30.345 9.200 30.505 9.720 ;
        RECT 36.910 9.720 47.090 9.890 ;
        RECT 36.325 9.305 36.695 9.675 ;
        RECT 31.460 9.200 31.785 9.265 ;
        RECT 30.345 9.030 31.785 9.200 ;
        RECT 16.175 8.535 16.455 8.875 ;
        RECT 24.590 7.415 24.870 7.440 ;
        RECT 24.590 7.095 24.880 7.415 ;
        RECT 24.590 7.065 24.870 7.095 ;
        RECT 25.640 7.065 25.920 7.440 ;
        RECT 27.000 7.325 27.260 7.415 ;
        RECT 26.380 7.185 27.260 7.325 ;
        RECT 24.960 6.045 25.240 6.420 ;
        RECT 24.280 3.655 24.560 4.035 ;
        RECT 25.020 4.015 25.160 6.045 ;
        RECT 25.700 5.285 25.840 7.065 ;
        RECT 26.380 5.400 26.520 7.185 ;
        RECT 27.000 7.095 27.260 7.185 ;
        RECT 28.020 6.075 28.280 6.395 ;
        RECT 25.700 5.145 26.180 5.285 ;
        RECT 25.620 4.345 25.900 4.720 ;
        RECT 24.960 3.695 25.220 4.015 ;
        RECT 26.040 3.695 26.180 5.145 ;
        RECT 26.320 5.025 26.600 5.400 ;
        RECT 26.320 4.005 26.600 4.380 ;
        RECT 28.080 4.355 28.220 6.075 ;
        RECT 28.405 4.695 28.730 4.805 ;
        RECT 28.405 4.510 29.235 4.695 ;
        RECT 28.405 4.480 28.730 4.510 ;
        RECT 28.020 4.035 28.280 4.355 ;
        RECT 25.980 3.355 26.240 3.695 ;
        RECT 29.065 3.615 29.235 4.510 ;
        RECT 30.345 3.860 30.505 9.030 ;
        RECT 31.460 8.940 31.785 9.030 ;
        RECT 33.850 9.145 34.175 9.270 ;
        RECT 36.910 9.225 37.080 9.720 ;
        RECT 33.850 9.140 34.685 9.145 ;
        RECT 36.855 9.140 37.135 9.225 ;
        RECT 33.850 8.975 37.135 9.140 ;
        RECT 33.850 8.945 34.175 8.975 ;
        RECT 34.685 8.970 37.135 8.975 ;
        RECT 30.660 8.565 30.980 8.890 ;
        RECT 36.855 8.885 37.135 8.970 ;
        RECT 46.930 9.200 47.090 9.720 ;
        RECT 53.495 9.720 63.675 9.890 ;
        RECT 52.910 9.280 53.280 9.675 ;
        RECT 48.045 9.200 48.370 9.265 ;
        RECT 46.930 9.030 48.370 9.200 ;
        RECT 30.690 8.330 30.860 8.565 ;
        RECT 30.690 8.155 30.865 8.330 ;
        RECT 30.690 7.980 31.665 8.155 ;
        RECT 30.660 3.860 30.980 3.980 ;
        RECT 30.345 3.690 30.980 3.860 ;
        RECT 30.660 3.660 30.980 3.690 ;
        RECT 28.990 3.290 29.315 3.615 ;
        RECT 31.490 3.610 31.665 7.980 ;
        RECT 41.175 7.415 41.455 7.440 ;
        RECT 41.175 7.095 41.465 7.415 ;
        RECT 41.175 7.065 41.455 7.095 ;
        RECT 42.225 7.065 42.505 7.440 ;
        RECT 43.585 7.325 43.845 7.415 ;
        RECT 42.965 7.185 43.845 7.325 ;
        RECT 41.545 6.045 41.825 6.420 ;
        RECT 40.865 3.655 41.145 4.035 ;
        RECT 41.605 4.015 41.745 6.045 ;
        RECT 42.285 5.285 42.425 7.065 ;
        RECT 42.965 5.400 43.105 7.185 ;
        RECT 43.585 7.095 43.845 7.185 ;
        RECT 44.605 6.075 44.865 6.395 ;
        RECT 42.285 5.145 42.765 5.285 ;
        RECT 42.205 4.345 42.485 4.720 ;
        RECT 41.545 3.695 41.805 4.015 ;
        RECT 42.625 3.695 42.765 5.145 ;
        RECT 42.905 5.025 43.185 5.400 ;
        RECT 42.905 4.005 43.185 4.380 ;
        RECT 44.665 4.355 44.805 6.075 ;
        RECT 44.990 4.695 45.315 4.805 ;
        RECT 44.990 4.510 45.820 4.695 ;
        RECT 44.990 4.480 45.315 4.510 ;
        RECT 44.605 4.035 44.865 4.355 ;
        RECT 31.435 3.260 31.785 3.610 ;
        RECT 42.565 3.355 42.825 3.695 ;
        RECT 45.650 3.615 45.820 4.510 ;
        RECT 46.930 3.860 47.090 9.030 ;
        RECT 48.045 8.940 48.370 9.030 ;
        RECT 50.435 9.145 50.760 9.270 ;
        RECT 53.495 9.225 53.665 9.720 ;
        RECT 50.435 9.140 51.050 9.145 ;
        RECT 53.440 9.140 53.720 9.225 ;
        RECT 50.435 8.975 53.720 9.140 ;
        RECT 50.435 8.945 50.760 8.975 ;
        RECT 51.050 8.970 53.720 8.975 ;
        RECT 47.245 8.565 47.565 8.890 ;
        RECT 53.440 8.885 53.720 8.970 ;
        RECT 63.515 9.200 63.675 9.720 ;
        RECT 70.080 9.720 80.260 9.890 ;
        RECT 69.495 9.280 69.865 9.675 ;
        RECT 64.630 9.200 64.955 9.265 ;
        RECT 63.515 9.030 64.955 9.200 ;
        RECT 47.275 8.330 47.445 8.565 ;
        RECT 47.275 8.155 47.450 8.330 ;
        RECT 47.275 7.980 48.250 8.155 ;
        RECT 47.245 3.860 47.565 3.980 ;
        RECT 46.930 3.690 47.565 3.860 ;
        RECT 47.245 3.660 47.565 3.690 ;
        RECT 45.575 3.290 45.900 3.615 ;
        RECT 48.075 3.610 48.250 7.980 ;
        RECT 57.760 7.415 58.040 7.440 ;
        RECT 57.760 7.095 58.050 7.415 ;
        RECT 57.760 7.065 58.040 7.095 ;
        RECT 58.810 7.065 59.090 7.440 ;
        RECT 60.170 7.325 60.430 7.415 ;
        RECT 59.550 7.185 60.430 7.325 ;
        RECT 58.130 6.045 58.410 6.420 ;
        RECT 57.450 3.655 57.730 4.035 ;
        RECT 58.190 4.015 58.330 6.045 ;
        RECT 58.870 5.285 59.010 7.065 ;
        RECT 59.550 5.400 59.690 7.185 ;
        RECT 60.170 7.095 60.430 7.185 ;
        RECT 61.190 6.075 61.450 6.395 ;
        RECT 58.870 5.145 59.350 5.285 ;
        RECT 58.790 4.345 59.070 4.720 ;
        RECT 58.130 3.695 58.390 4.015 ;
        RECT 59.210 3.695 59.350 5.145 ;
        RECT 59.490 5.025 59.770 5.400 ;
        RECT 59.490 4.005 59.770 4.380 ;
        RECT 61.250 4.355 61.390 6.075 ;
        RECT 61.575 4.695 61.900 4.805 ;
        RECT 61.575 4.510 62.405 4.695 ;
        RECT 61.575 4.480 61.900 4.510 ;
        RECT 61.190 4.035 61.450 4.355 ;
        RECT 48.020 3.260 48.370 3.610 ;
        RECT 59.150 3.355 59.410 3.695 ;
        RECT 62.235 3.615 62.405 4.510 ;
        RECT 63.515 3.860 63.675 9.030 ;
        RECT 64.630 8.940 64.955 9.030 ;
        RECT 67.020 9.145 67.345 9.270 ;
        RECT 70.080 9.225 70.250 9.720 ;
        RECT 67.020 9.140 67.865 9.145 ;
        RECT 70.025 9.140 70.305 9.225 ;
        RECT 67.020 8.975 70.305 9.140 ;
        RECT 67.020 8.945 67.345 8.975 ;
        RECT 67.865 8.970 70.305 8.975 ;
        RECT 63.830 8.565 64.150 8.890 ;
        RECT 70.025 8.885 70.305 8.970 ;
        RECT 80.100 9.200 80.260 9.720 ;
        RECT 86.660 9.720 96.840 9.890 ;
        RECT 86.075 9.650 86.445 9.675 ;
        RECT 86.075 9.305 86.450 9.650 ;
        RECT 86.080 9.280 86.450 9.305 ;
        RECT 81.215 9.200 81.540 9.265 ;
        RECT 80.100 9.030 81.540 9.200 ;
        RECT 63.860 8.330 64.030 8.565 ;
        RECT 63.860 8.155 64.035 8.330 ;
        RECT 63.860 7.980 64.835 8.155 ;
        RECT 63.830 3.860 64.150 3.980 ;
        RECT 63.515 3.690 64.150 3.860 ;
        RECT 63.830 3.660 64.150 3.690 ;
        RECT 62.160 3.290 62.485 3.615 ;
        RECT 64.660 3.610 64.835 7.980 ;
        RECT 74.345 7.415 74.625 7.440 ;
        RECT 74.345 7.095 74.635 7.415 ;
        RECT 74.345 7.065 74.625 7.095 ;
        RECT 75.395 7.065 75.675 7.440 ;
        RECT 76.755 7.325 77.015 7.415 ;
        RECT 76.135 7.185 77.015 7.325 ;
        RECT 74.715 6.045 74.995 6.420 ;
        RECT 74.035 3.655 74.315 4.035 ;
        RECT 74.775 4.015 74.915 6.045 ;
        RECT 75.455 5.285 75.595 7.065 ;
        RECT 76.135 5.400 76.275 7.185 ;
        RECT 76.755 7.095 77.015 7.185 ;
        RECT 77.775 6.075 78.035 6.395 ;
        RECT 75.455 5.145 75.935 5.285 ;
        RECT 75.375 4.345 75.655 4.720 ;
        RECT 74.715 3.695 74.975 4.015 ;
        RECT 75.795 3.695 75.935 5.145 ;
        RECT 76.075 5.025 76.355 5.400 ;
        RECT 76.075 4.005 76.355 4.380 ;
        RECT 77.835 4.355 77.975 6.075 ;
        RECT 78.160 4.695 78.485 4.805 ;
        RECT 78.160 4.510 78.990 4.695 ;
        RECT 78.160 4.480 78.485 4.510 ;
        RECT 77.775 4.035 78.035 4.355 ;
        RECT 64.605 3.260 64.955 3.610 ;
        RECT 75.735 3.355 75.995 3.695 ;
        RECT 78.820 3.615 78.990 4.510 ;
        RECT 80.100 3.860 80.260 9.030 ;
        RECT 81.215 8.940 81.540 9.030 ;
        RECT 83.605 9.145 83.930 9.270 ;
        RECT 86.660 9.225 86.830 9.720 ;
        RECT 83.605 9.140 84.310 9.145 ;
        RECT 86.605 9.140 86.885 9.225 ;
        RECT 83.605 8.975 86.885 9.140 ;
        RECT 83.605 8.945 83.930 8.975 ;
        RECT 84.310 8.970 86.885 8.975 ;
        RECT 80.415 8.565 80.735 8.890 ;
        RECT 86.605 8.885 86.885 8.970 ;
        RECT 96.680 9.200 96.840 9.720 ;
        RECT 100.150 9.585 100.475 9.910 ;
        RECT 97.795 9.200 98.120 9.265 ;
        RECT 96.680 9.030 98.120 9.200 ;
        RECT 80.445 8.330 80.615 8.565 ;
        RECT 80.445 8.155 80.620 8.330 ;
        RECT 80.445 7.980 81.420 8.155 ;
        RECT 80.415 3.860 80.735 3.980 ;
        RECT 80.100 3.690 80.735 3.860 ;
        RECT 80.415 3.660 80.735 3.690 ;
        RECT 78.745 3.290 79.070 3.615 ;
        RECT 81.245 3.610 81.420 7.980 ;
        RECT 90.925 7.415 91.205 7.440 ;
        RECT 90.925 7.095 91.215 7.415 ;
        RECT 90.925 7.065 91.205 7.095 ;
        RECT 91.975 7.065 92.255 7.440 ;
        RECT 93.335 7.325 93.595 7.415 ;
        RECT 92.715 7.185 93.595 7.325 ;
        RECT 91.295 6.045 91.575 6.420 ;
        RECT 90.615 3.655 90.895 4.035 ;
        RECT 91.355 4.015 91.495 6.045 ;
        RECT 92.035 5.285 92.175 7.065 ;
        RECT 92.715 5.400 92.855 7.185 ;
        RECT 93.335 7.095 93.595 7.185 ;
        RECT 94.355 6.075 94.615 6.395 ;
        RECT 92.035 5.145 92.515 5.285 ;
        RECT 91.955 4.345 92.235 4.720 ;
        RECT 91.295 3.695 91.555 4.015 ;
        RECT 92.375 3.695 92.515 5.145 ;
        RECT 92.655 5.025 92.935 5.400 ;
        RECT 92.655 4.005 92.935 4.380 ;
        RECT 94.415 4.355 94.555 6.075 ;
        RECT 94.740 4.695 95.065 4.805 ;
        RECT 94.740 4.510 95.570 4.695 ;
        RECT 94.740 4.480 95.065 4.510 ;
        RECT 94.355 4.035 94.615 4.355 ;
        RECT 81.190 3.260 81.540 3.610 ;
        RECT 92.315 3.355 92.575 3.695 ;
        RECT 95.400 3.615 95.570 4.510 ;
        RECT 96.680 3.860 96.840 9.030 ;
        RECT 97.795 8.940 98.120 9.030 ;
        RECT 96.995 8.565 97.315 8.890 ;
        RECT 97.025 8.330 97.195 8.565 ;
        RECT 97.025 8.155 97.200 8.330 ;
        RECT 97.025 7.980 98.000 8.155 ;
        RECT 96.995 3.860 97.315 3.980 ;
        RECT 96.680 3.690 97.315 3.860 ;
        RECT 96.995 3.660 97.315 3.690 ;
        RECT 95.325 3.290 95.650 3.615 ;
        RECT 97.825 3.610 98.000 7.980 ;
        RECT 97.770 3.260 98.120 3.610 ;
      LAYER met3 ;
        RECT 19.740 9.615 20.110 9.675 ;
        RECT 36.325 9.615 36.695 9.675 ;
        RECT 52.910 9.615 53.280 9.675 ;
        RECT 69.495 9.615 69.865 9.675 ;
        RECT 86.075 9.615 86.445 9.675 ;
        RECT 19.740 9.315 24.970 9.615 ;
        RECT 36.325 9.315 41.555 9.615 ;
        RECT 52.910 9.315 58.140 9.615 ;
        RECT 69.495 9.315 74.725 9.615 ;
        RECT 86.075 9.315 91.305 9.615 ;
        RECT 19.740 9.305 20.110 9.315 ;
        RECT 24.590 7.425 24.890 9.315 ;
        RECT 36.325 9.305 36.695 9.315 ;
        RECT 41.175 7.425 41.475 9.315 ;
        RECT 52.910 9.305 53.280 9.315 ;
        RECT 57.760 7.425 58.060 9.315 ;
        RECT 69.495 9.305 69.865 9.315 ;
        RECT 74.345 7.425 74.645 9.315 ;
        RECT 86.075 9.305 86.445 9.315 ;
        RECT 90.925 7.425 91.225 9.315 ;
        RECT 23.960 7.410 24.900 7.425 ;
        RECT 25.600 7.410 25.945 7.420 ;
        RECT 23.960 7.405 25.945 7.410 ;
        RECT 40.545 7.410 41.485 7.425 ;
        RECT 42.185 7.410 42.530 7.420 ;
        RECT 40.545 7.405 42.530 7.410 ;
        RECT 57.130 7.410 58.070 7.425 ;
        RECT 58.770 7.410 59.115 7.420 ;
        RECT 57.130 7.405 59.115 7.410 ;
        RECT 73.715 7.410 74.655 7.425 ;
        RECT 75.355 7.410 75.700 7.420 ;
        RECT 73.715 7.405 75.700 7.410 ;
        RECT 90.295 7.410 91.235 7.425 ;
        RECT 91.935 7.410 92.280 7.420 ;
        RECT 90.295 7.405 92.280 7.410 ;
        RECT 23.960 7.110 26.410 7.405 ;
        RECT 23.960 7.105 24.900 7.110 ;
        RECT 23.960 5.390 24.260 7.105 ;
        RECT 24.560 7.075 24.900 7.105 ;
        RECT 25.395 7.105 26.410 7.110 ;
        RECT 40.545 7.110 42.995 7.405 ;
        RECT 40.545 7.105 41.485 7.110 ;
        RECT 25.395 7.095 25.945 7.105 ;
        RECT 25.600 7.085 25.945 7.095 ;
        RECT 25.600 7.075 25.940 7.085 ;
        RECT 24.920 6.385 25.265 6.400 ;
        RECT 24.920 6.085 25.730 6.385 ;
        RECT 24.920 6.055 25.265 6.085 ;
        RECT 40.545 5.390 40.845 7.105 ;
        RECT 41.145 7.075 41.485 7.105 ;
        RECT 41.980 7.105 42.995 7.110 ;
        RECT 57.130 7.110 59.580 7.405 ;
        RECT 57.130 7.105 58.070 7.110 ;
        RECT 41.980 7.095 42.530 7.105 ;
        RECT 42.185 7.085 42.530 7.095 ;
        RECT 42.185 7.075 42.525 7.085 ;
        RECT 41.505 6.385 41.850 6.400 ;
        RECT 41.505 6.085 42.315 6.385 ;
        RECT 41.505 6.055 41.850 6.085 ;
        RECT 57.130 5.390 57.430 7.105 ;
        RECT 57.730 7.075 58.070 7.105 ;
        RECT 58.565 7.105 59.580 7.110 ;
        RECT 73.715 7.110 76.165 7.405 ;
        RECT 73.715 7.105 74.655 7.110 ;
        RECT 58.565 7.095 59.115 7.105 ;
        RECT 58.770 7.085 59.115 7.095 ;
        RECT 58.770 7.075 59.110 7.085 ;
        RECT 58.090 6.385 58.435 6.400 ;
        RECT 58.090 6.085 58.900 6.385 ;
        RECT 58.090 6.055 58.435 6.085 ;
        RECT 73.715 5.390 74.015 7.105 ;
        RECT 74.315 7.075 74.655 7.105 ;
        RECT 75.150 7.105 76.165 7.110 ;
        RECT 90.295 7.110 92.745 7.405 ;
        RECT 90.295 7.105 91.235 7.110 ;
        RECT 75.150 7.095 75.700 7.105 ;
        RECT 75.355 7.085 75.700 7.095 ;
        RECT 75.355 7.075 75.695 7.085 ;
        RECT 74.675 6.385 75.020 6.400 ;
        RECT 74.675 6.085 75.485 6.385 ;
        RECT 74.675 6.055 75.020 6.085 ;
        RECT 90.295 5.390 90.595 7.105 ;
        RECT 90.895 7.075 91.235 7.105 ;
        RECT 91.730 7.105 92.745 7.110 ;
        RECT 91.730 7.095 92.280 7.105 ;
        RECT 91.935 7.085 92.280 7.095 ;
        RECT 91.935 7.075 92.275 7.085 ;
        RECT 91.255 6.385 91.600 6.400 ;
        RECT 91.255 6.085 92.065 6.385 ;
        RECT 91.255 6.055 91.600 6.085 ;
        RECT 23.960 5.385 26.615 5.390 ;
        RECT 40.545 5.385 43.200 5.390 ;
        RECT 57.130 5.385 59.785 5.390 ;
        RECT 73.715 5.385 76.370 5.390 ;
        RECT 90.295 5.385 92.950 5.390 ;
        RECT 23.960 5.365 26.625 5.385 ;
        RECT 40.545 5.365 43.210 5.385 ;
        RECT 57.130 5.365 59.795 5.385 ;
        RECT 73.715 5.365 76.380 5.385 ;
        RECT 90.295 5.365 92.960 5.385 ;
        RECT 23.960 5.065 27.090 5.365 ;
        RECT 40.545 5.065 43.675 5.365 ;
        RECT 57.130 5.065 60.260 5.365 ;
        RECT 73.715 5.065 76.845 5.365 ;
        RECT 90.295 5.065 93.425 5.365 ;
        RECT 23.960 5.060 26.625 5.065 ;
        RECT 40.545 5.060 43.210 5.065 ;
        RECT 57.130 5.060 59.795 5.065 ;
        RECT 73.715 5.060 76.380 5.065 ;
        RECT 90.295 5.060 92.960 5.065 ;
        RECT 26.280 5.035 26.625 5.060 ;
        RECT 42.865 5.035 43.210 5.060 ;
        RECT 59.450 5.035 59.795 5.060 ;
        RECT 76.035 5.035 76.380 5.060 ;
        RECT 92.615 5.035 92.960 5.060 ;
        RECT 26.300 4.995 26.600 5.035 ;
        RECT 42.885 4.995 43.185 5.035 ;
        RECT 59.470 4.995 59.770 5.035 ;
        RECT 76.055 4.995 76.355 5.035 ;
        RECT 92.635 4.995 92.935 5.035 ;
        RECT 25.590 4.685 25.930 4.705 ;
        RECT 42.175 4.685 42.515 4.705 ;
        RECT 58.760 4.685 59.100 4.705 ;
        RECT 75.345 4.685 75.685 4.705 ;
        RECT 91.925 4.685 92.265 4.705 ;
        RECT 25.120 4.385 25.930 4.685 ;
        RECT 41.705 4.385 42.515 4.685 ;
        RECT 58.290 4.385 59.100 4.685 ;
        RECT 74.875 4.385 75.685 4.685 ;
        RECT 91.455 4.385 92.265 4.685 ;
        RECT 25.590 4.355 25.930 4.385 ;
        RECT 26.290 4.355 26.625 4.360 ;
        RECT 42.175 4.355 42.515 4.385 ;
        RECT 42.875 4.355 43.210 4.360 ;
        RECT 58.760 4.355 59.100 4.385 ;
        RECT 59.460 4.355 59.795 4.360 ;
        RECT 75.345 4.355 75.685 4.385 ;
        RECT 76.045 4.355 76.380 4.360 ;
        RECT 91.925 4.355 92.265 4.385 ;
        RECT 92.625 4.355 92.960 4.360 ;
        RECT 26.280 4.345 26.625 4.355 ;
        RECT 42.865 4.345 43.210 4.355 ;
        RECT 59.450 4.345 59.795 4.355 ;
        RECT 76.035 4.345 76.380 4.355 ;
        RECT 92.615 4.345 92.960 4.355 ;
        RECT 26.280 4.045 27.090 4.345 ;
        RECT 42.865 4.045 43.675 4.345 ;
        RECT 59.450 4.045 60.260 4.345 ;
        RECT 76.035 4.045 76.845 4.345 ;
        RECT 92.615 4.045 93.425 4.345 ;
        RECT 26.280 4.025 26.625 4.045 ;
        RECT 42.865 4.025 43.210 4.045 ;
        RECT 59.450 4.025 59.795 4.045 ;
        RECT 76.035 4.025 76.380 4.045 ;
        RECT 92.615 4.025 92.960 4.045 ;
        RECT 26.280 4.015 26.620 4.025 ;
        RECT 42.865 4.015 43.205 4.025 ;
        RECT 59.450 4.015 59.790 4.025 ;
        RECT 76.035 4.015 76.375 4.025 ;
        RECT 92.615 4.015 92.955 4.025 ;
        RECT 24.240 4.005 24.585 4.015 ;
        RECT 40.825 4.005 41.170 4.015 ;
        RECT 57.410 4.005 57.755 4.015 ;
        RECT 73.995 4.005 74.340 4.015 ;
        RECT 90.575 4.005 90.920 4.015 ;
        RECT 23.780 3.705 24.585 4.005 ;
        RECT 40.365 3.705 41.170 4.005 ;
        RECT 56.950 3.705 57.755 4.005 ;
        RECT 73.535 3.705 74.340 4.005 ;
        RECT 90.115 3.705 90.920 4.005 ;
        RECT 24.140 3.695 24.585 3.705 ;
        RECT 40.725 3.695 41.170 3.705 ;
        RECT 57.310 3.695 57.755 3.705 ;
        RECT 73.895 3.695 74.340 3.705 ;
        RECT 90.475 3.695 90.920 3.705 ;
        RECT 24.240 3.675 24.585 3.695 ;
        RECT 40.825 3.675 41.170 3.695 ;
        RECT 57.410 3.675 57.755 3.695 ;
        RECT 73.995 3.675 74.340 3.695 ;
        RECT 90.575 3.675 90.920 3.695 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r1
MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r1
  CLASS BLOCK ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ct_8_b0r1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 103.925 BY 12.460 ;
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 35.880 8.225 36.050 9.495 ;
        RECT 47.565 8.465 47.735 9.505 ;
        RECT 47.560 8.225 47.740 8.465 ;
        RECT 47.565 2.955 47.735 4.225 ;
      LAYER met1 ;
        RECT 35.785 8.400 36.125 8.495 ;
        RECT 35.785 8.395 36.140 8.400 ;
        RECT 35.785 8.365 36.280 8.395 ;
        RECT 38.105 8.365 38.445 8.455 ;
        RECT 35.785 8.200 38.445 8.365 ;
        RECT 35.785 8.155 36.125 8.200 ;
        RECT 38.105 8.175 38.445 8.200 ;
        RECT 47.490 8.405 47.815 8.465 ;
        RECT 47.490 8.235 47.965 8.405 ;
        RECT 47.490 8.140 47.815 8.235 ;
        RECT 47.490 4.790 47.815 5.115 ;
        RECT 47.570 4.255 47.740 4.790 ;
        RECT 47.505 4.225 47.795 4.255 ;
        RECT 47.505 4.055 47.965 4.225 ;
        RECT 47.505 4.025 47.795 4.055 ;
      LAYER met2 ;
        RECT 38.190 9.320 47.740 9.490 ;
        RECT 35.765 8.140 36.140 8.510 ;
        RECT 38.190 8.485 38.360 9.320 ;
        RECT 38.135 8.145 38.415 8.485 ;
        RECT 47.570 8.465 47.740 9.320 ;
        RECT 47.490 8.140 47.815 8.465 ;
        RECT 47.560 5.115 47.730 8.140 ;
        RECT 47.490 4.790 47.815 5.115 ;
      LAYER met3 ;
        RECT 35.790 8.510 36.120 12.445 ;
        RECT 35.765 8.140 36.140 8.510 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 53.100 8.225 53.270 9.495 ;
        RECT 64.785 8.465 64.955 9.505 ;
        RECT 64.780 8.225 64.960 8.465 ;
        RECT 64.785 2.955 64.955 4.225 ;
      LAYER met1 ;
        RECT 53.005 8.400 53.345 8.495 ;
        RECT 53.005 8.395 53.360 8.400 ;
        RECT 53.005 8.365 53.500 8.395 ;
        RECT 55.325 8.365 55.665 8.455 ;
        RECT 53.005 8.200 55.665 8.365 ;
        RECT 53.005 8.155 53.345 8.200 ;
        RECT 55.325 8.175 55.665 8.200 ;
        RECT 64.710 8.405 65.035 8.465 ;
        RECT 64.710 8.235 65.185 8.405 ;
        RECT 64.710 8.140 65.035 8.235 ;
        RECT 64.710 4.790 65.035 5.115 ;
        RECT 64.790 4.255 64.960 4.790 ;
        RECT 64.725 4.225 65.015 4.255 ;
        RECT 64.725 4.055 65.185 4.225 ;
        RECT 64.725 4.025 65.015 4.055 ;
      LAYER met2 ;
        RECT 55.410 9.320 64.960 9.490 ;
        RECT 52.985 8.140 53.360 8.510 ;
        RECT 55.410 8.485 55.580 9.320 ;
        RECT 55.355 8.145 55.635 8.485 ;
        RECT 64.790 8.465 64.960 9.320 ;
        RECT 64.710 8.140 65.035 8.465 ;
        RECT 64.780 5.115 64.950 8.140 ;
        RECT 64.710 4.790 65.035 5.115 ;
      LAYER met3 ;
        RECT 53.010 8.510 53.340 12.445 ;
        RECT 52.985 8.140 53.360 8.510 ;
    END
  END s3
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 103.375 4.010 103.550 5.155 ;
        RECT 103.375 3.575 103.545 4.010 ;
        RECT 103.380 1.865 103.550 2.375 ;
      LAYER met1 ;
        RECT 103.315 3.540 103.605 3.775 ;
        RECT 103.315 3.535 103.545 3.540 ;
        RECT 103.375 2.435 103.545 3.535 ;
        RECT 103.315 2.175 103.610 2.435 ;
    END
  END X5_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 86.155 4.010 86.330 5.155 ;
        RECT 86.155 3.575 86.325 4.010 ;
        RECT 86.160 1.865 86.330 2.375 ;
      LAYER met1 ;
        RECT 86.095 3.540 86.385 3.775 ;
        RECT 86.095 3.535 86.325 3.540 ;
        RECT 86.155 2.435 86.325 3.535 ;
        RECT 86.095 2.175 86.390 2.435 ;
    END
  END X4_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 68.935 4.010 69.110 5.155 ;
        RECT 68.935 3.575 69.105 4.010 ;
        RECT 68.940 1.865 69.110 2.375 ;
      LAYER met1 ;
        RECT 68.875 3.540 69.165 3.775 ;
        RECT 68.875 3.535 69.105 3.540 ;
        RECT 68.935 2.435 69.105 3.535 ;
        RECT 68.875 2.175 69.170 2.435 ;
    END
  END X3_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 51.715 4.010 51.890 5.155 ;
        RECT 51.715 3.575 51.885 4.010 ;
        RECT 51.720 1.865 51.890 2.375 ;
      LAYER met1 ;
        RECT 51.655 3.540 51.945 3.775 ;
        RECT 51.655 3.535 51.885 3.540 ;
        RECT 51.715 2.435 51.885 3.535 ;
        RECT 51.655 2.175 51.950 2.435 ;
    END
  END X2_Y1
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 34.495 4.010 34.670 5.155 ;
        RECT 34.495 3.575 34.665 4.010 ;
        RECT 34.500 1.865 34.670 2.375 ;
      LAYER met1 ;
        RECT 34.435 3.540 34.725 3.775 ;
        RECT 34.435 3.535 34.665 3.540 ;
        RECT 34.495 2.435 34.665 3.535 ;
        RECT 34.435 2.175 34.730 2.435 ;
    END
  END X1_Y1
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 87.540 8.225 87.710 9.495 ;
        RECT 99.225 8.465 99.395 9.505 ;
        RECT 99.220 8.225 99.400 8.465 ;
        RECT 99.225 2.955 99.395 4.225 ;
      LAYER met1 ;
        RECT 87.445 8.400 87.785 8.495 ;
        RECT 87.445 8.395 87.800 8.400 ;
        RECT 87.445 8.365 87.940 8.395 ;
        RECT 89.765 8.365 90.105 8.455 ;
        RECT 87.445 8.200 90.105 8.365 ;
        RECT 87.445 8.155 87.785 8.200 ;
        RECT 89.765 8.175 90.105 8.200 ;
        RECT 99.150 8.405 99.475 8.465 ;
        RECT 99.150 8.235 99.625 8.405 ;
        RECT 99.150 8.140 99.475 8.235 ;
        RECT 99.150 4.790 99.475 5.115 ;
        RECT 99.230 4.255 99.400 4.790 ;
        RECT 99.165 4.225 99.455 4.255 ;
        RECT 99.165 4.055 99.625 4.225 ;
        RECT 99.165 4.025 99.455 4.055 ;
      LAYER met2 ;
        RECT 89.850 9.320 99.400 9.490 ;
        RECT 87.425 8.140 87.800 8.510 ;
        RECT 89.850 8.485 90.020 9.320 ;
        RECT 89.795 8.145 90.075 8.485 ;
        RECT 99.230 8.465 99.400 9.320 ;
        RECT 99.150 8.140 99.475 8.465 ;
        RECT 99.220 5.115 99.390 8.140 ;
        RECT 99.150 4.790 99.475 5.115 ;
      LAYER met3 ;
        RECT 87.450 8.510 87.780 12.445 ;
        RECT 87.425 8.140 87.800 8.510 ;
    END
  END s5
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 70.320 8.225 70.490 9.495 ;
        RECT 82.005 8.465 82.175 9.505 ;
        RECT 82.000 8.225 82.180 8.465 ;
        RECT 82.005 2.955 82.175 4.225 ;
      LAYER met1 ;
        RECT 70.225 8.400 70.565 8.495 ;
        RECT 70.225 8.395 70.580 8.400 ;
        RECT 70.225 8.365 70.720 8.395 ;
        RECT 72.545 8.365 72.885 8.455 ;
        RECT 70.225 8.200 72.885 8.365 ;
        RECT 70.225 8.155 70.565 8.200 ;
        RECT 72.545 8.175 72.885 8.200 ;
        RECT 81.930 8.405 82.255 8.465 ;
        RECT 81.930 8.235 82.405 8.405 ;
        RECT 81.930 8.140 82.255 8.235 ;
        RECT 81.930 4.790 82.255 5.115 ;
        RECT 82.010 4.255 82.180 4.790 ;
        RECT 81.945 4.225 82.235 4.255 ;
        RECT 81.945 4.055 82.405 4.225 ;
        RECT 81.945 4.025 82.235 4.055 ;
      LAYER met2 ;
        RECT 72.630 9.320 82.180 9.490 ;
        RECT 70.205 8.140 70.580 8.510 ;
        RECT 72.630 8.485 72.800 9.320 ;
        RECT 72.575 8.145 72.855 8.485 ;
        RECT 82.010 8.465 82.180 9.320 ;
        RECT 81.930 8.140 82.255 8.465 ;
        RECT 82.000 5.115 82.170 8.140 ;
        RECT 81.930 4.790 82.255 5.115 ;
      LAYER met3 ;
        RECT 70.230 8.510 70.560 12.445 ;
        RECT 70.205 8.140 70.580 8.510 ;
    END
  END s4
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 15.250 8.235 15.420 9.505 ;
      LAYER met1 ;
        RECT 15.190 8.430 15.480 8.435 ;
        RECT 15.190 8.405 15.485 8.430 ;
        RECT 15.190 8.235 15.650 8.405 ;
        RECT 15.190 8.205 15.485 8.235 ;
        RECT 15.195 8.200 15.485 8.205 ;
    END
  END start
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 10.860 103.925 12.460 ;
        RECT 15.240 10.235 15.410 10.860 ;
        RECT 18.480 10.855 21.230 10.860 ;
        RECT 18.650 10.225 18.820 10.855 ;
        RECT 19.605 10.305 19.775 10.585 ;
        RECT 19.605 10.135 19.835 10.305 ;
        RECT 19.665 8.525 19.835 10.135 ;
        RECT 19.605 8.355 19.835 8.525 ;
        RECT 21.610 8.530 21.895 10.860 ;
        RECT 22.180 8.530 22.465 10.860 ;
        RECT 22.750 8.530 23.035 10.860 ;
        RECT 23.320 8.530 23.605 10.860 ;
        RECT 23.890 8.530 24.175 10.860 ;
        RECT 24.460 8.530 24.745 10.860 ;
        RECT 25.030 8.530 25.315 10.860 ;
        RECT 25.600 8.530 25.885 10.860 ;
        RECT 26.170 8.530 26.450 10.860 ;
        RECT 26.735 8.530 27.020 10.860 ;
        RECT 27.305 8.530 27.590 10.860 ;
        RECT 27.875 8.530 28.160 10.860 ;
        RECT 28.730 8.530 28.970 10.860 ;
        RECT 30.335 10.235 30.505 10.860 ;
        RECT 33.080 10.235 33.250 10.860 ;
        RECT 34.070 10.235 34.240 10.860 ;
        RECT 35.700 10.855 38.450 10.860 ;
        RECT 35.870 10.225 36.040 10.855 ;
        RECT 36.825 10.305 36.995 10.585 ;
        RECT 36.825 10.135 37.055 10.305 ;
        RECT 21.610 8.360 28.970 8.530 ;
        RECT 36.885 8.525 37.055 10.135 ;
        RECT 19.605 7.295 19.775 8.355 ;
        RECT 22.155 7.560 22.465 8.360 ;
        RECT 22.165 7.340 22.500 7.390 ;
        RECT 24.085 7.340 24.255 8.360 ;
        RECT 24.455 7.560 24.765 8.360 ;
        RECT 26.735 7.560 27.045 8.360 ;
        RECT 28.115 7.560 28.425 8.360 ;
        RECT 36.825 8.355 37.055 8.525 ;
        RECT 38.830 8.530 39.115 10.860 ;
        RECT 39.400 8.530 39.685 10.860 ;
        RECT 39.970 8.530 40.255 10.860 ;
        RECT 40.540 8.530 40.825 10.860 ;
        RECT 41.110 8.530 41.395 10.860 ;
        RECT 41.680 8.530 41.965 10.860 ;
        RECT 42.250 8.530 42.535 10.860 ;
        RECT 42.820 8.530 43.105 10.860 ;
        RECT 43.390 8.530 43.670 10.860 ;
        RECT 43.955 8.530 44.240 10.860 ;
        RECT 44.525 8.530 44.810 10.860 ;
        RECT 45.095 8.530 45.380 10.860 ;
        RECT 45.950 8.530 46.190 10.860 ;
        RECT 47.555 10.235 47.725 10.860 ;
        RECT 50.300 10.235 50.470 10.860 ;
        RECT 51.290 10.235 51.460 10.860 ;
        RECT 52.920 10.855 55.670 10.860 ;
        RECT 53.090 10.225 53.260 10.855 ;
        RECT 54.045 10.305 54.215 10.585 ;
        RECT 54.045 10.135 54.275 10.305 ;
        RECT 38.830 8.360 46.190 8.530 ;
        RECT 54.105 8.525 54.275 10.135 ;
        RECT 24.465 7.340 24.800 7.390 ;
        RECT 21.695 7.170 22.500 7.340 ;
        RECT 24.075 7.170 24.800 7.340 ;
        RECT 36.825 7.295 36.995 8.355 ;
        RECT 39.375 7.560 39.685 8.360 ;
        RECT 39.385 7.340 39.720 7.390 ;
        RECT 41.305 7.340 41.475 8.360 ;
        RECT 41.675 7.560 41.985 8.360 ;
        RECT 43.955 7.560 44.265 8.360 ;
        RECT 45.335 7.560 45.645 8.360 ;
        RECT 54.045 8.355 54.275 8.525 ;
        RECT 56.050 8.530 56.335 10.860 ;
        RECT 56.620 8.530 56.905 10.860 ;
        RECT 57.190 8.530 57.475 10.860 ;
        RECT 57.760 8.530 58.045 10.860 ;
        RECT 58.330 8.530 58.615 10.860 ;
        RECT 58.900 8.530 59.185 10.860 ;
        RECT 59.470 8.530 59.755 10.860 ;
        RECT 60.040 8.530 60.325 10.860 ;
        RECT 60.610 8.530 60.890 10.860 ;
        RECT 61.175 8.530 61.460 10.860 ;
        RECT 61.745 8.530 62.030 10.860 ;
        RECT 62.315 8.530 62.600 10.860 ;
        RECT 63.170 8.530 63.410 10.860 ;
        RECT 64.775 10.235 64.945 10.860 ;
        RECT 67.520 10.235 67.690 10.860 ;
        RECT 68.510 10.235 68.680 10.860 ;
        RECT 70.140 10.855 72.890 10.860 ;
        RECT 70.310 10.225 70.480 10.855 ;
        RECT 71.265 10.305 71.435 10.585 ;
        RECT 71.265 10.135 71.495 10.305 ;
        RECT 56.050 8.360 63.410 8.530 ;
        RECT 71.325 8.525 71.495 10.135 ;
        RECT 41.685 7.340 42.020 7.390 ;
        RECT 38.915 7.170 39.720 7.340 ;
        RECT 41.295 7.170 42.020 7.340 ;
        RECT 54.045 7.295 54.215 8.355 ;
        RECT 56.595 7.560 56.905 8.360 ;
        RECT 56.605 7.340 56.940 7.390 ;
        RECT 58.525 7.340 58.695 8.360 ;
        RECT 58.895 7.560 59.205 8.360 ;
        RECT 61.175 7.560 61.485 8.360 ;
        RECT 62.555 7.560 62.865 8.360 ;
        RECT 71.265 8.355 71.495 8.525 ;
        RECT 73.270 8.530 73.555 10.860 ;
        RECT 73.840 8.530 74.125 10.860 ;
        RECT 74.410 8.530 74.695 10.860 ;
        RECT 74.980 8.530 75.265 10.860 ;
        RECT 75.550 8.530 75.835 10.860 ;
        RECT 76.120 8.530 76.405 10.860 ;
        RECT 76.690 8.530 76.975 10.860 ;
        RECT 77.260 8.530 77.545 10.860 ;
        RECT 77.830 8.530 78.110 10.860 ;
        RECT 78.395 8.530 78.680 10.860 ;
        RECT 78.965 8.530 79.250 10.860 ;
        RECT 79.535 8.530 79.820 10.860 ;
        RECT 80.390 8.530 80.630 10.860 ;
        RECT 81.995 10.235 82.165 10.860 ;
        RECT 84.740 10.235 84.910 10.860 ;
        RECT 85.730 10.235 85.900 10.860 ;
        RECT 87.360 10.855 90.110 10.860 ;
        RECT 87.530 10.225 87.700 10.855 ;
        RECT 88.485 10.305 88.655 10.585 ;
        RECT 88.485 10.135 88.715 10.305 ;
        RECT 73.270 8.360 80.630 8.530 ;
        RECT 88.545 8.525 88.715 10.135 ;
        RECT 58.905 7.340 59.240 7.390 ;
        RECT 56.135 7.170 56.940 7.340 ;
        RECT 58.515 7.170 59.240 7.340 ;
        RECT 71.265 7.295 71.435 8.355 ;
        RECT 73.815 7.560 74.125 8.360 ;
        RECT 73.825 7.340 74.160 7.390 ;
        RECT 75.745 7.340 75.915 8.360 ;
        RECT 76.115 7.560 76.425 8.360 ;
        RECT 78.395 7.560 78.705 8.360 ;
        RECT 79.775 7.560 80.085 8.360 ;
        RECT 88.485 8.355 88.715 8.525 ;
        RECT 90.490 8.530 90.775 10.860 ;
        RECT 91.060 8.530 91.345 10.860 ;
        RECT 91.630 8.530 91.915 10.860 ;
        RECT 92.200 8.530 92.485 10.860 ;
        RECT 92.770 8.530 93.055 10.860 ;
        RECT 93.340 8.530 93.625 10.860 ;
        RECT 93.910 8.530 94.195 10.860 ;
        RECT 94.480 8.530 94.765 10.860 ;
        RECT 95.050 8.530 95.330 10.860 ;
        RECT 95.615 8.530 95.900 10.860 ;
        RECT 96.185 8.530 96.470 10.860 ;
        RECT 96.755 8.530 97.040 10.860 ;
        RECT 97.610 8.530 97.850 10.860 ;
        RECT 99.215 10.235 99.385 10.860 ;
        RECT 101.960 10.235 102.130 10.860 ;
        RECT 102.950 10.235 103.120 10.860 ;
        RECT 90.490 8.360 97.850 8.530 ;
        RECT 76.125 7.340 76.460 7.390 ;
        RECT 73.355 7.170 74.160 7.340 ;
        RECT 75.735 7.170 76.460 7.340 ;
        RECT 88.485 7.295 88.655 8.355 ;
        RECT 91.035 7.560 91.345 8.360 ;
        RECT 91.045 7.340 91.380 7.390 ;
        RECT 92.965 7.340 93.135 8.360 ;
        RECT 93.335 7.560 93.645 8.360 ;
        RECT 95.615 7.560 95.925 8.360 ;
        RECT 96.995 7.560 97.305 8.360 ;
        RECT 93.345 7.340 93.680 7.390 ;
        RECT 90.575 7.170 91.380 7.340 ;
        RECT 92.955 7.170 93.680 7.340 ;
        RECT 22.165 7.120 22.500 7.170 ;
        RECT 24.465 7.120 24.800 7.170 ;
        RECT 39.385 7.120 39.720 7.170 ;
        RECT 41.685 7.120 42.020 7.170 ;
        RECT 56.605 7.120 56.940 7.170 ;
        RECT 58.905 7.120 59.240 7.170 ;
        RECT 73.825 7.120 74.160 7.170 ;
        RECT 76.125 7.120 76.460 7.170 ;
        RECT 91.045 7.120 91.380 7.170 ;
        RECT 93.345 7.120 93.680 7.170 ;
      LAYER met1 ;
        RECT 0.000 10.860 103.925 12.460 ;
        RECT 18.480 10.855 21.230 10.860 ;
        RECT 19.200 8.775 19.370 10.855 ;
        RECT 19.605 8.775 19.895 8.805 ;
        RECT 19.200 8.595 19.895 8.775 ;
        RECT 19.605 8.575 19.895 8.595 ;
        RECT 21.610 8.685 21.895 10.860 ;
        RECT 22.180 8.685 22.465 10.860 ;
        RECT 22.750 8.685 23.035 10.860 ;
        RECT 23.320 8.685 23.605 10.860 ;
        RECT 23.890 8.685 24.175 10.860 ;
        RECT 24.460 8.685 24.745 10.860 ;
        RECT 25.030 8.685 25.315 10.860 ;
        RECT 25.600 8.685 25.885 10.860 ;
        RECT 26.170 8.685 26.450 10.860 ;
        RECT 26.735 8.685 27.020 10.860 ;
        RECT 27.305 8.685 27.590 10.860 ;
        RECT 27.875 8.685 28.160 10.860 ;
        RECT 28.730 8.685 28.970 10.860 ;
        RECT 35.700 10.855 38.450 10.860 ;
        RECT 21.610 8.330 28.970 8.685 ;
        RECT 36.420 8.775 36.590 10.855 ;
        RECT 36.825 8.775 37.115 8.805 ;
        RECT 36.420 8.595 37.115 8.775 ;
        RECT 36.825 8.575 37.115 8.595 ;
        RECT 38.830 8.685 39.115 10.860 ;
        RECT 39.400 8.685 39.685 10.860 ;
        RECT 39.970 8.685 40.255 10.860 ;
        RECT 40.540 8.685 40.825 10.860 ;
        RECT 41.110 8.685 41.395 10.860 ;
        RECT 41.680 8.685 41.965 10.860 ;
        RECT 42.250 8.685 42.535 10.860 ;
        RECT 42.820 8.685 43.105 10.860 ;
        RECT 43.390 8.685 43.670 10.860 ;
        RECT 43.955 8.685 44.240 10.860 ;
        RECT 44.525 8.685 44.810 10.860 ;
        RECT 45.095 8.685 45.380 10.860 ;
        RECT 45.950 8.685 46.190 10.860 ;
        RECT 52.920 10.855 55.670 10.860 ;
        RECT 38.830 8.330 46.190 8.685 ;
        RECT 53.640 8.775 53.810 10.855 ;
        RECT 54.045 8.775 54.335 8.805 ;
        RECT 53.640 8.595 54.335 8.775 ;
        RECT 54.045 8.575 54.335 8.595 ;
        RECT 56.050 8.685 56.335 10.860 ;
        RECT 56.620 8.685 56.905 10.860 ;
        RECT 57.190 8.685 57.475 10.860 ;
        RECT 57.760 8.685 58.045 10.860 ;
        RECT 58.330 8.685 58.615 10.860 ;
        RECT 58.900 8.685 59.185 10.860 ;
        RECT 59.470 8.685 59.755 10.860 ;
        RECT 60.040 8.685 60.325 10.860 ;
        RECT 60.610 8.685 60.890 10.860 ;
        RECT 61.175 8.685 61.460 10.860 ;
        RECT 61.745 8.685 62.030 10.860 ;
        RECT 62.315 8.685 62.600 10.860 ;
        RECT 63.170 8.685 63.410 10.860 ;
        RECT 70.140 10.855 72.890 10.860 ;
        RECT 56.050 8.330 63.410 8.685 ;
        RECT 70.860 8.775 71.030 10.855 ;
        RECT 71.265 8.775 71.555 8.805 ;
        RECT 70.860 8.595 71.555 8.775 ;
        RECT 71.265 8.575 71.555 8.595 ;
        RECT 73.270 8.685 73.555 10.860 ;
        RECT 73.840 8.685 74.125 10.860 ;
        RECT 74.410 8.685 74.695 10.860 ;
        RECT 74.980 8.685 75.265 10.860 ;
        RECT 75.550 8.685 75.835 10.860 ;
        RECT 76.120 8.685 76.405 10.860 ;
        RECT 76.690 8.685 76.975 10.860 ;
        RECT 77.260 8.685 77.545 10.860 ;
        RECT 77.830 8.685 78.110 10.860 ;
        RECT 78.395 8.685 78.680 10.860 ;
        RECT 78.965 8.685 79.250 10.860 ;
        RECT 79.535 8.685 79.820 10.860 ;
        RECT 80.390 8.685 80.630 10.860 ;
        RECT 87.360 10.855 90.110 10.860 ;
        RECT 73.270 8.330 80.630 8.685 ;
        RECT 88.080 8.775 88.250 10.855 ;
        RECT 88.485 8.775 88.775 8.805 ;
        RECT 88.080 8.595 88.775 8.775 ;
        RECT 88.485 8.575 88.775 8.595 ;
        RECT 90.490 8.685 90.775 10.860 ;
        RECT 91.060 8.685 91.345 10.860 ;
        RECT 91.630 8.685 91.915 10.860 ;
        RECT 92.200 8.685 92.485 10.860 ;
        RECT 92.770 8.685 93.055 10.860 ;
        RECT 93.340 8.685 93.625 10.860 ;
        RECT 93.910 8.685 94.195 10.860 ;
        RECT 94.480 8.685 94.765 10.860 ;
        RECT 95.050 8.685 95.330 10.860 ;
        RECT 95.615 8.685 95.900 10.860 ;
        RECT 96.185 8.685 96.470 10.860 ;
        RECT 96.755 8.685 97.040 10.860 ;
        RECT 97.610 8.685 97.850 10.860 ;
        RECT 90.490 8.330 97.850 8.685 ;
        RECT 21.635 7.325 21.925 7.370 ;
        RECT 24.000 7.325 24.320 7.385 ;
        RECT 21.635 7.185 24.320 7.325 ;
        RECT 21.635 7.140 21.925 7.185 ;
        RECT 24.000 7.125 24.320 7.185 ;
        RECT 38.855 7.325 39.145 7.370 ;
        RECT 41.220 7.325 41.540 7.385 ;
        RECT 38.855 7.185 41.540 7.325 ;
        RECT 38.855 7.140 39.145 7.185 ;
        RECT 41.220 7.125 41.540 7.185 ;
        RECT 56.075 7.325 56.365 7.370 ;
        RECT 58.440 7.325 58.760 7.385 ;
        RECT 56.075 7.185 58.760 7.325 ;
        RECT 56.075 7.140 56.365 7.185 ;
        RECT 58.440 7.125 58.760 7.185 ;
        RECT 73.295 7.325 73.585 7.370 ;
        RECT 75.660 7.325 75.980 7.385 ;
        RECT 73.295 7.185 75.980 7.325 ;
        RECT 73.295 7.140 73.585 7.185 ;
        RECT 75.660 7.125 75.980 7.185 ;
        RECT 90.515 7.325 90.805 7.370 ;
        RECT 92.880 7.325 93.200 7.385 ;
        RECT 90.515 7.185 93.200 7.325 ;
        RECT 90.515 7.140 90.805 7.185 ;
        RECT 92.880 7.125 93.200 7.185 ;
      LAYER met2 ;
        RECT 24.020 7.065 24.300 7.435 ;
        RECT 41.240 7.065 41.520 7.435 ;
        RECT 58.460 7.065 58.740 7.435 ;
        RECT 75.680 7.065 75.960 7.435 ;
        RECT 92.900 7.065 93.180 7.435 ;
      LAYER met3 ;
        RECT 23.995 7.400 24.325 7.415 ;
        RECT 41.215 7.400 41.545 7.415 ;
        RECT 58.435 7.400 58.765 7.415 ;
        RECT 75.655 7.400 75.985 7.415 ;
        RECT 92.875 7.400 93.205 7.415 ;
        RECT 23.525 7.100 24.325 7.400 ;
        RECT 40.745 7.100 41.545 7.400 ;
        RECT 57.965 7.100 58.765 7.400 ;
        RECT 75.185 7.100 75.985 7.400 ;
        RECT 92.405 7.100 93.205 7.400 ;
        RECT 23.995 7.085 24.325 7.100 ;
        RECT 41.215 7.085 41.545 7.100 ;
        RECT 58.435 7.085 58.765 7.100 ;
        RECT 75.655 7.085 75.985 7.100 ;
        RECT 92.875 7.085 93.205 7.100 ;
    END
    PORT
      LAYER li1 ;
        RECT 21.755 3.090 21.965 3.910 ;
        RECT 22.635 3.090 22.865 3.910 ;
        RECT 23.085 3.090 23.355 3.900 ;
        RECT 24.025 3.090 24.265 3.900 ;
        RECT 24.475 3.090 24.715 3.900 ;
        RECT 25.385 3.090 25.655 3.900 ;
        RECT 25.835 3.090 26.125 3.925 ;
        RECT 27.665 3.090 27.995 3.480 ;
        RECT 28.505 3.090 28.835 3.480 ;
        RECT 38.975 3.090 39.185 3.910 ;
        RECT 39.855 3.090 40.085 3.910 ;
        RECT 40.305 3.090 40.575 3.900 ;
        RECT 41.245 3.090 41.485 3.900 ;
        RECT 41.695 3.090 41.935 3.900 ;
        RECT 42.605 3.090 42.875 3.900 ;
        RECT 43.055 3.090 43.345 3.925 ;
        RECT 44.885 3.090 45.215 3.480 ;
        RECT 45.725 3.090 46.055 3.480 ;
        RECT 56.195 3.090 56.405 3.910 ;
        RECT 57.075 3.090 57.305 3.910 ;
        RECT 57.525 3.090 57.795 3.900 ;
        RECT 58.465 3.090 58.705 3.900 ;
        RECT 58.915 3.090 59.155 3.900 ;
        RECT 59.825 3.090 60.095 3.900 ;
        RECT 60.275 3.090 60.565 3.925 ;
        RECT 62.105 3.090 62.435 3.480 ;
        RECT 62.945 3.090 63.275 3.480 ;
        RECT 73.415 3.090 73.625 3.910 ;
        RECT 74.295 3.090 74.525 3.910 ;
        RECT 74.745 3.090 75.015 3.900 ;
        RECT 75.685 3.090 75.925 3.900 ;
        RECT 76.135 3.090 76.375 3.900 ;
        RECT 77.045 3.090 77.315 3.900 ;
        RECT 77.495 3.090 77.785 3.925 ;
        RECT 79.325 3.090 79.655 3.480 ;
        RECT 80.165 3.090 80.495 3.480 ;
        RECT 90.635 3.090 90.845 3.910 ;
        RECT 91.515 3.090 91.745 3.910 ;
        RECT 91.965 3.090 92.235 3.900 ;
        RECT 92.905 3.090 93.145 3.900 ;
        RECT 93.355 3.090 93.595 3.900 ;
        RECT 94.265 3.090 94.535 3.900 ;
        RECT 94.715 3.090 95.005 3.925 ;
        RECT 96.545 3.090 96.875 3.480 ;
        RECT 97.385 3.090 97.715 3.480 ;
        RECT 21.605 2.920 29.265 3.090 ;
        RECT 21.605 1.605 21.885 2.920 ;
        RECT 22.170 1.605 22.455 2.920 ;
        RECT 22.740 1.605 23.025 2.920 ;
        RECT 23.310 1.605 23.595 2.920 ;
        RECT 23.880 1.605 24.165 2.920 ;
        RECT 24.450 1.605 24.735 2.920 ;
        RECT 25.020 1.605 25.305 2.920 ;
        RECT 25.590 1.605 25.875 2.920 ;
        RECT 26.160 1.605 26.445 2.920 ;
        RECT 26.730 1.605 27.015 2.920 ;
        RECT 27.300 1.605 27.585 2.920 ;
        RECT 27.870 1.605 28.155 2.920 ;
        RECT 28.440 1.605 28.725 2.920 ;
        RECT 29.010 1.605 29.265 2.920 ;
        RECT 38.825 2.920 46.485 3.090 ;
        RECT 21.605 1.600 29.265 1.605 ;
        RECT 30.335 1.600 30.505 2.225 ;
        RECT 33.080 1.600 33.250 2.225 ;
        RECT 34.065 1.600 34.235 2.225 ;
        RECT 38.825 1.605 39.105 2.920 ;
        RECT 39.390 1.605 39.675 2.920 ;
        RECT 39.960 1.605 40.245 2.920 ;
        RECT 40.530 1.605 40.815 2.920 ;
        RECT 41.100 1.605 41.385 2.920 ;
        RECT 41.670 1.605 41.955 2.920 ;
        RECT 42.240 1.605 42.525 2.920 ;
        RECT 42.810 1.605 43.095 2.920 ;
        RECT 43.380 1.605 43.665 2.920 ;
        RECT 43.950 1.605 44.235 2.920 ;
        RECT 44.520 1.605 44.805 2.920 ;
        RECT 45.090 1.605 45.375 2.920 ;
        RECT 45.660 1.605 45.945 2.920 ;
        RECT 46.230 1.605 46.485 2.920 ;
        RECT 56.045 2.920 63.705 3.090 ;
        RECT 38.825 1.600 46.485 1.605 ;
        RECT 47.555 1.600 47.725 2.225 ;
        RECT 50.300 1.600 50.470 2.225 ;
        RECT 51.285 1.600 51.455 2.225 ;
        RECT 56.045 1.605 56.325 2.920 ;
        RECT 56.610 1.605 56.895 2.920 ;
        RECT 57.180 1.605 57.465 2.920 ;
        RECT 57.750 1.605 58.035 2.920 ;
        RECT 58.320 1.605 58.605 2.920 ;
        RECT 58.890 1.605 59.175 2.920 ;
        RECT 59.460 1.605 59.745 2.920 ;
        RECT 60.030 1.605 60.315 2.920 ;
        RECT 60.600 1.605 60.885 2.920 ;
        RECT 61.170 1.605 61.455 2.920 ;
        RECT 61.740 1.605 62.025 2.920 ;
        RECT 62.310 1.605 62.595 2.920 ;
        RECT 62.880 1.605 63.165 2.920 ;
        RECT 63.450 1.605 63.705 2.920 ;
        RECT 73.265 2.920 80.925 3.090 ;
        RECT 56.045 1.600 63.705 1.605 ;
        RECT 64.775 1.600 64.945 2.225 ;
        RECT 67.520 1.600 67.690 2.225 ;
        RECT 68.505 1.600 68.675 2.225 ;
        RECT 73.265 1.605 73.545 2.920 ;
        RECT 73.830 1.605 74.115 2.920 ;
        RECT 74.400 1.605 74.685 2.920 ;
        RECT 74.970 1.605 75.255 2.920 ;
        RECT 75.540 1.605 75.825 2.920 ;
        RECT 76.110 1.605 76.395 2.920 ;
        RECT 76.680 1.605 76.965 2.920 ;
        RECT 77.250 1.605 77.535 2.920 ;
        RECT 77.820 1.605 78.105 2.920 ;
        RECT 78.390 1.605 78.675 2.920 ;
        RECT 78.960 1.605 79.245 2.920 ;
        RECT 79.530 1.605 79.815 2.920 ;
        RECT 80.100 1.605 80.385 2.920 ;
        RECT 80.670 1.605 80.925 2.920 ;
        RECT 90.485 2.920 98.145 3.090 ;
        RECT 73.265 1.600 80.925 1.605 ;
        RECT 81.995 1.600 82.165 2.225 ;
        RECT 84.740 1.600 84.910 2.225 ;
        RECT 85.725 1.600 85.895 2.225 ;
        RECT 90.485 1.605 90.765 2.920 ;
        RECT 91.050 1.605 91.335 2.920 ;
        RECT 91.620 1.605 91.905 2.920 ;
        RECT 92.190 1.605 92.475 2.920 ;
        RECT 92.760 1.605 93.045 2.920 ;
        RECT 93.330 1.605 93.615 2.920 ;
        RECT 93.900 1.605 94.185 2.920 ;
        RECT 94.470 1.605 94.755 2.920 ;
        RECT 95.040 1.605 95.325 2.920 ;
        RECT 95.610 1.605 95.895 2.920 ;
        RECT 96.180 1.605 96.465 2.920 ;
        RECT 96.750 1.605 97.035 2.920 ;
        RECT 97.320 1.605 97.605 2.920 ;
        RECT 97.890 1.605 98.145 2.920 ;
        RECT 90.485 1.600 98.145 1.605 ;
        RECT 99.215 1.600 99.385 2.225 ;
        RECT 101.960 1.600 102.130 2.225 ;
        RECT 102.945 1.600 103.115 2.225 ;
        RECT 0.015 0.000 103.925 1.600 ;
      LAYER met1 ;
        RECT 21.605 2.765 29.265 3.120 ;
        RECT 21.605 1.605 21.885 2.765 ;
        RECT 22.170 1.605 22.455 2.765 ;
        RECT 22.740 1.605 23.025 2.765 ;
        RECT 23.310 1.605 23.595 2.765 ;
        RECT 23.880 1.605 24.165 2.765 ;
        RECT 24.450 1.605 24.735 2.765 ;
        RECT 25.020 1.605 25.305 2.765 ;
        RECT 25.590 1.605 25.875 2.765 ;
        RECT 26.160 1.605 26.445 2.765 ;
        RECT 26.730 1.605 27.015 2.765 ;
        RECT 27.300 1.605 27.585 2.765 ;
        RECT 27.870 1.605 28.155 2.765 ;
        RECT 28.440 1.605 28.725 2.765 ;
        RECT 29.010 1.605 29.265 2.765 ;
        RECT 21.605 1.600 29.265 1.605 ;
        RECT 38.825 2.765 46.485 3.120 ;
        RECT 38.825 1.605 39.105 2.765 ;
        RECT 39.390 1.605 39.675 2.765 ;
        RECT 39.960 1.605 40.245 2.765 ;
        RECT 40.530 1.605 40.815 2.765 ;
        RECT 41.100 1.605 41.385 2.765 ;
        RECT 41.670 1.605 41.955 2.765 ;
        RECT 42.240 1.605 42.525 2.765 ;
        RECT 42.810 1.605 43.095 2.765 ;
        RECT 43.380 1.605 43.665 2.765 ;
        RECT 43.950 1.605 44.235 2.765 ;
        RECT 44.520 1.605 44.805 2.765 ;
        RECT 45.090 1.605 45.375 2.765 ;
        RECT 45.660 1.605 45.945 2.765 ;
        RECT 46.230 1.605 46.485 2.765 ;
        RECT 38.825 1.600 46.485 1.605 ;
        RECT 56.045 2.765 63.705 3.120 ;
        RECT 56.045 1.605 56.325 2.765 ;
        RECT 56.610 1.605 56.895 2.765 ;
        RECT 57.180 1.605 57.465 2.765 ;
        RECT 57.750 1.605 58.035 2.765 ;
        RECT 58.320 1.605 58.605 2.765 ;
        RECT 58.890 1.605 59.175 2.765 ;
        RECT 59.460 1.605 59.745 2.765 ;
        RECT 60.030 1.605 60.315 2.765 ;
        RECT 60.600 1.605 60.885 2.765 ;
        RECT 61.170 1.605 61.455 2.765 ;
        RECT 61.740 1.605 62.025 2.765 ;
        RECT 62.310 1.605 62.595 2.765 ;
        RECT 62.880 1.605 63.165 2.765 ;
        RECT 63.450 1.605 63.705 2.765 ;
        RECT 56.045 1.600 63.705 1.605 ;
        RECT 73.265 2.765 80.925 3.120 ;
        RECT 73.265 1.605 73.545 2.765 ;
        RECT 73.830 1.605 74.115 2.765 ;
        RECT 74.400 1.605 74.685 2.765 ;
        RECT 74.970 1.605 75.255 2.765 ;
        RECT 75.540 1.605 75.825 2.765 ;
        RECT 76.110 1.605 76.395 2.765 ;
        RECT 76.680 1.605 76.965 2.765 ;
        RECT 77.250 1.605 77.535 2.765 ;
        RECT 77.820 1.605 78.105 2.765 ;
        RECT 78.390 1.605 78.675 2.765 ;
        RECT 78.960 1.605 79.245 2.765 ;
        RECT 79.530 1.605 79.815 2.765 ;
        RECT 80.100 1.605 80.385 2.765 ;
        RECT 80.670 1.605 80.925 2.765 ;
        RECT 73.265 1.600 80.925 1.605 ;
        RECT 90.485 2.765 98.145 3.120 ;
        RECT 90.485 1.605 90.765 2.765 ;
        RECT 91.050 1.605 91.335 2.765 ;
        RECT 91.620 1.605 91.905 2.765 ;
        RECT 92.190 1.605 92.475 2.765 ;
        RECT 92.760 1.605 93.045 2.765 ;
        RECT 93.330 1.605 93.615 2.765 ;
        RECT 93.900 1.605 94.185 2.765 ;
        RECT 94.470 1.605 94.755 2.765 ;
        RECT 95.040 1.605 95.325 2.765 ;
        RECT 95.610 1.605 95.895 2.765 ;
        RECT 96.180 1.605 96.465 2.765 ;
        RECT 96.750 1.605 97.035 2.765 ;
        RECT 97.320 1.605 97.605 2.765 ;
        RECT 97.890 1.605 98.145 2.765 ;
        RECT 90.485 1.600 98.145 1.605 ;
        RECT 0.015 0.000 103.925 1.600 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 15.015 8.745 16.010 9.015 ;
        RECT 15.015 8.740 18.495 8.745 ;
        RECT 30.115 8.740 35.680 8.745 ;
        RECT 47.335 8.740 53.030 8.745 ;
        RECT 64.555 8.740 70.105 8.745 ;
        RECT 81.775 8.740 87.320 8.745 ;
        RECT 98.995 8.740 103.775 8.745 ;
        RECT 15.015 7.145 21.410 8.740 ;
        RECT 29.350 8.130 38.465 8.740 ;
        RECT 46.570 8.130 55.685 8.740 ;
        RECT 63.790 8.130 72.905 8.740 ;
        RECT 81.010 8.130 90.125 8.740 ;
        RECT 98.230 8.130 103.925 8.740 ;
        RECT 29.155 7.145 38.465 8.130 ;
        RECT 46.375 7.145 55.685 8.130 ;
        RECT 63.595 7.145 72.905 8.130 ;
        RECT 80.815 7.145 90.125 8.130 ;
        RECT 15.015 7.140 21.455 7.145 ;
        RECT 29.155 7.140 38.675 7.145 ;
        RECT 46.375 7.140 55.895 7.145 ;
        RECT 63.595 7.140 73.115 7.145 ;
        RECT 80.815 7.140 90.335 7.145 ;
        RECT 98.035 7.140 103.925 8.130 ;
        RECT 15.015 4.310 103.925 7.140 ;
        RECT 15.015 3.710 21.410 4.310 ;
        RECT 29.350 3.720 38.630 4.310 ;
        RECT 46.570 3.720 55.850 4.310 ;
        RECT 63.790 3.720 73.070 4.310 ;
        RECT 81.010 3.720 90.290 4.310 ;
        RECT 98.230 3.720 103.925 4.310 ;
        RECT 30.115 3.715 38.630 3.720 ;
        RECT 47.335 3.715 55.850 3.720 ;
        RECT 64.555 3.715 73.070 3.720 ;
        RECT 81.775 3.715 90.290 3.720 ;
        RECT 98.995 3.715 103.770 3.720 ;
        RECT 35.035 3.710 38.630 3.715 ;
        RECT 52.255 3.710 55.850 3.715 ;
        RECT 69.475 3.710 73.070 3.715 ;
        RECT 86.695 3.710 90.290 3.715 ;
      LAYER li1 ;
        RECT 17.055 10.045 17.230 10.595 ;
        RECT 17.055 8.445 17.225 10.045 ;
        RECT 15.240 7.035 15.410 7.765 ;
        RECT 17.055 7.305 17.230 8.445 ;
        RECT 17.055 7.035 17.225 7.305 ;
        RECT 15.070 7.030 17.820 7.035 ;
        RECT 18.650 7.030 18.820 7.755 ;
        RECT 30.335 7.035 30.505 7.765 ;
        RECT 33.080 7.035 33.250 7.765 ;
        RECT 34.070 7.035 34.240 7.765 ;
        RECT 30.165 7.030 34.890 7.035 ;
        RECT 35.870 7.030 36.040 7.755 ;
        RECT 47.555 7.035 47.725 7.765 ;
        RECT 50.300 7.035 50.470 7.765 ;
        RECT 51.290 7.035 51.460 7.765 ;
        RECT 47.385 7.030 52.110 7.035 ;
        RECT 53.090 7.030 53.260 7.755 ;
        RECT 64.775 7.035 64.945 7.765 ;
        RECT 67.520 7.035 67.690 7.765 ;
        RECT 68.510 7.035 68.680 7.765 ;
        RECT 64.605 7.030 69.330 7.035 ;
        RECT 70.310 7.030 70.480 7.755 ;
        RECT 81.995 7.035 82.165 7.765 ;
        RECT 84.740 7.035 84.910 7.765 ;
        RECT 85.730 7.035 85.900 7.765 ;
        RECT 81.825 7.030 86.550 7.035 ;
        RECT 87.530 7.030 87.700 7.755 ;
        RECT 99.215 7.035 99.385 7.765 ;
        RECT 101.960 7.035 102.130 7.765 ;
        RECT 102.950 7.035 103.120 7.765 ;
        RECT 99.045 7.030 103.770 7.035 ;
        RECT 15.070 7.025 21.495 7.030 ;
        RECT 0.015 7.000 21.500 7.025 ;
        RECT 28.960 7.000 38.715 7.030 ;
        RECT 46.180 7.000 55.935 7.030 ;
        RECT 63.400 7.000 73.155 7.030 ;
        RECT 80.620 7.000 90.375 7.030 ;
        RECT 0.015 5.810 21.625 7.000 ;
        RECT 22.155 5.810 22.435 6.950 ;
        RECT 23.105 5.810 23.365 6.950 ;
        RECT 24.455 5.810 24.735 6.950 ;
        RECT 25.405 5.810 25.665 6.950 ;
        RECT 25.835 5.810 26.095 6.950 ;
        RECT 26.765 5.810 27.045 6.950 ;
        RECT 27.215 5.810 27.475 6.950 ;
        RECT 28.145 5.810 28.425 6.950 ;
        RECT 28.960 5.810 38.845 7.000 ;
        RECT 39.375 5.810 39.655 6.950 ;
        RECT 40.325 5.810 40.585 6.950 ;
        RECT 41.675 5.810 41.955 6.950 ;
        RECT 42.625 5.810 42.885 6.950 ;
        RECT 43.055 5.810 43.315 6.950 ;
        RECT 43.985 5.810 44.265 6.950 ;
        RECT 44.435 5.810 44.695 6.950 ;
        RECT 45.365 5.810 45.645 6.950 ;
        RECT 46.180 5.810 56.065 7.000 ;
        RECT 56.595 5.810 56.875 6.950 ;
        RECT 57.545 5.810 57.805 6.950 ;
        RECT 58.895 5.810 59.175 6.950 ;
        RECT 59.845 5.810 60.105 6.950 ;
        RECT 60.275 5.810 60.535 6.950 ;
        RECT 61.205 5.810 61.485 6.950 ;
        RECT 61.655 5.810 61.915 6.950 ;
        RECT 62.585 5.810 62.865 6.950 ;
        RECT 63.400 5.810 73.285 7.000 ;
        RECT 73.815 5.810 74.095 6.950 ;
        RECT 74.765 5.810 75.025 6.950 ;
        RECT 76.115 5.810 76.395 6.950 ;
        RECT 77.065 5.810 77.325 6.950 ;
        RECT 77.495 5.810 77.755 6.950 ;
        RECT 78.425 5.810 78.705 6.950 ;
        RECT 78.875 5.810 79.135 6.950 ;
        RECT 79.805 5.810 80.085 6.950 ;
        RECT 80.620 5.810 90.505 7.000 ;
        RECT 91.035 5.810 91.315 6.950 ;
        RECT 91.985 5.810 92.245 6.950 ;
        RECT 93.335 5.810 93.615 6.950 ;
        RECT 94.285 5.810 94.545 6.950 ;
        RECT 94.715 5.810 94.975 6.950 ;
        RECT 95.645 5.810 95.925 6.950 ;
        RECT 96.095 5.810 96.355 6.950 ;
        RECT 97.025 5.810 97.305 6.950 ;
        RECT 97.840 5.810 103.925 7.030 ;
        RECT 0.015 5.640 103.925 5.810 ;
        RECT 0.015 5.425 21.965 5.640 ;
        RECT 21.755 4.500 21.965 5.425 ;
        RECT 22.635 4.500 22.865 5.640 ;
        RECT 23.085 4.500 23.415 5.640 ;
        RECT 25.325 4.500 25.655 5.640 ;
        RECT 26.905 5.130 27.075 5.640 ;
        RECT 27.745 4.790 27.915 5.640 ;
        RECT 29.055 5.430 39.185 5.640 ;
        RECT 30.165 5.425 39.185 5.430 ;
        RECT 30.335 4.695 30.505 5.425 ;
        RECT 33.080 4.695 33.250 5.425 ;
        RECT 34.065 4.695 34.235 5.425 ;
        RECT 38.975 4.500 39.185 5.425 ;
        RECT 39.855 4.500 40.085 5.640 ;
        RECT 40.305 4.500 40.635 5.640 ;
        RECT 42.545 4.500 42.875 5.640 ;
        RECT 44.125 5.130 44.295 5.640 ;
        RECT 44.965 4.790 45.135 5.640 ;
        RECT 46.275 5.430 56.405 5.640 ;
        RECT 47.385 5.425 56.405 5.430 ;
        RECT 47.555 4.695 47.725 5.425 ;
        RECT 50.300 4.695 50.470 5.425 ;
        RECT 51.285 4.695 51.455 5.425 ;
        RECT 56.195 4.500 56.405 5.425 ;
        RECT 57.075 4.500 57.305 5.640 ;
        RECT 57.525 4.500 57.855 5.640 ;
        RECT 59.765 4.500 60.095 5.640 ;
        RECT 61.345 5.130 61.515 5.640 ;
        RECT 62.185 4.790 62.355 5.640 ;
        RECT 63.495 5.430 73.625 5.640 ;
        RECT 64.605 5.425 73.625 5.430 ;
        RECT 64.775 4.695 64.945 5.425 ;
        RECT 67.520 4.695 67.690 5.425 ;
        RECT 68.505 4.695 68.675 5.425 ;
        RECT 73.415 4.500 73.625 5.425 ;
        RECT 74.295 4.500 74.525 5.640 ;
        RECT 74.745 4.500 75.075 5.640 ;
        RECT 76.985 4.500 77.315 5.640 ;
        RECT 78.565 5.130 78.735 5.640 ;
        RECT 79.405 4.790 79.575 5.640 ;
        RECT 80.715 5.430 90.845 5.640 ;
        RECT 81.825 5.425 90.845 5.430 ;
        RECT 81.995 4.695 82.165 5.425 ;
        RECT 84.740 4.695 84.910 5.425 ;
        RECT 85.725 4.695 85.895 5.425 ;
        RECT 90.635 4.500 90.845 5.425 ;
        RECT 91.515 4.500 91.745 5.640 ;
        RECT 91.965 4.500 92.295 5.640 ;
        RECT 94.205 4.500 94.535 5.640 ;
        RECT 95.785 5.130 95.955 5.640 ;
        RECT 96.625 4.790 96.795 5.640 ;
        RECT 97.935 5.430 103.925 5.640 ;
        RECT 99.045 5.425 103.765 5.430 ;
        RECT 99.215 4.695 99.385 5.425 ;
        RECT 101.960 4.695 102.130 5.425 ;
        RECT 102.945 4.695 103.115 5.425 ;
      LAYER met1 ;
        RECT 16.995 9.145 17.285 9.175 ;
        RECT 16.825 8.975 17.285 9.145 ;
        RECT 16.995 8.945 17.285 8.975 ;
        RECT 15.070 7.030 17.820 7.035 ;
        RECT 30.165 7.030 34.890 7.035 ;
        RECT 47.385 7.030 52.110 7.035 ;
        RECT 64.605 7.030 69.330 7.035 ;
        RECT 81.825 7.030 86.550 7.035 ;
        RECT 99.045 7.030 103.770 7.035 ;
        RECT 15.070 7.025 21.495 7.030 ;
        RECT 0.015 7.000 21.500 7.025 ;
        RECT 28.960 7.000 38.715 7.030 ;
        RECT 46.180 7.000 55.935 7.030 ;
        RECT 63.400 7.000 73.155 7.030 ;
        RECT 80.620 7.000 90.375 7.030 ;
        RECT 0.015 5.965 21.625 7.000 ;
        RECT 28.960 5.965 38.845 7.000 ;
        RECT 46.180 5.965 56.065 7.000 ;
        RECT 63.400 5.965 73.285 7.000 ;
        RECT 80.620 5.965 90.505 7.000 ;
        RECT 97.840 5.965 103.925 7.030 ;
        RECT 0.015 5.485 103.925 5.965 ;
        RECT 0.015 5.425 21.785 5.485 ;
        RECT 29.055 5.430 39.005 5.485 ;
        RECT 46.275 5.430 56.225 5.485 ;
        RECT 63.495 5.430 73.445 5.485 ;
        RECT 80.715 5.430 90.665 5.485 ;
        RECT 97.935 5.430 103.925 5.485 ;
        RECT 30.165 5.425 39.005 5.430 ;
        RECT 47.385 5.425 56.225 5.430 ;
        RECT 64.605 5.425 73.445 5.430 ;
        RECT 81.825 5.425 90.665 5.430 ;
        RECT 99.045 5.425 103.765 5.430 ;
    END
  END vccd1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 18.660 8.225 18.830 9.495 ;
        RECT 30.345 8.465 30.515 9.505 ;
        RECT 30.340 8.225 30.520 8.465 ;
        RECT 30.345 2.955 30.515 4.225 ;
      LAYER met1 ;
        RECT 18.565 8.400 18.905 8.495 ;
        RECT 18.565 8.395 18.920 8.400 ;
        RECT 18.565 8.365 19.060 8.395 ;
        RECT 20.885 8.365 21.225 8.455 ;
        RECT 18.565 8.200 21.225 8.365 ;
        RECT 18.565 8.155 18.905 8.200 ;
        RECT 20.885 8.175 21.225 8.200 ;
        RECT 30.270 8.405 30.595 8.465 ;
        RECT 30.270 8.235 30.745 8.405 ;
        RECT 30.270 8.140 30.595 8.235 ;
        RECT 30.270 4.790 30.595 5.115 ;
        RECT 30.350 4.255 30.520 4.790 ;
        RECT 30.285 4.225 30.575 4.255 ;
        RECT 30.285 4.055 30.745 4.225 ;
        RECT 30.285 4.025 30.575 4.055 ;
      LAYER met2 ;
        RECT 20.970 9.320 30.520 9.490 ;
        RECT 18.545 8.140 18.920 8.510 ;
        RECT 20.970 8.485 21.140 9.320 ;
        RECT 20.915 8.145 21.195 8.485 ;
        RECT 30.350 8.465 30.520 9.320 ;
        RECT 30.270 8.140 30.595 8.465 ;
        RECT 30.340 5.115 30.510 8.140 ;
        RECT 30.270 4.790 30.595 5.115 ;
      LAYER met3 ;
        RECT 18.570 8.510 18.900 12.445 ;
        RECT 18.545 8.140 18.920 8.510 ;
    END
  END s1
  OBS
      LAYER pwell ;
        RECT 21.485 8.530 22.085 8.745 ;
        RECT 38.705 8.530 39.305 8.745 ;
        RECT 55.925 8.530 56.525 8.745 ;
        RECT 73.145 8.530 73.745 8.745 ;
        RECT 90.365 8.530 90.965 8.745 ;
        RECT 21.485 8.340 22.380 8.530 ;
        RECT 24.510 8.495 24.680 8.530 ;
        RECT 23.605 8.385 24.680 8.495 ;
        RECT 24.395 8.340 24.680 8.385 ;
        RECT 26.820 8.340 26.990 8.530 ;
        RECT 28.200 8.500 28.370 8.530 ;
        RECT 28.200 8.390 28.770 8.500 ;
        RECT 28.200 8.340 28.485 8.390 ;
        RECT 21.485 8.145 23.445 8.340 ;
        RECT 22.095 7.430 23.445 8.145 ;
        RECT 24.395 7.430 28.485 8.340 ;
        RECT 38.705 8.340 39.600 8.530 ;
        RECT 41.730 8.495 41.900 8.530 ;
        RECT 40.825 8.385 41.900 8.495 ;
        RECT 41.615 8.340 41.900 8.385 ;
        RECT 44.040 8.340 44.210 8.530 ;
        RECT 45.420 8.500 45.590 8.530 ;
        RECT 45.420 8.390 45.990 8.500 ;
        RECT 45.420 8.340 45.705 8.390 ;
        RECT 38.705 8.145 40.665 8.340 ;
        RECT 39.315 7.430 40.665 8.145 ;
        RECT 41.615 7.430 45.705 8.340 ;
        RECT 55.925 8.340 56.820 8.530 ;
        RECT 58.950 8.495 59.120 8.530 ;
        RECT 58.045 8.385 59.120 8.495 ;
        RECT 58.835 8.340 59.120 8.385 ;
        RECT 61.260 8.340 61.430 8.530 ;
        RECT 62.640 8.500 62.810 8.530 ;
        RECT 62.640 8.390 63.210 8.500 ;
        RECT 62.640 8.340 62.925 8.390 ;
        RECT 55.925 8.145 57.885 8.340 ;
        RECT 56.535 7.430 57.885 8.145 ;
        RECT 58.835 7.430 62.925 8.340 ;
        RECT 73.145 8.340 74.040 8.530 ;
        RECT 76.170 8.495 76.340 8.530 ;
        RECT 75.265 8.385 76.340 8.495 ;
        RECT 76.055 8.340 76.340 8.385 ;
        RECT 78.480 8.340 78.650 8.530 ;
        RECT 79.860 8.500 80.030 8.530 ;
        RECT 79.860 8.390 80.430 8.500 ;
        RECT 79.860 8.340 80.145 8.390 ;
        RECT 73.145 8.145 75.105 8.340 ;
        RECT 73.755 7.430 75.105 8.145 ;
        RECT 76.055 7.430 80.145 8.340 ;
        RECT 90.365 8.340 91.260 8.530 ;
        RECT 93.390 8.495 93.560 8.530 ;
        RECT 92.485 8.385 93.560 8.495 ;
        RECT 93.275 8.340 93.560 8.385 ;
        RECT 95.700 8.340 95.870 8.530 ;
        RECT 97.080 8.500 97.250 8.530 ;
        RECT 97.080 8.390 97.650 8.500 ;
        RECT 97.080 8.340 97.365 8.390 ;
        RECT 90.365 8.145 92.325 8.340 ;
        RECT 90.975 7.430 92.325 8.145 ;
        RECT 93.275 7.430 97.365 8.340 ;
        RECT 21.625 3.305 28.925 4.020 ;
        RECT 38.845 3.305 46.145 4.020 ;
        RECT 56.065 3.305 63.365 4.020 ;
        RECT 73.285 3.305 80.585 4.020 ;
        RECT 90.505 3.305 97.805 4.020 ;
        RECT 21.485 3.110 28.925 3.305 ;
        RECT 38.705 3.110 46.145 3.305 ;
        RECT 55.925 3.110 63.365 3.305 ;
        RECT 73.145 3.110 80.585 3.305 ;
        RECT 90.365 3.110 97.805 3.305 ;
        RECT 21.485 2.920 22.845 3.110 ;
        RECT 24.050 2.920 24.690 3.110 ;
        RECT 28.655 2.920 28.825 3.110 ;
        RECT 38.705 2.920 40.065 3.110 ;
        RECT 41.270 2.920 41.910 3.110 ;
        RECT 45.875 2.920 46.045 3.110 ;
        RECT 55.925 2.920 57.285 3.110 ;
        RECT 58.490 2.920 59.130 3.110 ;
        RECT 63.095 2.920 63.265 3.110 ;
        RECT 73.145 2.920 74.505 3.110 ;
        RECT 75.710 2.920 76.350 3.110 ;
        RECT 80.315 2.920 80.485 3.110 ;
        RECT 90.365 2.920 91.725 3.110 ;
        RECT 92.930 2.920 93.570 3.110 ;
        RECT 97.535 2.920 97.705 3.110 ;
        RECT 21.485 2.705 22.085 2.920 ;
        RECT 38.705 2.705 39.305 2.920 ;
        RECT 55.925 2.705 56.525 2.920 ;
        RECT 73.145 2.705 73.745 2.920 ;
        RECT 90.365 2.705 90.965 2.920 ;
      LAYER li1 ;
        RECT 15.670 10.105 15.845 10.595 ;
        RECT 16.195 10.315 16.365 10.595 ;
        RECT 16.195 10.145 16.425 10.315 ;
        RECT 15.670 9.935 15.840 10.105 ;
        RECT 15.670 9.605 16.080 9.935 ;
        RECT 15.670 9.095 15.840 9.605 ;
        RECT 15.670 8.765 16.080 9.095 ;
        RECT 15.670 8.565 15.840 8.765 ;
        RECT 15.670 7.305 15.845 8.565 ;
        RECT 16.255 8.535 16.425 10.145 ;
        RECT 16.625 10.085 16.800 10.595 ;
        RECT 19.080 10.095 19.255 10.585 ;
        RECT 19.080 9.925 19.250 10.095 ;
        RECT 20.035 10.075 20.210 10.585 ;
        RECT 20.465 10.035 20.640 10.585 ;
        RECT 30.765 10.105 30.940 10.595 ;
        RECT 31.290 10.315 31.460 10.595 ;
        RECT 31.290 10.145 31.520 10.315 ;
        RECT 19.080 9.595 19.490 9.925 ;
        RECT 16.195 8.365 16.425 8.535 ;
        RECT 16.625 8.565 16.795 9.515 ;
        RECT 19.080 9.085 19.250 9.595 ;
        RECT 19.080 8.755 19.490 9.085 ;
        RECT 16.195 7.305 16.365 8.365 ;
        RECT 16.625 7.305 16.800 8.565 ;
        RECT 19.080 8.555 19.250 8.755 ;
        RECT 20.035 8.555 20.205 9.505 ;
        RECT 19.080 7.295 19.255 8.555 ;
        RECT 20.035 7.295 20.210 8.555 ;
        RECT 20.465 8.435 20.635 10.035 ;
        RECT 30.765 9.935 30.935 10.105 ;
        RECT 30.765 9.605 31.175 9.935 ;
        RECT 30.765 9.095 30.935 9.605 ;
        RECT 30.765 8.765 31.175 9.095 ;
        RECT 30.765 8.565 30.935 8.765 ;
        RECT 20.465 7.295 20.640 8.435 ;
        RECT 22.670 7.560 23.365 8.190 ;
        RECT 22.670 6.960 22.840 7.560 ;
        RECT 23.010 7.340 23.345 7.370 ;
        RECT 23.735 7.340 23.905 8.020 ;
        RECT 23.010 7.170 23.905 7.340 ;
        RECT 24.970 7.560 25.665 8.190 ;
        RECT 25.835 7.560 26.530 8.190 ;
        RECT 27.215 7.560 27.910 8.190 ;
        RECT 23.010 7.120 23.345 7.170 ;
        RECT 24.970 6.960 25.140 7.560 ;
        RECT 25.310 7.340 25.645 7.370 ;
        RECT 25.855 7.340 26.190 7.370 ;
        RECT 25.310 7.170 26.190 7.340 ;
        RECT 25.310 7.120 25.645 7.170 ;
        RECT 25.855 7.120 26.190 7.170 ;
        RECT 26.360 6.960 26.530 7.560 ;
        RECT 26.700 7.120 27.035 7.390 ;
        RECT 27.235 7.120 27.570 7.370 ;
        RECT 27.740 6.960 27.910 7.560 ;
        RECT 28.080 7.120 28.415 7.390 ;
        RECT 30.765 7.305 30.940 8.565 ;
        RECT 31.350 8.535 31.520 10.145 ;
        RECT 31.720 10.085 31.895 10.595 ;
        RECT 32.150 10.045 32.325 10.595 ;
        RECT 33.515 10.085 33.685 10.595 ;
        RECT 34.505 10.085 34.675 10.595 ;
        RECT 36.300 10.095 36.475 10.585 ;
        RECT 31.290 8.365 31.520 8.535 ;
        RECT 31.720 8.565 31.890 9.515 ;
        RECT 31.290 7.305 31.460 8.365 ;
        RECT 31.720 7.305 31.895 8.565 ;
        RECT 32.150 8.445 32.320 10.045 ;
        RECT 36.300 9.925 36.470 10.095 ;
        RECT 37.255 10.075 37.430 10.585 ;
        RECT 37.685 10.035 37.860 10.585 ;
        RECT 47.985 10.105 48.160 10.595 ;
        RECT 48.510 10.315 48.680 10.595 ;
        RECT 48.510 10.145 48.740 10.315 ;
        RECT 33.080 9.425 33.310 9.610 ;
        RECT 36.300 9.595 36.710 9.925 ;
        RECT 33.080 9.380 33.610 9.425 ;
        RECT 33.140 9.255 33.610 9.380 ;
        RECT 34.130 9.255 34.600 9.425 ;
        RECT 33.140 8.565 33.310 9.255 ;
        RECT 33.510 8.780 33.680 8.885 ;
        RECT 34.130 8.780 34.300 9.255 ;
        RECT 36.300 9.085 36.470 9.595 ;
        RECT 33.510 8.605 34.300 8.780 ;
        RECT 32.150 7.305 32.325 8.445 ;
        RECT 33.510 7.305 33.685 8.605 ;
        RECT 34.130 8.565 34.300 8.605 ;
        RECT 34.500 8.450 34.670 8.885 ;
        RECT 36.300 8.755 36.710 9.085 ;
        RECT 36.300 8.555 36.470 8.755 ;
        RECT 37.255 8.555 37.425 9.505 ;
        RECT 34.500 7.305 34.675 8.450 ;
        RECT 36.300 7.295 36.475 8.555 ;
        RECT 37.255 7.295 37.430 8.555 ;
        RECT 37.685 8.435 37.855 10.035 ;
        RECT 47.985 9.935 48.155 10.105 ;
        RECT 47.985 9.605 48.395 9.935 ;
        RECT 47.985 9.095 48.155 9.605 ;
        RECT 47.985 8.765 48.395 9.095 ;
        RECT 47.985 8.565 48.155 8.765 ;
        RECT 37.685 7.295 37.860 8.435 ;
        RECT 39.890 7.560 40.585 8.190 ;
        RECT 39.890 6.960 40.060 7.560 ;
        RECT 40.230 7.340 40.565 7.370 ;
        RECT 40.955 7.340 41.125 8.020 ;
        RECT 40.230 7.170 41.125 7.340 ;
        RECT 42.190 7.560 42.885 8.190 ;
        RECT 43.055 7.560 43.750 8.190 ;
        RECT 44.435 7.560 45.130 8.190 ;
        RECT 40.230 7.120 40.565 7.170 ;
        RECT 42.190 6.960 42.360 7.560 ;
        RECT 42.530 7.340 42.865 7.370 ;
        RECT 43.075 7.340 43.410 7.370 ;
        RECT 42.530 7.170 43.410 7.340 ;
        RECT 42.530 7.120 42.865 7.170 ;
        RECT 43.075 7.120 43.410 7.170 ;
        RECT 43.580 6.960 43.750 7.560 ;
        RECT 43.920 7.120 44.255 7.390 ;
        RECT 44.455 7.120 44.790 7.370 ;
        RECT 44.960 6.960 45.130 7.560 ;
        RECT 45.300 7.120 45.635 7.390 ;
        RECT 47.985 7.305 48.160 8.565 ;
        RECT 48.570 8.535 48.740 10.145 ;
        RECT 48.940 10.085 49.115 10.595 ;
        RECT 49.370 10.045 49.545 10.595 ;
        RECT 50.735 10.085 50.905 10.595 ;
        RECT 51.725 10.085 51.895 10.595 ;
        RECT 53.520 10.095 53.695 10.585 ;
        RECT 48.510 8.365 48.740 8.535 ;
        RECT 48.940 8.565 49.110 9.515 ;
        RECT 48.510 7.305 48.680 8.365 ;
        RECT 48.940 7.305 49.115 8.565 ;
        RECT 49.370 8.445 49.540 10.045 ;
        RECT 53.520 9.925 53.690 10.095 ;
        RECT 54.475 10.075 54.650 10.585 ;
        RECT 54.905 10.035 55.080 10.585 ;
        RECT 65.205 10.105 65.380 10.595 ;
        RECT 65.730 10.315 65.900 10.595 ;
        RECT 65.730 10.145 65.960 10.315 ;
        RECT 50.300 9.425 50.530 9.610 ;
        RECT 53.520 9.595 53.930 9.925 ;
        RECT 50.300 9.380 50.830 9.425 ;
        RECT 50.360 9.255 50.830 9.380 ;
        RECT 51.350 9.255 51.820 9.425 ;
        RECT 50.360 8.565 50.530 9.255 ;
        RECT 50.730 8.780 50.900 8.885 ;
        RECT 51.350 8.780 51.520 9.255 ;
        RECT 53.520 9.085 53.690 9.595 ;
        RECT 50.730 8.605 51.520 8.780 ;
        RECT 49.370 7.305 49.545 8.445 ;
        RECT 50.730 7.305 50.905 8.605 ;
        RECT 51.350 8.565 51.520 8.605 ;
        RECT 51.720 8.450 51.890 8.885 ;
        RECT 53.520 8.755 53.930 9.085 ;
        RECT 53.520 8.555 53.690 8.755 ;
        RECT 54.475 8.555 54.645 9.505 ;
        RECT 51.720 7.305 51.895 8.450 ;
        RECT 53.520 7.295 53.695 8.555 ;
        RECT 54.475 7.295 54.650 8.555 ;
        RECT 54.905 8.435 55.075 10.035 ;
        RECT 65.205 9.935 65.375 10.105 ;
        RECT 65.205 9.605 65.615 9.935 ;
        RECT 65.205 9.095 65.375 9.605 ;
        RECT 65.205 8.765 65.615 9.095 ;
        RECT 65.205 8.565 65.375 8.765 ;
        RECT 54.905 7.295 55.080 8.435 ;
        RECT 57.110 7.560 57.805 8.190 ;
        RECT 57.110 6.960 57.280 7.560 ;
        RECT 57.450 7.340 57.785 7.370 ;
        RECT 58.175 7.340 58.345 8.020 ;
        RECT 57.450 7.170 58.345 7.340 ;
        RECT 59.410 7.560 60.105 8.190 ;
        RECT 60.275 7.560 60.970 8.190 ;
        RECT 61.655 7.560 62.350 8.190 ;
        RECT 57.450 7.120 57.785 7.170 ;
        RECT 59.410 6.960 59.580 7.560 ;
        RECT 59.750 7.340 60.085 7.370 ;
        RECT 60.295 7.340 60.630 7.370 ;
        RECT 59.750 7.170 60.630 7.340 ;
        RECT 59.750 7.120 60.085 7.170 ;
        RECT 60.295 7.120 60.630 7.170 ;
        RECT 60.800 6.960 60.970 7.560 ;
        RECT 61.140 7.120 61.475 7.390 ;
        RECT 61.675 7.120 62.010 7.370 ;
        RECT 62.180 6.960 62.350 7.560 ;
        RECT 62.520 7.120 62.855 7.390 ;
        RECT 65.205 7.305 65.380 8.565 ;
        RECT 65.790 8.535 65.960 10.145 ;
        RECT 66.160 10.085 66.335 10.595 ;
        RECT 66.590 10.045 66.765 10.595 ;
        RECT 67.955 10.085 68.125 10.595 ;
        RECT 68.945 10.085 69.115 10.595 ;
        RECT 70.740 10.095 70.915 10.585 ;
        RECT 65.730 8.365 65.960 8.535 ;
        RECT 66.160 8.565 66.330 9.515 ;
        RECT 65.730 7.305 65.900 8.365 ;
        RECT 66.160 7.305 66.335 8.565 ;
        RECT 66.590 8.445 66.760 10.045 ;
        RECT 70.740 9.925 70.910 10.095 ;
        RECT 71.695 10.075 71.870 10.585 ;
        RECT 72.125 10.035 72.300 10.585 ;
        RECT 82.425 10.105 82.600 10.595 ;
        RECT 82.950 10.315 83.120 10.595 ;
        RECT 82.950 10.145 83.180 10.315 ;
        RECT 67.520 9.425 67.750 9.610 ;
        RECT 70.740 9.595 71.150 9.925 ;
        RECT 67.520 9.380 68.050 9.425 ;
        RECT 67.580 9.255 68.050 9.380 ;
        RECT 68.570 9.255 69.040 9.425 ;
        RECT 67.580 8.565 67.750 9.255 ;
        RECT 67.950 8.780 68.120 8.885 ;
        RECT 68.570 8.780 68.740 9.255 ;
        RECT 70.740 9.085 70.910 9.595 ;
        RECT 67.950 8.605 68.740 8.780 ;
        RECT 66.590 7.305 66.765 8.445 ;
        RECT 67.950 7.305 68.125 8.605 ;
        RECT 68.570 8.565 68.740 8.605 ;
        RECT 68.940 8.450 69.110 8.885 ;
        RECT 70.740 8.755 71.150 9.085 ;
        RECT 70.740 8.555 70.910 8.755 ;
        RECT 71.695 8.555 71.865 9.505 ;
        RECT 68.940 7.305 69.115 8.450 ;
        RECT 70.740 7.295 70.915 8.555 ;
        RECT 71.695 7.295 71.870 8.555 ;
        RECT 72.125 8.435 72.295 10.035 ;
        RECT 82.425 9.935 82.595 10.105 ;
        RECT 82.425 9.605 82.835 9.935 ;
        RECT 82.425 9.095 82.595 9.605 ;
        RECT 82.425 8.765 82.835 9.095 ;
        RECT 82.425 8.565 82.595 8.765 ;
        RECT 72.125 7.295 72.300 8.435 ;
        RECT 74.330 7.560 75.025 8.190 ;
        RECT 74.330 6.960 74.500 7.560 ;
        RECT 74.670 7.340 75.005 7.370 ;
        RECT 75.395 7.340 75.565 8.020 ;
        RECT 74.670 7.170 75.565 7.340 ;
        RECT 76.630 7.560 77.325 8.190 ;
        RECT 77.495 7.560 78.190 8.190 ;
        RECT 78.875 7.560 79.570 8.190 ;
        RECT 74.670 7.120 75.005 7.170 ;
        RECT 76.630 6.960 76.800 7.560 ;
        RECT 76.970 7.340 77.305 7.370 ;
        RECT 77.515 7.340 77.850 7.370 ;
        RECT 76.970 7.170 77.850 7.340 ;
        RECT 76.970 7.120 77.305 7.170 ;
        RECT 77.515 7.120 77.850 7.170 ;
        RECT 78.020 6.960 78.190 7.560 ;
        RECT 78.360 7.120 78.695 7.390 ;
        RECT 78.895 7.120 79.230 7.370 ;
        RECT 79.400 6.960 79.570 7.560 ;
        RECT 79.740 7.120 80.075 7.390 ;
        RECT 82.425 7.305 82.600 8.565 ;
        RECT 83.010 8.535 83.180 10.145 ;
        RECT 83.380 10.085 83.555 10.595 ;
        RECT 83.810 10.045 83.985 10.595 ;
        RECT 85.175 10.085 85.345 10.595 ;
        RECT 86.165 10.085 86.335 10.595 ;
        RECT 87.960 10.095 88.135 10.585 ;
        RECT 82.950 8.365 83.180 8.535 ;
        RECT 83.380 8.565 83.550 9.515 ;
        RECT 82.950 7.305 83.120 8.365 ;
        RECT 83.380 7.305 83.555 8.565 ;
        RECT 83.810 8.445 83.980 10.045 ;
        RECT 87.960 9.925 88.130 10.095 ;
        RECT 88.915 10.075 89.090 10.585 ;
        RECT 89.345 10.035 89.520 10.585 ;
        RECT 99.645 10.105 99.820 10.595 ;
        RECT 100.170 10.315 100.340 10.595 ;
        RECT 100.170 10.145 100.400 10.315 ;
        RECT 84.740 9.425 84.970 9.610 ;
        RECT 87.960 9.595 88.370 9.925 ;
        RECT 84.740 9.380 85.270 9.425 ;
        RECT 84.800 9.255 85.270 9.380 ;
        RECT 85.790 9.255 86.260 9.425 ;
        RECT 84.800 8.565 84.970 9.255 ;
        RECT 85.170 8.780 85.340 8.885 ;
        RECT 85.790 8.780 85.960 9.255 ;
        RECT 87.960 9.085 88.130 9.595 ;
        RECT 85.170 8.605 85.960 8.780 ;
        RECT 83.810 7.305 83.985 8.445 ;
        RECT 85.170 7.305 85.345 8.605 ;
        RECT 85.790 8.565 85.960 8.605 ;
        RECT 86.160 8.450 86.330 8.885 ;
        RECT 87.960 8.755 88.370 9.085 ;
        RECT 87.960 8.555 88.130 8.755 ;
        RECT 88.915 8.555 89.085 9.505 ;
        RECT 86.160 7.305 86.335 8.450 ;
        RECT 87.960 7.295 88.135 8.555 ;
        RECT 88.915 7.295 89.090 8.555 ;
        RECT 89.345 8.435 89.515 10.035 ;
        RECT 99.645 9.935 99.815 10.105 ;
        RECT 99.645 9.605 100.055 9.935 ;
        RECT 99.645 9.095 99.815 9.605 ;
        RECT 99.645 8.765 100.055 9.095 ;
        RECT 99.645 8.565 99.815 8.765 ;
        RECT 89.345 7.295 89.520 8.435 ;
        RECT 91.550 7.560 92.245 8.190 ;
        RECT 91.550 6.960 91.720 7.560 ;
        RECT 91.890 7.340 92.225 7.370 ;
        RECT 92.615 7.340 92.785 8.020 ;
        RECT 91.890 7.170 92.785 7.340 ;
        RECT 93.850 7.560 94.545 8.190 ;
        RECT 94.715 7.560 95.410 8.190 ;
        RECT 96.095 7.560 96.790 8.190 ;
        RECT 91.890 7.120 92.225 7.170 ;
        RECT 93.850 6.960 94.020 7.560 ;
        RECT 94.190 7.340 94.525 7.370 ;
        RECT 94.735 7.340 95.070 7.370 ;
        RECT 94.190 7.170 95.070 7.340 ;
        RECT 94.190 7.120 94.525 7.170 ;
        RECT 94.735 7.120 95.070 7.170 ;
        RECT 95.240 6.960 95.410 7.560 ;
        RECT 95.580 7.120 95.915 7.390 ;
        RECT 96.115 7.120 96.450 7.370 ;
        RECT 96.620 6.960 96.790 7.560 ;
        RECT 96.960 7.120 97.295 7.390 ;
        RECT 99.645 7.305 99.820 8.565 ;
        RECT 100.230 8.535 100.400 10.145 ;
        RECT 100.600 10.085 100.775 10.595 ;
        RECT 101.030 10.045 101.205 10.595 ;
        RECT 102.395 10.085 102.565 10.595 ;
        RECT 103.385 10.085 103.555 10.595 ;
        RECT 100.170 8.365 100.400 8.535 ;
        RECT 100.600 8.565 100.770 9.515 ;
        RECT 100.170 7.305 100.340 8.365 ;
        RECT 100.600 7.305 100.775 8.565 ;
        RECT 101.030 8.445 101.200 10.045 ;
        RECT 101.960 9.425 102.190 9.610 ;
        RECT 101.960 9.380 102.490 9.425 ;
        RECT 102.020 9.255 102.490 9.380 ;
        RECT 103.010 9.255 103.480 9.425 ;
        RECT 102.020 8.565 102.190 9.255 ;
        RECT 102.390 8.780 102.560 8.885 ;
        RECT 103.010 8.780 103.180 9.255 ;
        RECT 102.390 8.605 103.180 8.780 ;
        RECT 101.030 7.305 101.205 8.445 ;
        RECT 102.390 7.305 102.565 8.605 ;
        RECT 103.010 8.565 103.180 8.605 ;
        RECT 103.380 8.450 103.550 8.885 ;
        RECT 103.380 7.305 103.555 8.450 ;
        RECT 22.605 5.980 22.935 6.960 ;
        RECT 24.905 5.980 25.235 6.960 ;
        RECT 26.265 5.980 26.595 6.960 ;
        RECT 27.645 5.980 27.975 6.960 ;
        RECT 39.825 5.980 40.155 6.960 ;
        RECT 42.125 5.980 42.455 6.960 ;
        RECT 43.485 5.980 43.815 6.960 ;
        RECT 44.865 5.980 45.195 6.960 ;
        RECT 57.045 5.980 57.375 6.960 ;
        RECT 59.345 5.980 59.675 6.960 ;
        RECT 60.705 5.980 61.035 6.960 ;
        RECT 62.085 5.980 62.415 6.960 ;
        RECT 74.265 5.980 74.595 6.960 ;
        RECT 76.565 5.980 76.895 6.960 ;
        RECT 77.925 5.980 78.255 6.960 ;
        RECT 79.305 5.980 79.635 6.960 ;
        RECT 91.485 5.980 91.815 6.960 ;
        RECT 93.785 5.980 94.115 6.960 ;
        RECT 95.145 5.980 95.475 6.960 ;
        RECT 96.525 5.980 96.855 6.960 ;
        RECT 22.135 4.490 22.465 5.470 ;
        RECT 23.945 4.670 24.275 5.455 ;
        RECT 23.595 4.500 24.275 4.670 ;
        RECT 24.465 4.670 24.795 5.455 ;
        RECT 24.465 4.500 25.145 4.670 ;
        RECT 22.135 3.890 22.385 4.490 ;
        RECT 22.555 4.280 22.885 4.330 ;
        RECT 23.075 4.280 23.425 4.330 ;
        RECT 22.555 4.110 23.425 4.280 ;
        RECT 22.555 4.080 22.885 4.110 ;
        RECT 23.075 4.080 23.425 4.110 ;
        RECT 23.595 3.900 23.765 4.500 ;
        RECT 23.935 4.080 24.285 4.330 ;
        RECT 24.455 4.080 24.805 4.330 ;
        RECT 24.975 3.900 25.145 4.500 ;
        RECT 25.835 4.620 26.155 5.470 ;
        RECT 26.335 4.960 26.735 5.470 ;
        RECT 27.245 4.960 27.575 5.470 ;
        RECT 26.335 4.790 27.575 4.960 ;
        RECT 28.155 4.620 28.325 5.300 ;
        RECT 28.505 4.790 28.885 5.470 ;
        RECT 25.835 4.540 26.285 4.620 ;
        RECT 25.835 4.370 26.465 4.540 ;
        RECT 25.315 4.080 25.665 4.330 ;
        RECT 22.135 3.260 22.465 3.890 ;
        RECT 23.525 3.260 23.855 3.900 ;
        RECT 24.885 3.260 25.215 3.900 ;
        RECT 26.295 3.490 26.465 4.370 ;
        RECT 27.240 4.450 28.545 4.620 ;
        RECT 26.635 3.830 26.865 4.330 ;
        RECT 27.240 4.250 27.410 4.450 ;
        RECT 27.035 4.080 27.410 4.250 ;
        RECT 27.580 4.080 28.130 4.280 ;
        RECT 28.300 4.000 28.545 4.450 ;
        RECT 28.715 3.830 28.885 4.790 ;
        RECT 26.635 3.660 28.885 3.830 ;
        RECT 30.765 3.895 30.940 5.155 ;
        RECT 31.290 4.095 31.460 5.155 ;
        RECT 31.290 3.925 31.520 4.095 ;
        RECT 30.765 3.695 30.935 3.895 ;
        RECT 26.295 3.320 27.250 3.490 ;
        RECT 28.165 3.340 28.335 3.660 ;
        RECT 30.765 3.365 31.175 3.695 ;
        RECT 30.765 2.855 30.935 3.365 ;
        RECT 30.765 2.525 31.175 2.855 ;
        RECT 30.765 2.355 30.935 2.525 ;
        RECT 30.765 1.865 30.940 2.355 ;
        RECT 31.350 2.315 31.520 3.925 ;
        RECT 31.720 3.895 31.895 5.155 ;
        RECT 32.150 4.015 32.325 5.155 ;
        RECT 31.720 2.945 31.890 3.895 ;
        RECT 32.150 2.415 32.320 4.015 ;
        RECT 33.510 4.010 33.685 5.155 ;
        RECT 39.355 4.490 39.685 5.470 ;
        RECT 41.165 4.670 41.495 5.455 ;
        RECT 40.815 4.500 41.495 4.670 ;
        RECT 41.685 4.670 42.015 5.455 ;
        RECT 41.685 4.500 42.365 4.670 ;
        RECT 33.140 3.205 33.310 3.895 ;
        RECT 33.510 3.805 33.680 4.010 ;
        RECT 34.125 3.805 34.295 3.895 ;
        RECT 33.510 3.625 34.295 3.805 ;
        RECT 33.510 3.575 33.680 3.625 ;
        RECT 34.125 3.205 34.295 3.625 ;
        RECT 39.355 3.890 39.605 4.490 ;
        RECT 39.775 4.280 40.105 4.330 ;
        RECT 40.295 4.280 40.645 4.330 ;
        RECT 39.775 4.110 40.645 4.280 ;
        RECT 39.775 4.080 40.105 4.110 ;
        RECT 40.295 4.080 40.645 4.110 ;
        RECT 40.815 3.900 40.985 4.500 ;
        RECT 41.155 4.080 41.505 4.330 ;
        RECT 41.675 4.080 42.025 4.330 ;
        RECT 42.195 3.900 42.365 4.500 ;
        RECT 43.055 4.620 43.375 5.470 ;
        RECT 43.555 4.960 43.955 5.470 ;
        RECT 44.465 4.960 44.795 5.470 ;
        RECT 43.555 4.790 44.795 4.960 ;
        RECT 45.375 4.620 45.545 5.300 ;
        RECT 45.725 4.790 46.105 5.470 ;
        RECT 43.055 4.540 43.505 4.620 ;
        RECT 43.055 4.370 43.685 4.540 ;
        RECT 42.535 4.080 42.885 4.330 ;
        RECT 39.355 3.260 39.685 3.890 ;
        RECT 40.745 3.260 41.075 3.900 ;
        RECT 42.105 3.260 42.435 3.900 ;
        RECT 43.515 3.490 43.685 4.370 ;
        RECT 44.460 4.450 45.765 4.620 ;
        RECT 43.855 3.830 44.085 4.330 ;
        RECT 44.460 4.250 44.630 4.450 ;
        RECT 44.255 4.080 44.630 4.250 ;
        RECT 44.800 4.080 45.350 4.280 ;
        RECT 45.520 4.000 45.765 4.450 ;
        RECT 45.935 3.830 46.105 4.790 ;
        RECT 43.855 3.660 46.105 3.830 ;
        RECT 47.985 3.895 48.160 5.155 ;
        RECT 48.510 4.095 48.680 5.155 ;
        RECT 48.510 3.925 48.740 4.095 ;
        RECT 47.985 3.695 48.155 3.895 ;
        RECT 43.515 3.320 44.470 3.490 ;
        RECT 45.385 3.340 45.555 3.660 ;
        RECT 47.985 3.365 48.395 3.695 ;
        RECT 33.140 3.175 33.610 3.205 ;
        RECT 33.095 3.035 33.610 3.175 ;
        RECT 34.125 3.035 34.595 3.205 ;
        RECT 33.095 2.945 33.325 3.035 ;
        RECT 47.985 2.855 48.155 3.365 ;
        RECT 47.985 2.525 48.395 2.855 ;
        RECT 31.290 2.145 31.520 2.315 ;
        RECT 31.290 1.865 31.460 2.145 ;
        RECT 31.720 1.865 31.895 2.375 ;
        RECT 32.150 1.865 32.325 2.415 ;
        RECT 33.515 1.865 33.685 2.375 ;
        RECT 47.985 2.355 48.155 2.525 ;
        RECT 47.985 1.865 48.160 2.355 ;
        RECT 48.570 2.315 48.740 3.925 ;
        RECT 48.940 3.895 49.115 5.155 ;
        RECT 49.370 4.015 49.545 5.155 ;
        RECT 48.940 2.945 49.110 3.895 ;
        RECT 49.370 2.415 49.540 4.015 ;
        RECT 50.730 4.010 50.905 5.155 ;
        RECT 56.575 4.490 56.905 5.470 ;
        RECT 58.385 4.670 58.715 5.455 ;
        RECT 58.035 4.500 58.715 4.670 ;
        RECT 58.905 4.670 59.235 5.455 ;
        RECT 58.905 4.500 59.585 4.670 ;
        RECT 50.360 3.205 50.530 3.895 ;
        RECT 50.730 3.805 50.900 4.010 ;
        RECT 51.345 3.805 51.515 3.895 ;
        RECT 50.730 3.625 51.515 3.805 ;
        RECT 50.730 3.575 50.900 3.625 ;
        RECT 51.345 3.205 51.515 3.625 ;
        RECT 56.575 3.890 56.825 4.490 ;
        RECT 56.995 4.280 57.325 4.330 ;
        RECT 57.515 4.280 57.865 4.330 ;
        RECT 56.995 4.110 57.865 4.280 ;
        RECT 56.995 4.080 57.325 4.110 ;
        RECT 57.515 4.080 57.865 4.110 ;
        RECT 58.035 3.900 58.205 4.500 ;
        RECT 58.375 4.080 58.725 4.330 ;
        RECT 58.895 4.080 59.245 4.330 ;
        RECT 59.415 3.900 59.585 4.500 ;
        RECT 60.275 4.620 60.595 5.470 ;
        RECT 60.775 4.960 61.175 5.470 ;
        RECT 61.685 4.960 62.015 5.470 ;
        RECT 60.775 4.790 62.015 4.960 ;
        RECT 62.595 4.620 62.765 5.300 ;
        RECT 62.945 4.790 63.325 5.470 ;
        RECT 60.275 4.540 60.725 4.620 ;
        RECT 60.275 4.370 60.905 4.540 ;
        RECT 59.755 4.080 60.105 4.330 ;
        RECT 56.575 3.260 56.905 3.890 ;
        RECT 57.965 3.260 58.295 3.900 ;
        RECT 59.325 3.260 59.655 3.900 ;
        RECT 60.735 3.490 60.905 4.370 ;
        RECT 61.680 4.450 62.985 4.620 ;
        RECT 61.075 3.830 61.305 4.330 ;
        RECT 61.680 4.250 61.850 4.450 ;
        RECT 61.475 4.080 61.850 4.250 ;
        RECT 62.020 4.080 62.570 4.280 ;
        RECT 62.740 4.000 62.985 4.450 ;
        RECT 63.155 3.830 63.325 4.790 ;
        RECT 61.075 3.660 63.325 3.830 ;
        RECT 65.205 3.895 65.380 5.155 ;
        RECT 65.730 4.095 65.900 5.155 ;
        RECT 65.730 3.925 65.960 4.095 ;
        RECT 65.205 3.695 65.375 3.895 ;
        RECT 60.735 3.320 61.690 3.490 ;
        RECT 62.605 3.340 62.775 3.660 ;
        RECT 65.205 3.365 65.615 3.695 ;
        RECT 50.360 3.175 50.830 3.205 ;
        RECT 50.315 3.035 50.830 3.175 ;
        RECT 51.345 3.035 51.815 3.205 ;
        RECT 50.315 2.945 50.545 3.035 ;
        RECT 65.205 2.855 65.375 3.365 ;
        RECT 65.205 2.525 65.615 2.855 ;
        RECT 48.510 2.145 48.740 2.315 ;
        RECT 48.510 1.865 48.680 2.145 ;
        RECT 48.940 1.865 49.115 2.375 ;
        RECT 49.370 1.865 49.545 2.415 ;
        RECT 50.735 1.865 50.905 2.375 ;
        RECT 65.205 2.355 65.375 2.525 ;
        RECT 65.205 1.865 65.380 2.355 ;
        RECT 65.790 2.315 65.960 3.925 ;
        RECT 66.160 3.895 66.335 5.155 ;
        RECT 66.590 4.015 66.765 5.155 ;
        RECT 66.160 2.945 66.330 3.895 ;
        RECT 66.590 2.415 66.760 4.015 ;
        RECT 67.950 4.010 68.125 5.155 ;
        RECT 73.795 4.490 74.125 5.470 ;
        RECT 75.605 4.670 75.935 5.455 ;
        RECT 75.255 4.500 75.935 4.670 ;
        RECT 76.125 4.670 76.455 5.455 ;
        RECT 76.125 4.500 76.805 4.670 ;
        RECT 67.580 3.205 67.750 3.895 ;
        RECT 67.950 3.805 68.120 4.010 ;
        RECT 68.565 3.805 68.735 3.895 ;
        RECT 67.950 3.625 68.735 3.805 ;
        RECT 67.950 3.575 68.120 3.625 ;
        RECT 68.565 3.205 68.735 3.625 ;
        RECT 73.795 3.890 74.045 4.490 ;
        RECT 74.215 4.280 74.545 4.330 ;
        RECT 74.735 4.280 75.085 4.330 ;
        RECT 74.215 4.110 75.085 4.280 ;
        RECT 74.215 4.080 74.545 4.110 ;
        RECT 74.735 4.080 75.085 4.110 ;
        RECT 75.255 3.900 75.425 4.500 ;
        RECT 75.595 4.080 75.945 4.330 ;
        RECT 76.115 4.080 76.465 4.330 ;
        RECT 76.635 3.900 76.805 4.500 ;
        RECT 77.495 4.620 77.815 5.470 ;
        RECT 77.995 4.960 78.395 5.470 ;
        RECT 78.905 4.960 79.235 5.470 ;
        RECT 77.995 4.790 79.235 4.960 ;
        RECT 79.815 4.620 79.985 5.300 ;
        RECT 80.165 4.790 80.545 5.470 ;
        RECT 77.495 4.540 77.945 4.620 ;
        RECT 77.495 4.370 78.125 4.540 ;
        RECT 76.975 4.080 77.325 4.330 ;
        RECT 73.795 3.260 74.125 3.890 ;
        RECT 75.185 3.260 75.515 3.900 ;
        RECT 76.545 3.260 76.875 3.900 ;
        RECT 77.955 3.490 78.125 4.370 ;
        RECT 78.900 4.450 80.205 4.620 ;
        RECT 78.295 3.830 78.525 4.330 ;
        RECT 78.900 4.250 79.070 4.450 ;
        RECT 78.695 4.080 79.070 4.250 ;
        RECT 79.240 4.080 79.790 4.280 ;
        RECT 79.960 4.000 80.205 4.450 ;
        RECT 80.375 3.830 80.545 4.790 ;
        RECT 78.295 3.660 80.545 3.830 ;
        RECT 82.425 3.895 82.600 5.155 ;
        RECT 82.950 4.095 83.120 5.155 ;
        RECT 82.950 3.925 83.180 4.095 ;
        RECT 82.425 3.695 82.595 3.895 ;
        RECT 77.955 3.320 78.910 3.490 ;
        RECT 79.825 3.340 79.995 3.660 ;
        RECT 82.425 3.365 82.835 3.695 ;
        RECT 67.580 3.175 68.050 3.205 ;
        RECT 67.535 3.035 68.050 3.175 ;
        RECT 68.565 3.035 69.035 3.205 ;
        RECT 67.535 2.945 67.765 3.035 ;
        RECT 82.425 2.855 82.595 3.365 ;
        RECT 82.425 2.525 82.835 2.855 ;
        RECT 65.730 2.145 65.960 2.315 ;
        RECT 65.730 1.865 65.900 2.145 ;
        RECT 66.160 1.865 66.335 2.375 ;
        RECT 66.590 1.865 66.765 2.415 ;
        RECT 67.955 1.865 68.125 2.375 ;
        RECT 82.425 2.355 82.595 2.525 ;
        RECT 82.425 1.865 82.600 2.355 ;
        RECT 83.010 2.315 83.180 3.925 ;
        RECT 83.380 3.895 83.555 5.155 ;
        RECT 83.810 4.015 83.985 5.155 ;
        RECT 83.380 2.945 83.550 3.895 ;
        RECT 83.810 2.415 83.980 4.015 ;
        RECT 85.170 4.010 85.345 5.155 ;
        RECT 91.015 4.490 91.345 5.470 ;
        RECT 92.825 4.670 93.155 5.455 ;
        RECT 92.475 4.500 93.155 4.670 ;
        RECT 93.345 4.670 93.675 5.455 ;
        RECT 93.345 4.500 94.025 4.670 ;
        RECT 84.800 3.205 84.970 3.895 ;
        RECT 85.170 3.805 85.340 4.010 ;
        RECT 85.785 3.805 85.955 3.895 ;
        RECT 85.170 3.625 85.955 3.805 ;
        RECT 85.170 3.575 85.340 3.625 ;
        RECT 85.785 3.205 85.955 3.625 ;
        RECT 91.015 3.890 91.265 4.490 ;
        RECT 91.435 4.280 91.765 4.330 ;
        RECT 91.955 4.280 92.305 4.330 ;
        RECT 91.435 4.110 92.305 4.280 ;
        RECT 91.435 4.080 91.765 4.110 ;
        RECT 91.955 4.080 92.305 4.110 ;
        RECT 92.475 3.900 92.645 4.500 ;
        RECT 92.815 4.080 93.165 4.330 ;
        RECT 93.335 4.080 93.685 4.330 ;
        RECT 93.855 3.900 94.025 4.500 ;
        RECT 94.715 4.620 95.035 5.470 ;
        RECT 95.215 4.960 95.615 5.470 ;
        RECT 96.125 4.960 96.455 5.470 ;
        RECT 95.215 4.790 96.455 4.960 ;
        RECT 97.035 4.620 97.205 5.300 ;
        RECT 97.385 4.790 97.765 5.470 ;
        RECT 94.715 4.540 95.165 4.620 ;
        RECT 94.715 4.370 95.345 4.540 ;
        RECT 94.195 4.080 94.545 4.330 ;
        RECT 91.015 3.260 91.345 3.890 ;
        RECT 92.405 3.260 92.735 3.900 ;
        RECT 93.765 3.260 94.095 3.900 ;
        RECT 95.175 3.490 95.345 4.370 ;
        RECT 96.120 4.450 97.425 4.620 ;
        RECT 95.515 3.830 95.745 4.330 ;
        RECT 96.120 4.250 96.290 4.450 ;
        RECT 95.915 4.080 96.290 4.250 ;
        RECT 96.460 4.080 97.010 4.280 ;
        RECT 97.180 4.000 97.425 4.450 ;
        RECT 97.595 3.830 97.765 4.790 ;
        RECT 95.515 3.660 97.765 3.830 ;
        RECT 99.645 3.895 99.820 5.155 ;
        RECT 100.170 4.095 100.340 5.155 ;
        RECT 100.170 3.925 100.400 4.095 ;
        RECT 99.645 3.695 99.815 3.895 ;
        RECT 95.175 3.320 96.130 3.490 ;
        RECT 97.045 3.340 97.215 3.660 ;
        RECT 99.645 3.365 100.055 3.695 ;
        RECT 84.800 3.175 85.270 3.205 ;
        RECT 84.755 3.035 85.270 3.175 ;
        RECT 85.785 3.035 86.255 3.205 ;
        RECT 84.755 2.945 84.985 3.035 ;
        RECT 99.645 2.855 99.815 3.365 ;
        RECT 99.645 2.525 100.055 2.855 ;
        RECT 82.950 2.145 83.180 2.315 ;
        RECT 82.950 1.865 83.120 2.145 ;
        RECT 83.380 1.865 83.555 2.375 ;
        RECT 83.810 1.865 83.985 2.415 ;
        RECT 85.175 1.865 85.345 2.375 ;
        RECT 99.645 2.355 99.815 2.525 ;
        RECT 99.645 1.865 99.820 2.355 ;
        RECT 100.230 2.315 100.400 3.925 ;
        RECT 100.600 3.895 100.775 5.155 ;
        RECT 101.030 4.015 101.205 5.155 ;
        RECT 100.600 2.945 100.770 3.895 ;
        RECT 101.030 2.415 101.200 4.015 ;
        RECT 102.390 4.010 102.565 5.155 ;
        RECT 102.020 3.205 102.190 3.895 ;
        RECT 102.390 3.805 102.560 4.010 ;
        RECT 103.005 3.805 103.175 3.895 ;
        RECT 102.390 3.625 103.175 3.805 ;
        RECT 102.390 3.575 102.560 3.625 ;
        RECT 103.005 3.205 103.175 3.625 ;
        RECT 102.020 3.175 102.490 3.205 ;
        RECT 101.975 3.035 102.490 3.175 ;
        RECT 103.005 3.035 103.475 3.205 ;
        RECT 101.975 2.945 102.205 3.035 ;
        RECT 100.170 2.145 100.400 2.315 ;
        RECT 100.170 1.865 100.340 2.145 ;
        RECT 100.600 1.865 100.775 2.375 ;
        RECT 101.030 1.865 101.205 2.415 ;
        RECT 102.395 1.865 102.565 2.375 ;
      LAYER met1 ;
        RECT 16.565 10.055 16.855 10.285 ;
        RECT 16.625 9.590 16.795 10.055 ;
        RECT 19.975 10.045 20.265 10.275 ;
        RECT 31.660 10.055 31.950 10.285 ;
        RECT 20.035 9.680 20.205 10.045 ;
        RECT 16.535 9.310 16.875 9.590 ;
        RECT 19.940 9.310 20.310 9.680 ;
        RECT 31.720 9.575 31.890 10.055 ;
        RECT 33.450 10.025 33.745 10.285 ;
        RECT 34.440 10.025 34.735 10.285 ;
        RECT 37.195 10.045 37.485 10.275 ;
        RECT 48.880 10.055 49.170 10.285 ;
        RECT 33.080 9.650 33.310 9.670 ;
        RECT 33.050 9.575 33.340 9.650 ;
        RECT 31.720 9.545 33.340 9.575 ;
        RECT 31.660 9.405 33.340 9.545 ;
        RECT 31.660 9.315 31.950 9.405 ;
        RECT 33.050 9.340 33.340 9.405 ;
        RECT 33.080 9.315 33.310 9.340 ;
        RECT 19.975 9.305 20.265 9.310 ;
        RECT 32.115 9.175 32.440 9.265 ;
        RECT 20.405 9.140 20.695 9.165 ;
        RECT 32.090 9.145 32.440 9.175 ;
        RECT 20.385 9.135 20.725 9.140 ;
        RECT 20.235 8.965 20.725 9.135 ;
        RECT 31.920 8.975 32.440 9.145 ;
        RECT 20.385 8.860 20.725 8.965 ;
        RECT 32.090 8.945 32.440 8.975 ;
        RECT 32.115 8.940 32.440 8.945 ;
        RECT 33.510 8.925 33.680 10.025 ;
        RECT 34.500 9.270 34.670 10.025 ;
        RECT 37.255 9.680 37.425 10.045 ;
        RECT 37.160 9.310 37.530 9.680 ;
        RECT 48.940 9.575 49.110 10.055 ;
        RECT 50.670 10.025 50.965 10.285 ;
        RECT 51.660 10.025 51.955 10.285 ;
        RECT 54.415 10.045 54.705 10.275 ;
        RECT 66.100 10.055 66.390 10.285 ;
        RECT 50.300 9.650 50.530 9.670 ;
        RECT 50.270 9.575 50.560 9.650 ;
        RECT 48.940 9.545 50.560 9.575 ;
        RECT 48.880 9.405 50.560 9.545 ;
        RECT 48.880 9.315 49.170 9.405 ;
        RECT 50.270 9.340 50.560 9.405 ;
        RECT 50.300 9.315 50.530 9.340 ;
        RECT 37.195 9.305 37.485 9.310 ;
        RECT 34.500 8.945 34.830 9.270 ;
        RECT 49.335 9.175 49.660 9.265 ;
        RECT 37.625 9.140 37.915 9.165 ;
        RECT 49.310 9.145 49.660 9.175 ;
        RECT 37.605 9.135 37.945 9.140 ;
        RECT 37.455 8.965 37.945 9.135 ;
        RECT 49.140 8.975 49.660 9.145 ;
        RECT 34.500 8.925 34.790 8.945 ;
        RECT 33.450 8.920 33.680 8.925 ;
        RECT 16.160 8.785 16.500 8.850 ;
        RECT 31.315 8.815 31.635 8.890 ;
        RECT 31.290 8.785 31.635 8.815 ;
        RECT 16.020 8.615 16.500 8.785 ;
        RECT 31.115 8.615 31.635 8.785 ;
        RECT 33.450 8.685 33.740 8.920 ;
        RECT 34.440 8.835 34.790 8.925 ;
        RECT 37.605 8.860 37.945 8.965 ;
        RECT 49.310 8.945 49.660 8.975 ;
        RECT 49.335 8.940 49.660 8.945 ;
        RECT 50.730 8.925 50.900 10.025 ;
        RECT 51.720 9.270 51.890 10.025 ;
        RECT 54.475 9.680 54.645 10.045 ;
        RECT 54.380 9.310 54.750 9.680 ;
        RECT 66.160 9.575 66.330 10.055 ;
        RECT 67.890 10.025 68.185 10.285 ;
        RECT 68.880 10.025 69.175 10.285 ;
        RECT 71.635 10.045 71.925 10.275 ;
        RECT 83.320 10.055 83.610 10.285 ;
        RECT 67.520 9.650 67.750 9.670 ;
        RECT 67.490 9.575 67.780 9.650 ;
        RECT 66.160 9.545 67.780 9.575 ;
        RECT 66.100 9.405 67.780 9.545 ;
        RECT 66.100 9.315 66.390 9.405 ;
        RECT 67.490 9.340 67.780 9.405 ;
        RECT 67.520 9.315 67.750 9.340 ;
        RECT 54.415 9.305 54.705 9.310 ;
        RECT 51.720 8.945 52.050 9.270 ;
        RECT 66.555 9.175 66.880 9.265 ;
        RECT 54.845 9.140 55.135 9.165 ;
        RECT 66.530 9.145 66.880 9.175 ;
        RECT 54.825 9.135 55.165 9.140 ;
        RECT 54.675 8.965 55.165 9.135 ;
        RECT 66.360 8.975 66.880 9.145 ;
        RECT 51.720 8.925 52.010 8.945 ;
        RECT 50.670 8.920 50.900 8.925 ;
        RECT 34.440 8.685 34.730 8.835 ;
        RECT 48.535 8.815 48.855 8.890 ;
        RECT 48.510 8.785 48.855 8.815 ;
        RECT 48.335 8.615 48.855 8.785 ;
        RECT 50.670 8.685 50.960 8.920 ;
        RECT 51.660 8.845 52.010 8.925 ;
        RECT 54.825 8.860 55.165 8.965 ;
        RECT 66.530 8.945 66.880 8.975 ;
        RECT 66.555 8.940 66.880 8.945 ;
        RECT 67.950 8.925 68.120 10.025 ;
        RECT 68.940 9.270 69.110 10.025 ;
        RECT 71.695 9.680 71.865 10.045 ;
        RECT 71.600 9.310 71.970 9.680 ;
        RECT 83.380 9.575 83.550 10.055 ;
        RECT 85.110 10.025 85.405 10.285 ;
        RECT 86.100 10.025 86.395 10.285 ;
        RECT 88.855 10.045 89.145 10.275 ;
        RECT 100.540 10.055 100.830 10.285 ;
        RECT 84.740 9.650 84.970 9.670 ;
        RECT 84.710 9.575 85.000 9.650 ;
        RECT 83.380 9.545 85.000 9.575 ;
        RECT 83.320 9.405 85.000 9.545 ;
        RECT 83.320 9.315 83.610 9.405 ;
        RECT 84.710 9.340 85.000 9.405 ;
        RECT 84.740 9.315 84.970 9.340 ;
        RECT 71.635 9.305 71.925 9.310 ;
        RECT 68.940 8.945 69.270 9.270 ;
        RECT 83.775 9.175 84.100 9.265 ;
        RECT 72.065 9.140 72.355 9.165 ;
        RECT 83.750 9.145 84.100 9.175 ;
        RECT 72.045 9.135 72.385 9.140 ;
        RECT 71.895 8.965 72.385 9.135 ;
        RECT 83.580 8.975 84.100 9.145 ;
        RECT 68.940 8.925 69.230 8.945 ;
        RECT 67.890 8.920 68.120 8.925 ;
        RECT 51.660 8.685 51.950 8.845 ;
        RECT 65.755 8.815 66.075 8.890 ;
        RECT 65.730 8.785 66.075 8.815 ;
        RECT 65.555 8.615 66.075 8.785 ;
        RECT 67.890 8.685 68.180 8.920 ;
        RECT 68.880 8.825 69.230 8.925 ;
        RECT 72.045 8.860 72.385 8.965 ;
        RECT 83.750 8.945 84.100 8.975 ;
        RECT 83.775 8.940 84.100 8.945 ;
        RECT 85.170 8.925 85.340 10.025 ;
        RECT 86.160 9.270 86.330 10.025 ;
        RECT 88.915 9.680 89.085 10.045 ;
        RECT 88.820 9.310 89.190 9.680 ;
        RECT 100.600 9.575 100.770 10.055 ;
        RECT 102.330 10.025 102.625 10.285 ;
        RECT 103.320 10.025 103.615 10.285 ;
        RECT 101.960 9.650 102.190 9.670 ;
        RECT 101.930 9.575 102.220 9.650 ;
        RECT 100.600 9.545 102.220 9.575 ;
        RECT 100.540 9.405 102.220 9.545 ;
        RECT 100.540 9.315 100.830 9.405 ;
        RECT 101.930 9.340 102.220 9.405 ;
        RECT 101.960 9.315 102.190 9.340 ;
        RECT 88.855 9.305 89.145 9.310 ;
        RECT 86.160 8.945 86.490 9.270 ;
        RECT 100.995 9.175 101.320 9.265 ;
        RECT 89.285 9.140 89.575 9.165 ;
        RECT 100.970 9.145 101.320 9.175 ;
        RECT 89.265 9.135 89.605 9.140 ;
        RECT 89.115 8.965 89.605 9.135 ;
        RECT 100.800 8.975 101.320 9.145 ;
        RECT 86.160 8.925 86.450 8.945 ;
        RECT 85.110 8.920 85.340 8.925 ;
        RECT 68.880 8.685 69.170 8.825 ;
        RECT 82.975 8.815 83.295 8.890 ;
        RECT 82.950 8.785 83.295 8.815 ;
        RECT 82.775 8.615 83.295 8.785 ;
        RECT 85.110 8.685 85.400 8.920 ;
        RECT 86.100 8.805 86.450 8.925 ;
        RECT 89.265 8.860 89.605 8.965 ;
        RECT 100.970 8.945 101.320 8.975 ;
        RECT 100.995 8.940 101.320 8.945 ;
        RECT 102.390 8.925 102.560 10.025 ;
        RECT 103.350 10.010 103.615 10.025 ;
        RECT 103.350 9.585 103.675 10.010 ;
        RECT 103.380 8.925 103.550 9.585 ;
        RECT 102.330 8.920 102.560 8.925 ;
        RECT 103.320 8.920 103.550 8.925 ;
        RECT 100.195 8.815 100.515 8.890 ;
        RECT 86.100 8.685 86.390 8.805 ;
        RECT 100.170 8.785 100.515 8.815 ;
        RECT 99.995 8.615 100.515 8.785 ;
        RECT 102.330 8.685 102.620 8.920 ;
        RECT 103.320 8.685 103.610 8.920 ;
        RECT 16.160 8.570 16.500 8.615 ;
        RECT 31.290 8.585 31.635 8.615 ;
        RECT 48.510 8.585 48.855 8.615 ;
        RECT 65.730 8.585 66.075 8.615 ;
        RECT 82.950 8.585 83.295 8.615 ;
        RECT 100.170 8.585 100.515 8.615 ;
        RECT 31.315 8.565 31.635 8.585 ;
        RECT 48.535 8.565 48.855 8.585 ;
        RECT 65.755 8.565 66.075 8.585 ;
        RECT 82.975 8.565 83.295 8.585 ;
        RECT 100.195 8.565 100.515 8.585 ;
        RECT 23.675 8.005 23.965 8.050 ;
        RECT 24.680 8.005 25.000 8.035 ;
        RECT 26.040 8.005 26.360 8.050 ;
        RECT 23.675 7.865 25.590 8.005 ;
        RECT 23.675 7.820 23.965 7.865 ;
        RECT 24.675 7.835 25.005 7.865 ;
        RECT 24.680 7.775 25.000 7.835 ;
        RECT 25.450 7.650 25.590 7.865 ;
        RECT 26.040 7.865 26.635 8.005 ;
        RECT 26.040 7.790 26.360 7.865 ;
        RECT 27.415 7.805 28.060 8.050 ;
        RECT 40.895 8.005 41.185 8.050 ;
        RECT 41.900 8.005 42.220 8.035 ;
        RECT 43.260 8.005 43.580 8.050 ;
        RECT 40.895 7.865 42.810 8.005 ;
        RECT 40.895 7.820 41.185 7.865 ;
        RECT 41.895 7.835 42.225 7.865 ;
        RECT 27.740 7.775 28.060 7.805 ;
        RECT 41.900 7.775 42.220 7.835 ;
        RECT 42.670 7.650 42.810 7.865 ;
        RECT 43.260 7.865 43.855 8.005 ;
        RECT 43.260 7.790 43.580 7.865 ;
        RECT 44.635 7.805 45.280 8.050 ;
        RECT 58.115 8.005 58.405 8.050 ;
        RECT 59.120 8.005 59.440 8.035 ;
        RECT 60.480 8.005 60.800 8.050 ;
        RECT 58.115 7.865 60.030 8.005 ;
        RECT 58.115 7.820 58.405 7.865 ;
        RECT 59.115 7.835 59.445 7.865 ;
        RECT 44.960 7.775 45.280 7.805 ;
        RECT 59.120 7.775 59.440 7.835 ;
        RECT 59.890 7.650 60.030 7.865 ;
        RECT 60.480 7.865 61.075 8.005 ;
        RECT 60.480 7.790 60.800 7.865 ;
        RECT 61.855 7.805 62.500 8.050 ;
        RECT 75.335 8.005 75.625 8.050 ;
        RECT 76.340 8.005 76.660 8.035 ;
        RECT 77.700 8.005 78.020 8.050 ;
        RECT 75.335 7.865 77.250 8.005 ;
        RECT 75.335 7.820 75.625 7.865 ;
        RECT 76.335 7.835 76.665 7.865 ;
        RECT 62.180 7.775 62.500 7.805 ;
        RECT 76.340 7.775 76.660 7.835 ;
        RECT 77.110 7.650 77.250 7.865 ;
        RECT 77.700 7.865 78.295 8.005 ;
        RECT 77.700 7.790 78.020 7.865 ;
        RECT 79.075 7.805 79.720 8.050 ;
        RECT 92.555 8.005 92.845 8.050 ;
        RECT 93.560 8.005 93.880 8.035 ;
        RECT 94.920 8.005 95.240 8.050 ;
        RECT 92.555 7.865 94.470 8.005 ;
        RECT 92.555 7.820 92.845 7.865 ;
        RECT 93.555 7.835 93.885 7.865 ;
        RECT 79.400 7.775 79.720 7.805 ;
        RECT 93.560 7.775 93.880 7.835 ;
        RECT 94.330 7.650 94.470 7.865 ;
        RECT 94.920 7.865 95.515 8.005 ;
        RECT 94.920 7.790 95.240 7.865 ;
        RECT 96.295 7.805 96.940 8.050 ;
        RECT 96.620 7.775 96.940 7.805 ;
        RECT 25.450 7.510 27.460 7.650 ;
        RECT 42.670 7.510 44.680 7.650 ;
        RECT 59.890 7.510 61.900 7.650 ;
        RECT 77.110 7.510 79.120 7.650 ;
        RECT 94.330 7.510 96.340 7.650 ;
        RECT 27.320 7.370 27.460 7.510 ;
        RECT 44.540 7.370 44.680 7.510 ;
        RECT 61.760 7.370 61.900 7.510 ;
        RECT 78.980 7.370 79.120 7.510 ;
        RECT 96.200 7.370 96.340 7.510 ;
        RECT 25.365 7.125 26.010 7.370 ;
        RECT 25.690 7.110 26.010 7.125 ;
        RECT 26.720 7.110 27.040 7.370 ;
        RECT 27.245 7.140 27.535 7.370 ;
        RECT 28.095 7.140 28.385 7.370 ;
        RECT 26.810 6.970 26.950 7.110 ;
        RECT 28.170 6.970 28.310 7.140 ;
        RECT 42.585 7.125 43.230 7.370 ;
        RECT 42.910 7.110 43.230 7.125 ;
        RECT 43.940 7.110 44.260 7.370 ;
        RECT 44.465 7.140 44.755 7.370 ;
        RECT 45.315 7.140 45.605 7.370 ;
        RECT 26.810 6.830 28.310 6.970 ;
        RECT 44.030 6.970 44.170 7.110 ;
        RECT 45.390 6.970 45.530 7.140 ;
        RECT 59.805 7.125 60.450 7.370 ;
        RECT 60.130 7.110 60.450 7.125 ;
        RECT 61.160 7.110 61.480 7.370 ;
        RECT 61.685 7.140 61.975 7.370 ;
        RECT 62.535 7.140 62.825 7.370 ;
        RECT 44.030 6.830 45.530 6.970 ;
        RECT 61.250 6.970 61.390 7.110 ;
        RECT 62.610 6.970 62.750 7.140 ;
        RECT 77.025 7.125 77.670 7.370 ;
        RECT 77.350 7.110 77.670 7.125 ;
        RECT 78.380 7.110 78.700 7.370 ;
        RECT 78.905 7.140 79.195 7.370 ;
        RECT 79.755 7.140 80.045 7.370 ;
        RECT 61.250 6.830 62.750 6.970 ;
        RECT 78.470 6.970 78.610 7.110 ;
        RECT 79.830 6.970 79.970 7.140 ;
        RECT 94.245 7.125 94.890 7.370 ;
        RECT 94.570 7.110 94.890 7.125 ;
        RECT 95.600 7.110 95.920 7.370 ;
        RECT 96.125 7.140 96.415 7.370 ;
        RECT 96.975 7.140 97.265 7.370 ;
        RECT 78.470 6.830 79.970 6.970 ;
        RECT 95.690 6.970 95.830 7.110 ;
        RECT 97.050 6.970 97.190 7.140 ;
        RECT 95.690 6.830 97.190 6.970 ;
        RECT 22.640 6.305 22.960 6.365 ;
        RECT 22.365 6.165 22.960 6.305 ;
        RECT 22.640 6.105 22.960 6.165 ;
        RECT 24.915 6.305 25.205 6.350 ;
        RECT 27.060 6.305 27.380 6.365 ;
        RECT 39.860 6.305 40.180 6.365 ;
        RECT 24.915 6.165 27.380 6.305 ;
        RECT 39.585 6.165 40.180 6.305 ;
        RECT 24.915 6.120 25.205 6.165 ;
        RECT 27.060 6.105 27.380 6.165 ;
        RECT 39.860 6.105 40.180 6.165 ;
        RECT 42.135 6.305 42.425 6.350 ;
        RECT 44.280 6.305 44.600 6.365 ;
        RECT 57.080 6.305 57.400 6.365 ;
        RECT 42.135 6.165 44.600 6.305 ;
        RECT 56.805 6.165 57.400 6.305 ;
        RECT 42.135 6.120 42.425 6.165 ;
        RECT 44.280 6.105 44.600 6.165 ;
        RECT 57.080 6.105 57.400 6.165 ;
        RECT 59.355 6.305 59.645 6.350 ;
        RECT 61.500 6.305 61.820 6.365 ;
        RECT 74.300 6.305 74.620 6.365 ;
        RECT 59.355 6.165 61.820 6.305 ;
        RECT 74.025 6.165 74.620 6.305 ;
        RECT 59.355 6.120 59.645 6.165 ;
        RECT 61.500 6.105 61.820 6.165 ;
        RECT 74.300 6.105 74.620 6.165 ;
        RECT 76.575 6.305 76.865 6.350 ;
        RECT 78.720 6.305 79.040 6.365 ;
        RECT 91.520 6.305 91.840 6.365 ;
        RECT 76.575 6.165 79.040 6.305 ;
        RECT 91.245 6.165 91.840 6.305 ;
        RECT 76.575 6.120 76.865 6.165 ;
        RECT 78.720 6.105 79.040 6.165 ;
        RECT 91.520 6.105 91.840 6.165 ;
        RECT 93.795 6.305 94.085 6.350 ;
        RECT 95.940 6.305 96.260 6.365 ;
        RECT 93.795 6.165 96.260 6.305 ;
        RECT 93.795 6.120 94.085 6.165 ;
        RECT 95.940 6.105 96.260 6.165 ;
        RECT 24.015 5.285 24.305 5.330 ;
        RECT 26.380 5.285 26.700 5.345 ;
        RECT 24.015 5.145 26.700 5.285 ;
        RECT 24.015 5.100 24.305 5.145 ;
        RECT 26.380 5.085 26.700 5.145 ;
        RECT 27.060 5.285 27.380 5.345 ;
        RECT 28.095 5.285 28.385 5.330 ;
        RECT 27.060 5.145 28.385 5.285 ;
        RECT 27.060 5.085 27.380 5.145 ;
        RECT 28.095 5.100 28.385 5.145 ;
        RECT 41.235 5.285 41.525 5.330 ;
        RECT 43.600 5.285 43.920 5.345 ;
        RECT 41.235 5.145 43.920 5.285 ;
        RECT 41.235 5.100 41.525 5.145 ;
        RECT 43.600 5.085 43.920 5.145 ;
        RECT 44.280 5.285 44.600 5.345 ;
        RECT 45.315 5.285 45.605 5.330 ;
        RECT 44.280 5.145 45.605 5.285 ;
        RECT 44.280 5.085 44.600 5.145 ;
        RECT 45.315 5.100 45.605 5.145 ;
        RECT 58.455 5.285 58.745 5.330 ;
        RECT 60.820 5.285 61.140 5.345 ;
        RECT 58.455 5.145 61.140 5.285 ;
        RECT 58.455 5.100 58.745 5.145 ;
        RECT 60.820 5.085 61.140 5.145 ;
        RECT 61.500 5.285 61.820 5.345 ;
        RECT 62.535 5.285 62.825 5.330 ;
        RECT 61.500 5.145 62.825 5.285 ;
        RECT 61.500 5.085 61.820 5.145 ;
        RECT 62.535 5.100 62.825 5.145 ;
        RECT 75.675 5.285 75.965 5.330 ;
        RECT 78.040 5.285 78.360 5.345 ;
        RECT 75.675 5.145 78.360 5.285 ;
        RECT 75.675 5.100 75.965 5.145 ;
        RECT 78.040 5.085 78.360 5.145 ;
        RECT 78.720 5.285 79.040 5.345 ;
        RECT 79.755 5.285 80.045 5.330 ;
        RECT 78.720 5.145 80.045 5.285 ;
        RECT 78.720 5.085 79.040 5.145 ;
        RECT 79.755 5.100 80.045 5.145 ;
        RECT 92.895 5.285 93.185 5.330 ;
        RECT 95.260 5.285 95.580 5.345 ;
        RECT 92.895 5.145 95.580 5.285 ;
        RECT 92.895 5.100 93.185 5.145 ;
        RECT 95.260 5.085 95.580 5.145 ;
        RECT 95.940 5.285 96.260 5.345 ;
        RECT 96.975 5.285 97.265 5.330 ;
        RECT 95.940 5.145 97.265 5.285 ;
        RECT 95.940 5.085 96.260 5.145 ;
        RECT 96.975 5.100 97.265 5.145 ;
        RECT 22.145 4.945 22.435 4.990 ;
        RECT 25.020 4.945 25.340 5.005 ;
        RECT 22.145 4.805 25.340 4.945 ;
        RECT 22.145 4.760 22.435 4.805 ;
        RECT 22.640 4.265 22.960 4.325 ;
        RECT 24.600 4.315 24.740 4.805 ;
        RECT 25.020 4.745 25.340 4.805 ;
        RECT 39.365 4.945 39.655 4.990 ;
        RECT 42.240 4.945 42.560 5.005 ;
        RECT 39.365 4.805 42.560 4.945 ;
        RECT 39.365 4.760 39.655 4.805 ;
        RECT 26.040 4.605 26.360 4.665 ;
        RECT 25.765 4.465 26.360 4.605 ;
        RECT 26.040 4.405 26.360 4.465 ;
        RECT 24.015 4.270 24.305 4.315 ;
        RECT 22.365 4.125 22.960 4.265 ;
        RECT 22.640 4.065 22.960 4.125 ;
        RECT 23.410 4.130 24.305 4.270 ;
        RECT 23.410 3.985 23.550 4.130 ;
        RECT 24.015 4.085 24.305 4.130 ;
        RECT 24.525 4.085 24.815 4.315 ;
        RECT 25.360 4.265 25.680 4.325 ;
        RECT 27.740 4.265 28.060 4.325 ;
        RECT 39.860 4.265 40.180 4.325 ;
        RECT 41.820 4.315 41.960 4.805 ;
        RECT 42.240 4.745 42.560 4.805 ;
        RECT 56.585 4.945 56.875 4.990 ;
        RECT 59.460 4.945 59.780 5.005 ;
        RECT 56.585 4.805 59.780 4.945 ;
        RECT 56.585 4.760 56.875 4.805 ;
        RECT 43.260 4.605 43.580 4.665 ;
        RECT 42.985 4.465 43.580 4.605 ;
        RECT 43.260 4.405 43.580 4.465 ;
        RECT 41.235 4.270 41.525 4.315 ;
        RECT 25.085 4.125 25.680 4.265 ;
        RECT 27.465 4.125 28.060 4.265 ;
        RECT 39.585 4.125 40.180 4.265 ;
        RECT 25.360 4.065 25.680 4.125 ;
        RECT 27.740 4.065 28.060 4.125 ;
        RECT 39.860 4.065 40.180 4.125 ;
        RECT 40.630 4.130 41.525 4.270 ;
        RECT 40.630 3.985 40.770 4.130 ;
        RECT 41.235 4.085 41.525 4.130 ;
        RECT 41.745 4.085 42.035 4.315 ;
        RECT 42.580 4.265 42.900 4.325 ;
        RECT 44.960 4.265 45.280 4.325 ;
        RECT 57.080 4.265 57.400 4.325 ;
        RECT 59.040 4.315 59.180 4.805 ;
        RECT 59.460 4.745 59.780 4.805 ;
        RECT 73.805 4.945 74.095 4.990 ;
        RECT 76.680 4.945 77.000 5.005 ;
        RECT 73.805 4.805 77.000 4.945 ;
        RECT 73.805 4.760 74.095 4.805 ;
        RECT 60.480 4.605 60.800 4.665 ;
        RECT 60.205 4.465 60.800 4.605 ;
        RECT 60.480 4.405 60.800 4.465 ;
        RECT 58.455 4.270 58.745 4.315 ;
        RECT 42.305 4.125 42.900 4.265 ;
        RECT 44.685 4.125 45.280 4.265 ;
        RECT 56.805 4.125 57.400 4.265 ;
        RECT 42.580 4.065 42.900 4.125 ;
        RECT 44.960 4.065 45.280 4.125 ;
        RECT 57.080 4.065 57.400 4.125 ;
        RECT 57.850 4.130 58.745 4.270 ;
        RECT 57.850 3.985 57.990 4.130 ;
        RECT 58.455 4.085 58.745 4.130 ;
        RECT 58.965 4.085 59.255 4.315 ;
        RECT 59.800 4.265 60.120 4.325 ;
        RECT 62.180 4.265 62.500 4.325 ;
        RECT 74.300 4.265 74.620 4.325 ;
        RECT 76.260 4.315 76.400 4.805 ;
        RECT 76.680 4.745 77.000 4.805 ;
        RECT 91.025 4.945 91.315 4.990 ;
        RECT 93.900 4.945 94.220 5.005 ;
        RECT 91.025 4.805 94.220 4.945 ;
        RECT 91.025 4.760 91.315 4.805 ;
        RECT 77.700 4.605 78.020 4.665 ;
        RECT 77.425 4.465 78.020 4.605 ;
        RECT 77.700 4.405 78.020 4.465 ;
        RECT 75.675 4.270 75.965 4.315 ;
        RECT 59.525 4.125 60.120 4.265 ;
        RECT 61.905 4.125 62.500 4.265 ;
        RECT 74.025 4.125 74.620 4.265 ;
        RECT 59.800 4.065 60.120 4.125 ;
        RECT 62.180 4.065 62.500 4.125 ;
        RECT 74.300 4.065 74.620 4.125 ;
        RECT 75.070 4.130 75.965 4.270 ;
        RECT 75.070 3.985 75.210 4.130 ;
        RECT 75.675 4.085 75.965 4.130 ;
        RECT 76.185 4.085 76.475 4.315 ;
        RECT 77.020 4.265 77.340 4.325 ;
        RECT 79.400 4.265 79.720 4.325 ;
        RECT 91.520 4.265 91.840 4.325 ;
        RECT 93.480 4.315 93.620 4.805 ;
        RECT 93.900 4.745 94.220 4.805 ;
        RECT 94.920 4.605 95.240 4.665 ;
        RECT 94.645 4.465 95.240 4.605 ;
        RECT 94.920 4.405 95.240 4.465 ;
        RECT 92.895 4.270 93.185 4.315 ;
        RECT 76.745 4.125 77.340 4.265 ;
        RECT 79.125 4.125 79.720 4.265 ;
        RECT 91.245 4.125 91.840 4.265 ;
        RECT 77.020 4.065 77.340 4.125 ;
        RECT 79.400 4.065 79.720 4.125 ;
        RECT 91.520 4.065 91.840 4.125 ;
        RECT 92.290 4.130 93.185 4.270 ;
        RECT 92.290 3.985 92.430 4.130 ;
        RECT 92.895 4.085 93.185 4.130 ;
        RECT 93.405 4.085 93.695 4.315 ;
        RECT 94.240 4.265 94.560 4.325 ;
        RECT 96.620 4.265 96.940 4.325 ;
        RECT 93.965 4.125 94.560 4.265 ;
        RECT 96.345 4.125 96.940 4.265 ;
        RECT 94.240 4.065 94.560 4.125 ;
        RECT 96.620 4.065 96.940 4.125 ;
        RECT 23.320 3.725 23.640 3.985 ;
        RECT 31.315 3.875 31.635 3.980 ;
        RECT 31.290 3.860 31.635 3.875 ;
        RECT 24.680 3.800 25.000 3.815 ;
        RECT 24.680 3.755 25.185 3.800 ;
        RECT 24.590 3.615 25.185 3.755 ;
        RECT 31.000 3.690 31.635 3.860 ;
        RECT 31.115 3.675 31.635 3.690 ;
        RECT 31.290 3.660 31.635 3.675 ;
        RECT 31.290 3.645 31.580 3.660 ;
        RECT 24.680 3.570 25.185 3.615 ;
        RECT 24.680 3.555 25.000 3.570 ;
        RECT 29.645 3.290 29.970 3.615 ;
        RECT 32.090 3.485 32.440 3.610 ;
        RECT 33.450 3.540 33.740 3.775 ;
        RECT 40.540 3.725 40.860 3.985 ;
        RECT 48.535 3.875 48.855 3.980 ;
        RECT 48.510 3.860 48.855 3.875 ;
        RECT 41.900 3.800 42.220 3.815 ;
        RECT 41.900 3.755 42.405 3.800 ;
        RECT 41.810 3.615 42.405 3.755 ;
        RECT 48.220 3.690 48.855 3.860 ;
        RECT 48.335 3.675 48.855 3.690 ;
        RECT 48.510 3.660 48.855 3.675 ;
        RECT 48.510 3.645 48.800 3.660 ;
        RECT 41.900 3.570 42.405 3.615 ;
        RECT 41.900 3.555 42.220 3.570 ;
        RECT 33.450 3.535 33.680 3.540 ;
        RECT 31.920 3.315 32.440 3.485 ;
        RECT 32.090 3.260 32.440 3.315 ;
        RECT 33.090 3.225 33.325 3.235 ;
        RECT 31.660 3.120 31.950 3.145 ;
        RECT 33.030 3.120 33.370 3.225 ;
        RECT 31.660 2.950 33.370 3.120 ;
        RECT 31.660 2.915 31.950 2.950 ;
        RECT 31.720 2.405 31.890 2.915 ;
        RECT 33.030 2.910 33.370 2.950 ;
        RECT 33.090 2.885 33.325 2.910 ;
        RECT 33.510 2.435 33.680 3.535 ;
        RECT 46.865 3.290 47.190 3.615 ;
        RECT 49.310 3.485 49.660 3.610 ;
        RECT 50.670 3.540 50.960 3.775 ;
        RECT 57.760 3.725 58.080 3.985 ;
        RECT 65.755 3.875 66.075 3.980 ;
        RECT 65.730 3.860 66.075 3.875 ;
        RECT 59.120 3.800 59.440 3.815 ;
        RECT 59.120 3.755 59.625 3.800 ;
        RECT 59.030 3.615 59.625 3.755 ;
        RECT 65.440 3.690 66.075 3.860 ;
        RECT 65.555 3.675 66.075 3.690 ;
        RECT 65.730 3.660 66.075 3.675 ;
        RECT 65.730 3.645 66.020 3.660 ;
        RECT 59.120 3.570 59.625 3.615 ;
        RECT 59.120 3.555 59.440 3.570 ;
        RECT 50.670 3.535 50.900 3.540 ;
        RECT 49.140 3.315 49.660 3.485 ;
        RECT 49.310 3.260 49.660 3.315 ;
        RECT 50.310 3.225 50.545 3.235 ;
        RECT 48.880 3.120 49.170 3.145 ;
        RECT 50.250 3.120 50.590 3.225 ;
        RECT 48.880 2.950 50.590 3.120 ;
        RECT 48.880 2.915 49.170 2.950 ;
        RECT 31.660 2.175 31.950 2.405 ;
        RECT 33.450 2.175 33.745 2.435 ;
        RECT 48.940 2.405 49.110 2.915 ;
        RECT 50.250 2.910 50.590 2.950 ;
        RECT 50.310 2.885 50.545 2.910 ;
        RECT 50.730 2.435 50.900 3.535 ;
        RECT 64.085 3.290 64.410 3.615 ;
        RECT 66.530 3.485 66.880 3.610 ;
        RECT 67.890 3.540 68.180 3.775 ;
        RECT 74.980 3.725 75.300 3.985 ;
        RECT 82.975 3.875 83.295 3.980 ;
        RECT 82.950 3.860 83.295 3.875 ;
        RECT 76.340 3.800 76.660 3.815 ;
        RECT 76.340 3.755 76.845 3.800 ;
        RECT 76.250 3.615 76.845 3.755 ;
        RECT 82.660 3.690 83.295 3.860 ;
        RECT 82.775 3.675 83.295 3.690 ;
        RECT 82.950 3.660 83.295 3.675 ;
        RECT 82.950 3.645 83.240 3.660 ;
        RECT 76.340 3.570 76.845 3.615 ;
        RECT 76.340 3.555 76.660 3.570 ;
        RECT 67.890 3.535 68.120 3.540 ;
        RECT 66.360 3.315 66.880 3.485 ;
        RECT 66.530 3.260 66.880 3.315 ;
        RECT 67.530 3.225 67.765 3.235 ;
        RECT 66.100 3.120 66.390 3.145 ;
        RECT 67.470 3.120 67.810 3.225 ;
        RECT 66.100 2.950 67.810 3.120 ;
        RECT 66.100 2.915 66.390 2.950 ;
        RECT 48.880 2.175 49.170 2.405 ;
        RECT 50.670 2.175 50.965 2.435 ;
        RECT 66.160 2.405 66.330 2.915 ;
        RECT 67.470 2.910 67.810 2.950 ;
        RECT 67.530 2.885 67.765 2.910 ;
        RECT 67.950 2.435 68.120 3.535 ;
        RECT 81.305 3.290 81.630 3.615 ;
        RECT 83.750 3.485 84.100 3.610 ;
        RECT 85.110 3.540 85.400 3.775 ;
        RECT 92.200 3.725 92.520 3.985 ;
        RECT 100.195 3.875 100.515 3.980 ;
        RECT 100.170 3.860 100.515 3.875 ;
        RECT 93.560 3.800 93.880 3.815 ;
        RECT 93.560 3.755 94.065 3.800 ;
        RECT 93.470 3.615 94.065 3.755 ;
        RECT 99.880 3.690 100.515 3.860 ;
        RECT 99.995 3.675 100.515 3.690 ;
        RECT 100.170 3.660 100.515 3.675 ;
        RECT 100.170 3.645 100.460 3.660 ;
        RECT 93.560 3.570 94.065 3.615 ;
        RECT 93.560 3.555 93.880 3.570 ;
        RECT 85.110 3.535 85.340 3.540 ;
        RECT 83.580 3.315 84.100 3.485 ;
        RECT 83.750 3.260 84.100 3.315 ;
        RECT 84.750 3.225 84.985 3.235 ;
        RECT 83.320 3.120 83.610 3.145 ;
        RECT 84.690 3.120 85.030 3.225 ;
        RECT 83.320 2.950 85.030 3.120 ;
        RECT 83.320 2.915 83.610 2.950 ;
        RECT 66.100 2.175 66.390 2.405 ;
        RECT 67.890 2.175 68.185 2.435 ;
        RECT 83.380 2.405 83.550 2.915 ;
        RECT 84.690 2.910 85.030 2.950 ;
        RECT 84.750 2.885 84.985 2.910 ;
        RECT 85.170 2.435 85.340 3.535 ;
        RECT 98.525 3.290 98.850 3.615 ;
        RECT 100.970 3.485 101.320 3.610 ;
        RECT 102.330 3.540 102.620 3.775 ;
        RECT 102.330 3.535 102.560 3.540 ;
        RECT 100.800 3.315 101.320 3.485 ;
        RECT 100.970 3.260 101.320 3.315 ;
        RECT 101.970 3.225 102.205 3.235 ;
        RECT 100.540 3.120 100.830 3.145 ;
        RECT 101.910 3.120 102.250 3.225 ;
        RECT 100.540 2.950 102.250 3.120 ;
        RECT 100.540 2.915 100.830 2.950 ;
        RECT 83.320 2.175 83.610 2.405 ;
        RECT 85.110 2.175 85.405 2.435 ;
        RECT 100.600 2.405 100.770 2.915 ;
        RECT 101.910 2.910 102.250 2.950 ;
        RECT 101.970 2.885 102.205 2.910 ;
        RECT 102.390 2.435 102.560 3.535 ;
        RECT 100.540 2.175 100.830 2.405 ;
        RECT 102.330 2.175 102.625 2.435 ;
      LAYER met2 ;
        RECT 16.245 10.065 103.555 10.235 ;
        RECT 16.245 8.880 16.415 10.065 ;
        RECT 103.385 9.910 103.555 10.065 ;
        RECT 16.565 9.515 16.845 9.620 ;
        RECT 16.565 9.345 17.775 9.515 ;
        RECT 16.565 9.280 16.845 9.345 ;
        RECT 17.605 9.140 17.775 9.345 ;
        RECT 19.940 9.310 20.310 9.680 ;
        RECT 20.465 9.650 31.160 9.820 ;
        RECT 20.465 9.170 20.635 9.650 ;
        RECT 31.000 9.200 31.160 9.650 ;
        RECT 37.160 9.310 37.530 9.680 ;
        RECT 37.685 9.650 48.380 9.820 ;
        RECT 32.115 9.200 32.440 9.265 ;
        RECT 20.415 9.140 20.695 9.170 ;
        RECT 17.605 8.970 20.695 9.140 ;
        RECT 16.190 8.540 16.470 8.880 ;
        RECT 20.415 8.830 20.695 8.970 ;
        RECT 31.000 9.030 32.440 9.200 ;
        RECT 24.700 7.725 24.980 8.095 ;
        RECT 26.070 8.050 26.330 8.095 ;
        RECT 26.040 7.805 26.360 8.050 ;
        RECT 26.070 7.760 26.330 7.805 ;
        RECT 27.770 7.760 28.030 8.095 ;
        RECT 25.710 7.065 25.990 7.435 ;
        RECT 26.130 6.645 26.270 7.760 ;
        RECT 26.750 7.065 27.030 7.435 ;
        RECT 25.450 6.505 26.270 6.645 ;
        RECT 22.670 6.075 22.930 6.395 ;
        RECT 22.730 4.355 22.870 6.075 ;
        RECT 25.450 5.800 25.590 6.505 ;
        RECT 27.090 6.075 27.350 6.395 ;
        RECT 23.340 5.430 23.620 5.800 ;
        RECT 25.380 5.430 25.660 5.800 ;
        RECT 22.670 4.035 22.930 4.355 ;
        RECT 23.410 4.015 23.550 5.430 ;
        RECT 25.030 4.690 25.310 5.060 ;
        RECT 25.450 4.355 25.590 5.430 ;
        RECT 26.400 5.030 26.680 5.400 ;
        RECT 27.150 5.375 27.290 6.075 ;
        RECT 27.090 5.055 27.350 5.375 ;
        RECT 25.390 4.035 25.650 4.355 ;
        RECT 26.060 4.350 26.340 4.720 ;
        RECT 27.830 4.355 27.970 7.760 ;
        RECT 23.350 3.695 23.610 4.015 ;
        RECT 24.700 3.500 24.980 3.870 ;
        RECT 26.130 3.815 26.305 4.350 ;
        RECT 27.770 4.035 28.030 4.355 ;
        RECT 31.000 3.860 31.160 9.030 ;
        RECT 32.115 8.940 32.440 9.030 ;
        RECT 34.505 9.145 34.830 9.270 ;
        RECT 37.685 9.170 37.855 9.650 ;
        RECT 48.220 9.200 48.380 9.650 ;
        RECT 54.380 9.310 54.750 9.680 ;
        RECT 54.905 9.650 65.600 9.820 ;
        RECT 49.335 9.200 49.660 9.265 ;
        RECT 34.505 9.140 35.415 9.145 ;
        RECT 37.635 9.140 37.915 9.170 ;
        RECT 34.505 8.975 37.915 9.140 ;
        RECT 34.505 8.945 34.830 8.975 ;
        RECT 35.415 8.970 37.915 8.975 ;
        RECT 31.315 8.565 31.635 8.890 ;
        RECT 37.635 8.830 37.915 8.970 ;
        RECT 48.220 9.030 49.660 9.200 ;
        RECT 31.345 8.330 31.515 8.565 ;
        RECT 31.345 8.155 31.520 8.330 ;
        RECT 31.345 7.980 32.320 8.155 ;
        RECT 31.315 3.860 31.635 3.980 ;
        RECT 26.130 3.640 29.350 3.815 ;
        RECT 31.000 3.690 31.635 3.860 ;
        RECT 31.315 3.660 31.635 3.690 ;
        RECT 29.175 3.490 29.350 3.640 ;
        RECT 29.645 3.490 29.970 3.615 ;
        RECT 32.145 3.610 32.320 7.980 ;
        RECT 41.920 7.725 42.200 8.095 ;
        RECT 43.290 8.050 43.550 8.095 ;
        RECT 43.260 7.805 43.580 8.050 ;
        RECT 43.290 7.760 43.550 7.805 ;
        RECT 44.990 7.760 45.250 8.095 ;
        RECT 42.930 7.065 43.210 7.435 ;
        RECT 43.350 6.645 43.490 7.760 ;
        RECT 43.970 7.065 44.250 7.435 ;
        RECT 42.670 6.505 43.490 6.645 ;
        RECT 39.890 6.075 40.150 6.395 ;
        RECT 39.950 4.355 40.090 6.075 ;
        RECT 42.670 5.800 42.810 6.505 ;
        RECT 44.310 6.075 44.570 6.395 ;
        RECT 40.560 5.430 40.840 5.800 ;
        RECT 42.600 5.430 42.880 5.800 ;
        RECT 39.890 4.035 40.150 4.355 ;
        RECT 40.630 4.015 40.770 5.430 ;
        RECT 42.250 4.690 42.530 5.060 ;
        RECT 42.670 4.355 42.810 5.430 ;
        RECT 43.620 5.030 43.900 5.400 ;
        RECT 44.370 5.375 44.510 6.075 ;
        RECT 44.310 5.055 44.570 5.375 ;
        RECT 42.610 4.035 42.870 4.355 ;
        RECT 43.280 4.350 43.560 4.720 ;
        RECT 45.050 4.355 45.190 7.760 ;
        RECT 40.570 3.695 40.830 4.015 ;
        RECT 32.090 3.490 32.440 3.610 ;
        RECT 41.920 3.500 42.200 3.870 ;
        RECT 43.350 3.815 43.525 4.350 ;
        RECT 44.990 4.035 45.250 4.355 ;
        RECT 48.220 3.860 48.380 9.030 ;
        RECT 49.335 8.940 49.660 9.030 ;
        RECT 51.725 9.145 52.050 9.270 ;
        RECT 54.905 9.170 55.075 9.650 ;
        RECT 65.440 9.200 65.600 9.650 ;
        RECT 71.600 9.310 71.970 9.680 ;
        RECT 72.125 9.650 82.820 9.820 ;
        RECT 66.555 9.200 66.880 9.265 ;
        RECT 51.725 9.140 52.650 9.145 ;
        RECT 54.855 9.140 55.135 9.170 ;
        RECT 51.725 8.975 55.145 9.140 ;
        RECT 51.725 8.945 52.050 8.975 ;
        RECT 53.675 8.970 55.145 8.975 ;
        RECT 65.440 9.030 66.880 9.200 ;
        RECT 48.535 8.565 48.855 8.890 ;
        RECT 54.855 8.830 55.135 8.970 ;
        RECT 48.565 8.330 48.735 8.565 ;
        RECT 48.565 8.155 48.740 8.330 ;
        RECT 48.565 7.980 49.540 8.155 ;
        RECT 48.535 3.860 48.855 3.980 ;
        RECT 43.350 3.640 46.570 3.815 ;
        RECT 48.220 3.690 48.855 3.860 ;
        RECT 48.535 3.660 48.855 3.690 ;
        RECT 29.175 3.320 32.440 3.490 ;
        RECT 46.395 3.490 46.570 3.640 ;
        RECT 46.865 3.490 47.190 3.615 ;
        RECT 49.365 3.610 49.540 7.980 ;
        RECT 59.140 7.725 59.420 8.095 ;
        RECT 60.510 8.050 60.770 8.095 ;
        RECT 60.480 7.805 60.800 8.050 ;
        RECT 60.510 7.760 60.770 7.805 ;
        RECT 62.210 7.760 62.470 8.095 ;
        RECT 60.150 7.065 60.430 7.435 ;
        RECT 60.570 6.645 60.710 7.760 ;
        RECT 61.190 7.065 61.470 7.435 ;
        RECT 59.890 6.505 60.710 6.645 ;
        RECT 57.110 6.075 57.370 6.395 ;
        RECT 57.170 4.355 57.310 6.075 ;
        RECT 59.890 5.800 60.030 6.505 ;
        RECT 61.530 6.075 61.790 6.395 ;
        RECT 57.780 5.430 58.060 5.800 ;
        RECT 59.820 5.430 60.100 5.800 ;
        RECT 57.110 4.035 57.370 4.355 ;
        RECT 57.850 4.015 57.990 5.430 ;
        RECT 59.470 4.690 59.750 5.060 ;
        RECT 59.890 4.355 60.030 5.430 ;
        RECT 60.840 5.030 61.120 5.400 ;
        RECT 61.590 5.375 61.730 6.075 ;
        RECT 61.530 5.055 61.790 5.375 ;
        RECT 59.830 4.035 60.090 4.355 ;
        RECT 60.500 4.350 60.780 4.720 ;
        RECT 62.270 4.355 62.410 7.760 ;
        RECT 57.790 3.695 58.050 4.015 ;
        RECT 49.310 3.490 49.660 3.610 ;
        RECT 59.140 3.500 59.420 3.870 ;
        RECT 60.570 3.815 60.745 4.350 ;
        RECT 62.210 4.035 62.470 4.355 ;
        RECT 65.440 3.860 65.600 9.030 ;
        RECT 66.555 8.940 66.880 9.030 ;
        RECT 68.945 9.145 69.270 9.270 ;
        RECT 72.125 9.170 72.295 9.650 ;
        RECT 82.660 9.200 82.820 9.650 ;
        RECT 88.820 9.310 89.190 9.680 ;
        RECT 89.345 9.650 100.040 9.820 ;
        RECT 83.775 9.200 84.100 9.265 ;
        RECT 68.945 9.140 69.890 9.145 ;
        RECT 72.075 9.140 72.355 9.170 ;
        RECT 68.945 8.975 72.355 9.140 ;
        RECT 68.945 8.945 69.270 8.975 ;
        RECT 69.890 8.970 72.355 8.975 ;
        RECT 65.755 8.565 66.075 8.890 ;
        RECT 72.075 8.830 72.355 8.970 ;
        RECT 82.660 9.030 84.100 9.200 ;
        RECT 65.785 8.330 65.955 8.565 ;
        RECT 65.785 8.155 65.960 8.330 ;
        RECT 65.785 7.980 66.760 8.155 ;
        RECT 65.755 3.860 66.075 3.980 ;
        RECT 60.570 3.640 63.790 3.815 ;
        RECT 65.440 3.690 66.075 3.860 ;
        RECT 65.755 3.660 66.075 3.690 ;
        RECT 46.395 3.320 49.660 3.490 ;
        RECT 63.615 3.490 63.790 3.640 ;
        RECT 64.085 3.490 64.410 3.615 ;
        RECT 66.585 3.610 66.760 7.980 ;
        RECT 76.360 7.725 76.640 8.095 ;
        RECT 77.730 8.050 77.990 8.095 ;
        RECT 77.700 7.805 78.020 8.050 ;
        RECT 77.730 7.760 77.990 7.805 ;
        RECT 79.430 7.760 79.690 8.095 ;
        RECT 77.370 7.065 77.650 7.435 ;
        RECT 77.790 6.645 77.930 7.760 ;
        RECT 78.410 7.065 78.690 7.435 ;
        RECT 77.110 6.505 77.930 6.645 ;
        RECT 74.330 6.075 74.590 6.395 ;
        RECT 74.390 4.355 74.530 6.075 ;
        RECT 77.110 5.800 77.250 6.505 ;
        RECT 78.750 6.075 79.010 6.395 ;
        RECT 75.000 5.430 75.280 5.800 ;
        RECT 77.040 5.430 77.320 5.800 ;
        RECT 74.330 4.035 74.590 4.355 ;
        RECT 75.070 4.015 75.210 5.430 ;
        RECT 76.690 4.690 76.970 5.060 ;
        RECT 77.110 4.355 77.250 5.430 ;
        RECT 78.060 5.030 78.340 5.400 ;
        RECT 78.810 5.375 78.950 6.075 ;
        RECT 78.750 5.055 79.010 5.375 ;
        RECT 77.050 4.035 77.310 4.355 ;
        RECT 77.720 4.350 78.000 4.720 ;
        RECT 79.490 4.355 79.630 7.760 ;
        RECT 75.010 3.695 75.270 4.015 ;
        RECT 66.530 3.490 66.880 3.610 ;
        RECT 76.360 3.500 76.640 3.870 ;
        RECT 77.790 3.815 77.965 4.350 ;
        RECT 79.430 4.035 79.690 4.355 ;
        RECT 82.660 3.860 82.820 9.030 ;
        RECT 83.775 8.940 84.100 9.030 ;
        RECT 86.165 9.145 86.490 9.270 ;
        RECT 89.345 9.170 89.515 9.650 ;
        RECT 99.880 9.200 100.040 9.650 ;
        RECT 103.350 9.585 103.675 9.910 ;
        RECT 100.995 9.200 101.320 9.265 ;
        RECT 86.165 9.140 87.155 9.145 ;
        RECT 89.295 9.140 89.575 9.170 ;
        RECT 86.165 8.975 89.575 9.140 ;
        RECT 86.165 8.945 86.490 8.975 ;
        RECT 87.155 8.970 89.575 8.975 ;
        RECT 82.975 8.565 83.295 8.890 ;
        RECT 89.295 8.830 89.575 8.970 ;
        RECT 99.880 9.030 101.320 9.200 ;
        RECT 83.005 8.330 83.175 8.565 ;
        RECT 83.005 8.155 83.180 8.330 ;
        RECT 83.005 7.980 83.980 8.155 ;
        RECT 82.975 3.860 83.295 3.980 ;
        RECT 77.790 3.640 81.010 3.815 ;
        RECT 82.660 3.690 83.295 3.860 ;
        RECT 82.975 3.660 83.295 3.690 ;
        RECT 63.615 3.320 66.880 3.490 ;
        RECT 80.835 3.490 81.010 3.640 ;
        RECT 81.305 3.490 81.630 3.615 ;
        RECT 83.805 3.610 83.980 7.980 ;
        RECT 93.580 7.725 93.860 8.095 ;
        RECT 94.950 8.050 95.210 8.095 ;
        RECT 94.920 7.805 95.240 8.050 ;
        RECT 94.950 7.760 95.210 7.805 ;
        RECT 96.650 7.760 96.910 8.095 ;
        RECT 94.590 7.065 94.870 7.435 ;
        RECT 95.010 6.645 95.150 7.760 ;
        RECT 95.630 7.065 95.910 7.435 ;
        RECT 94.330 6.505 95.150 6.645 ;
        RECT 91.550 6.075 91.810 6.395 ;
        RECT 91.610 4.355 91.750 6.075 ;
        RECT 94.330 5.800 94.470 6.505 ;
        RECT 95.970 6.075 96.230 6.395 ;
        RECT 92.220 5.430 92.500 5.800 ;
        RECT 94.260 5.430 94.540 5.800 ;
        RECT 91.550 4.035 91.810 4.355 ;
        RECT 92.290 4.015 92.430 5.430 ;
        RECT 93.910 4.690 94.190 5.060 ;
        RECT 94.330 4.355 94.470 5.430 ;
        RECT 95.280 5.030 95.560 5.400 ;
        RECT 96.030 5.375 96.170 6.075 ;
        RECT 95.970 5.055 96.230 5.375 ;
        RECT 94.270 4.035 94.530 4.355 ;
        RECT 94.940 4.350 95.220 4.720 ;
        RECT 96.710 4.355 96.850 7.760 ;
        RECT 92.230 3.695 92.490 4.015 ;
        RECT 83.750 3.490 84.100 3.610 ;
        RECT 93.580 3.500 93.860 3.870 ;
        RECT 95.010 3.815 95.185 4.350 ;
        RECT 96.650 4.035 96.910 4.355 ;
        RECT 99.880 3.860 100.040 9.030 ;
        RECT 100.995 8.940 101.320 9.030 ;
        RECT 100.195 8.565 100.515 8.890 ;
        RECT 100.225 8.330 100.395 8.565 ;
        RECT 100.225 8.155 100.400 8.330 ;
        RECT 100.225 7.980 101.200 8.155 ;
        RECT 100.195 3.860 100.515 3.980 ;
        RECT 95.010 3.640 98.230 3.815 ;
        RECT 99.880 3.690 100.515 3.860 ;
        RECT 100.195 3.660 100.515 3.690 ;
        RECT 80.835 3.320 84.100 3.490 ;
        RECT 98.055 3.490 98.230 3.640 ;
        RECT 98.525 3.490 98.850 3.615 ;
        RECT 101.025 3.610 101.200 7.980 ;
        RECT 100.970 3.490 101.320 3.610 ;
        RECT 98.055 3.320 101.320 3.490 ;
        RECT 29.645 3.290 29.970 3.320 ;
        RECT 32.090 3.260 32.440 3.320 ;
        RECT 46.865 3.290 47.190 3.320 ;
        RECT 49.310 3.260 49.660 3.320 ;
        RECT 64.085 3.290 64.410 3.320 ;
        RECT 66.530 3.260 66.880 3.320 ;
        RECT 81.305 3.290 81.630 3.320 ;
        RECT 83.750 3.260 84.100 3.320 ;
        RECT 98.525 3.290 98.850 3.320 ;
        RECT 100.970 3.260 101.320 3.320 ;
      LAYER met3 ;
        RECT 19.940 9.620 20.310 9.680 ;
        RECT 37.160 9.620 37.530 9.680 ;
        RECT 54.380 9.620 54.750 9.680 ;
        RECT 71.600 9.620 71.970 9.680 ;
        RECT 88.820 9.620 89.190 9.680 ;
        RECT 19.940 9.320 27.090 9.620 ;
        RECT 19.940 9.310 20.310 9.320 ;
        RECT 24.705 8.090 25.005 9.320 ;
        RECT 24.205 7.790 25.005 8.090 ;
        RECT 24.585 7.745 25.005 7.790 ;
        RECT 24.585 7.720 24.885 7.745 ;
        RECT 25.735 7.430 26.035 9.320 ;
        RECT 26.790 7.465 27.090 9.320 ;
        RECT 37.160 9.320 44.310 9.620 ;
        RECT 37.160 9.310 37.530 9.320 ;
        RECT 41.925 8.090 42.225 9.320 ;
        RECT 41.425 7.790 42.225 8.090 ;
        RECT 41.805 7.745 42.225 7.790 ;
        RECT 41.805 7.720 42.105 7.745 ;
        RECT 25.695 7.415 26.035 7.430 ;
        RECT 25.685 7.400 26.035 7.415 ;
        RECT 25.215 7.100 26.035 7.400 ;
        RECT 26.715 7.400 27.090 7.465 ;
        RECT 42.955 7.430 43.255 9.320 ;
        RECT 44.010 7.465 44.310 9.320 ;
        RECT 54.380 9.320 61.530 9.620 ;
        RECT 54.380 9.310 54.750 9.320 ;
        RECT 59.145 8.090 59.445 9.320 ;
        RECT 58.645 7.790 59.445 8.090 ;
        RECT 59.025 7.745 59.445 7.790 ;
        RECT 59.025 7.720 59.325 7.745 ;
        RECT 42.915 7.415 43.255 7.430 ;
        RECT 42.905 7.400 43.255 7.415 ;
        RECT 26.715 7.100 27.525 7.400 ;
        RECT 42.435 7.100 43.255 7.400 ;
        RECT 43.935 7.400 44.310 7.465 ;
        RECT 60.175 7.430 60.475 9.320 ;
        RECT 61.230 7.465 61.530 9.320 ;
        RECT 71.600 9.320 78.750 9.620 ;
        RECT 71.600 9.310 71.970 9.320 ;
        RECT 76.365 8.090 76.665 9.320 ;
        RECT 75.865 7.790 76.665 8.090 ;
        RECT 76.245 7.745 76.665 7.790 ;
        RECT 76.245 7.720 76.545 7.745 ;
        RECT 60.135 7.415 60.475 7.430 ;
        RECT 60.125 7.400 60.475 7.415 ;
        RECT 43.935 7.100 44.745 7.400 ;
        RECT 59.655 7.100 60.475 7.400 ;
        RECT 61.155 7.400 61.530 7.465 ;
        RECT 77.395 7.430 77.695 9.320 ;
        RECT 78.450 7.465 78.750 9.320 ;
        RECT 88.820 9.320 95.970 9.620 ;
        RECT 88.820 9.310 89.190 9.320 ;
        RECT 93.585 8.090 93.885 9.320 ;
        RECT 93.085 7.790 93.885 8.090 ;
        RECT 93.465 7.745 93.885 7.790 ;
        RECT 93.465 7.720 93.765 7.745 ;
        RECT 77.355 7.415 77.695 7.430 ;
        RECT 77.345 7.400 77.695 7.415 ;
        RECT 61.155 7.100 61.965 7.400 ;
        RECT 76.875 7.100 77.695 7.400 ;
        RECT 78.375 7.400 78.750 7.465 ;
        RECT 94.615 7.430 94.915 9.320 ;
        RECT 95.670 7.465 95.970 9.320 ;
        RECT 94.575 7.415 94.915 7.430 ;
        RECT 94.565 7.400 94.915 7.415 ;
        RECT 78.375 7.100 79.185 7.400 ;
        RECT 94.095 7.100 94.915 7.400 ;
        RECT 95.595 7.400 95.970 7.465 ;
        RECT 95.595 7.100 96.405 7.400 ;
        RECT 25.685 7.085 26.035 7.100 ;
        RECT 26.725 7.085 27.080 7.100 ;
        RECT 42.905 7.085 43.255 7.100 ;
        RECT 43.945 7.085 44.300 7.100 ;
        RECT 60.125 7.085 60.475 7.100 ;
        RECT 61.165 7.085 61.520 7.100 ;
        RECT 77.345 7.085 77.695 7.100 ;
        RECT 78.385 7.085 78.740 7.100 ;
        RECT 94.565 7.085 94.915 7.100 ;
        RECT 95.605 7.085 95.960 7.100 ;
        RECT 25.695 7.080 26.035 7.085 ;
        RECT 25.710 7.040 26.010 7.080 ;
        RECT 26.780 7.060 27.080 7.085 ;
        RECT 42.915 7.080 43.255 7.085 ;
        RECT 42.930 7.040 43.230 7.080 ;
        RECT 44.000 7.060 44.300 7.085 ;
        RECT 60.135 7.080 60.475 7.085 ;
        RECT 60.150 7.040 60.450 7.080 ;
        RECT 61.220 7.060 61.520 7.085 ;
        RECT 77.355 7.080 77.695 7.085 ;
        RECT 77.370 7.040 77.670 7.080 ;
        RECT 78.440 7.060 78.740 7.085 ;
        RECT 94.575 7.080 94.915 7.085 ;
        RECT 94.590 7.040 94.890 7.080 ;
        RECT 95.660 7.060 95.960 7.085 ;
        RECT 23.315 5.765 23.645 5.780 ;
        RECT 25.355 5.765 25.685 5.780 ;
        RECT 23.315 5.465 25.685 5.765 ;
        RECT 23.315 5.450 23.645 5.465 ;
        RECT 25.355 5.450 25.685 5.465 ;
        RECT 40.535 5.765 40.865 5.780 ;
        RECT 42.575 5.765 42.905 5.780 ;
        RECT 40.535 5.465 42.905 5.765 ;
        RECT 40.535 5.450 40.865 5.465 ;
        RECT 42.575 5.450 42.905 5.465 ;
        RECT 57.755 5.765 58.085 5.780 ;
        RECT 59.795 5.765 60.125 5.780 ;
        RECT 57.755 5.465 60.125 5.765 ;
        RECT 57.755 5.450 58.085 5.465 ;
        RECT 59.795 5.450 60.125 5.465 ;
        RECT 74.975 5.765 75.305 5.780 ;
        RECT 77.015 5.765 77.345 5.780 ;
        RECT 74.975 5.465 77.345 5.765 ;
        RECT 74.975 5.450 75.305 5.465 ;
        RECT 77.015 5.450 77.345 5.465 ;
        RECT 92.195 5.765 92.525 5.780 ;
        RECT 94.235 5.765 94.565 5.780 ;
        RECT 92.195 5.465 94.565 5.765 ;
        RECT 92.195 5.450 92.525 5.465 ;
        RECT 94.235 5.450 94.565 5.465 ;
        RECT 26.375 5.365 26.705 5.380 ;
        RECT 43.595 5.365 43.925 5.380 ;
        RECT 60.815 5.365 61.145 5.380 ;
        RECT 78.035 5.365 78.365 5.380 ;
        RECT 95.255 5.365 95.585 5.380 ;
        RECT 26.375 5.065 27.175 5.365 ;
        RECT 43.595 5.065 44.395 5.365 ;
        RECT 60.815 5.065 61.615 5.365 ;
        RECT 78.035 5.065 78.835 5.365 ;
        RECT 95.255 5.065 96.055 5.365 ;
        RECT 26.375 5.050 26.705 5.065 ;
        RECT 43.595 5.050 43.925 5.065 ;
        RECT 60.815 5.050 61.145 5.065 ;
        RECT 78.035 5.050 78.365 5.065 ;
        RECT 95.255 5.050 95.585 5.065 ;
        RECT 25.005 5.025 25.335 5.040 ;
        RECT 24.545 4.725 25.345 5.025 ;
        RECT 26.390 5.020 26.690 5.050 ;
        RECT 42.225 5.025 42.555 5.040 ;
        RECT 41.765 4.725 42.565 5.025 ;
        RECT 43.610 5.020 43.910 5.050 ;
        RECT 59.445 5.025 59.775 5.040 ;
        RECT 58.985 4.725 59.785 5.025 ;
        RECT 60.830 5.020 61.130 5.050 ;
        RECT 76.665 5.025 76.995 5.040 ;
        RECT 76.205 4.725 77.005 5.025 ;
        RECT 78.050 5.020 78.350 5.050 ;
        RECT 93.885 5.025 94.215 5.040 ;
        RECT 93.425 4.725 94.225 5.025 ;
        RECT 95.270 5.020 95.570 5.050 ;
        RECT 25.005 4.710 25.335 4.725 ;
        RECT 42.225 4.710 42.555 4.725 ;
        RECT 59.445 4.710 59.775 4.725 ;
        RECT 76.665 4.710 76.995 4.725 ;
        RECT 93.885 4.710 94.215 4.725 ;
        RECT 26.035 4.685 26.365 4.700 ;
        RECT 43.255 4.685 43.585 4.700 ;
        RECT 60.475 4.685 60.805 4.700 ;
        RECT 77.695 4.685 78.025 4.700 ;
        RECT 94.915 4.685 95.245 4.700 ;
        RECT 26.035 4.385 26.835 4.685 ;
        RECT 43.255 4.385 44.055 4.685 ;
        RECT 60.475 4.385 61.275 4.685 ;
        RECT 77.695 4.385 78.495 4.685 ;
        RECT 94.915 4.385 95.715 4.685 ;
        RECT 26.035 4.370 26.420 4.385 ;
        RECT 43.255 4.370 43.640 4.385 ;
        RECT 60.475 4.370 60.860 4.385 ;
        RECT 77.695 4.370 78.080 4.385 ;
        RECT 94.915 4.370 95.300 4.385 ;
        RECT 26.120 4.360 26.420 4.370 ;
        RECT 43.340 4.360 43.640 4.370 ;
        RECT 60.560 4.360 60.860 4.370 ;
        RECT 77.780 4.360 78.080 4.370 ;
        RECT 95.000 4.360 95.300 4.370 ;
        RECT 24.675 3.835 25.005 3.850 ;
        RECT 41.895 3.835 42.225 3.850 ;
        RECT 59.115 3.835 59.445 3.850 ;
        RECT 76.335 3.835 76.665 3.850 ;
        RECT 93.555 3.835 93.885 3.850 ;
        RECT 24.205 3.535 25.005 3.835 ;
        RECT 41.425 3.535 42.225 3.835 ;
        RECT 58.645 3.535 59.445 3.835 ;
        RECT 75.865 3.535 76.665 3.835 ;
        RECT 93.085 3.535 93.885 3.835 ;
        RECT 24.665 3.530 25.005 3.535 ;
        RECT 41.885 3.530 42.225 3.535 ;
        RECT 59.105 3.530 59.445 3.535 ;
        RECT 76.325 3.530 76.665 3.535 ;
        RECT 93.545 3.530 93.885 3.535 ;
        RECT 24.675 3.520 25.005 3.530 ;
        RECT 41.895 3.520 42.225 3.530 ;
        RECT 59.115 3.520 59.445 3.530 ;
        RECT 76.335 3.520 76.665 3.530 ;
        RECT 93.555 3.520 93.885 3.530 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r1
MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r1
  CLASS BLOCK ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ea_8_b0r1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 99.430 BY 12.460 ;
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 23.810 8.235 23.980 9.505 ;
        RECT 29.425 8.235 29.595 9.505 ;
        RECT 29.425 2.955 29.595 4.225 ;
      LAYER met1 ;
        RECT 23.735 8.405 24.055 8.465 ;
        RECT 29.345 8.405 29.685 8.475 ;
        RECT 23.735 8.375 24.210 8.405 ;
        RECT 29.345 8.400 29.825 8.405 ;
        RECT 29.330 8.375 29.825 8.400 ;
        RECT 23.735 8.235 29.825 8.375 ;
        RECT 23.735 8.205 29.685 8.235 ;
        RECT 23.735 8.175 24.055 8.205 ;
        RECT 29.345 8.125 29.685 8.205 ;
        RECT 29.355 4.225 29.695 4.370 ;
        RECT 29.355 4.055 29.825 4.225 ;
        RECT 29.355 4.015 29.695 4.055 ;
      LAYER met2 ;
        RECT 29.345 8.125 29.685 8.475 ;
        RECT 29.430 4.370 29.600 8.125 ;
        RECT 29.355 4.020 29.695 4.370 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 40.135 8.235 40.305 9.505 ;
        RECT 45.750 8.235 45.920 9.505 ;
        RECT 45.750 2.955 45.920 4.225 ;
      LAYER met1 ;
        RECT 40.035 8.405 40.405 8.505 ;
        RECT 45.670 8.405 46.010 8.475 ;
        RECT 40.035 8.375 40.535 8.405 ;
        RECT 45.670 8.400 46.150 8.405 ;
        RECT 45.655 8.375 46.150 8.400 ;
        RECT 40.035 8.235 46.150 8.375 ;
        RECT 40.035 8.205 46.010 8.235 ;
        RECT 40.035 8.135 40.405 8.205 ;
        RECT 45.670 8.125 46.010 8.205 ;
        RECT 45.680 4.225 46.020 4.370 ;
        RECT 45.680 4.055 46.150 4.225 ;
        RECT 45.680 4.015 46.020 4.055 ;
      LAYER met2 ;
        RECT 40.035 8.135 40.405 8.505 ;
        RECT 45.670 8.125 46.010 8.475 ;
        RECT 45.755 4.370 45.925 8.125 ;
        RECT 45.680 4.020 46.020 4.370 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 56.460 8.235 56.630 9.505 ;
        RECT 62.075 8.235 62.245 9.505 ;
        RECT 62.075 2.955 62.245 4.225 ;
      LAYER met1 ;
        RECT 56.385 8.405 56.705 8.465 ;
        RECT 61.995 8.405 62.335 8.475 ;
        RECT 56.385 8.375 56.860 8.405 ;
        RECT 61.995 8.400 62.475 8.405 ;
        RECT 61.980 8.375 62.475 8.400 ;
        RECT 56.385 8.235 62.475 8.375 ;
        RECT 56.385 8.205 62.335 8.235 ;
        RECT 56.385 8.175 56.705 8.205 ;
        RECT 61.995 8.125 62.335 8.205 ;
        RECT 62.005 4.225 62.345 4.370 ;
        RECT 62.005 4.055 62.475 4.225 ;
        RECT 62.005 4.015 62.345 4.055 ;
      LAYER met2 ;
        RECT 61.995 8.125 62.335 8.475 ;
        RECT 62.080 4.370 62.250 8.125 ;
        RECT 62.005 4.020 62.345 4.370 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 72.785 8.235 72.955 9.505 ;
        RECT 78.400 8.235 78.570 9.505 ;
        RECT 78.400 2.955 78.570 4.225 ;
      LAYER met1 ;
        RECT 72.710 8.405 73.030 8.465 ;
        RECT 78.320 8.405 78.660 8.475 ;
        RECT 72.710 8.375 73.185 8.405 ;
        RECT 78.320 8.400 78.800 8.405 ;
        RECT 78.305 8.375 78.800 8.400 ;
        RECT 72.710 8.235 78.800 8.375 ;
        RECT 72.710 8.205 78.660 8.235 ;
        RECT 72.710 8.175 73.030 8.205 ;
        RECT 78.320 8.125 78.660 8.205 ;
        RECT 78.330 4.225 78.670 4.370 ;
        RECT 78.330 4.055 78.800 4.225 ;
        RECT 78.330 4.015 78.670 4.055 ;
      LAYER met2 ;
        RECT 78.320 8.125 78.660 8.475 ;
        RECT 78.405 4.370 78.575 8.125 ;
        RECT 78.330 4.020 78.670 4.370 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 89.110 8.235 89.280 9.505 ;
        RECT 94.725 8.235 94.895 9.505 ;
        RECT 94.725 2.955 94.895 4.225 ;
      LAYER met1 ;
        RECT 89.035 8.405 89.355 8.465 ;
        RECT 94.645 8.405 94.985 8.475 ;
        RECT 89.035 8.375 89.510 8.405 ;
        RECT 94.645 8.400 95.125 8.405 ;
        RECT 94.630 8.375 95.125 8.400 ;
        RECT 89.035 8.235 95.125 8.375 ;
        RECT 89.035 8.205 94.985 8.235 ;
        RECT 89.035 8.175 89.355 8.205 ;
        RECT 94.645 8.125 94.985 8.205 ;
        RECT 94.655 4.225 94.995 4.370 ;
        RECT 94.655 4.055 95.125 4.225 ;
        RECT 94.655 4.015 94.995 4.055 ;
      LAYER met2 ;
        RECT 94.645 8.125 94.985 8.475 ;
        RECT 94.730 4.370 94.900 8.125 ;
        RECT 94.655 4.020 94.995 4.370 ;
    END
  END s5
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 33.580 4.015 33.755 5.160 ;
        RECT 33.580 3.580 33.750 4.015 ;
        RECT 33.585 1.870 33.755 2.380 ;
      LAYER met1 ;
        RECT 33.520 3.545 33.810 3.780 ;
        RECT 33.520 3.540 33.750 3.545 ;
        RECT 33.580 2.440 33.750 3.540 ;
        RECT 33.520 2.180 33.815 2.440 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 49.905 4.015 50.080 5.160 ;
        RECT 49.905 3.580 50.075 4.015 ;
        RECT 49.910 1.870 50.080 2.380 ;
      LAYER met1 ;
        RECT 49.845 3.545 50.135 3.780 ;
        RECT 49.845 3.540 50.075 3.545 ;
        RECT 49.905 2.440 50.075 3.540 ;
        RECT 49.845 2.180 50.140 2.440 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 66.230 4.015 66.405 5.160 ;
        RECT 66.230 3.580 66.400 4.015 ;
        RECT 66.235 1.870 66.405 2.380 ;
      LAYER met1 ;
        RECT 66.170 3.545 66.460 3.780 ;
        RECT 66.170 3.540 66.400 3.545 ;
        RECT 66.230 2.440 66.400 3.540 ;
        RECT 66.170 2.180 66.465 2.440 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 82.555 4.015 82.730 5.160 ;
        RECT 82.555 3.580 82.725 4.015 ;
        RECT 82.560 1.870 82.730 2.380 ;
      LAYER met1 ;
        RECT 82.495 3.545 82.785 3.780 ;
        RECT 82.495 3.540 82.725 3.545 ;
        RECT 82.555 2.440 82.725 3.540 ;
        RECT 82.495 2.180 82.790 2.440 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 98.880 4.015 99.055 5.160 ;
        RECT 98.880 3.580 99.050 4.015 ;
        RECT 98.885 1.870 99.055 2.380 ;
      LAYER met1 ;
        RECT 98.820 3.545 99.110 3.780 ;
        RECT 98.820 3.540 99.050 3.545 ;
        RECT 98.880 2.440 99.050 3.540 ;
        RECT 98.820 2.180 99.115 2.440 ;
    END
  END X5_Y1
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 15.230 8.235 15.400 9.505 ;
      LAYER met1 ;
        RECT 15.170 8.430 15.460 8.435 ;
        RECT 15.170 8.405 15.465 8.430 ;
        RECT 15.170 8.235 15.630 8.405 ;
        RECT 15.170 8.205 15.465 8.235 ;
        RECT 15.175 8.200 15.465 8.205 ;
    END
  END start
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.050 10.860 99.430 12.460 ;
        RECT 15.220 10.235 15.390 10.860 ;
        RECT 23.800 10.235 23.970 10.860 ;
        RECT 24.755 10.315 24.925 10.595 ;
        RECT 24.755 10.145 24.985 10.315 ;
        RECT 29.415 10.235 29.585 10.860 ;
        RECT 32.160 10.235 32.330 10.860 ;
        RECT 33.155 10.230 33.325 10.860 ;
        RECT 40.125 10.235 40.295 10.860 ;
        RECT 41.080 10.315 41.250 10.595 ;
        RECT 41.080 10.145 41.310 10.315 ;
        RECT 45.740 10.235 45.910 10.860 ;
        RECT 48.485 10.235 48.655 10.860 ;
        RECT 49.480 10.230 49.650 10.860 ;
        RECT 56.450 10.235 56.620 10.860 ;
        RECT 57.405 10.315 57.575 10.595 ;
        RECT 57.405 10.145 57.635 10.315 ;
        RECT 62.065 10.235 62.235 10.860 ;
        RECT 64.810 10.235 64.980 10.860 ;
        RECT 65.805 10.230 65.975 10.860 ;
        RECT 72.775 10.235 72.945 10.860 ;
        RECT 73.730 10.315 73.900 10.595 ;
        RECT 73.730 10.145 73.960 10.315 ;
        RECT 78.390 10.235 78.560 10.860 ;
        RECT 81.135 10.235 81.305 10.860 ;
        RECT 82.130 10.230 82.300 10.860 ;
        RECT 89.100 10.235 89.270 10.860 ;
        RECT 90.055 10.315 90.225 10.595 ;
        RECT 90.055 10.145 90.285 10.315 ;
        RECT 94.715 10.235 94.885 10.860 ;
        RECT 97.460 10.235 97.630 10.860 ;
        RECT 98.455 10.230 98.625 10.860 ;
        RECT 24.815 8.535 24.985 10.145 ;
        RECT 41.140 8.535 41.310 10.145 ;
        RECT 57.465 8.535 57.635 10.145 ;
        RECT 73.790 8.535 73.960 10.145 ;
        RECT 90.115 8.535 90.285 10.145 ;
        RECT 24.755 8.365 24.985 8.535 ;
        RECT 41.080 8.365 41.310 8.535 ;
        RECT 57.405 8.365 57.635 8.535 ;
        RECT 73.730 8.365 73.960 8.535 ;
        RECT 90.055 8.365 90.285 8.535 ;
        RECT 24.755 7.305 24.925 8.365 ;
        RECT 41.080 7.305 41.250 8.365 ;
        RECT 57.405 7.305 57.575 8.365 ;
        RECT 73.730 7.305 73.900 8.365 ;
        RECT 90.055 7.305 90.225 8.365 ;
      LAYER met1 ;
        RECT 0.050 10.860 99.430 12.460 ;
        RECT 24.375 8.785 24.550 10.860 ;
        RECT 24.755 8.785 25.045 8.815 ;
        RECT 24.375 8.600 25.045 8.785 ;
        RECT 40.700 8.785 40.875 10.860 ;
        RECT 41.080 8.785 41.370 8.815 ;
        RECT 40.700 8.600 41.370 8.785 ;
        RECT 57.025 8.785 57.200 10.860 ;
        RECT 57.405 8.785 57.695 8.815 ;
        RECT 57.025 8.600 57.695 8.785 ;
        RECT 73.350 8.785 73.525 10.860 ;
        RECT 73.730 8.785 74.020 8.815 ;
        RECT 73.350 8.600 74.020 8.785 ;
        RECT 89.675 8.785 89.850 10.860 ;
        RECT 90.055 8.785 90.345 8.815 ;
        RECT 89.675 8.600 90.345 8.785 ;
        RECT 24.755 8.585 25.045 8.600 ;
        RECT 41.080 8.585 41.370 8.600 ;
        RECT 57.405 8.585 57.695 8.600 ;
        RECT 73.730 8.585 74.020 8.600 ;
        RECT 90.055 8.585 90.345 8.600 ;
    END
    PORT
      LAYER li1 ;
        RECT 25.670 4.035 25.840 4.235 ;
        RECT 27.630 4.035 27.800 4.235 ;
        RECT 41.995 4.035 42.165 4.235 ;
        RECT 43.955 4.035 44.125 4.235 ;
        RECT 58.320 4.035 58.490 4.235 ;
        RECT 60.280 4.035 60.450 4.235 ;
        RECT 74.645 4.035 74.815 4.235 ;
        RECT 76.605 4.035 76.775 4.235 ;
        RECT 90.970 4.035 91.140 4.235 ;
        RECT 92.930 4.035 93.100 4.235 ;
        RECT 25.350 3.865 25.840 4.035 ;
        RECT 27.310 3.865 27.800 4.035 ;
        RECT 41.675 3.865 42.165 4.035 ;
        RECT 43.635 3.865 44.125 4.035 ;
        RECT 58.000 3.865 58.490 4.035 ;
        RECT 59.960 3.865 60.450 4.035 ;
        RECT 74.325 3.865 74.815 4.035 ;
        RECT 76.285 3.865 76.775 4.035 ;
        RECT 90.650 3.865 91.140 4.035 ;
        RECT 92.610 3.865 93.100 4.035 ;
        RECT 18.870 2.890 19.040 3.375 ;
        RECT 18.665 2.875 19.040 2.890 ;
        RECT 19.830 2.875 20.000 3.375 ;
        RECT 20.790 2.890 20.960 3.375 ;
        RECT 21.310 2.890 21.480 3.375 ;
        RECT 20.790 2.875 21.480 2.890 ;
        RECT 22.270 2.875 22.440 3.375 ;
        RECT 24.710 2.890 24.880 3.375 ;
        RECT 23.090 2.875 23.285 2.890 ;
        RECT 24.640 2.875 24.880 2.890 ;
        RECT 26.670 2.875 26.840 3.375 ;
        RECT 35.195 2.890 35.365 3.375 ;
        RECT 28.165 2.875 28.355 2.880 ;
        RECT 34.990 2.875 35.365 2.890 ;
        RECT 36.155 2.875 36.325 3.375 ;
        RECT 37.115 2.890 37.285 3.375 ;
        RECT 37.635 2.890 37.805 3.375 ;
        RECT 37.115 2.875 37.805 2.890 ;
        RECT 38.595 2.875 38.765 3.375 ;
        RECT 41.035 2.890 41.205 3.375 ;
        RECT 39.415 2.875 39.610 2.890 ;
        RECT 40.965 2.875 41.205 2.890 ;
        RECT 42.995 2.875 43.165 3.375 ;
        RECT 51.520 2.890 51.690 3.375 ;
        RECT 44.490 2.875 44.680 2.880 ;
        RECT 51.315 2.875 51.690 2.890 ;
        RECT 52.480 2.875 52.650 3.375 ;
        RECT 53.440 2.890 53.610 3.375 ;
        RECT 53.960 2.890 54.130 3.375 ;
        RECT 53.440 2.875 54.130 2.890 ;
        RECT 54.920 2.875 55.090 3.375 ;
        RECT 57.360 2.890 57.530 3.375 ;
        RECT 55.740 2.875 55.935 2.890 ;
        RECT 57.290 2.875 57.530 2.890 ;
        RECT 59.320 2.875 59.490 3.375 ;
        RECT 67.845 2.890 68.015 3.375 ;
        RECT 60.815 2.875 61.005 2.880 ;
        RECT 67.640 2.875 68.015 2.890 ;
        RECT 68.805 2.875 68.975 3.375 ;
        RECT 69.765 2.890 69.935 3.375 ;
        RECT 70.285 2.890 70.455 3.375 ;
        RECT 69.765 2.875 70.455 2.890 ;
        RECT 71.245 2.875 71.415 3.375 ;
        RECT 73.685 2.890 73.855 3.375 ;
        RECT 72.065 2.875 72.260 2.890 ;
        RECT 73.615 2.875 73.855 2.890 ;
        RECT 75.645 2.875 75.815 3.375 ;
        RECT 84.170 2.890 84.340 3.375 ;
        RECT 77.140 2.875 77.330 2.880 ;
        RECT 83.965 2.875 84.340 2.890 ;
        RECT 85.130 2.875 85.300 3.375 ;
        RECT 86.090 2.890 86.260 3.375 ;
        RECT 86.610 2.890 86.780 3.375 ;
        RECT 86.090 2.875 86.780 2.890 ;
        RECT 87.570 2.875 87.740 3.375 ;
        RECT 90.010 2.890 90.180 3.375 ;
        RECT 88.390 2.875 88.585 2.890 ;
        RECT 89.940 2.875 90.180 2.890 ;
        RECT 91.970 2.875 92.140 3.375 ;
        RECT 93.465 2.875 93.655 2.880 ;
        RECT 18.540 1.600 28.355 2.875 ;
        RECT 29.415 1.600 29.585 2.225 ;
        RECT 32.160 1.600 32.330 2.225 ;
        RECT 33.150 1.600 33.320 2.230 ;
        RECT 34.865 1.600 44.680 2.875 ;
        RECT 45.740 1.600 45.910 2.225 ;
        RECT 48.485 1.600 48.655 2.225 ;
        RECT 49.475 1.600 49.645 2.230 ;
        RECT 51.190 1.600 61.005 2.875 ;
        RECT 62.065 1.600 62.235 2.225 ;
        RECT 64.810 1.600 64.980 2.225 ;
        RECT 65.800 1.600 65.970 2.230 ;
        RECT 67.515 1.600 77.330 2.875 ;
        RECT 78.390 1.600 78.560 2.225 ;
        RECT 81.135 1.600 81.305 2.225 ;
        RECT 82.125 1.600 82.295 2.230 ;
        RECT 83.840 1.600 93.655 2.875 ;
        RECT 94.715 1.600 94.885 2.225 ;
        RECT 97.460 1.600 97.630 2.225 ;
        RECT 98.450 1.600 98.620 2.230 ;
        RECT 0.000 0.000 99.425 1.600 ;
      LAYER met1 ;
        RECT 25.940 4.350 27.540 4.365 ;
        RECT 42.265 4.350 43.865 4.365 ;
        RECT 58.590 4.350 60.190 4.365 ;
        RECT 74.915 4.350 76.515 4.365 ;
        RECT 91.240 4.350 92.840 4.365 ;
        RECT 25.940 4.285 27.710 4.350 ;
        RECT 42.265 4.285 44.035 4.350 ;
        RECT 58.590 4.285 60.360 4.350 ;
        RECT 74.915 4.285 76.685 4.350 ;
        RECT 91.240 4.285 93.010 4.350 ;
        RECT 25.940 4.265 27.750 4.285 ;
        RECT 42.265 4.265 44.075 4.285 ;
        RECT 58.590 4.265 60.400 4.285 ;
        RECT 74.915 4.265 76.725 4.285 ;
        RECT 91.240 4.265 93.050 4.285 ;
        RECT 25.610 4.240 27.860 4.265 ;
        RECT 41.935 4.240 44.185 4.265 ;
        RECT 58.260 4.240 60.510 4.265 ;
        RECT 74.585 4.240 76.835 4.265 ;
        RECT 90.910 4.240 93.160 4.265 ;
        RECT 25.610 4.225 28.355 4.240 ;
        RECT 25.610 4.085 26.080 4.225 ;
        RECT 27.400 4.085 28.355 4.225 ;
        RECT 25.610 4.035 25.900 4.085 ;
        RECT 27.430 4.055 28.355 4.085 ;
        RECT 27.430 4.035 27.860 4.055 ;
        RECT 27.430 4.025 27.750 4.035 ;
        RECT 28.170 2.905 28.355 4.055 ;
        RECT 41.935 4.225 44.680 4.240 ;
        RECT 41.935 4.085 42.405 4.225 ;
        RECT 43.725 4.085 44.680 4.225 ;
        RECT 41.935 4.035 42.225 4.085 ;
        RECT 43.755 4.055 44.680 4.085 ;
        RECT 43.755 4.035 44.185 4.055 ;
        RECT 43.755 4.025 44.075 4.035 ;
        RECT 44.495 2.905 44.680 4.055 ;
        RECT 58.260 4.225 61.005 4.240 ;
        RECT 58.260 4.085 58.730 4.225 ;
        RECT 60.050 4.085 61.005 4.225 ;
        RECT 58.260 4.035 58.550 4.085 ;
        RECT 60.080 4.055 61.005 4.085 ;
        RECT 60.080 4.035 60.510 4.055 ;
        RECT 60.080 4.025 60.400 4.035 ;
        RECT 60.820 2.905 61.005 4.055 ;
        RECT 74.585 4.225 77.330 4.240 ;
        RECT 74.585 4.085 75.055 4.225 ;
        RECT 76.375 4.085 77.330 4.225 ;
        RECT 74.585 4.035 74.875 4.085 ;
        RECT 76.405 4.055 77.330 4.085 ;
        RECT 76.405 4.035 76.835 4.055 ;
        RECT 76.405 4.025 76.725 4.035 ;
        RECT 77.145 2.905 77.330 4.055 ;
        RECT 90.910 4.225 93.655 4.240 ;
        RECT 90.910 4.085 91.380 4.225 ;
        RECT 92.700 4.085 93.655 4.225 ;
        RECT 90.910 4.035 91.200 4.085 ;
        RECT 92.730 4.055 93.655 4.085 ;
        RECT 92.730 4.035 93.160 4.055 ;
        RECT 92.730 4.025 93.050 4.035 ;
        RECT 93.470 2.905 93.655 4.055 ;
        RECT 18.540 1.600 28.355 2.905 ;
        RECT 34.865 1.600 44.680 2.905 ;
        RECT 51.190 1.600 61.005 2.905 ;
        RECT 67.515 1.600 77.330 2.905 ;
        RECT 83.840 1.600 93.655 2.905 ;
        RECT 0.000 0.000 99.425 1.600 ;
      LAYER met2 ;
        RECT 27.450 4.245 27.730 4.620 ;
        RECT 43.775 4.245 44.055 4.620 ;
        RECT 60.100 4.245 60.380 4.620 ;
        RECT 76.425 4.245 76.705 4.620 ;
        RECT 92.750 4.245 93.030 4.620 ;
        RECT 27.460 3.995 27.720 4.245 ;
        RECT 43.785 3.995 44.045 4.245 ;
        RECT 60.110 3.995 60.370 4.245 ;
        RECT 76.435 3.995 76.695 4.245 ;
        RECT 92.760 3.995 93.020 4.245 ;
      LAYER met3 ;
        RECT 27.430 4.595 27.760 4.995 ;
        RECT 43.755 4.595 44.085 4.995 ;
        RECT 60.080 4.595 60.410 4.995 ;
        RECT 76.405 4.595 76.735 4.995 ;
        RECT 92.730 4.595 93.060 4.995 ;
        RECT 27.425 4.265 27.760 4.595 ;
        RECT 43.750 4.265 44.085 4.595 ;
        RECT 60.075 4.265 60.410 4.595 ;
        RECT 76.400 4.265 76.735 4.595 ;
        RECT 92.725 4.265 93.060 4.595 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 15.000 8.740 17.810 8.745 ;
        RECT 23.580 8.740 26.390 8.745 ;
        RECT 29.195 8.740 32.985 8.745 ;
        RECT 39.905 8.740 42.715 8.745 ;
        RECT 45.520 8.740 49.310 8.745 ;
        RECT 56.230 8.740 59.040 8.745 ;
        RECT 61.845 8.740 65.635 8.745 ;
        RECT 72.555 8.740 75.365 8.745 ;
        RECT 78.170 8.740 81.960 8.745 ;
        RECT 88.880 8.740 91.690 8.745 ;
        RECT 94.495 8.740 98.285 8.745 ;
        RECT 15.000 4.100 99.425 8.740 ;
        RECT 17.790 4.095 99.425 4.100 ;
        RECT 28.175 4.020 34.125 4.095 ;
        RECT 44.500 4.020 50.450 4.095 ;
        RECT 60.825 4.020 66.775 4.095 ;
        RECT 77.150 4.020 83.100 4.095 ;
        RECT 93.475 4.020 99.425 4.095 ;
        RECT 28.180 3.720 34.125 4.020 ;
        RECT 44.505 3.720 50.450 4.020 ;
        RECT 60.830 3.720 66.775 4.020 ;
        RECT 77.155 3.720 83.100 4.020 ;
        RECT 93.480 3.720 99.425 4.020 ;
        RECT 29.195 3.715 32.985 3.720 ;
        RECT 45.520 3.715 49.310 3.720 ;
        RECT 61.845 3.715 65.635 3.720 ;
        RECT 78.170 3.715 81.960 3.720 ;
        RECT 94.495 3.715 98.285 3.720 ;
      LAYER li1 ;
        RECT 17.035 10.045 17.210 10.595 ;
        RECT 17.035 8.445 17.205 10.045 ;
        RECT 15.220 7.035 15.390 7.765 ;
        RECT 17.035 7.305 17.210 8.445 ;
        RECT 17.035 7.035 17.205 7.305 ;
        RECT 23.800 7.035 23.970 7.765 ;
        RECT 29.415 7.035 29.585 7.765 ;
        RECT 32.160 7.035 32.330 7.765 ;
        RECT 15.050 7.030 17.800 7.035 ;
        RECT 23.630 7.030 26.380 7.035 ;
        RECT 29.245 7.030 32.980 7.035 ;
        RECT 33.155 7.030 33.325 7.760 ;
        RECT 40.125 7.035 40.295 7.765 ;
        RECT 45.740 7.035 45.910 7.765 ;
        RECT 48.485 7.035 48.655 7.765 ;
        RECT 39.955 7.030 42.705 7.035 ;
        RECT 45.570 7.030 49.305 7.035 ;
        RECT 49.480 7.030 49.650 7.760 ;
        RECT 56.450 7.035 56.620 7.765 ;
        RECT 62.065 7.035 62.235 7.765 ;
        RECT 64.810 7.035 64.980 7.765 ;
        RECT 56.280 7.030 59.030 7.035 ;
        RECT 61.895 7.030 65.630 7.035 ;
        RECT 65.805 7.030 65.975 7.760 ;
        RECT 72.775 7.035 72.945 7.765 ;
        RECT 78.390 7.035 78.560 7.765 ;
        RECT 81.135 7.035 81.305 7.765 ;
        RECT 72.605 7.030 75.355 7.035 ;
        RECT 78.220 7.030 81.955 7.035 ;
        RECT 82.130 7.030 82.300 7.760 ;
        RECT 89.100 7.035 89.270 7.765 ;
        RECT 94.715 7.035 94.885 7.765 ;
        RECT 97.460 7.035 97.630 7.765 ;
        RECT 88.930 7.030 91.680 7.035 ;
        RECT 94.545 7.030 98.280 7.035 ;
        RECT 98.455 7.030 98.625 7.760 ;
        RECT 0.005 5.430 99.425 7.030 ;
        RECT 18.540 5.425 28.200 5.430 ;
        RECT 29.245 5.425 32.980 5.430 ;
        RECT 19.830 4.925 20.000 5.425 ;
        RECT 22.270 4.925 22.440 5.425 ;
        RECT 23.230 4.925 23.400 5.425 ;
        RECT 24.230 4.925 24.400 5.425 ;
        RECT 26.670 4.925 26.840 5.425 ;
        RECT 27.630 4.925 27.800 5.425 ;
        RECT 29.415 4.695 29.585 5.425 ;
        RECT 32.160 4.695 32.330 5.425 ;
        RECT 33.150 4.700 33.320 5.430 ;
        RECT 34.865 5.425 44.525 5.430 ;
        RECT 45.570 5.425 49.305 5.430 ;
        RECT 36.155 4.925 36.325 5.425 ;
        RECT 38.595 4.925 38.765 5.425 ;
        RECT 39.555 4.925 39.725 5.425 ;
        RECT 40.555 4.925 40.725 5.425 ;
        RECT 42.995 4.925 43.165 5.425 ;
        RECT 43.955 4.925 44.125 5.425 ;
        RECT 45.740 4.695 45.910 5.425 ;
        RECT 48.485 4.695 48.655 5.425 ;
        RECT 49.475 4.700 49.645 5.430 ;
        RECT 51.190 5.425 60.850 5.430 ;
        RECT 61.895 5.425 65.630 5.430 ;
        RECT 52.480 4.925 52.650 5.425 ;
        RECT 54.920 4.925 55.090 5.425 ;
        RECT 55.880 4.925 56.050 5.425 ;
        RECT 56.880 4.925 57.050 5.425 ;
        RECT 59.320 4.925 59.490 5.425 ;
        RECT 60.280 4.925 60.450 5.425 ;
        RECT 62.065 4.695 62.235 5.425 ;
        RECT 64.810 4.695 64.980 5.425 ;
        RECT 65.800 4.700 65.970 5.430 ;
        RECT 67.515 5.425 77.175 5.430 ;
        RECT 78.220 5.425 81.955 5.430 ;
        RECT 68.805 4.925 68.975 5.425 ;
        RECT 71.245 4.925 71.415 5.425 ;
        RECT 72.205 4.925 72.375 5.425 ;
        RECT 73.205 4.925 73.375 5.425 ;
        RECT 75.645 4.925 75.815 5.425 ;
        RECT 76.605 4.925 76.775 5.425 ;
        RECT 78.390 4.695 78.560 5.425 ;
        RECT 81.135 4.695 81.305 5.425 ;
        RECT 82.125 4.700 82.295 5.430 ;
        RECT 83.840 5.425 93.500 5.430 ;
        RECT 94.545 5.425 98.280 5.430 ;
        RECT 85.130 4.925 85.300 5.425 ;
        RECT 87.570 4.925 87.740 5.425 ;
        RECT 88.530 4.925 88.700 5.425 ;
        RECT 89.530 4.925 89.700 5.425 ;
        RECT 91.970 4.925 92.140 5.425 ;
        RECT 92.930 4.925 93.100 5.425 ;
        RECT 94.715 4.695 94.885 5.425 ;
        RECT 97.460 4.695 97.630 5.425 ;
        RECT 98.450 4.700 98.620 5.430 ;
      LAYER met1 ;
        RECT 16.975 9.145 17.265 9.175 ;
        RECT 16.805 8.975 17.265 9.145 ;
        RECT 16.975 8.945 17.265 8.975 ;
        RECT 15.050 7.030 17.800 7.035 ;
        RECT 23.630 7.030 26.380 7.035 ;
        RECT 29.245 7.030 32.980 7.035 ;
        RECT 39.955 7.030 42.705 7.035 ;
        RECT 45.570 7.030 49.305 7.035 ;
        RECT 56.280 7.030 59.030 7.035 ;
        RECT 61.895 7.030 65.630 7.035 ;
        RECT 72.605 7.030 75.355 7.035 ;
        RECT 78.220 7.030 81.955 7.035 ;
        RECT 88.930 7.030 91.680 7.035 ;
        RECT 94.545 7.030 98.280 7.035 ;
        RECT 0.005 5.430 99.425 7.030 ;
        RECT 18.540 5.395 28.200 5.430 ;
        RECT 29.245 5.425 32.980 5.430 ;
        RECT 34.865 5.395 44.525 5.430 ;
        RECT 45.570 5.425 49.305 5.430 ;
        RECT 51.190 5.395 60.850 5.430 ;
        RECT 61.895 5.425 65.630 5.430 ;
        RECT 67.515 5.395 77.175 5.430 ;
        RECT 78.220 5.425 81.955 5.430 ;
        RECT 83.840 5.395 93.500 5.430 ;
        RECT 94.545 5.425 98.280 5.430 ;
    END
  END vccd1
  OBS
      LAYER pwell ;
        RECT 18.700 2.735 18.870 2.875 ;
        RECT 18.680 2.715 18.870 2.735 ;
        RECT 21.140 2.715 21.310 2.875 ;
        RECT 23.580 2.715 23.750 2.875 ;
        RECT 26.020 2.735 26.190 2.875 ;
        RECT 35.025 2.735 35.195 2.875 ;
        RECT 26.020 2.715 26.210 2.735 ;
        RECT 18.680 2.705 18.850 2.715 ;
        RECT 26.040 2.705 26.210 2.715 ;
        RECT 35.005 2.715 35.195 2.735 ;
        RECT 37.465 2.715 37.635 2.875 ;
        RECT 39.905 2.715 40.075 2.875 ;
        RECT 42.345 2.735 42.515 2.875 ;
        RECT 51.350 2.735 51.520 2.875 ;
        RECT 42.345 2.715 42.535 2.735 ;
        RECT 35.005 2.705 35.175 2.715 ;
        RECT 42.365 2.705 42.535 2.715 ;
        RECT 51.330 2.715 51.520 2.735 ;
        RECT 53.790 2.715 53.960 2.875 ;
        RECT 56.230 2.715 56.400 2.875 ;
        RECT 58.670 2.735 58.840 2.875 ;
        RECT 67.675 2.735 67.845 2.875 ;
        RECT 58.670 2.715 58.860 2.735 ;
        RECT 51.330 2.705 51.500 2.715 ;
        RECT 58.690 2.705 58.860 2.715 ;
        RECT 67.655 2.715 67.845 2.735 ;
        RECT 70.115 2.715 70.285 2.875 ;
        RECT 72.555 2.715 72.725 2.875 ;
        RECT 74.995 2.735 75.165 2.875 ;
        RECT 84.000 2.735 84.170 2.875 ;
        RECT 74.995 2.715 75.185 2.735 ;
        RECT 67.655 2.705 67.825 2.715 ;
        RECT 75.015 2.705 75.185 2.715 ;
        RECT 83.980 2.715 84.170 2.735 ;
        RECT 86.440 2.715 86.610 2.875 ;
        RECT 88.880 2.715 89.050 2.875 ;
        RECT 91.320 2.735 91.490 2.875 ;
        RECT 91.320 2.715 91.510 2.735 ;
        RECT 83.980 2.705 84.150 2.715 ;
        RECT 91.340 2.705 91.510 2.715 ;
      LAYER li1 ;
        RECT 15.650 10.105 15.825 10.595 ;
        RECT 16.175 10.315 16.345 10.595 ;
        RECT 16.175 10.145 16.405 10.315 ;
        RECT 15.650 9.935 15.820 10.105 ;
        RECT 15.650 9.605 16.060 9.935 ;
        RECT 15.650 9.095 15.820 9.605 ;
        RECT 15.650 8.765 16.060 9.095 ;
        RECT 15.650 8.565 15.820 8.765 ;
        RECT 15.650 7.305 15.825 8.565 ;
        RECT 16.235 8.535 16.405 10.145 ;
        RECT 16.605 10.085 16.780 10.595 ;
        RECT 24.230 10.105 24.405 10.595 ;
        RECT 24.230 9.935 24.400 10.105 ;
        RECT 25.185 10.085 25.360 10.595 ;
        RECT 25.615 10.045 25.790 10.595 ;
        RECT 29.845 10.105 30.020 10.595 ;
        RECT 30.370 10.315 30.540 10.595 ;
        RECT 30.370 10.145 30.600 10.315 ;
        RECT 24.230 9.605 24.640 9.935 ;
        RECT 16.175 8.365 16.405 8.535 ;
        RECT 16.605 8.565 16.775 9.515 ;
        RECT 24.230 9.095 24.400 9.605 ;
        RECT 24.230 8.765 24.640 9.095 ;
        RECT 24.230 8.565 24.400 8.765 ;
        RECT 25.185 8.565 25.355 9.515 ;
        RECT 16.175 7.305 16.345 8.365 ;
        RECT 16.605 7.305 16.780 8.565 ;
        RECT 24.230 7.305 24.405 8.565 ;
        RECT 25.185 7.305 25.360 8.565 ;
        RECT 25.615 8.445 25.785 10.045 ;
        RECT 29.845 9.935 30.015 10.105 ;
        RECT 29.845 9.605 30.255 9.935 ;
        RECT 29.845 9.095 30.015 9.605 ;
        RECT 29.845 8.765 30.255 9.095 ;
        RECT 29.845 8.565 30.015 8.765 ;
        RECT 25.615 7.305 25.790 8.445 ;
        RECT 29.845 7.305 30.020 8.565 ;
        RECT 30.430 8.535 30.600 10.145 ;
        RECT 30.800 10.085 30.975 10.595 ;
        RECT 31.230 10.045 31.405 10.595 ;
        RECT 32.595 10.085 32.765 10.595 ;
        RECT 33.590 10.080 33.760 10.590 ;
        RECT 40.555 10.105 40.730 10.595 ;
        RECT 30.370 8.365 30.600 8.535 ;
        RECT 30.800 8.565 30.970 9.515 ;
        RECT 30.370 7.305 30.540 8.365 ;
        RECT 30.800 7.305 30.975 8.565 ;
        RECT 31.230 8.445 31.400 10.045 ;
        RECT 40.555 9.935 40.725 10.105 ;
        RECT 41.510 10.085 41.685 10.595 ;
        RECT 41.940 10.045 42.115 10.595 ;
        RECT 46.170 10.105 46.345 10.595 ;
        RECT 46.695 10.315 46.865 10.595 ;
        RECT 46.695 10.145 46.925 10.315 ;
        RECT 40.555 9.605 40.965 9.935 ;
        RECT 31.770 9.425 32.000 9.575 ;
        RECT 31.770 9.255 32.690 9.425 ;
        RECT 32.220 8.565 32.390 9.255 ;
        RECT 33.215 9.250 33.685 9.420 ;
        RECT 32.590 8.775 32.760 8.885 ;
        RECT 33.215 8.775 33.385 9.250 ;
        RECT 40.555 9.095 40.725 9.605 ;
        RECT 32.590 8.605 33.385 8.775 ;
        RECT 31.230 7.305 31.405 8.445 ;
        RECT 32.590 7.305 32.765 8.605 ;
        RECT 33.215 8.560 33.385 8.605 ;
        RECT 33.585 8.445 33.755 8.880 ;
        RECT 40.555 8.765 40.965 9.095 ;
        RECT 40.555 8.565 40.725 8.765 ;
        RECT 41.510 8.565 41.680 9.515 ;
        RECT 33.585 7.300 33.760 8.445 ;
        RECT 40.555 7.305 40.730 8.565 ;
        RECT 41.510 7.305 41.685 8.565 ;
        RECT 41.940 8.445 42.110 10.045 ;
        RECT 46.170 9.935 46.340 10.105 ;
        RECT 46.170 9.605 46.580 9.935 ;
        RECT 46.170 9.095 46.340 9.605 ;
        RECT 46.170 8.765 46.580 9.095 ;
        RECT 46.170 8.565 46.340 8.765 ;
        RECT 41.940 7.305 42.115 8.445 ;
        RECT 46.170 7.305 46.345 8.565 ;
        RECT 46.755 8.535 46.925 10.145 ;
        RECT 47.125 10.085 47.300 10.595 ;
        RECT 47.555 10.045 47.730 10.595 ;
        RECT 48.920 10.085 49.090 10.595 ;
        RECT 49.915 10.080 50.085 10.590 ;
        RECT 56.880 10.105 57.055 10.595 ;
        RECT 46.695 8.365 46.925 8.535 ;
        RECT 47.125 8.565 47.295 9.515 ;
        RECT 46.695 7.305 46.865 8.365 ;
        RECT 47.125 7.305 47.300 8.565 ;
        RECT 47.555 8.445 47.725 10.045 ;
        RECT 56.880 9.935 57.050 10.105 ;
        RECT 57.835 10.085 58.010 10.595 ;
        RECT 58.265 10.045 58.440 10.595 ;
        RECT 62.495 10.105 62.670 10.595 ;
        RECT 63.020 10.315 63.190 10.595 ;
        RECT 63.020 10.145 63.250 10.315 ;
        RECT 56.880 9.605 57.290 9.935 ;
        RECT 48.095 9.425 48.325 9.575 ;
        RECT 48.095 9.255 49.015 9.425 ;
        RECT 48.545 8.565 48.715 9.255 ;
        RECT 49.540 9.250 50.010 9.420 ;
        RECT 48.915 8.775 49.085 8.885 ;
        RECT 49.540 8.775 49.710 9.250 ;
        RECT 56.880 9.095 57.050 9.605 ;
        RECT 48.915 8.605 49.710 8.775 ;
        RECT 47.555 7.305 47.730 8.445 ;
        RECT 48.915 7.305 49.090 8.605 ;
        RECT 49.540 8.560 49.710 8.605 ;
        RECT 49.910 8.445 50.080 8.880 ;
        RECT 56.880 8.765 57.290 9.095 ;
        RECT 56.880 8.565 57.050 8.765 ;
        RECT 57.835 8.565 58.005 9.515 ;
        RECT 49.910 7.300 50.085 8.445 ;
        RECT 56.880 7.305 57.055 8.565 ;
        RECT 57.835 7.305 58.010 8.565 ;
        RECT 58.265 8.445 58.435 10.045 ;
        RECT 62.495 9.935 62.665 10.105 ;
        RECT 62.495 9.605 62.905 9.935 ;
        RECT 62.495 9.095 62.665 9.605 ;
        RECT 62.495 8.765 62.905 9.095 ;
        RECT 62.495 8.565 62.665 8.765 ;
        RECT 58.265 7.305 58.440 8.445 ;
        RECT 62.495 7.305 62.670 8.565 ;
        RECT 63.080 8.535 63.250 10.145 ;
        RECT 63.450 10.085 63.625 10.595 ;
        RECT 63.880 10.045 64.055 10.595 ;
        RECT 65.245 10.085 65.415 10.595 ;
        RECT 66.240 10.080 66.410 10.590 ;
        RECT 73.205 10.105 73.380 10.595 ;
        RECT 63.020 8.365 63.250 8.535 ;
        RECT 63.450 8.565 63.620 9.515 ;
        RECT 63.020 7.305 63.190 8.365 ;
        RECT 63.450 7.305 63.625 8.565 ;
        RECT 63.880 8.445 64.050 10.045 ;
        RECT 73.205 9.935 73.375 10.105 ;
        RECT 74.160 10.085 74.335 10.595 ;
        RECT 74.590 10.045 74.765 10.595 ;
        RECT 78.820 10.105 78.995 10.595 ;
        RECT 79.345 10.315 79.515 10.595 ;
        RECT 79.345 10.145 79.575 10.315 ;
        RECT 73.205 9.605 73.615 9.935 ;
        RECT 64.420 9.425 64.650 9.575 ;
        RECT 64.420 9.255 65.340 9.425 ;
        RECT 64.870 8.565 65.040 9.255 ;
        RECT 65.865 9.250 66.335 9.420 ;
        RECT 65.240 8.775 65.410 8.885 ;
        RECT 65.865 8.775 66.035 9.250 ;
        RECT 73.205 9.095 73.375 9.605 ;
        RECT 65.240 8.605 66.035 8.775 ;
        RECT 63.880 7.305 64.055 8.445 ;
        RECT 65.240 7.305 65.415 8.605 ;
        RECT 65.865 8.560 66.035 8.605 ;
        RECT 66.235 8.445 66.405 8.880 ;
        RECT 73.205 8.765 73.615 9.095 ;
        RECT 73.205 8.565 73.375 8.765 ;
        RECT 74.160 8.565 74.330 9.515 ;
        RECT 66.235 7.300 66.410 8.445 ;
        RECT 73.205 7.305 73.380 8.565 ;
        RECT 74.160 7.305 74.335 8.565 ;
        RECT 74.590 8.445 74.760 10.045 ;
        RECT 78.820 9.935 78.990 10.105 ;
        RECT 78.820 9.605 79.230 9.935 ;
        RECT 78.820 9.095 78.990 9.605 ;
        RECT 78.820 8.765 79.230 9.095 ;
        RECT 78.820 8.565 78.990 8.765 ;
        RECT 74.590 7.305 74.765 8.445 ;
        RECT 78.820 7.305 78.995 8.565 ;
        RECT 79.405 8.535 79.575 10.145 ;
        RECT 79.775 10.085 79.950 10.595 ;
        RECT 80.205 10.045 80.380 10.595 ;
        RECT 81.570 10.085 81.740 10.595 ;
        RECT 82.565 10.080 82.735 10.590 ;
        RECT 89.530 10.105 89.705 10.595 ;
        RECT 79.345 8.365 79.575 8.535 ;
        RECT 79.775 8.565 79.945 9.515 ;
        RECT 79.345 7.305 79.515 8.365 ;
        RECT 79.775 7.305 79.950 8.565 ;
        RECT 80.205 8.445 80.375 10.045 ;
        RECT 89.530 9.935 89.700 10.105 ;
        RECT 90.485 10.085 90.660 10.595 ;
        RECT 90.915 10.045 91.090 10.595 ;
        RECT 95.145 10.105 95.320 10.595 ;
        RECT 95.670 10.315 95.840 10.595 ;
        RECT 95.670 10.145 95.900 10.315 ;
        RECT 89.530 9.605 89.940 9.935 ;
        RECT 80.745 9.425 80.975 9.575 ;
        RECT 80.745 9.255 81.665 9.425 ;
        RECT 81.195 8.565 81.365 9.255 ;
        RECT 82.190 9.250 82.660 9.420 ;
        RECT 81.565 8.775 81.735 8.885 ;
        RECT 82.190 8.775 82.360 9.250 ;
        RECT 89.530 9.095 89.700 9.605 ;
        RECT 81.565 8.605 82.360 8.775 ;
        RECT 80.205 7.305 80.380 8.445 ;
        RECT 81.565 7.305 81.740 8.605 ;
        RECT 82.190 8.560 82.360 8.605 ;
        RECT 82.560 8.445 82.730 8.880 ;
        RECT 89.530 8.765 89.940 9.095 ;
        RECT 89.530 8.565 89.700 8.765 ;
        RECT 90.485 8.565 90.655 9.515 ;
        RECT 82.560 7.300 82.735 8.445 ;
        RECT 89.530 7.305 89.705 8.565 ;
        RECT 90.485 7.305 90.660 8.565 ;
        RECT 90.915 8.445 91.085 10.045 ;
        RECT 95.145 9.935 95.315 10.105 ;
        RECT 95.145 9.605 95.555 9.935 ;
        RECT 95.145 9.095 95.315 9.605 ;
        RECT 95.145 8.765 95.555 9.095 ;
        RECT 95.145 8.565 95.315 8.765 ;
        RECT 90.915 7.305 91.090 8.445 ;
        RECT 95.145 7.305 95.320 8.565 ;
        RECT 95.730 8.535 95.900 10.145 ;
        RECT 96.100 10.085 96.275 10.595 ;
        RECT 96.530 10.045 96.705 10.595 ;
        RECT 97.895 10.085 98.065 10.595 ;
        RECT 98.890 10.080 99.060 10.590 ;
        RECT 95.670 8.365 95.900 8.535 ;
        RECT 96.100 8.565 96.270 9.515 ;
        RECT 95.670 7.305 95.840 8.365 ;
        RECT 96.100 7.305 96.275 8.565 ;
        RECT 96.530 8.445 96.700 10.045 ;
        RECT 97.070 9.425 97.300 9.575 ;
        RECT 97.070 9.255 97.990 9.425 ;
        RECT 97.520 8.565 97.690 9.255 ;
        RECT 98.515 9.250 98.985 9.420 ;
        RECT 97.890 8.775 98.060 8.885 ;
        RECT 98.515 8.775 98.685 9.250 ;
        RECT 97.890 8.605 98.685 8.775 ;
        RECT 96.530 7.305 96.705 8.445 ;
        RECT 97.890 7.305 98.065 8.605 ;
        RECT 98.515 8.560 98.685 8.605 ;
        RECT 98.885 8.445 99.055 8.880 ;
        RECT 98.885 7.300 99.060 8.445 ;
        RECT 19.230 4.905 19.520 5.075 ;
        RECT 18.870 4.345 19.040 4.765 ;
        RECT 19.230 4.035 19.400 4.905 ;
        RECT 20.550 4.625 20.960 4.795 ;
        RECT 19.030 3.865 19.400 4.035 ;
        RECT 19.590 4.345 20.240 4.515 ;
        RECT 20.790 4.435 20.960 4.625 ;
        RECT 21.310 4.345 21.480 4.765 ;
        RECT 21.670 4.625 21.960 4.795 ;
        RECT 19.590 3.785 19.760 4.345 ;
        RECT 20.070 3.785 20.240 4.115 ;
        RECT 21.670 4.035 21.840 4.625 ;
        RECT 22.750 4.435 22.920 4.795 ;
        RECT 25.190 4.775 25.360 5.105 ;
        RECT 26.190 4.775 26.360 5.105 ;
        RECT 23.670 4.605 24.960 4.685 ;
        RECT 25.590 4.605 25.920 4.685 ;
        RECT 23.670 4.515 25.920 4.605 ;
        RECT 27.070 4.515 27.400 4.685 ;
        RECT 24.710 4.435 25.840 4.515 ;
        RECT 26.310 4.345 27.320 4.515 ;
        RECT 20.470 3.865 20.960 4.035 ;
        RECT 21.470 3.865 21.840 4.035 ;
        RECT 20.790 3.785 20.960 3.865 ;
        RECT 22.030 3.785 22.200 4.115 ;
        RECT 22.510 3.785 22.680 4.235 ;
        RECT 22.910 3.865 24.240 4.035 ;
        RECT 23.990 3.785 24.160 3.865 ;
        RECT 24.470 3.785 24.640 4.115 ;
        RECT 24.950 3.785 25.120 4.235 ;
        RECT 26.310 4.115 26.480 4.345 ;
        RECT 26.310 3.865 26.600 4.115 ;
        RECT 26.430 3.785 26.600 3.865 ;
        RECT 26.910 3.785 27.080 4.115 ;
        RECT 29.845 3.895 30.020 5.155 ;
        RECT 30.370 4.095 30.540 5.155 ;
        RECT 30.370 3.925 30.600 4.095 ;
        RECT 29.845 3.695 30.015 3.895 ;
        RECT 22.990 3.635 23.160 3.675 ;
        RECT 22.990 3.465 23.480 3.635 ;
        RECT 25.430 3.505 25.840 3.675 ;
        RECT 19.350 3.045 19.520 3.395 ;
        RECT 20.310 3.045 20.480 3.395 ;
        RECT 21.790 3.045 21.960 3.395 ;
        RECT 23.750 3.045 23.920 3.395 ;
        RECT 25.670 3.045 25.840 3.505 ;
        RECT 26.190 3.045 26.360 3.395 ;
        RECT 27.150 3.295 27.320 3.395 ;
        RECT 29.845 3.365 30.255 3.695 ;
        RECT 27.150 3.125 27.880 3.295 ;
        RECT 29.845 2.855 30.015 3.365 ;
        RECT 29.845 2.525 30.255 2.855 ;
        RECT 29.845 2.355 30.015 2.525 ;
        RECT 29.845 1.865 30.020 2.355 ;
        RECT 30.430 2.315 30.600 3.925 ;
        RECT 30.800 3.895 30.975 5.155 ;
        RECT 31.230 4.015 31.405 5.155 ;
        RECT 30.800 2.945 30.970 3.895 ;
        RECT 31.230 2.415 31.400 4.015 ;
        RECT 32.590 4.010 32.765 5.155 ;
        RECT 35.555 4.905 35.845 5.075 ;
        RECT 35.195 4.345 35.365 4.765 ;
        RECT 35.555 4.035 35.725 4.905 ;
        RECT 36.875 4.625 37.285 4.795 ;
        RECT 32.220 3.205 32.390 3.895 ;
        RECT 32.590 3.795 32.760 4.010 ;
        RECT 33.210 3.795 33.380 3.900 ;
        RECT 35.355 3.865 35.725 4.035 ;
        RECT 35.915 4.345 36.565 4.515 ;
        RECT 37.115 4.435 37.285 4.625 ;
        RECT 37.635 4.345 37.805 4.765 ;
        RECT 37.995 4.625 38.285 4.795 ;
        RECT 32.590 3.625 33.380 3.795 ;
        RECT 35.915 3.785 36.085 4.345 ;
        RECT 36.395 3.785 36.565 4.115 ;
        RECT 37.995 4.035 38.165 4.625 ;
        RECT 39.075 4.435 39.245 4.795 ;
        RECT 41.515 4.775 41.685 5.105 ;
        RECT 42.515 4.775 42.685 5.105 ;
        RECT 39.995 4.605 41.285 4.685 ;
        RECT 41.915 4.605 42.245 4.685 ;
        RECT 39.995 4.515 42.245 4.605 ;
        RECT 43.395 4.515 43.725 4.685 ;
        RECT 41.035 4.435 42.165 4.515 ;
        RECT 42.635 4.345 43.645 4.515 ;
        RECT 36.795 3.865 37.285 4.035 ;
        RECT 37.795 3.865 38.165 4.035 ;
        RECT 37.115 3.785 37.285 3.865 ;
        RECT 38.355 3.785 38.525 4.115 ;
        RECT 38.835 3.785 39.005 4.235 ;
        RECT 39.235 3.865 40.565 4.035 ;
        RECT 40.315 3.785 40.485 3.865 ;
        RECT 40.795 3.785 40.965 4.115 ;
        RECT 41.275 3.785 41.445 4.235 ;
        RECT 42.635 4.115 42.805 4.345 ;
        RECT 42.635 3.865 42.925 4.115 ;
        RECT 42.755 3.785 42.925 3.865 ;
        RECT 43.235 3.785 43.405 4.115 ;
        RECT 46.170 3.895 46.345 5.155 ;
        RECT 46.695 4.095 46.865 5.155 ;
        RECT 46.695 3.925 46.925 4.095 ;
        RECT 46.170 3.695 46.340 3.895 ;
        RECT 32.590 3.575 32.760 3.625 ;
        RECT 33.210 3.210 33.380 3.625 ;
        RECT 39.315 3.635 39.485 3.675 ;
        RECT 39.315 3.465 39.805 3.635 ;
        RECT 41.755 3.505 42.165 3.675 ;
        RECT 31.770 3.035 32.690 3.205 ;
        RECT 33.210 3.040 33.680 3.210 ;
        RECT 35.675 3.045 35.845 3.395 ;
        RECT 36.635 3.045 36.805 3.395 ;
        RECT 38.115 3.045 38.285 3.395 ;
        RECT 40.075 3.045 40.245 3.395 ;
        RECT 41.995 3.045 42.165 3.505 ;
        RECT 42.515 3.045 42.685 3.395 ;
        RECT 43.475 3.295 43.645 3.395 ;
        RECT 46.170 3.365 46.580 3.695 ;
        RECT 43.475 3.125 44.205 3.295 ;
        RECT 31.770 2.885 32.000 3.035 ;
        RECT 46.170 2.855 46.340 3.365 ;
        RECT 46.170 2.525 46.580 2.855 ;
        RECT 30.370 2.145 30.600 2.315 ;
        RECT 30.370 1.865 30.540 2.145 ;
        RECT 30.800 1.865 30.975 2.375 ;
        RECT 31.230 1.865 31.405 2.415 ;
        RECT 32.595 1.865 32.765 2.375 ;
        RECT 46.170 2.355 46.340 2.525 ;
        RECT 46.170 1.865 46.345 2.355 ;
        RECT 46.755 2.315 46.925 3.925 ;
        RECT 47.125 3.895 47.300 5.155 ;
        RECT 47.555 4.015 47.730 5.155 ;
        RECT 47.125 2.945 47.295 3.895 ;
        RECT 47.555 2.415 47.725 4.015 ;
        RECT 48.915 4.010 49.090 5.155 ;
        RECT 51.880 4.905 52.170 5.075 ;
        RECT 51.520 4.345 51.690 4.765 ;
        RECT 51.880 4.035 52.050 4.905 ;
        RECT 53.200 4.625 53.610 4.795 ;
        RECT 48.545 3.205 48.715 3.895 ;
        RECT 48.915 3.795 49.085 4.010 ;
        RECT 49.535 3.795 49.705 3.900 ;
        RECT 51.680 3.865 52.050 4.035 ;
        RECT 52.240 4.345 52.890 4.515 ;
        RECT 53.440 4.435 53.610 4.625 ;
        RECT 53.960 4.345 54.130 4.765 ;
        RECT 54.320 4.625 54.610 4.795 ;
        RECT 48.915 3.625 49.705 3.795 ;
        RECT 52.240 3.785 52.410 4.345 ;
        RECT 52.720 3.785 52.890 4.115 ;
        RECT 54.320 4.035 54.490 4.625 ;
        RECT 55.400 4.435 55.570 4.795 ;
        RECT 57.840 4.775 58.010 5.105 ;
        RECT 58.840 4.775 59.010 5.105 ;
        RECT 56.320 4.605 57.610 4.685 ;
        RECT 58.240 4.605 58.570 4.685 ;
        RECT 56.320 4.515 58.570 4.605 ;
        RECT 59.720 4.515 60.050 4.685 ;
        RECT 57.360 4.435 58.490 4.515 ;
        RECT 58.960 4.345 59.970 4.515 ;
        RECT 53.120 3.865 53.610 4.035 ;
        RECT 54.120 3.865 54.490 4.035 ;
        RECT 53.440 3.785 53.610 3.865 ;
        RECT 54.680 3.785 54.850 4.115 ;
        RECT 55.160 3.785 55.330 4.235 ;
        RECT 55.560 3.865 56.890 4.035 ;
        RECT 56.640 3.785 56.810 3.865 ;
        RECT 57.120 3.785 57.290 4.115 ;
        RECT 57.600 3.785 57.770 4.235 ;
        RECT 58.960 4.115 59.130 4.345 ;
        RECT 58.960 3.865 59.250 4.115 ;
        RECT 59.080 3.785 59.250 3.865 ;
        RECT 59.560 3.785 59.730 4.115 ;
        RECT 62.495 3.895 62.670 5.155 ;
        RECT 63.020 4.095 63.190 5.155 ;
        RECT 63.020 3.925 63.250 4.095 ;
        RECT 62.495 3.695 62.665 3.895 ;
        RECT 48.915 3.575 49.085 3.625 ;
        RECT 49.535 3.210 49.705 3.625 ;
        RECT 55.640 3.635 55.810 3.675 ;
        RECT 55.640 3.465 56.130 3.635 ;
        RECT 58.080 3.505 58.490 3.675 ;
        RECT 48.095 3.035 49.015 3.205 ;
        RECT 49.535 3.040 50.005 3.210 ;
        RECT 52.000 3.045 52.170 3.395 ;
        RECT 52.960 3.045 53.130 3.395 ;
        RECT 54.440 3.045 54.610 3.395 ;
        RECT 56.400 3.045 56.570 3.395 ;
        RECT 58.320 3.045 58.490 3.505 ;
        RECT 58.840 3.045 59.010 3.395 ;
        RECT 59.800 3.295 59.970 3.395 ;
        RECT 62.495 3.365 62.905 3.695 ;
        RECT 59.800 3.125 60.530 3.295 ;
        RECT 48.095 2.885 48.325 3.035 ;
        RECT 62.495 2.855 62.665 3.365 ;
        RECT 62.495 2.525 62.905 2.855 ;
        RECT 46.695 2.145 46.925 2.315 ;
        RECT 46.695 1.865 46.865 2.145 ;
        RECT 47.125 1.865 47.300 2.375 ;
        RECT 47.555 1.865 47.730 2.415 ;
        RECT 48.920 1.865 49.090 2.375 ;
        RECT 62.495 2.355 62.665 2.525 ;
        RECT 62.495 1.865 62.670 2.355 ;
        RECT 63.080 2.315 63.250 3.925 ;
        RECT 63.450 3.895 63.625 5.155 ;
        RECT 63.880 4.015 64.055 5.155 ;
        RECT 63.450 2.945 63.620 3.895 ;
        RECT 63.880 2.415 64.050 4.015 ;
        RECT 65.240 4.010 65.415 5.155 ;
        RECT 68.205 4.905 68.495 5.075 ;
        RECT 67.845 4.345 68.015 4.765 ;
        RECT 68.205 4.035 68.375 4.905 ;
        RECT 69.525 4.625 69.935 4.795 ;
        RECT 64.870 3.205 65.040 3.895 ;
        RECT 65.240 3.795 65.410 4.010 ;
        RECT 65.860 3.795 66.030 3.900 ;
        RECT 68.005 3.865 68.375 4.035 ;
        RECT 68.565 4.345 69.215 4.515 ;
        RECT 69.765 4.435 69.935 4.625 ;
        RECT 70.285 4.345 70.455 4.765 ;
        RECT 70.645 4.625 70.935 4.795 ;
        RECT 65.240 3.625 66.030 3.795 ;
        RECT 68.565 3.785 68.735 4.345 ;
        RECT 69.045 3.785 69.215 4.115 ;
        RECT 70.645 4.035 70.815 4.625 ;
        RECT 71.725 4.435 71.895 4.795 ;
        RECT 74.165 4.775 74.335 5.105 ;
        RECT 75.165 4.775 75.335 5.105 ;
        RECT 72.645 4.605 73.935 4.685 ;
        RECT 74.565 4.605 74.895 4.685 ;
        RECT 72.645 4.515 74.895 4.605 ;
        RECT 76.045 4.515 76.375 4.685 ;
        RECT 73.685 4.435 74.815 4.515 ;
        RECT 75.285 4.345 76.295 4.515 ;
        RECT 69.445 3.865 69.935 4.035 ;
        RECT 70.445 3.865 70.815 4.035 ;
        RECT 69.765 3.785 69.935 3.865 ;
        RECT 71.005 3.785 71.175 4.115 ;
        RECT 71.485 3.785 71.655 4.235 ;
        RECT 71.885 3.865 73.215 4.035 ;
        RECT 72.965 3.785 73.135 3.865 ;
        RECT 73.445 3.785 73.615 4.115 ;
        RECT 73.925 3.785 74.095 4.235 ;
        RECT 75.285 4.115 75.455 4.345 ;
        RECT 75.285 3.865 75.575 4.115 ;
        RECT 75.405 3.785 75.575 3.865 ;
        RECT 75.885 3.785 76.055 4.115 ;
        RECT 78.820 3.895 78.995 5.155 ;
        RECT 79.345 4.095 79.515 5.155 ;
        RECT 79.345 3.925 79.575 4.095 ;
        RECT 78.820 3.695 78.990 3.895 ;
        RECT 65.240 3.575 65.410 3.625 ;
        RECT 65.860 3.210 66.030 3.625 ;
        RECT 71.965 3.635 72.135 3.675 ;
        RECT 71.965 3.465 72.455 3.635 ;
        RECT 74.405 3.505 74.815 3.675 ;
        RECT 64.420 3.035 65.340 3.205 ;
        RECT 65.860 3.040 66.330 3.210 ;
        RECT 68.325 3.045 68.495 3.395 ;
        RECT 69.285 3.045 69.455 3.395 ;
        RECT 70.765 3.045 70.935 3.395 ;
        RECT 72.725 3.045 72.895 3.395 ;
        RECT 74.645 3.045 74.815 3.505 ;
        RECT 75.165 3.045 75.335 3.395 ;
        RECT 76.125 3.295 76.295 3.395 ;
        RECT 78.820 3.365 79.230 3.695 ;
        RECT 76.125 3.125 76.855 3.295 ;
        RECT 64.420 2.885 64.650 3.035 ;
        RECT 78.820 2.855 78.990 3.365 ;
        RECT 78.820 2.525 79.230 2.855 ;
        RECT 63.020 2.145 63.250 2.315 ;
        RECT 63.020 1.865 63.190 2.145 ;
        RECT 63.450 1.865 63.625 2.375 ;
        RECT 63.880 1.865 64.055 2.415 ;
        RECT 65.245 1.865 65.415 2.375 ;
        RECT 78.820 2.355 78.990 2.525 ;
        RECT 78.820 1.865 78.995 2.355 ;
        RECT 79.405 2.315 79.575 3.925 ;
        RECT 79.775 3.895 79.950 5.155 ;
        RECT 80.205 4.015 80.380 5.155 ;
        RECT 79.775 2.945 79.945 3.895 ;
        RECT 80.205 2.415 80.375 4.015 ;
        RECT 81.565 4.010 81.740 5.155 ;
        RECT 84.530 4.905 84.820 5.075 ;
        RECT 84.170 4.345 84.340 4.765 ;
        RECT 84.530 4.035 84.700 4.905 ;
        RECT 85.850 4.625 86.260 4.795 ;
        RECT 81.195 3.205 81.365 3.895 ;
        RECT 81.565 3.795 81.735 4.010 ;
        RECT 82.185 3.795 82.355 3.900 ;
        RECT 84.330 3.865 84.700 4.035 ;
        RECT 84.890 4.345 85.540 4.515 ;
        RECT 86.090 4.435 86.260 4.625 ;
        RECT 86.610 4.345 86.780 4.765 ;
        RECT 86.970 4.625 87.260 4.795 ;
        RECT 81.565 3.625 82.355 3.795 ;
        RECT 84.890 3.785 85.060 4.345 ;
        RECT 85.370 3.785 85.540 4.115 ;
        RECT 86.970 4.035 87.140 4.625 ;
        RECT 88.050 4.435 88.220 4.795 ;
        RECT 90.490 4.775 90.660 5.105 ;
        RECT 91.490 4.775 91.660 5.105 ;
        RECT 88.970 4.605 90.260 4.685 ;
        RECT 90.890 4.605 91.220 4.685 ;
        RECT 88.970 4.515 91.220 4.605 ;
        RECT 92.370 4.515 92.700 4.685 ;
        RECT 90.010 4.435 91.140 4.515 ;
        RECT 91.610 4.345 92.620 4.515 ;
        RECT 85.770 3.865 86.260 4.035 ;
        RECT 86.770 3.865 87.140 4.035 ;
        RECT 86.090 3.785 86.260 3.865 ;
        RECT 87.330 3.785 87.500 4.115 ;
        RECT 87.810 3.785 87.980 4.235 ;
        RECT 88.210 3.865 89.540 4.035 ;
        RECT 89.290 3.785 89.460 3.865 ;
        RECT 89.770 3.785 89.940 4.115 ;
        RECT 90.250 3.785 90.420 4.235 ;
        RECT 91.610 4.115 91.780 4.345 ;
        RECT 91.610 3.865 91.900 4.115 ;
        RECT 91.730 3.785 91.900 3.865 ;
        RECT 92.210 3.785 92.380 4.115 ;
        RECT 95.145 3.895 95.320 5.155 ;
        RECT 95.670 4.095 95.840 5.155 ;
        RECT 95.670 3.925 95.900 4.095 ;
        RECT 95.145 3.695 95.315 3.895 ;
        RECT 81.565 3.575 81.735 3.625 ;
        RECT 82.185 3.210 82.355 3.625 ;
        RECT 88.290 3.635 88.460 3.675 ;
        RECT 88.290 3.465 88.780 3.635 ;
        RECT 90.730 3.505 91.140 3.675 ;
        RECT 80.745 3.035 81.665 3.205 ;
        RECT 82.185 3.040 82.655 3.210 ;
        RECT 84.650 3.045 84.820 3.395 ;
        RECT 85.610 3.045 85.780 3.395 ;
        RECT 87.090 3.045 87.260 3.395 ;
        RECT 89.050 3.045 89.220 3.395 ;
        RECT 90.970 3.045 91.140 3.505 ;
        RECT 91.490 3.045 91.660 3.395 ;
        RECT 92.450 3.295 92.620 3.395 ;
        RECT 95.145 3.365 95.555 3.695 ;
        RECT 92.450 3.125 93.180 3.295 ;
        RECT 80.745 2.885 80.975 3.035 ;
        RECT 95.145 2.855 95.315 3.365 ;
        RECT 95.145 2.525 95.555 2.855 ;
        RECT 79.345 2.145 79.575 2.315 ;
        RECT 79.345 1.865 79.515 2.145 ;
        RECT 79.775 1.865 79.950 2.375 ;
        RECT 80.205 1.865 80.380 2.415 ;
        RECT 81.570 1.865 81.740 2.375 ;
        RECT 95.145 2.355 95.315 2.525 ;
        RECT 95.145 1.865 95.320 2.355 ;
        RECT 95.730 2.315 95.900 3.925 ;
        RECT 96.100 3.895 96.275 5.155 ;
        RECT 96.530 4.015 96.705 5.155 ;
        RECT 96.100 2.945 96.270 3.895 ;
        RECT 96.530 2.415 96.700 4.015 ;
        RECT 97.890 4.010 98.065 5.155 ;
        RECT 97.520 3.205 97.690 3.895 ;
        RECT 97.890 3.795 98.060 4.010 ;
        RECT 98.510 3.795 98.680 3.900 ;
        RECT 97.890 3.625 98.680 3.795 ;
        RECT 97.890 3.575 98.060 3.625 ;
        RECT 98.510 3.210 98.680 3.625 ;
        RECT 97.070 3.035 97.990 3.205 ;
        RECT 98.510 3.040 98.980 3.210 ;
        RECT 97.070 2.885 97.300 3.035 ;
        RECT 95.670 2.145 95.900 2.315 ;
        RECT 95.670 1.865 95.840 2.145 ;
        RECT 96.100 1.865 96.275 2.375 ;
        RECT 96.530 1.865 96.705 2.415 ;
        RECT 97.895 1.865 98.065 2.375 ;
      LAYER met1 ;
        RECT 16.545 10.055 16.835 10.285 ;
        RECT 25.125 10.055 25.415 10.285 ;
        RECT 30.740 10.055 31.030 10.285 ;
        RECT 16.605 9.605 16.775 10.055 ;
        RECT 25.185 9.710 25.355 10.055 ;
        RECT 16.515 9.315 16.865 9.605 ;
        RECT 25.105 9.360 25.475 9.710 ;
        RECT 30.800 9.575 30.970 10.055 ;
        RECT 32.530 10.025 32.825 10.285 ;
        RECT 31.710 9.575 32.060 9.605 ;
        RECT 30.800 9.545 32.060 9.575 ;
        RECT 30.740 9.405 32.060 9.545 ;
        RECT 25.105 9.340 25.415 9.360 ;
        RECT 25.125 9.315 25.415 9.340 ;
        RECT 30.740 9.315 31.030 9.405 ;
        RECT 31.710 9.315 32.060 9.405 ;
        RECT 25.555 9.145 25.845 9.175 ;
        RECT 25.385 9.140 25.845 9.145 ;
        RECT 26.590 9.140 26.940 9.240 ;
        RECT 31.195 9.175 31.520 9.265 ;
        RECT 31.170 9.145 31.520 9.175 ;
        RECT 31.000 9.140 31.520 9.145 ;
        RECT 25.385 8.975 31.520 9.140 ;
        RECT 25.555 8.970 31.520 8.975 ;
        RECT 25.555 8.945 25.845 8.970 ;
        RECT 26.590 8.890 26.940 8.970 ;
        RECT 31.170 8.945 31.520 8.970 ;
        RECT 31.195 8.940 31.520 8.945 ;
        RECT 32.590 8.925 32.760 10.025 ;
        RECT 33.525 10.020 33.820 10.280 ;
        RECT 41.450 10.055 41.740 10.285 ;
        RECT 47.065 10.055 47.355 10.285 ;
        RECT 33.585 9.290 33.755 10.020 ;
        RECT 41.510 9.710 41.680 10.055 ;
        RECT 41.430 9.360 41.800 9.710 ;
        RECT 47.125 9.575 47.295 10.055 ;
        RECT 48.855 10.025 49.150 10.285 ;
        RECT 48.035 9.575 48.385 9.605 ;
        RECT 47.125 9.545 48.385 9.575 ;
        RECT 47.065 9.405 48.385 9.545 ;
        RECT 41.430 9.340 41.740 9.360 ;
        RECT 41.450 9.315 41.740 9.340 ;
        RECT 47.065 9.315 47.355 9.405 ;
        RECT 48.035 9.315 48.385 9.405 ;
        RECT 32.530 8.920 32.760 8.925 ;
        RECT 33.575 8.940 33.925 9.290 ;
        RECT 42.080 9.175 42.430 9.245 ;
        RECT 47.520 9.175 47.845 9.265 ;
        RECT 41.880 9.145 42.430 9.175 ;
        RECT 47.495 9.145 47.845 9.175 ;
        RECT 41.710 9.140 42.430 9.145 ;
        RECT 47.325 9.140 47.845 9.145 ;
        RECT 41.710 8.975 47.845 9.140 ;
        RECT 41.880 8.970 47.845 8.975 ;
        RECT 41.880 8.945 42.430 8.970 ;
        RECT 47.495 8.945 47.845 8.970 ;
        RECT 33.575 8.920 33.875 8.940 ;
        RECT 16.140 8.785 16.490 8.860 ;
        RECT 30.395 8.815 30.715 8.830 ;
        RECT 30.370 8.785 30.715 8.815 ;
        RECT 16.000 8.615 16.490 8.785 ;
        RECT 30.195 8.615 30.715 8.785 ;
        RECT 32.530 8.685 32.820 8.920 ;
        RECT 33.525 8.835 33.875 8.920 ;
        RECT 42.080 8.895 42.430 8.945 ;
        RECT 47.520 8.940 47.845 8.945 ;
        RECT 48.915 8.925 49.085 10.025 ;
        RECT 49.850 10.020 50.145 10.280 ;
        RECT 57.775 10.055 58.065 10.285 ;
        RECT 63.390 10.055 63.680 10.285 ;
        RECT 49.910 9.300 50.080 10.020 ;
        RECT 57.835 9.710 58.005 10.055 ;
        RECT 57.755 9.360 58.125 9.710 ;
        RECT 63.450 9.575 63.620 10.055 ;
        RECT 65.180 10.025 65.475 10.285 ;
        RECT 64.360 9.575 64.710 9.605 ;
        RECT 63.450 9.545 64.710 9.575 ;
        RECT 63.390 9.405 64.710 9.545 ;
        RECT 57.755 9.340 58.065 9.360 ;
        RECT 57.775 9.315 58.065 9.340 ;
        RECT 63.390 9.315 63.680 9.405 ;
        RECT 64.360 9.315 64.710 9.405 ;
        RECT 48.855 8.920 49.085 8.925 ;
        RECT 49.895 8.945 50.250 9.300 ;
        RECT 58.405 9.175 58.755 9.250 ;
        RECT 63.845 9.175 64.170 9.265 ;
        RECT 58.205 9.145 58.755 9.175 ;
        RECT 63.820 9.145 64.170 9.175 ;
        RECT 58.035 9.140 58.755 9.145 ;
        RECT 63.650 9.140 64.170 9.145 ;
        RECT 58.035 8.975 64.170 9.140 ;
        RECT 58.205 8.970 64.170 8.975 ;
        RECT 58.205 8.945 58.755 8.970 ;
        RECT 63.820 8.945 64.170 8.970 ;
        RECT 49.895 8.920 50.200 8.945 ;
        RECT 33.525 8.680 33.815 8.835 ;
        RECT 46.720 8.815 47.040 8.830 ;
        RECT 46.695 8.785 47.040 8.815 ;
        RECT 46.520 8.615 47.040 8.785 ;
        RECT 48.855 8.685 49.145 8.920 ;
        RECT 49.850 8.840 50.200 8.920 ;
        RECT 58.405 8.900 58.755 8.945 ;
        RECT 63.845 8.940 64.170 8.945 ;
        RECT 65.240 8.925 65.410 10.025 ;
        RECT 66.175 10.020 66.470 10.280 ;
        RECT 74.100 10.055 74.390 10.285 ;
        RECT 79.715 10.055 80.005 10.285 ;
        RECT 66.235 9.290 66.405 10.020 ;
        RECT 74.160 9.710 74.330 10.055 ;
        RECT 74.080 9.360 74.450 9.710 ;
        RECT 79.775 9.575 79.945 10.055 ;
        RECT 81.505 10.025 81.800 10.285 ;
        RECT 80.685 9.575 81.035 9.605 ;
        RECT 79.775 9.545 81.035 9.575 ;
        RECT 79.715 9.405 81.035 9.545 ;
        RECT 74.080 9.340 74.390 9.360 ;
        RECT 74.100 9.315 74.390 9.340 ;
        RECT 79.715 9.315 80.005 9.405 ;
        RECT 80.685 9.315 81.035 9.405 ;
        RECT 65.180 8.920 65.410 8.925 ;
        RECT 66.180 8.940 66.530 9.290 ;
        RECT 74.730 9.175 75.080 9.245 ;
        RECT 80.170 9.175 80.495 9.265 ;
        RECT 74.530 9.145 75.080 9.175 ;
        RECT 80.145 9.145 80.495 9.175 ;
        RECT 74.360 9.140 75.080 9.145 ;
        RECT 79.975 9.140 80.495 9.145 ;
        RECT 74.360 8.975 80.495 9.140 ;
        RECT 74.530 8.970 80.495 8.975 ;
        RECT 74.530 8.945 75.080 8.970 ;
        RECT 80.145 8.945 80.495 8.970 ;
        RECT 66.180 8.920 66.525 8.940 ;
        RECT 49.850 8.680 50.140 8.840 ;
        RECT 63.045 8.815 63.365 8.830 ;
        RECT 63.020 8.785 63.365 8.815 ;
        RECT 62.845 8.615 63.365 8.785 ;
        RECT 65.180 8.685 65.470 8.920 ;
        RECT 66.175 8.840 66.525 8.920 ;
        RECT 74.730 8.895 75.080 8.945 ;
        RECT 80.170 8.940 80.495 8.945 ;
        RECT 81.565 8.925 81.735 10.025 ;
        RECT 82.500 10.020 82.795 10.280 ;
        RECT 90.425 10.055 90.715 10.285 ;
        RECT 96.040 10.055 96.330 10.285 ;
        RECT 82.560 9.290 82.730 10.020 ;
        RECT 90.485 9.710 90.655 10.055 ;
        RECT 90.405 9.360 90.775 9.710 ;
        RECT 96.100 9.575 96.270 10.055 ;
        RECT 97.830 10.025 98.125 10.285 ;
        RECT 97.010 9.575 97.360 9.605 ;
        RECT 96.100 9.545 97.360 9.575 ;
        RECT 96.040 9.405 97.360 9.545 ;
        RECT 90.405 9.340 90.715 9.360 ;
        RECT 90.425 9.315 90.715 9.340 ;
        RECT 96.040 9.315 96.330 9.405 ;
        RECT 97.010 9.315 97.360 9.405 ;
        RECT 81.505 8.920 81.735 8.925 ;
        RECT 82.505 8.940 82.855 9.290 ;
        RECT 91.060 9.175 91.410 9.245 ;
        RECT 96.495 9.175 96.820 9.265 ;
        RECT 90.855 9.145 91.410 9.175 ;
        RECT 96.470 9.145 96.820 9.175 ;
        RECT 90.685 9.140 91.410 9.145 ;
        RECT 96.300 9.140 96.820 9.145 ;
        RECT 90.685 8.975 96.820 9.140 ;
        RECT 90.855 8.970 96.820 8.975 ;
        RECT 90.855 8.945 91.410 8.970 ;
        RECT 96.470 8.945 96.820 8.970 ;
        RECT 82.505 8.920 82.850 8.940 ;
        RECT 66.175 8.680 66.465 8.840 ;
        RECT 79.370 8.815 79.690 8.830 ;
        RECT 79.345 8.785 79.690 8.815 ;
        RECT 79.170 8.615 79.690 8.785 ;
        RECT 81.505 8.685 81.795 8.920 ;
        RECT 82.500 8.845 82.850 8.920 ;
        RECT 91.060 8.895 91.410 8.945 ;
        RECT 96.495 8.940 96.820 8.945 ;
        RECT 97.890 8.925 98.060 10.025 ;
        RECT 98.825 10.020 99.120 10.280 ;
        RECT 98.855 10.005 99.120 10.020 ;
        RECT 98.855 9.910 99.180 10.005 ;
        RECT 98.855 9.560 99.205 9.910 ;
        RECT 97.830 8.920 98.060 8.925 ;
        RECT 98.885 8.920 99.055 9.560 ;
        RECT 82.500 8.680 82.790 8.845 ;
        RECT 95.695 8.815 96.015 8.830 ;
        RECT 95.670 8.785 96.015 8.815 ;
        RECT 95.495 8.615 96.015 8.785 ;
        RECT 97.830 8.685 98.120 8.920 ;
        RECT 98.825 8.915 99.055 8.920 ;
        RECT 98.825 8.680 99.115 8.915 ;
        RECT 16.140 8.570 16.490 8.615 ;
        RECT 30.370 8.585 30.715 8.615 ;
        RECT 46.695 8.585 47.040 8.615 ;
        RECT 63.020 8.585 63.365 8.615 ;
        RECT 79.345 8.585 79.690 8.615 ;
        RECT 95.670 8.585 96.015 8.615 ;
        RECT 30.395 8.540 30.715 8.585 ;
        RECT 46.720 8.540 47.040 8.585 ;
        RECT 63.045 8.540 63.365 8.585 ;
        RECT 79.370 8.540 79.690 8.585 ;
        RECT 95.695 8.540 96.015 8.585 ;
        RECT 19.290 5.065 19.580 5.105 ;
        RECT 19.990 5.065 20.310 5.125 ;
        RECT 19.290 4.925 20.310 5.065 ;
        RECT 19.290 4.875 19.620 4.925 ;
        RECT 19.990 4.865 20.310 4.925 ;
        RECT 25.130 5.065 25.420 5.105 ;
        RECT 25.130 4.875 25.460 5.065 ;
        RECT 20.490 4.785 20.780 4.825 ;
        RECT 21.710 4.785 22.030 4.845 ;
        RECT 22.550 4.825 22.870 4.845 ;
        RECT 22.550 4.785 22.980 4.825 ;
        RECT 20.490 4.595 20.940 4.785 ;
        RECT 18.790 4.305 19.110 4.565 ;
        RECT 19.750 4.545 20.070 4.565 ;
        RECT 19.750 4.315 20.300 4.545 ;
        RECT 20.800 4.365 20.940 4.595 ;
        RECT 21.710 4.645 22.980 4.785 ;
        RECT 21.710 4.585 22.030 4.645 ;
        RECT 22.550 4.595 22.980 4.645 ;
        RECT 22.550 4.585 22.870 4.595 ;
        RECT 19.750 4.305 20.070 4.315 ;
        RECT 18.880 3.385 19.020 4.305 ;
        RECT 20.440 4.225 20.940 4.365 ;
        RECT 21.250 4.315 21.540 4.545 ;
        RECT 19.750 3.985 20.070 4.005 ;
        RECT 19.750 3.755 20.300 3.985 ;
        RECT 19.750 3.745 20.070 3.755 ;
        RECT 20.440 3.445 20.580 4.225 ;
        RECT 21.320 4.005 21.460 4.315 ;
        RECT 22.520 4.265 25.100 4.365 ;
        RECT 22.450 4.225 25.180 4.265 ;
        RECT 22.450 4.035 23.110 4.225 ;
        RECT 24.890 4.035 25.180 4.225 ;
        RECT 22.790 4.025 23.110 4.035 ;
        RECT 20.970 3.985 21.460 4.005 ;
        RECT 20.730 3.755 21.460 3.985 ;
        RECT 20.970 3.745 21.460 3.755 ;
        RECT 21.950 3.745 22.270 4.005 ;
        RECT 23.790 3.985 24.110 4.005 ;
        RECT 23.790 3.755 24.220 3.985 ;
        RECT 23.790 3.745 24.110 3.755 ;
        RECT 24.390 3.745 24.710 4.005 ;
        RECT 19.290 3.385 19.580 3.425 ;
        RECT 18.880 3.245 19.580 3.385 ;
        RECT 19.290 3.195 19.580 3.245 ;
        RECT 20.230 3.245 20.580 3.445 ;
        RECT 21.320 3.385 21.460 3.745 ;
        RECT 22.430 3.665 22.750 3.725 ;
        RECT 25.320 3.705 25.460 4.875 ;
        RECT 26.130 4.845 26.420 5.105 ;
        RECT 35.615 5.065 35.905 5.105 ;
        RECT 36.315 5.065 36.635 5.125 ;
        RECT 35.615 4.925 36.635 5.065 ;
        RECT 35.615 4.875 35.945 4.925 ;
        RECT 36.315 4.865 36.635 4.925 ;
        RECT 41.455 5.065 41.745 5.105 ;
        RECT 41.455 4.875 41.785 5.065 ;
        RECT 26.110 4.585 26.430 4.845 ;
        RECT 36.815 4.785 37.105 4.825 ;
        RECT 38.035 4.785 38.355 4.845 ;
        RECT 38.875 4.825 39.195 4.845 ;
        RECT 38.875 4.785 39.305 4.825 ;
        RECT 36.815 4.595 37.265 4.785 ;
        RECT 35.115 4.305 35.435 4.565 ;
        RECT 36.075 4.545 36.395 4.565 ;
        RECT 36.075 4.315 36.625 4.545 ;
        RECT 37.125 4.365 37.265 4.595 ;
        RECT 38.035 4.645 39.305 4.785 ;
        RECT 38.035 4.585 38.355 4.645 ;
        RECT 38.875 4.595 39.305 4.645 ;
        RECT 38.875 4.585 39.195 4.595 ;
        RECT 36.075 4.305 36.395 4.315 ;
        RECT 26.230 3.985 26.550 4.005 ;
        RECT 26.230 3.745 26.700 3.985 ;
        RECT 26.850 3.945 27.140 3.985 ;
        RECT 26.850 3.805 27.300 3.945 ;
        RECT 30.395 3.875 30.715 3.945 ;
        RECT 30.370 3.845 30.715 3.875 ;
        RECT 26.850 3.755 27.780 3.805 ;
        RECT 22.930 3.665 23.220 3.705 ;
        RECT 25.320 3.665 25.660 3.705 ;
        RECT 22.430 3.525 23.220 3.665 ;
        RECT 22.430 3.465 22.750 3.525 ;
        RECT 22.930 3.475 23.220 3.525 ;
        RECT 24.960 3.525 25.660 3.665 ;
        RECT 24.960 3.505 25.100 3.525 ;
        RECT 23.500 3.445 25.100 3.505 ;
        RECT 25.370 3.475 25.660 3.525 ;
        RECT 26.560 3.505 26.700 3.745 ;
        RECT 27.160 3.725 27.780 3.755 ;
        RECT 27.160 3.665 27.870 3.725 ;
        RECT 30.195 3.675 30.715 3.845 ;
        RECT 21.730 3.385 22.020 3.425 ;
        RECT 21.320 3.245 22.020 3.385 ;
        RECT 20.230 3.185 20.550 3.245 ;
        RECT 21.730 3.195 22.020 3.245 ;
        RECT 23.410 3.365 25.100 3.445 ;
        RECT 25.850 3.425 26.170 3.445 ;
        RECT 23.410 3.195 23.980 3.365 ;
        RECT 25.850 3.195 26.420 3.425 ;
        RECT 26.560 3.385 26.820 3.505 ;
        RECT 27.550 3.465 27.870 3.665 ;
        RECT 30.370 3.645 30.715 3.675 ;
        RECT 31.170 3.490 31.520 3.610 ;
        RECT 32.530 3.540 32.820 3.775 ;
        RECT 32.530 3.535 32.760 3.540 ;
        RECT 27.090 3.385 27.380 3.425 ;
        RECT 26.560 3.365 27.380 3.385 ;
        RECT 26.680 3.245 27.380 3.365 ;
        RECT 27.090 3.195 27.380 3.245 ;
        RECT 28.865 3.320 31.520 3.490 ;
        RECT 23.410 3.185 23.730 3.195 ;
        RECT 25.850 3.185 26.170 3.195 ;
        RECT 28.865 3.105 29.035 3.320 ;
        RECT 31.000 3.315 31.520 3.320 ;
        RECT 31.170 3.260 31.520 3.315 ;
        RECT 30.740 3.120 31.030 3.145 ;
        RECT 31.710 3.120 32.060 3.145 ;
        RECT 28.775 2.755 29.115 3.105 ;
        RECT 30.740 2.950 32.060 3.120 ;
        RECT 30.740 2.915 31.030 2.950 ;
        RECT 30.800 2.405 30.970 2.915 ;
        RECT 31.710 2.855 32.060 2.950 ;
        RECT 32.590 2.435 32.760 3.535 ;
        RECT 35.205 3.385 35.345 4.305 ;
        RECT 36.765 4.225 37.265 4.365 ;
        RECT 37.575 4.315 37.865 4.545 ;
        RECT 36.075 3.985 36.395 4.005 ;
        RECT 36.075 3.755 36.625 3.985 ;
        RECT 36.075 3.745 36.395 3.755 ;
        RECT 36.765 3.445 36.905 4.225 ;
        RECT 37.645 4.005 37.785 4.315 ;
        RECT 38.845 4.265 41.425 4.365 ;
        RECT 38.775 4.225 41.505 4.265 ;
        RECT 38.775 4.035 39.435 4.225 ;
        RECT 41.215 4.035 41.505 4.225 ;
        RECT 39.115 4.025 39.435 4.035 ;
        RECT 37.295 3.985 37.785 4.005 ;
        RECT 37.055 3.755 37.785 3.985 ;
        RECT 37.295 3.745 37.785 3.755 ;
        RECT 38.275 3.745 38.595 4.005 ;
        RECT 40.115 3.985 40.435 4.005 ;
        RECT 40.115 3.755 40.545 3.985 ;
        RECT 40.115 3.745 40.435 3.755 ;
        RECT 40.715 3.745 41.035 4.005 ;
        RECT 35.615 3.385 35.905 3.425 ;
        RECT 35.205 3.245 35.905 3.385 ;
        RECT 35.615 3.195 35.905 3.245 ;
        RECT 36.555 3.245 36.905 3.445 ;
        RECT 37.645 3.385 37.785 3.745 ;
        RECT 38.755 3.665 39.075 3.725 ;
        RECT 41.645 3.705 41.785 4.875 ;
        RECT 42.455 4.845 42.745 5.105 ;
        RECT 51.940 5.065 52.230 5.105 ;
        RECT 52.640 5.065 52.960 5.125 ;
        RECT 51.940 4.925 52.960 5.065 ;
        RECT 51.940 4.875 52.270 4.925 ;
        RECT 52.640 4.865 52.960 4.925 ;
        RECT 57.780 5.065 58.070 5.105 ;
        RECT 57.780 4.875 58.110 5.065 ;
        RECT 42.435 4.585 42.755 4.845 ;
        RECT 53.140 4.785 53.430 4.825 ;
        RECT 54.360 4.785 54.680 4.845 ;
        RECT 55.200 4.825 55.520 4.845 ;
        RECT 55.200 4.785 55.630 4.825 ;
        RECT 53.140 4.595 53.590 4.785 ;
        RECT 51.440 4.305 51.760 4.565 ;
        RECT 52.400 4.545 52.720 4.565 ;
        RECT 52.400 4.315 52.950 4.545 ;
        RECT 53.450 4.365 53.590 4.595 ;
        RECT 54.360 4.645 55.630 4.785 ;
        RECT 54.360 4.585 54.680 4.645 ;
        RECT 55.200 4.595 55.630 4.645 ;
        RECT 55.200 4.585 55.520 4.595 ;
        RECT 52.400 4.305 52.720 4.315 ;
        RECT 42.555 3.985 42.875 4.005 ;
        RECT 42.555 3.745 43.025 3.985 ;
        RECT 43.175 3.945 43.465 3.985 ;
        RECT 43.175 3.805 43.625 3.945 ;
        RECT 46.720 3.875 47.040 3.945 ;
        RECT 46.695 3.845 47.040 3.875 ;
        RECT 43.175 3.755 44.105 3.805 ;
        RECT 39.255 3.665 39.545 3.705 ;
        RECT 41.645 3.665 41.985 3.705 ;
        RECT 38.755 3.525 39.545 3.665 ;
        RECT 38.755 3.465 39.075 3.525 ;
        RECT 39.255 3.475 39.545 3.525 ;
        RECT 41.285 3.525 41.985 3.665 ;
        RECT 41.285 3.505 41.425 3.525 ;
        RECT 39.825 3.445 41.425 3.505 ;
        RECT 41.695 3.475 41.985 3.525 ;
        RECT 42.885 3.505 43.025 3.745 ;
        RECT 43.485 3.725 44.105 3.755 ;
        RECT 43.485 3.665 44.195 3.725 ;
        RECT 46.520 3.675 47.040 3.845 ;
        RECT 38.055 3.385 38.345 3.425 ;
        RECT 37.645 3.245 38.345 3.385 ;
        RECT 36.555 3.185 36.875 3.245 ;
        RECT 38.055 3.195 38.345 3.245 ;
        RECT 39.735 3.365 41.425 3.445 ;
        RECT 42.175 3.425 42.495 3.445 ;
        RECT 39.735 3.195 40.305 3.365 ;
        RECT 42.175 3.195 42.745 3.425 ;
        RECT 42.885 3.385 43.145 3.505 ;
        RECT 43.875 3.465 44.195 3.665 ;
        RECT 46.695 3.645 47.040 3.675 ;
        RECT 47.495 3.490 47.845 3.610 ;
        RECT 48.855 3.540 49.145 3.775 ;
        RECT 48.855 3.535 49.085 3.540 ;
        RECT 43.415 3.385 43.705 3.425 ;
        RECT 42.885 3.365 43.705 3.385 ;
        RECT 43.005 3.245 43.705 3.365 ;
        RECT 43.415 3.195 43.705 3.245 ;
        RECT 45.190 3.320 47.845 3.490 ;
        RECT 39.735 3.185 40.055 3.195 ;
        RECT 42.175 3.185 42.495 3.195 ;
        RECT 45.190 3.105 45.360 3.320 ;
        RECT 47.325 3.315 47.845 3.320 ;
        RECT 47.495 3.260 47.845 3.315 ;
        RECT 47.065 3.120 47.355 3.145 ;
        RECT 48.035 3.120 48.385 3.145 ;
        RECT 45.100 2.755 45.440 3.105 ;
        RECT 47.065 2.950 48.385 3.120 ;
        RECT 47.065 2.915 47.355 2.950 ;
        RECT 30.740 2.175 31.030 2.405 ;
        RECT 32.530 2.175 32.825 2.435 ;
        RECT 47.125 2.405 47.295 2.915 ;
        RECT 48.035 2.855 48.385 2.950 ;
        RECT 48.915 2.435 49.085 3.535 ;
        RECT 51.530 3.385 51.670 4.305 ;
        RECT 53.090 4.225 53.590 4.365 ;
        RECT 53.900 4.315 54.190 4.545 ;
        RECT 52.400 3.985 52.720 4.005 ;
        RECT 52.400 3.755 52.950 3.985 ;
        RECT 52.400 3.745 52.720 3.755 ;
        RECT 53.090 3.445 53.230 4.225 ;
        RECT 53.970 4.005 54.110 4.315 ;
        RECT 55.170 4.265 57.750 4.365 ;
        RECT 55.100 4.225 57.830 4.265 ;
        RECT 55.100 4.035 55.760 4.225 ;
        RECT 57.540 4.035 57.830 4.225 ;
        RECT 55.440 4.025 55.760 4.035 ;
        RECT 53.620 3.985 54.110 4.005 ;
        RECT 53.380 3.755 54.110 3.985 ;
        RECT 53.620 3.745 54.110 3.755 ;
        RECT 54.600 3.745 54.920 4.005 ;
        RECT 56.440 3.985 56.760 4.005 ;
        RECT 56.440 3.755 56.870 3.985 ;
        RECT 56.440 3.745 56.760 3.755 ;
        RECT 57.040 3.745 57.360 4.005 ;
        RECT 51.940 3.385 52.230 3.425 ;
        RECT 51.530 3.245 52.230 3.385 ;
        RECT 51.940 3.195 52.230 3.245 ;
        RECT 52.880 3.245 53.230 3.445 ;
        RECT 53.970 3.385 54.110 3.745 ;
        RECT 55.080 3.665 55.400 3.725 ;
        RECT 57.970 3.705 58.110 4.875 ;
        RECT 58.780 4.845 59.070 5.105 ;
        RECT 68.265 5.065 68.555 5.105 ;
        RECT 68.965 5.065 69.285 5.125 ;
        RECT 68.265 4.925 69.285 5.065 ;
        RECT 68.265 4.875 68.595 4.925 ;
        RECT 68.965 4.865 69.285 4.925 ;
        RECT 74.105 5.065 74.395 5.105 ;
        RECT 74.105 4.875 74.435 5.065 ;
        RECT 58.760 4.585 59.080 4.845 ;
        RECT 69.465 4.785 69.755 4.825 ;
        RECT 70.685 4.785 71.005 4.845 ;
        RECT 71.525 4.825 71.845 4.845 ;
        RECT 71.525 4.785 71.955 4.825 ;
        RECT 69.465 4.595 69.915 4.785 ;
        RECT 67.765 4.305 68.085 4.565 ;
        RECT 68.725 4.545 69.045 4.565 ;
        RECT 68.725 4.315 69.275 4.545 ;
        RECT 69.775 4.365 69.915 4.595 ;
        RECT 70.685 4.645 71.955 4.785 ;
        RECT 70.685 4.585 71.005 4.645 ;
        RECT 71.525 4.595 71.955 4.645 ;
        RECT 71.525 4.585 71.845 4.595 ;
        RECT 68.725 4.305 69.045 4.315 ;
        RECT 58.880 3.985 59.200 4.005 ;
        RECT 58.880 3.745 59.350 3.985 ;
        RECT 59.500 3.945 59.790 3.985 ;
        RECT 59.500 3.805 59.950 3.945 ;
        RECT 63.045 3.875 63.365 3.945 ;
        RECT 63.020 3.845 63.365 3.875 ;
        RECT 59.500 3.755 60.430 3.805 ;
        RECT 55.580 3.665 55.870 3.705 ;
        RECT 57.970 3.665 58.310 3.705 ;
        RECT 55.080 3.525 55.870 3.665 ;
        RECT 55.080 3.465 55.400 3.525 ;
        RECT 55.580 3.475 55.870 3.525 ;
        RECT 57.610 3.525 58.310 3.665 ;
        RECT 57.610 3.505 57.750 3.525 ;
        RECT 56.150 3.445 57.750 3.505 ;
        RECT 58.020 3.475 58.310 3.525 ;
        RECT 59.210 3.505 59.350 3.745 ;
        RECT 59.810 3.725 60.430 3.755 ;
        RECT 59.810 3.665 60.520 3.725 ;
        RECT 62.845 3.675 63.365 3.845 ;
        RECT 54.380 3.385 54.670 3.425 ;
        RECT 53.970 3.245 54.670 3.385 ;
        RECT 52.880 3.185 53.200 3.245 ;
        RECT 54.380 3.195 54.670 3.245 ;
        RECT 56.060 3.365 57.750 3.445 ;
        RECT 58.500 3.425 58.820 3.445 ;
        RECT 56.060 3.195 56.630 3.365 ;
        RECT 58.500 3.195 59.070 3.425 ;
        RECT 59.210 3.385 59.470 3.505 ;
        RECT 60.200 3.465 60.520 3.665 ;
        RECT 63.020 3.645 63.365 3.675 ;
        RECT 63.820 3.490 64.170 3.610 ;
        RECT 65.180 3.540 65.470 3.775 ;
        RECT 65.180 3.535 65.410 3.540 ;
        RECT 59.740 3.385 60.030 3.425 ;
        RECT 59.210 3.365 60.030 3.385 ;
        RECT 59.330 3.245 60.030 3.365 ;
        RECT 59.740 3.195 60.030 3.245 ;
        RECT 61.515 3.320 64.170 3.490 ;
        RECT 56.060 3.185 56.380 3.195 ;
        RECT 58.500 3.185 58.820 3.195 ;
        RECT 61.515 3.105 61.685 3.320 ;
        RECT 63.650 3.315 64.170 3.320 ;
        RECT 63.820 3.260 64.170 3.315 ;
        RECT 63.390 3.120 63.680 3.145 ;
        RECT 64.360 3.120 64.710 3.145 ;
        RECT 61.425 2.755 61.765 3.105 ;
        RECT 63.390 2.950 64.710 3.120 ;
        RECT 63.390 2.915 63.680 2.950 ;
        RECT 47.065 2.175 47.355 2.405 ;
        RECT 48.855 2.175 49.150 2.435 ;
        RECT 63.450 2.405 63.620 2.915 ;
        RECT 64.360 2.855 64.710 2.950 ;
        RECT 65.240 2.435 65.410 3.535 ;
        RECT 67.855 3.385 67.995 4.305 ;
        RECT 69.415 4.225 69.915 4.365 ;
        RECT 70.225 4.315 70.515 4.545 ;
        RECT 68.725 3.985 69.045 4.005 ;
        RECT 68.725 3.755 69.275 3.985 ;
        RECT 68.725 3.745 69.045 3.755 ;
        RECT 69.415 3.445 69.555 4.225 ;
        RECT 70.295 4.005 70.435 4.315 ;
        RECT 71.495 4.265 74.075 4.365 ;
        RECT 71.425 4.225 74.155 4.265 ;
        RECT 71.425 4.035 72.085 4.225 ;
        RECT 73.865 4.035 74.155 4.225 ;
        RECT 71.765 4.025 72.085 4.035 ;
        RECT 69.945 3.985 70.435 4.005 ;
        RECT 69.705 3.755 70.435 3.985 ;
        RECT 69.945 3.745 70.435 3.755 ;
        RECT 70.925 3.745 71.245 4.005 ;
        RECT 72.765 3.985 73.085 4.005 ;
        RECT 72.765 3.755 73.195 3.985 ;
        RECT 72.765 3.745 73.085 3.755 ;
        RECT 73.365 3.745 73.685 4.005 ;
        RECT 68.265 3.385 68.555 3.425 ;
        RECT 67.855 3.245 68.555 3.385 ;
        RECT 68.265 3.195 68.555 3.245 ;
        RECT 69.205 3.245 69.555 3.445 ;
        RECT 70.295 3.385 70.435 3.745 ;
        RECT 71.405 3.665 71.725 3.725 ;
        RECT 74.295 3.705 74.435 4.875 ;
        RECT 75.105 4.845 75.395 5.105 ;
        RECT 84.590 5.065 84.880 5.105 ;
        RECT 85.290 5.065 85.610 5.125 ;
        RECT 84.590 4.925 85.610 5.065 ;
        RECT 84.590 4.875 84.920 4.925 ;
        RECT 85.290 4.865 85.610 4.925 ;
        RECT 90.430 5.065 90.720 5.105 ;
        RECT 90.430 4.875 90.760 5.065 ;
        RECT 75.085 4.585 75.405 4.845 ;
        RECT 85.790 4.785 86.080 4.825 ;
        RECT 87.010 4.785 87.330 4.845 ;
        RECT 87.850 4.825 88.170 4.845 ;
        RECT 87.850 4.785 88.280 4.825 ;
        RECT 85.790 4.595 86.240 4.785 ;
        RECT 84.090 4.305 84.410 4.565 ;
        RECT 85.050 4.545 85.370 4.565 ;
        RECT 85.050 4.315 85.600 4.545 ;
        RECT 86.100 4.365 86.240 4.595 ;
        RECT 87.010 4.645 88.280 4.785 ;
        RECT 87.010 4.585 87.330 4.645 ;
        RECT 87.850 4.595 88.280 4.645 ;
        RECT 87.850 4.585 88.170 4.595 ;
        RECT 85.050 4.305 85.370 4.315 ;
        RECT 75.205 3.985 75.525 4.005 ;
        RECT 75.205 3.745 75.675 3.985 ;
        RECT 75.825 3.945 76.115 3.985 ;
        RECT 75.825 3.805 76.275 3.945 ;
        RECT 79.370 3.875 79.690 3.945 ;
        RECT 79.345 3.845 79.690 3.875 ;
        RECT 75.825 3.755 76.755 3.805 ;
        RECT 71.905 3.665 72.195 3.705 ;
        RECT 74.295 3.665 74.635 3.705 ;
        RECT 71.405 3.525 72.195 3.665 ;
        RECT 71.405 3.465 71.725 3.525 ;
        RECT 71.905 3.475 72.195 3.525 ;
        RECT 73.935 3.525 74.635 3.665 ;
        RECT 73.935 3.505 74.075 3.525 ;
        RECT 72.475 3.445 74.075 3.505 ;
        RECT 74.345 3.475 74.635 3.525 ;
        RECT 75.535 3.505 75.675 3.745 ;
        RECT 76.135 3.725 76.755 3.755 ;
        RECT 76.135 3.665 76.845 3.725 ;
        RECT 79.170 3.675 79.690 3.845 ;
        RECT 70.705 3.385 70.995 3.425 ;
        RECT 70.295 3.245 70.995 3.385 ;
        RECT 69.205 3.185 69.525 3.245 ;
        RECT 70.705 3.195 70.995 3.245 ;
        RECT 72.385 3.365 74.075 3.445 ;
        RECT 74.825 3.425 75.145 3.445 ;
        RECT 72.385 3.195 72.955 3.365 ;
        RECT 74.825 3.195 75.395 3.425 ;
        RECT 75.535 3.385 75.795 3.505 ;
        RECT 76.525 3.465 76.845 3.665 ;
        RECT 79.345 3.645 79.690 3.675 ;
        RECT 80.145 3.490 80.495 3.610 ;
        RECT 81.505 3.540 81.795 3.775 ;
        RECT 81.505 3.535 81.735 3.540 ;
        RECT 76.065 3.385 76.355 3.425 ;
        RECT 75.535 3.365 76.355 3.385 ;
        RECT 75.655 3.245 76.355 3.365 ;
        RECT 76.065 3.195 76.355 3.245 ;
        RECT 77.840 3.320 80.495 3.490 ;
        RECT 72.385 3.185 72.705 3.195 ;
        RECT 74.825 3.185 75.145 3.195 ;
        RECT 77.840 3.105 78.010 3.320 ;
        RECT 79.975 3.315 80.495 3.320 ;
        RECT 80.145 3.260 80.495 3.315 ;
        RECT 79.715 3.120 80.005 3.145 ;
        RECT 80.685 3.120 81.035 3.145 ;
        RECT 77.750 2.755 78.090 3.105 ;
        RECT 79.715 2.950 81.035 3.120 ;
        RECT 79.715 2.915 80.005 2.950 ;
        RECT 63.390 2.175 63.680 2.405 ;
        RECT 65.180 2.175 65.475 2.435 ;
        RECT 79.775 2.405 79.945 2.915 ;
        RECT 80.685 2.855 81.035 2.950 ;
        RECT 81.565 2.435 81.735 3.535 ;
        RECT 84.180 3.385 84.320 4.305 ;
        RECT 85.740 4.225 86.240 4.365 ;
        RECT 86.550 4.315 86.840 4.545 ;
        RECT 85.050 3.985 85.370 4.005 ;
        RECT 85.050 3.755 85.600 3.985 ;
        RECT 85.050 3.745 85.370 3.755 ;
        RECT 85.740 3.445 85.880 4.225 ;
        RECT 86.620 4.005 86.760 4.315 ;
        RECT 87.820 4.265 90.400 4.365 ;
        RECT 87.750 4.225 90.480 4.265 ;
        RECT 87.750 4.035 88.410 4.225 ;
        RECT 90.190 4.035 90.480 4.225 ;
        RECT 88.090 4.025 88.410 4.035 ;
        RECT 86.270 3.985 86.760 4.005 ;
        RECT 86.030 3.755 86.760 3.985 ;
        RECT 86.270 3.745 86.760 3.755 ;
        RECT 87.250 3.745 87.570 4.005 ;
        RECT 89.090 3.985 89.410 4.005 ;
        RECT 89.090 3.755 89.520 3.985 ;
        RECT 89.090 3.745 89.410 3.755 ;
        RECT 89.690 3.745 90.010 4.005 ;
        RECT 84.590 3.385 84.880 3.425 ;
        RECT 84.180 3.245 84.880 3.385 ;
        RECT 84.590 3.195 84.880 3.245 ;
        RECT 85.530 3.245 85.880 3.445 ;
        RECT 86.620 3.385 86.760 3.745 ;
        RECT 87.730 3.665 88.050 3.725 ;
        RECT 90.620 3.705 90.760 4.875 ;
        RECT 91.430 4.845 91.720 5.105 ;
        RECT 91.410 4.585 91.730 4.845 ;
        RECT 91.530 3.985 91.850 4.005 ;
        RECT 91.530 3.745 92.000 3.985 ;
        RECT 92.150 3.945 92.440 3.985 ;
        RECT 92.150 3.805 92.600 3.945 ;
        RECT 95.695 3.875 96.015 3.945 ;
        RECT 95.670 3.845 96.015 3.875 ;
        RECT 92.150 3.755 93.080 3.805 ;
        RECT 88.230 3.665 88.520 3.705 ;
        RECT 90.620 3.665 90.960 3.705 ;
        RECT 87.730 3.525 88.520 3.665 ;
        RECT 87.730 3.465 88.050 3.525 ;
        RECT 88.230 3.475 88.520 3.525 ;
        RECT 90.260 3.525 90.960 3.665 ;
        RECT 90.260 3.505 90.400 3.525 ;
        RECT 88.800 3.445 90.400 3.505 ;
        RECT 90.670 3.475 90.960 3.525 ;
        RECT 91.860 3.505 92.000 3.745 ;
        RECT 92.460 3.725 93.080 3.755 ;
        RECT 92.460 3.665 93.170 3.725 ;
        RECT 95.495 3.675 96.015 3.845 ;
        RECT 87.030 3.385 87.320 3.425 ;
        RECT 86.620 3.245 87.320 3.385 ;
        RECT 85.530 3.185 85.850 3.245 ;
        RECT 87.030 3.195 87.320 3.245 ;
        RECT 88.710 3.365 90.400 3.445 ;
        RECT 91.150 3.425 91.470 3.445 ;
        RECT 88.710 3.195 89.280 3.365 ;
        RECT 91.150 3.195 91.720 3.425 ;
        RECT 91.860 3.385 92.120 3.505 ;
        RECT 92.850 3.465 93.170 3.665 ;
        RECT 95.670 3.645 96.015 3.675 ;
        RECT 96.470 3.490 96.820 3.610 ;
        RECT 97.830 3.540 98.120 3.775 ;
        RECT 97.830 3.535 98.060 3.540 ;
        RECT 92.390 3.385 92.680 3.425 ;
        RECT 91.860 3.365 92.680 3.385 ;
        RECT 91.980 3.245 92.680 3.365 ;
        RECT 92.390 3.195 92.680 3.245 ;
        RECT 94.165 3.320 96.820 3.490 ;
        RECT 88.710 3.185 89.030 3.195 ;
        RECT 91.150 3.185 91.470 3.195 ;
        RECT 94.165 3.105 94.335 3.320 ;
        RECT 96.300 3.315 96.820 3.320 ;
        RECT 96.470 3.260 96.820 3.315 ;
        RECT 96.040 3.120 96.330 3.145 ;
        RECT 97.010 3.120 97.360 3.145 ;
        RECT 94.075 2.755 94.415 3.105 ;
        RECT 96.040 2.950 97.360 3.120 ;
        RECT 96.040 2.915 96.330 2.950 ;
        RECT 79.715 2.175 80.005 2.405 ;
        RECT 81.505 2.175 81.800 2.435 ;
        RECT 96.100 2.405 96.270 2.915 ;
        RECT 97.010 2.855 97.360 2.950 ;
        RECT 97.890 2.435 98.060 3.535 ;
        RECT 96.040 2.175 96.330 2.405 ;
        RECT 97.830 2.175 98.125 2.435 ;
      LAYER met2 ;
        RECT 16.230 10.685 99.055 10.855 ;
        RECT 16.230 8.890 16.400 10.685 ;
        RECT 98.885 9.910 99.055 10.685 ;
        RECT 16.545 9.515 16.835 9.635 ;
        RECT 16.545 9.510 16.920 9.515 ;
        RECT 16.545 9.335 17.830 9.510 ;
        RECT 25.105 9.340 25.475 9.710 ;
        RECT 41.430 9.340 41.800 9.710 ;
        RECT 57.755 9.340 58.125 9.710 ;
        RECT 74.080 9.340 74.450 9.710 ;
        RECT 90.405 9.340 90.775 9.710 ;
        RECT 98.855 9.560 99.205 9.910 ;
        RECT 16.545 9.285 16.835 9.335 ;
        RECT 17.655 9.145 17.830 9.335 ;
        RECT 26.590 9.145 26.940 9.240 ;
        RECT 31.195 9.200 31.520 9.265 ;
        RECT 17.655 8.970 26.940 9.145 ;
        RECT 26.590 8.890 26.940 8.970 ;
        RECT 30.080 9.030 31.520 9.200 ;
        RECT 16.170 8.540 16.460 8.890 ;
        RECT 19.600 5.295 23.260 5.435 ;
        RECT 18.810 4.245 19.090 4.620 ;
        RECT 19.600 4.615 19.740 5.295 ;
        RECT 20.020 5.065 20.280 5.155 ;
        RECT 20.020 4.925 21.700 5.065 ;
        RECT 20.020 4.835 20.280 4.925 ;
        RECT 21.560 4.875 21.700 4.925 ;
        RECT 21.560 4.645 22.000 4.875 ;
        RECT 19.600 4.365 20.050 4.615 ;
        RECT 21.740 4.555 22.000 4.645 ;
        RECT 22.520 4.555 22.840 4.875 ;
        RECT 23.120 4.615 23.260 5.295 ;
        RECT 23.430 5.065 23.710 5.180 ;
        RECT 24.510 5.065 26.690 5.175 ;
        RECT 23.430 5.015 26.690 5.065 ;
        RECT 23.430 4.925 24.650 5.015 ;
        RECT 23.430 4.805 23.710 4.925 ;
        RECT 25.350 4.615 25.650 4.620 ;
        RECT 19.770 4.245 20.050 4.365 ;
        RECT 21.060 4.060 21.460 4.225 ;
        RECT 21.060 4.035 21.530 4.060 ;
        RECT 19.780 3.945 20.040 4.035 ;
        RECT 19.780 3.805 20.820 3.945 ;
        RECT 19.780 3.715 20.040 3.805 ;
        RECT 20.250 3.125 20.530 3.500 ;
        RECT 20.680 3.155 20.820 3.805 ;
        RECT 21.000 3.715 21.530 4.035 ;
        RECT 21.250 3.685 21.530 3.715 ;
        RECT 21.970 3.685 22.250 4.060 ;
        RECT 22.520 3.755 22.660 4.555 ;
        RECT 23.120 4.505 25.650 4.615 ;
        RECT 26.140 4.555 26.400 4.875 ;
        RECT 26.140 4.505 26.340 4.555 ;
        RECT 23.120 4.475 26.340 4.505 ;
        RECT 25.370 4.365 26.340 4.475 ;
        RECT 22.820 4.225 23.080 4.315 ;
        RECT 25.370 4.245 25.650 4.365 ;
        RECT 22.820 4.060 23.140 4.225 ;
        RECT 22.820 3.995 23.210 4.060 ;
        RECT 22.460 3.435 22.720 3.755 ;
        RECT 22.930 3.685 23.210 3.995 ;
        RECT 23.810 3.685 24.090 4.060 ;
        RECT 24.420 3.715 24.680 4.035 ;
        RECT 23.440 3.155 23.700 3.475 ;
        RECT 20.290 2.735 20.460 3.125 ;
        RECT 20.680 3.015 23.640 3.155 ;
        RECT 24.480 3.015 24.620 3.715 ;
        RECT 25.490 3.685 25.770 4.055 ;
        RECT 25.560 3.015 25.700 3.685 ;
        RECT 25.940 3.475 26.080 4.365 ;
        RECT 26.540 4.035 26.690 5.015 ;
        RECT 26.260 3.895 26.690 4.035 ;
        RECT 26.260 3.715 26.520 3.895 ;
        RECT 26.970 3.665 27.250 3.895 ;
        RECT 30.080 3.825 30.240 9.030 ;
        RECT 31.195 8.940 31.520 9.030 ;
        RECT 33.575 9.170 33.925 9.290 ;
        RECT 42.080 9.170 42.430 9.245 ;
        RECT 47.520 9.200 47.845 9.265 ;
        RECT 33.575 8.970 42.430 9.170 ;
        RECT 33.575 8.940 33.925 8.970 ;
        RECT 42.080 8.895 42.430 8.970 ;
        RECT 46.405 9.030 47.845 9.200 ;
        RECT 30.395 8.505 30.715 8.830 ;
        RECT 30.425 8.330 30.595 8.505 ;
        RECT 30.425 8.155 30.600 8.330 ;
        RECT 30.425 7.980 31.400 8.155 ;
        RECT 30.395 3.825 30.715 3.945 ;
        RECT 27.580 3.665 27.840 3.755 ;
        RECT 26.680 3.525 27.840 3.665 ;
        RECT 30.080 3.655 30.715 3.825 ;
        RECT 30.395 3.625 30.715 3.655 ;
        RECT 31.225 3.610 31.400 7.980 ;
        RECT 35.925 5.295 39.585 5.435 ;
        RECT 35.135 4.245 35.415 4.620 ;
        RECT 35.925 4.615 36.065 5.295 ;
        RECT 36.345 5.065 36.605 5.155 ;
        RECT 36.345 4.925 38.025 5.065 ;
        RECT 36.345 4.835 36.605 4.925 ;
        RECT 37.885 4.875 38.025 4.925 ;
        RECT 37.885 4.645 38.325 4.875 ;
        RECT 35.925 4.365 36.375 4.615 ;
        RECT 38.065 4.555 38.325 4.645 ;
        RECT 38.845 4.555 39.165 4.875 ;
        RECT 39.445 4.615 39.585 5.295 ;
        RECT 39.755 5.065 40.035 5.180 ;
        RECT 40.835 5.065 43.015 5.175 ;
        RECT 39.755 5.015 43.015 5.065 ;
        RECT 39.755 4.925 40.975 5.015 ;
        RECT 39.755 4.805 40.035 4.925 ;
        RECT 41.675 4.615 41.975 4.620 ;
        RECT 36.095 4.245 36.375 4.365 ;
        RECT 37.385 4.060 37.785 4.225 ;
        RECT 37.385 4.035 37.855 4.060 ;
        RECT 36.105 3.945 36.365 4.035 ;
        RECT 36.105 3.805 37.145 3.945 ;
        RECT 36.105 3.715 36.365 3.805 ;
        RECT 25.880 3.155 26.140 3.475 ;
        RECT 26.680 3.015 26.820 3.525 ;
        RECT 27.580 3.435 27.840 3.525 ;
        RECT 31.170 3.260 31.520 3.610 ;
        RECT 36.575 3.125 36.855 3.500 ;
        RECT 37.005 3.155 37.145 3.805 ;
        RECT 37.325 3.715 37.855 4.035 ;
        RECT 37.575 3.685 37.855 3.715 ;
        RECT 38.295 3.685 38.575 4.060 ;
        RECT 38.845 3.755 38.985 4.555 ;
        RECT 39.445 4.505 41.975 4.615 ;
        RECT 42.465 4.555 42.725 4.875 ;
        RECT 42.465 4.505 42.665 4.555 ;
        RECT 39.445 4.475 42.665 4.505 ;
        RECT 41.695 4.365 42.665 4.475 ;
        RECT 39.145 4.225 39.405 4.315 ;
        RECT 41.695 4.245 41.975 4.365 ;
        RECT 39.145 4.060 39.465 4.225 ;
        RECT 39.145 3.995 39.535 4.060 ;
        RECT 38.785 3.435 39.045 3.755 ;
        RECT 39.255 3.685 39.535 3.995 ;
        RECT 40.135 3.685 40.415 4.060 ;
        RECT 40.745 3.715 41.005 4.035 ;
        RECT 39.765 3.155 40.025 3.475 ;
        RECT 28.865 3.105 29.035 3.110 ;
        RECT 24.480 2.875 26.820 3.015 ;
        RECT 28.775 2.755 29.115 3.105 ;
        RECT 28.775 2.735 29.035 2.755 ;
        RECT 20.290 2.565 29.035 2.735 ;
        RECT 36.615 2.735 36.785 3.125 ;
        RECT 37.005 3.015 39.965 3.155 ;
        RECT 40.805 3.015 40.945 3.715 ;
        RECT 41.815 3.685 42.095 4.055 ;
        RECT 41.885 3.015 42.025 3.685 ;
        RECT 42.265 3.475 42.405 4.365 ;
        RECT 42.865 4.035 43.015 5.015 ;
        RECT 42.585 3.895 43.015 4.035 ;
        RECT 42.585 3.715 42.845 3.895 ;
        RECT 43.295 3.665 43.575 3.895 ;
        RECT 46.405 3.825 46.565 9.030 ;
        RECT 47.520 8.940 47.845 9.030 ;
        RECT 49.900 9.175 50.250 9.295 ;
        RECT 58.405 9.175 58.755 9.250 ;
        RECT 63.845 9.200 64.170 9.265 ;
        RECT 49.900 8.975 58.755 9.175 ;
        RECT 49.900 8.945 50.250 8.975 ;
        RECT 58.405 8.900 58.755 8.975 ;
        RECT 62.730 9.030 64.170 9.200 ;
        RECT 46.720 8.505 47.040 8.830 ;
        RECT 46.750 8.330 46.920 8.505 ;
        RECT 46.750 8.155 46.925 8.330 ;
        RECT 46.750 7.980 47.725 8.155 ;
        RECT 46.720 3.825 47.040 3.945 ;
        RECT 43.905 3.665 44.165 3.755 ;
        RECT 43.005 3.525 44.165 3.665 ;
        RECT 46.405 3.655 47.040 3.825 ;
        RECT 46.720 3.625 47.040 3.655 ;
        RECT 47.550 3.610 47.725 7.980 ;
        RECT 52.250 5.295 55.910 5.435 ;
        RECT 51.460 4.245 51.740 4.620 ;
        RECT 52.250 4.615 52.390 5.295 ;
        RECT 52.670 5.065 52.930 5.155 ;
        RECT 52.670 4.925 54.350 5.065 ;
        RECT 52.670 4.835 52.930 4.925 ;
        RECT 54.210 4.875 54.350 4.925 ;
        RECT 54.210 4.645 54.650 4.875 ;
        RECT 52.250 4.365 52.700 4.615 ;
        RECT 54.390 4.555 54.650 4.645 ;
        RECT 55.170 4.555 55.490 4.875 ;
        RECT 55.770 4.615 55.910 5.295 ;
        RECT 56.080 5.065 56.360 5.180 ;
        RECT 57.160 5.065 59.340 5.175 ;
        RECT 56.080 5.015 59.340 5.065 ;
        RECT 56.080 4.925 57.300 5.015 ;
        RECT 56.080 4.805 56.360 4.925 ;
        RECT 58.000 4.615 58.300 4.620 ;
        RECT 52.420 4.245 52.700 4.365 ;
        RECT 53.710 4.060 54.110 4.225 ;
        RECT 53.710 4.035 54.180 4.060 ;
        RECT 52.430 3.945 52.690 4.035 ;
        RECT 52.430 3.805 53.470 3.945 ;
        RECT 52.430 3.715 52.690 3.805 ;
        RECT 42.205 3.155 42.465 3.475 ;
        RECT 43.005 3.015 43.145 3.525 ;
        RECT 43.905 3.435 44.165 3.525 ;
        RECT 47.495 3.260 47.845 3.610 ;
        RECT 52.900 3.125 53.180 3.500 ;
        RECT 53.330 3.155 53.470 3.805 ;
        RECT 53.650 3.715 54.180 4.035 ;
        RECT 53.900 3.685 54.180 3.715 ;
        RECT 54.620 3.685 54.900 4.060 ;
        RECT 55.170 3.755 55.310 4.555 ;
        RECT 55.770 4.505 58.300 4.615 ;
        RECT 58.790 4.555 59.050 4.875 ;
        RECT 58.790 4.505 58.990 4.555 ;
        RECT 55.770 4.475 58.990 4.505 ;
        RECT 58.020 4.365 58.990 4.475 ;
        RECT 55.470 4.225 55.730 4.315 ;
        RECT 58.020 4.245 58.300 4.365 ;
        RECT 55.470 4.060 55.790 4.225 ;
        RECT 55.470 3.995 55.860 4.060 ;
        RECT 55.110 3.435 55.370 3.755 ;
        RECT 55.580 3.685 55.860 3.995 ;
        RECT 56.460 3.685 56.740 4.060 ;
        RECT 57.070 3.715 57.330 4.035 ;
        RECT 56.090 3.155 56.350 3.475 ;
        RECT 45.190 3.105 45.360 3.110 ;
        RECT 40.805 2.875 43.145 3.015 ;
        RECT 45.100 2.755 45.440 3.105 ;
        RECT 45.100 2.735 45.360 2.755 ;
        RECT 36.615 2.565 45.360 2.735 ;
        RECT 52.940 2.735 53.110 3.125 ;
        RECT 53.330 3.015 56.290 3.155 ;
        RECT 57.130 3.015 57.270 3.715 ;
        RECT 58.140 3.685 58.420 4.055 ;
        RECT 58.210 3.015 58.350 3.685 ;
        RECT 58.590 3.475 58.730 4.365 ;
        RECT 59.190 4.035 59.340 5.015 ;
        RECT 58.910 3.895 59.340 4.035 ;
        RECT 58.910 3.715 59.170 3.895 ;
        RECT 59.620 3.665 59.900 3.895 ;
        RECT 62.730 3.825 62.890 9.030 ;
        RECT 63.845 8.940 64.170 9.030 ;
        RECT 66.180 9.170 66.530 9.290 ;
        RECT 74.730 9.170 75.080 9.245 ;
        RECT 80.170 9.200 80.495 9.265 ;
        RECT 66.180 8.970 75.080 9.170 ;
        RECT 66.180 8.940 66.530 8.970 ;
        RECT 74.730 8.895 75.080 8.970 ;
        RECT 79.055 9.030 80.495 9.200 ;
        RECT 63.045 8.505 63.365 8.830 ;
        RECT 63.075 8.330 63.245 8.505 ;
        RECT 63.075 8.155 63.250 8.330 ;
        RECT 63.075 7.980 64.050 8.155 ;
        RECT 63.045 3.825 63.365 3.945 ;
        RECT 60.230 3.665 60.490 3.755 ;
        RECT 59.330 3.525 60.490 3.665 ;
        RECT 62.730 3.655 63.365 3.825 ;
        RECT 63.045 3.625 63.365 3.655 ;
        RECT 63.875 3.610 64.050 7.980 ;
        RECT 68.575 5.295 72.235 5.435 ;
        RECT 67.785 4.245 68.065 4.620 ;
        RECT 68.575 4.615 68.715 5.295 ;
        RECT 68.995 5.065 69.255 5.155 ;
        RECT 68.995 4.925 70.675 5.065 ;
        RECT 68.995 4.835 69.255 4.925 ;
        RECT 70.535 4.875 70.675 4.925 ;
        RECT 70.535 4.645 70.975 4.875 ;
        RECT 68.575 4.365 69.025 4.615 ;
        RECT 70.715 4.555 70.975 4.645 ;
        RECT 71.495 4.555 71.815 4.875 ;
        RECT 72.095 4.615 72.235 5.295 ;
        RECT 72.405 5.065 72.685 5.180 ;
        RECT 73.485 5.065 75.665 5.175 ;
        RECT 72.405 5.015 75.665 5.065 ;
        RECT 72.405 4.925 73.625 5.015 ;
        RECT 72.405 4.805 72.685 4.925 ;
        RECT 74.325 4.615 74.625 4.620 ;
        RECT 68.745 4.245 69.025 4.365 ;
        RECT 70.035 4.060 70.435 4.225 ;
        RECT 70.035 4.035 70.505 4.060 ;
        RECT 68.755 3.945 69.015 4.035 ;
        RECT 68.755 3.805 69.795 3.945 ;
        RECT 68.755 3.715 69.015 3.805 ;
        RECT 58.530 3.155 58.790 3.475 ;
        RECT 59.330 3.015 59.470 3.525 ;
        RECT 60.230 3.435 60.490 3.525 ;
        RECT 63.820 3.260 64.170 3.610 ;
        RECT 69.225 3.125 69.505 3.500 ;
        RECT 69.655 3.155 69.795 3.805 ;
        RECT 69.975 3.715 70.505 4.035 ;
        RECT 70.225 3.685 70.505 3.715 ;
        RECT 70.945 3.685 71.225 4.060 ;
        RECT 71.495 3.755 71.635 4.555 ;
        RECT 72.095 4.505 74.625 4.615 ;
        RECT 75.115 4.555 75.375 4.875 ;
        RECT 75.115 4.505 75.315 4.555 ;
        RECT 72.095 4.475 75.315 4.505 ;
        RECT 74.345 4.365 75.315 4.475 ;
        RECT 71.795 4.225 72.055 4.315 ;
        RECT 74.345 4.245 74.625 4.365 ;
        RECT 71.795 4.060 72.115 4.225 ;
        RECT 71.795 3.995 72.185 4.060 ;
        RECT 71.435 3.435 71.695 3.755 ;
        RECT 71.905 3.685 72.185 3.995 ;
        RECT 72.785 3.685 73.065 4.060 ;
        RECT 73.395 3.715 73.655 4.035 ;
        RECT 72.415 3.155 72.675 3.475 ;
        RECT 61.515 3.105 61.685 3.110 ;
        RECT 57.130 2.875 59.470 3.015 ;
        RECT 61.425 2.755 61.765 3.105 ;
        RECT 61.425 2.735 61.685 2.755 ;
        RECT 52.940 2.565 61.685 2.735 ;
        RECT 69.265 2.735 69.435 3.125 ;
        RECT 69.655 3.015 72.615 3.155 ;
        RECT 73.455 3.015 73.595 3.715 ;
        RECT 74.465 3.685 74.745 4.055 ;
        RECT 74.535 3.015 74.675 3.685 ;
        RECT 74.915 3.475 75.055 4.365 ;
        RECT 75.515 4.035 75.665 5.015 ;
        RECT 75.235 3.895 75.665 4.035 ;
        RECT 75.235 3.715 75.495 3.895 ;
        RECT 75.945 3.665 76.225 3.895 ;
        RECT 79.055 3.825 79.215 9.030 ;
        RECT 80.170 8.940 80.495 9.030 ;
        RECT 82.505 9.170 82.855 9.290 ;
        RECT 91.060 9.170 91.410 9.245 ;
        RECT 96.495 9.200 96.820 9.265 ;
        RECT 82.505 8.970 91.410 9.170 ;
        RECT 82.505 8.940 82.855 8.970 ;
        RECT 91.060 8.895 91.410 8.970 ;
        RECT 95.380 9.030 96.820 9.200 ;
        RECT 79.370 8.505 79.690 8.830 ;
        RECT 79.400 8.330 79.570 8.505 ;
        RECT 79.400 8.155 79.575 8.330 ;
        RECT 79.400 7.980 80.375 8.155 ;
        RECT 79.370 3.825 79.690 3.945 ;
        RECT 76.555 3.665 76.815 3.755 ;
        RECT 75.655 3.525 76.815 3.665 ;
        RECT 79.055 3.655 79.690 3.825 ;
        RECT 79.370 3.625 79.690 3.655 ;
        RECT 80.200 3.610 80.375 7.980 ;
        RECT 84.900 5.295 88.560 5.435 ;
        RECT 84.110 4.245 84.390 4.620 ;
        RECT 84.900 4.615 85.040 5.295 ;
        RECT 85.320 5.065 85.580 5.155 ;
        RECT 85.320 4.925 87.000 5.065 ;
        RECT 85.320 4.835 85.580 4.925 ;
        RECT 86.860 4.875 87.000 4.925 ;
        RECT 86.860 4.645 87.300 4.875 ;
        RECT 84.900 4.365 85.350 4.615 ;
        RECT 87.040 4.555 87.300 4.645 ;
        RECT 87.820 4.555 88.140 4.875 ;
        RECT 88.420 4.615 88.560 5.295 ;
        RECT 88.730 5.065 89.010 5.180 ;
        RECT 89.810 5.065 91.990 5.175 ;
        RECT 88.730 5.015 91.990 5.065 ;
        RECT 88.730 4.925 89.950 5.015 ;
        RECT 88.730 4.805 89.010 4.925 ;
        RECT 90.650 4.615 90.950 4.620 ;
        RECT 85.070 4.245 85.350 4.365 ;
        RECT 86.360 4.060 86.760 4.225 ;
        RECT 86.360 4.035 86.830 4.060 ;
        RECT 85.080 3.945 85.340 4.035 ;
        RECT 85.080 3.805 86.120 3.945 ;
        RECT 85.080 3.715 85.340 3.805 ;
        RECT 74.855 3.155 75.115 3.475 ;
        RECT 75.655 3.015 75.795 3.525 ;
        RECT 76.555 3.435 76.815 3.525 ;
        RECT 80.145 3.260 80.495 3.610 ;
        RECT 85.550 3.125 85.830 3.500 ;
        RECT 85.980 3.155 86.120 3.805 ;
        RECT 86.300 3.715 86.830 4.035 ;
        RECT 86.550 3.685 86.830 3.715 ;
        RECT 87.270 3.685 87.550 4.060 ;
        RECT 87.820 3.755 87.960 4.555 ;
        RECT 88.420 4.505 90.950 4.615 ;
        RECT 91.440 4.555 91.700 4.875 ;
        RECT 91.440 4.505 91.640 4.555 ;
        RECT 88.420 4.475 91.640 4.505 ;
        RECT 90.670 4.365 91.640 4.475 ;
        RECT 88.120 4.225 88.380 4.315 ;
        RECT 90.670 4.245 90.950 4.365 ;
        RECT 88.120 4.060 88.440 4.225 ;
        RECT 88.120 3.995 88.510 4.060 ;
        RECT 87.760 3.435 88.020 3.755 ;
        RECT 88.230 3.685 88.510 3.995 ;
        RECT 89.110 3.685 89.390 4.060 ;
        RECT 89.720 3.715 89.980 4.035 ;
        RECT 88.740 3.155 89.000 3.475 ;
        RECT 77.840 3.105 78.010 3.110 ;
        RECT 73.455 2.875 75.795 3.015 ;
        RECT 77.750 2.755 78.090 3.105 ;
        RECT 77.750 2.735 78.010 2.755 ;
        RECT 69.265 2.565 78.010 2.735 ;
        RECT 85.590 2.735 85.760 3.125 ;
        RECT 85.980 3.015 88.940 3.155 ;
        RECT 89.780 3.015 89.920 3.715 ;
        RECT 90.790 3.685 91.070 4.055 ;
        RECT 90.860 3.015 91.000 3.685 ;
        RECT 91.240 3.475 91.380 4.365 ;
        RECT 91.840 4.035 91.990 5.015 ;
        RECT 91.560 3.895 91.990 4.035 ;
        RECT 91.560 3.715 91.820 3.895 ;
        RECT 92.270 3.665 92.550 3.895 ;
        RECT 95.380 3.825 95.540 9.030 ;
        RECT 96.495 8.940 96.820 9.030 ;
        RECT 95.695 8.505 96.015 8.830 ;
        RECT 95.725 8.330 95.895 8.505 ;
        RECT 95.725 8.155 95.900 8.330 ;
        RECT 95.725 7.980 96.700 8.155 ;
        RECT 95.695 3.825 96.015 3.945 ;
        RECT 92.880 3.665 93.140 3.755 ;
        RECT 91.980 3.525 93.140 3.665 ;
        RECT 95.380 3.655 96.015 3.825 ;
        RECT 95.695 3.625 96.015 3.655 ;
        RECT 96.525 3.610 96.700 7.980 ;
        RECT 91.180 3.155 91.440 3.475 ;
        RECT 91.980 3.015 92.120 3.525 ;
        RECT 92.880 3.435 93.140 3.525 ;
        RECT 96.470 3.260 96.820 3.610 ;
        RECT 94.165 3.105 94.335 3.110 ;
        RECT 89.780 2.875 92.120 3.015 ;
        RECT 94.075 2.755 94.415 3.105 ;
        RECT 94.075 2.735 94.335 2.755 ;
        RECT 85.590 2.565 94.335 2.735 ;
      LAYER met3 ;
        RECT 25.105 9.675 25.475 9.710 ;
        RECT 41.430 9.675 41.800 9.710 ;
        RECT 57.755 9.675 58.125 9.710 ;
        RECT 74.080 9.675 74.450 9.710 ;
        RECT 90.405 9.675 90.775 9.710 ;
        RECT 25.105 9.375 27.090 9.675 ;
        RECT 25.105 9.340 25.475 9.375 ;
        RECT 23.405 5.145 23.740 5.165 ;
        RECT 22.200 4.845 23.740 5.145 ;
        RECT 18.785 3.865 19.120 4.600 ;
        RECT 21.230 4.040 21.560 4.435 ;
        RECT 22.200 4.040 22.500 4.845 ;
        RECT 23.405 4.825 23.740 4.845 ;
        RECT 25.345 4.275 25.680 4.600 ;
        RECT 20.230 3.470 20.560 3.875 ;
        RECT 21.225 3.705 21.560 4.040 ;
        RECT 21.945 3.725 22.500 4.040 ;
        RECT 22.905 3.875 23.240 4.040 ;
        RECT 23.785 3.875 24.120 4.040 ;
        RECT 21.945 3.705 22.280 3.725 ;
        RECT 22.905 3.710 25.050 3.875 ;
        RECT 25.350 3.865 25.680 4.275 ;
        RECT 26.790 3.875 27.090 9.375 ;
        RECT 41.430 9.375 43.415 9.675 ;
        RECT 41.430 9.340 41.800 9.375 ;
        RECT 39.730 5.145 40.065 5.165 ;
        RECT 38.525 4.845 40.065 5.145 ;
        RECT 20.225 3.145 20.560 3.470 ;
        RECT 22.910 3.575 25.050 3.710 ;
        RECT 22.910 3.305 23.240 3.575 ;
        RECT 23.790 3.305 24.120 3.575 ;
        RECT 24.750 3.565 25.050 3.575 ;
        RECT 25.990 3.575 27.280 3.875 ;
        RECT 35.110 3.865 35.445 4.600 ;
        RECT 37.555 4.040 37.885 4.435 ;
        RECT 38.525 4.040 38.825 4.845 ;
        RECT 39.730 4.825 40.065 4.845 ;
        RECT 41.670 4.275 42.005 4.600 ;
        RECT 25.990 3.565 26.295 3.575 ;
        RECT 24.750 3.275 26.295 3.565 ;
        RECT 26.945 3.525 27.280 3.575 ;
        RECT 24.750 3.260 26.110 3.275 ;
        RECT 26.950 3.145 27.280 3.525 ;
        RECT 36.555 3.470 36.885 3.875 ;
        RECT 37.550 3.705 37.885 4.040 ;
        RECT 38.270 3.725 38.825 4.040 ;
        RECT 39.230 3.875 39.565 4.040 ;
        RECT 40.110 3.875 40.445 4.040 ;
        RECT 38.270 3.705 38.605 3.725 ;
        RECT 39.230 3.710 41.375 3.875 ;
        RECT 41.675 3.865 42.005 4.275 ;
        RECT 43.115 3.875 43.415 9.375 ;
        RECT 57.755 9.375 59.740 9.675 ;
        RECT 57.755 9.340 58.125 9.375 ;
        RECT 56.055 5.145 56.390 5.165 ;
        RECT 54.850 4.845 56.390 5.145 ;
        RECT 36.550 3.145 36.885 3.470 ;
        RECT 39.235 3.575 41.375 3.710 ;
        RECT 39.235 3.305 39.565 3.575 ;
        RECT 40.115 3.305 40.445 3.575 ;
        RECT 41.075 3.565 41.375 3.575 ;
        RECT 42.315 3.575 43.605 3.875 ;
        RECT 51.435 3.865 51.770 4.600 ;
        RECT 53.880 4.040 54.210 4.435 ;
        RECT 54.850 4.040 55.150 4.845 ;
        RECT 56.055 4.825 56.390 4.845 ;
        RECT 57.995 4.275 58.330 4.600 ;
        RECT 42.315 3.565 42.620 3.575 ;
        RECT 41.075 3.275 42.620 3.565 ;
        RECT 43.270 3.525 43.605 3.575 ;
        RECT 41.075 3.260 42.435 3.275 ;
        RECT 43.275 3.145 43.605 3.525 ;
        RECT 52.880 3.470 53.210 3.875 ;
        RECT 53.875 3.705 54.210 4.040 ;
        RECT 54.595 3.725 55.150 4.040 ;
        RECT 55.555 3.875 55.890 4.040 ;
        RECT 56.435 3.875 56.770 4.040 ;
        RECT 54.595 3.705 54.930 3.725 ;
        RECT 55.555 3.710 57.700 3.875 ;
        RECT 58.000 3.865 58.330 4.275 ;
        RECT 59.440 3.875 59.740 9.375 ;
        RECT 74.080 9.375 76.065 9.675 ;
        RECT 74.080 9.340 74.450 9.375 ;
        RECT 72.380 5.145 72.715 5.165 ;
        RECT 71.175 4.845 72.715 5.145 ;
        RECT 52.875 3.145 53.210 3.470 ;
        RECT 55.560 3.575 57.700 3.710 ;
        RECT 55.560 3.305 55.890 3.575 ;
        RECT 56.440 3.305 56.770 3.575 ;
        RECT 57.400 3.565 57.700 3.575 ;
        RECT 58.640 3.575 59.930 3.875 ;
        RECT 67.760 3.865 68.095 4.600 ;
        RECT 70.205 4.040 70.535 4.435 ;
        RECT 71.175 4.040 71.475 4.845 ;
        RECT 72.380 4.825 72.715 4.845 ;
        RECT 74.320 4.275 74.655 4.600 ;
        RECT 58.640 3.565 58.945 3.575 ;
        RECT 57.400 3.275 58.945 3.565 ;
        RECT 59.595 3.525 59.930 3.575 ;
        RECT 57.400 3.260 58.760 3.275 ;
        RECT 59.600 3.145 59.930 3.525 ;
        RECT 69.205 3.470 69.535 3.875 ;
        RECT 70.200 3.705 70.535 4.040 ;
        RECT 70.920 3.725 71.475 4.040 ;
        RECT 71.880 3.875 72.215 4.040 ;
        RECT 72.760 3.875 73.095 4.040 ;
        RECT 70.920 3.705 71.255 3.725 ;
        RECT 71.880 3.710 74.025 3.875 ;
        RECT 74.325 3.865 74.655 4.275 ;
        RECT 75.765 3.875 76.065 9.375 ;
        RECT 90.405 9.375 92.390 9.675 ;
        RECT 90.405 9.340 90.775 9.375 ;
        RECT 88.705 5.145 89.040 5.165 ;
        RECT 87.500 4.845 89.040 5.145 ;
        RECT 69.200 3.145 69.535 3.470 ;
        RECT 71.885 3.575 74.025 3.710 ;
        RECT 71.885 3.305 72.215 3.575 ;
        RECT 72.765 3.305 73.095 3.575 ;
        RECT 73.725 3.565 74.025 3.575 ;
        RECT 74.965 3.575 76.255 3.875 ;
        RECT 84.085 3.865 84.420 4.600 ;
        RECT 86.530 4.040 86.860 4.435 ;
        RECT 87.500 4.040 87.800 4.845 ;
        RECT 88.705 4.825 89.040 4.845 ;
        RECT 90.645 4.275 90.980 4.600 ;
        RECT 74.965 3.565 75.270 3.575 ;
        RECT 73.725 3.275 75.270 3.565 ;
        RECT 75.920 3.525 76.255 3.575 ;
        RECT 73.725 3.260 75.085 3.275 ;
        RECT 75.925 3.145 76.255 3.525 ;
        RECT 85.530 3.470 85.860 3.875 ;
        RECT 86.525 3.705 86.860 4.040 ;
        RECT 87.245 3.725 87.800 4.040 ;
        RECT 88.205 3.875 88.540 4.040 ;
        RECT 89.085 3.875 89.420 4.040 ;
        RECT 87.245 3.705 87.580 3.725 ;
        RECT 88.205 3.710 90.350 3.875 ;
        RECT 90.650 3.865 90.980 4.275 ;
        RECT 92.090 3.875 92.390 9.375 ;
        RECT 85.525 3.145 85.860 3.470 ;
        RECT 88.210 3.575 90.350 3.710 ;
        RECT 88.210 3.305 88.540 3.575 ;
        RECT 89.090 3.305 89.420 3.575 ;
        RECT 90.050 3.565 90.350 3.575 ;
        RECT 91.290 3.575 92.580 3.875 ;
        RECT 91.290 3.565 91.595 3.575 ;
        RECT 90.050 3.275 91.595 3.565 ;
        RECT 92.245 3.525 92.580 3.575 ;
        RECT 90.050 3.260 91.410 3.275 ;
        RECT 92.250 3.145 92.580 3.525 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r1
MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r1
  CLASS BLOCK ;
  FOREIGN sky130_osu_ring_oscillator_mpr2et_8_b0r1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.615 BY 12.465 ;
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 26.045 8.240 26.215 9.510 ;
        RECT 31.660 8.240 31.830 9.510 ;
        RECT 31.660 2.955 31.830 4.225 ;
      LAYER met1 ;
        RECT 25.960 8.410 26.310 8.500 ;
        RECT 31.580 8.410 31.920 8.485 ;
        RECT 25.960 8.380 26.445 8.410 ;
        RECT 31.580 8.405 32.060 8.410 ;
        RECT 31.565 8.380 32.065 8.405 ;
        RECT 25.960 8.235 32.065 8.380 ;
        RECT 25.960 8.200 31.920 8.235 ;
        RECT 25.960 8.150 26.310 8.200 ;
        RECT 31.580 8.135 31.920 8.200 ;
        RECT 31.590 4.225 31.930 4.350 ;
        RECT 31.590 4.055 32.060 4.225 ;
        RECT 31.590 4.000 31.930 4.055 ;
      LAYER met2 ;
        RECT 25.945 8.135 26.325 8.515 ;
        RECT 31.580 8.135 31.920 8.485 ;
        RECT 31.665 4.350 31.835 8.135 ;
        RECT 31.590 4.000 31.930 4.350 ;
      LAYER met3 ;
        RECT 25.970 8.515 26.295 12.360 ;
        RECT 25.945 8.135 26.325 8.515 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 44.605 8.240 44.775 9.510 ;
        RECT 50.220 8.240 50.390 9.510 ;
        RECT 50.220 2.955 50.390 4.225 ;
      LAYER met1 ;
        RECT 44.520 8.410 44.870 8.500 ;
        RECT 50.140 8.410 50.480 8.485 ;
        RECT 44.520 8.380 45.005 8.410 ;
        RECT 50.140 8.405 50.620 8.410 ;
        RECT 50.125 8.380 50.625 8.405 ;
        RECT 44.520 8.235 50.625 8.380 ;
        RECT 44.520 8.200 50.480 8.235 ;
        RECT 44.520 8.150 44.870 8.200 ;
        RECT 50.140 8.135 50.480 8.200 ;
        RECT 50.150 4.225 50.490 4.350 ;
        RECT 50.150 4.055 50.620 4.225 ;
        RECT 50.150 4.000 50.490 4.055 ;
      LAYER met2 ;
        RECT 44.505 8.135 44.885 8.515 ;
        RECT 50.140 8.135 50.480 8.485 ;
        RECT 50.225 4.350 50.395 8.135 ;
        RECT 50.150 4.000 50.490 4.350 ;
      LAYER met3 ;
        RECT 44.530 8.515 44.855 12.360 ;
        RECT 44.505 8.135 44.885 8.515 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 63.165 8.240 63.335 9.510 ;
        RECT 68.780 8.240 68.950 9.510 ;
        RECT 68.780 2.955 68.950 4.225 ;
      LAYER met1 ;
        RECT 63.080 8.410 63.430 8.500 ;
        RECT 68.700 8.410 69.040 8.485 ;
        RECT 63.080 8.380 63.565 8.410 ;
        RECT 68.700 8.405 69.180 8.410 ;
        RECT 68.685 8.380 69.185 8.405 ;
        RECT 63.080 8.235 69.185 8.380 ;
        RECT 63.080 8.200 69.040 8.235 ;
        RECT 63.080 8.150 63.430 8.200 ;
        RECT 68.700 8.135 69.040 8.200 ;
        RECT 68.710 4.225 69.050 4.350 ;
        RECT 68.710 4.055 69.180 4.225 ;
        RECT 68.710 4.000 69.050 4.055 ;
      LAYER met2 ;
        RECT 63.065 8.135 63.445 8.515 ;
        RECT 68.700 8.135 69.040 8.485 ;
        RECT 68.785 4.350 68.955 8.135 ;
        RECT 68.710 4.000 69.050 4.350 ;
      LAYER met3 ;
        RECT 63.090 8.515 63.415 12.360 ;
        RECT 63.065 8.135 63.445 8.515 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 81.725 8.240 81.895 9.510 ;
        RECT 87.340 8.240 87.510 9.510 ;
        RECT 87.340 2.955 87.510 4.225 ;
      LAYER met1 ;
        RECT 81.640 8.410 81.990 8.500 ;
        RECT 87.260 8.410 87.600 8.485 ;
        RECT 81.640 8.380 82.125 8.410 ;
        RECT 87.260 8.405 87.740 8.410 ;
        RECT 87.245 8.380 87.745 8.405 ;
        RECT 81.640 8.235 87.745 8.380 ;
        RECT 81.640 8.200 87.600 8.235 ;
        RECT 81.640 8.150 81.990 8.200 ;
        RECT 87.260 8.135 87.600 8.200 ;
        RECT 87.270 4.225 87.610 4.350 ;
        RECT 87.270 4.055 87.740 4.225 ;
        RECT 87.270 4.000 87.610 4.055 ;
      LAYER met2 ;
        RECT 81.625 8.135 82.005 8.515 ;
        RECT 87.260 8.135 87.600 8.485 ;
        RECT 87.345 4.350 87.515 8.135 ;
        RECT 87.270 4.000 87.610 4.350 ;
      LAYER met3 ;
        RECT 81.650 8.515 81.975 12.360 ;
        RECT 81.625 8.135 82.005 8.515 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 100.285 8.240 100.455 9.510 ;
        RECT 105.900 8.240 106.070 9.510 ;
        RECT 105.900 2.955 106.070 4.225 ;
      LAYER met1 ;
        RECT 100.200 8.410 100.550 8.500 ;
        RECT 105.820 8.410 106.160 8.485 ;
        RECT 100.200 8.380 100.685 8.410 ;
        RECT 105.820 8.405 106.300 8.410 ;
        RECT 105.805 8.380 106.305 8.405 ;
        RECT 100.200 8.235 106.305 8.380 ;
        RECT 100.200 8.200 106.160 8.235 ;
        RECT 100.200 8.150 100.550 8.200 ;
        RECT 105.820 8.135 106.160 8.200 ;
        RECT 105.830 4.225 106.170 4.350 ;
        RECT 105.830 4.055 106.300 4.225 ;
        RECT 105.830 4.000 106.170 4.055 ;
      LAYER met2 ;
        RECT 100.185 8.135 100.565 8.515 ;
        RECT 105.820 8.135 106.160 8.485 ;
        RECT 105.905 4.350 106.075 8.135 ;
        RECT 105.830 4.000 106.170 4.350 ;
      LAYER met3 ;
        RECT 100.210 8.515 100.535 12.360 ;
        RECT 100.185 8.135 100.565 8.515 ;
    END
  END s5
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 35.810 4.015 35.985 5.160 ;
        RECT 35.810 3.580 35.980 4.015 ;
        RECT 35.815 1.870 35.985 2.380 ;
      LAYER met1 ;
        RECT 35.750 3.545 36.040 3.780 ;
        RECT 35.750 3.540 35.980 3.545 ;
        RECT 35.810 2.440 35.980 3.540 ;
        RECT 35.750 2.180 36.045 2.440 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 54.370 4.015 54.545 5.160 ;
        RECT 54.370 3.580 54.540 4.015 ;
        RECT 54.375 1.870 54.545 2.380 ;
      LAYER met1 ;
        RECT 54.310 3.545 54.600 3.780 ;
        RECT 54.310 3.540 54.540 3.545 ;
        RECT 54.370 2.440 54.540 3.540 ;
        RECT 54.310 2.180 54.605 2.440 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 72.930 4.015 73.105 5.160 ;
        RECT 72.930 3.580 73.100 4.015 ;
        RECT 72.935 1.870 73.105 2.380 ;
      LAYER met1 ;
        RECT 72.870 3.545 73.160 3.780 ;
        RECT 72.870 3.540 73.100 3.545 ;
        RECT 72.930 2.440 73.100 3.540 ;
        RECT 72.870 2.180 73.165 2.440 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 91.490 4.015 91.665 5.160 ;
        RECT 91.490 3.580 91.660 4.015 ;
        RECT 91.495 1.870 91.665 2.380 ;
      LAYER met1 ;
        RECT 91.430 3.545 91.720 3.780 ;
        RECT 91.430 3.540 91.660 3.545 ;
        RECT 91.490 2.440 91.660 3.540 ;
        RECT 91.430 2.180 91.725 2.440 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 110.050 4.015 110.225 5.160 ;
        RECT 110.050 3.580 110.220 4.015 ;
        RECT 110.055 1.870 110.225 2.380 ;
      LAYER met1 ;
        RECT 109.990 3.545 110.280 3.780 ;
        RECT 109.990 3.540 110.220 3.545 ;
        RECT 110.050 2.440 110.220 3.540 ;
        RECT 109.990 2.180 110.285 2.440 ;
    END
  END X5_Y1
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 15.230 8.240 15.400 9.510 ;
      LAYER met1 ;
        RECT 15.170 8.435 15.460 8.440 ;
        RECT 15.170 8.410 15.465 8.435 ;
        RECT 15.170 8.240 15.630 8.410 ;
        RECT 15.170 8.210 15.465 8.240 ;
        RECT 15.175 8.205 15.465 8.210 ;
    END
  END start
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.005 10.865 110.605 12.465 ;
        RECT 15.220 10.240 15.390 10.865 ;
        RECT 26.035 10.240 26.205 10.865 ;
        RECT 26.990 10.320 27.160 10.600 ;
        RECT 26.990 10.150 27.220 10.320 ;
        RECT 31.650 10.240 31.820 10.865 ;
        RECT 34.395 10.235 34.565 10.865 ;
        RECT 35.385 10.235 35.555 10.865 ;
        RECT 44.595 10.240 44.765 10.865 ;
        RECT 45.550 10.320 45.720 10.600 ;
        RECT 45.550 10.150 45.780 10.320 ;
        RECT 50.210 10.240 50.380 10.865 ;
        RECT 52.955 10.235 53.125 10.865 ;
        RECT 53.945 10.235 54.115 10.865 ;
        RECT 63.155 10.240 63.325 10.865 ;
        RECT 64.110 10.320 64.280 10.600 ;
        RECT 64.110 10.150 64.340 10.320 ;
        RECT 68.770 10.240 68.940 10.865 ;
        RECT 71.515 10.235 71.685 10.865 ;
        RECT 72.505 10.235 72.675 10.865 ;
        RECT 81.715 10.240 81.885 10.865 ;
        RECT 82.670 10.320 82.840 10.600 ;
        RECT 82.670 10.150 82.900 10.320 ;
        RECT 87.330 10.240 87.500 10.865 ;
        RECT 90.075 10.235 90.245 10.865 ;
        RECT 91.065 10.235 91.235 10.865 ;
        RECT 100.275 10.240 100.445 10.865 ;
        RECT 101.230 10.320 101.400 10.600 ;
        RECT 101.230 10.150 101.460 10.320 ;
        RECT 105.890 10.240 106.060 10.865 ;
        RECT 108.635 10.235 108.805 10.865 ;
        RECT 109.625 10.235 109.795 10.865 ;
        RECT 27.050 8.540 27.220 10.150 ;
        RECT 45.610 8.540 45.780 10.150 ;
        RECT 64.170 8.540 64.340 10.150 ;
        RECT 82.730 8.540 82.900 10.150 ;
        RECT 101.290 8.540 101.460 10.150 ;
        RECT 26.990 8.370 27.220 8.540 ;
        RECT 45.550 8.370 45.780 8.540 ;
        RECT 64.110 8.370 64.340 8.540 ;
        RECT 82.670 8.370 82.900 8.540 ;
        RECT 101.230 8.370 101.460 8.540 ;
        RECT 26.990 7.310 27.160 8.370 ;
        RECT 45.550 7.310 45.720 8.370 ;
        RECT 64.110 7.310 64.280 8.370 ;
        RECT 82.670 7.310 82.840 8.370 ;
        RECT 101.230 7.310 101.400 8.370 ;
      LAYER met1 ;
        RECT 0.005 10.865 110.605 12.465 ;
        RECT 26.550 8.790 26.720 10.865 ;
        RECT 26.990 8.790 27.280 8.820 ;
        RECT 26.550 8.605 27.280 8.790 ;
        RECT 45.110 8.790 45.280 10.865 ;
        RECT 45.550 8.790 45.840 8.820 ;
        RECT 45.110 8.605 45.840 8.790 ;
        RECT 63.670 8.790 63.840 10.865 ;
        RECT 64.110 8.790 64.400 8.820 ;
        RECT 63.670 8.605 64.400 8.790 ;
        RECT 82.230 8.790 82.400 10.865 ;
        RECT 82.670 8.790 82.960 8.820 ;
        RECT 82.230 8.605 82.960 8.790 ;
        RECT 100.790 8.790 100.960 10.865 ;
        RECT 101.230 8.790 101.520 8.820 ;
        RECT 100.790 8.605 101.520 8.790 ;
        RECT 26.990 8.590 27.280 8.605 ;
        RECT 45.550 8.590 45.840 8.605 ;
        RECT 64.110 8.590 64.400 8.605 ;
        RECT 82.670 8.590 82.960 8.605 ;
        RECT 101.230 8.590 101.520 8.605 ;
    END
    PORT
      LAYER li1 ;
        RECT 20.195 4.345 20.485 4.515 ;
        RECT 38.755 4.345 39.045 4.515 ;
        RECT 57.315 4.345 57.605 4.515 ;
        RECT 75.875 4.345 76.165 4.515 ;
        RECT 94.435 4.345 94.725 4.515 ;
        RECT 20.195 4.035 20.365 4.345 ;
        RECT 19.995 3.865 20.365 4.035 ;
        RECT 22.035 3.785 22.205 4.115 ;
        RECT 38.755 4.035 38.925 4.345 ;
        RECT 38.555 3.865 38.925 4.035 ;
        RECT 40.595 3.785 40.765 4.115 ;
        RECT 57.315 4.035 57.485 4.345 ;
        RECT 57.115 3.865 57.485 4.035 ;
        RECT 59.155 3.785 59.325 4.115 ;
        RECT 75.875 4.035 76.045 4.345 ;
        RECT 75.675 3.865 76.045 4.035 ;
        RECT 77.715 3.785 77.885 4.115 ;
        RECT 94.435 4.035 94.605 4.345 ;
        RECT 94.235 3.865 94.605 4.035 ;
        RECT 96.275 3.785 96.445 4.115 ;
        RECT 19.355 2.875 19.525 3.375 ;
        RECT 20.835 2.875 21.005 3.375 ;
        RECT 22.755 2.875 22.925 3.375 ;
        RECT 24.235 2.875 24.405 3.375 ;
        RECT 25.195 2.875 25.365 3.375 ;
        RECT 26.195 2.875 26.365 3.375 ;
        RECT 27.155 2.875 27.325 3.375 ;
        RECT 27.675 2.875 27.845 3.375 ;
        RECT 28.635 2.875 28.805 3.375 ;
        RECT 29.595 2.875 29.765 3.375 ;
        RECT 37.915 2.875 38.085 3.375 ;
        RECT 39.395 2.875 39.565 3.375 ;
        RECT 41.315 2.875 41.485 3.375 ;
        RECT 42.795 2.875 42.965 3.375 ;
        RECT 43.755 2.875 43.925 3.375 ;
        RECT 44.755 2.875 44.925 3.375 ;
        RECT 45.715 2.875 45.885 3.375 ;
        RECT 46.235 2.875 46.405 3.375 ;
        RECT 47.195 2.875 47.365 3.375 ;
        RECT 48.155 2.875 48.325 3.375 ;
        RECT 56.475 2.875 56.645 3.375 ;
        RECT 57.955 2.875 58.125 3.375 ;
        RECT 59.875 2.875 60.045 3.375 ;
        RECT 61.355 2.875 61.525 3.375 ;
        RECT 62.315 2.875 62.485 3.375 ;
        RECT 63.315 2.875 63.485 3.375 ;
        RECT 64.275 2.875 64.445 3.375 ;
        RECT 64.795 2.875 64.965 3.375 ;
        RECT 65.755 2.875 65.925 3.375 ;
        RECT 66.715 2.875 66.885 3.375 ;
        RECT 75.035 2.875 75.205 3.375 ;
        RECT 76.515 2.875 76.685 3.375 ;
        RECT 78.435 2.875 78.605 3.375 ;
        RECT 79.915 2.875 80.085 3.375 ;
        RECT 80.875 2.875 81.045 3.375 ;
        RECT 81.875 2.875 82.045 3.375 ;
        RECT 82.835 2.875 83.005 3.375 ;
        RECT 83.355 2.875 83.525 3.375 ;
        RECT 84.315 2.875 84.485 3.375 ;
        RECT 85.275 2.875 85.445 3.375 ;
        RECT 93.595 2.875 93.765 3.375 ;
        RECT 95.075 2.875 95.245 3.375 ;
        RECT 96.995 2.875 97.165 3.375 ;
        RECT 98.475 2.875 98.645 3.375 ;
        RECT 99.435 2.875 99.605 3.375 ;
        RECT 100.435 2.875 100.605 3.375 ;
        RECT 101.395 2.875 101.565 3.375 ;
        RECT 101.915 2.875 102.085 3.375 ;
        RECT 102.875 2.875 103.045 3.375 ;
        RECT 103.835 2.875 104.005 3.375 ;
        RECT 18.545 1.600 30.590 2.875 ;
        RECT 31.650 1.600 31.820 2.225 ;
        RECT 34.395 1.600 34.565 2.230 ;
        RECT 35.380 1.600 35.550 2.230 ;
        RECT 37.105 1.600 49.150 2.875 ;
        RECT 50.210 1.600 50.380 2.225 ;
        RECT 52.955 1.600 53.125 2.230 ;
        RECT 53.940 1.600 54.110 2.230 ;
        RECT 55.665 1.600 67.710 2.875 ;
        RECT 68.770 1.600 68.940 2.225 ;
        RECT 71.515 1.600 71.685 2.230 ;
        RECT 72.500 1.600 72.670 2.230 ;
        RECT 74.225 1.600 86.270 2.875 ;
        RECT 87.330 1.600 87.500 2.225 ;
        RECT 90.075 1.600 90.245 2.230 ;
        RECT 91.060 1.600 91.230 2.230 ;
        RECT 92.785 1.600 104.830 2.875 ;
        RECT 105.890 1.600 106.060 2.225 ;
        RECT 108.635 1.600 108.805 2.230 ;
        RECT 109.620 1.600 109.790 2.230 ;
        RECT 0.005 0.000 110.600 1.600 ;
      LAYER met1 ;
        RECT 20.235 4.305 20.555 4.565 ;
        RECT 38.795 4.305 39.115 4.565 ;
        RECT 57.355 4.305 57.675 4.565 ;
        RECT 75.915 4.305 76.235 4.565 ;
        RECT 94.475 4.305 94.795 4.565 ;
        RECT 21.975 3.805 22.265 4.035 ;
        RECT 40.535 3.805 40.825 4.035 ;
        RECT 59.095 3.805 59.385 4.035 ;
        RECT 77.655 3.805 77.945 4.035 ;
        RECT 96.215 3.805 96.505 4.035 ;
        RECT 21.205 3.665 22.265 3.805 ;
        RECT 39.765 3.665 40.825 3.805 ;
        RECT 58.325 3.665 59.385 3.805 ;
        RECT 76.885 3.665 77.945 3.805 ;
        RECT 95.445 3.665 96.505 3.805 ;
        RECT 18.545 1.600 30.590 2.905 ;
        RECT 37.105 1.600 49.150 2.905 ;
        RECT 55.665 1.600 67.710 2.905 ;
        RECT 74.225 1.600 86.270 2.905 ;
        RECT 92.785 1.600 104.830 2.905 ;
        RECT 0.005 0.000 110.605 1.600 ;
      LAYER met2 ;
        RECT 20.265 4.505 20.525 4.595 ;
        RECT 38.825 4.505 39.085 4.595 ;
        RECT 57.385 4.505 57.645 4.595 ;
        RECT 75.945 4.505 76.205 4.595 ;
        RECT 94.505 4.505 94.765 4.595 ;
        RECT 20.205 4.275 20.525 4.505 ;
        RECT 38.765 4.275 39.085 4.505 ;
        RECT 57.325 4.275 57.645 4.505 ;
        RECT 75.885 4.275 76.205 4.505 ;
        RECT 94.445 4.275 94.765 4.505 ;
        RECT 20.205 3.945 20.345 4.275 ;
        RECT 20.515 3.945 20.795 4.060 ;
        RECT 21.985 3.945 22.245 4.035 ;
        RECT 20.205 3.805 22.245 3.945 ;
        RECT 38.765 3.945 38.905 4.275 ;
        RECT 39.075 3.945 39.355 4.060 ;
        RECT 40.545 3.945 40.805 4.035 ;
        RECT 38.765 3.805 40.805 3.945 ;
        RECT 57.325 3.945 57.465 4.275 ;
        RECT 57.635 3.945 57.915 4.060 ;
        RECT 59.105 3.945 59.365 4.035 ;
        RECT 57.325 3.805 59.365 3.945 ;
        RECT 75.885 3.945 76.025 4.275 ;
        RECT 76.195 3.945 76.475 4.060 ;
        RECT 77.665 3.945 77.925 4.035 ;
        RECT 75.885 3.805 77.925 3.945 ;
        RECT 94.445 3.945 94.585 4.275 ;
        RECT 94.755 3.945 95.035 4.060 ;
        RECT 96.225 3.945 96.485 4.035 ;
        RECT 94.445 3.805 96.485 3.945 ;
        RECT 20.515 3.685 20.795 3.805 ;
        RECT 21.985 3.715 22.245 3.805 ;
        RECT 39.075 3.685 39.355 3.805 ;
        RECT 40.545 3.715 40.805 3.805 ;
        RECT 57.635 3.685 57.915 3.805 ;
        RECT 59.105 3.715 59.365 3.805 ;
        RECT 76.195 3.685 76.475 3.805 ;
        RECT 77.665 3.715 77.925 3.805 ;
        RECT 94.755 3.685 95.035 3.805 ;
        RECT 96.225 3.715 96.485 3.805 ;
        RECT 20.615 2.635 20.785 3.685 ;
        RECT 39.175 2.635 39.345 3.685 ;
        RECT 57.735 2.635 57.905 3.685 ;
        RECT 76.295 2.635 76.465 3.685 ;
        RECT 94.855 2.635 95.025 3.685 ;
        RECT 20.590 2.295 20.930 2.635 ;
        RECT 39.150 2.295 39.490 2.635 ;
        RECT 57.710 2.295 58.050 2.635 ;
        RECT 76.270 2.295 76.610 2.635 ;
        RECT 94.830 2.295 95.170 2.635 ;
      LAYER met3 ;
        RECT 20.495 4.035 20.820 4.040 ;
        RECT 39.055 4.035 39.380 4.040 ;
        RECT 57.615 4.035 57.940 4.040 ;
        RECT 76.175 4.035 76.500 4.040 ;
        RECT 94.735 4.035 95.060 4.040 ;
        RECT 20.155 3.705 20.885 4.035 ;
        RECT 38.715 3.705 39.445 4.035 ;
        RECT 57.275 3.705 58.005 4.035 ;
        RECT 75.835 3.705 76.565 4.035 ;
        RECT 94.395 3.705 95.125 4.035 ;
        RECT 20.495 3.700 20.820 3.705 ;
        RECT 39.055 3.700 39.380 3.705 ;
        RECT 57.615 3.700 57.940 3.705 ;
        RECT 76.175 3.700 76.500 3.705 ;
        RECT 94.735 3.700 95.060 3.705 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 15.000 8.745 20.165 8.750 ;
        RECT 25.815 8.745 28.625 8.750 ;
        RECT 31.430 8.745 34.240 8.750 ;
        RECT 36.360 8.745 38.725 8.750 ;
        RECT 44.375 8.745 47.185 8.750 ;
        RECT 49.990 8.745 52.800 8.750 ;
        RECT 54.920 8.745 57.285 8.750 ;
        RECT 62.935 8.745 65.745 8.750 ;
        RECT 68.550 8.745 71.360 8.750 ;
        RECT 73.480 8.745 75.845 8.750 ;
        RECT 81.495 8.745 84.305 8.750 ;
        RECT 87.110 8.745 89.920 8.750 ;
        RECT 92.040 8.745 94.405 8.750 ;
        RECT 100.055 8.745 102.865 8.750 ;
        RECT 105.670 8.745 108.480 8.750 ;
        RECT 15.000 5.450 110.600 8.745 ;
        RECT 15.005 5.095 110.600 5.450 ;
        RECT 17.800 4.100 110.600 5.095 ;
        RECT 18.305 4.095 110.600 4.100 ;
        RECT 30.410 3.720 36.360 4.095 ;
        RECT 48.970 3.720 54.920 4.095 ;
        RECT 67.530 4.090 74.800 4.095 ;
        RECT 67.530 3.720 73.480 4.090 ;
        RECT 86.090 3.720 92.040 4.095 ;
        RECT 104.650 3.720 110.600 4.095 ;
        RECT 31.430 3.715 34.240 3.720 ;
        RECT 49.990 3.715 52.800 3.720 ;
        RECT 68.550 3.715 71.360 3.720 ;
        RECT 87.110 3.715 89.920 3.720 ;
        RECT 105.670 3.715 108.480 3.720 ;
      LAYER li1 ;
        RECT 17.035 10.050 17.210 10.600 ;
        RECT 17.035 8.450 17.205 10.050 ;
        RECT 15.220 7.050 15.390 7.770 ;
        RECT 17.035 7.310 17.210 8.450 ;
        RECT 17.035 7.050 17.205 7.310 ;
        RECT 26.035 7.050 26.205 7.770 ;
        RECT 31.650 7.050 31.820 7.770 ;
        RECT 34.395 7.050 34.565 7.765 ;
        RECT 35.385 7.050 35.555 7.765 ;
        RECT 44.595 7.050 44.765 7.770 ;
        RECT 50.210 7.050 50.380 7.770 ;
        RECT 52.955 7.050 53.125 7.765 ;
        RECT 53.945 7.050 54.115 7.765 ;
        RECT 63.155 7.050 63.325 7.770 ;
        RECT 68.770 7.050 68.940 7.770 ;
        RECT 71.515 7.050 71.685 7.765 ;
        RECT 72.505 7.050 72.675 7.765 ;
        RECT 81.715 7.050 81.885 7.770 ;
        RECT 87.330 7.050 87.500 7.770 ;
        RECT 90.075 7.050 90.245 7.765 ;
        RECT 91.065 7.050 91.235 7.765 ;
        RECT 100.275 7.050 100.445 7.770 ;
        RECT 105.890 7.050 106.060 7.770 ;
        RECT 108.635 7.050 108.805 7.765 ;
        RECT 109.625 7.050 109.795 7.765 ;
        RECT 0.000 5.450 110.600 7.050 ;
        RECT 17.800 5.435 110.600 5.450 ;
        RECT 18.545 5.430 36.360 5.435 ;
        RECT 37.105 5.430 54.920 5.435 ;
        RECT 55.665 5.430 73.480 5.435 ;
        RECT 74.225 5.430 92.040 5.435 ;
        RECT 92.785 5.430 110.600 5.435 ;
        RECT 18.545 5.425 30.505 5.430 ;
        RECT 31.480 5.425 34.565 5.430 ;
        RECT 19.355 4.925 19.525 5.425 ;
        RECT 20.315 4.925 20.485 5.425 ;
        RECT 21.315 4.925 21.485 5.425 ;
        RECT 23.275 4.925 23.445 5.425 ;
        RECT 24.235 4.925 24.405 5.425 ;
        RECT 26.195 4.925 26.365 5.425 ;
        RECT 28.635 4.925 28.805 5.425 ;
        RECT 31.650 4.695 31.820 5.425 ;
        RECT 34.395 4.700 34.565 5.425 ;
        RECT 35.380 4.700 35.550 5.430 ;
        RECT 37.105 5.425 49.065 5.430 ;
        RECT 50.040 5.425 53.125 5.430 ;
        RECT 37.915 4.925 38.085 5.425 ;
        RECT 38.875 4.925 39.045 5.425 ;
        RECT 39.875 4.925 40.045 5.425 ;
        RECT 41.835 4.925 42.005 5.425 ;
        RECT 42.795 4.925 42.965 5.425 ;
        RECT 44.755 4.925 44.925 5.425 ;
        RECT 47.195 4.925 47.365 5.425 ;
        RECT 50.210 4.695 50.380 5.425 ;
        RECT 52.955 4.700 53.125 5.425 ;
        RECT 53.940 4.700 54.110 5.430 ;
        RECT 55.665 5.425 67.625 5.430 ;
        RECT 68.600 5.425 71.685 5.430 ;
        RECT 56.475 4.925 56.645 5.425 ;
        RECT 57.435 4.925 57.605 5.425 ;
        RECT 58.435 4.925 58.605 5.425 ;
        RECT 60.395 4.925 60.565 5.425 ;
        RECT 61.355 4.925 61.525 5.425 ;
        RECT 63.315 4.925 63.485 5.425 ;
        RECT 65.755 4.925 65.925 5.425 ;
        RECT 68.770 4.695 68.940 5.425 ;
        RECT 71.515 4.700 71.685 5.425 ;
        RECT 72.500 4.700 72.670 5.430 ;
        RECT 74.225 5.425 86.185 5.430 ;
        RECT 87.160 5.425 90.245 5.430 ;
        RECT 75.035 4.925 75.205 5.425 ;
        RECT 75.995 4.925 76.165 5.425 ;
        RECT 76.995 4.925 77.165 5.425 ;
        RECT 78.955 4.925 79.125 5.425 ;
        RECT 79.915 4.925 80.085 5.425 ;
        RECT 81.875 4.925 82.045 5.425 ;
        RECT 84.315 4.925 84.485 5.425 ;
        RECT 87.330 4.695 87.500 5.425 ;
        RECT 90.075 4.700 90.245 5.425 ;
        RECT 91.060 4.700 91.230 5.430 ;
        RECT 92.785 5.425 104.745 5.430 ;
        RECT 105.720 5.425 108.805 5.430 ;
        RECT 93.595 4.925 93.765 5.425 ;
        RECT 94.555 4.925 94.725 5.425 ;
        RECT 95.555 4.925 95.725 5.425 ;
        RECT 97.515 4.925 97.685 5.425 ;
        RECT 98.475 4.925 98.645 5.425 ;
        RECT 100.435 4.925 100.605 5.425 ;
        RECT 102.875 4.925 103.045 5.425 ;
        RECT 105.890 4.695 106.060 5.425 ;
        RECT 108.635 4.700 108.805 5.425 ;
        RECT 109.620 4.700 109.790 5.430 ;
      LAYER met1 ;
        RECT 16.975 9.150 17.265 9.180 ;
        RECT 16.805 8.980 17.265 9.150 ;
        RECT 16.975 8.950 17.265 8.980 ;
        RECT 0.000 7.025 110.600 7.050 ;
        RECT 0.000 5.450 110.615 7.025 ;
        RECT 17.815 5.425 110.615 5.450 ;
        RECT 18.545 5.395 30.505 5.425 ;
        RECT 37.105 5.395 49.065 5.425 ;
        RECT 55.665 5.395 67.625 5.425 ;
        RECT 74.225 5.395 86.185 5.425 ;
        RECT 92.785 5.395 104.745 5.425 ;
    END
  END vccd1
  OBS
      LAYER pwell ;
        RECT 18.705 2.735 18.875 2.875 ;
        RECT 18.685 2.715 18.875 2.735 ;
        RECT 18.685 2.705 18.855 2.715 ;
        RECT 20.665 2.705 20.835 2.875 ;
        RECT 23.105 2.705 23.275 2.875 ;
        RECT 25.545 2.705 25.715 2.875 ;
        RECT 27.505 2.705 27.675 2.875 ;
        RECT 37.265 2.735 37.435 2.875 ;
        RECT 37.245 2.715 37.435 2.735 ;
        RECT 37.245 2.705 37.415 2.715 ;
        RECT 39.225 2.705 39.395 2.875 ;
        RECT 41.665 2.705 41.835 2.875 ;
        RECT 44.105 2.705 44.275 2.875 ;
        RECT 46.065 2.705 46.235 2.875 ;
        RECT 55.825 2.735 55.995 2.875 ;
        RECT 55.805 2.715 55.995 2.735 ;
        RECT 55.805 2.705 55.975 2.715 ;
        RECT 57.785 2.705 57.955 2.875 ;
        RECT 60.225 2.705 60.395 2.875 ;
        RECT 62.665 2.705 62.835 2.875 ;
        RECT 64.625 2.705 64.795 2.875 ;
        RECT 74.385 2.735 74.555 2.875 ;
        RECT 74.365 2.715 74.555 2.735 ;
        RECT 74.365 2.705 74.535 2.715 ;
        RECT 76.345 2.705 76.515 2.875 ;
        RECT 78.785 2.705 78.955 2.875 ;
        RECT 81.225 2.705 81.395 2.875 ;
        RECT 83.185 2.705 83.355 2.875 ;
        RECT 92.945 2.735 93.115 2.875 ;
        RECT 92.925 2.715 93.115 2.735 ;
        RECT 92.925 2.705 93.095 2.715 ;
        RECT 94.905 2.705 95.075 2.875 ;
        RECT 97.345 2.705 97.515 2.875 ;
        RECT 99.785 2.705 99.955 2.875 ;
        RECT 101.745 2.705 101.915 2.875 ;
      LAYER li1 ;
        RECT 15.650 10.110 15.825 10.600 ;
        RECT 16.175 10.320 16.345 10.600 ;
        RECT 16.175 10.150 16.405 10.320 ;
        RECT 15.650 9.940 15.820 10.110 ;
        RECT 15.650 9.610 16.060 9.940 ;
        RECT 15.650 9.100 15.820 9.610 ;
        RECT 15.650 8.770 16.060 9.100 ;
        RECT 15.650 8.570 15.820 8.770 ;
        RECT 15.650 7.310 15.825 8.570 ;
        RECT 16.235 8.540 16.405 10.150 ;
        RECT 16.605 10.090 16.780 10.600 ;
        RECT 26.465 10.110 26.640 10.600 ;
        RECT 26.465 9.940 26.635 10.110 ;
        RECT 27.420 10.090 27.595 10.600 ;
        RECT 27.850 10.050 28.025 10.600 ;
        RECT 32.080 10.110 32.255 10.600 ;
        RECT 32.605 10.320 32.775 10.600 ;
        RECT 32.605 10.150 32.835 10.320 ;
        RECT 26.465 9.610 26.875 9.940 ;
        RECT 16.175 8.370 16.405 8.540 ;
        RECT 16.605 8.570 16.775 9.520 ;
        RECT 26.465 9.100 26.635 9.610 ;
        RECT 26.465 8.770 26.875 9.100 ;
        RECT 26.465 8.570 26.635 8.770 ;
        RECT 27.420 8.570 27.590 9.520 ;
        RECT 16.175 7.310 16.345 8.370 ;
        RECT 16.605 7.310 16.780 8.570 ;
        RECT 26.465 7.310 26.640 8.570 ;
        RECT 27.420 7.310 27.595 8.570 ;
        RECT 27.850 8.450 28.020 10.050 ;
        RECT 32.080 9.940 32.250 10.110 ;
        RECT 32.080 9.610 32.490 9.940 ;
        RECT 32.080 9.100 32.250 9.610 ;
        RECT 32.080 8.770 32.490 9.100 ;
        RECT 32.080 8.570 32.250 8.770 ;
        RECT 27.850 7.310 28.025 8.450 ;
        RECT 32.080 7.310 32.255 8.570 ;
        RECT 32.665 8.540 32.835 10.150 ;
        RECT 33.035 10.090 33.210 10.600 ;
        RECT 33.465 10.050 33.640 10.600 ;
        RECT 34.830 10.085 35.000 10.595 ;
        RECT 35.820 10.085 35.990 10.595 ;
        RECT 45.025 10.110 45.200 10.600 ;
        RECT 32.605 8.370 32.835 8.540 ;
        RECT 33.035 8.570 33.205 9.520 ;
        RECT 32.605 7.310 32.775 8.370 ;
        RECT 33.035 7.310 33.210 8.570 ;
        RECT 33.465 8.450 33.635 10.050 ;
        RECT 45.025 9.940 45.195 10.110 ;
        RECT 45.980 10.090 46.155 10.600 ;
        RECT 46.410 10.050 46.585 10.600 ;
        RECT 50.640 10.110 50.815 10.600 ;
        RECT 51.165 10.320 51.335 10.600 ;
        RECT 51.165 10.150 51.395 10.320 ;
        RECT 34.395 9.425 34.625 9.625 ;
        RECT 45.025 9.610 45.435 9.940 ;
        RECT 34.395 9.395 34.925 9.425 ;
        RECT 34.455 9.255 34.925 9.395 ;
        RECT 35.445 9.255 35.915 9.425 ;
        RECT 34.455 8.565 34.625 9.255 ;
        RECT 34.825 8.790 34.995 8.885 ;
        RECT 35.445 8.790 35.615 9.255 ;
        RECT 45.025 9.100 45.195 9.610 ;
        RECT 34.825 8.610 35.615 8.790 ;
        RECT 33.465 7.310 33.640 8.450 ;
        RECT 34.825 7.305 35.000 8.610 ;
        RECT 35.445 8.565 35.615 8.610 ;
        RECT 35.815 8.450 35.985 8.885 ;
        RECT 45.025 8.770 45.435 9.100 ;
        RECT 45.025 8.570 45.195 8.770 ;
        RECT 45.980 8.570 46.150 9.520 ;
        RECT 35.815 7.305 35.990 8.450 ;
        RECT 45.025 7.310 45.200 8.570 ;
        RECT 45.980 7.310 46.155 8.570 ;
        RECT 46.410 8.450 46.580 10.050 ;
        RECT 50.640 9.940 50.810 10.110 ;
        RECT 50.640 9.610 51.050 9.940 ;
        RECT 50.640 9.100 50.810 9.610 ;
        RECT 50.640 8.770 51.050 9.100 ;
        RECT 50.640 8.570 50.810 8.770 ;
        RECT 46.410 7.310 46.585 8.450 ;
        RECT 50.640 7.310 50.815 8.570 ;
        RECT 51.225 8.540 51.395 10.150 ;
        RECT 51.595 10.090 51.770 10.600 ;
        RECT 52.025 10.050 52.200 10.600 ;
        RECT 53.390 10.085 53.560 10.595 ;
        RECT 54.380 10.085 54.550 10.595 ;
        RECT 63.585 10.110 63.760 10.600 ;
        RECT 51.165 8.370 51.395 8.540 ;
        RECT 51.595 8.570 51.765 9.520 ;
        RECT 51.165 7.310 51.335 8.370 ;
        RECT 51.595 7.310 51.770 8.570 ;
        RECT 52.025 8.450 52.195 10.050 ;
        RECT 63.585 9.940 63.755 10.110 ;
        RECT 64.540 10.090 64.715 10.600 ;
        RECT 64.970 10.050 65.145 10.600 ;
        RECT 69.200 10.110 69.375 10.600 ;
        RECT 69.725 10.320 69.895 10.600 ;
        RECT 69.725 10.150 69.955 10.320 ;
        RECT 52.955 9.425 53.185 9.625 ;
        RECT 63.585 9.610 63.995 9.940 ;
        RECT 52.955 9.395 53.485 9.425 ;
        RECT 53.015 9.255 53.485 9.395 ;
        RECT 54.005 9.255 54.475 9.425 ;
        RECT 53.015 8.565 53.185 9.255 ;
        RECT 53.385 8.790 53.555 8.885 ;
        RECT 54.005 8.790 54.175 9.255 ;
        RECT 63.585 9.100 63.755 9.610 ;
        RECT 53.385 8.610 54.175 8.790 ;
        RECT 52.025 7.310 52.200 8.450 ;
        RECT 53.385 7.305 53.560 8.610 ;
        RECT 54.005 8.565 54.175 8.610 ;
        RECT 54.375 8.450 54.545 8.885 ;
        RECT 63.585 8.770 63.995 9.100 ;
        RECT 63.585 8.570 63.755 8.770 ;
        RECT 64.540 8.570 64.710 9.520 ;
        RECT 54.375 7.305 54.550 8.450 ;
        RECT 63.585 7.310 63.760 8.570 ;
        RECT 64.540 7.310 64.715 8.570 ;
        RECT 64.970 8.450 65.140 10.050 ;
        RECT 69.200 9.940 69.370 10.110 ;
        RECT 69.200 9.610 69.610 9.940 ;
        RECT 69.200 9.100 69.370 9.610 ;
        RECT 69.200 8.770 69.610 9.100 ;
        RECT 69.200 8.570 69.370 8.770 ;
        RECT 64.970 7.310 65.145 8.450 ;
        RECT 69.200 7.310 69.375 8.570 ;
        RECT 69.785 8.540 69.955 10.150 ;
        RECT 70.155 10.090 70.330 10.600 ;
        RECT 70.585 10.050 70.760 10.600 ;
        RECT 71.950 10.085 72.120 10.595 ;
        RECT 72.940 10.085 73.110 10.595 ;
        RECT 82.145 10.110 82.320 10.600 ;
        RECT 69.725 8.370 69.955 8.540 ;
        RECT 70.155 8.570 70.325 9.520 ;
        RECT 69.725 7.310 69.895 8.370 ;
        RECT 70.155 7.310 70.330 8.570 ;
        RECT 70.585 8.450 70.755 10.050 ;
        RECT 82.145 9.940 82.315 10.110 ;
        RECT 83.100 10.090 83.275 10.600 ;
        RECT 83.530 10.050 83.705 10.600 ;
        RECT 87.760 10.110 87.935 10.600 ;
        RECT 88.285 10.320 88.455 10.600 ;
        RECT 88.285 10.150 88.515 10.320 ;
        RECT 71.515 9.425 71.745 9.625 ;
        RECT 82.145 9.610 82.555 9.940 ;
        RECT 71.515 9.395 72.045 9.425 ;
        RECT 71.575 9.255 72.045 9.395 ;
        RECT 72.565 9.255 73.035 9.425 ;
        RECT 71.575 8.565 71.745 9.255 ;
        RECT 71.945 8.790 72.115 8.885 ;
        RECT 72.565 8.790 72.735 9.255 ;
        RECT 82.145 9.100 82.315 9.610 ;
        RECT 71.945 8.610 72.735 8.790 ;
        RECT 70.585 7.310 70.760 8.450 ;
        RECT 71.945 7.305 72.120 8.610 ;
        RECT 72.565 8.565 72.735 8.610 ;
        RECT 72.935 8.450 73.105 8.885 ;
        RECT 82.145 8.770 82.555 9.100 ;
        RECT 82.145 8.570 82.315 8.770 ;
        RECT 83.100 8.570 83.270 9.520 ;
        RECT 72.935 7.305 73.110 8.450 ;
        RECT 82.145 7.310 82.320 8.570 ;
        RECT 83.100 7.310 83.275 8.570 ;
        RECT 83.530 8.450 83.700 10.050 ;
        RECT 87.760 9.940 87.930 10.110 ;
        RECT 87.760 9.610 88.170 9.940 ;
        RECT 87.760 9.100 87.930 9.610 ;
        RECT 87.760 8.770 88.170 9.100 ;
        RECT 87.760 8.570 87.930 8.770 ;
        RECT 83.530 7.310 83.705 8.450 ;
        RECT 87.760 7.310 87.935 8.570 ;
        RECT 88.345 8.540 88.515 10.150 ;
        RECT 88.715 10.090 88.890 10.600 ;
        RECT 89.145 10.050 89.320 10.600 ;
        RECT 90.510 10.085 90.680 10.595 ;
        RECT 91.500 10.085 91.670 10.595 ;
        RECT 100.705 10.110 100.880 10.600 ;
        RECT 88.285 8.370 88.515 8.540 ;
        RECT 88.715 8.570 88.885 9.520 ;
        RECT 88.285 7.310 88.455 8.370 ;
        RECT 88.715 7.310 88.890 8.570 ;
        RECT 89.145 8.450 89.315 10.050 ;
        RECT 100.705 9.940 100.875 10.110 ;
        RECT 101.660 10.090 101.835 10.600 ;
        RECT 102.090 10.050 102.265 10.600 ;
        RECT 106.320 10.110 106.495 10.600 ;
        RECT 106.845 10.320 107.015 10.600 ;
        RECT 106.845 10.150 107.075 10.320 ;
        RECT 90.075 9.425 90.305 9.625 ;
        RECT 100.705 9.610 101.115 9.940 ;
        RECT 90.075 9.395 90.605 9.425 ;
        RECT 90.135 9.255 90.605 9.395 ;
        RECT 91.125 9.255 91.595 9.425 ;
        RECT 90.135 8.565 90.305 9.255 ;
        RECT 90.505 8.790 90.675 8.885 ;
        RECT 91.125 8.790 91.295 9.255 ;
        RECT 100.705 9.100 100.875 9.610 ;
        RECT 90.505 8.610 91.295 8.790 ;
        RECT 89.145 7.310 89.320 8.450 ;
        RECT 90.505 7.305 90.680 8.610 ;
        RECT 91.125 8.565 91.295 8.610 ;
        RECT 91.495 8.450 91.665 8.885 ;
        RECT 100.705 8.770 101.115 9.100 ;
        RECT 100.705 8.570 100.875 8.770 ;
        RECT 101.660 8.570 101.830 9.520 ;
        RECT 91.495 7.305 91.670 8.450 ;
        RECT 100.705 7.310 100.880 8.570 ;
        RECT 101.660 7.310 101.835 8.570 ;
        RECT 102.090 8.450 102.260 10.050 ;
        RECT 106.320 9.940 106.490 10.110 ;
        RECT 106.320 9.610 106.730 9.940 ;
        RECT 106.320 9.100 106.490 9.610 ;
        RECT 106.320 8.770 106.730 9.100 ;
        RECT 106.320 8.570 106.490 8.770 ;
        RECT 102.090 7.310 102.265 8.450 ;
        RECT 106.320 7.310 106.495 8.570 ;
        RECT 106.905 8.540 107.075 10.150 ;
        RECT 107.275 10.090 107.450 10.600 ;
        RECT 107.705 10.050 107.880 10.600 ;
        RECT 109.070 10.085 109.240 10.595 ;
        RECT 110.060 10.085 110.230 10.595 ;
        RECT 106.845 8.370 107.075 8.540 ;
        RECT 107.275 8.570 107.445 9.520 ;
        RECT 106.845 7.310 107.015 8.370 ;
        RECT 107.275 7.310 107.450 8.570 ;
        RECT 107.705 8.450 107.875 10.050 ;
        RECT 108.635 9.425 108.865 9.625 ;
        RECT 108.635 9.395 109.165 9.425 ;
        RECT 108.695 9.255 109.165 9.395 ;
        RECT 109.685 9.255 110.155 9.425 ;
        RECT 108.695 8.565 108.865 9.255 ;
        RECT 109.065 8.790 109.235 8.885 ;
        RECT 109.685 8.790 109.855 9.255 ;
        RECT 109.065 8.610 109.855 8.790 ;
        RECT 107.705 7.310 107.880 8.450 ;
        RECT 109.065 7.305 109.240 8.610 ;
        RECT 109.685 8.565 109.855 8.610 ;
        RECT 110.055 8.450 110.225 8.885 ;
        RECT 110.055 7.305 110.230 8.450 ;
        RECT 18.875 4.575 19.045 4.935 ;
        RECT 19.835 4.605 20.005 4.765 ;
        RECT 21.795 4.685 21.965 4.795 ;
        RECT 19.215 4.435 20.005 4.605 ;
        RECT 20.755 4.515 22.045 4.685 ;
        RECT 19.215 4.375 19.385 4.435 ;
        RECT 19.115 4.205 19.385 4.375 ;
        RECT 19.835 4.345 20.005 4.435 ;
        RECT 22.275 4.345 22.445 4.765 ;
        RECT 22.755 4.435 22.925 4.795 ;
        RECT 23.675 4.515 24.165 4.685 ;
        RECT 19.115 4.135 19.285 4.205 ;
        RECT 18.875 3.865 19.285 4.135 ;
        RECT 19.115 3.785 19.285 3.865 ;
        RECT 19.595 3.785 19.765 4.115 ;
        RECT 20.745 3.865 21.325 4.035 ;
        RECT 20.745 3.785 20.915 3.865 ;
        RECT 21.555 3.785 21.725 4.235 ;
        RECT 23.275 4.035 23.445 4.515 ;
        RECT 23.995 4.345 25.005 4.515 ;
        RECT 25.195 4.435 25.365 5.075 ;
        RECT 25.715 4.775 25.885 5.105 ;
        RECT 26.675 4.905 27.325 5.075 ;
        RECT 27.035 4.515 27.325 4.905 ;
        RECT 28.035 4.905 28.325 5.075 ;
        RECT 24.835 4.115 25.005 4.345 ;
        RECT 25.715 4.375 25.885 4.515 ;
        RECT 27.155 4.435 27.325 4.515 ;
        RECT 25.715 4.205 26.605 4.375 ;
        RECT 27.675 4.345 27.845 4.765 ;
        RECT 28.035 4.515 28.205 4.905 ;
        RECT 28.875 4.515 29.845 4.685 ;
        RECT 28.035 4.345 28.325 4.515 ;
        RECT 28.875 4.345 29.045 4.515 ;
        RECT 22.435 3.865 22.925 4.035 ;
        RECT 23.275 3.865 23.765 4.035 ;
        RECT 22.755 3.785 22.925 3.865 ;
        RECT 23.995 3.785 24.165 4.115 ;
        RECT 24.475 3.785 24.645 4.115 ;
        RECT 24.835 3.865 25.125 4.115 ;
        RECT 24.955 3.785 25.125 3.865 ;
        RECT 25.715 3.865 26.205 4.035 ;
        RECT 25.715 3.785 25.885 3.865 ;
        RECT 26.435 3.785 26.605 4.205 ;
        RECT 27.155 4.135 27.325 4.235 ;
        RECT 26.915 4.035 27.325 4.135 ;
        RECT 28.035 4.035 28.205 4.345 ;
        RECT 26.835 3.965 27.325 4.035 ;
        RECT 26.835 3.865 27.165 3.965 ;
        RECT 27.835 3.865 28.205 4.035 ;
        RECT 28.395 4.035 28.565 4.115 ;
        RECT 28.395 3.865 29.125 4.035 ;
        RECT 28.395 3.785 28.565 3.865 ;
        RECT 29.355 3.785 29.525 4.235 ;
        RECT 32.080 3.895 32.255 5.155 ;
        RECT 32.605 4.095 32.775 5.155 ;
        RECT 32.605 3.925 32.835 4.095 ;
        RECT 32.080 3.695 32.250 3.895 ;
        RECT 18.875 3.045 19.045 3.395 ;
        RECT 19.835 3.295 20.005 3.395 ;
        RECT 22.275 3.295 22.445 3.395 ;
        RECT 23.755 3.295 23.925 3.395 ;
        RECT 19.835 3.125 20.565 3.295 ;
        RECT 21.715 3.125 22.445 3.295 ;
        RECT 23.195 3.125 23.925 3.295 ;
        RECT 24.715 3.045 24.885 3.395 ;
        RECT 25.715 3.045 25.885 3.395 ;
        RECT 26.675 3.045 26.845 3.395 ;
        RECT 28.155 3.045 28.325 3.395 ;
        RECT 29.115 3.045 29.285 3.395 ;
        RECT 32.080 3.365 32.490 3.695 ;
        RECT 32.080 2.855 32.250 3.365 ;
        RECT 32.080 2.525 32.490 2.855 ;
        RECT 32.080 2.355 32.250 2.525 ;
        RECT 32.080 1.865 32.255 2.355 ;
        RECT 32.665 2.315 32.835 3.925 ;
        RECT 33.035 3.895 33.210 5.155 ;
        RECT 33.465 4.015 33.640 5.155 ;
        RECT 33.035 2.945 33.205 3.895 ;
        RECT 33.465 2.415 33.635 4.015 ;
        RECT 34.455 3.210 34.625 3.900 ;
        RECT 34.825 3.860 35.000 5.160 ;
        RECT 37.435 4.575 37.605 4.935 ;
        RECT 38.395 4.605 38.565 4.765 ;
        RECT 40.355 4.685 40.525 4.795 ;
        RECT 37.775 4.435 38.565 4.605 ;
        RECT 39.315 4.515 40.605 4.685 ;
        RECT 37.775 4.375 37.945 4.435 ;
        RECT 37.675 4.205 37.945 4.375 ;
        RECT 38.395 4.345 38.565 4.435 ;
        RECT 40.835 4.345 41.005 4.765 ;
        RECT 41.315 4.435 41.485 4.795 ;
        RECT 42.235 4.515 42.725 4.685 ;
        RECT 37.675 4.135 37.845 4.205 ;
        RECT 35.440 3.860 35.610 3.900 ;
        RECT 37.435 3.865 37.845 4.135 ;
        RECT 34.825 3.665 35.610 3.860 ;
        RECT 37.675 3.785 37.845 3.865 ;
        RECT 38.155 3.785 38.325 4.115 ;
        RECT 39.305 3.865 39.885 4.035 ;
        RECT 39.305 3.785 39.475 3.865 ;
        RECT 40.115 3.785 40.285 4.235 ;
        RECT 41.835 4.035 42.005 4.515 ;
        RECT 42.555 4.345 43.565 4.515 ;
        RECT 43.755 4.435 43.925 5.075 ;
        RECT 44.275 4.775 44.445 5.105 ;
        RECT 45.235 4.905 45.885 5.075 ;
        RECT 45.595 4.515 45.885 4.905 ;
        RECT 46.595 4.905 46.885 5.075 ;
        RECT 43.395 4.115 43.565 4.345 ;
        RECT 44.275 4.375 44.445 4.515 ;
        RECT 45.715 4.435 45.885 4.515 ;
        RECT 44.275 4.205 45.165 4.375 ;
        RECT 46.235 4.345 46.405 4.765 ;
        RECT 46.595 4.515 46.765 4.905 ;
        RECT 47.435 4.515 48.405 4.685 ;
        RECT 46.595 4.345 46.885 4.515 ;
        RECT 47.435 4.345 47.605 4.515 ;
        RECT 40.995 3.865 41.485 4.035 ;
        RECT 41.835 3.865 42.325 4.035 ;
        RECT 41.315 3.785 41.485 3.865 ;
        RECT 42.555 3.785 42.725 4.115 ;
        RECT 43.035 3.785 43.205 4.115 ;
        RECT 43.395 3.865 43.685 4.115 ;
        RECT 43.515 3.785 43.685 3.865 ;
        RECT 44.275 3.865 44.765 4.035 ;
        RECT 44.275 3.785 44.445 3.865 ;
        RECT 44.995 3.785 45.165 4.205 ;
        RECT 45.715 4.135 45.885 4.235 ;
        RECT 45.475 4.035 45.885 4.135 ;
        RECT 46.595 4.035 46.765 4.345 ;
        RECT 45.395 3.965 45.885 4.035 ;
        RECT 45.395 3.865 45.725 3.965 ;
        RECT 46.395 3.865 46.765 4.035 ;
        RECT 46.955 4.035 47.125 4.115 ;
        RECT 46.955 3.865 47.685 4.035 ;
        RECT 46.955 3.785 47.125 3.865 ;
        RECT 47.915 3.785 48.085 4.235 ;
        RECT 50.640 3.895 50.815 5.155 ;
        RECT 51.165 4.095 51.335 5.155 ;
        RECT 51.165 3.925 51.395 4.095 ;
        RECT 34.825 3.580 34.995 3.665 ;
        RECT 35.440 3.210 35.610 3.665 ;
        RECT 50.640 3.695 50.810 3.895 ;
        RECT 34.455 3.185 34.925 3.210 ;
        RECT 34.400 3.040 34.925 3.185 ;
        RECT 35.440 3.040 35.910 3.210 ;
        RECT 37.435 3.045 37.605 3.395 ;
        RECT 38.395 3.295 38.565 3.395 ;
        RECT 40.835 3.295 41.005 3.395 ;
        RECT 42.315 3.295 42.485 3.395 ;
        RECT 38.395 3.125 39.125 3.295 ;
        RECT 40.275 3.125 41.005 3.295 ;
        RECT 41.755 3.125 42.485 3.295 ;
        RECT 43.275 3.045 43.445 3.395 ;
        RECT 44.275 3.045 44.445 3.395 ;
        RECT 45.235 3.045 45.405 3.395 ;
        RECT 46.715 3.045 46.885 3.395 ;
        RECT 47.675 3.045 47.845 3.395 ;
        RECT 50.640 3.365 51.050 3.695 ;
        RECT 34.400 2.955 34.630 3.040 ;
        RECT 50.640 2.855 50.810 3.365 ;
        RECT 50.640 2.525 51.050 2.855 ;
        RECT 32.605 2.145 32.835 2.315 ;
        RECT 32.605 1.865 32.775 2.145 ;
        RECT 33.035 1.865 33.210 2.375 ;
        RECT 33.465 1.865 33.640 2.415 ;
        RECT 34.830 1.870 35.000 2.380 ;
        RECT 50.640 2.355 50.810 2.525 ;
        RECT 50.640 1.865 50.815 2.355 ;
        RECT 51.225 2.315 51.395 3.925 ;
        RECT 51.595 3.895 51.770 5.155 ;
        RECT 52.025 4.015 52.200 5.155 ;
        RECT 51.595 2.945 51.765 3.895 ;
        RECT 52.025 2.415 52.195 4.015 ;
        RECT 53.015 3.210 53.185 3.900 ;
        RECT 53.385 3.860 53.560 5.160 ;
        RECT 55.995 4.575 56.165 4.935 ;
        RECT 56.955 4.605 57.125 4.765 ;
        RECT 58.915 4.685 59.085 4.795 ;
        RECT 56.335 4.435 57.125 4.605 ;
        RECT 57.875 4.515 59.165 4.685 ;
        RECT 56.335 4.375 56.505 4.435 ;
        RECT 56.235 4.205 56.505 4.375 ;
        RECT 56.955 4.345 57.125 4.435 ;
        RECT 59.395 4.345 59.565 4.765 ;
        RECT 59.875 4.435 60.045 4.795 ;
        RECT 60.795 4.515 61.285 4.685 ;
        RECT 56.235 4.135 56.405 4.205 ;
        RECT 54.000 3.860 54.170 3.900 ;
        RECT 55.995 3.865 56.405 4.135 ;
        RECT 53.385 3.665 54.170 3.860 ;
        RECT 56.235 3.785 56.405 3.865 ;
        RECT 56.715 3.785 56.885 4.115 ;
        RECT 57.865 3.865 58.445 4.035 ;
        RECT 57.865 3.785 58.035 3.865 ;
        RECT 58.675 3.785 58.845 4.235 ;
        RECT 60.395 4.035 60.565 4.515 ;
        RECT 61.115 4.345 62.125 4.515 ;
        RECT 62.315 4.435 62.485 5.075 ;
        RECT 62.835 4.775 63.005 5.105 ;
        RECT 63.795 4.905 64.445 5.075 ;
        RECT 64.155 4.515 64.445 4.905 ;
        RECT 65.155 4.905 65.445 5.075 ;
        RECT 61.955 4.115 62.125 4.345 ;
        RECT 62.835 4.375 63.005 4.515 ;
        RECT 64.275 4.435 64.445 4.515 ;
        RECT 62.835 4.205 63.725 4.375 ;
        RECT 64.795 4.345 64.965 4.765 ;
        RECT 65.155 4.515 65.325 4.905 ;
        RECT 65.995 4.515 66.965 4.685 ;
        RECT 65.155 4.345 65.445 4.515 ;
        RECT 65.995 4.345 66.165 4.515 ;
        RECT 59.555 3.865 60.045 4.035 ;
        RECT 60.395 3.865 60.885 4.035 ;
        RECT 59.875 3.785 60.045 3.865 ;
        RECT 61.115 3.785 61.285 4.115 ;
        RECT 61.595 3.785 61.765 4.115 ;
        RECT 61.955 3.865 62.245 4.115 ;
        RECT 62.075 3.785 62.245 3.865 ;
        RECT 62.835 3.865 63.325 4.035 ;
        RECT 62.835 3.785 63.005 3.865 ;
        RECT 63.555 3.785 63.725 4.205 ;
        RECT 64.275 4.135 64.445 4.235 ;
        RECT 64.035 4.035 64.445 4.135 ;
        RECT 65.155 4.035 65.325 4.345 ;
        RECT 63.955 3.965 64.445 4.035 ;
        RECT 63.955 3.865 64.285 3.965 ;
        RECT 64.955 3.865 65.325 4.035 ;
        RECT 65.515 4.035 65.685 4.115 ;
        RECT 65.515 3.865 66.245 4.035 ;
        RECT 65.515 3.785 65.685 3.865 ;
        RECT 66.475 3.785 66.645 4.235 ;
        RECT 69.200 3.895 69.375 5.155 ;
        RECT 69.725 4.095 69.895 5.155 ;
        RECT 69.725 3.925 69.955 4.095 ;
        RECT 53.385 3.580 53.555 3.665 ;
        RECT 54.000 3.210 54.170 3.665 ;
        RECT 69.200 3.695 69.370 3.895 ;
        RECT 53.015 3.185 53.485 3.210 ;
        RECT 52.960 3.040 53.485 3.185 ;
        RECT 54.000 3.040 54.470 3.210 ;
        RECT 55.995 3.045 56.165 3.395 ;
        RECT 56.955 3.295 57.125 3.395 ;
        RECT 59.395 3.295 59.565 3.395 ;
        RECT 60.875 3.295 61.045 3.395 ;
        RECT 56.955 3.125 57.685 3.295 ;
        RECT 58.835 3.125 59.565 3.295 ;
        RECT 60.315 3.125 61.045 3.295 ;
        RECT 61.835 3.045 62.005 3.395 ;
        RECT 62.835 3.045 63.005 3.395 ;
        RECT 63.795 3.045 63.965 3.395 ;
        RECT 65.275 3.045 65.445 3.395 ;
        RECT 66.235 3.045 66.405 3.395 ;
        RECT 69.200 3.365 69.610 3.695 ;
        RECT 52.960 2.955 53.190 3.040 ;
        RECT 69.200 2.855 69.370 3.365 ;
        RECT 69.200 2.525 69.610 2.855 ;
        RECT 51.165 2.145 51.395 2.315 ;
        RECT 51.165 1.865 51.335 2.145 ;
        RECT 51.595 1.865 51.770 2.375 ;
        RECT 52.025 1.865 52.200 2.415 ;
        RECT 53.390 1.870 53.560 2.380 ;
        RECT 69.200 2.355 69.370 2.525 ;
        RECT 69.200 1.865 69.375 2.355 ;
        RECT 69.785 2.315 69.955 3.925 ;
        RECT 70.155 3.895 70.330 5.155 ;
        RECT 70.585 4.015 70.760 5.155 ;
        RECT 70.155 2.945 70.325 3.895 ;
        RECT 70.585 2.415 70.755 4.015 ;
        RECT 71.575 3.210 71.745 3.900 ;
        RECT 71.945 3.860 72.120 5.160 ;
        RECT 74.555 4.575 74.725 4.935 ;
        RECT 75.515 4.605 75.685 4.765 ;
        RECT 77.475 4.685 77.645 4.795 ;
        RECT 74.895 4.435 75.685 4.605 ;
        RECT 76.435 4.515 77.725 4.685 ;
        RECT 74.895 4.375 75.065 4.435 ;
        RECT 74.795 4.205 75.065 4.375 ;
        RECT 75.515 4.345 75.685 4.435 ;
        RECT 77.955 4.345 78.125 4.765 ;
        RECT 78.435 4.435 78.605 4.795 ;
        RECT 79.355 4.515 79.845 4.685 ;
        RECT 74.795 4.135 74.965 4.205 ;
        RECT 72.560 3.860 72.730 3.900 ;
        RECT 74.555 3.865 74.965 4.135 ;
        RECT 71.945 3.665 72.730 3.860 ;
        RECT 74.795 3.785 74.965 3.865 ;
        RECT 75.275 3.785 75.445 4.115 ;
        RECT 76.425 3.865 77.005 4.035 ;
        RECT 76.425 3.785 76.595 3.865 ;
        RECT 77.235 3.785 77.405 4.235 ;
        RECT 78.955 4.035 79.125 4.515 ;
        RECT 79.675 4.345 80.685 4.515 ;
        RECT 80.875 4.435 81.045 5.075 ;
        RECT 81.395 4.775 81.565 5.105 ;
        RECT 82.355 4.905 83.005 5.075 ;
        RECT 82.715 4.515 83.005 4.905 ;
        RECT 83.715 4.905 84.005 5.075 ;
        RECT 80.515 4.115 80.685 4.345 ;
        RECT 81.395 4.375 81.565 4.515 ;
        RECT 82.835 4.435 83.005 4.515 ;
        RECT 81.395 4.205 82.285 4.375 ;
        RECT 83.355 4.345 83.525 4.765 ;
        RECT 83.715 4.515 83.885 4.905 ;
        RECT 84.555 4.515 85.525 4.685 ;
        RECT 83.715 4.345 84.005 4.515 ;
        RECT 84.555 4.345 84.725 4.515 ;
        RECT 78.115 3.865 78.605 4.035 ;
        RECT 78.955 3.865 79.445 4.035 ;
        RECT 78.435 3.785 78.605 3.865 ;
        RECT 79.675 3.785 79.845 4.115 ;
        RECT 80.155 3.785 80.325 4.115 ;
        RECT 80.515 3.865 80.805 4.115 ;
        RECT 80.635 3.785 80.805 3.865 ;
        RECT 81.395 3.865 81.885 4.035 ;
        RECT 81.395 3.785 81.565 3.865 ;
        RECT 82.115 3.785 82.285 4.205 ;
        RECT 82.835 4.135 83.005 4.235 ;
        RECT 82.595 4.035 83.005 4.135 ;
        RECT 83.715 4.035 83.885 4.345 ;
        RECT 82.515 3.965 83.005 4.035 ;
        RECT 82.515 3.865 82.845 3.965 ;
        RECT 83.515 3.865 83.885 4.035 ;
        RECT 84.075 4.035 84.245 4.115 ;
        RECT 84.075 3.865 84.805 4.035 ;
        RECT 84.075 3.785 84.245 3.865 ;
        RECT 85.035 3.785 85.205 4.235 ;
        RECT 87.760 3.895 87.935 5.155 ;
        RECT 88.285 4.095 88.455 5.155 ;
        RECT 88.285 3.925 88.515 4.095 ;
        RECT 71.945 3.580 72.115 3.665 ;
        RECT 72.560 3.210 72.730 3.665 ;
        RECT 87.760 3.695 87.930 3.895 ;
        RECT 71.575 3.185 72.045 3.210 ;
        RECT 71.520 3.040 72.045 3.185 ;
        RECT 72.560 3.040 73.030 3.210 ;
        RECT 74.555 3.045 74.725 3.395 ;
        RECT 75.515 3.295 75.685 3.395 ;
        RECT 77.955 3.295 78.125 3.395 ;
        RECT 79.435 3.295 79.605 3.395 ;
        RECT 75.515 3.125 76.245 3.295 ;
        RECT 77.395 3.125 78.125 3.295 ;
        RECT 78.875 3.125 79.605 3.295 ;
        RECT 80.395 3.045 80.565 3.395 ;
        RECT 81.395 3.045 81.565 3.395 ;
        RECT 82.355 3.045 82.525 3.395 ;
        RECT 83.835 3.045 84.005 3.395 ;
        RECT 84.795 3.045 84.965 3.395 ;
        RECT 87.760 3.365 88.170 3.695 ;
        RECT 71.520 2.955 71.750 3.040 ;
        RECT 87.760 2.855 87.930 3.365 ;
        RECT 87.760 2.525 88.170 2.855 ;
        RECT 69.725 2.145 69.955 2.315 ;
        RECT 69.725 1.865 69.895 2.145 ;
        RECT 70.155 1.865 70.330 2.375 ;
        RECT 70.585 1.865 70.760 2.415 ;
        RECT 71.950 1.870 72.120 2.380 ;
        RECT 87.760 2.355 87.930 2.525 ;
        RECT 87.760 1.865 87.935 2.355 ;
        RECT 88.345 2.315 88.515 3.925 ;
        RECT 88.715 3.895 88.890 5.155 ;
        RECT 89.145 4.015 89.320 5.155 ;
        RECT 88.715 2.945 88.885 3.895 ;
        RECT 89.145 2.415 89.315 4.015 ;
        RECT 90.135 3.210 90.305 3.900 ;
        RECT 90.505 3.860 90.680 5.160 ;
        RECT 93.115 4.575 93.285 4.935 ;
        RECT 94.075 4.605 94.245 4.765 ;
        RECT 96.035 4.685 96.205 4.795 ;
        RECT 93.455 4.435 94.245 4.605 ;
        RECT 94.995 4.515 96.285 4.685 ;
        RECT 93.455 4.375 93.625 4.435 ;
        RECT 93.355 4.205 93.625 4.375 ;
        RECT 94.075 4.345 94.245 4.435 ;
        RECT 96.515 4.345 96.685 4.765 ;
        RECT 96.995 4.435 97.165 4.795 ;
        RECT 97.915 4.515 98.405 4.685 ;
        RECT 93.355 4.135 93.525 4.205 ;
        RECT 91.120 3.860 91.290 3.900 ;
        RECT 93.115 3.865 93.525 4.135 ;
        RECT 90.505 3.665 91.290 3.860 ;
        RECT 93.355 3.785 93.525 3.865 ;
        RECT 93.835 3.785 94.005 4.115 ;
        RECT 94.985 3.865 95.565 4.035 ;
        RECT 94.985 3.785 95.155 3.865 ;
        RECT 95.795 3.785 95.965 4.235 ;
        RECT 97.515 4.035 97.685 4.515 ;
        RECT 98.235 4.345 99.245 4.515 ;
        RECT 99.435 4.435 99.605 5.075 ;
        RECT 99.955 4.775 100.125 5.105 ;
        RECT 100.915 4.905 101.565 5.075 ;
        RECT 101.275 4.515 101.565 4.905 ;
        RECT 102.275 4.905 102.565 5.075 ;
        RECT 99.075 4.115 99.245 4.345 ;
        RECT 99.955 4.375 100.125 4.515 ;
        RECT 101.395 4.435 101.565 4.515 ;
        RECT 99.955 4.205 100.845 4.375 ;
        RECT 101.915 4.345 102.085 4.765 ;
        RECT 102.275 4.515 102.445 4.905 ;
        RECT 103.115 4.515 104.085 4.685 ;
        RECT 102.275 4.345 102.565 4.515 ;
        RECT 103.115 4.345 103.285 4.515 ;
        RECT 96.675 3.865 97.165 4.035 ;
        RECT 97.515 3.865 98.005 4.035 ;
        RECT 96.995 3.785 97.165 3.865 ;
        RECT 98.235 3.785 98.405 4.115 ;
        RECT 98.715 3.785 98.885 4.115 ;
        RECT 99.075 3.865 99.365 4.115 ;
        RECT 99.195 3.785 99.365 3.865 ;
        RECT 99.955 3.865 100.445 4.035 ;
        RECT 99.955 3.785 100.125 3.865 ;
        RECT 100.675 3.785 100.845 4.205 ;
        RECT 101.395 4.135 101.565 4.235 ;
        RECT 101.155 4.035 101.565 4.135 ;
        RECT 102.275 4.035 102.445 4.345 ;
        RECT 101.075 3.965 101.565 4.035 ;
        RECT 101.075 3.865 101.405 3.965 ;
        RECT 102.075 3.865 102.445 4.035 ;
        RECT 102.635 4.035 102.805 4.115 ;
        RECT 102.635 3.865 103.365 4.035 ;
        RECT 102.635 3.785 102.805 3.865 ;
        RECT 103.595 3.785 103.765 4.235 ;
        RECT 106.320 3.895 106.495 5.155 ;
        RECT 106.845 4.095 107.015 5.155 ;
        RECT 106.845 3.925 107.075 4.095 ;
        RECT 90.505 3.580 90.675 3.665 ;
        RECT 91.120 3.210 91.290 3.665 ;
        RECT 106.320 3.695 106.490 3.895 ;
        RECT 90.135 3.185 90.605 3.210 ;
        RECT 90.080 3.040 90.605 3.185 ;
        RECT 91.120 3.040 91.590 3.210 ;
        RECT 93.115 3.045 93.285 3.395 ;
        RECT 94.075 3.295 94.245 3.395 ;
        RECT 96.515 3.295 96.685 3.395 ;
        RECT 97.995 3.295 98.165 3.395 ;
        RECT 94.075 3.125 94.805 3.295 ;
        RECT 95.955 3.125 96.685 3.295 ;
        RECT 97.435 3.125 98.165 3.295 ;
        RECT 98.955 3.045 99.125 3.395 ;
        RECT 99.955 3.045 100.125 3.395 ;
        RECT 100.915 3.045 101.085 3.395 ;
        RECT 102.395 3.045 102.565 3.395 ;
        RECT 103.355 3.045 103.525 3.395 ;
        RECT 106.320 3.365 106.730 3.695 ;
        RECT 90.080 2.955 90.310 3.040 ;
        RECT 106.320 2.855 106.490 3.365 ;
        RECT 106.320 2.525 106.730 2.855 ;
        RECT 88.285 2.145 88.515 2.315 ;
        RECT 88.285 1.865 88.455 2.145 ;
        RECT 88.715 1.865 88.890 2.375 ;
        RECT 89.145 1.865 89.320 2.415 ;
        RECT 90.510 1.870 90.680 2.380 ;
        RECT 106.320 2.355 106.490 2.525 ;
        RECT 106.320 1.865 106.495 2.355 ;
        RECT 106.905 2.315 107.075 3.925 ;
        RECT 107.275 3.895 107.450 5.155 ;
        RECT 107.705 4.015 107.880 5.155 ;
        RECT 107.275 2.945 107.445 3.895 ;
        RECT 107.705 2.415 107.875 4.015 ;
        RECT 108.695 3.210 108.865 3.900 ;
        RECT 109.065 3.860 109.240 5.160 ;
        RECT 109.680 3.860 109.850 3.900 ;
        RECT 109.065 3.665 109.850 3.860 ;
        RECT 109.065 3.580 109.235 3.665 ;
        RECT 109.680 3.210 109.850 3.665 ;
        RECT 108.695 3.185 109.165 3.210 ;
        RECT 108.640 3.040 109.165 3.185 ;
        RECT 109.680 3.040 110.150 3.210 ;
        RECT 108.640 2.955 108.870 3.040 ;
        RECT 106.845 2.145 107.075 2.315 ;
        RECT 106.845 1.865 107.015 2.145 ;
        RECT 107.275 1.865 107.450 2.375 ;
        RECT 107.705 1.865 107.880 2.415 ;
        RECT 109.070 1.870 109.240 2.380 ;
      LAYER met1 ;
        RECT 16.545 10.060 16.835 10.290 ;
        RECT 27.360 10.060 27.650 10.290 ;
        RECT 32.975 10.060 33.265 10.290 ;
        RECT 16.605 9.610 16.775 10.060 ;
        RECT 27.420 9.715 27.590 10.060 ;
        RECT 16.515 9.320 16.865 9.610 ;
        RECT 27.320 9.345 27.700 9.715 ;
        RECT 33.035 9.580 33.205 10.060 ;
        RECT 34.765 10.025 35.060 10.285 ;
        RECT 35.755 10.025 36.050 10.285 ;
        RECT 45.920 10.060 46.210 10.290 ;
        RECT 51.535 10.060 51.825 10.290 ;
        RECT 34.395 9.655 34.625 9.685 ;
        RECT 34.365 9.580 34.655 9.655 ;
        RECT 33.035 9.550 34.655 9.580 ;
        RECT 32.975 9.410 34.655 9.550 ;
        RECT 27.360 9.320 27.650 9.345 ;
        RECT 32.975 9.320 33.265 9.410 ;
        RECT 34.365 9.350 34.655 9.410 ;
        RECT 34.395 9.335 34.625 9.350 ;
        RECT 27.995 9.180 28.345 9.245 ;
        RECT 33.430 9.180 33.755 9.270 ;
        RECT 27.790 9.150 28.345 9.180 ;
        RECT 33.405 9.150 33.755 9.180 ;
        RECT 27.620 9.145 28.345 9.150 ;
        RECT 33.235 9.145 33.755 9.150 ;
        RECT 27.620 8.975 33.755 9.145 ;
        RECT 27.790 8.950 28.345 8.975 ;
        RECT 33.405 8.950 33.755 8.975 ;
        RECT 27.995 8.895 28.345 8.950 ;
        RECT 33.430 8.945 33.755 8.950 ;
        RECT 34.825 8.925 34.995 10.025 ;
        RECT 35.815 9.295 35.985 10.025 ;
        RECT 45.980 9.715 46.150 10.060 ;
        RECT 45.880 9.345 46.260 9.715 ;
        RECT 51.595 9.580 51.765 10.060 ;
        RECT 53.325 10.025 53.620 10.285 ;
        RECT 54.315 10.025 54.610 10.285 ;
        RECT 64.480 10.060 64.770 10.290 ;
        RECT 70.095 10.060 70.385 10.290 ;
        RECT 52.955 9.655 53.185 9.685 ;
        RECT 52.925 9.580 53.215 9.655 ;
        RECT 51.595 9.550 53.215 9.580 ;
        RECT 51.535 9.410 53.215 9.550 ;
        RECT 45.920 9.320 46.210 9.345 ;
        RECT 51.535 9.320 51.825 9.410 ;
        RECT 52.925 9.350 53.215 9.410 ;
        RECT 52.955 9.335 53.185 9.350 ;
        RECT 35.810 8.945 36.160 9.295 ;
        RECT 46.555 9.180 46.905 9.250 ;
        RECT 51.990 9.180 52.315 9.270 ;
        RECT 46.350 9.150 46.905 9.180 ;
        RECT 51.965 9.150 52.315 9.180 ;
        RECT 46.180 9.145 46.905 9.150 ;
        RECT 51.795 9.145 52.315 9.150 ;
        RECT 46.180 8.975 52.315 9.145 ;
        RECT 46.350 8.950 46.905 8.975 ;
        RECT 51.965 8.950 52.315 8.975 ;
        RECT 35.810 8.925 36.105 8.945 ;
        RECT 34.765 8.920 34.995 8.925 ;
        RECT 16.140 8.790 16.490 8.865 ;
        RECT 32.630 8.820 32.950 8.835 ;
        RECT 32.605 8.790 32.950 8.820 ;
        RECT 16.000 8.620 16.490 8.790 ;
        RECT 32.430 8.620 32.950 8.790 ;
        RECT 34.765 8.685 35.055 8.920 ;
        RECT 35.755 8.855 36.105 8.925 ;
        RECT 46.555 8.900 46.905 8.950 ;
        RECT 51.990 8.945 52.315 8.950 ;
        RECT 53.385 8.925 53.555 10.025 ;
        RECT 54.375 9.305 54.545 10.025 ;
        RECT 64.540 9.715 64.710 10.060 ;
        RECT 64.440 9.345 64.820 9.715 ;
        RECT 70.155 9.580 70.325 10.060 ;
        RECT 71.885 10.025 72.180 10.285 ;
        RECT 72.875 10.025 73.170 10.285 ;
        RECT 83.040 10.060 83.330 10.290 ;
        RECT 88.655 10.060 88.945 10.290 ;
        RECT 71.515 9.655 71.745 9.685 ;
        RECT 71.485 9.580 71.775 9.655 ;
        RECT 70.155 9.550 71.775 9.580 ;
        RECT 70.095 9.410 71.775 9.550 ;
        RECT 64.480 9.320 64.770 9.345 ;
        RECT 70.095 9.320 70.385 9.410 ;
        RECT 71.485 9.350 71.775 9.410 ;
        RECT 71.515 9.335 71.745 9.350 ;
        RECT 54.365 8.950 54.720 9.305 ;
        RECT 65.110 9.180 65.460 9.255 ;
        RECT 70.550 9.180 70.875 9.270 ;
        RECT 64.910 9.150 65.460 9.180 ;
        RECT 70.525 9.150 70.875 9.180 ;
        RECT 64.740 9.145 65.460 9.150 ;
        RECT 70.355 9.145 70.875 9.150 ;
        RECT 64.740 8.975 70.875 9.145 ;
        RECT 64.910 8.950 65.460 8.975 ;
        RECT 70.525 8.950 70.875 8.975 ;
        RECT 54.365 8.925 54.665 8.950 ;
        RECT 53.325 8.920 53.555 8.925 ;
        RECT 35.755 8.685 36.045 8.855 ;
        RECT 51.190 8.820 51.510 8.835 ;
        RECT 51.165 8.790 51.510 8.820 ;
        RECT 50.990 8.620 51.510 8.790 ;
        RECT 53.325 8.685 53.615 8.920 ;
        RECT 54.315 8.855 54.665 8.925 ;
        RECT 65.110 8.905 65.460 8.950 ;
        RECT 70.550 8.945 70.875 8.950 ;
        RECT 71.945 8.925 72.115 10.025 ;
        RECT 72.935 9.295 73.105 10.025 ;
        RECT 83.100 9.715 83.270 10.060 ;
        RECT 83.000 9.345 83.380 9.715 ;
        RECT 88.715 9.580 88.885 10.060 ;
        RECT 90.445 10.025 90.740 10.285 ;
        RECT 91.435 10.025 91.730 10.285 ;
        RECT 101.600 10.060 101.890 10.290 ;
        RECT 107.215 10.060 107.505 10.290 ;
        RECT 90.075 9.655 90.305 9.685 ;
        RECT 90.045 9.580 90.335 9.655 ;
        RECT 88.715 9.550 90.335 9.580 ;
        RECT 88.655 9.410 90.335 9.550 ;
        RECT 83.040 9.320 83.330 9.345 ;
        RECT 88.655 9.320 88.945 9.410 ;
        RECT 90.045 9.350 90.335 9.410 ;
        RECT 90.075 9.335 90.305 9.350 ;
        RECT 72.885 8.945 73.235 9.295 ;
        RECT 83.670 9.180 84.020 9.250 ;
        RECT 89.110 9.180 89.435 9.270 ;
        RECT 83.470 9.150 84.020 9.180 ;
        RECT 89.085 9.150 89.435 9.180 ;
        RECT 83.300 9.145 84.020 9.150 ;
        RECT 88.915 9.145 89.435 9.150 ;
        RECT 83.300 8.975 89.435 9.145 ;
        RECT 83.470 8.950 84.020 8.975 ;
        RECT 89.085 8.950 89.435 8.975 ;
        RECT 72.885 8.925 73.225 8.945 ;
        RECT 71.885 8.920 72.115 8.925 ;
        RECT 54.315 8.685 54.605 8.855 ;
        RECT 69.750 8.820 70.070 8.835 ;
        RECT 69.725 8.790 70.070 8.820 ;
        RECT 69.550 8.620 70.070 8.790 ;
        RECT 71.885 8.685 72.175 8.920 ;
        RECT 72.875 8.855 73.225 8.925 ;
        RECT 83.670 8.900 84.020 8.950 ;
        RECT 89.110 8.945 89.435 8.950 ;
        RECT 90.505 8.925 90.675 10.025 ;
        RECT 91.495 9.295 91.665 10.025 ;
        RECT 101.660 9.715 101.830 10.060 ;
        RECT 101.560 9.345 101.940 9.715 ;
        RECT 107.275 9.580 107.445 10.060 ;
        RECT 109.005 10.025 109.300 10.285 ;
        RECT 109.995 10.025 110.290 10.285 ;
        RECT 108.635 9.655 108.865 9.685 ;
        RECT 108.605 9.580 108.895 9.655 ;
        RECT 107.275 9.550 108.895 9.580 ;
        RECT 107.215 9.410 108.895 9.550 ;
        RECT 101.600 9.320 101.890 9.345 ;
        RECT 107.215 9.320 107.505 9.410 ;
        RECT 108.605 9.350 108.895 9.410 ;
        RECT 108.635 9.335 108.865 9.350 ;
        RECT 91.445 8.945 91.795 9.295 ;
        RECT 102.230 9.180 102.580 9.250 ;
        RECT 107.670 9.180 107.995 9.270 ;
        RECT 102.030 9.150 102.580 9.180 ;
        RECT 107.645 9.150 107.995 9.180 ;
        RECT 101.860 9.145 102.580 9.150 ;
        RECT 107.475 9.145 107.995 9.150 ;
        RECT 101.860 8.975 107.995 9.145 ;
        RECT 102.030 8.950 102.580 8.975 ;
        RECT 107.645 8.950 107.995 8.975 ;
        RECT 91.445 8.925 91.785 8.945 ;
        RECT 90.445 8.920 90.675 8.925 ;
        RECT 72.875 8.685 73.165 8.855 ;
        RECT 88.310 8.820 88.630 8.835 ;
        RECT 88.285 8.790 88.630 8.820 ;
        RECT 88.110 8.620 88.630 8.790 ;
        RECT 90.445 8.685 90.735 8.920 ;
        RECT 91.435 8.855 91.785 8.925 ;
        RECT 102.230 8.900 102.580 8.950 ;
        RECT 107.670 8.945 107.995 8.950 ;
        RECT 109.065 8.925 109.235 10.025 ;
        RECT 110.030 10.000 110.290 10.025 ;
        RECT 110.030 9.915 110.350 10.000 ;
        RECT 110.030 9.565 110.380 9.915 ;
        RECT 110.055 8.925 110.225 9.565 ;
        RECT 109.005 8.920 109.235 8.925 ;
        RECT 109.995 8.920 110.225 8.925 ;
        RECT 91.435 8.685 91.725 8.855 ;
        RECT 106.870 8.820 107.190 8.835 ;
        RECT 106.845 8.790 107.190 8.820 ;
        RECT 106.670 8.620 107.190 8.790 ;
        RECT 109.005 8.685 109.295 8.920 ;
        RECT 109.995 8.685 110.285 8.920 ;
        RECT 16.140 8.575 16.490 8.620 ;
        RECT 32.605 8.590 32.950 8.620 ;
        RECT 51.165 8.590 51.510 8.620 ;
        RECT 69.725 8.590 70.070 8.620 ;
        RECT 88.285 8.590 88.630 8.620 ;
        RECT 106.845 8.590 107.190 8.620 ;
        RECT 32.630 8.545 32.950 8.590 ;
        RECT 51.190 8.545 51.510 8.590 ;
        RECT 69.750 8.545 70.070 8.590 ;
        RECT 88.310 8.545 88.630 8.590 ;
        RECT 106.870 8.545 107.190 8.590 ;
        RECT 23.555 5.065 23.875 5.125 ;
        RECT 18.795 4.555 19.115 4.965 ;
        RECT 23.555 4.925 24.625 5.065 ;
        RECT 21.805 4.825 22.905 4.895 ;
        RECT 23.555 4.865 23.875 4.925 ;
        RECT 21.735 4.755 22.985 4.825 ;
        RECT 21.735 4.595 22.025 4.755 ;
        RECT 22.695 4.595 22.985 4.755 ;
        RECT 18.875 3.425 19.035 4.555 ;
        RECT 19.755 4.305 20.075 4.565 ;
        RECT 20.875 4.445 21.195 4.565 ;
        RECT 22.215 4.505 22.505 4.545 ;
        RECT 20.875 4.305 21.705 4.445 ;
        RECT 22.215 4.315 22.545 4.505 ;
        RECT 21.495 4.265 21.705 4.305 ;
        RECT 21.495 4.035 21.785 4.265 ;
        RECT 19.275 3.985 19.595 4.005 ;
        RECT 19.275 3.845 20.225 3.985 ;
        RECT 20.685 3.945 20.975 3.985 ;
        RECT 19.275 3.755 19.825 3.845 ;
        RECT 20.085 3.805 20.225 3.845 ;
        RECT 20.585 3.805 20.975 3.945 ;
        RECT 20.085 3.755 20.975 3.805 ;
        RECT 19.275 3.745 19.595 3.755 ;
        RECT 20.085 3.665 20.725 3.755 ;
        RECT 18.815 3.195 19.105 3.425 ;
        RECT 19.755 3.385 20.075 3.445 ;
        RECT 21.715 3.385 22.035 3.445 ;
        RECT 22.405 3.425 22.545 4.315 ;
        RECT 23.195 4.305 23.515 4.565 ;
        RECT 23.915 4.305 24.235 4.565 ;
        RECT 24.485 4.505 24.625 4.925 ;
        RECT 25.115 4.865 25.435 5.125 ;
        RECT 25.655 5.065 25.945 5.105 ;
        RECT 26.115 5.065 26.435 5.125 ;
        RECT 25.655 4.925 26.435 5.065 ;
        RECT 25.655 4.875 25.945 4.925 ;
        RECT 26.115 4.865 26.435 4.925 ;
        RECT 26.595 4.865 26.915 5.125 ;
        RECT 27.075 4.865 27.395 5.125 ;
        RECT 28.075 4.895 28.395 5.125 ;
        RECT 42.115 5.065 42.435 5.125 ;
        RECT 28.075 4.865 29.505 4.895 ;
        RECT 28.165 4.755 29.505 4.865 ;
        RECT 25.655 4.505 25.945 4.545 ;
        RECT 24.485 4.365 25.945 4.505 ;
        RECT 25.655 4.315 25.945 4.365 ;
        RECT 27.595 4.305 27.915 4.565 ;
        RECT 28.165 4.545 28.305 4.755 ;
        RECT 28.095 4.315 28.385 4.545 ;
        RECT 28.815 4.505 29.105 4.545 ;
        RECT 28.815 4.315 29.145 4.505 ;
        RECT 27.095 4.225 27.385 4.265 ;
        RECT 27.595 4.225 27.825 4.305 ;
        RECT 27.095 4.085 27.825 4.225 ;
        RECT 27.095 4.035 27.385 4.085 ;
        RECT 22.935 3.985 23.255 4.005 ;
        RECT 22.695 3.945 23.255 3.985 ;
        RECT 23.935 3.945 24.225 3.985 ;
        RECT 22.695 3.805 24.225 3.945 ;
        RECT 22.695 3.755 23.255 3.805 ;
        RECT 23.935 3.755 24.225 3.805 ;
        RECT 24.415 3.945 24.705 3.985 ;
        RECT 24.415 3.805 25.345 3.945 ;
        RECT 24.415 3.755 24.705 3.805 ;
        RECT 22.935 3.745 23.255 3.755 ;
        RECT 19.755 3.245 22.035 3.385 ;
        RECT 19.755 3.185 20.075 3.245 ;
        RECT 21.715 3.185 22.035 3.245 ;
        RECT 22.215 3.385 22.545 3.425 ;
        RECT 23.195 3.385 23.515 3.445 ;
        RECT 23.915 3.425 24.235 3.445 ;
        RECT 22.215 3.245 23.515 3.385 ;
        RECT 22.215 3.195 22.505 3.245 ;
        RECT 23.195 3.185 23.515 3.245 ;
        RECT 23.695 3.195 24.235 3.425 ;
        RECT 23.915 3.185 24.235 3.195 ;
        RECT 24.635 3.185 24.955 3.445 ;
        RECT 25.205 3.385 25.345 3.805 ;
        RECT 25.635 3.805 25.955 4.005 ;
        RECT 28.335 3.805 28.625 3.985 ;
        RECT 25.635 3.755 28.625 3.805 ;
        RECT 25.635 3.745 28.545 3.755 ;
        RECT 25.725 3.665 28.545 3.745 ;
        RECT 29.005 3.445 29.145 4.315 ;
        RECT 29.365 4.265 29.505 4.755 ;
        RECT 31.025 4.445 31.365 4.795 ;
        RECT 37.355 4.555 37.675 4.965 ;
        RECT 42.115 4.925 43.185 5.065 ;
        RECT 40.365 4.825 41.465 4.895 ;
        RECT 42.115 4.865 42.435 4.925 ;
        RECT 40.295 4.755 41.545 4.825 ;
        RECT 40.295 4.595 40.585 4.755 ;
        RECT 41.255 4.595 41.545 4.755 ;
        RECT 29.295 4.035 29.585 4.265 ;
        RECT 31.115 3.490 31.285 4.445 ;
        RECT 32.630 3.875 32.950 3.980 ;
        RECT 32.605 3.860 32.950 3.875 ;
        RECT 32.600 3.845 32.950 3.860 ;
        RECT 32.430 3.675 32.950 3.845 ;
        RECT 32.605 3.660 32.950 3.675 ;
        RECT 32.605 3.645 32.895 3.660 ;
        RECT 33.405 3.490 33.755 3.610 ;
        RECT 34.765 3.545 35.055 3.780 ;
        RECT 34.765 3.540 34.995 3.545 ;
        RECT 25.875 3.425 26.195 3.445 ;
        RECT 25.655 3.385 26.195 3.425 ;
        RECT 25.205 3.245 26.195 3.385 ;
        RECT 25.655 3.195 26.195 3.245 ;
        RECT 25.875 3.185 26.195 3.195 ;
        RECT 26.475 3.185 27.155 3.445 ;
        RECT 27.595 3.385 27.915 3.445 ;
        RECT 28.095 3.385 28.385 3.425 ;
        RECT 27.595 3.245 28.385 3.385 ;
        RECT 29.005 3.245 29.355 3.445 ;
        RECT 31.115 3.320 33.755 3.490 ;
        RECT 33.235 3.315 33.755 3.320 ;
        RECT 33.405 3.260 33.755 3.315 ;
        RECT 27.595 3.185 27.915 3.245 ;
        RECT 28.095 3.195 28.385 3.245 ;
        RECT 29.035 3.185 29.355 3.245 ;
        RECT 34.400 3.225 34.630 3.245 ;
        RECT 32.975 3.120 33.265 3.145 ;
        RECT 34.370 3.120 34.660 3.225 ;
        RECT 32.975 2.950 34.660 3.120 ;
        RECT 32.975 2.915 33.265 2.950 ;
        RECT 34.370 2.915 34.660 2.950 ;
        RECT 33.035 2.405 33.205 2.915 ;
        RECT 34.400 2.895 34.630 2.915 ;
        RECT 34.825 2.440 34.995 3.540 ;
        RECT 37.435 3.425 37.595 4.555 ;
        RECT 38.315 4.305 38.635 4.565 ;
        RECT 39.435 4.445 39.755 4.565 ;
        RECT 40.775 4.505 41.065 4.545 ;
        RECT 39.435 4.305 40.265 4.445 ;
        RECT 40.775 4.315 41.105 4.505 ;
        RECT 40.055 4.265 40.265 4.305 ;
        RECT 40.055 4.035 40.345 4.265 ;
        RECT 37.835 3.985 38.155 4.005 ;
        RECT 37.835 3.845 38.785 3.985 ;
        RECT 39.245 3.945 39.535 3.985 ;
        RECT 37.835 3.755 38.385 3.845 ;
        RECT 38.645 3.805 38.785 3.845 ;
        RECT 39.145 3.805 39.535 3.945 ;
        RECT 38.645 3.755 39.535 3.805 ;
        RECT 37.835 3.745 38.155 3.755 ;
        RECT 38.645 3.665 39.285 3.755 ;
        RECT 37.375 3.195 37.665 3.425 ;
        RECT 38.315 3.385 38.635 3.445 ;
        RECT 40.275 3.385 40.595 3.445 ;
        RECT 40.965 3.425 41.105 4.315 ;
        RECT 41.755 4.305 42.075 4.565 ;
        RECT 42.475 4.305 42.795 4.565 ;
        RECT 43.045 4.505 43.185 4.925 ;
        RECT 43.675 4.865 43.995 5.125 ;
        RECT 44.215 5.065 44.505 5.105 ;
        RECT 44.675 5.065 44.995 5.125 ;
        RECT 44.215 4.925 44.995 5.065 ;
        RECT 44.215 4.875 44.505 4.925 ;
        RECT 44.675 4.865 44.995 4.925 ;
        RECT 45.155 4.865 45.475 5.125 ;
        RECT 45.635 4.865 45.955 5.125 ;
        RECT 46.635 4.895 46.955 5.125 ;
        RECT 60.675 5.065 60.995 5.125 ;
        RECT 46.635 4.865 48.065 4.895 ;
        RECT 46.725 4.755 48.065 4.865 ;
        RECT 44.215 4.505 44.505 4.545 ;
        RECT 43.045 4.365 44.505 4.505 ;
        RECT 44.215 4.315 44.505 4.365 ;
        RECT 46.155 4.305 46.475 4.565 ;
        RECT 46.725 4.545 46.865 4.755 ;
        RECT 46.655 4.315 46.945 4.545 ;
        RECT 47.375 4.505 47.665 4.545 ;
        RECT 47.375 4.315 47.705 4.505 ;
        RECT 45.655 4.225 45.945 4.265 ;
        RECT 46.155 4.225 46.385 4.305 ;
        RECT 45.655 4.085 46.385 4.225 ;
        RECT 45.655 4.035 45.945 4.085 ;
        RECT 41.495 3.985 41.815 4.005 ;
        RECT 41.255 3.945 41.815 3.985 ;
        RECT 42.495 3.945 42.785 3.985 ;
        RECT 41.255 3.805 42.785 3.945 ;
        RECT 41.255 3.755 41.815 3.805 ;
        RECT 42.495 3.755 42.785 3.805 ;
        RECT 42.975 3.945 43.265 3.985 ;
        RECT 42.975 3.805 43.905 3.945 ;
        RECT 42.975 3.755 43.265 3.805 ;
        RECT 41.495 3.745 41.815 3.755 ;
        RECT 38.315 3.245 40.595 3.385 ;
        RECT 38.315 3.185 38.635 3.245 ;
        RECT 40.275 3.185 40.595 3.245 ;
        RECT 40.775 3.385 41.105 3.425 ;
        RECT 41.755 3.385 42.075 3.445 ;
        RECT 42.475 3.425 42.795 3.445 ;
        RECT 40.775 3.245 42.075 3.385 ;
        RECT 40.775 3.195 41.065 3.245 ;
        RECT 41.755 3.185 42.075 3.245 ;
        RECT 42.255 3.195 42.795 3.425 ;
        RECT 42.475 3.185 42.795 3.195 ;
        RECT 43.195 3.185 43.515 3.445 ;
        RECT 43.765 3.385 43.905 3.805 ;
        RECT 44.195 3.805 44.515 4.005 ;
        RECT 46.895 3.805 47.185 3.985 ;
        RECT 44.195 3.755 47.185 3.805 ;
        RECT 44.195 3.745 47.105 3.755 ;
        RECT 44.285 3.665 47.105 3.745 ;
        RECT 47.565 3.445 47.705 4.315 ;
        RECT 47.925 4.265 48.065 4.755 ;
        RECT 49.585 4.445 49.925 4.795 ;
        RECT 55.915 4.555 56.235 4.965 ;
        RECT 60.675 4.925 61.745 5.065 ;
        RECT 58.925 4.825 60.025 4.895 ;
        RECT 60.675 4.865 60.995 4.925 ;
        RECT 58.855 4.755 60.105 4.825 ;
        RECT 58.855 4.595 59.145 4.755 ;
        RECT 59.815 4.595 60.105 4.755 ;
        RECT 47.855 4.035 48.145 4.265 ;
        RECT 49.675 3.490 49.845 4.445 ;
        RECT 51.190 3.875 51.510 3.980 ;
        RECT 51.165 3.860 51.510 3.875 ;
        RECT 51.160 3.845 51.510 3.860 ;
        RECT 50.990 3.675 51.510 3.845 ;
        RECT 51.165 3.660 51.510 3.675 ;
        RECT 51.165 3.645 51.455 3.660 ;
        RECT 51.965 3.490 52.315 3.610 ;
        RECT 53.325 3.545 53.615 3.780 ;
        RECT 53.325 3.540 53.555 3.545 ;
        RECT 44.435 3.425 44.755 3.445 ;
        RECT 44.215 3.385 44.755 3.425 ;
        RECT 43.765 3.245 44.755 3.385 ;
        RECT 44.215 3.195 44.755 3.245 ;
        RECT 44.435 3.185 44.755 3.195 ;
        RECT 45.035 3.185 45.715 3.445 ;
        RECT 46.155 3.385 46.475 3.445 ;
        RECT 46.655 3.385 46.945 3.425 ;
        RECT 46.155 3.245 46.945 3.385 ;
        RECT 47.565 3.245 47.915 3.445 ;
        RECT 49.675 3.320 52.315 3.490 ;
        RECT 51.795 3.315 52.315 3.320 ;
        RECT 51.965 3.260 52.315 3.315 ;
        RECT 46.155 3.185 46.475 3.245 ;
        RECT 46.655 3.195 46.945 3.245 ;
        RECT 47.595 3.185 47.915 3.245 ;
        RECT 52.960 3.225 53.190 3.245 ;
        RECT 51.535 3.120 51.825 3.145 ;
        RECT 52.930 3.120 53.220 3.225 ;
        RECT 51.535 2.950 53.220 3.120 ;
        RECT 51.535 2.915 51.825 2.950 ;
        RECT 52.930 2.915 53.220 2.950 ;
        RECT 32.975 2.175 33.265 2.405 ;
        RECT 34.765 2.180 35.060 2.440 ;
        RECT 51.595 2.405 51.765 2.915 ;
        RECT 52.960 2.895 53.190 2.915 ;
        RECT 53.385 2.440 53.555 3.540 ;
        RECT 55.995 3.425 56.155 4.555 ;
        RECT 56.875 4.305 57.195 4.565 ;
        RECT 57.995 4.445 58.315 4.565 ;
        RECT 59.335 4.505 59.625 4.545 ;
        RECT 57.995 4.305 58.825 4.445 ;
        RECT 59.335 4.315 59.665 4.505 ;
        RECT 58.615 4.265 58.825 4.305 ;
        RECT 58.615 4.035 58.905 4.265 ;
        RECT 56.395 3.985 56.715 4.005 ;
        RECT 56.395 3.845 57.345 3.985 ;
        RECT 57.805 3.945 58.095 3.985 ;
        RECT 56.395 3.755 56.945 3.845 ;
        RECT 57.205 3.805 57.345 3.845 ;
        RECT 57.705 3.805 58.095 3.945 ;
        RECT 57.205 3.755 58.095 3.805 ;
        RECT 56.395 3.745 56.715 3.755 ;
        RECT 57.205 3.665 57.845 3.755 ;
        RECT 55.935 3.195 56.225 3.425 ;
        RECT 56.875 3.385 57.195 3.445 ;
        RECT 58.835 3.385 59.155 3.445 ;
        RECT 59.525 3.425 59.665 4.315 ;
        RECT 60.315 4.305 60.635 4.565 ;
        RECT 61.035 4.305 61.355 4.565 ;
        RECT 61.605 4.505 61.745 4.925 ;
        RECT 62.235 4.865 62.555 5.125 ;
        RECT 62.775 5.065 63.065 5.105 ;
        RECT 63.235 5.065 63.555 5.125 ;
        RECT 62.775 4.925 63.555 5.065 ;
        RECT 62.775 4.875 63.065 4.925 ;
        RECT 63.235 4.865 63.555 4.925 ;
        RECT 63.715 4.865 64.035 5.125 ;
        RECT 64.195 4.865 64.515 5.125 ;
        RECT 65.195 4.895 65.515 5.125 ;
        RECT 79.235 5.065 79.555 5.125 ;
        RECT 65.195 4.865 66.625 4.895 ;
        RECT 65.285 4.755 66.625 4.865 ;
        RECT 62.775 4.505 63.065 4.545 ;
        RECT 61.605 4.365 63.065 4.505 ;
        RECT 62.775 4.315 63.065 4.365 ;
        RECT 64.715 4.305 65.035 4.565 ;
        RECT 65.285 4.545 65.425 4.755 ;
        RECT 65.215 4.315 65.505 4.545 ;
        RECT 65.935 4.505 66.225 4.545 ;
        RECT 65.935 4.315 66.265 4.505 ;
        RECT 64.215 4.225 64.505 4.265 ;
        RECT 64.715 4.225 64.945 4.305 ;
        RECT 64.215 4.085 64.945 4.225 ;
        RECT 64.215 4.035 64.505 4.085 ;
        RECT 60.055 3.985 60.375 4.005 ;
        RECT 59.815 3.945 60.375 3.985 ;
        RECT 61.055 3.945 61.345 3.985 ;
        RECT 59.815 3.805 61.345 3.945 ;
        RECT 59.815 3.755 60.375 3.805 ;
        RECT 61.055 3.755 61.345 3.805 ;
        RECT 61.535 3.945 61.825 3.985 ;
        RECT 61.535 3.805 62.465 3.945 ;
        RECT 61.535 3.755 61.825 3.805 ;
        RECT 60.055 3.745 60.375 3.755 ;
        RECT 56.875 3.245 59.155 3.385 ;
        RECT 56.875 3.185 57.195 3.245 ;
        RECT 58.835 3.185 59.155 3.245 ;
        RECT 59.335 3.385 59.665 3.425 ;
        RECT 60.315 3.385 60.635 3.445 ;
        RECT 61.035 3.425 61.355 3.445 ;
        RECT 59.335 3.245 60.635 3.385 ;
        RECT 59.335 3.195 59.625 3.245 ;
        RECT 60.315 3.185 60.635 3.245 ;
        RECT 60.815 3.195 61.355 3.425 ;
        RECT 61.035 3.185 61.355 3.195 ;
        RECT 61.755 3.185 62.075 3.445 ;
        RECT 62.325 3.385 62.465 3.805 ;
        RECT 62.755 3.805 63.075 4.005 ;
        RECT 65.455 3.805 65.745 3.985 ;
        RECT 62.755 3.755 65.745 3.805 ;
        RECT 62.755 3.745 65.665 3.755 ;
        RECT 62.845 3.665 65.665 3.745 ;
        RECT 66.125 3.445 66.265 4.315 ;
        RECT 66.485 4.265 66.625 4.755 ;
        RECT 68.145 4.445 68.485 4.795 ;
        RECT 74.475 4.555 74.795 4.965 ;
        RECT 79.235 4.925 80.305 5.065 ;
        RECT 77.485 4.825 78.585 4.895 ;
        RECT 79.235 4.865 79.555 4.925 ;
        RECT 77.415 4.755 78.665 4.825 ;
        RECT 77.415 4.595 77.705 4.755 ;
        RECT 78.375 4.595 78.665 4.755 ;
        RECT 66.415 4.035 66.705 4.265 ;
        RECT 68.235 3.490 68.405 4.445 ;
        RECT 69.750 3.875 70.070 3.980 ;
        RECT 69.725 3.860 70.070 3.875 ;
        RECT 69.720 3.845 70.070 3.860 ;
        RECT 69.550 3.675 70.070 3.845 ;
        RECT 69.725 3.660 70.070 3.675 ;
        RECT 69.725 3.645 70.015 3.660 ;
        RECT 70.525 3.490 70.875 3.610 ;
        RECT 71.885 3.545 72.175 3.780 ;
        RECT 71.885 3.540 72.115 3.545 ;
        RECT 62.995 3.425 63.315 3.445 ;
        RECT 62.775 3.385 63.315 3.425 ;
        RECT 62.325 3.245 63.315 3.385 ;
        RECT 62.775 3.195 63.315 3.245 ;
        RECT 62.995 3.185 63.315 3.195 ;
        RECT 63.595 3.185 64.275 3.445 ;
        RECT 64.715 3.385 65.035 3.445 ;
        RECT 65.215 3.385 65.505 3.425 ;
        RECT 64.715 3.245 65.505 3.385 ;
        RECT 66.125 3.245 66.475 3.445 ;
        RECT 68.235 3.320 70.875 3.490 ;
        RECT 70.355 3.315 70.875 3.320 ;
        RECT 70.525 3.260 70.875 3.315 ;
        RECT 64.715 3.185 65.035 3.245 ;
        RECT 65.215 3.195 65.505 3.245 ;
        RECT 66.155 3.185 66.475 3.245 ;
        RECT 71.520 3.225 71.750 3.245 ;
        RECT 70.095 3.120 70.385 3.145 ;
        RECT 71.490 3.120 71.780 3.225 ;
        RECT 70.095 2.950 71.780 3.120 ;
        RECT 70.095 2.915 70.385 2.950 ;
        RECT 71.490 2.915 71.780 2.950 ;
        RECT 51.535 2.175 51.825 2.405 ;
        RECT 53.325 2.180 53.620 2.440 ;
        RECT 70.155 2.405 70.325 2.915 ;
        RECT 71.520 2.895 71.750 2.915 ;
        RECT 71.945 2.440 72.115 3.540 ;
        RECT 74.555 3.425 74.715 4.555 ;
        RECT 75.435 4.305 75.755 4.565 ;
        RECT 76.555 4.445 76.875 4.565 ;
        RECT 77.895 4.505 78.185 4.545 ;
        RECT 76.555 4.305 77.385 4.445 ;
        RECT 77.895 4.315 78.225 4.505 ;
        RECT 77.175 4.265 77.385 4.305 ;
        RECT 77.175 4.035 77.465 4.265 ;
        RECT 74.955 3.985 75.275 4.005 ;
        RECT 74.955 3.845 75.905 3.985 ;
        RECT 76.365 3.945 76.655 3.985 ;
        RECT 74.955 3.755 75.505 3.845 ;
        RECT 75.765 3.805 75.905 3.845 ;
        RECT 76.265 3.805 76.655 3.945 ;
        RECT 75.765 3.755 76.655 3.805 ;
        RECT 74.955 3.745 75.275 3.755 ;
        RECT 75.765 3.665 76.405 3.755 ;
        RECT 74.495 3.195 74.785 3.425 ;
        RECT 75.435 3.385 75.755 3.445 ;
        RECT 77.395 3.385 77.715 3.445 ;
        RECT 78.085 3.425 78.225 4.315 ;
        RECT 78.875 4.305 79.195 4.565 ;
        RECT 79.595 4.305 79.915 4.565 ;
        RECT 80.165 4.505 80.305 4.925 ;
        RECT 80.795 4.865 81.115 5.125 ;
        RECT 81.335 5.065 81.625 5.105 ;
        RECT 81.795 5.065 82.115 5.125 ;
        RECT 81.335 4.925 82.115 5.065 ;
        RECT 81.335 4.875 81.625 4.925 ;
        RECT 81.795 4.865 82.115 4.925 ;
        RECT 82.275 4.865 82.595 5.125 ;
        RECT 82.755 4.865 83.075 5.125 ;
        RECT 83.755 4.895 84.075 5.125 ;
        RECT 97.795 5.065 98.115 5.125 ;
        RECT 83.755 4.865 85.185 4.895 ;
        RECT 83.845 4.755 85.185 4.865 ;
        RECT 81.335 4.505 81.625 4.545 ;
        RECT 80.165 4.365 81.625 4.505 ;
        RECT 81.335 4.315 81.625 4.365 ;
        RECT 83.275 4.305 83.595 4.565 ;
        RECT 83.845 4.545 83.985 4.755 ;
        RECT 83.775 4.315 84.065 4.545 ;
        RECT 84.495 4.505 84.785 4.545 ;
        RECT 84.495 4.315 84.825 4.505 ;
        RECT 82.775 4.225 83.065 4.265 ;
        RECT 83.275 4.225 83.505 4.305 ;
        RECT 82.775 4.085 83.505 4.225 ;
        RECT 82.775 4.035 83.065 4.085 ;
        RECT 78.615 3.985 78.935 4.005 ;
        RECT 78.375 3.945 78.935 3.985 ;
        RECT 79.615 3.945 79.905 3.985 ;
        RECT 78.375 3.805 79.905 3.945 ;
        RECT 78.375 3.755 78.935 3.805 ;
        RECT 79.615 3.755 79.905 3.805 ;
        RECT 80.095 3.945 80.385 3.985 ;
        RECT 80.095 3.805 81.025 3.945 ;
        RECT 80.095 3.755 80.385 3.805 ;
        RECT 78.615 3.745 78.935 3.755 ;
        RECT 75.435 3.245 77.715 3.385 ;
        RECT 75.435 3.185 75.755 3.245 ;
        RECT 77.395 3.185 77.715 3.245 ;
        RECT 77.895 3.385 78.225 3.425 ;
        RECT 78.875 3.385 79.195 3.445 ;
        RECT 79.595 3.425 79.915 3.445 ;
        RECT 77.895 3.245 79.195 3.385 ;
        RECT 77.895 3.195 78.185 3.245 ;
        RECT 78.875 3.185 79.195 3.245 ;
        RECT 79.375 3.195 79.915 3.425 ;
        RECT 79.595 3.185 79.915 3.195 ;
        RECT 80.315 3.185 80.635 3.445 ;
        RECT 80.885 3.385 81.025 3.805 ;
        RECT 81.315 3.805 81.635 4.005 ;
        RECT 84.015 3.805 84.305 3.985 ;
        RECT 81.315 3.755 84.305 3.805 ;
        RECT 81.315 3.745 84.225 3.755 ;
        RECT 81.405 3.665 84.225 3.745 ;
        RECT 84.685 3.445 84.825 4.315 ;
        RECT 85.045 4.265 85.185 4.755 ;
        RECT 86.705 4.445 87.045 4.795 ;
        RECT 93.035 4.555 93.355 4.965 ;
        RECT 97.795 4.925 98.865 5.065 ;
        RECT 96.045 4.825 97.145 4.895 ;
        RECT 97.795 4.865 98.115 4.925 ;
        RECT 95.975 4.755 97.225 4.825 ;
        RECT 95.975 4.595 96.265 4.755 ;
        RECT 96.935 4.595 97.225 4.755 ;
        RECT 84.975 4.035 85.265 4.265 ;
        RECT 86.795 3.490 86.965 4.445 ;
        RECT 88.310 3.875 88.630 3.980 ;
        RECT 88.285 3.860 88.630 3.875 ;
        RECT 88.280 3.845 88.630 3.860 ;
        RECT 88.110 3.675 88.630 3.845 ;
        RECT 88.285 3.660 88.630 3.675 ;
        RECT 88.285 3.645 88.575 3.660 ;
        RECT 89.085 3.490 89.435 3.610 ;
        RECT 90.445 3.545 90.735 3.780 ;
        RECT 90.445 3.540 90.675 3.545 ;
        RECT 81.555 3.425 81.875 3.445 ;
        RECT 81.335 3.385 81.875 3.425 ;
        RECT 80.885 3.245 81.875 3.385 ;
        RECT 81.335 3.195 81.875 3.245 ;
        RECT 81.555 3.185 81.875 3.195 ;
        RECT 82.155 3.185 82.835 3.445 ;
        RECT 83.275 3.385 83.595 3.445 ;
        RECT 83.775 3.385 84.065 3.425 ;
        RECT 83.275 3.245 84.065 3.385 ;
        RECT 84.685 3.245 85.035 3.445 ;
        RECT 86.795 3.320 89.435 3.490 ;
        RECT 88.915 3.315 89.435 3.320 ;
        RECT 89.085 3.260 89.435 3.315 ;
        RECT 83.275 3.185 83.595 3.245 ;
        RECT 83.775 3.195 84.065 3.245 ;
        RECT 84.715 3.185 85.035 3.245 ;
        RECT 90.080 3.225 90.310 3.245 ;
        RECT 88.655 3.120 88.945 3.145 ;
        RECT 90.050 3.120 90.340 3.225 ;
        RECT 88.655 2.950 90.340 3.120 ;
        RECT 88.655 2.915 88.945 2.950 ;
        RECT 90.050 2.915 90.340 2.950 ;
        RECT 70.095 2.175 70.385 2.405 ;
        RECT 71.885 2.180 72.180 2.440 ;
        RECT 88.715 2.405 88.885 2.915 ;
        RECT 90.080 2.895 90.310 2.915 ;
        RECT 90.505 2.440 90.675 3.540 ;
        RECT 93.115 3.425 93.275 4.555 ;
        RECT 93.995 4.305 94.315 4.565 ;
        RECT 95.115 4.445 95.435 4.565 ;
        RECT 96.455 4.505 96.745 4.545 ;
        RECT 95.115 4.305 95.945 4.445 ;
        RECT 96.455 4.315 96.785 4.505 ;
        RECT 95.735 4.265 95.945 4.305 ;
        RECT 95.735 4.035 96.025 4.265 ;
        RECT 93.515 3.985 93.835 4.005 ;
        RECT 93.515 3.845 94.465 3.985 ;
        RECT 94.925 3.945 95.215 3.985 ;
        RECT 93.515 3.755 94.065 3.845 ;
        RECT 94.325 3.805 94.465 3.845 ;
        RECT 94.825 3.805 95.215 3.945 ;
        RECT 94.325 3.755 95.215 3.805 ;
        RECT 93.515 3.745 93.835 3.755 ;
        RECT 94.325 3.665 94.965 3.755 ;
        RECT 93.055 3.195 93.345 3.425 ;
        RECT 93.995 3.385 94.315 3.445 ;
        RECT 95.955 3.385 96.275 3.445 ;
        RECT 96.645 3.425 96.785 4.315 ;
        RECT 97.435 4.305 97.755 4.565 ;
        RECT 98.155 4.305 98.475 4.565 ;
        RECT 98.725 4.505 98.865 4.925 ;
        RECT 99.355 4.865 99.675 5.125 ;
        RECT 99.895 5.065 100.185 5.105 ;
        RECT 100.355 5.065 100.675 5.125 ;
        RECT 99.895 4.925 100.675 5.065 ;
        RECT 99.895 4.875 100.185 4.925 ;
        RECT 100.355 4.865 100.675 4.925 ;
        RECT 100.835 4.865 101.155 5.125 ;
        RECT 101.315 4.865 101.635 5.125 ;
        RECT 102.315 4.895 102.635 5.125 ;
        RECT 102.315 4.865 103.745 4.895 ;
        RECT 102.405 4.755 103.745 4.865 ;
        RECT 99.895 4.505 100.185 4.545 ;
        RECT 98.725 4.365 100.185 4.505 ;
        RECT 99.895 4.315 100.185 4.365 ;
        RECT 101.835 4.305 102.155 4.565 ;
        RECT 102.405 4.545 102.545 4.755 ;
        RECT 102.335 4.315 102.625 4.545 ;
        RECT 103.055 4.505 103.345 4.545 ;
        RECT 103.055 4.315 103.385 4.505 ;
        RECT 101.335 4.225 101.625 4.265 ;
        RECT 101.835 4.225 102.065 4.305 ;
        RECT 101.335 4.085 102.065 4.225 ;
        RECT 101.335 4.035 101.625 4.085 ;
        RECT 97.175 3.985 97.495 4.005 ;
        RECT 96.935 3.945 97.495 3.985 ;
        RECT 98.175 3.945 98.465 3.985 ;
        RECT 96.935 3.805 98.465 3.945 ;
        RECT 96.935 3.755 97.495 3.805 ;
        RECT 98.175 3.755 98.465 3.805 ;
        RECT 98.655 3.945 98.945 3.985 ;
        RECT 98.655 3.805 99.585 3.945 ;
        RECT 98.655 3.755 98.945 3.805 ;
        RECT 97.175 3.745 97.495 3.755 ;
        RECT 93.995 3.245 96.275 3.385 ;
        RECT 93.995 3.185 94.315 3.245 ;
        RECT 95.955 3.185 96.275 3.245 ;
        RECT 96.455 3.385 96.785 3.425 ;
        RECT 97.435 3.385 97.755 3.445 ;
        RECT 98.155 3.425 98.475 3.445 ;
        RECT 96.455 3.245 97.755 3.385 ;
        RECT 96.455 3.195 96.745 3.245 ;
        RECT 97.435 3.185 97.755 3.245 ;
        RECT 97.935 3.195 98.475 3.425 ;
        RECT 98.155 3.185 98.475 3.195 ;
        RECT 98.875 3.185 99.195 3.445 ;
        RECT 99.445 3.385 99.585 3.805 ;
        RECT 99.875 3.805 100.195 4.005 ;
        RECT 102.575 3.805 102.865 3.985 ;
        RECT 99.875 3.755 102.865 3.805 ;
        RECT 99.875 3.745 102.785 3.755 ;
        RECT 99.965 3.665 102.785 3.745 ;
        RECT 103.245 3.445 103.385 4.315 ;
        RECT 103.605 4.265 103.745 4.755 ;
        RECT 105.265 4.445 105.605 4.795 ;
        RECT 103.535 4.035 103.825 4.265 ;
        RECT 105.355 3.490 105.525 4.445 ;
        RECT 106.870 3.875 107.190 3.980 ;
        RECT 106.845 3.860 107.190 3.875 ;
        RECT 106.840 3.845 107.190 3.860 ;
        RECT 106.670 3.675 107.190 3.845 ;
        RECT 106.845 3.660 107.190 3.675 ;
        RECT 106.845 3.645 107.135 3.660 ;
        RECT 107.645 3.490 107.995 3.610 ;
        RECT 109.005 3.545 109.295 3.780 ;
        RECT 109.005 3.540 109.235 3.545 ;
        RECT 100.115 3.425 100.435 3.445 ;
        RECT 99.895 3.385 100.435 3.425 ;
        RECT 99.445 3.245 100.435 3.385 ;
        RECT 99.895 3.195 100.435 3.245 ;
        RECT 100.115 3.185 100.435 3.195 ;
        RECT 100.715 3.185 101.395 3.445 ;
        RECT 101.835 3.385 102.155 3.445 ;
        RECT 102.335 3.385 102.625 3.425 ;
        RECT 101.835 3.245 102.625 3.385 ;
        RECT 103.245 3.245 103.595 3.445 ;
        RECT 105.355 3.320 107.995 3.490 ;
        RECT 107.475 3.315 107.995 3.320 ;
        RECT 107.645 3.260 107.995 3.315 ;
        RECT 101.835 3.185 102.155 3.245 ;
        RECT 102.335 3.195 102.625 3.245 ;
        RECT 103.275 3.185 103.595 3.245 ;
        RECT 108.640 3.225 108.870 3.245 ;
        RECT 107.215 3.120 107.505 3.145 ;
        RECT 108.610 3.120 108.900 3.225 ;
        RECT 107.215 2.950 108.900 3.120 ;
        RECT 107.215 2.915 107.505 2.950 ;
        RECT 108.610 2.915 108.900 2.950 ;
        RECT 88.655 2.175 88.945 2.405 ;
        RECT 90.445 2.180 90.740 2.440 ;
        RECT 107.275 2.405 107.445 2.915 ;
        RECT 108.640 2.895 108.870 2.915 ;
        RECT 109.065 2.440 109.235 3.540 ;
        RECT 107.215 2.175 107.505 2.405 ;
        RECT 109.005 2.180 109.300 2.440 ;
      LAYER met2 ;
        RECT 16.235 10.690 110.230 10.860 ;
        RECT 16.235 8.895 16.405 10.690 ;
        RECT 110.060 9.915 110.230 10.690 ;
        RECT 16.545 9.515 16.835 9.640 ;
        RECT 16.545 9.510 16.865 9.515 ;
        RECT 16.545 9.340 17.860 9.510 ;
        RECT 27.320 9.345 27.695 9.715 ;
        RECT 45.880 9.345 46.255 9.715 ;
        RECT 64.440 9.345 64.815 9.715 ;
        RECT 83.000 9.345 83.375 9.715 ;
        RECT 101.560 9.345 101.935 9.715 ;
        RECT 110.030 9.565 110.380 9.915 ;
        RECT 16.545 9.290 16.835 9.340 ;
        RECT 17.690 9.145 17.860 9.340 ;
        RECT 27.995 9.145 28.345 9.245 ;
        RECT 33.430 9.205 33.755 9.270 ;
        RECT 17.690 8.975 28.345 9.145 ;
        RECT 27.995 8.895 28.345 8.975 ;
        RECT 32.315 9.035 33.755 9.205 ;
        RECT 16.170 8.545 16.460 8.895 ;
        RECT 27.150 5.430 31.285 5.620 ;
        RECT 27.150 5.180 27.340 5.430 ;
        RECT 18.815 4.805 19.095 5.180 ;
        RECT 23.585 4.835 23.845 5.155 ;
        RECT 18.825 4.555 19.085 4.805 ;
        RECT 21.255 4.595 21.535 4.620 ;
        RECT 19.785 4.275 20.045 4.595 ;
        RECT 20.905 4.505 21.535 4.595 ;
        RECT 23.225 4.505 23.485 4.595 ;
        RECT 20.905 4.365 23.485 4.505 ;
        RECT 20.905 4.275 21.535 4.365 ;
        RECT 23.225 4.275 23.485 4.365 ;
        RECT 19.295 3.685 19.575 4.060 ;
        RECT 19.845 3.475 19.985 4.275 ;
        RECT 21.255 4.245 21.535 4.275 ;
        RECT 22.695 4.035 22.975 4.060 ;
        RECT 22.695 3.715 23.225 4.035 ;
        RECT 22.695 3.685 22.975 3.715 ;
        RECT 19.785 3.155 20.045 3.475 ;
        RECT 21.745 3.385 22.005 3.475 ;
        RECT 23.225 3.385 23.485 3.475 ;
        RECT 23.645 3.385 23.785 4.835 ;
        RECT 25.135 4.805 25.415 5.180 ;
        RECT 26.145 4.835 26.405 5.155 ;
        RECT 26.625 4.835 26.885 5.155 ;
        RECT 23.935 4.245 24.215 4.620 ;
        RECT 25.205 4.615 25.345 4.805 ;
        RECT 25.015 4.505 25.345 4.615 ;
        RECT 24.725 4.365 25.345 4.505 ;
        RECT 24.005 3.475 24.145 4.245 ;
        RECT 24.725 3.475 24.865 4.365 ;
        RECT 25.015 4.245 25.295 4.365 ;
        RECT 25.665 3.945 25.925 4.035 ;
        RECT 25.085 3.805 25.925 3.945 ;
        RECT 21.745 3.245 22.785 3.385 ;
        RECT 21.745 3.155 22.005 3.245 ;
        RECT 22.645 3.005 22.785 3.245 ;
        RECT 23.225 3.245 23.785 3.385 ;
        RECT 23.225 3.155 23.485 3.245 ;
        RECT 23.945 3.155 24.205 3.475 ;
        RECT 24.665 3.155 24.925 3.475 ;
        RECT 25.085 3.005 25.225 3.805 ;
        RECT 25.665 3.715 25.925 3.805 ;
        RECT 26.205 3.475 26.345 4.835 ;
        RECT 26.625 4.785 26.825 4.835 ;
        RECT 27.095 4.805 27.375 5.180 ;
        RECT 28.095 4.805 28.375 5.180 ;
        RECT 31.095 4.795 31.285 5.430 ;
        RECT 26.565 4.615 26.825 4.785 ;
        RECT 26.565 4.245 27.065 4.615 ;
        RECT 27.625 4.275 27.885 4.595 ;
        RECT 31.025 4.445 31.365 4.795 ;
        RECT 31.115 4.440 31.285 4.445 ;
        RECT 26.565 3.475 26.705 4.245 ;
        RECT 27.685 3.475 27.825 4.275 ;
        RECT 32.315 3.860 32.475 9.035 ;
        RECT 33.430 8.945 33.755 9.035 ;
        RECT 35.810 9.175 36.160 9.295 ;
        RECT 46.555 9.175 46.905 9.250 ;
        RECT 51.990 9.205 52.315 9.270 ;
        RECT 35.810 8.975 46.905 9.175 ;
        RECT 35.810 8.945 36.160 8.975 ;
        RECT 46.555 8.900 46.905 8.975 ;
        RECT 50.875 9.035 52.315 9.205 ;
        RECT 32.630 8.510 32.950 8.835 ;
        RECT 32.660 8.335 32.830 8.510 ;
        RECT 32.660 8.160 32.835 8.335 ;
        RECT 32.660 7.985 33.635 8.160 ;
        RECT 32.630 3.860 32.950 3.980 ;
        RECT 32.315 3.690 32.950 3.860 ;
        RECT 32.630 3.660 32.950 3.690 ;
        RECT 33.460 3.610 33.635 7.985 ;
        RECT 45.710 5.430 49.845 5.620 ;
        RECT 45.710 5.180 45.900 5.430 ;
        RECT 37.375 4.805 37.655 5.180 ;
        RECT 42.145 4.835 42.405 5.155 ;
        RECT 37.385 4.555 37.645 4.805 ;
        RECT 39.815 4.595 40.095 4.620 ;
        RECT 38.345 4.275 38.605 4.595 ;
        RECT 39.465 4.505 40.095 4.595 ;
        RECT 41.785 4.505 42.045 4.595 ;
        RECT 39.465 4.365 42.045 4.505 ;
        RECT 39.465 4.275 40.095 4.365 ;
        RECT 41.785 4.275 42.045 4.365 ;
        RECT 37.855 3.685 38.135 4.060 ;
        RECT 25.905 3.245 26.345 3.475 ;
        RECT 25.905 3.155 26.165 3.245 ;
        RECT 26.505 3.155 26.765 3.475 ;
        RECT 27.625 3.155 27.885 3.475 ;
        RECT 29.055 3.125 29.335 3.500 ;
        RECT 33.405 3.260 33.755 3.610 ;
        RECT 38.405 3.475 38.545 4.275 ;
        RECT 39.815 4.245 40.095 4.275 ;
        RECT 41.255 4.035 41.535 4.060 ;
        RECT 41.255 3.715 41.785 4.035 ;
        RECT 41.255 3.685 41.535 3.715 ;
        RECT 38.345 3.155 38.605 3.475 ;
        RECT 40.305 3.385 40.565 3.475 ;
        RECT 41.785 3.385 42.045 3.475 ;
        RECT 42.205 3.385 42.345 4.835 ;
        RECT 43.695 4.805 43.975 5.180 ;
        RECT 44.705 4.835 44.965 5.155 ;
        RECT 45.185 4.835 45.445 5.155 ;
        RECT 42.495 4.245 42.775 4.620 ;
        RECT 43.765 4.615 43.905 4.805 ;
        RECT 43.575 4.505 43.905 4.615 ;
        RECT 43.285 4.365 43.905 4.505 ;
        RECT 42.565 3.475 42.705 4.245 ;
        RECT 43.285 3.475 43.425 4.365 ;
        RECT 43.575 4.245 43.855 4.365 ;
        RECT 44.225 3.945 44.485 4.035 ;
        RECT 43.645 3.805 44.485 3.945 ;
        RECT 40.305 3.245 41.345 3.385 ;
        RECT 40.305 3.155 40.565 3.245 ;
        RECT 22.645 2.865 25.225 3.005 ;
        RECT 41.205 3.005 41.345 3.245 ;
        RECT 41.785 3.245 42.345 3.385 ;
        RECT 41.785 3.155 42.045 3.245 ;
        RECT 42.505 3.155 42.765 3.475 ;
        RECT 43.225 3.155 43.485 3.475 ;
        RECT 43.645 3.005 43.785 3.805 ;
        RECT 44.225 3.715 44.485 3.805 ;
        RECT 44.765 3.475 44.905 4.835 ;
        RECT 45.185 4.785 45.385 4.835 ;
        RECT 45.655 4.805 45.935 5.180 ;
        RECT 46.655 4.805 46.935 5.180 ;
        RECT 49.655 4.795 49.845 5.430 ;
        RECT 45.125 4.615 45.385 4.785 ;
        RECT 45.125 4.245 45.625 4.615 ;
        RECT 46.185 4.275 46.445 4.595 ;
        RECT 49.585 4.445 49.925 4.795 ;
        RECT 49.675 4.440 49.845 4.445 ;
        RECT 45.125 3.475 45.265 4.245 ;
        RECT 46.245 3.475 46.385 4.275 ;
        RECT 50.875 3.860 51.035 9.035 ;
        RECT 51.990 8.945 52.315 9.035 ;
        RECT 54.370 9.180 54.720 9.300 ;
        RECT 65.110 9.180 65.460 9.255 ;
        RECT 70.550 9.205 70.875 9.270 ;
        RECT 54.370 8.980 65.460 9.180 ;
        RECT 54.370 8.950 54.720 8.980 ;
        RECT 65.110 8.905 65.460 8.980 ;
        RECT 69.435 9.035 70.875 9.205 ;
        RECT 51.190 8.510 51.510 8.835 ;
        RECT 51.220 8.335 51.390 8.510 ;
        RECT 51.220 8.160 51.395 8.335 ;
        RECT 51.220 7.985 52.195 8.160 ;
        RECT 51.190 3.860 51.510 3.980 ;
        RECT 50.875 3.690 51.510 3.860 ;
        RECT 51.190 3.660 51.510 3.690 ;
        RECT 52.020 3.610 52.195 7.985 ;
        RECT 64.270 5.430 68.405 5.620 ;
        RECT 64.270 5.180 64.460 5.430 ;
        RECT 55.935 4.805 56.215 5.180 ;
        RECT 60.705 4.835 60.965 5.155 ;
        RECT 55.945 4.555 56.205 4.805 ;
        RECT 58.375 4.595 58.655 4.620 ;
        RECT 56.905 4.275 57.165 4.595 ;
        RECT 58.025 4.505 58.655 4.595 ;
        RECT 60.345 4.505 60.605 4.595 ;
        RECT 58.025 4.365 60.605 4.505 ;
        RECT 58.025 4.275 58.655 4.365 ;
        RECT 60.345 4.275 60.605 4.365 ;
        RECT 56.415 3.685 56.695 4.060 ;
        RECT 44.465 3.245 44.905 3.475 ;
        RECT 44.465 3.155 44.725 3.245 ;
        RECT 45.065 3.155 45.325 3.475 ;
        RECT 46.185 3.155 46.445 3.475 ;
        RECT 47.615 3.125 47.895 3.500 ;
        RECT 51.965 3.260 52.315 3.610 ;
        RECT 56.965 3.475 57.105 4.275 ;
        RECT 58.375 4.245 58.655 4.275 ;
        RECT 59.815 4.035 60.095 4.060 ;
        RECT 59.815 3.715 60.345 4.035 ;
        RECT 59.815 3.685 60.095 3.715 ;
        RECT 56.905 3.155 57.165 3.475 ;
        RECT 58.865 3.385 59.125 3.475 ;
        RECT 60.345 3.385 60.605 3.475 ;
        RECT 60.765 3.385 60.905 4.835 ;
        RECT 62.255 4.805 62.535 5.180 ;
        RECT 63.265 4.835 63.525 5.155 ;
        RECT 63.745 4.835 64.005 5.155 ;
        RECT 61.055 4.245 61.335 4.620 ;
        RECT 62.325 4.615 62.465 4.805 ;
        RECT 62.135 4.505 62.465 4.615 ;
        RECT 61.845 4.365 62.465 4.505 ;
        RECT 61.125 3.475 61.265 4.245 ;
        RECT 61.845 3.475 61.985 4.365 ;
        RECT 62.135 4.245 62.415 4.365 ;
        RECT 62.785 3.945 63.045 4.035 ;
        RECT 62.205 3.805 63.045 3.945 ;
        RECT 58.865 3.245 59.905 3.385 ;
        RECT 58.865 3.155 59.125 3.245 ;
        RECT 41.205 2.865 43.785 3.005 ;
        RECT 59.765 3.005 59.905 3.245 ;
        RECT 60.345 3.245 60.905 3.385 ;
        RECT 60.345 3.155 60.605 3.245 ;
        RECT 61.065 3.155 61.325 3.475 ;
        RECT 61.785 3.155 62.045 3.475 ;
        RECT 62.205 3.005 62.345 3.805 ;
        RECT 62.785 3.715 63.045 3.805 ;
        RECT 63.325 3.475 63.465 4.835 ;
        RECT 63.745 4.785 63.945 4.835 ;
        RECT 64.215 4.805 64.495 5.180 ;
        RECT 65.215 4.805 65.495 5.180 ;
        RECT 68.215 4.795 68.405 5.430 ;
        RECT 63.685 4.615 63.945 4.785 ;
        RECT 63.685 4.245 64.185 4.615 ;
        RECT 64.745 4.275 65.005 4.595 ;
        RECT 68.145 4.445 68.485 4.795 ;
        RECT 68.235 4.440 68.405 4.445 ;
        RECT 63.685 3.475 63.825 4.245 ;
        RECT 64.805 3.475 64.945 4.275 ;
        RECT 69.435 3.860 69.595 9.035 ;
        RECT 70.550 8.945 70.875 9.035 ;
        RECT 72.885 9.175 73.235 9.295 ;
        RECT 83.670 9.175 84.020 9.250 ;
        RECT 89.110 9.205 89.435 9.270 ;
        RECT 72.885 8.975 84.020 9.175 ;
        RECT 72.885 8.945 73.235 8.975 ;
        RECT 83.670 8.900 84.020 8.975 ;
        RECT 87.995 9.035 89.435 9.205 ;
        RECT 69.750 8.510 70.070 8.835 ;
        RECT 69.780 8.335 69.950 8.510 ;
        RECT 69.780 8.160 69.955 8.335 ;
        RECT 69.780 7.985 70.755 8.160 ;
        RECT 69.750 3.860 70.070 3.980 ;
        RECT 69.435 3.690 70.070 3.860 ;
        RECT 69.750 3.660 70.070 3.690 ;
        RECT 70.580 3.610 70.755 7.985 ;
        RECT 82.830 5.430 86.965 5.620 ;
        RECT 82.830 5.180 83.020 5.430 ;
        RECT 74.495 4.805 74.775 5.180 ;
        RECT 79.265 4.835 79.525 5.155 ;
        RECT 74.505 4.555 74.765 4.805 ;
        RECT 76.935 4.595 77.215 4.620 ;
        RECT 75.465 4.275 75.725 4.595 ;
        RECT 76.585 4.505 77.215 4.595 ;
        RECT 78.905 4.505 79.165 4.595 ;
        RECT 76.585 4.365 79.165 4.505 ;
        RECT 76.585 4.275 77.215 4.365 ;
        RECT 78.905 4.275 79.165 4.365 ;
        RECT 74.975 3.685 75.255 4.060 ;
        RECT 63.025 3.245 63.465 3.475 ;
        RECT 63.025 3.155 63.285 3.245 ;
        RECT 63.625 3.155 63.885 3.475 ;
        RECT 64.745 3.155 65.005 3.475 ;
        RECT 66.175 3.125 66.455 3.500 ;
        RECT 70.525 3.260 70.875 3.610 ;
        RECT 75.525 3.475 75.665 4.275 ;
        RECT 76.935 4.245 77.215 4.275 ;
        RECT 78.375 4.035 78.655 4.060 ;
        RECT 78.375 3.715 78.905 4.035 ;
        RECT 78.375 3.685 78.655 3.715 ;
        RECT 75.465 3.155 75.725 3.475 ;
        RECT 77.425 3.385 77.685 3.475 ;
        RECT 78.905 3.385 79.165 3.475 ;
        RECT 79.325 3.385 79.465 4.835 ;
        RECT 80.815 4.805 81.095 5.180 ;
        RECT 81.825 4.835 82.085 5.155 ;
        RECT 82.305 4.835 82.565 5.155 ;
        RECT 79.615 4.245 79.895 4.620 ;
        RECT 80.885 4.615 81.025 4.805 ;
        RECT 80.695 4.505 81.025 4.615 ;
        RECT 80.405 4.365 81.025 4.505 ;
        RECT 79.685 3.475 79.825 4.245 ;
        RECT 80.405 3.475 80.545 4.365 ;
        RECT 80.695 4.245 80.975 4.365 ;
        RECT 81.345 3.945 81.605 4.035 ;
        RECT 80.765 3.805 81.605 3.945 ;
        RECT 77.425 3.245 78.465 3.385 ;
        RECT 77.425 3.155 77.685 3.245 ;
        RECT 59.765 2.865 62.345 3.005 ;
        RECT 78.325 3.005 78.465 3.245 ;
        RECT 78.905 3.245 79.465 3.385 ;
        RECT 78.905 3.155 79.165 3.245 ;
        RECT 79.625 3.155 79.885 3.475 ;
        RECT 80.345 3.155 80.605 3.475 ;
        RECT 80.765 3.005 80.905 3.805 ;
        RECT 81.345 3.715 81.605 3.805 ;
        RECT 81.885 3.475 82.025 4.835 ;
        RECT 82.305 4.785 82.505 4.835 ;
        RECT 82.775 4.805 83.055 5.180 ;
        RECT 83.775 4.805 84.055 5.180 ;
        RECT 86.775 4.795 86.965 5.430 ;
        RECT 82.245 4.615 82.505 4.785 ;
        RECT 82.245 4.245 82.745 4.615 ;
        RECT 83.305 4.275 83.565 4.595 ;
        RECT 86.705 4.445 87.045 4.795 ;
        RECT 86.795 4.440 86.965 4.445 ;
        RECT 82.245 3.475 82.385 4.245 ;
        RECT 83.365 3.475 83.505 4.275 ;
        RECT 87.995 3.860 88.155 9.035 ;
        RECT 89.110 8.945 89.435 9.035 ;
        RECT 91.445 9.175 91.795 9.295 ;
        RECT 102.230 9.175 102.580 9.250 ;
        RECT 107.670 9.205 107.995 9.270 ;
        RECT 91.445 8.975 102.580 9.175 ;
        RECT 91.445 8.945 91.795 8.975 ;
        RECT 102.230 8.900 102.580 8.975 ;
        RECT 106.555 9.035 107.995 9.205 ;
        RECT 88.310 8.510 88.630 8.835 ;
        RECT 88.340 8.335 88.510 8.510 ;
        RECT 88.340 8.160 88.515 8.335 ;
        RECT 88.340 7.985 89.315 8.160 ;
        RECT 88.310 3.860 88.630 3.980 ;
        RECT 87.995 3.690 88.630 3.860 ;
        RECT 88.310 3.660 88.630 3.690 ;
        RECT 89.140 3.610 89.315 7.985 ;
        RECT 101.390 5.430 105.525 5.620 ;
        RECT 101.390 5.180 101.580 5.430 ;
        RECT 93.055 4.805 93.335 5.180 ;
        RECT 97.825 4.835 98.085 5.155 ;
        RECT 93.065 4.555 93.325 4.805 ;
        RECT 95.495 4.595 95.775 4.620 ;
        RECT 94.025 4.275 94.285 4.595 ;
        RECT 95.145 4.505 95.775 4.595 ;
        RECT 97.465 4.505 97.725 4.595 ;
        RECT 95.145 4.365 97.725 4.505 ;
        RECT 95.145 4.275 95.775 4.365 ;
        RECT 97.465 4.275 97.725 4.365 ;
        RECT 93.535 3.685 93.815 4.060 ;
        RECT 81.585 3.245 82.025 3.475 ;
        RECT 81.585 3.155 81.845 3.245 ;
        RECT 82.185 3.155 82.445 3.475 ;
        RECT 83.305 3.155 83.565 3.475 ;
        RECT 84.735 3.125 85.015 3.500 ;
        RECT 89.085 3.260 89.435 3.610 ;
        RECT 94.085 3.475 94.225 4.275 ;
        RECT 95.495 4.245 95.775 4.275 ;
        RECT 96.935 4.035 97.215 4.060 ;
        RECT 96.935 3.715 97.465 4.035 ;
        RECT 96.935 3.685 97.215 3.715 ;
        RECT 94.025 3.155 94.285 3.475 ;
        RECT 95.985 3.385 96.245 3.475 ;
        RECT 97.465 3.385 97.725 3.475 ;
        RECT 97.885 3.385 98.025 4.835 ;
        RECT 99.375 4.805 99.655 5.180 ;
        RECT 100.385 4.835 100.645 5.155 ;
        RECT 100.865 4.835 101.125 5.155 ;
        RECT 98.175 4.245 98.455 4.620 ;
        RECT 99.445 4.615 99.585 4.805 ;
        RECT 99.255 4.505 99.585 4.615 ;
        RECT 98.965 4.365 99.585 4.505 ;
        RECT 98.245 3.475 98.385 4.245 ;
        RECT 98.965 3.475 99.105 4.365 ;
        RECT 99.255 4.245 99.535 4.365 ;
        RECT 99.905 3.945 100.165 4.035 ;
        RECT 99.325 3.805 100.165 3.945 ;
        RECT 95.985 3.245 97.025 3.385 ;
        RECT 95.985 3.155 96.245 3.245 ;
        RECT 78.325 2.865 80.905 3.005 ;
        RECT 96.885 3.005 97.025 3.245 ;
        RECT 97.465 3.245 98.025 3.385 ;
        RECT 97.465 3.155 97.725 3.245 ;
        RECT 98.185 3.155 98.445 3.475 ;
        RECT 98.905 3.155 99.165 3.475 ;
        RECT 99.325 3.005 99.465 3.805 ;
        RECT 99.905 3.715 100.165 3.805 ;
        RECT 100.445 3.475 100.585 4.835 ;
        RECT 100.865 4.785 101.065 4.835 ;
        RECT 101.335 4.805 101.615 5.180 ;
        RECT 102.335 4.805 102.615 5.180 ;
        RECT 105.335 4.795 105.525 5.430 ;
        RECT 100.805 4.615 101.065 4.785 ;
        RECT 100.805 4.245 101.305 4.615 ;
        RECT 101.865 4.275 102.125 4.595 ;
        RECT 105.265 4.445 105.605 4.795 ;
        RECT 105.355 4.440 105.525 4.445 ;
        RECT 100.805 3.475 100.945 4.245 ;
        RECT 101.925 3.475 102.065 4.275 ;
        RECT 106.555 3.860 106.715 9.035 ;
        RECT 107.670 8.945 107.995 9.035 ;
        RECT 106.870 8.510 107.190 8.835 ;
        RECT 106.900 8.335 107.070 8.510 ;
        RECT 106.900 8.160 107.075 8.335 ;
        RECT 106.900 7.985 107.875 8.160 ;
        RECT 106.870 3.860 107.190 3.980 ;
        RECT 106.555 3.690 107.190 3.860 ;
        RECT 106.870 3.660 107.190 3.690 ;
        RECT 107.700 3.610 107.875 7.985 ;
        RECT 100.145 3.245 100.585 3.475 ;
        RECT 100.145 3.155 100.405 3.245 ;
        RECT 100.745 3.155 101.005 3.475 ;
        RECT 101.865 3.155 102.125 3.475 ;
        RECT 103.295 3.125 103.575 3.500 ;
        RECT 107.645 3.260 107.995 3.610 ;
        RECT 96.885 2.865 99.465 3.005 ;
      LAYER met3 ;
        RECT 27.320 9.685 27.695 9.715 ;
        RECT 45.880 9.685 46.255 9.715 ;
        RECT 64.440 9.685 64.815 9.715 ;
        RECT 83.000 9.685 83.375 9.715 ;
        RECT 101.560 9.685 101.935 9.715 ;
        RECT 27.320 9.385 28.325 9.685 ;
        RECT 27.320 9.345 27.695 9.385 ;
        RECT 28.025 6.995 28.325 9.385 ;
        RECT 45.880 9.385 46.885 9.685 ;
        RECT 45.880 9.345 46.255 9.385 ;
        RECT 46.585 6.995 46.885 9.385 ;
        RECT 64.440 9.385 65.445 9.685 ;
        RECT 64.440 9.345 64.815 9.385 ;
        RECT 65.145 6.995 65.445 9.385 ;
        RECT 83.000 9.385 84.005 9.685 ;
        RECT 83.000 9.345 83.375 9.385 ;
        RECT 83.705 6.995 84.005 9.385 ;
        RECT 101.560 9.385 102.565 9.685 ;
        RECT 101.560 9.345 101.935 9.385 ;
        RECT 102.265 6.995 102.565 9.385 ;
        RECT 18.190 5.925 28.325 6.995 ;
        RECT 36.750 5.925 46.885 6.995 ;
        RECT 55.310 5.925 65.445 6.995 ;
        RECT 73.870 5.925 84.005 6.995 ;
        RECT 92.430 5.925 102.565 6.995 ;
        RECT 17.800 5.700 28.325 5.925 ;
        RECT 36.360 5.700 46.885 5.925 ;
        RECT 54.920 5.700 65.445 5.925 ;
        RECT 73.480 5.700 84.005 5.925 ;
        RECT 92.040 5.700 102.565 5.925 ;
        RECT 17.800 5.435 18.640 5.700 ;
        RECT 18.190 4.015 18.490 5.435 ;
        RECT 18.790 5.155 19.120 5.160 ;
        RECT 18.790 4.825 19.525 5.155 ;
        RECT 18.790 4.820 19.115 4.825 ;
        RECT 21.265 4.600 21.565 5.700 ;
        RECT 21.230 4.595 21.565 4.600 ;
        RECT 21.230 4.265 21.965 4.595 ;
        RECT 21.230 4.260 21.560 4.265 ;
        RECT 22.700 4.040 23.000 5.700 ;
        RECT 36.360 5.435 37.200 5.700 ;
        RECT 28.075 5.160 28.395 5.180 ;
        RECT 25.110 5.155 25.445 5.160 ;
        RECT 27.075 5.155 27.400 5.160 ;
        RECT 28.075 5.155 28.400 5.160 ;
        RECT 25.110 4.825 25.845 5.155 ;
        RECT 26.815 4.825 27.545 5.155 ;
        RECT 27.845 4.825 28.405 5.155 ;
        RECT 25.110 4.820 25.445 4.825 ;
        RECT 27.075 4.820 27.400 4.825 ;
        RECT 23.910 4.595 24.235 4.600 ;
        RECT 23.910 4.260 24.465 4.595 ;
        RECT 19.125 4.035 19.645 4.040 ;
        RECT 22.670 4.035 23.000 4.040 ;
        RECT 19.125 4.015 19.855 4.035 ;
        RECT 18.190 3.715 19.855 4.015 ;
        RECT 19.125 3.705 19.855 3.715 ;
        RECT 22.670 3.705 23.405 4.035 ;
        RECT 22.670 3.700 22.995 3.705 ;
        RECT 24.165 3.465 24.465 4.260 ;
        RECT 27.845 3.465 28.145 4.825 ;
        RECT 36.750 4.015 37.050 5.435 ;
        RECT 37.350 5.155 37.680 5.160 ;
        RECT 37.350 4.825 38.085 5.155 ;
        RECT 37.350 4.820 37.675 4.825 ;
        RECT 39.825 4.600 40.125 5.700 ;
        RECT 39.790 4.595 40.125 4.600 ;
        RECT 39.790 4.265 40.525 4.595 ;
        RECT 39.790 4.260 40.120 4.265 ;
        RECT 41.260 4.040 41.560 5.700 ;
        RECT 54.920 5.435 55.760 5.700 ;
        RECT 46.635 5.160 46.955 5.180 ;
        RECT 43.670 5.155 44.005 5.160 ;
        RECT 45.635 5.155 45.960 5.160 ;
        RECT 46.635 5.155 46.960 5.160 ;
        RECT 43.670 4.825 44.405 5.155 ;
        RECT 45.375 4.825 46.105 5.155 ;
        RECT 46.405 4.825 46.965 5.155 ;
        RECT 43.670 4.820 44.005 4.825 ;
        RECT 45.635 4.820 45.960 4.825 ;
        RECT 42.470 4.595 42.795 4.600 ;
        RECT 42.470 4.260 43.025 4.595 ;
        RECT 37.685 4.035 38.205 4.040 ;
        RECT 41.230 4.035 41.560 4.040 ;
        RECT 37.685 4.015 38.415 4.035 ;
        RECT 36.750 3.715 38.415 4.015 ;
        RECT 37.685 3.705 38.415 3.715 ;
        RECT 41.230 3.705 41.965 4.035 ;
        RECT 41.230 3.700 41.555 3.705 ;
        RECT 24.165 3.165 28.145 3.465 ;
        RECT 29.030 3.475 29.355 3.500 ;
        RECT 29.030 3.145 29.765 3.475 ;
        RECT 42.725 3.465 43.025 4.260 ;
        RECT 46.405 3.465 46.705 4.825 ;
        RECT 55.310 4.015 55.610 5.435 ;
        RECT 55.910 5.155 56.240 5.160 ;
        RECT 55.910 4.825 56.645 5.155 ;
        RECT 55.910 4.820 56.235 4.825 ;
        RECT 58.385 4.600 58.685 5.700 ;
        RECT 58.350 4.595 58.685 4.600 ;
        RECT 58.350 4.265 59.085 4.595 ;
        RECT 58.350 4.260 58.680 4.265 ;
        RECT 59.820 4.040 60.120 5.700 ;
        RECT 73.480 5.435 74.320 5.700 ;
        RECT 65.195 5.160 65.515 5.180 ;
        RECT 62.230 5.155 62.565 5.160 ;
        RECT 64.195 5.155 64.520 5.160 ;
        RECT 65.195 5.155 65.520 5.160 ;
        RECT 62.230 4.825 62.965 5.155 ;
        RECT 63.935 4.825 64.665 5.155 ;
        RECT 64.965 4.825 65.525 5.155 ;
        RECT 62.230 4.820 62.565 4.825 ;
        RECT 64.195 4.820 64.520 4.825 ;
        RECT 61.030 4.595 61.355 4.600 ;
        RECT 61.030 4.260 61.585 4.595 ;
        RECT 56.245 4.035 56.765 4.040 ;
        RECT 59.790 4.035 60.120 4.040 ;
        RECT 56.245 4.015 56.975 4.035 ;
        RECT 55.310 3.715 56.975 4.015 ;
        RECT 56.245 3.705 56.975 3.715 ;
        RECT 59.790 3.705 60.525 4.035 ;
        RECT 59.790 3.700 60.115 3.705 ;
        RECT 42.725 3.165 46.705 3.465 ;
        RECT 47.590 3.475 47.915 3.500 ;
        RECT 47.590 3.145 48.325 3.475 ;
        RECT 61.285 3.465 61.585 4.260 ;
        RECT 64.965 3.465 65.265 4.825 ;
        RECT 73.870 4.015 74.170 5.435 ;
        RECT 74.470 5.155 74.800 5.160 ;
        RECT 74.470 4.825 75.205 5.155 ;
        RECT 74.470 4.820 74.795 4.825 ;
        RECT 76.945 4.600 77.245 5.700 ;
        RECT 76.910 4.595 77.245 4.600 ;
        RECT 76.910 4.265 77.645 4.595 ;
        RECT 76.910 4.260 77.240 4.265 ;
        RECT 78.380 4.040 78.680 5.700 ;
        RECT 92.040 5.435 92.880 5.700 ;
        RECT 83.755 5.160 84.075 5.180 ;
        RECT 80.790 5.155 81.125 5.160 ;
        RECT 82.755 5.155 83.080 5.160 ;
        RECT 83.755 5.155 84.080 5.160 ;
        RECT 80.790 4.825 81.525 5.155 ;
        RECT 82.495 4.825 83.225 5.155 ;
        RECT 83.525 4.825 84.085 5.155 ;
        RECT 80.790 4.820 81.125 4.825 ;
        RECT 82.755 4.820 83.080 4.825 ;
        RECT 79.590 4.595 79.915 4.600 ;
        RECT 79.590 4.260 80.145 4.595 ;
        RECT 74.805 4.035 75.325 4.040 ;
        RECT 78.350 4.035 78.680 4.040 ;
        RECT 74.805 4.015 75.535 4.035 ;
        RECT 73.870 3.715 75.535 4.015 ;
        RECT 74.805 3.705 75.535 3.715 ;
        RECT 78.350 3.705 79.085 4.035 ;
        RECT 78.350 3.700 78.675 3.705 ;
        RECT 61.285 3.165 65.265 3.465 ;
        RECT 66.150 3.475 66.475 3.500 ;
        RECT 66.150 3.145 66.885 3.475 ;
        RECT 79.845 3.465 80.145 4.260 ;
        RECT 83.525 3.465 83.825 4.825 ;
        RECT 92.430 4.015 92.730 5.435 ;
        RECT 93.030 5.155 93.360 5.160 ;
        RECT 93.030 4.825 93.765 5.155 ;
        RECT 93.030 4.820 93.355 4.825 ;
        RECT 95.505 4.600 95.805 5.700 ;
        RECT 95.470 4.595 95.805 4.600 ;
        RECT 95.470 4.265 96.205 4.595 ;
        RECT 95.470 4.260 95.800 4.265 ;
        RECT 96.940 4.040 97.240 5.700 ;
        RECT 102.315 5.160 102.635 5.180 ;
        RECT 99.350 5.155 99.685 5.160 ;
        RECT 101.315 5.155 101.640 5.160 ;
        RECT 102.315 5.155 102.640 5.160 ;
        RECT 99.350 4.825 100.085 5.155 ;
        RECT 101.055 4.825 101.785 5.155 ;
        RECT 102.085 4.825 102.645 5.155 ;
        RECT 99.350 4.820 99.685 4.825 ;
        RECT 101.315 4.820 101.640 4.825 ;
        RECT 98.150 4.595 98.475 4.600 ;
        RECT 98.150 4.260 98.705 4.595 ;
        RECT 93.365 4.035 93.885 4.040 ;
        RECT 96.910 4.035 97.240 4.040 ;
        RECT 93.365 4.015 94.095 4.035 ;
        RECT 92.430 3.715 94.095 4.015 ;
        RECT 93.365 3.705 94.095 3.715 ;
        RECT 96.910 3.705 97.645 4.035 ;
        RECT 96.910 3.700 97.235 3.705 ;
        RECT 79.845 3.165 83.825 3.465 ;
        RECT 84.710 3.475 85.035 3.500 ;
        RECT 84.710 3.145 85.445 3.475 ;
        RECT 98.405 3.465 98.705 4.260 ;
        RECT 102.085 3.465 102.385 4.825 ;
        RECT 98.405 3.165 102.385 3.465 ;
        RECT 103.270 3.475 103.595 3.500 ;
        RECT 103.270 3.145 104.005 3.475 ;
        RECT 29.030 3.140 29.355 3.145 ;
        RECT 47.590 3.140 47.915 3.145 ;
        RECT 66.150 3.140 66.475 3.145 ;
        RECT 84.710 3.140 85.035 3.145 ;
        RECT 103.270 3.140 103.595 3.145 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r1
MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r2
  CLASS BLOCK ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 101.085 BY 12.470 ;
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 18.825 8.225 18.995 9.495 ;
        RECT 30.050 8.230 30.220 9.500 ;
        RECT 30.050 2.960 30.220 4.230 ;
      LAYER met1 ;
        RECT 18.740 8.395 19.080 8.455 ;
        RECT 18.740 8.365 19.225 8.395 ;
        RECT 21.050 8.365 21.390 8.455 ;
        RECT 18.740 8.195 21.390 8.365 ;
        RECT 18.740 8.175 19.080 8.195 ;
        RECT 21.050 8.175 21.390 8.195 ;
        RECT 29.980 8.400 30.305 8.475 ;
        RECT 29.980 8.230 30.450 8.400 ;
        RECT 29.980 8.150 30.305 8.230 ;
        RECT 29.975 4.930 30.300 5.255 ;
        RECT 30.050 4.260 30.230 4.930 ;
        RECT 29.990 4.230 30.280 4.260 ;
        RECT 29.990 4.060 30.450 4.230 ;
        RECT 29.990 4.030 30.280 4.060 ;
      LAYER met2 ;
        RECT 21.135 9.300 30.220 9.470 ;
        RECT 18.770 8.130 19.050 8.500 ;
        RECT 21.135 8.485 21.305 9.300 ;
        RECT 21.080 8.145 21.360 8.485 ;
        RECT 30.045 8.475 30.220 9.300 ;
        RECT 29.980 8.150 30.305 8.475 ;
        RECT 30.045 5.255 30.220 8.150 ;
        RECT 29.975 4.930 30.300 5.255 ;
      LAYER met3 ;
        RECT 18.740 8.130 19.080 12.460 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 35.410 8.225 35.580 9.495 ;
        RECT 46.635 8.230 46.805 9.500 ;
        RECT 46.635 2.960 46.805 4.230 ;
      LAYER met1 ;
        RECT 35.325 8.395 35.665 8.455 ;
        RECT 35.325 8.365 35.810 8.395 ;
        RECT 37.635 8.365 37.975 8.455 ;
        RECT 35.325 8.195 37.975 8.365 ;
        RECT 35.325 8.175 35.665 8.195 ;
        RECT 37.635 8.175 37.975 8.195 ;
        RECT 46.565 8.400 46.890 8.475 ;
        RECT 46.565 8.230 47.035 8.400 ;
        RECT 46.565 8.150 46.890 8.230 ;
        RECT 46.560 4.930 46.885 5.255 ;
        RECT 46.635 4.260 46.815 4.930 ;
        RECT 46.575 4.230 46.865 4.260 ;
        RECT 46.575 4.060 47.035 4.230 ;
        RECT 46.575 4.030 46.865 4.060 ;
      LAYER met2 ;
        RECT 37.720 9.300 46.805 9.470 ;
        RECT 35.355 8.130 35.635 8.500 ;
        RECT 37.720 8.485 37.890 9.300 ;
        RECT 37.665 8.145 37.945 8.485 ;
        RECT 46.630 8.475 46.805 9.300 ;
        RECT 46.565 8.150 46.890 8.475 ;
        RECT 46.630 5.255 46.805 8.150 ;
        RECT 46.560 4.930 46.885 5.255 ;
      LAYER met3 ;
        RECT 35.325 8.130 35.665 12.460 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 51.995 8.230 52.165 9.500 ;
        RECT 63.220 8.235 63.390 9.505 ;
        RECT 63.220 2.965 63.390 4.235 ;
      LAYER met1 ;
        RECT 51.910 8.400 52.250 8.460 ;
        RECT 51.910 8.370 52.395 8.400 ;
        RECT 54.220 8.370 54.560 8.460 ;
        RECT 51.910 8.200 54.560 8.370 ;
        RECT 51.910 8.180 52.250 8.200 ;
        RECT 54.220 8.180 54.560 8.200 ;
        RECT 63.150 8.405 63.475 8.480 ;
        RECT 63.150 8.235 63.620 8.405 ;
        RECT 63.150 8.155 63.475 8.235 ;
        RECT 63.145 4.935 63.470 5.260 ;
        RECT 63.220 4.265 63.400 4.935 ;
        RECT 63.160 4.235 63.450 4.265 ;
        RECT 63.160 4.065 63.620 4.235 ;
        RECT 63.160 4.035 63.450 4.065 ;
      LAYER met2 ;
        RECT 54.305 9.305 63.390 9.475 ;
        RECT 51.940 8.135 52.220 8.505 ;
        RECT 54.305 8.490 54.475 9.305 ;
        RECT 54.250 8.150 54.530 8.490 ;
        RECT 63.215 8.480 63.390 9.305 ;
        RECT 63.150 8.155 63.475 8.480 ;
        RECT 63.215 5.260 63.390 8.155 ;
        RECT 63.145 4.935 63.470 5.260 ;
      LAYER met3 ;
        RECT 51.910 8.135 52.250 12.465 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 68.580 8.235 68.750 9.505 ;
        RECT 79.805 8.240 79.975 9.510 ;
        RECT 79.805 2.970 79.975 4.240 ;
      LAYER met1 ;
        RECT 68.495 8.405 68.835 8.465 ;
        RECT 68.495 8.375 68.980 8.405 ;
        RECT 70.805 8.375 71.145 8.465 ;
        RECT 68.495 8.205 71.145 8.375 ;
        RECT 68.495 8.185 68.835 8.205 ;
        RECT 70.805 8.185 71.145 8.205 ;
        RECT 79.735 8.410 80.060 8.485 ;
        RECT 79.735 8.240 80.205 8.410 ;
        RECT 79.735 8.160 80.060 8.240 ;
        RECT 79.730 4.940 80.055 5.265 ;
        RECT 79.805 4.270 79.985 4.940 ;
        RECT 79.745 4.240 80.035 4.270 ;
        RECT 79.745 4.070 80.205 4.240 ;
        RECT 79.745 4.040 80.035 4.070 ;
      LAYER met2 ;
        RECT 70.890 9.310 79.975 9.480 ;
        RECT 68.525 8.140 68.805 8.510 ;
        RECT 70.890 8.495 71.060 9.310 ;
        RECT 70.835 8.155 71.115 8.495 ;
        RECT 79.800 8.485 79.975 9.310 ;
        RECT 79.735 8.160 80.060 8.485 ;
        RECT 79.800 5.265 79.975 8.160 ;
        RECT 79.730 4.940 80.055 5.265 ;
      LAYER met3 ;
        RECT 68.495 8.140 68.835 12.470 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 85.160 8.235 85.330 9.505 ;
        RECT 96.385 8.240 96.555 9.510 ;
        RECT 96.385 2.970 96.555 4.240 ;
      LAYER met1 ;
        RECT 85.075 8.405 85.415 8.465 ;
        RECT 85.075 8.375 85.560 8.405 ;
        RECT 87.385 8.375 87.725 8.465 ;
        RECT 85.075 8.205 87.725 8.375 ;
        RECT 85.075 8.185 85.415 8.205 ;
        RECT 87.385 8.185 87.725 8.205 ;
        RECT 96.315 8.410 96.640 8.485 ;
        RECT 96.315 8.240 96.785 8.410 ;
        RECT 96.315 8.160 96.640 8.240 ;
        RECT 96.310 4.940 96.635 5.265 ;
        RECT 96.385 4.270 96.565 4.940 ;
        RECT 96.325 4.240 96.615 4.270 ;
        RECT 96.325 4.070 96.785 4.240 ;
        RECT 96.325 4.040 96.615 4.070 ;
      LAYER met2 ;
        RECT 87.470 9.310 96.555 9.480 ;
        RECT 85.105 8.140 85.385 8.510 ;
        RECT 87.470 8.495 87.640 9.310 ;
        RECT 87.415 8.155 87.695 8.495 ;
        RECT 96.380 8.485 96.555 9.310 ;
        RECT 96.315 8.160 96.640 8.485 ;
        RECT 96.380 5.265 96.555 8.160 ;
        RECT 96.310 4.940 96.635 5.265 ;
      LAYER met3 ;
        RECT 85.075 8.140 85.415 12.470 ;
    END
  END s5
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 100.540 4.025 100.715 5.170 ;
        RECT 100.540 3.590 100.710 4.025 ;
        RECT 100.545 1.880 100.715 2.390 ;
      LAYER met1 ;
        RECT 100.480 3.555 100.770 3.790 ;
        RECT 100.480 3.550 100.710 3.555 ;
        RECT 100.540 2.450 100.710 3.550 ;
        RECT 100.480 2.190 100.775 2.450 ;
    END
  END X5_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 83.960 4.025 84.135 5.170 ;
        RECT 83.960 3.590 84.130 4.025 ;
        RECT 83.965 1.880 84.135 2.390 ;
      LAYER met1 ;
        RECT 83.900 3.555 84.190 3.790 ;
        RECT 83.900 3.550 84.130 3.555 ;
        RECT 83.960 2.450 84.130 3.550 ;
        RECT 83.900 2.190 84.195 2.450 ;
    END
  END X4_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 67.375 4.020 67.550 5.165 ;
        RECT 67.375 3.585 67.545 4.020 ;
        RECT 67.380 1.875 67.550 2.385 ;
      LAYER met1 ;
        RECT 67.315 3.550 67.605 3.785 ;
        RECT 67.315 3.545 67.545 3.550 ;
        RECT 67.375 2.445 67.545 3.545 ;
        RECT 67.315 2.185 67.610 2.445 ;
    END
  END X3_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 50.790 4.015 50.965 5.160 ;
        RECT 50.790 3.580 50.960 4.015 ;
        RECT 50.795 1.870 50.965 2.380 ;
      LAYER met1 ;
        RECT 50.730 3.545 51.020 3.780 ;
        RECT 50.730 3.540 50.960 3.545 ;
        RECT 50.790 2.440 50.960 3.540 ;
        RECT 50.730 2.180 51.025 2.440 ;
    END
  END X2_Y1
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 34.205 4.015 34.380 5.160 ;
        RECT 34.205 3.580 34.375 4.015 ;
        RECT 34.210 1.870 34.380 2.380 ;
      LAYER met1 ;
        RECT 34.145 3.545 34.435 3.780 ;
        RECT 34.145 3.540 34.375 3.545 ;
        RECT 34.205 2.440 34.375 3.540 ;
        RECT 34.145 2.180 34.440 2.440 ;
    END
  END X1_Y1
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 15.595 8.225 15.765 9.495 ;
      LAYER met1 ;
        RECT 15.540 8.425 15.830 8.430 ;
        RECT 15.535 8.395 15.830 8.425 ;
        RECT 15.535 8.225 15.995 8.395 ;
        RECT 15.535 8.200 15.830 8.225 ;
        RECT 15.535 8.195 15.825 8.200 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 67.750 8.745 71.425 8.750 ;
        RECT 51.180 8.740 54.840 8.745 ;
        RECT 15.205 8.130 21.670 8.740 ;
        RECT 28.895 8.130 38.255 8.740 ;
        RECT 45.480 8.135 54.840 8.740 ;
        RECT 62.065 8.140 71.425 8.745 ;
        RECT 78.650 8.140 88.005 8.750 ;
        RECT 15.205 7.135 21.690 8.130 ;
        RECT 28.895 7.135 38.275 8.130 ;
        RECT 45.480 7.140 54.860 8.135 ;
        RECT 62.065 7.145 71.445 8.140 ;
        RECT 78.650 7.145 88.025 8.140 ;
        RECT 95.230 7.145 101.085 8.750 ;
        RECT 62.065 7.140 101.085 7.145 ;
        RECT 45.480 7.135 101.085 7.140 ;
        RECT 15.205 4.705 101.085 7.135 ;
        RECT 15.210 4.315 101.085 4.705 ;
        RECT 15.210 4.310 71.115 4.315 ;
        RECT 15.210 4.305 54.530 4.310 ;
        RECT 15.210 4.225 21.670 4.305 ;
        RECT 15.210 3.715 21.360 4.225 ;
        RECT 29.055 3.720 37.945 4.305 ;
        RECT 45.640 3.720 54.530 4.305 ;
        RECT 62.225 3.725 71.115 4.310 ;
        RECT 78.810 3.730 87.695 4.315 ;
        RECT 95.390 3.730 101.085 4.315 ;
        RECT 67.915 3.720 71.115 3.725 ;
        RECT 84.495 3.720 87.695 3.730 ;
        RECT 18.160 3.710 21.360 3.715 ;
        RECT 34.745 3.710 37.945 3.720 ;
        RECT 51.330 3.715 54.530 3.720 ;
      LAYER li1 ;
        RECT 17.400 10.035 17.575 10.585 ;
        RECT 17.400 8.435 17.570 10.035 ;
        RECT 15.585 7.025 15.755 7.755 ;
        RECT 17.400 7.295 17.575 8.435 ;
        RECT 17.400 7.025 17.570 7.295 ;
        RECT 18.815 7.025 18.985 7.755 ;
        RECT 30.040 7.040 30.210 7.760 ;
        RECT 32.785 7.040 32.955 7.760 ;
        RECT 33.775 7.040 33.945 7.760 ;
        RECT 28.810 7.030 34.750 7.040 ;
        RECT 35.400 7.030 35.570 7.755 ;
        RECT 46.625 7.040 46.795 7.760 ;
        RECT 49.370 7.040 49.540 7.760 ;
        RECT 50.360 7.040 50.530 7.760 ;
        RECT 45.395 7.030 51.335 7.040 ;
        RECT 51.985 7.030 52.155 7.760 ;
        RECT 63.210 7.045 63.380 7.765 ;
        RECT 65.955 7.045 66.125 7.765 ;
        RECT 66.945 7.045 67.115 7.765 ;
        RECT 61.980 7.035 67.920 7.045 ;
        RECT 68.570 7.035 68.740 7.765 ;
        RECT 79.795 7.050 79.965 7.770 ;
        RECT 82.540 7.050 82.710 7.770 ;
        RECT 83.530 7.050 83.700 7.770 ;
        RECT 78.565 7.035 84.505 7.050 ;
        RECT 85.150 7.035 85.320 7.765 ;
        RECT 96.375 7.050 96.545 7.770 ;
        RECT 99.120 7.050 99.290 7.770 ;
        RECT 100.110 7.050 100.280 7.770 ;
        RECT 61.980 7.030 71.495 7.035 ;
        RECT 78.565 7.030 88.075 7.035 ;
        RECT 0.000 5.805 21.965 7.025 ;
        RECT 23.070 5.805 23.400 6.525 ;
        RECT 24.085 5.805 24.365 6.265 ;
        RECT 25.230 5.805 25.500 6.585 ;
        RECT 26.050 5.805 26.420 6.185 ;
        RECT 28.810 5.965 38.575 7.030 ;
        RECT 28.680 5.805 38.575 5.965 ;
        RECT 39.655 5.805 39.985 6.525 ;
        RECT 40.670 5.805 40.950 6.265 ;
        RECT 41.815 5.805 42.085 6.585 ;
        RECT 42.635 5.805 43.005 6.185 ;
        RECT 45.395 5.965 55.160 7.030 ;
        RECT 45.265 5.810 55.160 5.965 ;
        RECT 56.240 5.810 56.570 6.530 ;
        RECT 57.255 5.810 57.535 6.270 ;
        RECT 58.400 5.810 58.670 6.590 ;
        RECT 59.220 5.810 59.590 6.190 ;
        RECT 61.980 5.970 71.745 7.030 ;
        RECT 61.850 5.815 71.745 5.970 ;
        RECT 72.825 5.815 73.155 6.535 ;
        RECT 73.840 5.815 74.120 6.275 ;
        RECT 74.985 5.815 75.255 6.595 ;
        RECT 75.805 5.815 76.175 6.195 ;
        RECT 78.565 5.975 88.330 7.030 ;
        RECT 78.435 5.815 88.330 5.975 ;
        RECT 89.405 5.815 89.735 6.535 ;
        RECT 90.420 5.815 90.700 6.275 ;
        RECT 91.565 5.815 91.835 6.595 ;
        RECT 92.385 5.815 92.755 6.195 ;
        RECT 95.145 5.975 101.085 7.050 ;
        RECT 95.015 5.815 101.085 5.975 ;
        RECT 61.850 5.810 101.085 5.815 ;
        RECT 45.265 5.805 101.085 5.810 ;
        RECT 0.000 5.645 101.085 5.805 ;
        RECT 0.000 5.640 71.745 5.645 ;
        RECT 0.000 5.635 55.160 5.640 ;
        RECT 0.000 5.425 21.965 5.635 ;
        RECT 21.655 5.125 21.915 5.425 ;
        RECT 22.880 5.135 23.500 5.635 ;
        RECT 23.300 4.955 23.500 5.135 ;
        RECT 24.310 5.095 24.530 5.635 ;
        RECT 25.180 4.985 25.790 5.635 ;
        RECT 26.610 5.095 26.870 5.635 ;
        RECT 28.350 5.430 38.575 5.635 ;
        RECT 25.610 4.955 25.800 4.985 ;
        RECT 23.300 4.765 23.630 4.955 ;
        RECT 25.610 4.715 25.940 4.955 ;
        RECT 28.350 4.495 28.680 5.430 ;
        RECT 30.040 4.700 30.210 5.430 ;
        RECT 32.785 4.700 32.955 5.430 ;
        RECT 33.775 4.700 33.945 5.430 ;
        RECT 34.750 5.425 38.500 5.430 ;
        RECT 38.240 5.125 38.500 5.425 ;
        RECT 39.465 5.135 40.085 5.635 ;
        RECT 39.885 4.955 40.085 5.135 ;
        RECT 40.895 5.095 41.115 5.635 ;
        RECT 41.765 4.985 42.375 5.635 ;
        RECT 43.195 5.095 43.455 5.635 ;
        RECT 44.935 5.430 55.160 5.635 ;
        RECT 42.195 4.955 42.385 4.985 ;
        RECT 39.885 4.765 40.215 4.955 ;
        RECT 42.195 4.715 42.525 4.955 ;
        RECT 44.935 4.495 45.265 5.430 ;
        RECT 46.625 4.700 46.795 5.430 ;
        RECT 49.370 4.700 49.540 5.430 ;
        RECT 50.360 4.700 50.530 5.430 ;
        RECT 54.825 5.130 55.085 5.430 ;
        RECT 56.050 5.140 56.670 5.640 ;
        RECT 56.470 4.960 56.670 5.140 ;
        RECT 57.480 5.100 57.700 5.640 ;
        RECT 58.350 4.990 58.960 5.640 ;
        RECT 59.780 5.100 60.040 5.640 ;
        RECT 61.520 5.430 71.745 5.640 ;
        RECT 58.780 4.960 58.970 4.990 ;
        RECT 56.470 4.770 56.800 4.960 ;
        RECT 58.780 4.720 59.110 4.960 ;
        RECT 61.520 4.500 61.850 5.430 ;
        RECT 63.210 4.705 63.380 5.430 ;
        RECT 65.955 4.705 66.125 5.430 ;
        RECT 66.945 4.705 67.115 5.430 ;
        RECT 71.410 5.135 71.670 5.430 ;
        RECT 72.635 5.145 73.255 5.645 ;
        RECT 73.055 4.965 73.255 5.145 ;
        RECT 74.065 5.105 74.285 5.645 ;
        RECT 74.935 4.995 75.545 5.645 ;
        RECT 76.365 5.105 76.625 5.645 ;
        RECT 78.105 5.430 88.330 5.645 ;
        RECT 75.365 4.965 75.555 4.995 ;
        RECT 73.055 4.775 73.385 4.965 ;
        RECT 75.365 4.725 75.695 4.965 ;
        RECT 78.105 4.505 78.435 5.430 ;
        RECT 79.795 4.710 79.965 5.430 ;
        RECT 82.540 4.710 82.710 5.430 ;
        RECT 83.530 4.710 83.700 5.430 ;
        RECT 87.990 5.135 88.250 5.430 ;
        RECT 89.215 5.145 89.835 5.645 ;
        RECT 89.635 4.965 89.835 5.145 ;
        RECT 90.645 5.105 90.865 5.645 ;
        RECT 91.515 4.995 92.125 5.645 ;
        RECT 92.945 5.105 93.205 5.645 ;
        RECT 94.685 5.430 101.085 5.645 ;
        RECT 91.945 4.965 92.135 4.995 ;
        RECT 89.635 4.775 89.965 4.965 ;
        RECT 91.945 4.725 92.275 4.965 ;
        RECT 94.685 4.505 95.015 5.430 ;
        RECT 96.375 4.710 96.545 5.430 ;
        RECT 99.120 4.710 99.290 5.430 ;
        RECT 100.110 4.710 100.280 5.430 ;
      LAYER met1 ;
        RECT 17.340 9.135 17.630 9.165 ;
        RECT 17.170 8.965 17.630 9.135 ;
        RECT 17.340 8.935 17.630 8.965 ;
        RECT 28.810 7.030 34.750 7.040 ;
        RECT 45.395 7.030 51.335 7.040 ;
        RECT 61.980 7.035 67.920 7.045 ;
        RECT 78.565 7.035 84.505 7.050 ;
        RECT 61.980 7.030 71.495 7.035 ;
        RECT 78.565 7.030 88.075 7.035 ;
        RECT 0.000 5.965 21.965 7.025 ;
        RECT 23.490 5.965 23.640 5.970 ;
        RECT 28.810 5.965 38.575 7.030 ;
        RECT 45.395 5.970 55.160 7.030 ;
        RECT 61.980 5.975 71.745 7.030 ;
        RECT 73.245 5.975 73.395 5.980 ;
        RECT 78.565 5.975 88.330 7.030 ;
        RECT 89.825 5.975 89.975 5.980 ;
        RECT 95.145 5.975 101.085 7.050 ;
        RECT 56.660 5.970 56.810 5.975 ;
        RECT 61.980 5.970 101.085 5.975 ;
        RECT 40.075 5.965 40.225 5.970 ;
        RECT 45.395 5.965 101.085 5.970 ;
        RECT 0.000 5.495 101.085 5.965 ;
        RECT 0.000 5.490 71.745 5.495 ;
        RECT 0.000 5.485 55.160 5.490 ;
        RECT 0.000 5.425 21.965 5.485 ;
        RECT 28.680 5.445 38.575 5.485 ;
        RECT 45.265 5.445 55.160 5.485 ;
        RECT 61.850 5.450 71.745 5.490 ;
        RECT 78.435 5.455 88.330 5.495 ;
        RECT 95.015 5.455 101.085 5.495 ;
        RECT 28.685 5.430 38.575 5.445 ;
        RECT 45.270 5.430 55.160 5.445 ;
        RECT 61.855 5.435 71.745 5.450 ;
        RECT 78.440 5.440 88.330 5.455 ;
        RECT 95.020 5.440 101.085 5.455 ;
        RECT 61.980 5.430 71.745 5.435 ;
        RECT 78.565 5.430 88.330 5.440 ;
        RECT 95.145 5.430 101.085 5.440 ;
        RECT 34.750 5.425 38.475 5.430 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 67.920 12.465 101.085 12.470 ;
        RECT 51.335 12.460 101.085 12.465 ;
        RECT 0.000 10.860 101.085 12.460 ;
        RECT 15.415 10.855 18.165 10.860 ;
        RECT 18.645 10.855 22.170 10.860 ;
        RECT 15.585 10.225 15.755 10.855 ;
        RECT 18.815 10.225 18.985 10.855 ;
        RECT 19.770 10.305 19.940 10.585 ;
        RECT 19.770 10.135 20.000 10.305 ;
        RECT 19.830 8.525 20.000 10.135 ;
        RECT 21.880 8.525 22.170 10.855 ;
        RECT 22.450 8.525 22.730 10.860 ;
        RECT 23.010 8.525 23.290 10.860 ;
        RECT 23.570 8.525 23.850 10.860 ;
        RECT 24.130 8.525 24.410 10.860 ;
        RECT 24.690 8.525 24.970 10.860 ;
        RECT 25.250 8.525 25.530 10.860 ;
        RECT 25.810 8.525 26.090 10.860 ;
        RECT 26.370 8.525 26.650 10.860 ;
        RECT 26.930 8.525 27.210 10.860 ;
        RECT 27.490 8.525 27.770 10.860 ;
        RECT 28.050 8.525 28.330 10.860 ;
        RECT 28.610 8.525 28.785 10.860 ;
        RECT 30.040 10.230 30.210 10.860 ;
        RECT 32.785 10.230 32.955 10.860 ;
        RECT 33.775 10.230 33.945 10.860 ;
        RECT 35.230 10.855 38.755 10.860 ;
        RECT 35.400 10.225 35.570 10.855 ;
        RECT 36.355 10.305 36.525 10.585 ;
        RECT 36.355 10.135 36.585 10.305 ;
        RECT 36.415 8.525 36.585 10.135 ;
        RECT 38.465 8.525 38.755 10.855 ;
        RECT 39.035 8.525 39.315 10.860 ;
        RECT 39.595 8.525 39.875 10.860 ;
        RECT 40.155 8.525 40.435 10.860 ;
        RECT 40.715 8.525 40.995 10.860 ;
        RECT 41.275 8.525 41.555 10.860 ;
        RECT 41.835 8.525 42.115 10.860 ;
        RECT 42.395 8.525 42.675 10.860 ;
        RECT 42.955 8.525 43.235 10.860 ;
        RECT 43.515 8.525 43.795 10.860 ;
        RECT 44.075 8.525 44.355 10.860 ;
        RECT 44.635 8.525 44.915 10.860 ;
        RECT 45.195 8.525 45.370 10.860 ;
        RECT 46.625 10.230 46.795 10.860 ;
        RECT 49.370 10.230 49.540 10.860 ;
        RECT 50.360 10.230 50.530 10.860 ;
        RECT 51.985 10.230 52.155 10.860 ;
        RECT 52.940 10.310 53.110 10.590 ;
        RECT 52.940 10.140 53.170 10.310 ;
        RECT 53.000 8.530 53.170 10.140 ;
        RECT 55.050 8.530 55.340 10.860 ;
        RECT 55.620 8.530 55.900 10.860 ;
        RECT 56.180 8.530 56.460 10.860 ;
        RECT 56.740 8.530 57.020 10.860 ;
        RECT 57.300 8.530 57.580 10.860 ;
        RECT 57.860 8.530 58.140 10.860 ;
        RECT 58.420 8.530 58.700 10.860 ;
        RECT 58.980 8.530 59.260 10.860 ;
        RECT 59.540 8.530 59.820 10.860 ;
        RECT 60.100 8.530 60.380 10.860 ;
        RECT 60.660 8.530 60.940 10.860 ;
        RECT 61.220 8.530 61.500 10.860 ;
        RECT 61.780 8.530 61.955 10.860 ;
        RECT 63.210 10.235 63.380 10.860 ;
        RECT 65.955 10.235 66.125 10.860 ;
        RECT 66.945 10.235 67.115 10.860 ;
        RECT 68.570 10.235 68.740 10.860 ;
        RECT 69.525 10.315 69.695 10.595 ;
        RECT 69.525 10.145 69.755 10.315 ;
        RECT 69.585 8.535 69.755 10.145 ;
        RECT 71.635 8.535 71.925 10.860 ;
        RECT 72.205 8.535 72.485 10.860 ;
        RECT 72.765 8.535 73.045 10.860 ;
        RECT 73.325 8.535 73.605 10.860 ;
        RECT 73.885 8.535 74.165 10.860 ;
        RECT 74.445 8.535 74.725 10.860 ;
        RECT 75.005 8.535 75.285 10.860 ;
        RECT 75.565 8.535 75.845 10.860 ;
        RECT 76.125 8.535 76.405 10.860 ;
        RECT 76.685 8.535 76.965 10.860 ;
        RECT 77.245 8.535 77.525 10.860 ;
        RECT 77.805 8.535 78.085 10.860 ;
        RECT 78.365 8.535 78.540 10.860 ;
        RECT 79.795 10.240 79.965 10.860 ;
        RECT 82.540 10.240 82.710 10.860 ;
        RECT 83.530 10.240 83.700 10.860 ;
        RECT 85.150 10.235 85.320 10.860 ;
        RECT 86.105 10.315 86.275 10.595 ;
        RECT 86.105 10.145 86.335 10.315 ;
        RECT 86.165 8.535 86.335 10.145 ;
        RECT 88.215 8.535 88.505 10.860 ;
        RECT 88.785 8.535 89.065 10.860 ;
        RECT 89.345 8.535 89.625 10.860 ;
        RECT 89.905 8.535 90.185 10.860 ;
        RECT 90.465 8.535 90.745 10.860 ;
        RECT 91.025 8.535 91.305 10.860 ;
        RECT 91.585 8.535 91.865 10.860 ;
        RECT 92.145 8.535 92.425 10.860 ;
        RECT 92.705 8.535 92.985 10.860 ;
        RECT 93.265 8.535 93.545 10.860 ;
        RECT 93.825 8.535 94.105 10.860 ;
        RECT 94.385 8.535 94.665 10.860 ;
        RECT 94.945 8.535 95.120 10.860 ;
        RECT 96.375 10.240 96.545 10.860 ;
        RECT 99.120 10.240 99.290 10.860 ;
        RECT 100.110 10.240 100.280 10.860 ;
        RECT 19.770 8.355 20.000 8.525 ;
        RECT 21.740 8.355 28.785 8.525 ;
        RECT 36.355 8.355 36.585 8.525 ;
        RECT 38.325 8.355 45.370 8.525 ;
        RECT 52.940 8.360 53.170 8.530 ;
        RECT 54.910 8.360 61.955 8.530 ;
        RECT 69.525 8.365 69.755 8.535 ;
        RECT 71.495 8.365 78.540 8.535 ;
        RECT 86.105 8.365 86.335 8.535 ;
        RECT 88.075 8.365 95.120 8.535 ;
        RECT 19.770 7.295 19.940 8.355 ;
        RECT 23.150 7.895 23.400 8.355 ;
        RECT 25.220 7.955 25.550 8.355 ;
        RECT 27.310 7.845 27.760 8.355 ;
        RECT 23.300 7.115 23.640 7.365 ;
        RECT 25.520 7.115 25.850 7.445 ;
        RECT 36.355 7.295 36.525 8.355 ;
        RECT 39.735 7.895 39.985 8.355 ;
        RECT 41.805 7.955 42.135 8.355 ;
        RECT 43.895 7.845 44.345 8.355 ;
        RECT 39.885 7.115 40.225 7.365 ;
        RECT 42.105 7.115 42.435 7.445 ;
        RECT 52.940 7.300 53.110 8.360 ;
        RECT 56.320 7.900 56.570 8.360 ;
        RECT 58.390 7.960 58.720 8.360 ;
        RECT 60.480 7.850 60.930 8.360 ;
        RECT 56.470 7.120 56.810 7.370 ;
        RECT 58.690 7.120 59.020 7.450 ;
        RECT 69.525 7.305 69.695 8.365 ;
        RECT 72.905 7.905 73.155 8.365 ;
        RECT 74.975 7.965 75.305 8.365 ;
        RECT 77.065 7.855 77.515 8.365 ;
        RECT 73.055 7.125 73.395 7.375 ;
        RECT 75.275 7.125 75.605 7.455 ;
        RECT 86.105 7.305 86.275 8.365 ;
        RECT 89.485 7.905 89.735 8.365 ;
        RECT 91.555 7.965 91.885 8.365 ;
        RECT 93.645 7.855 94.095 8.365 ;
        RECT 89.635 7.125 89.975 7.375 ;
        RECT 91.855 7.125 92.185 7.455 ;
      LAYER met1 ;
        RECT 67.920 12.465 101.085 12.470 ;
        RECT 51.335 12.460 101.085 12.465 ;
        RECT 0.000 10.860 101.085 12.460 ;
        RECT 15.415 10.855 18.165 10.860 ;
        RECT 18.645 10.855 22.170 10.860 ;
        RECT 19.605 10.850 19.780 10.855 ;
        RECT 19.605 8.805 19.775 10.850 ;
        RECT 19.605 8.775 20.060 8.805 ;
        RECT 19.595 8.605 20.060 8.775 ;
        RECT 21.880 8.685 22.170 10.855 ;
        RECT 22.450 8.685 22.730 10.860 ;
        RECT 23.010 8.685 23.290 10.860 ;
        RECT 23.570 8.685 23.850 10.860 ;
        RECT 24.130 8.685 24.410 10.860 ;
        RECT 24.690 8.685 24.970 10.860 ;
        RECT 25.250 8.685 25.530 10.860 ;
        RECT 25.810 8.685 26.090 10.860 ;
        RECT 26.370 8.685 26.650 10.860 ;
        RECT 26.930 8.685 27.210 10.860 ;
        RECT 27.490 8.685 27.770 10.860 ;
        RECT 28.050 8.685 28.330 10.860 ;
        RECT 28.610 8.685 28.785 10.860 ;
        RECT 35.230 10.855 38.755 10.860 ;
        RECT 36.190 10.850 36.365 10.855 ;
        RECT 36.190 8.805 36.360 10.850 ;
        RECT 36.190 8.775 36.645 8.805 ;
        RECT 19.605 8.600 20.060 8.605 ;
        RECT 19.770 8.575 20.060 8.600 ;
        RECT 21.740 8.325 28.785 8.685 ;
        RECT 36.180 8.605 36.645 8.775 ;
        RECT 38.465 8.685 38.755 10.855 ;
        RECT 39.035 8.685 39.315 10.860 ;
        RECT 39.595 8.685 39.875 10.860 ;
        RECT 40.155 8.685 40.435 10.860 ;
        RECT 40.715 8.685 40.995 10.860 ;
        RECT 41.275 8.685 41.555 10.860 ;
        RECT 41.835 8.685 42.115 10.860 ;
        RECT 42.395 8.685 42.675 10.860 ;
        RECT 42.955 8.685 43.235 10.860 ;
        RECT 43.515 8.685 43.795 10.860 ;
        RECT 44.075 8.685 44.355 10.860 ;
        RECT 44.635 8.685 44.915 10.860 ;
        RECT 45.195 8.685 45.370 10.860 ;
        RECT 52.775 10.855 52.950 10.860 ;
        RECT 52.775 8.810 52.945 10.855 ;
        RECT 52.775 8.780 53.230 8.810 ;
        RECT 36.190 8.600 36.645 8.605 ;
        RECT 36.355 8.575 36.645 8.600 ;
        RECT 38.325 8.325 45.370 8.685 ;
        RECT 52.765 8.610 53.230 8.780 ;
        RECT 55.050 8.690 55.340 10.860 ;
        RECT 55.620 8.690 55.900 10.860 ;
        RECT 56.180 8.690 56.460 10.860 ;
        RECT 56.740 8.690 57.020 10.860 ;
        RECT 57.300 8.690 57.580 10.860 ;
        RECT 57.860 8.690 58.140 10.860 ;
        RECT 58.420 8.690 58.700 10.860 ;
        RECT 58.980 8.690 59.260 10.860 ;
        RECT 59.540 8.690 59.820 10.860 ;
        RECT 60.100 8.690 60.380 10.860 ;
        RECT 60.660 8.690 60.940 10.860 ;
        RECT 61.220 8.690 61.500 10.860 ;
        RECT 61.780 8.690 61.955 10.860 ;
        RECT 69.360 8.815 69.530 10.860 ;
        RECT 69.360 8.785 69.815 8.815 ;
        RECT 52.775 8.605 53.230 8.610 ;
        RECT 52.940 8.580 53.230 8.605 ;
        RECT 54.910 8.330 61.955 8.690 ;
        RECT 69.350 8.615 69.815 8.785 ;
        RECT 71.635 8.695 71.925 10.860 ;
        RECT 72.205 8.695 72.485 10.860 ;
        RECT 72.765 8.695 73.045 10.860 ;
        RECT 73.325 8.695 73.605 10.860 ;
        RECT 73.885 8.695 74.165 10.860 ;
        RECT 74.445 8.695 74.725 10.860 ;
        RECT 75.005 8.695 75.285 10.860 ;
        RECT 75.565 8.695 75.845 10.860 ;
        RECT 76.125 8.695 76.405 10.860 ;
        RECT 76.685 8.695 76.965 10.860 ;
        RECT 77.245 8.695 77.525 10.860 ;
        RECT 77.805 8.695 78.085 10.860 ;
        RECT 78.365 8.695 78.540 10.860 ;
        RECT 85.940 8.815 86.110 10.860 ;
        RECT 85.940 8.785 86.395 8.815 ;
        RECT 69.360 8.610 69.815 8.615 ;
        RECT 69.525 8.585 69.815 8.610 ;
        RECT 71.495 8.335 78.540 8.695 ;
        RECT 85.930 8.615 86.395 8.785 ;
        RECT 88.215 8.695 88.505 10.860 ;
        RECT 88.785 8.695 89.065 10.860 ;
        RECT 89.345 8.695 89.625 10.860 ;
        RECT 89.905 8.695 90.185 10.860 ;
        RECT 90.465 8.695 90.745 10.860 ;
        RECT 91.025 8.695 91.305 10.860 ;
        RECT 91.585 8.695 91.865 10.860 ;
        RECT 92.145 8.695 92.425 10.860 ;
        RECT 92.705 8.695 92.985 10.860 ;
        RECT 93.265 8.695 93.545 10.860 ;
        RECT 93.825 8.695 94.105 10.860 ;
        RECT 94.385 8.695 94.665 10.860 ;
        RECT 94.945 8.695 95.120 10.860 ;
        RECT 85.940 8.610 86.395 8.615 ;
        RECT 86.105 8.585 86.395 8.610 ;
        RECT 88.075 8.335 95.120 8.695 ;
        RECT 24.305 8.045 24.565 8.325 ;
        RECT 40.890 8.045 41.150 8.325 ;
        RECT 57.475 8.050 57.735 8.330 ;
        RECT 74.060 8.055 74.320 8.335 ;
        RECT 90.640 8.055 90.900 8.335 ;
        RECT 24.270 7.945 24.700 8.045 ;
        RECT 40.855 7.945 41.285 8.045 ;
        RECT 57.440 7.950 57.870 8.050 ;
        RECT 74.025 7.955 74.455 8.055 ;
        RECT 90.605 7.955 91.035 8.055 ;
        RECT 23.340 7.805 25.690 7.945 ;
        RECT 23.340 7.365 23.480 7.805 ;
        RECT 24.280 7.775 24.560 7.805 ;
        RECT 24.300 7.745 24.560 7.775 ;
        RECT 25.550 7.365 25.690 7.805 ;
        RECT 39.925 7.805 42.275 7.945 ;
        RECT 39.925 7.365 40.065 7.805 ;
        RECT 40.865 7.775 41.145 7.805 ;
        RECT 40.885 7.745 41.145 7.775 ;
        RECT 42.135 7.365 42.275 7.805 ;
        RECT 56.510 7.810 58.860 7.950 ;
        RECT 56.510 7.370 56.650 7.810 ;
        RECT 57.450 7.780 57.730 7.810 ;
        RECT 57.470 7.750 57.730 7.780 ;
        RECT 58.720 7.370 58.860 7.810 ;
        RECT 73.095 7.815 75.445 7.955 ;
        RECT 73.095 7.375 73.235 7.815 ;
        RECT 74.035 7.785 74.315 7.815 ;
        RECT 74.055 7.755 74.315 7.785 ;
        RECT 75.305 7.375 75.445 7.815 ;
        RECT 89.675 7.815 92.025 7.955 ;
        RECT 89.675 7.375 89.815 7.815 ;
        RECT 90.615 7.785 90.895 7.815 ;
        RECT 90.635 7.755 90.895 7.785 ;
        RECT 91.885 7.375 92.025 7.815 ;
        RECT 23.260 7.135 23.550 7.365 ;
        RECT 25.470 7.135 25.760 7.365 ;
        RECT 39.845 7.135 40.135 7.365 ;
        RECT 42.055 7.135 42.345 7.365 ;
        RECT 56.430 7.140 56.720 7.370 ;
        RECT 58.640 7.140 58.930 7.370 ;
        RECT 73.015 7.145 73.305 7.375 ;
        RECT 75.225 7.145 75.515 7.375 ;
        RECT 89.595 7.145 89.885 7.375 ;
        RECT 91.805 7.145 92.095 7.375 ;
      LAYER met2 ;
        RECT 24.280 7.715 24.560 8.095 ;
        RECT 40.865 7.715 41.145 8.095 ;
        RECT 57.450 7.720 57.730 8.100 ;
        RECT 74.035 7.725 74.315 8.105 ;
        RECT 90.615 7.725 90.895 8.105 ;
      LAYER met3 ;
        RECT 24.220 8.095 24.560 8.195 ;
        RECT 40.805 8.095 41.145 8.195 ;
        RECT 57.390 8.100 57.730 8.200 ;
        RECT 73.975 8.105 74.315 8.205 ;
        RECT 90.555 8.105 90.895 8.205 ;
        RECT 24.220 8.085 24.580 8.095 ;
        RECT 40.805 8.085 41.165 8.095 ;
        RECT 57.390 8.090 57.750 8.100 ;
        RECT 73.975 8.095 74.335 8.105 ;
        RECT 90.555 8.095 90.915 8.105 ;
        RECT 23.780 8.065 24.580 8.085 ;
        RECT 40.365 8.065 41.165 8.085 ;
        RECT 56.950 8.070 57.750 8.090 ;
        RECT 73.535 8.075 74.335 8.095 ;
        RECT 90.115 8.075 90.915 8.095 ;
        RECT 23.780 7.785 24.585 8.065 ;
        RECT 40.365 7.785 41.170 8.065 ;
        RECT 56.950 7.790 57.755 8.070 ;
        RECT 73.535 7.795 74.340 8.075 ;
        RECT 90.115 7.795 90.920 8.075 ;
        RECT 24.240 7.755 24.585 7.785 ;
        RECT 40.825 7.755 41.170 7.785 ;
        RECT 57.410 7.760 57.755 7.790 ;
        RECT 73.995 7.765 74.340 7.795 ;
        RECT 90.575 7.765 90.920 7.795 ;
        RECT 24.250 7.725 24.585 7.755 ;
        RECT 40.835 7.725 41.170 7.755 ;
        RECT 57.420 7.730 57.755 7.760 ;
        RECT 74.005 7.735 74.340 7.765 ;
        RECT 90.585 7.735 90.920 7.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 21.660 3.355 21.915 3.905 ;
        RECT 21.660 3.095 21.920 3.355 ;
        RECT 24.250 3.095 24.580 3.545 ;
        RECT 26.630 3.095 26.880 3.625 ;
        RECT 27.500 3.095 27.740 3.895 ;
        RECT 28.410 3.095 28.680 3.895 ;
        RECT 38.245 3.355 38.500 3.905 ;
        RECT 38.245 3.095 38.505 3.355 ;
        RECT 40.835 3.095 41.165 3.545 ;
        RECT 43.215 3.095 43.465 3.625 ;
        RECT 44.085 3.095 44.325 3.895 ;
        RECT 44.995 3.095 45.265 3.895 ;
        RECT 54.830 3.360 55.085 3.910 ;
        RECT 54.830 3.100 55.090 3.360 ;
        RECT 57.420 3.100 57.750 3.550 ;
        RECT 59.800 3.100 60.050 3.630 ;
        RECT 60.670 3.100 60.910 3.900 ;
        RECT 61.580 3.100 61.850 3.900 ;
        RECT 71.415 3.365 71.670 3.915 ;
        RECT 71.415 3.105 71.675 3.365 ;
        RECT 74.005 3.105 74.335 3.555 ;
        RECT 76.385 3.105 76.635 3.635 ;
        RECT 77.255 3.105 77.495 3.905 ;
        RECT 78.165 3.105 78.435 3.905 ;
        RECT 87.995 3.365 88.250 3.915 ;
        RECT 87.995 3.105 88.255 3.365 ;
        RECT 90.585 3.105 90.915 3.555 ;
        RECT 92.965 3.105 93.215 3.635 ;
        RECT 93.835 3.105 94.075 3.905 ;
        RECT 94.745 3.105 95.015 3.905 ;
        RECT 21.580 2.925 28.970 3.095 ;
        RECT 38.165 2.925 45.555 3.095 ;
        RECT 54.750 2.930 62.140 3.100 ;
        RECT 71.335 2.935 78.725 3.105 ;
        RECT 87.915 2.935 95.305 3.105 ;
        RECT 21.625 1.605 21.920 2.925 ;
        RECT 22.210 1.605 22.500 2.925 ;
        RECT 22.790 1.605 23.080 2.925 ;
        RECT 23.370 1.605 23.660 2.925 ;
        RECT 23.950 1.605 24.240 2.925 ;
        RECT 24.530 1.605 24.815 2.925 ;
        RECT 25.105 1.605 25.395 2.925 ;
        RECT 25.685 1.605 25.975 2.925 ;
        RECT 26.265 1.605 26.555 2.925 ;
        RECT 26.845 1.605 27.130 2.925 ;
        RECT 27.420 1.605 27.710 2.925 ;
        RECT 28.000 1.605 28.290 2.925 ;
        RECT 28.580 1.605 28.970 2.925 ;
        RECT 21.625 1.600 28.970 1.605 ;
        RECT 30.040 1.600 30.210 2.230 ;
        RECT 32.785 1.600 32.955 2.230 ;
        RECT 33.775 1.600 33.945 2.230 ;
        RECT 38.210 1.605 38.505 2.925 ;
        RECT 38.795 1.605 39.085 2.925 ;
        RECT 39.375 1.605 39.665 2.925 ;
        RECT 39.955 1.605 40.245 2.925 ;
        RECT 40.535 1.605 40.825 2.925 ;
        RECT 41.115 1.605 41.400 2.925 ;
        RECT 41.690 1.605 41.980 2.925 ;
        RECT 42.270 1.605 42.560 2.925 ;
        RECT 42.850 1.605 43.140 2.925 ;
        RECT 43.430 1.605 43.715 2.925 ;
        RECT 44.005 1.605 44.295 2.925 ;
        RECT 44.585 1.605 44.875 2.925 ;
        RECT 45.165 1.605 45.555 2.925 ;
        RECT 38.210 1.600 45.555 1.605 ;
        RECT 46.625 1.600 46.795 2.230 ;
        RECT 49.370 1.600 49.540 2.230 ;
        RECT 50.360 1.600 50.530 2.230 ;
        RECT 54.795 1.610 55.090 2.930 ;
        RECT 55.380 1.610 55.670 2.930 ;
        RECT 55.960 1.610 56.250 2.930 ;
        RECT 56.540 1.610 56.830 2.930 ;
        RECT 57.120 1.610 57.410 2.930 ;
        RECT 57.700 1.610 57.985 2.930 ;
        RECT 58.275 1.610 58.565 2.930 ;
        RECT 58.855 1.610 59.145 2.930 ;
        RECT 59.435 1.610 59.725 2.930 ;
        RECT 60.015 1.610 60.300 2.930 ;
        RECT 60.590 1.610 60.880 2.930 ;
        RECT 61.170 1.610 61.460 2.930 ;
        RECT 61.750 1.610 62.140 2.930 ;
        RECT 54.795 1.605 62.140 1.610 ;
        RECT 63.210 1.605 63.380 2.235 ;
        RECT 65.955 1.605 66.125 2.235 ;
        RECT 66.945 1.605 67.115 2.235 ;
        RECT 71.380 1.615 71.675 2.935 ;
        RECT 71.965 1.615 72.255 2.935 ;
        RECT 72.545 1.615 72.835 2.935 ;
        RECT 73.125 1.615 73.415 2.935 ;
        RECT 73.705 1.615 73.995 2.935 ;
        RECT 74.285 1.615 74.570 2.935 ;
        RECT 74.860 1.615 75.150 2.935 ;
        RECT 75.440 1.615 75.730 2.935 ;
        RECT 76.020 1.615 76.310 2.935 ;
        RECT 76.600 1.615 76.885 2.935 ;
        RECT 77.175 1.615 77.465 2.935 ;
        RECT 77.755 1.615 78.045 2.935 ;
        RECT 78.335 1.615 78.725 2.935 ;
        RECT 71.380 1.610 78.725 1.615 ;
        RECT 79.795 1.610 79.965 2.240 ;
        RECT 82.540 1.610 82.710 2.240 ;
        RECT 83.530 1.610 83.700 2.240 ;
        RECT 87.960 1.615 88.255 2.935 ;
        RECT 88.545 1.615 88.835 2.935 ;
        RECT 89.125 1.615 89.415 2.935 ;
        RECT 89.705 1.615 89.995 2.935 ;
        RECT 90.285 1.615 90.575 2.935 ;
        RECT 90.865 1.615 91.150 2.935 ;
        RECT 91.440 1.615 91.730 2.935 ;
        RECT 92.020 1.615 92.310 2.935 ;
        RECT 92.600 1.615 92.890 2.935 ;
        RECT 93.180 1.615 93.465 2.935 ;
        RECT 93.755 1.615 94.045 2.935 ;
        RECT 94.335 1.615 94.625 2.935 ;
        RECT 94.915 1.615 95.305 2.935 ;
        RECT 87.960 1.610 95.305 1.615 ;
        RECT 96.375 1.610 96.545 2.240 ;
        RECT 99.120 1.610 99.290 2.240 ;
        RECT 100.110 1.610 100.280 2.240 ;
        RECT 67.920 1.605 101.085 1.610 ;
        RECT 51.335 1.600 101.085 1.605 ;
        RECT 0.000 0.000 101.085 1.600 ;
      LAYER met1 ;
        RECT 21.580 2.765 28.970 3.125 ;
        RECT 38.165 2.765 45.555 3.125 ;
        RECT 54.750 2.770 62.140 3.130 ;
        RECT 71.335 2.775 78.725 3.135 ;
        RECT 87.915 2.775 95.305 3.135 ;
        RECT 21.625 1.605 21.920 2.765 ;
        RECT 22.210 1.605 22.500 2.765 ;
        RECT 22.790 1.605 23.080 2.765 ;
        RECT 23.370 1.605 23.660 2.765 ;
        RECT 23.950 1.605 24.240 2.765 ;
        RECT 24.530 1.605 24.815 2.765 ;
        RECT 25.105 1.605 25.395 2.765 ;
        RECT 25.685 1.605 25.975 2.765 ;
        RECT 26.265 1.605 26.555 2.765 ;
        RECT 26.845 1.605 27.130 2.765 ;
        RECT 27.420 1.605 27.710 2.765 ;
        RECT 28.000 1.605 28.290 2.765 ;
        RECT 28.580 1.605 28.970 2.765 ;
        RECT 21.625 1.600 28.970 1.605 ;
        RECT 38.210 1.605 38.505 2.765 ;
        RECT 38.795 1.605 39.085 2.765 ;
        RECT 39.375 1.605 39.665 2.765 ;
        RECT 39.955 1.605 40.245 2.765 ;
        RECT 40.535 1.605 40.825 2.765 ;
        RECT 41.115 1.605 41.400 2.765 ;
        RECT 41.690 1.605 41.980 2.765 ;
        RECT 42.270 1.605 42.560 2.765 ;
        RECT 42.850 1.605 43.140 2.765 ;
        RECT 43.430 1.605 43.715 2.765 ;
        RECT 44.005 1.605 44.295 2.765 ;
        RECT 44.585 1.605 44.875 2.765 ;
        RECT 45.165 1.605 45.555 2.765 ;
        RECT 54.795 1.610 55.090 2.770 ;
        RECT 55.380 1.610 55.670 2.770 ;
        RECT 55.960 1.610 56.250 2.770 ;
        RECT 56.540 1.610 56.830 2.770 ;
        RECT 57.120 1.610 57.410 2.770 ;
        RECT 57.700 1.610 57.985 2.770 ;
        RECT 58.275 1.610 58.565 2.770 ;
        RECT 58.855 1.610 59.145 2.770 ;
        RECT 59.435 1.610 59.725 2.770 ;
        RECT 60.015 1.610 60.300 2.770 ;
        RECT 60.590 1.610 60.880 2.770 ;
        RECT 61.170 1.610 61.460 2.770 ;
        RECT 61.750 1.610 62.140 2.770 ;
        RECT 71.380 1.615 71.675 2.775 ;
        RECT 71.965 1.615 72.255 2.775 ;
        RECT 72.545 1.615 72.835 2.775 ;
        RECT 73.125 1.615 73.415 2.775 ;
        RECT 73.705 1.615 73.995 2.775 ;
        RECT 74.285 1.615 74.570 2.775 ;
        RECT 74.860 1.615 75.150 2.775 ;
        RECT 75.440 1.615 75.730 2.775 ;
        RECT 76.020 1.615 76.310 2.775 ;
        RECT 76.600 1.615 76.885 2.775 ;
        RECT 77.175 1.615 77.465 2.775 ;
        RECT 77.755 1.615 78.045 2.775 ;
        RECT 78.335 1.615 78.725 2.775 ;
        RECT 71.380 1.610 78.725 1.615 ;
        RECT 87.960 1.615 88.255 2.775 ;
        RECT 88.545 1.615 88.835 2.775 ;
        RECT 89.125 1.615 89.415 2.775 ;
        RECT 89.705 1.615 89.995 2.775 ;
        RECT 90.285 1.615 90.575 2.775 ;
        RECT 90.865 1.615 91.150 2.775 ;
        RECT 91.440 1.615 91.730 2.775 ;
        RECT 92.020 1.615 92.310 2.775 ;
        RECT 92.600 1.615 92.890 2.775 ;
        RECT 93.180 1.615 93.465 2.775 ;
        RECT 93.755 1.615 94.045 2.775 ;
        RECT 94.335 1.615 94.625 2.775 ;
        RECT 94.915 1.615 95.305 2.775 ;
        RECT 87.960 1.610 95.305 1.615 ;
        RECT 54.795 1.605 62.140 1.610 ;
        RECT 67.920 1.605 101.085 1.610 ;
        RECT 38.210 1.600 45.555 1.605 ;
        RECT 51.335 1.600 101.085 1.605 ;
        RECT 0.000 0.000 101.085 1.600 ;
    END
  END vssd1
  OBS
      LAYER pwell ;
        RECT 21.680 8.335 22.410 8.745 ;
        RECT 24.320 8.495 24.490 8.525 ;
        RECT 27.540 8.495 27.710 8.525 ;
        RECT 24.320 8.335 24.900 8.495 ;
        RECT 27.540 8.385 28.170 8.495 ;
        RECT 27.540 8.335 27.850 8.385 ;
        RECT 21.680 8.145 27.850 8.335 ;
        RECT 38.265 8.335 38.995 8.745 ;
        RECT 40.905 8.495 41.075 8.525 ;
        RECT 44.125 8.495 44.295 8.525 ;
        RECT 40.905 8.335 41.485 8.495 ;
        RECT 44.125 8.385 44.755 8.495 ;
        RECT 44.125 8.335 44.435 8.385 ;
        RECT 38.265 8.145 44.435 8.335 ;
        RECT 54.850 8.340 55.580 8.750 ;
        RECT 57.490 8.500 57.660 8.530 ;
        RECT 60.710 8.500 60.880 8.530 ;
        RECT 57.490 8.340 58.070 8.500 ;
        RECT 60.710 8.390 61.340 8.500 ;
        RECT 60.710 8.340 61.020 8.390 ;
        RECT 54.850 8.150 61.020 8.340 ;
        RECT 71.435 8.345 72.165 8.755 ;
        RECT 74.075 8.505 74.245 8.535 ;
        RECT 77.295 8.505 77.465 8.535 ;
        RECT 74.075 8.345 74.655 8.505 ;
        RECT 77.295 8.395 77.925 8.505 ;
        RECT 77.295 8.345 77.605 8.395 ;
        RECT 71.435 8.155 77.605 8.345 ;
        RECT 88.015 8.345 88.745 8.755 ;
        RECT 90.655 8.505 90.825 8.535 ;
        RECT 93.875 8.505 94.045 8.535 ;
        RECT 90.655 8.345 91.235 8.505 ;
        RECT 93.875 8.395 94.505 8.505 ;
        RECT 93.875 8.345 94.185 8.395 ;
        RECT 88.015 8.155 94.185 8.345 ;
        RECT 22.540 7.515 27.850 8.145 ;
        RECT 22.540 7.425 23.490 7.515 ;
        RECT 25.100 7.425 27.850 7.515 ;
        RECT 39.125 7.515 44.435 8.145 ;
        RECT 39.125 7.425 40.075 7.515 ;
        RECT 41.685 7.425 44.435 7.515 ;
        RECT 55.710 7.520 61.020 8.150 ;
        RECT 55.710 7.430 56.660 7.520 ;
        RECT 58.270 7.430 61.020 7.520 ;
        RECT 72.295 7.525 77.605 8.155 ;
        RECT 72.295 7.435 73.245 7.525 ;
        RECT 74.855 7.435 77.605 7.525 ;
        RECT 88.875 7.525 94.185 8.155 ;
        RECT 88.875 7.435 89.825 7.525 ;
        RECT 91.435 7.435 94.185 7.525 ;
        RECT 21.580 3.815 22.810 4.015 ;
        RECT 24.140 3.815 25.090 4.015 ;
        RECT 21.580 3.790 25.090 3.815 ;
        RECT 26.470 3.790 28.750 4.015 ;
        RECT 21.580 3.305 28.750 3.790 ;
        RECT 38.165 3.815 39.395 4.015 ;
        RECT 40.725 3.815 41.675 4.015 ;
        RECT 38.165 3.790 41.675 3.815 ;
        RECT 43.055 3.790 45.335 4.015 ;
        RECT 38.165 3.305 45.335 3.790 ;
        RECT 54.750 3.820 55.980 4.020 ;
        RECT 57.310 3.820 58.260 4.020 ;
        RECT 54.750 3.795 58.260 3.820 ;
        RECT 59.640 3.795 61.920 4.020 ;
        RECT 54.750 3.310 61.920 3.795 ;
        RECT 71.335 3.825 72.565 4.025 ;
        RECT 73.895 3.825 74.845 4.025 ;
        RECT 71.335 3.800 74.845 3.825 ;
        RECT 76.225 3.800 78.505 4.025 ;
        RECT 71.335 3.315 78.505 3.800 ;
        RECT 87.915 3.825 89.145 4.025 ;
        RECT 90.475 3.825 91.425 4.025 ;
        RECT 87.915 3.800 91.425 3.825 ;
        RECT 92.805 3.800 95.085 4.025 ;
        RECT 87.915 3.315 95.085 3.800 ;
        RECT 21.520 3.135 28.750 3.305 ;
        RECT 21.520 2.705 22.110 3.135 ;
        RECT 24.160 3.110 28.750 3.135 ;
        RECT 38.105 3.135 45.335 3.305 ;
        RECT 25.240 2.925 25.410 3.105 ;
        RECT 27.550 3.095 27.720 3.105 ;
        RECT 27.540 3.085 27.720 3.095 ;
        RECT 27.550 2.925 27.720 3.085 ;
        RECT 38.105 2.705 38.695 3.135 ;
        RECT 40.745 3.110 45.335 3.135 ;
        RECT 54.690 3.140 61.920 3.310 ;
        RECT 41.825 2.925 41.995 3.105 ;
        RECT 44.135 3.095 44.305 3.105 ;
        RECT 44.125 3.085 44.305 3.095 ;
        RECT 44.135 2.925 44.305 3.085 ;
        RECT 54.690 2.710 55.280 3.140 ;
        RECT 57.330 3.115 61.920 3.140 ;
        RECT 71.275 3.145 78.505 3.315 ;
        RECT 58.410 2.930 58.580 3.110 ;
        RECT 60.720 3.100 60.890 3.110 ;
        RECT 60.710 3.090 60.890 3.100 ;
        RECT 60.720 2.930 60.890 3.090 ;
        RECT 71.275 2.715 71.865 3.145 ;
        RECT 73.915 3.120 78.505 3.145 ;
        RECT 87.855 3.145 95.085 3.315 ;
        RECT 74.995 2.935 75.165 3.115 ;
        RECT 77.305 3.105 77.475 3.115 ;
        RECT 77.295 3.095 77.475 3.105 ;
        RECT 77.305 2.935 77.475 3.095 ;
        RECT 87.855 2.715 88.445 3.145 ;
        RECT 90.495 3.120 95.085 3.145 ;
        RECT 91.575 2.935 91.745 3.115 ;
        RECT 93.885 3.105 94.055 3.115 ;
        RECT 93.875 3.095 94.055 3.105 ;
        RECT 93.885 2.935 94.055 3.095 ;
      LAYER li1 ;
        RECT 16.015 10.095 16.190 10.585 ;
        RECT 16.540 10.305 16.710 10.585 ;
        RECT 16.540 10.135 16.770 10.305 ;
        RECT 16.015 9.925 16.185 10.095 ;
        RECT 16.015 9.595 16.425 9.925 ;
        RECT 16.015 9.085 16.185 9.595 ;
        RECT 16.015 8.755 16.425 9.085 ;
        RECT 16.015 8.555 16.185 8.755 ;
        RECT 16.015 7.295 16.190 8.555 ;
        RECT 16.600 8.525 16.770 10.135 ;
        RECT 16.970 10.075 17.145 10.585 ;
        RECT 19.245 10.095 19.420 10.585 ;
        RECT 19.245 9.925 19.415 10.095 ;
        RECT 20.200 10.075 20.375 10.585 ;
        RECT 20.630 10.035 20.805 10.585 ;
        RECT 30.470 10.100 30.645 10.590 ;
        RECT 30.995 10.310 31.165 10.590 ;
        RECT 30.995 10.140 31.225 10.310 ;
        RECT 19.245 9.595 19.655 9.925 ;
        RECT 16.540 8.355 16.770 8.525 ;
        RECT 16.970 8.555 17.140 9.505 ;
        RECT 19.245 9.085 19.415 9.595 ;
        RECT 19.245 8.755 19.655 9.085 ;
        RECT 19.245 8.555 19.415 8.755 ;
        RECT 20.200 8.555 20.370 9.505 ;
        RECT 16.540 7.295 16.710 8.355 ;
        RECT 16.970 7.295 17.145 8.555 ;
        RECT 19.245 7.295 19.420 8.555 ;
        RECT 20.200 7.295 20.375 8.555 ;
        RECT 20.630 8.435 20.800 10.035 ;
        RECT 30.470 9.930 30.640 10.100 ;
        RECT 30.470 9.600 30.880 9.930 ;
        RECT 30.470 9.090 30.640 9.600 ;
        RECT 30.470 8.760 30.880 9.090 ;
        RECT 30.470 8.560 30.640 8.760 ;
        RECT 20.630 7.295 20.805 8.435 ;
        RECT 22.420 7.895 22.980 8.185 ;
        RECT 24.020 8.055 24.280 8.085 ;
        RECT 22.420 6.525 22.670 7.895 ;
        RECT 24.020 7.725 24.350 8.055 ;
        RECT 25.730 7.935 27.040 8.185 ;
        RECT 25.730 7.785 25.910 7.935 ;
        RECT 22.960 7.535 24.350 7.725 ;
        RECT 25.180 7.615 25.910 7.785 ;
        RECT 22.960 7.445 23.130 7.535 ;
        RECT 22.840 7.115 23.130 7.445 ;
        RECT 23.860 7.115 24.540 7.365 ;
        RECT 22.960 6.865 23.130 7.115 ;
        RECT 22.960 6.695 23.905 6.865 ;
        RECT 24.270 6.755 24.540 7.115 ;
        RECT 25.180 6.945 25.350 7.615 ;
        RECT 26.160 7.365 26.370 7.765 ;
        RECT 26.020 7.165 26.370 7.365 ;
        RECT 26.620 7.365 26.870 7.765 ;
        RECT 26.620 7.165 27.090 7.365 ;
        RECT 27.280 7.165 27.730 7.675 ;
        RECT 30.470 7.300 30.645 8.560 ;
        RECT 31.055 8.530 31.225 10.140 ;
        RECT 31.425 10.080 31.600 10.590 ;
        RECT 31.855 10.040 32.030 10.590 ;
        RECT 33.220 10.080 33.390 10.590 ;
        RECT 34.210 10.080 34.380 10.590 ;
        RECT 35.830 10.095 36.005 10.585 ;
        RECT 30.995 8.360 31.225 8.530 ;
        RECT 31.425 8.560 31.595 9.510 ;
        RECT 30.995 7.300 31.165 8.360 ;
        RECT 31.425 7.300 31.600 8.560 ;
        RECT 31.855 8.440 32.025 10.040 ;
        RECT 35.830 9.925 36.000 10.095 ;
        RECT 36.785 10.075 36.960 10.585 ;
        RECT 37.215 10.035 37.390 10.585 ;
        RECT 47.055 10.100 47.230 10.590 ;
        RECT 47.580 10.310 47.750 10.590 ;
        RECT 47.580 10.140 47.810 10.310 ;
        RECT 35.830 9.595 36.240 9.925 ;
        RECT 32.395 9.420 32.625 9.570 ;
        RECT 32.395 9.250 33.315 9.420 ;
        RECT 33.835 9.250 34.305 9.420 ;
        RECT 32.845 8.560 33.015 9.250 ;
        RECT 33.215 8.770 33.385 8.880 ;
        RECT 33.835 8.770 34.005 9.250 ;
        RECT 35.830 9.085 36.000 9.595 ;
        RECT 33.215 8.600 34.005 8.770 ;
        RECT 31.855 7.300 32.030 8.440 ;
        RECT 33.215 7.300 33.390 8.600 ;
        RECT 33.835 8.560 34.005 8.600 ;
        RECT 34.205 8.445 34.375 8.880 ;
        RECT 35.830 8.755 36.240 9.085 ;
        RECT 35.830 8.555 36.000 8.755 ;
        RECT 36.785 8.555 36.955 9.505 ;
        RECT 34.205 7.300 34.380 8.445 ;
        RECT 35.830 7.295 36.005 8.555 ;
        RECT 36.785 7.295 36.960 8.555 ;
        RECT 37.215 8.435 37.385 10.035 ;
        RECT 47.055 9.930 47.225 10.100 ;
        RECT 47.055 9.600 47.465 9.930 ;
        RECT 47.055 9.090 47.225 9.600 ;
        RECT 47.055 8.760 47.465 9.090 ;
        RECT 47.055 8.560 47.225 8.760 ;
        RECT 37.215 7.295 37.390 8.435 ;
        RECT 39.005 7.895 39.565 8.185 ;
        RECT 40.605 8.055 40.865 8.085 ;
        RECT 26.020 6.945 27.760 6.995 ;
        RECT 25.180 6.815 27.760 6.945 ;
        RECT 25.180 6.775 26.240 6.815 ;
        RECT 22.420 5.975 22.880 6.525 ;
        RECT 23.600 5.975 23.905 6.695 ;
        RECT 26.380 6.605 27.260 6.645 ;
        RECT 25.730 6.405 27.260 6.605 ;
        RECT 25.730 6.275 25.900 6.405 ;
        RECT 26.650 6.355 27.260 6.405 ;
        RECT 27.030 6.315 27.260 6.355 ;
        RECT 27.430 6.315 27.760 6.815 ;
        RECT 39.005 6.525 39.255 7.895 ;
        RECT 40.605 7.725 40.935 8.055 ;
        RECT 42.315 7.935 43.625 8.185 ;
        RECT 42.315 7.785 42.495 7.935 ;
        RECT 39.545 7.535 40.935 7.725 ;
        RECT 41.765 7.615 42.495 7.785 ;
        RECT 39.545 7.445 39.715 7.535 ;
        RECT 39.425 7.115 39.715 7.445 ;
        RECT 40.445 7.115 41.125 7.365 ;
        RECT 39.545 6.865 39.715 7.115 ;
        RECT 39.545 6.695 40.490 6.865 ;
        RECT 40.855 6.755 41.125 7.115 ;
        RECT 41.765 6.945 41.935 7.615 ;
        RECT 42.745 7.365 42.955 7.765 ;
        RECT 42.605 7.165 42.955 7.365 ;
        RECT 43.205 7.365 43.455 7.765 ;
        RECT 43.205 7.165 43.675 7.365 ;
        RECT 43.865 7.165 44.315 7.675 ;
        RECT 47.055 7.300 47.230 8.560 ;
        RECT 47.640 8.530 47.810 10.140 ;
        RECT 48.010 10.080 48.185 10.590 ;
        RECT 48.440 10.040 48.615 10.590 ;
        RECT 49.805 10.080 49.975 10.590 ;
        RECT 50.795 10.080 50.965 10.590 ;
        RECT 52.415 10.100 52.590 10.590 ;
        RECT 47.580 8.360 47.810 8.530 ;
        RECT 48.010 8.560 48.180 9.510 ;
        RECT 47.580 7.300 47.750 8.360 ;
        RECT 48.010 7.300 48.185 8.560 ;
        RECT 48.440 8.440 48.610 10.040 ;
        RECT 52.415 9.930 52.585 10.100 ;
        RECT 53.370 10.080 53.545 10.590 ;
        RECT 53.800 10.040 53.975 10.590 ;
        RECT 63.640 10.105 63.815 10.595 ;
        RECT 64.165 10.315 64.335 10.595 ;
        RECT 64.165 10.145 64.395 10.315 ;
        RECT 52.415 9.600 52.825 9.930 ;
        RECT 48.980 9.420 49.210 9.570 ;
        RECT 48.980 9.250 49.900 9.420 ;
        RECT 50.420 9.250 50.890 9.420 ;
        RECT 49.430 8.560 49.600 9.250 ;
        RECT 49.800 8.770 49.970 8.880 ;
        RECT 50.420 8.770 50.590 9.250 ;
        RECT 52.415 9.090 52.585 9.600 ;
        RECT 49.800 8.600 50.590 8.770 ;
        RECT 48.440 7.300 48.615 8.440 ;
        RECT 49.800 7.300 49.975 8.600 ;
        RECT 50.420 8.560 50.590 8.600 ;
        RECT 50.790 8.445 50.960 8.880 ;
        RECT 52.415 8.760 52.825 9.090 ;
        RECT 52.415 8.560 52.585 8.760 ;
        RECT 53.370 8.560 53.540 9.510 ;
        RECT 50.790 7.300 50.965 8.445 ;
        RECT 52.415 7.300 52.590 8.560 ;
        RECT 53.370 7.300 53.545 8.560 ;
        RECT 53.800 8.440 53.970 10.040 ;
        RECT 63.640 9.935 63.810 10.105 ;
        RECT 63.640 9.605 64.050 9.935 ;
        RECT 63.640 9.095 63.810 9.605 ;
        RECT 63.640 8.765 64.050 9.095 ;
        RECT 63.640 8.565 63.810 8.765 ;
        RECT 53.800 7.300 53.975 8.440 ;
        RECT 55.590 7.900 56.150 8.190 ;
        RECT 57.190 8.060 57.450 8.090 ;
        RECT 42.605 6.945 44.345 6.995 ;
        RECT 41.765 6.815 44.345 6.945 ;
        RECT 41.765 6.775 42.825 6.815 ;
        RECT 26.590 6.145 26.920 6.185 ;
        RECT 27.430 6.145 28.250 6.315 ;
        RECT 26.590 5.975 27.760 6.145 ;
        RECT 39.005 5.975 39.465 6.525 ;
        RECT 40.185 5.975 40.490 6.695 ;
        RECT 42.965 6.605 43.845 6.645 ;
        RECT 42.315 6.405 43.845 6.605 ;
        RECT 42.315 6.275 42.485 6.405 ;
        RECT 43.235 6.355 43.845 6.405 ;
        RECT 43.615 6.315 43.845 6.355 ;
        RECT 44.015 6.315 44.345 6.815 ;
        RECT 55.590 6.530 55.840 7.900 ;
        RECT 57.190 7.730 57.520 8.060 ;
        RECT 58.900 7.940 60.210 8.190 ;
        RECT 58.900 7.790 59.080 7.940 ;
        RECT 56.130 7.540 57.520 7.730 ;
        RECT 58.350 7.620 59.080 7.790 ;
        RECT 56.130 7.450 56.300 7.540 ;
        RECT 56.010 7.120 56.300 7.450 ;
        RECT 57.030 7.120 57.710 7.370 ;
        RECT 56.130 6.870 56.300 7.120 ;
        RECT 56.130 6.700 57.075 6.870 ;
        RECT 57.440 6.760 57.710 7.120 ;
        RECT 58.350 6.950 58.520 7.620 ;
        RECT 59.330 7.370 59.540 7.770 ;
        RECT 59.190 7.170 59.540 7.370 ;
        RECT 59.790 7.370 60.040 7.770 ;
        RECT 59.790 7.170 60.260 7.370 ;
        RECT 60.450 7.170 60.900 7.680 ;
        RECT 63.640 7.305 63.815 8.565 ;
        RECT 64.225 8.535 64.395 10.145 ;
        RECT 64.595 10.085 64.770 10.595 ;
        RECT 65.025 10.045 65.200 10.595 ;
        RECT 66.390 10.085 66.560 10.595 ;
        RECT 67.380 10.085 67.550 10.595 ;
        RECT 69.000 10.105 69.175 10.595 ;
        RECT 64.165 8.365 64.395 8.535 ;
        RECT 64.595 8.565 64.765 9.515 ;
        RECT 64.165 7.305 64.335 8.365 ;
        RECT 64.595 7.305 64.770 8.565 ;
        RECT 65.025 8.445 65.195 10.045 ;
        RECT 69.000 9.935 69.170 10.105 ;
        RECT 69.955 10.085 70.130 10.595 ;
        RECT 70.385 10.045 70.560 10.595 ;
        RECT 80.225 10.110 80.400 10.600 ;
        RECT 80.750 10.320 80.920 10.600 ;
        RECT 80.750 10.150 80.980 10.320 ;
        RECT 69.000 9.605 69.410 9.935 ;
        RECT 65.565 9.425 65.795 9.575 ;
        RECT 65.565 9.255 66.485 9.425 ;
        RECT 67.005 9.255 67.475 9.425 ;
        RECT 66.015 8.565 66.185 9.255 ;
        RECT 66.385 8.775 66.555 8.885 ;
        RECT 67.005 8.775 67.175 9.255 ;
        RECT 69.000 9.095 69.170 9.605 ;
        RECT 66.385 8.605 67.175 8.775 ;
        RECT 65.025 7.305 65.200 8.445 ;
        RECT 66.385 7.305 66.560 8.605 ;
        RECT 67.005 8.565 67.175 8.605 ;
        RECT 67.375 8.450 67.545 8.885 ;
        RECT 69.000 8.765 69.410 9.095 ;
        RECT 69.000 8.565 69.170 8.765 ;
        RECT 69.955 8.565 70.125 9.515 ;
        RECT 67.375 7.305 67.550 8.450 ;
        RECT 69.000 7.305 69.175 8.565 ;
        RECT 69.955 7.305 70.130 8.565 ;
        RECT 70.385 8.445 70.555 10.045 ;
        RECT 80.225 9.940 80.395 10.110 ;
        RECT 80.225 9.610 80.635 9.940 ;
        RECT 80.225 9.100 80.395 9.610 ;
        RECT 80.225 8.770 80.635 9.100 ;
        RECT 80.225 8.570 80.395 8.770 ;
        RECT 70.385 7.305 70.560 8.445 ;
        RECT 72.175 7.905 72.735 8.195 ;
        RECT 73.775 8.065 74.035 8.095 ;
        RECT 59.190 6.950 60.930 7.000 ;
        RECT 58.350 6.820 60.930 6.950 ;
        RECT 58.350 6.780 59.410 6.820 ;
        RECT 43.175 6.145 43.505 6.185 ;
        RECT 44.015 6.145 44.835 6.315 ;
        RECT 43.175 5.975 44.345 6.145 ;
        RECT 55.590 5.980 56.050 6.530 ;
        RECT 56.770 5.980 57.075 6.700 ;
        RECT 59.550 6.610 60.430 6.650 ;
        RECT 58.900 6.410 60.430 6.610 ;
        RECT 58.900 6.280 59.070 6.410 ;
        RECT 59.820 6.360 60.430 6.410 ;
        RECT 60.200 6.320 60.430 6.360 ;
        RECT 60.600 6.320 60.930 6.820 ;
        RECT 72.175 6.535 72.425 7.905 ;
        RECT 73.775 7.735 74.105 8.065 ;
        RECT 75.485 7.945 76.795 8.195 ;
        RECT 75.485 7.795 75.665 7.945 ;
        RECT 72.715 7.545 74.105 7.735 ;
        RECT 74.935 7.625 75.665 7.795 ;
        RECT 72.715 7.455 72.885 7.545 ;
        RECT 72.595 7.125 72.885 7.455 ;
        RECT 73.615 7.125 74.295 7.375 ;
        RECT 72.715 6.875 72.885 7.125 ;
        RECT 72.715 6.705 73.660 6.875 ;
        RECT 74.025 6.765 74.295 7.125 ;
        RECT 74.935 6.955 75.105 7.625 ;
        RECT 75.915 7.375 76.125 7.775 ;
        RECT 75.775 7.175 76.125 7.375 ;
        RECT 76.375 7.375 76.625 7.775 ;
        RECT 76.375 7.175 76.845 7.375 ;
        RECT 77.035 7.175 77.485 7.685 ;
        RECT 80.225 7.310 80.400 8.570 ;
        RECT 80.810 8.540 80.980 10.150 ;
        RECT 81.180 10.090 81.355 10.600 ;
        RECT 81.610 10.050 81.785 10.600 ;
        RECT 82.975 10.090 83.145 10.600 ;
        RECT 83.965 10.090 84.135 10.600 ;
        RECT 85.580 10.105 85.755 10.595 ;
        RECT 80.750 8.370 80.980 8.540 ;
        RECT 81.180 8.570 81.350 9.520 ;
        RECT 80.750 7.310 80.920 8.370 ;
        RECT 81.180 7.310 81.355 8.570 ;
        RECT 81.610 8.450 81.780 10.050 ;
        RECT 85.580 9.935 85.750 10.105 ;
        RECT 86.535 10.085 86.710 10.595 ;
        RECT 86.965 10.045 87.140 10.595 ;
        RECT 96.805 10.110 96.980 10.600 ;
        RECT 97.330 10.320 97.500 10.600 ;
        RECT 97.330 10.150 97.560 10.320 ;
        RECT 85.580 9.605 85.990 9.935 ;
        RECT 82.150 9.430 82.380 9.580 ;
        RECT 82.150 9.260 83.070 9.430 ;
        RECT 83.590 9.260 84.060 9.430 ;
        RECT 82.600 8.570 82.770 9.260 ;
        RECT 82.970 8.780 83.140 8.890 ;
        RECT 83.590 8.780 83.760 9.260 ;
        RECT 85.580 9.095 85.750 9.605 ;
        RECT 82.970 8.610 83.760 8.780 ;
        RECT 81.610 7.310 81.785 8.450 ;
        RECT 82.970 7.310 83.145 8.610 ;
        RECT 83.590 8.570 83.760 8.610 ;
        RECT 83.960 8.455 84.130 8.890 ;
        RECT 85.580 8.765 85.990 9.095 ;
        RECT 85.580 8.565 85.750 8.765 ;
        RECT 86.535 8.565 86.705 9.515 ;
        RECT 83.960 7.310 84.135 8.455 ;
        RECT 85.580 7.305 85.755 8.565 ;
        RECT 86.535 7.305 86.710 8.565 ;
        RECT 86.965 8.445 87.135 10.045 ;
        RECT 96.805 9.940 96.975 10.110 ;
        RECT 96.805 9.610 97.215 9.940 ;
        RECT 96.805 9.100 96.975 9.610 ;
        RECT 96.805 8.770 97.215 9.100 ;
        RECT 96.805 8.570 96.975 8.770 ;
        RECT 86.965 7.305 87.140 8.445 ;
        RECT 88.755 7.905 89.315 8.195 ;
        RECT 90.355 8.065 90.615 8.095 ;
        RECT 75.775 6.955 77.515 7.005 ;
        RECT 74.935 6.825 77.515 6.955 ;
        RECT 74.935 6.785 75.995 6.825 ;
        RECT 59.760 6.150 60.090 6.190 ;
        RECT 60.600 6.150 61.420 6.320 ;
        RECT 59.760 5.980 60.930 6.150 ;
        RECT 72.175 5.985 72.635 6.535 ;
        RECT 73.355 5.985 73.660 6.705 ;
        RECT 76.135 6.615 77.015 6.655 ;
        RECT 75.485 6.415 77.015 6.615 ;
        RECT 75.485 6.285 75.655 6.415 ;
        RECT 76.405 6.365 77.015 6.415 ;
        RECT 76.785 6.325 77.015 6.365 ;
        RECT 77.185 6.325 77.515 6.825 ;
        RECT 88.755 6.535 89.005 7.905 ;
        RECT 90.355 7.735 90.685 8.065 ;
        RECT 92.065 7.945 93.375 8.195 ;
        RECT 92.065 7.795 92.245 7.945 ;
        RECT 89.295 7.545 90.685 7.735 ;
        RECT 91.515 7.625 92.245 7.795 ;
        RECT 89.295 7.455 89.465 7.545 ;
        RECT 89.175 7.125 89.465 7.455 ;
        RECT 90.195 7.125 90.875 7.375 ;
        RECT 89.295 6.875 89.465 7.125 ;
        RECT 89.295 6.705 90.240 6.875 ;
        RECT 90.605 6.765 90.875 7.125 ;
        RECT 91.515 6.955 91.685 7.625 ;
        RECT 92.495 7.375 92.705 7.775 ;
        RECT 92.355 7.175 92.705 7.375 ;
        RECT 92.955 7.375 93.205 7.775 ;
        RECT 92.955 7.175 93.425 7.375 ;
        RECT 93.615 7.175 94.065 7.685 ;
        RECT 96.805 7.310 96.980 8.570 ;
        RECT 97.390 8.540 97.560 10.150 ;
        RECT 97.760 10.090 97.935 10.600 ;
        RECT 98.190 10.050 98.365 10.600 ;
        RECT 99.555 10.090 99.725 10.600 ;
        RECT 100.545 10.090 100.715 10.600 ;
        RECT 97.330 8.370 97.560 8.540 ;
        RECT 97.760 8.570 97.930 9.520 ;
        RECT 97.330 7.310 97.500 8.370 ;
        RECT 97.760 7.310 97.935 8.570 ;
        RECT 98.190 8.450 98.360 10.050 ;
        RECT 98.730 9.430 98.960 9.580 ;
        RECT 98.730 9.260 99.650 9.430 ;
        RECT 100.170 9.260 100.640 9.430 ;
        RECT 99.180 8.570 99.350 9.260 ;
        RECT 99.550 8.780 99.720 8.890 ;
        RECT 100.170 8.780 100.340 9.260 ;
        RECT 99.550 8.610 100.340 8.780 ;
        RECT 98.190 7.310 98.365 8.450 ;
        RECT 99.550 7.310 99.725 8.610 ;
        RECT 100.170 8.570 100.340 8.610 ;
        RECT 100.540 8.455 100.710 8.890 ;
        RECT 100.540 7.310 100.715 8.455 ;
        RECT 92.355 6.955 94.095 7.005 ;
        RECT 91.515 6.825 94.095 6.955 ;
        RECT 91.515 6.785 92.575 6.825 ;
        RECT 76.345 6.155 76.675 6.195 ;
        RECT 77.185 6.155 78.005 6.325 ;
        RECT 76.345 5.985 77.515 6.155 ;
        RECT 88.755 5.985 89.215 6.535 ;
        RECT 89.935 5.985 90.240 6.705 ;
        RECT 92.715 6.615 93.595 6.655 ;
        RECT 92.065 6.415 93.595 6.615 ;
        RECT 92.065 6.285 92.235 6.415 ;
        RECT 92.985 6.365 93.595 6.415 ;
        RECT 93.365 6.325 93.595 6.365 ;
        RECT 93.765 6.325 94.095 6.825 ;
        RECT 92.925 6.155 93.255 6.195 ;
        RECT 93.765 6.155 94.585 6.325 ;
        RECT 92.925 5.985 94.095 6.155 ;
        RECT 22.175 5.125 22.345 5.465 ;
        RECT 23.670 5.125 24.140 5.465 ;
        RECT 22.170 5.065 22.345 5.125 ;
        RECT 21.660 4.075 22.000 4.955 ;
        RECT 22.170 4.245 22.340 5.065 ;
        RECT 22.880 4.595 23.130 4.965 ;
        RECT 23.850 4.595 24.570 4.895 ;
        RECT 24.740 4.765 25.010 5.465 ;
        RECT 25.960 5.125 26.440 5.465 ;
        RECT 22.880 4.425 24.670 4.595 ;
        RECT 22.170 3.995 23.270 4.245 ;
        RECT 22.170 3.905 22.420 3.995 ;
        RECT 22.120 3.485 22.420 3.905 ;
        RECT 23.440 3.575 23.690 4.425 ;
        RECT 22.900 3.305 23.690 3.575 ;
        RECT 23.860 3.725 24.270 4.245 ;
        RECT 24.440 3.995 24.670 4.425 ;
        RECT 24.840 3.735 25.010 4.765 ;
        RECT 25.180 4.365 25.440 4.815 ;
        RECT 26.110 4.635 26.870 4.885 ;
        RECT 27.040 4.765 27.310 5.465 ;
        RECT 26.100 4.605 26.870 4.635 ;
        RECT 26.080 4.595 26.870 4.605 ;
        RECT 26.080 4.575 26.970 4.595 ;
        RECT 26.060 4.565 26.970 4.575 ;
        RECT 26.040 4.555 26.970 4.565 ;
        RECT 26.010 4.545 26.970 4.555 ;
        RECT 25.940 4.515 26.970 4.545 ;
        RECT 25.920 4.485 26.970 4.515 ;
        RECT 25.900 4.455 26.970 4.485 ;
        RECT 25.870 4.425 26.970 4.455 ;
        RECT 25.840 4.395 26.970 4.425 ;
        RECT 25.810 4.385 26.970 4.395 ;
        RECT 25.810 4.375 26.170 4.385 ;
        RECT 25.810 4.365 26.160 4.375 ;
        RECT 25.180 4.355 26.140 4.365 ;
        RECT 25.180 4.345 26.130 4.355 ;
        RECT 25.180 4.325 26.110 4.345 ;
        RECT 25.180 4.315 26.100 4.325 ;
        RECT 25.180 4.195 26.070 4.315 ;
        RECT 23.860 3.305 24.060 3.725 ;
        RECT 24.750 3.265 25.010 3.735 ;
        RECT 25.180 3.635 25.730 4.025 ;
        RECT 25.900 3.465 26.070 4.195 ;
        RECT 25.180 3.295 26.070 3.465 ;
        RECT 26.240 3.795 26.570 4.215 ;
        RECT 26.740 3.995 26.970 4.385 ;
        RECT 27.140 4.275 27.310 4.765 ;
        RECT 27.490 4.665 27.820 5.455 ;
        RECT 27.490 4.495 28.170 4.665 ;
        RECT 27.480 4.275 27.830 4.325 ;
        RECT 27.140 4.105 27.830 4.275 ;
        RECT 26.240 3.305 26.460 3.795 ;
        RECT 27.140 3.735 27.310 4.105 ;
        RECT 27.480 4.075 27.830 4.105 ;
        RECT 28.000 3.895 28.170 4.495 ;
        RECT 28.340 4.075 28.690 4.325 ;
        RECT 30.470 3.900 30.645 5.160 ;
        RECT 30.995 4.100 31.165 5.160 ;
        RECT 30.995 3.930 31.225 4.100 ;
        RECT 27.050 3.265 27.310 3.735 ;
        RECT 27.910 3.265 28.240 3.895 ;
        RECT 30.470 3.700 30.640 3.900 ;
        RECT 30.470 3.370 30.880 3.700 ;
        RECT 30.470 2.860 30.640 3.370 ;
        RECT 30.470 2.530 30.880 2.860 ;
        RECT 30.470 2.360 30.640 2.530 ;
        RECT 30.470 1.870 30.645 2.360 ;
        RECT 31.055 2.320 31.225 3.930 ;
        RECT 31.425 3.900 31.600 5.160 ;
        RECT 31.855 4.020 32.030 5.160 ;
        RECT 31.425 2.950 31.595 3.900 ;
        RECT 31.855 2.420 32.025 4.020 ;
        RECT 33.215 4.015 33.390 5.160 ;
        RECT 38.760 5.125 38.930 5.465 ;
        RECT 40.255 5.125 40.725 5.465 ;
        RECT 38.755 5.065 38.930 5.125 ;
        RECT 38.245 4.075 38.585 4.955 ;
        RECT 38.755 4.245 38.925 5.065 ;
        RECT 39.465 4.595 39.715 4.965 ;
        RECT 40.435 4.595 41.155 4.895 ;
        RECT 41.325 4.765 41.595 5.465 ;
        RECT 42.545 5.125 43.025 5.465 ;
        RECT 39.465 4.425 41.255 4.595 ;
        RECT 32.845 3.210 33.015 3.900 ;
        RECT 33.215 3.800 33.385 4.015 ;
        RECT 38.755 3.995 39.855 4.245 ;
        RECT 38.755 3.905 39.005 3.995 ;
        RECT 33.835 3.800 34.005 3.900 ;
        RECT 33.215 3.630 34.005 3.800 ;
        RECT 33.215 3.580 33.385 3.630 ;
        RECT 33.835 3.210 34.005 3.630 ;
        RECT 38.705 3.485 39.005 3.905 ;
        RECT 40.025 3.575 40.275 4.425 ;
        RECT 39.485 3.305 40.275 3.575 ;
        RECT 40.445 3.725 40.855 4.245 ;
        RECT 41.025 3.995 41.255 4.425 ;
        RECT 41.425 3.735 41.595 4.765 ;
        RECT 41.765 4.365 42.025 4.815 ;
        RECT 42.695 4.635 43.455 4.885 ;
        RECT 43.625 4.765 43.895 5.465 ;
        RECT 42.685 4.605 43.455 4.635 ;
        RECT 42.665 4.595 43.455 4.605 ;
        RECT 42.665 4.575 43.555 4.595 ;
        RECT 42.645 4.565 43.555 4.575 ;
        RECT 42.625 4.555 43.555 4.565 ;
        RECT 42.595 4.545 43.555 4.555 ;
        RECT 42.525 4.515 43.555 4.545 ;
        RECT 42.505 4.485 43.555 4.515 ;
        RECT 42.485 4.455 43.555 4.485 ;
        RECT 42.455 4.425 43.555 4.455 ;
        RECT 42.425 4.395 43.555 4.425 ;
        RECT 42.395 4.385 43.555 4.395 ;
        RECT 42.395 4.375 42.755 4.385 ;
        RECT 42.395 4.365 42.745 4.375 ;
        RECT 41.765 4.355 42.725 4.365 ;
        RECT 41.765 4.345 42.715 4.355 ;
        RECT 41.765 4.325 42.695 4.345 ;
        RECT 41.765 4.315 42.685 4.325 ;
        RECT 41.765 4.195 42.655 4.315 ;
        RECT 40.445 3.305 40.645 3.725 ;
        RECT 41.335 3.265 41.595 3.735 ;
        RECT 41.765 3.635 42.315 4.025 ;
        RECT 42.485 3.465 42.655 4.195 ;
        RECT 41.765 3.295 42.655 3.465 ;
        RECT 42.825 3.795 43.155 4.215 ;
        RECT 43.325 3.995 43.555 4.385 ;
        RECT 43.725 4.275 43.895 4.765 ;
        RECT 44.075 4.665 44.405 5.455 ;
        RECT 44.075 4.495 44.755 4.665 ;
        RECT 44.065 4.275 44.415 4.325 ;
        RECT 43.725 4.105 44.415 4.275 ;
        RECT 42.825 3.305 43.045 3.795 ;
        RECT 43.725 3.735 43.895 4.105 ;
        RECT 44.065 4.075 44.415 4.105 ;
        RECT 44.585 3.895 44.755 4.495 ;
        RECT 44.925 4.075 45.275 4.325 ;
        RECT 47.055 3.900 47.230 5.160 ;
        RECT 47.580 4.100 47.750 5.160 ;
        RECT 47.580 3.930 47.810 4.100 ;
        RECT 43.635 3.265 43.895 3.735 ;
        RECT 44.495 3.265 44.825 3.895 ;
        RECT 47.055 3.700 47.225 3.900 ;
        RECT 47.055 3.370 47.465 3.700 ;
        RECT 32.395 3.040 33.315 3.210 ;
        RECT 33.835 3.040 34.305 3.210 ;
        RECT 32.395 2.890 32.625 3.040 ;
        RECT 47.055 2.860 47.225 3.370 ;
        RECT 47.055 2.530 47.465 2.860 ;
        RECT 30.995 2.150 31.225 2.320 ;
        RECT 30.995 1.870 31.165 2.150 ;
        RECT 31.425 1.870 31.600 2.380 ;
        RECT 31.855 1.870 32.030 2.420 ;
        RECT 33.220 1.870 33.390 2.380 ;
        RECT 47.055 2.360 47.225 2.530 ;
        RECT 47.055 1.870 47.230 2.360 ;
        RECT 47.640 2.320 47.810 3.930 ;
        RECT 48.010 3.900 48.185 5.160 ;
        RECT 48.440 4.020 48.615 5.160 ;
        RECT 48.010 2.950 48.180 3.900 ;
        RECT 48.440 2.420 48.610 4.020 ;
        RECT 49.800 4.015 49.975 5.160 ;
        RECT 55.345 5.130 55.515 5.470 ;
        RECT 56.840 5.130 57.310 5.470 ;
        RECT 55.340 5.070 55.515 5.130 ;
        RECT 54.830 4.080 55.170 4.960 ;
        RECT 55.340 4.250 55.510 5.070 ;
        RECT 56.050 4.600 56.300 4.970 ;
        RECT 57.020 4.600 57.740 4.900 ;
        RECT 57.910 4.770 58.180 5.470 ;
        RECT 59.130 5.130 59.610 5.470 ;
        RECT 56.050 4.430 57.840 4.600 ;
        RECT 49.430 3.210 49.600 3.900 ;
        RECT 49.800 3.800 49.970 4.015 ;
        RECT 55.340 4.000 56.440 4.250 ;
        RECT 55.340 3.910 55.590 4.000 ;
        RECT 50.420 3.800 50.590 3.900 ;
        RECT 49.800 3.630 50.590 3.800 ;
        RECT 49.800 3.580 49.970 3.630 ;
        RECT 50.420 3.210 50.590 3.630 ;
        RECT 55.290 3.490 55.590 3.910 ;
        RECT 56.610 3.580 56.860 4.430 ;
        RECT 56.070 3.310 56.860 3.580 ;
        RECT 57.030 3.730 57.440 4.250 ;
        RECT 57.610 4.000 57.840 4.430 ;
        RECT 58.010 3.740 58.180 4.770 ;
        RECT 58.350 4.370 58.610 4.820 ;
        RECT 59.280 4.640 60.040 4.890 ;
        RECT 60.210 4.770 60.480 5.470 ;
        RECT 59.270 4.610 60.040 4.640 ;
        RECT 59.250 4.600 60.040 4.610 ;
        RECT 59.250 4.580 60.140 4.600 ;
        RECT 59.230 4.570 60.140 4.580 ;
        RECT 59.210 4.560 60.140 4.570 ;
        RECT 59.180 4.550 60.140 4.560 ;
        RECT 59.110 4.520 60.140 4.550 ;
        RECT 59.090 4.490 60.140 4.520 ;
        RECT 59.070 4.460 60.140 4.490 ;
        RECT 59.040 4.430 60.140 4.460 ;
        RECT 59.010 4.400 60.140 4.430 ;
        RECT 58.980 4.390 60.140 4.400 ;
        RECT 58.980 4.380 59.340 4.390 ;
        RECT 58.980 4.370 59.330 4.380 ;
        RECT 58.350 4.360 59.310 4.370 ;
        RECT 58.350 4.350 59.300 4.360 ;
        RECT 58.350 4.330 59.280 4.350 ;
        RECT 58.350 4.320 59.270 4.330 ;
        RECT 58.350 4.200 59.240 4.320 ;
        RECT 57.030 3.310 57.230 3.730 ;
        RECT 57.920 3.270 58.180 3.740 ;
        RECT 58.350 3.640 58.900 4.030 ;
        RECT 59.070 3.470 59.240 4.200 ;
        RECT 58.350 3.300 59.240 3.470 ;
        RECT 59.410 3.800 59.740 4.220 ;
        RECT 59.910 4.000 60.140 4.390 ;
        RECT 60.310 4.280 60.480 4.770 ;
        RECT 60.660 4.670 60.990 5.460 ;
        RECT 60.660 4.500 61.340 4.670 ;
        RECT 60.650 4.280 61.000 4.330 ;
        RECT 60.310 4.110 61.000 4.280 ;
        RECT 59.410 3.310 59.630 3.800 ;
        RECT 60.310 3.740 60.480 4.110 ;
        RECT 60.650 4.080 61.000 4.110 ;
        RECT 61.170 3.900 61.340 4.500 ;
        RECT 61.510 4.080 61.860 4.330 ;
        RECT 63.640 3.905 63.815 5.165 ;
        RECT 64.165 4.105 64.335 5.165 ;
        RECT 64.165 3.935 64.395 4.105 ;
        RECT 60.220 3.270 60.480 3.740 ;
        RECT 61.080 3.270 61.410 3.900 ;
        RECT 63.640 3.705 63.810 3.905 ;
        RECT 63.640 3.375 64.050 3.705 ;
        RECT 48.980 3.040 49.900 3.210 ;
        RECT 50.420 3.040 50.890 3.210 ;
        RECT 48.980 2.890 49.210 3.040 ;
        RECT 63.640 2.865 63.810 3.375 ;
        RECT 63.640 2.535 64.050 2.865 ;
        RECT 47.580 2.150 47.810 2.320 ;
        RECT 47.580 1.870 47.750 2.150 ;
        RECT 48.010 1.870 48.185 2.380 ;
        RECT 48.440 1.870 48.615 2.420 ;
        RECT 49.805 1.870 49.975 2.380 ;
        RECT 63.640 2.365 63.810 2.535 ;
        RECT 63.640 1.875 63.815 2.365 ;
        RECT 64.225 2.325 64.395 3.935 ;
        RECT 64.595 3.905 64.770 5.165 ;
        RECT 65.025 4.025 65.200 5.165 ;
        RECT 64.595 2.955 64.765 3.905 ;
        RECT 65.025 2.425 65.195 4.025 ;
        RECT 66.385 4.020 66.560 5.165 ;
        RECT 71.930 5.135 72.100 5.475 ;
        RECT 73.425 5.135 73.895 5.475 ;
        RECT 71.925 5.075 72.100 5.135 ;
        RECT 71.415 4.085 71.755 4.965 ;
        RECT 71.925 4.255 72.095 5.075 ;
        RECT 72.635 4.605 72.885 4.975 ;
        RECT 73.605 4.605 74.325 4.905 ;
        RECT 74.495 4.775 74.765 5.475 ;
        RECT 75.715 5.135 76.195 5.475 ;
        RECT 72.635 4.435 74.425 4.605 ;
        RECT 66.015 3.215 66.185 3.905 ;
        RECT 66.385 3.805 66.555 4.020 ;
        RECT 71.925 4.005 73.025 4.255 ;
        RECT 71.925 3.915 72.175 4.005 ;
        RECT 67.005 3.805 67.175 3.905 ;
        RECT 66.385 3.635 67.175 3.805 ;
        RECT 66.385 3.585 66.555 3.635 ;
        RECT 67.005 3.215 67.175 3.635 ;
        RECT 71.875 3.495 72.175 3.915 ;
        RECT 73.195 3.585 73.445 4.435 ;
        RECT 72.655 3.315 73.445 3.585 ;
        RECT 73.615 3.735 74.025 4.255 ;
        RECT 74.195 4.005 74.425 4.435 ;
        RECT 74.595 3.745 74.765 4.775 ;
        RECT 74.935 4.375 75.195 4.825 ;
        RECT 75.865 4.645 76.625 4.895 ;
        RECT 76.795 4.775 77.065 5.475 ;
        RECT 75.855 4.615 76.625 4.645 ;
        RECT 75.835 4.605 76.625 4.615 ;
        RECT 75.835 4.585 76.725 4.605 ;
        RECT 75.815 4.575 76.725 4.585 ;
        RECT 75.795 4.565 76.725 4.575 ;
        RECT 75.765 4.555 76.725 4.565 ;
        RECT 75.695 4.525 76.725 4.555 ;
        RECT 75.675 4.495 76.725 4.525 ;
        RECT 75.655 4.465 76.725 4.495 ;
        RECT 75.625 4.435 76.725 4.465 ;
        RECT 75.595 4.405 76.725 4.435 ;
        RECT 75.565 4.395 76.725 4.405 ;
        RECT 75.565 4.385 75.925 4.395 ;
        RECT 75.565 4.375 75.915 4.385 ;
        RECT 74.935 4.365 75.895 4.375 ;
        RECT 74.935 4.355 75.885 4.365 ;
        RECT 74.935 4.335 75.865 4.355 ;
        RECT 74.935 4.325 75.855 4.335 ;
        RECT 74.935 4.205 75.825 4.325 ;
        RECT 73.615 3.315 73.815 3.735 ;
        RECT 74.505 3.275 74.765 3.745 ;
        RECT 74.935 3.645 75.485 4.035 ;
        RECT 75.655 3.475 75.825 4.205 ;
        RECT 74.935 3.305 75.825 3.475 ;
        RECT 75.995 3.805 76.325 4.225 ;
        RECT 76.495 4.005 76.725 4.395 ;
        RECT 76.895 4.285 77.065 4.775 ;
        RECT 77.245 4.675 77.575 5.465 ;
        RECT 77.245 4.505 77.925 4.675 ;
        RECT 77.235 4.285 77.585 4.335 ;
        RECT 76.895 4.115 77.585 4.285 ;
        RECT 75.995 3.315 76.215 3.805 ;
        RECT 76.895 3.745 77.065 4.115 ;
        RECT 77.235 4.085 77.585 4.115 ;
        RECT 77.755 3.905 77.925 4.505 ;
        RECT 78.095 4.085 78.445 4.335 ;
        RECT 80.225 3.910 80.400 5.170 ;
        RECT 80.750 4.110 80.920 5.170 ;
        RECT 80.750 3.940 80.980 4.110 ;
        RECT 76.805 3.275 77.065 3.745 ;
        RECT 77.665 3.275 77.995 3.905 ;
        RECT 80.225 3.710 80.395 3.910 ;
        RECT 80.225 3.380 80.635 3.710 ;
        RECT 65.565 3.045 66.485 3.215 ;
        RECT 67.005 3.045 67.475 3.215 ;
        RECT 65.565 2.895 65.795 3.045 ;
        RECT 80.225 2.870 80.395 3.380 ;
        RECT 80.225 2.540 80.635 2.870 ;
        RECT 64.165 2.155 64.395 2.325 ;
        RECT 64.165 1.875 64.335 2.155 ;
        RECT 64.595 1.875 64.770 2.385 ;
        RECT 65.025 1.875 65.200 2.425 ;
        RECT 66.390 1.875 66.560 2.385 ;
        RECT 80.225 2.370 80.395 2.540 ;
        RECT 80.225 1.880 80.400 2.370 ;
        RECT 80.810 2.330 80.980 3.940 ;
        RECT 81.180 3.910 81.355 5.170 ;
        RECT 81.610 4.030 81.785 5.170 ;
        RECT 81.180 2.960 81.350 3.910 ;
        RECT 81.610 2.430 81.780 4.030 ;
        RECT 82.970 4.025 83.145 5.170 ;
        RECT 88.510 5.135 88.680 5.475 ;
        RECT 90.005 5.135 90.475 5.475 ;
        RECT 88.505 5.075 88.680 5.135 ;
        RECT 87.995 4.085 88.335 4.965 ;
        RECT 88.505 4.255 88.675 5.075 ;
        RECT 89.215 4.605 89.465 4.975 ;
        RECT 90.185 4.605 90.905 4.905 ;
        RECT 91.075 4.775 91.345 5.475 ;
        RECT 92.295 5.135 92.775 5.475 ;
        RECT 89.215 4.435 91.005 4.605 ;
        RECT 82.600 3.220 82.770 3.910 ;
        RECT 82.970 3.810 83.140 4.025 ;
        RECT 88.505 4.005 89.605 4.255 ;
        RECT 88.505 3.915 88.755 4.005 ;
        RECT 83.590 3.810 83.760 3.910 ;
        RECT 82.970 3.640 83.760 3.810 ;
        RECT 82.970 3.590 83.140 3.640 ;
        RECT 83.590 3.220 83.760 3.640 ;
        RECT 88.455 3.495 88.755 3.915 ;
        RECT 89.775 3.585 90.025 4.435 ;
        RECT 89.235 3.315 90.025 3.585 ;
        RECT 90.195 3.735 90.605 4.255 ;
        RECT 90.775 4.005 91.005 4.435 ;
        RECT 91.175 3.745 91.345 4.775 ;
        RECT 91.515 4.375 91.775 4.825 ;
        RECT 92.445 4.645 93.205 4.895 ;
        RECT 93.375 4.775 93.645 5.475 ;
        RECT 92.435 4.615 93.205 4.645 ;
        RECT 92.415 4.605 93.205 4.615 ;
        RECT 92.415 4.585 93.305 4.605 ;
        RECT 92.395 4.575 93.305 4.585 ;
        RECT 92.375 4.565 93.305 4.575 ;
        RECT 92.345 4.555 93.305 4.565 ;
        RECT 92.275 4.525 93.305 4.555 ;
        RECT 92.255 4.495 93.305 4.525 ;
        RECT 92.235 4.465 93.305 4.495 ;
        RECT 92.205 4.435 93.305 4.465 ;
        RECT 92.175 4.405 93.305 4.435 ;
        RECT 92.145 4.395 93.305 4.405 ;
        RECT 92.145 4.385 92.505 4.395 ;
        RECT 92.145 4.375 92.495 4.385 ;
        RECT 91.515 4.365 92.475 4.375 ;
        RECT 91.515 4.355 92.465 4.365 ;
        RECT 91.515 4.335 92.445 4.355 ;
        RECT 91.515 4.325 92.435 4.335 ;
        RECT 91.515 4.205 92.405 4.325 ;
        RECT 90.195 3.315 90.395 3.735 ;
        RECT 91.085 3.275 91.345 3.745 ;
        RECT 91.515 3.645 92.065 4.035 ;
        RECT 92.235 3.475 92.405 4.205 ;
        RECT 91.515 3.305 92.405 3.475 ;
        RECT 92.575 3.805 92.905 4.225 ;
        RECT 93.075 4.005 93.305 4.395 ;
        RECT 93.475 4.285 93.645 4.775 ;
        RECT 93.825 4.675 94.155 5.465 ;
        RECT 93.825 4.505 94.505 4.675 ;
        RECT 93.815 4.285 94.165 4.335 ;
        RECT 93.475 4.115 94.165 4.285 ;
        RECT 92.575 3.315 92.795 3.805 ;
        RECT 93.475 3.745 93.645 4.115 ;
        RECT 93.815 4.085 94.165 4.115 ;
        RECT 94.335 3.905 94.505 4.505 ;
        RECT 94.675 4.085 95.025 4.335 ;
        RECT 96.805 3.910 96.980 5.170 ;
        RECT 97.330 4.110 97.500 5.170 ;
        RECT 97.330 3.940 97.560 4.110 ;
        RECT 93.385 3.275 93.645 3.745 ;
        RECT 94.245 3.275 94.575 3.905 ;
        RECT 96.805 3.710 96.975 3.910 ;
        RECT 96.805 3.380 97.215 3.710 ;
        RECT 82.150 3.050 83.070 3.220 ;
        RECT 83.590 3.050 84.060 3.220 ;
        RECT 82.150 2.900 82.380 3.050 ;
        RECT 96.805 2.870 96.975 3.380 ;
        RECT 96.805 2.540 97.215 2.870 ;
        RECT 80.750 2.160 80.980 2.330 ;
        RECT 80.750 1.880 80.920 2.160 ;
        RECT 81.180 1.880 81.355 2.390 ;
        RECT 81.610 1.880 81.785 2.430 ;
        RECT 82.975 1.880 83.145 2.390 ;
        RECT 96.805 2.370 96.975 2.540 ;
        RECT 96.805 1.880 96.980 2.370 ;
        RECT 97.390 2.330 97.560 3.940 ;
        RECT 97.760 3.910 97.935 5.170 ;
        RECT 98.190 4.030 98.365 5.170 ;
        RECT 97.760 2.960 97.930 3.910 ;
        RECT 98.190 2.430 98.360 4.030 ;
        RECT 99.550 4.025 99.725 5.170 ;
        RECT 99.180 3.220 99.350 3.910 ;
        RECT 99.550 3.810 99.720 4.025 ;
        RECT 100.170 3.810 100.340 3.910 ;
        RECT 99.550 3.640 100.340 3.810 ;
        RECT 99.550 3.590 99.720 3.640 ;
        RECT 100.170 3.220 100.340 3.640 ;
        RECT 98.730 3.050 99.650 3.220 ;
        RECT 100.170 3.050 100.640 3.220 ;
        RECT 98.730 2.900 98.960 3.050 ;
        RECT 97.330 2.160 97.560 2.330 ;
        RECT 97.330 1.880 97.500 2.160 ;
        RECT 97.760 1.880 97.935 2.390 ;
        RECT 98.190 1.880 98.365 2.430 ;
        RECT 99.555 1.880 99.725 2.390 ;
      LAYER met1 ;
        RECT 16.910 10.045 17.200 10.275 ;
        RECT 20.140 10.045 20.430 10.275 ;
        RECT 31.365 10.050 31.655 10.280 ;
        RECT 16.970 9.590 17.140 10.045 ;
        RECT 20.200 9.675 20.370 10.045 ;
        RECT 16.890 9.310 17.230 9.590 ;
        RECT 16.910 9.305 17.200 9.310 ;
        RECT 20.100 9.305 20.470 9.675 ;
        RECT 31.425 9.575 31.595 10.050 ;
        RECT 33.155 10.020 33.450 10.280 ;
        RECT 34.145 10.020 34.440 10.280 ;
        RECT 36.725 10.045 37.015 10.275 ;
        RECT 47.950 10.050 48.240 10.280 ;
        RECT 32.335 9.575 32.685 9.600 ;
        RECT 31.425 9.540 32.685 9.575 ;
        RECT 31.365 9.405 32.685 9.540 ;
        RECT 31.365 9.310 31.655 9.405 ;
        RECT 32.335 9.310 32.685 9.405 ;
        RECT 20.600 9.165 20.940 9.195 ;
        RECT 31.820 9.170 32.145 9.265 ;
        RECT 20.570 9.135 20.940 9.165 ;
        RECT 31.795 9.140 32.145 9.170 ;
        RECT 20.400 8.965 20.940 9.135 ;
        RECT 31.625 8.970 32.145 9.140 ;
        RECT 20.570 8.935 20.940 8.965 ;
        RECT 31.795 8.940 32.145 8.970 ;
        RECT 20.600 8.915 20.940 8.935 ;
        RECT 33.215 8.920 33.385 10.020 ;
        RECT 34.205 9.270 34.375 10.020 ;
        RECT 36.785 9.675 36.955 10.045 ;
        RECT 36.685 9.305 37.055 9.675 ;
        RECT 48.010 9.575 48.180 10.050 ;
        RECT 49.740 10.020 50.035 10.280 ;
        RECT 50.730 10.020 51.025 10.280 ;
        RECT 53.310 10.050 53.600 10.280 ;
        RECT 64.535 10.055 64.825 10.285 ;
        RECT 48.920 9.575 49.270 9.600 ;
        RECT 48.010 9.540 49.270 9.575 ;
        RECT 47.950 9.405 49.270 9.540 ;
        RECT 47.950 9.310 48.240 9.405 ;
        RECT 48.920 9.310 49.270 9.405 ;
        RECT 34.205 8.945 34.535 9.270 ;
        RECT 37.185 9.165 37.525 9.195 ;
        RECT 48.405 9.170 48.730 9.265 ;
        RECT 37.155 9.135 37.525 9.165 ;
        RECT 48.380 9.140 48.730 9.170 ;
        RECT 36.985 8.965 37.525 9.135 ;
        RECT 48.210 8.970 48.730 9.140 ;
        RECT 34.205 8.920 34.495 8.945 ;
        RECT 37.155 8.935 37.525 8.965 ;
        RECT 48.380 8.940 48.730 8.970 ;
        RECT 33.155 8.915 33.385 8.920 ;
        RECT 16.505 8.775 16.845 8.850 ;
        RECT 31.020 8.810 31.340 8.890 ;
        RECT 30.995 8.780 31.340 8.810 ;
        RECT 16.365 8.605 16.845 8.775 ;
        RECT 30.820 8.610 31.340 8.780 ;
        RECT 33.155 8.680 33.445 8.915 ;
        RECT 34.145 8.805 34.495 8.920 ;
        RECT 37.185 8.915 37.525 8.935 ;
        RECT 49.800 8.920 49.970 10.020 ;
        RECT 50.790 9.270 50.960 10.020 ;
        RECT 53.370 9.680 53.540 10.050 ;
        RECT 53.270 9.310 53.640 9.680 ;
        RECT 64.595 9.580 64.765 10.055 ;
        RECT 66.325 10.025 66.620 10.285 ;
        RECT 67.315 10.025 67.610 10.285 ;
        RECT 69.895 10.055 70.185 10.285 ;
        RECT 81.120 10.060 81.410 10.290 ;
        RECT 65.505 9.580 65.855 9.605 ;
        RECT 64.595 9.545 65.855 9.580 ;
        RECT 64.535 9.410 65.855 9.545 ;
        RECT 64.535 9.315 64.825 9.410 ;
        RECT 65.505 9.315 65.855 9.410 ;
        RECT 50.790 8.945 51.120 9.270 ;
        RECT 53.800 9.200 54.080 9.230 ;
        RECT 53.770 9.170 54.110 9.200 ;
        RECT 64.990 9.175 65.315 9.270 ;
        RECT 53.740 9.140 54.110 9.170 ;
        RECT 64.965 9.145 65.315 9.175 ;
        RECT 53.570 8.970 54.110 9.140 ;
        RECT 64.795 8.975 65.315 9.145 ;
        RECT 50.790 8.920 51.080 8.945 ;
        RECT 49.740 8.915 49.970 8.920 ;
        RECT 47.605 8.810 47.925 8.890 ;
        RECT 34.145 8.680 34.435 8.805 ;
        RECT 47.580 8.780 47.925 8.810 ;
        RECT 47.405 8.610 47.925 8.780 ;
        RECT 49.740 8.680 50.030 8.915 ;
        RECT 50.730 8.815 51.080 8.920 ;
        RECT 53.740 8.885 54.110 8.970 ;
        RECT 64.965 8.945 65.315 8.975 ;
        RECT 66.385 8.925 66.555 10.025 ;
        RECT 67.375 9.275 67.545 10.025 ;
        RECT 69.955 9.685 70.125 10.055 ;
        RECT 69.855 9.315 70.225 9.685 ;
        RECT 81.180 9.585 81.350 10.060 ;
        RECT 82.910 10.030 83.205 10.290 ;
        RECT 83.900 10.030 84.195 10.290 ;
        RECT 86.475 10.055 86.765 10.285 ;
        RECT 97.700 10.060 97.990 10.290 ;
        RECT 82.090 9.585 82.440 9.610 ;
        RECT 81.180 9.550 82.440 9.585 ;
        RECT 81.120 9.415 82.440 9.550 ;
        RECT 81.120 9.320 81.410 9.415 ;
        RECT 82.090 9.320 82.440 9.415 ;
        RECT 67.375 8.950 67.705 9.275 ;
        RECT 70.355 9.175 70.695 9.205 ;
        RECT 81.575 9.180 81.900 9.275 ;
        RECT 70.325 9.145 70.695 9.175 ;
        RECT 81.550 9.150 81.900 9.180 ;
        RECT 70.155 8.975 70.695 9.145 ;
        RECT 81.380 8.980 81.900 9.150 ;
        RECT 67.375 8.925 67.665 8.950 ;
        RECT 70.325 8.945 70.695 8.975 ;
        RECT 81.550 8.950 81.900 8.980 ;
        RECT 70.355 8.925 70.695 8.945 ;
        RECT 82.970 8.930 83.140 10.030 ;
        RECT 83.960 9.280 84.130 10.030 ;
        RECT 86.535 9.685 86.705 10.055 ;
        RECT 86.435 9.315 86.805 9.685 ;
        RECT 97.760 9.585 97.930 10.060 ;
        RECT 99.490 10.030 99.785 10.290 ;
        RECT 100.480 10.030 100.775 10.290 ;
        RECT 98.670 9.585 99.020 9.610 ;
        RECT 97.760 9.550 99.020 9.585 ;
        RECT 97.700 9.415 99.020 9.550 ;
        RECT 97.700 9.320 97.990 9.415 ;
        RECT 98.670 9.320 99.020 9.415 ;
        RECT 83.960 8.955 84.290 9.280 ;
        RECT 86.935 9.175 87.275 9.205 ;
        RECT 98.155 9.180 98.480 9.275 ;
        RECT 86.905 9.145 87.275 9.175 ;
        RECT 98.130 9.150 98.480 9.180 ;
        RECT 86.735 8.975 87.275 9.145 ;
        RECT 97.960 8.980 98.480 9.150 ;
        RECT 83.960 8.930 84.250 8.955 ;
        RECT 86.905 8.945 87.275 8.975 ;
        RECT 98.130 8.950 98.480 8.980 ;
        RECT 82.910 8.925 83.140 8.930 ;
        RECT 66.325 8.920 66.555 8.925 ;
        RECT 64.190 8.815 64.510 8.895 ;
        RECT 50.730 8.680 51.020 8.815 ;
        RECT 64.165 8.785 64.510 8.815 ;
        RECT 63.990 8.615 64.510 8.785 ;
        RECT 66.325 8.685 66.615 8.920 ;
        RECT 67.315 8.820 67.665 8.925 ;
        RECT 80.775 8.820 81.095 8.900 ;
        RECT 67.315 8.685 67.605 8.820 ;
        RECT 80.750 8.790 81.095 8.820 ;
        RECT 80.575 8.620 81.095 8.790 ;
        RECT 82.910 8.690 83.200 8.925 ;
        RECT 83.900 8.815 84.250 8.930 ;
        RECT 86.935 8.925 87.275 8.945 ;
        RECT 99.550 8.930 99.720 10.030 ;
        RECT 100.510 10.000 100.775 10.030 ;
        RECT 100.510 9.585 100.835 10.000 ;
        RECT 100.540 8.930 100.710 9.585 ;
        RECT 99.490 8.925 99.720 8.930 ;
        RECT 100.480 8.925 100.710 8.930 ;
        RECT 97.355 8.820 97.675 8.900 ;
        RECT 83.900 8.690 84.190 8.815 ;
        RECT 97.330 8.790 97.675 8.820 ;
        RECT 97.155 8.620 97.675 8.790 ;
        RECT 99.490 8.690 99.780 8.925 ;
        RECT 100.480 8.690 100.770 8.925 ;
        RECT 16.505 8.570 16.845 8.605 ;
        RECT 30.995 8.580 31.340 8.610 ;
        RECT 47.580 8.580 47.925 8.610 ;
        RECT 64.165 8.585 64.510 8.615 ;
        RECT 80.750 8.590 81.095 8.620 ;
        RECT 97.330 8.590 97.675 8.620 ;
        RECT 31.020 8.565 31.340 8.580 ;
        RECT 47.605 8.565 47.925 8.580 ;
        RECT 64.190 8.570 64.510 8.585 ;
        RECT 80.775 8.575 81.095 8.590 ;
        RECT 97.355 8.575 97.675 8.590 ;
        RECT 24.280 7.325 24.570 7.365 ;
        RECT 24.950 7.325 25.270 7.385 ;
        RECT 24.280 7.185 25.270 7.325 ;
        RECT 24.280 7.135 24.570 7.185 ;
        RECT 24.950 7.125 25.270 7.185 ;
        RECT 25.970 7.125 26.290 7.385 ;
        RECT 26.660 7.135 26.950 7.365 ;
        RECT 27.330 7.325 27.650 7.385 ;
        RECT 40.865 7.325 41.155 7.365 ;
        RECT 41.535 7.325 41.855 7.385 ;
        RECT 27.330 7.185 27.920 7.325 ;
        RECT 40.865 7.185 41.855 7.325 ;
        RECT 25.040 6.985 25.180 7.125 ;
        RECT 26.740 6.985 26.880 7.135 ;
        RECT 27.330 7.125 27.650 7.185 ;
        RECT 40.865 7.135 41.155 7.185 ;
        RECT 41.535 7.125 41.855 7.185 ;
        RECT 42.555 7.125 42.875 7.385 ;
        RECT 43.245 7.135 43.535 7.365 ;
        RECT 43.915 7.325 44.235 7.385 ;
        RECT 57.450 7.330 57.740 7.370 ;
        RECT 58.120 7.330 58.440 7.390 ;
        RECT 43.915 7.185 44.505 7.325 ;
        RECT 57.450 7.190 58.440 7.330 ;
        RECT 25.040 6.845 26.880 6.985 ;
        RECT 41.625 6.985 41.765 7.125 ;
        RECT 43.325 6.985 43.465 7.135 ;
        RECT 43.915 7.125 44.235 7.185 ;
        RECT 57.450 7.140 57.740 7.190 ;
        RECT 58.120 7.130 58.440 7.190 ;
        RECT 59.140 7.130 59.460 7.390 ;
        RECT 59.830 7.140 60.120 7.370 ;
        RECT 60.500 7.330 60.820 7.390 ;
        RECT 74.035 7.335 74.325 7.375 ;
        RECT 74.705 7.335 75.025 7.395 ;
        RECT 60.500 7.190 61.090 7.330 ;
        RECT 74.035 7.195 75.025 7.335 ;
        RECT 41.625 6.845 43.465 6.985 ;
        RECT 58.210 6.990 58.350 7.130 ;
        RECT 59.910 6.990 60.050 7.140 ;
        RECT 60.500 7.130 60.820 7.190 ;
        RECT 74.035 7.145 74.325 7.195 ;
        RECT 74.705 7.135 75.025 7.195 ;
        RECT 75.725 7.135 76.045 7.395 ;
        RECT 76.415 7.145 76.705 7.375 ;
        RECT 77.085 7.335 77.405 7.395 ;
        RECT 90.615 7.335 90.905 7.375 ;
        RECT 91.285 7.335 91.605 7.395 ;
        RECT 77.085 7.195 77.675 7.335 ;
        RECT 90.615 7.195 91.605 7.335 ;
        RECT 58.210 6.850 60.050 6.990 ;
        RECT 74.795 6.995 74.935 7.135 ;
        RECT 76.495 6.995 76.635 7.145 ;
        RECT 77.085 7.135 77.405 7.195 ;
        RECT 90.615 7.145 90.905 7.195 ;
        RECT 91.285 7.135 91.605 7.195 ;
        RECT 92.305 7.135 92.625 7.395 ;
        RECT 92.995 7.145 93.285 7.375 ;
        RECT 93.665 7.335 93.985 7.395 ;
        RECT 93.665 7.195 94.255 7.335 ;
        RECT 74.795 6.855 76.635 6.995 ;
        RECT 91.375 6.995 91.515 7.135 ;
        RECT 93.075 6.995 93.215 7.145 ;
        RECT 93.665 7.135 93.985 7.195 ;
        RECT 91.375 6.855 93.215 6.995 ;
        RECT 22.580 6.305 22.870 6.345 ;
        RECT 25.290 6.305 25.610 6.365 ;
        RECT 22.580 6.165 25.610 6.305 ;
        RECT 22.580 6.115 22.870 6.165 ;
        RECT 25.290 6.105 25.610 6.165 ;
        RECT 28.020 6.105 28.670 6.365 ;
        RECT 39.165 6.305 39.455 6.345 ;
        RECT 41.875 6.305 42.195 6.365 ;
        RECT 39.165 6.165 42.195 6.305 ;
        RECT 39.165 6.115 39.455 6.165 ;
        RECT 41.875 6.105 42.195 6.165 ;
        RECT 44.605 6.105 45.255 6.365 ;
        RECT 55.750 6.310 56.040 6.350 ;
        RECT 58.460 6.310 58.780 6.370 ;
        RECT 55.750 6.170 58.780 6.310 ;
        RECT 55.750 6.120 56.040 6.170 ;
        RECT 58.460 6.110 58.780 6.170 ;
        RECT 61.190 6.110 61.840 6.370 ;
        RECT 72.335 6.315 72.625 6.355 ;
        RECT 75.045 6.315 75.365 6.375 ;
        RECT 72.335 6.175 75.365 6.315 ;
        RECT 72.335 6.125 72.625 6.175 ;
        RECT 75.045 6.115 75.365 6.175 ;
        RECT 77.775 6.115 78.425 6.375 ;
        RECT 88.915 6.315 89.205 6.355 ;
        RECT 91.625 6.315 91.945 6.375 ;
        RECT 88.915 6.175 91.945 6.315 ;
        RECT 88.915 6.125 89.205 6.175 ;
        RECT 91.625 6.115 91.945 6.175 ;
        RECT 94.355 6.115 95.005 6.375 ;
        RECT 23.770 5.285 24.060 5.325 ;
        RECT 25.980 5.285 26.270 5.325 ;
        RECT 26.650 5.285 26.970 5.345 ;
        RECT 23.770 5.145 26.970 5.285 ;
        RECT 23.770 5.095 24.060 5.145 ;
        RECT 25.980 5.095 26.270 5.145 ;
        RECT 26.650 5.085 26.970 5.145 ;
        RECT 40.355 5.285 40.645 5.325 ;
        RECT 42.565 5.285 42.855 5.325 ;
        RECT 43.235 5.285 43.555 5.345 ;
        RECT 40.355 5.145 43.555 5.285 ;
        RECT 40.355 5.095 40.645 5.145 ;
        RECT 42.565 5.095 42.855 5.145 ;
        RECT 43.235 5.085 43.555 5.145 ;
        RECT 56.940 5.290 57.230 5.330 ;
        RECT 59.150 5.290 59.440 5.330 ;
        RECT 59.820 5.290 60.140 5.350 ;
        RECT 56.940 5.150 60.140 5.290 ;
        RECT 56.940 5.100 57.230 5.150 ;
        RECT 59.150 5.100 59.440 5.150 ;
        RECT 59.820 5.090 60.140 5.150 ;
        RECT 73.525 5.295 73.815 5.335 ;
        RECT 75.735 5.295 76.025 5.335 ;
        RECT 76.405 5.295 76.725 5.355 ;
        RECT 73.525 5.155 76.725 5.295 ;
        RECT 73.525 5.105 73.815 5.155 ;
        RECT 75.735 5.105 76.025 5.155 ;
        RECT 76.405 5.095 76.725 5.155 ;
        RECT 90.105 5.295 90.395 5.335 ;
        RECT 92.315 5.295 92.605 5.335 ;
        RECT 92.985 5.295 93.305 5.355 ;
        RECT 90.105 5.155 93.305 5.295 ;
        RECT 90.105 5.105 90.395 5.155 ;
        RECT 92.315 5.105 92.605 5.155 ;
        RECT 92.985 5.095 93.305 5.155 ;
        RECT 25.970 4.605 26.290 4.665 ;
        RECT 27.940 4.605 28.230 4.645 ;
        RECT 42.555 4.605 42.875 4.665 ;
        RECT 44.525 4.605 44.815 4.645 ;
        RECT 59.140 4.610 59.460 4.670 ;
        RECT 61.110 4.610 61.400 4.650 ;
        RECT 75.725 4.615 76.045 4.675 ;
        RECT 77.695 4.615 77.985 4.655 ;
        RECT 92.305 4.615 92.625 4.675 ;
        RECT 94.275 4.615 94.565 4.655 ;
        RECT 25.970 4.465 28.235 4.605 ;
        RECT 42.555 4.465 44.820 4.605 ;
        RECT 59.140 4.470 61.405 4.610 ;
        RECT 75.725 4.475 77.990 4.615 ;
        RECT 92.305 4.475 94.570 4.615 ;
        RECT 25.970 4.405 26.290 4.465 ;
        RECT 27.940 4.415 28.230 4.465 ;
        RECT 42.555 4.405 42.875 4.465 ;
        RECT 44.525 4.415 44.815 4.465 ;
        RECT 59.140 4.410 59.460 4.470 ;
        RECT 61.110 4.420 61.400 4.470 ;
        RECT 75.725 4.415 76.045 4.475 ;
        RECT 77.695 4.425 77.985 4.475 ;
        RECT 92.305 4.415 92.625 4.475 ;
        RECT 94.275 4.425 94.565 4.475 ;
        RECT 21.610 4.265 21.900 4.305 ;
        RECT 24.345 4.265 25.215 4.295 ;
        RECT 26.650 4.265 26.970 4.325 ;
        RECT 28.350 4.265 28.670 4.325 ;
        RECT 21.610 4.155 26.970 4.265 ;
        RECT 21.610 4.125 24.485 4.155 ;
        RECT 25.075 4.125 26.970 4.155 ;
        RECT 28.070 4.125 28.670 4.265 ;
        RECT 21.610 4.075 21.900 4.125 ;
        RECT 26.650 4.065 26.970 4.125 ;
        RECT 28.350 4.065 28.670 4.125 ;
        RECT 38.195 4.265 38.485 4.305 ;
        RECT 40.930 4.265 41.800 4.295 ;
        RECT 43.235 4.265 43.555 4.325 ;
        RECT 44.935 4.265 45.255 4.325 ;
        RECT 38.195 4.155 43.555 4.265 ;
        RECT 38.195 4.125 41.070 4.155 ;
        RECT 41.660 4.125 43.555 4.155 ;
        RECT 44.655 4.125 45.255 4.265 ;
        RECT 38.195 4.075 38.485 4.125 ;
        RECT 43.235 4.065 43.555 4.125 ;
        RECT 44.935 4.065 45.255 4.125 ;
        RECT 54.780 4.270 55.070 4.310 ;
        RECT 57.515 4.270 58.385 4.300 ;
        RECT 59.820 4.270 60.140 4.330 ;
        RECT 61.520 4.270 61.840 4.330 ;
        RECT 54.780 4.160 60.140 4.270 ;
        RECT 54.780 4.130 57.655 4.160 ;
        RECT 58.245 4.130 60.140 4.160 ;
        RECT 61.240 4.130 61.840 4.270 ;
        RECT 54.780 4.080 55.070 4.130 ;
        RECT 59.820 4.070 60.140 4.130 ;
        RECT 61.520 4.070 61.840 4.130 ;
        RECT 71.365 4.275 71.655 4.315 ;
        RECT 74.100 4.275 74.970 4.305 ;
        RECT 76.405 4.275 76.725 4.335 ;
        RECT 78.105 4.275 78.425 4.335 ;
        RECT 71.365 4.165 76.725 4.275 ;
        RECT 71.365 4.135 74.240 4.165 ;
        RECT 74.830 4.135 76.725 4.165 ;
        RECT 77.825 4.135 78.425 4.275 ;
        RECT 71.365 4.085 71.655 4.135 ;
        RECT 76.405 4.075 76.725 4.135 ;
        RECT 78.105 4.075 78.425 4.135 ;
        RECT 87.945 4.275 88.235 4.315 ;
        RECT 90.680 4.275 91.550 4.305 ;
        RECT 92.985 4.275 93.305 4.335 ;
        RECT 94.685 4.275 95.005 4.335 ;
        RECT 87.945 4.165 93.305 4.275 ;
        RECT 87.945 4.135 90.820 4.165 ;
        RECT 91.410 4.135 93.305 4.165 ;
        RECT 94.405 4.135 95.005 4.275 ;
        RECT 87.945 4.085 88.235 4.135 ;
        RECT 92.985 4.075 93.305 4.135 ;
        RECT 94.685 4.075 95.005 4.135 ;
        RECT 24.610 3.965 24.930 3.975 ;
        RECT 23.940 3.735 24.230 3.965 ;
        RECT 24.610 3.925 25.070 3.965 ;
        RECT 25.290 3.925 25.610 3.985 ;
        RECT 26.740 3.925 26.880 4.065 ;
        RECT 24.610 3.785 25.090 3.925 ;
        RECT 25.290 3.785 25.880 3.925 ;
        RECT 26.740 3.785 27.220 3.925 ;
        RECT 31.020 3.880 31.340 3.980 ;
        RECT 41.195 3.965 41.515 3.975 ;
        RECT 30.995 3.860 31.340 3.880 ;
        RECT 24.610 3.735 25.070 3.785 ;
        RECT 24.020 3.535 24.160 3.735 ;
        RECT 24.610 3.715 24.930 3.735 ;
        RECT 25.290 3.725 25.610 3.785 ;
        RECT 26.340 3.665 26.600 3.695 ;
        RECT 26.310 3.645 26.630 3.665 ;
        RECT 27.080 3.645 27.220 3.785 ;
        RECT 30.705 3.690 31.340 3.860 ;
        RECT 30.820 3.680 31.340 3.690 ;
        RECT 30.995 3.660 31.340 3.680 ;
        RECT 30.995 3.650 31.285 3.660 ;
        RECT 26.210 3.535 26.630 3.645 ;
        RECT 24.020 3.405 26.630 3.535 ;
        RECT 27.000 3.415 27.290 3.645 ;
        RECT 29.350 3.490 29.675 3.615 ;
        RECT 31.795 3.490 32.145 3.610 ;
        RECT 33.155 3.545 33.445 3.780 ;
        RECT 40.525 3.735 40.815 3.965 ;
        RECT 41.195 3.925 41.655 3.965 ;
        RECT 41.875 3.925 42.195 3.985 ;
        RECT 43.325 3.925 43.465 4.065 ;
        RECT 41.195 3.785 41.675 3.925 ;
        RECT 41.875 3.785 42.465 3.925 ;
        RECT 43.325 3.785 43.805 3.925 ;
        RECT 47.605 3.880 47.925 3.980 ;
        RECT 57.780 3.970 58.100 3.980 ;
        RECT 47.580 3.860 47.925 3.880 ;
        RECT 41.195 3.735 41.655 3.785 ;
        RECT 33.155 3.540 33.385 3.545 ;
        RECT 24.020 3.395 26.270 3.405 ;
        RECT 29.350 3.320 32.145 3.490 ;
        RECT 29.350 3.290 29.675 3.320 ;
        RECT 31.795 3.260 32.145 3.320 ;
        RECT 31.365 3.120 31.655 3.150 ;
        RECT 32.335 3.120 32.685 3.150 ;
        RECT 31.365 2.950 32.685 3.120 ;
        RECT 31.365 2.920 31.655 2.950 ;
        RECT 31.425 2.410 31.595 2.920 ;
        RECT 32.335 2.860 32.685 2.950 ;
        RECT 33.215 2.440 33.385 3.540 ;
        RECT 40.605 3.535 40.745 3.735 ;
        RECT 41.195 3.715 41.515 3.735 ;
        RECT 41.875 3.725 42.195 3.785 ;
        RECT 42.925 3.665 43.185 3.695 ;
        RECT 42.895 3.645 43.215 3.665 ;
        RECT 43.665 3.645 43.805 3.785 ;
        RECT 47.290 3.690 47.925 3.860 ;
        RECT 47.405 3.680 47.925 3.690 ;
        RECT 47.580 3.660 47.925 3.680 ;
        RECT 47.580 3.650 47.870 3.660 ;
        RECT 42.795 3.535 43.215 3.645 ;
        RECT 40.605 3.405 43.215 3.535 ;
        RECT 43.585 3.415 43.875 3.645 ;
        RECT 45.935 3.490 46.260 3.615 ;
        RECT 48.380 3.490 48.730 3.610 ;
        RECT 49.740 3.545 50.030 3.780 ;
        RECT 57.110 3.740 57.400 3.970 ;
        RECT 57.780 3.930 58.240 3.970 ;
        RECT 58.460 3.930 58.780 3.990 ;
        RECT 59.910 3.930 60.050 4.070 ;
        RECT 57.780 3.790 58.260 3.930 ;
        RECT 58.460 3.790 59.050 3.930 ;
        RECT 59.910 3.790 60.390 3.930 ;
        RECT 64.190 3.885 64.510 3.985 ;
        RECT 74.365 3.975 74.685 3.985 ;
        RECT 64.165 3.865 64.510 3.885 ;
        RECT 57.780 3.740 58.240 3.790 ;
        RECT 49.740 3.540 49.970 3.545 ;
        RECT 40.605 3.395 42.855 3.405 ;
        RECT 45.935 3.320 48.730 3.490 ;
        RECT 45.935 3.290 46.260 3.320 ;
        RECT 48.380 3.260 48.730 3.320 ;
        RECT 47.950 3.120 48.240 3.150 ;
        RECT 48.920 3.120 49.270 3.150 ;
        RECT 47.950 2.950 49.270 3.120 ;
        RECT 47.950 2.920 48.240 2.950 ;
        RECT 31.365 2.180 31.655 2.410 ;
        RECT 33.155 2.180 33.450 2.440 ;
        RECT 48.010 2.410 48.180 2.920 ;
        RECT 48.920 2.860 49.270 2.950 ;
        RECT 49.800 2.440 49.970 3.540 ;
        RECT 57.190 3.540 57.330 3.740 ;
        RECT 57.780 3.720 58.100 3.740 ;
        RECT 58.460 3.730 58.780 3.790 ;
        RECT 59.510 3.670 59.770 3.700 ;
        RECT 59.480 3.650 59.800 3.670 ;
        RECT 60.250 3.650 60.390 3.790 ;
        RECT 63.875 3.695 64.510 3.865 ;
        RECT 63.990 3.685 64.510 3.695 ;
        RECT 64.165 3.665 64.510 3.685 ;
        RECT 64.165 3.655 64.455 3.665 ;
        RECT 59.380 3.540 59.800 3.650 ;
        RECT 57.190 3.410 59.800 3.540 ;
        RECT 60.170 3.420 60.460 3.650 ;
        RECT 62.520 3.495 62.845 3.620 ;
        RECT 64.965 3.495 65.315 3.615 ;
        RECT 66.325 3.550 66.615 3.785 ;
        RECT 73.695 3.745 73.985 3.975 ;
        RECT 74.365 3.935 74.825 3.975 ;
        RECT 75.045 3.935 75.365 3.995 ;
        RECT 76.495 3.935 76.635 4.075 ;
        RECT 74.365 3.795 74.845 3.935 ;
        RECT 75.045 3.795 75.635 3.935 ;
        RECT 76.495 3.795 76.975 3.935 ;
        RECT 80.775 3.890 81.095 3.990 ;
        RECT 90.945 3.975 91.265 3.985 ;
        RECT 80.750 3.870 81.095 3.890 ;
        RECT 74.365 3.745 74.825 3.795 ;
        RECT 66.325 3.545 66.555 3.550 ;
        RECT 57.190 3.400 59.440 3.410 ;
        RECT 62.520 3.325 65.315 3.495 ;
        RECT 62.520 3.295 62.845 3.325 ;
        RECT 64.965 3.265 65.315 3.325 ;
        RECT 64.535 3.125 64.825 3.155 ;
        RECT 65.505 3.125 65.855 3.155 ;
        RECT 64.535 2.955 65.855 3.125 ;
        RECT 64.535 2.925 64.825 2.955 ;
        RECT 47.950 2.180 48.240 2.410 ;
        RECT 49.740 2.180 50.035 2.440 ;
        RECT 64.595 2.415 64.765 2.925 ;
        RECT 65.505 2.865 65.855 2.955 ;
        RECT 66.385 2.445 66.555 3.545 ;
        RECT 73.775 3.545 73.915 3.745 ;
        RECT 74.365 3.725 74.685 3.745 ;
        RECT 75.045 3.735 75.365 3.795 ;
        RECT 76.095 3.675 76.355 3.705 ;
        RECT 76.065 3.655 76.385 3.675 ;
        RECT 76.835 3.655 76.975 3.795 ;
        RECT 80.460 3.700 81.095 3.870 ;
        RECT 80.575 3.690 81.095 3.700 ;
        RECT 80.750 3.670 81.095 3.690 ;
        RECT 80.750 3.660 81.040 3.670 ;
        RECT 75.965 3.545 76.385 3.655 ;
        RECT 73.775 3.415 76.385 3.545 ;
        RECT 76.755 3.425 77.045 3.655 ;
        RECT 79.105 3.500 79.430 3.625 ;
        RECT 81.550 3.500 81.900 3.620 ;
        RECT 82.910 3.555 83.200 3.790 ;
        RECT 90.275 3.745 90.565 3.975 ;
        RECT 90.945 3.935 91.405 3.975 ;
        RECT 91.625 3.935 91.945 3.995 ;
        RECT 93.075 3.935 93.215 4.075 ;
        RECT 90.945 3.795 91.425 3.935 ;
        RECT 91.625 3.795 92.215 3.935 ;
        RECT 93.075 3.795 93.555 3.935 ;
        RECT 97.355 3.890 97.675 3.990 ;
        RECT 97.330 3.870 97.675 3.890 ;
        RECT 90.945 3.745 91.405 3.795 ;
        RECT 82.910 3.550 83.140 3.555 ;
        RECT 73.775 3.405 76.025 3.415 ;
        RECT 79.105 3.330 81.900 3.500 ;
        RECT 79.105 3.300 79.430 3.330 ;
        RECT 81.550 3.270 81.900 3.330 ;
        RECT 81.120 3.130 81.410 3.160 ;
        RECT 82.090 3.130 82.440 3.160 ;
        RECT 81.120 2.960 82.440 3.130 ;
        RECT 81.120 2.930 81.410 2.960 ;
        RECT 64.535 2.185 64.825 2.415 ;
        RECT 66.325 2.185 66.620 2.445 ;
        RECT 81.180 2.420 81.350 2.930 ;
        RECT 82.090 2.870 82.440 2.960 ;
        RECT 82.970 2.450 83.140 3.550 ;
        RECT 90.355 3.545 90.495 3.745 ;
        RECT 90.945 3.725 91.265 3.745 ;
        RECT 91.625 3.735 91.945 3.795 ;
        RECT 92.675 3.675 92.935 3.705 ;
        RECT 92.645 3.655 92.965 3.675 ;
        RECT 93.415 3.655 93.555 3.795 ;
        RECT 97.040 3.700 97.675 3.870 ;
        RECT 97.155 3.690 97.675 3.700 ;
        RECT 97.330 3.670 97.675 3.690 ;
        RECT 97.330 3.660 97.620 3.670 ;
        RECT 92.545 3.545 92.965 3.655 ;
        RECT 90.355 3.415 92.965 3.545 ;
        RECT 93.335 3.425 93.625 3.655 ;
        RECT 95.685 3.500 96.010 3.625 ;
        RECT 98.130 3.500 98.480 3.620 ;
        RECT 99.490 3.555 99.780 3.790 ;
        RECT 99.490 3.550 99.720 3.555 ;
        RECT 90.355 3.405 92.605 3.415 ;
        RECT 95.685 3.330 98.480 3.500 ;
        RECT 95.685 3.300 96.010 3.330 ;
        RECT 98.130 3.270 98.480 3.330 ;
        RECT 97.700 3.130 97.990 3.160 ;
        RECT 98.670 3.130 99.020 3.160 ;
        RECT 97.700 2.960 99.020 3.130 ;
        RECT 97.700 2.930 97.990 2.960 ;
        RECT 81.120 2.190 81.410 2.420 ;
        RECT 82.910 2.190 83.205 2.450 ;
        RECT 97.760 2.420 97.930 2.930 ;
        RECT 98.670 2.870 99.020 2.960 ;
        RECT 99.550 2.450 99.720 3.550 ;
        RECT 97.700 2.190 97.990 2.420 ;
        RECT 99.490 2.190 99.785 2.450 ;
      LAYER met2 ;
        RECT 16.575 10.065 100.715 10.235 ;
        RECT 16.575 8.880 16.745 10.065 ;
        RECT 100.545 9.910 100.715 10.065 ;
        RECT 20.685 9.705 30.865 9.875 ;
        RECT 16.920 9.515 17.200 9.620 ;
        RECT 16.920 9.345 18.110 9.515 ;
        RECT 16.920 9.280 17.200 9.345 ;
        RECT 17.940 9.140 18.110 9.345 ;
        RECT 20.100 9.305 20.470 9.675 ;
        RECT 20.685 9.225 20.855 9.705 ;
        RECT 20.630 9.140 20.910 9.225 ;
        RECT 17.940 8.970 20.910 9.140 ;
        RECT 20.630 8.885 20.910 8.970 ;
        RECT 30.705 9.200 30.865 9.705 ;
        RECT 37.270 9.705 47.450 9.875 ;
        RECT 36.685 9.305 37.055 9.675 ;
        RECT 31.820 9.200 32.145 9.265 ;
        RECT 30.705 9.030 32.145 9.200 ;
        RECT 16.535 8.540 16.815 8.880 ;
        RECT 24.950 7.415 25.230 7.440 ;
        RECT 24.950 7.095 25.240 7.415 ;
        RECT 24.950 7.065 25.230 7.095 ;
        RECT 26.000 7.065 26.280 7.440 ;
        RECT 27.360 7.325 27.620 7.415 ;
        RECT 26.740 7.185 27.620 7.325 ;
        RECT 25.320 6.045 25.600 6.420 ;
        RECT 24.640 3.655 24.920 4.035 ;
        RECT 25.380 4.015 25.520 6.045 ;
        RECT 26.060 5.285 26.200 7.065 ;
        RECT 26.740 5.400 26.880 7.185 ;
        RECT 27.360 7.095 27.620 7.185 ;
        RECT 28.380 6.075 28.640 6.395 ;
        RECT 26.060 5.145 26.540 5.285 ;
        RECT 25.980 4.345 26.260 4.720 ;
        RECT 25.320 3.695 25.580 4.015 ;
        RECT 26.400 3.695 26.540 5.145 ;
        RECT 26.680 5.025 26.960 5.400 ;
        RECT 26.680 4.005 26.960 4.380 ;
        RECT 28.440 4.355 28.580 6.075 ;
        RECT 28.380 4.035 28.640 4.355 ;
        RECT 30.705 3.860 30.865 9.030 ;
        RECT 31.820 8.940 32.145 9.030 ;
        RECT 34.210 9.145 34.535 9.270 ;
        RECT 37.270 9.225 37.440 9.705 ;
        RECT 34.210 9.140 35.260 9.145 ;
        RECT 37.215 9.140 37.495 9.225 ;
        RECT 34.210 8.975 37.495 9.140 ;
        RECT 34.210 8.945 34.535 8.975 ;
        RECT 35.260 8.970 37.495 8.975 ;
        RECT 31.020 8.565 31.340 8.890 ;
        RECT 37.215 8.885 37.495 8.970 ;
        RECT 47.290 9.200 47.450 9.705 ;
        RECT 53.855 9.710 64.035 9.880 ;
        RECT 53.270 9.280 53.640 9.680 ;
        RECT 48.405 9.200 48.730 9.265 ;
        RECT 47.290 9.030 48.730 9.200 ;
        RECT 31.050 8.330 31.220 8.565 ;
        RECT 31.050 8.155 31.225 8.330 ;
        RECT 31.050 7.980 32.025 8.155 ;
        RECT 31.020 3.860 31.340 3.980 ;
        RECT 24.685 3.070 24.855 3.655 ;
        RECT 26.340 3.355 26.600 3.695 ;
        RECT 30.705 3.690 31.340 3.860 ;
        RECT 31.020 3.660 31.340 3.690 ;
        RECT 29.350 3.290 29.675 3.615 ;
        RECT 31.850 3.610 32.025 7.980 ;
        RECT 41.535 7.415 41.815 7.440 ;
        RECT 41.535 7.095 41.825 7.415 ;
        RECT 41.535 7.065 41.815 7.095 ;
        RECT 42.585 7.065 42.865 7.440 ;
        RECT 43.945 7.325 44.205 7.415 ;
        RECT 43.325 7.185 44.205 7.325 ;
        RECT 41.905 6.045 42.185 6.420 ;
        RECT 41.225 3.655 41.505 4.035 ;
        RECT 41.965 4.015 42.105 6.045 ;
        RECT 42.645 5.285 42.785 7.065 ;
        RECT 43.325 5.400 43.465 7.185 ;
        RECT 43.945 7.095 44.205 7.185 ;
        RECT 44.965 6.075 45.225 6.395 ;
        RECT 42.645 5.145 43.125 5.285 ;
        RECT 42.565 4.345 42.845 4.720 ;
        RECT 41.905 3.695 42.165 4.015 ;
        RECT 42.985 3.695 43.125 5.145 ;
        RECT 43.265 5.025 43.545 5.400 ;
        RECT 43.265 4.005 43.545 4.380 ;
        RECT 45.025 4.355 45.165 6.075 ;
        RECT 44.965 4.035 45.225 4.355 ;
        RECT 47.290 3.860 47.450 9.030 ;
        RECT 48.405 8.940 48.730 9.030 ;
        RECT 50.795 9.145 51.120 9.270 ;
        RECT 53.855 9.230 54.025 9.710 ;
        RECT 50.795 9.140 52.075 9.145 ;
        RECT 53.800 9.140 54.080 9.230 ;
        RECT 50.795 8.975 54.080 9.140 ;
        RECT 50.795 8.945 51.120 8.975 ;
        RECT 52.075 8.970 54.080 8.975 ;
        RECT 53.800 8.890 54.080 8.970 ;
        RECT 63.875 9.205 64.035 9.710 ;
        RECT 70.440 9.715 80.620 9.885 ;
        RECT 69.855 9.280 70.225 9.685 ;
        RECT 64.990 9.205 65.315 9.270 ;
        RECT 63.875 9.035 65.315 9.205 ;
        RECT 47.605 8.565 47.925 8.890 ;
        RECT 47.635 8.330 47.805 8.565 ;
        RECT 47.635 8.155 47.810 8.330 ;
        RECT 47.635 7.980 48.610 8.155 ;
        RECT 47.605 3.860 47.925 3.980 ;
        RECT 29.425 3.070 29.595 3.290 ;
        RECT 31.795 3.260 32.145 3.610 ;
        RECT 24.685 2.900 29.595 3.070 ;
        RECT 41.270 3.070 41.440 3.655 ;
        RECT 42.925 3.355 43.185 3.695 ;
        RECT 47.290 3.690 47.925 3.860 ;
        RECT 47.605 3.660 47.925 3.690 ;
        RECT 45.935 3.290 46.260 3.615 ;
        RECT 48.435 3.610 48.610 7.980 ;
        RECT 58.120 7.420 58.400 7.445 ;
        RECT 58.120 7.100 58.410 7.420 ;
        RECT 58.120 7.070 58.400 7.100 ;
        RECT 59.170 7.070 59.450 7.445 ;
        RECT 60.530 7.330 60.790 7.420 ;
        RECT 59.910 7.190 60.790 7.330 ;
        RECT 58.490 6.050 58.770 6.425 ;
        RECT 57.810 3.660 58.090 4.040 ;
        RECT 58.550 4.020 58.690 6.050 ;
        RECT 59.230 5.290 59.370 7.070 ;
        RECT 59.910 5.405 60.050 7.190 ;
        RECT 60.530 7.100 60.790 7.190 ;
        RECT 61.550 6.080 61.810 6.400 ;
        RECT 59.230 5.150 59.710 5.290 ;
        RECT 59.150 4.350 59.430 4.725 ;
        RECT 58.490 3.700 58.750 4.020 ;
        RECT 59.570 3.700 59.710 5.150 ;
        RECT 59.850 5.030 60.130 5.405 ;
        RECT 59.850 4.010 60.130 4.385 ;
        RECT 61.610 4.360 61.750 6.080 ;
        RECT 61.550 4.040 61.810 4.360 ;
        RECT 63.875 3.865 64.035 9.035 ;
        RECT 64.990 8.945 65.315 9.035 ;
        RECT 67.380 9.150 67.705 9.275 ;
        RECT 70.440 9.235 70.610 9.715 ;
        RECT 67.380 9.140 68.305 9.150 ;
        RECT 70.385 9.140 70.665 9.235 ;
        RECT 67.380 8.980 70.665 9.140 ;
        RECT 67.380 8.950 67.705 8.980 ;
        RECT 68.305 8.970 70.665 8.980 ;
        RECT 70.385 8.895 70.665 8.970 ;
        RECT 80.460 9.210 80.620 9.715 ;
        RECT 87.020 9.715 97.200 9.885 ;
        RECT 86.435 9.660 86.805 9.685 ;
        RECT 86.435 9.315 86.810 9.660 ;
        RECT 86.440 9.280 86.810 9.315 ;
        RECT 81.575 9.210 81.900 9.275 ;
        RECT 80.460 9.040 81.900 9.210 ;
        RECT 64.190 8.570 64.510 8.895 ;
        RECT 64.220 8.335 64.390 8.570 ;
        RECT 64.220 8.160 64.395 8.335 ;
        RECT 64.220 7.985 65.195 8.160 ;
        RECT 64.190 3.865 64.510 3.985 ;
        RECT 46.010 3.070 46.180 3.290 ;
        RECT 48.380 3.260 48.730 3.610 ;
        RECT 41.270 2.900 46.180 3.070 ;
        RECT 57.855 3.075 58.025 3.660 ;
        RECT 59.510 3.360 59.770 3.700 ;
        RECT 63.875 3.695 64.510 3.865 ;
        RECT 64.190 3.665 64.510 3.695 ;
        RECT 62.520 3.295 62.845 3.620 ;
        RECT 65.020 3.615 65.195 7.985 ;
        RECT 74.705 7.425 74.985 7.450 ;
        RECT 74.705 7.105 74.995 7.425 ;
        RECT 74.705 7.075 74.985 7.105 ;
        RECT 75.755 7.075 76.035 7.450 ;
        RECT 77.115 7.335 77.375 7.425 ;
        RECT 76.495 7.195 77.375 7.335 ;
        RECT 75.075 6.055 75.355 6.430 ;
        RECT 74.395 3.665 74.675 4.045 ;
        RECT 75.135 4.025 75.275 6.055 ;
        RECT 75.815 5.295 75.955 7.075 ;
        RECT 76.495 5.410 76.635 7.195 ;
        RECT 77.115 7.105 77.375 7.195 ;
        RECT 78.135 6.085 78.395 6.405 ;
        RECT 75.815 5.155 76.295 5.295 ;
        RECT 75.735 4.355 76.015 4.730 ;
        RECT 75.075 3.705 75.335 4.025 ;
        RECT 76.155 3.705 76.295 5.155 ;
        RECT 76.435 5.035 76.715 5.410 ;
        RECT 76.435 4.015 76.715 4.390 ;
        RECT 78.195 4.365 78.335 6.085 ;
        RECT 78.135 4.045 78.395 4.365 ;
        RECT 80.460 3.870 80.620 9.040 ;
        RECT 81.575 8.950 81.900 9.040 ;
        RECT 83.965 9.155 84.290 9.280 ;
        RECT 87.020 9.235 87.190 9.715 ;
        RECT 83.965 9.140 84.840 9.155 ;
        RECT 86.965 9.140 87.245 9.235 ;
        RECT 83.965 8.985 87.245 9.140 ;
        RECT 83.965 8.955 84.290 8.985 ;
        RECT 84.840 8.970 87.245 8.985 ;
        RECT 80.775 8.575 81.095 8.900 ;
        RECT 86.965 8.895 87.245 8.970 ;
        RECT 97.040 9.210 97.200 9.715 ;
        RECT 100.510 9.585 100.835 9.910 ;
        RECT 98.155 9.210 98.480 9.275 ;
        RECT 97.040 9.040 98.480 9.210 ;
        RECT 80.805 8.340 80.975 8.575 ;
        RECT 80.805 8.165 80.980 8.340 ;
        RECT 80.805 7.990 81.780 8.165 ;
        RECT 80.775 3.870 81.095 3.990 ;
        RECT 62.595 3.075 62.765 3.295 ;
        RECT 64.965 3.265 65.315 3.615 ;
        RECT 57.855 2.905 62.765 3.075 ;
        RECT 74.440 3.080 74.610 3.665 ;
        RECT 76.095 3.365 76.355 3.705 ;
        RECT 80.460 3.700 81.095 3.870 ;
        RECT 80.775 3.670 81.095 3.700 ;
        RECT 79.105 3.300 79.430 3.625 ;
        RECT 81.605 3.620 81.780 7.990 ;
        RECT 91.285 7.425 91.565 7.450 ;
        RECT 91.285 7.105 91.575 7.425 ;
        RECT 91.285 7.075 91.565 7.105 ;
        RECT 92.335 7.075 92.615 7.450 ;
        RECT 93.695 7.335 93.955 7.425 ;
        RECT 93.075 7.195 93.955 7.335 ;
        RECT 91.655 6.055 91.935 6.430 ;
        RECT 90.975 3.665 91.255 4.045 ;
        RECT 91.715 4.025 91.855 6.055 ;
        RECT 92.395 5.295 92.535 7.075 ;
        RECT 93.075 5.410 93.215 7.195 ;
        RECT 93.695 7.105 93.955 7.195 ;
        RECT 94.715 6.085 94.975 6.405 ;
        RECT 92.395 5.155 92.875 5.295 ;
        RECT 92.315 4.355 92.595 4.730 ;
        RECT 91.655 3.705 91.915 4.025 ;
        RECT 92.735 3.705 92.875 5.155 ;
        RECT 93.015 5.035 93.295 5.410 ;
        RECT 93.015 4.015 93.295 4.390 ;
        RECT 94.775 4.365 94.915 6.085 ;
        RECT 94.715 4.045 94.975 4.365 ;
        RECT 97.040 3.870 97.200 9.040 ;
        RECT 98.155 8.950 98.480 9.040 ;
        RECT 97.355 8.575 97.675 8.900 ;
        RECT 97.385 8.340 97.555 8.575 ;
        RECT 97.385 8.165 97.560 8.340 ;
        RECT 97.385 7.990 98.360 8.165 ;
        RECT 97.355 3.870 97.675 3.990 ;
        RECT 79.180 3.080 79.350 3.300 ;
        RECT 81.550 3.270 81.900 3.620 ;
        RECT 74.440 2.910 79.350 3.080 ;
        RECT 91.020 3.080 91.190 3.665 ;
        RECT 92.675 3.365 92.935 3.705 ;
        RECT 97.040 3.700 97.675 3.870 ;
        RECT 97.355 3.670 97.675 3.700 ;
        RECT 95.685 3.300 96.010 3.625 ;
        RECT 98.185 3.620 98.360 7.990 ;
        RECT 95.760 3.080 95.930 3.300 ;
        RECT 98.130 3.270 98.480 3.620 ;
        RECT 91.020 2.910 95.930 3.080 ;
      LAYER met3 ;
        RECT 20.100 9.615 20.470 9.675 ;
        RECT 36.685 9.615 37.055 9.675 ;
        RECT 53.270 9.620 53.640 9.680 ;
        RECT 69.855 9.625 70.225 9.685 ;
        RECT 86.435 9.625 86.805 9.685 ;
        RECT 20.100 9.315 25.255 9.615 ;
        RECT 36.685 9.315 41.840 9.615 ;
        RECT 53.270 9.320 58.425 9.620 ;
        RECT 69.855 9.325 75.010 9.625 ;
        RECT 86.435 9.325 91.590 9.625 ;
        RECT 20.100 9.305 20.470 9.315 ;
        RECT 24.950 7.420 25.250 9.315 ;
        RECT 36.685 9.305 37.055 9.315 ;
        RECT 41.535 7.420 41.835 9.315 ;
        RECT 53.270 9.310 53.640 9.320 ;
        RECT 58.120 7.425 58.420 9.320 ;
        RECT 69.855 9.315 70.225 9.325 ;
        RECT 74.705 7.430 75.005 9.325 ;
        RECT 86.435 9.315 86.805 9.325 ;
        RECT 91.285 7.430 91.585 9.325 ;
        RECT 24.320 7.405 25.260 7.420 ;
        RECT 25.960 7.405 26.305 7.420 ;
        RECT 40.905 7.405 41.845 7.420 ;
        RECT 42.545 7.405 42.890 7.420 ;
        RECT 57.490 7.410 58.430 7.425 ;
        RECT 59.130 7.410 59.475 7.425 ;
        RECT 74.075 7.415 75.015 7.430 ;
        RECT 75.715 7.415 76.060 7.430 ;
        RECT 90.655 7.415 91.595 7.430 ;
        RECT 92.295 7.415 92.640 7.430 ;
        RECT 24.320 7.105 26.770 7.405 ;
        RECT 40.905 7.105 43.355 7.405 ;
        RECT 57.490 7.110 59.940 7.410 ;
        RECT 74.075 7.115 76.525 7.415 ;
        RECT 90.655 7.115 93.105 7.415 ;
        RECT 24.320 7.090 26.305 7.105 ;
        RECT 24.320 7.080 25.260 7.090 ;
        RECT 24.320 5.390 24.620 7.080 ;
        RECT 24.920 7.075 25.260 7.080 ;
        RECT 25.960 7.085 26.305 7.090 ;
        RECT 40.905 7.090 42.890 7.105 ;
        RECT 25.960 7.075 26.300 7.085 ;
        RECT 40.905 7.080 41.845 7.090 ;
        RECT 25.280 6.385 25.625 6.400 ;
        RECT 25.280 6.085 26.090 6.385 ;
        RECT 25.280 6.055 25.625 6.085 ;
        RECT 40.905 5.390 41.205 7.080 ;
        RECT 41.505 7.075 41.845 7.080 ;
        RECT 42.545 7.085 42.890 7.090 ;
        RECT 57.490 7.095 59.475 7.110 ;
        RECT 57.490 7.085 58.430 7.095 ;
        RECT 42.545 7.075 42.885 7.085 ;
        RECT 41.865 6.385 42.210 6.400 ;
        RECT 41.865 6.085 42.675 6.385 ;
        RECT 41.865 6.055 42.210 6.085 ;
        RECT 57.490 5.395 57.790 7.085 ;
        RECT 58.090 7.080 58.430 7.085 ;
        RECT 59.130 7.090 59.475 7.095 ;
        RECT 74.075 7.100 76.060 7.115 ;
        RECT 74.075 7.090 75.015 7.100 ;
        RECT 59.130 7.080 59.470 7.090 ;
        RECT 58.450 6.390 58.795 6.405 ;
        RECT 58.450 6.090 59.260 6.390 ;
        RECT 58.450 6.060 58.795 6.090 ;
        RECT 74.075 5.400 74.375 7.090 ;
        RECT 74.675 7.085 75.015 7.090 ;
        RECT 75.715 7.095 76.060 7.100 ;
        RECT 90.655 7.100 92.640 7.115 ;
        RECT 75.715 7.085 76.055 7.095 ;
        RECT 90.655 7.090 91.595 7.100 ;
        RECT 75.035 6.395 75.380 6.410 ;
        RECT 75.035 6.095 75.845 6.395 ;
        RECT 75.035 6.065 75.380 6.095 ;
        RECT 90.655 5.400 90.955 7.090 ;
        RECT 91.255 7.085 91.595 7.090 ;
        RECT 92.295 7.095 92.640 7.100 ;
        RECT 92.295 7.085 92.635 7.095 ;
        RECT 91.615 6.395 91.960 6.410 ;
        RECT 91.615 6.095 92.425 6.395 ;
        RECT 91.615 6.065 91.960 6.095 ;
        RECT 74.075 5.395 76.730 5.400 ;
        RECT 90.655 5.395 93.310 5.400 ;
        RECT 57.490 5.390 60.145 5.395 ;
        RECT 24.320 5.385 26.975 5.390 ;
        RECT 40.905 5.385 43.560 5.390 ;
        RECT 24.320 5.365 26.985 5.385 ;
        RECT 40.905 5.365 43.570 5.385 ;
        RECT 57.490 5.370 60.155 5.390 ;
        RECT 74.075 5.375 76.740 5.395 ;
        RECT 90.655 5.375 93.320 5.395 ;
        RECT 24.320 5.065 27.450 5.365 ;
        RECT 40.905 5.065 44.035 5.365 ;
        RECT 57.490 5.070 60.620 5.370 ;
        RECT 74.075 5.075 77.205 5.375 ;
        RECT 90.655 5.075 93.785 5.375 ;
        RECT 74.075 5.070 76.740 5.075 ;
        RECT 90.655 5.070 93.320 5.075 ;
        RECT 57.490 5.065 60.155 5.070 ;
        RECT 24.320 5.060 26.985 5.065 ;
        RECT 40.905 5.060 43.570 5.065 ;
        RECT 26.640 5.035 26.985 5.060 ;
        RECT 43.225 5.035 43.570 5.060 ;
        RECT 59.810 5.040 60.155 5.065 ;
        RECT 76.395 5.045 76.740 5.070 ;
        RECT 92.975 5.045 93.320 5.070 ;
        RECT 26.660 4.995 26.960 5.035 ;
        RECT 43.245 4.995 43.545 5.035 ;
        RECT 59.830 5.000 60.130 5.040 ;
        RECT 76.415 5.005 76.715 5.045 ;
        RECT 92.995 5.005 93.295 5.045 ;
        RECT 25.950 4.685 26.290 4.705 ;
        RECT 42.535 4.685 42.875 4.705 ;
        RECT 59.120 4.690 59.460 4.710 ;
        RECT 75.705 4.695 76.045 4.715 ;
        RECT 92.285 4.695 92.625 4.715 ;
        RECT 25.480 4.385 26.290 4.685 ;
        RECT 42.065 4.385 42.875 4.685 ;
        RECT 58.650 4.390 59.460 4.690 ;
        RECT 75.235 4.395 76.045 4.695 ;
        RECT 91.815 4.395 92.625 4.695 ;
        RECT 25.950 4.355 26.290 4.385 ;
        RECT 26.650 4.355 26.985 4.360 ;
        RECT 42.535 4.355 42.875 4.385 ;
        RECT 59.120 4.360 59.460 4.390 ;
        RECT 75.705 4.365 76.045 4.395 ;
        RECT 76.405 4.365 76.740 4.370 ;
        RECT 92.285 4.365 92.625 4.395 ;
        RECT 92.985 4.365 93.320 4.370 ;
        RECT 59.820 4.360 60.155 4.365 ;
        RECT 43.235 4.355 43.570 4.360 ;
        RECT 26.640 4.345 26.985 4.355 ;
        RECT 43.225 4.345 43.570 4.355 ;
        RECT 59.810 4.350 60.155 4.360 ;
        RECT 76.395 4.355 76.740 4.365 ;
        RECT 92.975 4.355 93.320 4.365 ;
        RECT 26.640 4.045 27.450 4.345 ;
        RECT 43.225 4.045 44.035 4.345 ;
        RECT 59.810 4.050 60.620 4.350 ;
        RECT 76.395 4.055 77.205 4.355 ;
        RECT 92.975 4.055 93.785 4.355 ;
        RECT 26.640 4.025 26.985 4.045 ;
        RECT 43.225 4.025 43.570 4.045 ;
        RECT 59.810 4.030 60.155 4.050 ;
        RECT 76.395 4.035 76.740 4.055 ;
        RECT 92.975 4.035 93.320 4.055 ;
        RECT 26.640 4.015 26.980 4.025 ;
        RECT 43.225 4.015 43.565 4.025 ;
        RECT 59.810 4.020 60.150 4.030 ;
        RECT 76.395 4.025 76.735 4.035 ;
        RECT 92.975 4.025 93.315 4.035 ;
        RECT 24.600 4.005 24.945 4.015 ;
        RECT 41.185 4.005 41.530 4.015 ;
        RECT 57.770 4.010 58.115 4.020 ;
        RECT 74.355 4.015 74.700 4.025 ;
        RECT 90.935 4.015 91.280 4.025 ;
        RECT 24.140 3.705 24.945 4.005 ;
        RECT 40.725 3.705 41.530 4.005 ;
        RECT 57.310 3.710 58.115 4.010 ;
        RECT 73.895 3.715 74.700 4.015 ;
        RECT 90.475 3.715 91.280 4.015 ;
        RECT 24.500 3.695 24.945 3.705 ;
        RECT 41.085 3.695 41.530 3.705 ;
        RECT 57.670 3.700 58.115 3.710 ;
        RECT 74.255 3.705 74.700 3.715 ;
        RECT 90.835 3.705 91.280 3.715 ;
        RECT 24.600 3.675 24.945 3.695 ;
        RECT 41.185 3.675 41.530 3.695 ;
        RECT 57.770 3.680 58.115 3.700 ;
        RECT 74.355 3.685 74.700 3.705 ;
        RECT 90.935 3.685 91.280 3.705 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r2
MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r1
  CLASS BLOCK ;
  FOREIGN sky130_osu_ring_oscillator_mpr2xa_8_b0r1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 104.045 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 42.455 4.010 42.630 5.155 ;
        RECT 42.455 3.575 42.625 4.010 ;
        RECT 42.460 1.865 42.630 2.375 ;
      LAYER met1 ;
        RECT 42.395 3.540 42.685 3.775 ;
        RECT 42.395 3.535 42.625 3.540 ;
        RECT 42.455 2.435 42.625 3.535 ;
        RECT 42.395 2.175 42.690 2.435 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 57.715 4.010 57.890 5.155 ;
        RECT 57.715 3.575 57.885 4.010 ;
        RECT 57.720 1.865 57.890 2.375 ;
      LAYER met1 ;
        RECT 57.655 3.540 57.945 3.775 ;
        RECT 57.655 3.535 57.885 3.540 ;
        RECT 57.715 2.435 57.885 3.535 ;
        RECT 57.655 2.175 57.950 2.435 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 72.975 4.010 73.150 5.155 ;
        RECT 72.975 3.575 73.145 4.010 ;
        RECT 72.980 1.865 73.150 2.375 ;
      LAYER met1 ;
        RECT 72.915 3.540 73.205 3.775 ;
        RECT 72.915 3.535 73.145 3.540 ;
        RECT 72.975 2.435 73.145 3.535 ;
        RECT 72.915 2.175 73.210 2.435 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 88.235 4.010 88.410 5.155 ;
        RECT 88.235 3.575 88.405 4.010 ;
        RECT 88.240 1.865 88.410 2.375 ;
      LAYER met1 ;
        RECT 88.175 3.540 88.465 3.775 ;
        RECT 88.175 3.535 88.405 3.540 ;
        RECT 88.235 2.435 88.405 3.535 ;
        RECT 88.175 2.175 88.470 2.435 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 103.495 4.010 103.670 5.155 ;
        RECT 103.495 3.575 103.665 4.010 ;
        RECT 103.500 1.865 103.670 2.375 ;
      LAYER met1 ;
        RECT 103.435 3.540 103.725 3.775 ;
        RECT 103.435 3.535 103.665 3.540 ;
        RECT 103.495 2.435 103.665 3.535 ;
        RECT 103.435 2.175 103.730 2.435 ;
    END
  END X5_Y1
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 25.175 8.240 25.345 9.510 ;
      LAYER met1 ;
        RECT 25.115 8.435 25.405 8.440 ;
        RECT 25.115 8.410 25.410 8.435 ;
        RECT 25.115 8.240 25.575 8.410 ;
        RECT 25.115 8.210 25.410 8.240 ;
        RECT 25.120 8.205 25.410 8.210 ;
    END
  END start
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 10.865 104.045 12.465 ;
        RECT 25.165 10.240 25.335 10.865 ;
        RECT 32.680 10.240 32.850 10.865 ;
        RECT 33.635 10.320 33.805 10.600 ;
        RECT 33.635 10.150 33.865 10.320 ;
        RECT 38.295 10.240 38.465 10.865 ;
        RECT 41.040 10.240 41.210 10.865 ;
        RECT 42.030 10.240 42.200 10.865 ;
        RECT 47.940 10.240 48.110 10.865 ;
        RECT 48.895 10.320 49.065 10.600 ;
        RECT 48.895 10.150 49.125 10.320 ;
        RECT 53.555 10.240 53.725 10.865 ;
        RECT 56.300 10.240 56.470 10.865 ;
        RECT 57.290 10.240 57.460 10.865 ;
        RECT 63.200 10.240 63.370 10.865 ;
        RECT 64.155 10.320 64.325 10.600 ;
        RECT 64.155 10.150 64.385 10.320 ;
        RECT 68.815 10.240 68.985 10.865 ;
        RECT 71.560 10.240 71.730 10.865 ;
        RECT 72.550 10.240 72.720 10.865 ;
        RECT 78.460 10.240 78.630 10.865 ;
        RECT 79.415 10.320 79.585 10.600 ;
        RECT 79.415 10.150 79.645 10.320 ;
        RECT 84.075 10.240 84.245 10.865 ;
        RECT 86.820 10.240 86.990 10.865 ;
        RECT 87.810 10.240 87.980 10.865 ;
        RECT 93.720 10.240 93.890 10.865 ;
        RECT 94.675 10.320 94.845 10.600 ;
        RECT 94.675 10.150 94.905 10.320 ;
        RECT 99.335 10.240 99.505 10.865 ;
        RECT 102.080 10.240 102.250 10.865 ;
        RECT 103.070 10.240 103.240 10.865 ;
        RECT 33.695 8.540 33.865 10.150 ;
        RECT 48.955 8.540 49.125 10.150 ;
        RECT 64.215 8.540 64.385 10.150 ;
        RECT 79.475 8.540 79.645 10.150 ;
        RECT 94.735 8.540 94.905 10.150 ;
        RECT 33.635 8.370 33.865 8.540 ;
        RECT 48.895 8.370 49.125 8.540 ;
        RECT 64.155 8.370 64.385 8.540 ;
        RECT 79.415 8.370 79.645 8.540 ;
        RECT 94.675 8.370 94.905 8.540 ;
        RECT 33.635 7.310 33.805 8.370 ;
        RECT 48.895 7.310 49.065 8.370 ;
        RECT 64.155 7.310 64.325 8.370 ;
        RECT 79.415 7.310 79.585 8.370 ;
        RECT 94.675 7.310 94.845 8.370 ;
      LAYER met1 ;
        RECT 0.000 10.865 104.045 12.465 ;
        RECT 33.465 8.820 33.635 10.865 ;
        RECT 48.725 8.820 48.895 10.865 ;
        RECT 63.985 8.820 64.155 10.865 ;
        RECT 79.245 8.820 79.415 10.865 ;
        RECT 94.505 8.820 94.675 10.865 ;
        RECT 33.465 8.790 33.925 8.820 ;
        RECT 48.725 8.790 49.185 8.820 ;
        RECT 63.985 8.790 64.445 8.820 ;
        RECT 79.245 8.790 79.705 8.820 ;
        RECT 94.505 8.790 94.965 8.820 ;
        RECT 33.460 8.620 33.925 8.790 ;
        RECT 48.720 8.620 49.185 8.790 ;
        RECT 63.980 8.620 64.445 8.790 ;
        RECT 79.240 8.620 79.705 8.790 ;
        RECT 94.500 8.620 94.965 8.790 ;
        RECT 33.465 8.605 33.925 8.620 ;
        RECT 48.725 8.605 49.185 8.620 ;
        RECT 63.985 8.605 64.445 8.620 ;
        RECT 79.245 8.605 79.705 8.620 ;
        RECT 94.505 8.605 94.965 8.620 ;
        RECT 33.635 8.590 33.925 8.605 ;
        RECT 48.895 8.590 49.185 8.605 ;
        RECT 64.155 8.590 64.445 8.605 ;
        RECT 79.415 8.590 79.705 8.605 ;
        RECT 94.675 8.590 94.965 8.605 ;
    END
    PORT
      LAYER li1 ;
        RECT 29.045 3.785 29.215 4.235 ;
        RECT 30.365 3.865 30.735 4.035 ;
        RECT 30.365 3.395 30.535 3.865 ;
        RECT 44.305 3.785 44.475 4.235 ;
        RECT 45.625 3.865 45.995 4.035 ;
        RECT 45.625 3.395 45.795 3.865 ;
        RECT 59.565 3.785 59.735 4.235 ;
        RECT 60.885 3.865 61.255 4.035 ;
        RECT 60.885 3.395 61.055 3.865 ;
        RECT 74.825 3.785 74.995 4.235 ;
        RECT 76.145 3.865 76.515 4.035 ;
        RECT 76.145 3.395 76.315 3.865 ;
        RECT 90.085 3.785 90.255 4.235 ;
        RECT 91.405 3.865 91.775 4.035 ;
        RECT 91.405 3.395 91.575 3.865 ;
        RECT 29.765 2.890 29.935 3.375 ;
        RECT 30.245 3.225 30.535 3.395 ;
        RECT 29.765 2.875 30.040 2.890 ;
        RECT 31.685 2.875 31.855 3.375 ;
        RECT 32.645 2.875 32.815 3.375 ;
        RECT 33.520 2.875 33.715 2.890 ;
        RECT 34.565 2.875 34.735 3.375 ;
        RECT 35.525 2.880 35.695 3.375 ;
        RECT 35.370 2.875 35.695 2.880 ;
        RECT 36.465 2.875 36.635 3.375 ;
        RECT 45.025 2.890 45.195 3.375 ;
        RECT 45.505 3.225 45.795 3.395 ;
        RECT 37.040 2.875 37.235 2.880 ;
        RECT 45.025 2.875 45.300 2.890 ;
        RECT 46.945 2.875 47.115 3.375 ;
        RECT 47.905 2.875 48.075 3.375 ;
        RECT 48.780 2.875 48.975 2.890 ;
        RECT 49.825 2.875 49.995 3.375 ;
        RECT 50.785 2.880 50.955 3.375 ;
        RECT 50.630 2.875 50.955 2.880 ;
        RECT 51.725 2.875 51.895 3.375 ;
        RECT 60.285 2.890 60.455 3.375 ;
        RECT 60.765 3.225 61.055 3.395 ;
        RECT 52.300 2.875 52.495 2.880 ;
        RECT 60.285 2.875 60.560 2.890 ;
        RECT 62.205 2.875 62.375 3.375 ;
        RECT 63.165 2.875 63.335 3.375 ;
        RECT 64.040 2.875 64.235 2.890 ;
        RECT 65.085 2.875 65.255 3.375 ;
        RECT 66.045 2.880 66.215 3.375 ;
        RECT 65.890 2.875 66.215 2.880 ;
        RECT 66.985 2.875 67.155 3.375 ;
        RECT 75.545 2.890 75.715 3.375 ;
        RECT 76.025 3.225 76.315 3.395 ;
        RECT 67.560 2.875 67.755 2.880 ;
        RECT 75.545 2.875 75.820 2.890 ;
        RECT 77.465 2.875 77.635 3.375 ;
        RECT 78.425 2.875 78.595 3.375 ;
        RECT 79.300 2.875 79.495 2.890 ;
        RECT 80.345 2.875 80.515 3.375 ;
        RECT 81.305 2.880 81.475 3.375 ;
        RECT 81.150 2.875 81.475 2.880 ;
        RECT 82.245 2.875 82.415 3.375 ;
        RECT 90.805 2.890 90.975 3.375 ;
        RECT 91.285 3.225 91.575 3.395 ;
        RECT 82.820 2.875 83.015 2.880 ;
        RECT 90.805 2.875 91.080 2.890 ;
        RECT 92.725 2.875 92.895 3.375 ;
        RECT 93.685 2.875 93.855 3.375 ;
        RECT 94.560 2.875 94.755 2.890 ;
        RECT 95.605 2.875 95.775 3.375 ;
        RECT 96.565 2.880 96.735 3.375 ;
        RECT 96.410 2.875 96.735 2.880 ;
        RECT 97.505 2.875 97.675 3.375 ;
        RECT 98.080 2.875 98.275 2.880 ;
        RECT 28.495 1.600 37.235 2.875 ;
        RECT 38.295 1.600 38.465 2.225 ;
        RECT 41.040 1.600 41.210 2.225 ;
        RECT 42.025 1.600 42.195 2.225 ;
        RECT 43.755 1.600 52.495 2.875 ;
        RECT 53.555 1.600 53.725 2.225 ;
        RECT 56.300 1.600 56.470 2.225 ;
        RECT 57.285 1.600 57.455 2.225 ;
        RECT 59.015 1.600 67.755 2.875 ;
        RECT 68.815 1.600 68.985 2.225 ;
        RECT 71.560 1.600 71.730 2.225 ;
        RECT 72.545 1.600 72.715 2.225 ;
        RECT 74.275 1.600 83.015 2.875 ;
        RECT 84.075 1.600 84.245 2.225 ;
        RECT 86.820 1.600 86.990 2.225 ;
        RECT 87.805 1.600 87.975 2.225 ;
        RECT 89.535 1.600 98.275 2.875 ;
        RECT 99.335 1.600 99.505 2.225 ;
        RECT 102.080 1.600 102.250 2.225 ;
        RECT 103.065 1.600 103.235 2.225 ;
        RECT 0.000 0.000 104.045 1.600 ;
      LAYER met1 ;
        RECT 28.985 4.035 29.275 4.265 ;
        RECT 44.245 4.035 44.535 4.265 ;
        RECT 59.505 4.035 59.795 4.265 ;
        RECT 74.765 4.035 75.055 4.265 ;
        RECT 90.025 4.035 90.315 4.265 ;
        RECT 29.055 3.805 29.195 4.035 ;
        RECT 44.315 3.805 44.455 4.035 ;
        RECT 59.575 3.805 59.715 4.035 ;
        RECT 74.835 3.805 74.975 4.035 ;
        RECT 90.095 3.805 90.235 4.035 ;
        RECT 29.055 3.665 29.675 3.805 ;
        RECT 44.315 3.665 44.935 3.805 ;
        RECT 59.575 3.665 60.195 3.805 ;
        RECT 74.835 3.665 75.455 3.805 ;
        RECT 90.095 3.665 90.715 3.805 ;
        RECT 29.535 3.505 29.675 3.665 ;
        RECT 44.795 3.505 44.935 3.665 ;
        RECT 60.055 3.505 60.195 3.665 ;
        RECT 75.315 3.505 75.455 3.665 ;
        RECT 90.575 3.505 90.715 3.665 ;
        RECT 29.295 3.445 29.675 3.505 ;
        RECT 44.555 3.445 44.935 3.505 ;
        RECT 59.815 3.445 60.195 3.505 ;
        RECT 75.075 3.445 75.455 3.505 ;
        RECT 90.335 3.445 90.715 3.505 ;
        RECT 29.295 3.385 29.885 3.445 ;
        RECT 30.185 3.385 30.475 3.425 ;
        RECT 29.295 3.245 30.475 3.385 ;
        RECT 44.555 3.385 45.145 3.445 ;
        RECT 45.445 3.385 45.735 3.425 ;
        RECT 44.555 3.245 45.735 3.385 ;
        RECT 59.815 3.385 60.405 3.445 ;
        RECT 60.705 3.385 60.995 3.425 ;
        RECT 59.815 3.245 60.995 3.385 ;
        RECT 75.075 3.385 75.665 3.445 ;
        RECT 75.965 3.385 76.255 3.425 ;
        RECT 75.075 3.245 76.255 3.385 ;
        RECT 90.335 3.385 90.925 3.445 ;
        RECT 91.225 3.385 91.515 3.425 ;
        RECT 90.335 3.245 91.515 3.385 ;
        RECT 29.480 3.185 29.885 3.245 ;
        RECT 30.185 3.195 30.475 3.245 ;
        RECT 44.740 3.185 45.145 3.245 ;
        RECT 45.445 3.195 45.735 3.245 ;
        RECT 60.000 3.185 60.405 3.245 ;
        RECT 60.705 3.195 60.995 3.245 ;
        RECT 75.260 3.185 75.665 3.245 ;
        RECT 75.965 3.195 76.255 3.245 ;
        RECT 90.520 3.185 90.925 3.245 ;
        RECT 91.225 3.195 91.515 3.245 ;
        RECT 29.480 2.915 29.770 3.185 ;
        RECT 37.040 2.915 37.235 2.920 ;
        RECT 44.740 2.915 45.030 3.185 ;
        RECT 52.300 2.915 52.495 2.920 ;
        RECT 60.000 2.915 60.290 3.185 ;
        RECT 67.560 2.915 67.755 2.920 ;
        RECT 75.260 2.915 75.550 3.185 ;
        RECT 82.820 2.915 83.015 2.920 ;
        RECT 90.520 2.915 90.810 3.185 ;
        RECT 98.080 2.915 98.275 2.920 ;
        RECT 28.495 1.600 37.235 2.915 ;
        RECT 43.755 1.600 52.495 2.915 ;
        RECT 59.015 1.600 67.755 2.915 ;
        RECT 74.275 1.600 83.015 2.915 ;
        RECT 89.535 1.600 98.275 2.915 ;
        RECT 0.000 0.000 104.045 1.600 ;
      LAYER met2 ;
        RECT 29.465 3.475 29.745 3.500 ;
        RECT 44.725 3.475 45.005 3.500 ;
        RECT 59.985 3.475 60.265 3.500 ;
        RECT 75.245 3.475 75.525 3.500 ;
        RECT 90.505 3.475 90.785 3.500 ;
        RECT 29.465 3.155 29.855 3.475 ;
        RECT 44.725 3.155 45.115 3.475 ;
        RECT 59.985 3.155 60.375 3.475 ;
        RECT 75.245 3.155 75.635 3.475 ;
        RECT 90.505 3.155 90.895 3.475 ;
        RECT 29.465 3.125 29.745 3.155 ;
        RECT 44.725 3.125 45.005 3.155 ;
        RECT 59.985 3.125 60.265 3.155 ;
        RECT 75.245 3.125 75.525 3.155 ;
        RECT 90.505 3.125 90.785 3.155 ;
      LAYER met3 ;
        RECT 29.425 3.475 29.780 3.480 ;
        RECT 44.685 3.475 45.040 3.480 ;
        RECT 59.945 3.475 60.300 3.480 ;
        RECT 75.205 3.475 75.560 3.480 ;
        RECT 90.465 3.475 90.820 3.480 ;
        RECT 29.325 3.145 30.055 3.475 ;
        RECT 44.585 3.145 45.315 3.475 ;
        RECT 59.845 3.145 60.575 3.475 ;
        RECT 75.105 3.145 75.835 3.475 ;
        RECT 90.365 3.145 91.095 3.475 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 24.945 8.745 27.755 8.750 ;
        RECT 32.460 8.745 35.270 8.750 ;
        RECT 38.075 8.745 42.855 8.750 ;
        RECT 47.720 8.745 50.530 8.750 ;
        RECT 53.335 8.745 58.115 8.750 ;
        RECT 62.980 8.745 65.790 8.750 ;
        RECT 68.595 8.745 73.375 8.750 ;
        RECT 78.240 8.745 81.050 8.750 ;
        RECT 83.855 8.745 88.635 8.750 ;
        RECT 93.500 8.745 96.310 8.750 ;
        RECT 99.115 8.745 103.895 8.750 ;
        RECT 24.945 6.660 104.045 8.745 ;
        RECT 24.980 4.100 104.045 6.660 ;
        RECT 27.745 4.095 104.045 4.100 ;
        RECT 37.055 3.720 43.005 4.095 ;
        RECT 52.315 3.720 58.265 4.095 ;
        RECT 67.575 3.720 73.525 4.095 ;
        RECT 82.835 3.720 88.785 4.095 ;
        RECT 98.095 3.720 104.045 4.095 ;
        RECT 38.075 3.715 42.850 3.720 ;
        RECT 53.335 3.715 58.110 3.720 ;
        RECT 68.595 3.715 73.370 3.720 ;
        RECT 83.855 3.715 88.630 3.720 ;
        RECT 99.115 3.715 103.890 3.720 ;
      LAYER li1 ;
        RECT 26.980 10.050 27.155 10.600 ;
        RECT 26.980 8.450 27.150 10.050 ;
        RECT 25.165 7.040 25.335 7.770 ;
        RECT 26.980 7.310 27.155 8.450 ;
        RECT 26.980 7.040 27.150 7.310 ;
        RECT 32.680 7.040 32.850 7.770 ;
        RECT 38.295 7.040 38.465 7.770 ;
        RECT 41.040 7.040 41.210 7.770 ;
        RECT 42.030 7.040 42.200 7.770 ;
        RECT 47.940 7.040 48.110 7.770 ;
        RECT 53.555 7.040 53.725 7.770 ;
        RECT 56.300 7.040 56.470 7.770 ;
        RECT 57.290 7.040 57.460 7.770 ;
        RECT 63.200 7.040 63.370 7.770 ;
        RECT 68.815 7.040 68.985 7.770 ;
        RECT 71.560 7.040 71.730 7.770 ;
        RECT 72.550 7.040 72.720 7.770 ;
        RECT 78.460 7.040 78.630 7.770 ;
        RECT 84.075 7.040 84.245 7.770 ;
        RECT 86.820 7.040 86.990 7.770 ;
        RECT 87.810 7.040 87.980 7.770 ;
        RECT 93.720 7.040 93.890 7.770 ;
        RECT 99.335 7.040 99.505 7.770 ;
        RECT 102.080 7.040 102.250 7.770 ;
        RECT 103.070 7.040 103.240 7.770 ;
        RECT 24.995 7.035 27.745 7.040 ;
        RECT 32.510 7.035 35.260 7.040 ;
        RECT 38.125 7.035 42.850 7.040 ;
        RECT 47.770 7.035 50.520 7.040 ;
        RECT 53.385 7.035 58.110 7.040 ;
        RECT 63.030 7.035 65.780 7.040 ;
        RECT 68.645 7.035 73.370 7.040 ;
        RECT 78.290 7.035 81.040 7.040 ;
        RECT 83.905 7.035 88.630 7.040 ;
        RECT 93.550 7.035 96.300 7.040 ;
        RECT 99.165 7.035 103.890 7.040 ;
        RECT 0.000 5.435 104.045 7.035 ;
        RECT 28.495 5.430 43.005 5.435 ;
        RECT 43.755 5.430 58.265 5.435 ;
        RECT 59.015 5.430 73.525 5.435 ;
        RECT 74.275 5.430 88.785 5.435 ;
        RECT 89.535 5.430 104.045 5.435 ;
        RECT 28.495 5.425 37.235 5.430 ;
        RECT 38.125 5.425 42.845 5.430 ;
        RECT 43.755 5.425 52.495 5.430 ;
        RECT 53.385 5.425 58.105 5.430 ;
        RECT 59.015 5.425 67.755 5.430 ;
        RECT 68.645 5.425 73.365 5.430 ;
        RECT 74.275 5.425 83.015 5.430 ;
        RECT 83.905 5.425 88.625 5.430 ;
        RECT 89.535 5.425 98.275 5.430 ;
        RECT 99.165 5.425 103.885 5.430 ;
        RECT 29.285 4.925 29.455 5.425 ;
        RECT 31.205 4.925 31.375 5.425 ;
        RECT 32.665 4.925 32.835 5.425 ;
        RECT 33.605 4.925 33.775 5.425 ;
        RECT 35.525 4.925 35.695 5.425 ;
        RECT 38.295 4.695 38.465 5.425 ;
        RECT 41.040 4.695 41.210 5.425 ;
        RECT 42.025 4.695 42.195 5.425 ;
        RECT 44.545 4.925 44.715 5.425 ;
        RECT 46.465 4.925 46.635 5.425 ;
        RECT 47.925 4.925 48.095 5.425 ;
        RECT 48.865 4.925 49.035 5.425 ;
        RECT 50.785 4.925 50.955 5.425 ;
        RECT 53.555 4.695 53.725 5.425 ;
        RECT 56.300 4.695 56.470 5.425 ;
        RECT 57.285 4.695 57.455 5.425 ;
        RECT 59.805 4.925 59.975 5.425 ;
        RECT 61.725 4.925 61.895 5.425 ;
        RECT 63.185 4.925 63.355 5.425 ;
        RECT 64.125 4.925 64.295 5.425 ;
        RECT 66.045 4.925 66.215 5.425 ;
        RECT 68.815 4.695 68.985 5.425 ;
        RECT 71.560 4.695 71.730 5.425 ;
        RECT 72.545 4.695 72.715 5.425 ;
        RECT 75.065 4.925 75.235 5.425 ;
        RECT 76.985 4.925 77.155 5.425 ;
        RECT 78.445 4.925 78.615 5.425 ;
        RECT 79.385 4.925 79.555 5.425 ;
        RECT 81.305 4.925 81.475 5.425 ;
        RECT 84.075 4.695 84.245 5.425 ;
        RECT 86.820 4.695 86.990 5.425 ;
        RECT 87.805 4.695 87.975 5.425 ;
        RECT 90.325 4.925 90.495 5.425 ;
        RECT 92.245 4.925 92.415 5.425 ;
        RECT 93.705 4.925 93.875 5.425 ;
        RECT 94.645 4.925 94.815 5.425 ;
        RECT 96.565 4.925 96.735 5.425 ;
        RECT 99.335 4.695 99.505 5.425 ;
        RECT 102.080 4.695 102.250 5.425 ;
        RECT 103.065 4.695 103.235 5.425 ;
      LAYER met1 ;
        RECT 26.920 9.150 27.210 9.180 ;
        RECT 26.750 8.980 27.210 9.150 ;
        RECT 26.920 8.950 27.210 8.980 ;
        RECT 24.995 7.035 27.745 7.040 ;
        RECT 32.510 7.035 35.260 7.040 ;
        RECT 38.125 7.035 42.850 7.040 ;
        RECT 47.770 7.035 50.520 7.040 ;
        RECT 53.385 7.035 58.110 7.040 ;
        RECT 63.030 7.035 65.780 7.040 ;
        RECT 68.645 7.035 73.370 7.040 ;
        RECT 78.290 7.035 81.040 7.040 ;
        RECT 83.905 7.035 88.630 7.040 ;
        RECT 93.550 7.035 96.300 7.040 ;
        RECT 99.165 7.035 103.890 7.040 ;
        RECT 0.000 5.435 104.045 7.035 ;
        RECT 28.495 5.430 43.005 5.435 ;
        RECT 43.755 5.430 58.265 5.435 ;
        RECT 59.015 5.430 73.525 5.435 ;
        RECT 74.275 5.430 88.785 5.435 ;
        RECT 89.535 5.430 104.045 5.435 ;
        RECT 28.495 5.395 37.235 5.430 ;
        RECT 38.125 5.425 42.845 5.430 ;
        RECT 43.755 5.395 52.495 5.430 ;
        RECT 53.385 5.425 58.105 5.430 ;
        RECT 59.015 5.395 67.755 5.430 ;
        RECT 68.645 5.425 73.365 5.430 ;
        RECT 74.275 5.395 83.015 5.430 ;
        RECT 83.905 5.425 88.625 5.430 ;
        RECT 89.535 5.395 98.275 5.430 ;
        RECT 99.165 5.425 103.885 5.430 ;
    END
  END vccd1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 32.690 8.240 32.860 9.510 ;
        RECT 38.305 8.240 38.475 9.510 ;
        RECT 38.305 2.955 38.475 4.225 ;
      LAYER met1 ;
        RECT 32.600 8.410 32.950 8.470 ;
        RECT 38.230 8.410 38.570 8.500 ;
        RECT 32.600 8.370 33.090 8.410 ;
        RECT 38.230 8.405 38.705 8.410 ;
        RECT 38.210 8.370 38.705 8.405 ;
        RECT 32.600 8.240 38.705 8.370 ;
        RECT 32.600 8.205 38.570 8.240 ;
        RECT 32.600 8.180 32.950 8.205 ;
        RECT 38.230 8.150 38.570 8.205 ;
        RECT 38.230 4.225 38.570 4.350 ;
        RECT 38.230 4.055 38.705 4.225 ;
        RECT 38.230 4.000 38.570 4.055 ;
      LAYER met2 ;
        RECT 38.230 8.150 38.570 8.500 ;
        RECT 38.310 4.350 38.480 8.150 ;
        RECT 38.230 4.000 38.570 4.350 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 47.950 8.240 48.120 9.510 ;
        RECT 53.565 8.240 53.735 9.510 ;
        RECT 53.565 2.955 53.735 4.225 ;
      LAYER met1 ;
        RECT 47.860 8.410 48.210 8.470 ;
        RECT 53.490 8.410 53.830 8.500 ;
        RECT 47.860 8.370 48.350 8.410 ;
        RECT 53.490 8.405 53.965 8.410 ;
        RECT 53.470 8.370 53.965 8.405 ;
        RECT 47.860 8.240 53.965 8.370 ;
        RECT 47.860 8.205 53.830 8.240 ;
        RECT 47.860 8.180 48.210 8.205 ;
        RECT 53.490 8.150 53.830 8.205 ;
        RECT 53.490 4.225 53.830 4.350 ;
        RECT 53.490 4.055 53.965 4.225 ;
        RECT 53.490 4.000 53.830 4.055 ;
      LAYER met2 ;
        RECT 53.490 8.150 53.830 8.500 ;
        RECT 53.570 4.350 53.740 8.150 ;
        RECT 53.490 4.000 53.830 4.350 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 63.210 8.240 63.380 9.510 ;
        RECT 68.825 8.240 68.995 9.510 ;
        RECT 68.825 2.955 68.995 4.225 ;
      LAYER met1 ;
        RECT 63.120 8.410 63.470 8.470 ;
        RECT 68.750 8.410 69.090 8.500 ;
        RECT 63.120 8.370 63.610 8.410 ;
        RECT 68.750 8.405 69.225 8.410 ;
        RECT 68.730 8.370 69.225 8.405 ;
        RECT 63.120 8.240 69.225 8.370 ;
        RECT 63.120 8.205 69.090 8.240 ;
        RECT 63.120 8.180 63.470 8.205 ;
        RECT 68.750 8.150 69.090 8.205 ;
        RECT 68.750 4.225 69.090 4.350 ;
        RECT 68.750 4.055 69.225 4.225 ;
        RECT 68.750 4.000 69.090 4.055 ;
      LAYER met2 ;
        RECT 68.750 8.150 69.090 8.500 ;
        RECT 68.830 4.350 69.000 8.150 ;
        RECT 68.750 4.000 69.090 4.350 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 78.470 8.240 78.640 9.510 ;
        RECT 84.085 8.240 84.255 9.510 ;
        RECT 84.085 2.955 84.255 4.225 ;
      LAYER met1 ;
        RECT 78.380 8.410 78.730 8.470 ;
        RECT 84.010 8.410 84.350 8.500 ;
        RECT 78.380 8.370 78.870 8.410 ;
        RECT 84.010 8.405 84.485 8.410 ;
        RECT 83.990 8.370 84.485 8.405 ;
        RECT 78.380 8.240 84.485 8.370 ;
        RECT 78.380 8.205 84.350 8.240 ;
        RECT 78.380 8.180 78.730 8.205 ;
        RECT 84.010 8.150 84.350 8.205 ;
        RECT 84.010 4.225 84.350 4.350 ;
        RECT 84.010 4.055 84.485 4.225 ;
        RECT 84.010 4.000 84.350 4.055 ;
      LAYER met2 ;
        RECT 84.010 8.150 84.350 8.500 ;
        RECT 84.090 4.350 84.260 8.150 ;
        RECT 84.010 4.000 84.350 4.350 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 93.730 8.240 93.900 9.510 ;
        RECT 99.345 8.240 99.515 9.510 ;
        RECT 99.345 2.955 99.515 4.225 ;
      LAYER met1 ;
        RECT 93.640 8.410 93.990 8.470 ;
        RECT 99.270 8.410 99.610 8.500 ;
        RECT 93.640 8.370 94.130 8.410 ;
        RECT 99.270 8.405 99.745 8.410 ;
        RECT 99.250 8.370 99.745 8.405 ;
        RECT 93.640 8.240 99.745 8.370 ;
        RECT 93.640 8.205 99.610 8.240 ;
        RECT 93.640 8.180 93.990 8.205 ;
        RECT 99.270 8.150 99.610 8.205 ;
        RECT 99.270 4.225 99.610 4.350 ;
        RECT 99.270 4.055 99.745 4.225 ;
        RECT 99.270 4.000 99.610 4.055 ;
      LAYER met2 ;
        RECT 99.270 8.150 99.610 8.500 ;
        RECT 99.350 4.350 99.520 8.150 ;
        RECT 99.270 4.000 99.610 4.350 ;
    END
  END s5
  OBS
      LAYER pwell ;
        RECT 28.875 2.715 29.045 2.875 ;
        RECT 44.135 2.715 44.305 2.875 ;
        RECT 59.395 2.715 59.565 2.875 ;
        RECT 74.655 2.715 74.825 2.875 ;
        RECT 89.915 2.715 90.085 2.875 ;
      LAYER li1 ;
        RECT 25.595 10.110 25.770 10.600 ;
        RECT 26.120 10.320 26.290 10.600 ;
        RECT 26.120 10.150 26.350 10.320 ;
        RECT 25.595 9.940 25.765 10.110 ;
        RECT 25.595 9.610 26.005 9.940 ;
        RECT 25.595 9.100 25.765 9.610 ;
        RECT 25.595 8.770 26.005 9.100 ;
        RECT 25.595 8.570 25.765 8.770 ;
        RECT 25.595 7.310 25.770 8.570 ;
        RECT 26.180 8.540 26.350 10.150 ;
        RECT 26.550 10.090 26.725 10.600 ;
        RECT 33.110 10.110 33.285 10.600 ;
        RECT 33.110 9.940 33.280 10.110 ;
        RECT 34.065 10.090 34.240 10.600 ;
        RECT 34.495 10.050 34.670 10.600 ;
        RECT 38.725 10.110 38.900 10.600 ;
        RECT 39.250 10.320 39.420 10.600 ;
        RECT 39.250 10.150 39.480 10.320 ;
        RECT 33.110 9.610 33.520 9.940 ;
        RECT 26.120 8.370 26.350 8.540 ;
        RECT 26.550 8.570 26.720 9.520 ;
        RECT 33.110 9.100 33.280 9.610 ;
        RECT 33.110 8.770 33.520 9.100 ;
        RECT 33.110 8.570 33.280 8.770 ;
        RECT 34.065 8.570 34.235 9.520 ;
        RECT 26.120 7.310 26.290 8.370 ;
        RECT 26.550 7.310 26.725 8.570 ;
        RECT 33.110 7.310 33.285 8.570 ;
        RECT 34.065 7.310 34.240 8.570 ;
        RECT 34.495 8.450 34.665 10.050 ;
        RECT 38.725 9.940 38.895 10.110 ;
        RECT 38.725 9.610 39.135 9.940 ;
        RECT 38.725 9.100 38.895 9.610 ;
        RECT 38.725 8.770 39.135 9.100 ;
        RECT 38.725 8.570 38.895 8.770 ;
        RECT 34.495 7.310 34.670 8.450 ;
        RECT 38.725 7.310 38.900 8.570 ;
        RECT 39.310 8.540 39.480 10.150 ;
        RECT 39.680 10.090 39.855 10.600 ;
        RECT 40.110 10.050 40.285 10.600 ;
        RECT 41.475 10.090 41.645 10.600 ;
        RECT 42.465 10.090 42.635 10.600 ;
        RECT 48.370 10.110 48.545 10.600 ;
        RECT 39.250 8.370 39.480 8.540 ;
        RECT 39.680 8.570 39.850 9.520 ;
        RECT 39.250 7.310 39.420 8.370 ;
        RECT 39.680 7.310 39.855 8.570 ;
        RECT 40.110 8.450 40.280 10.050 ;
        RECT 48.370 9.940 48.540 10.110 ;
        RECT 49.325 10.090 49.500 10.600 ;
        RECT 49.755 10.050 49.930 10.600 ;
        RECT 53.985 10.110 54.160 10.600 ;
        RECT 54.510 10.320 54.680 10.600 ;
        RECT 54.510 10.150 54.740 10.320 ;
        RECT 48.370 9.610 48.780 9.940 ;
        RECT 40.650 9.430 40.880 9.580 ;
        RECT 40.650 9.260 41.570 9.430 ;
        RECT 42.090 9.260 42.560 9.430 ;
        RECT 41.100 8.570 41.270 9.260 ;
        RECT 41.470 8.780 41.640 8.890 ;
        RECT 42.090 8.780 42.260 9.260 ;
        RECT 48.370 9.100 48.540 9.610 ;
        RECT 41.470 8.610 42.260 8.780 ;
        RECT 40.110 7.310 40.285 8.450 ;
        RECT 41.470 7.310 41.645 8.610 ;
        RECT 42.090 8.570 42.260 8.610 ;
        RECT 42.460 8.455 42.630 8.890 ;
        RECT 48.370 8.770 48.780 9.100 ;
        RECT 48.370 8.570 48.540 8.770 ;
        RECT 49.325 8.570 49.495 9.520 ;
        RECT 42.460 7.310 42.635 8.455 ;
        RECT 48.370 7.310 48.545 8.570 ;
        RECT 49.325 7.310 49.500 8.570 ;
        RECT 49.755 8.450 49.925 10.050 ;
        RECT 53.985 9.940 54.155 10.110 ;
        RECT 53.985 9.610 54.395 9.940 ;
        RECT 53.985 9.100 54.155 9.610 ;
        RECT 53.985 8.770 54.395 9.100 ;
        RECT 53.985 8.570 54.155 8.770 ;
        RECT 49.755 7.310 49.930 8.450 ;
        RECT 53.985 7.310 54.160 8.570 ;
        RECT 54.570 8.540 54.740 10.150 ;
        RECT 54.940 10.090 55.115 10.600 ;
        RECT 55.370 10.050 55.545 10.600 ;
        RECT 56.735 10.090 56.905 10.600 ;
        RECT 57.725 10.090 57.895 10.600 ;
        RECT 63.630 10.110 63.805 10.600 ;
        RECT 54.510 8.370 54.740 8.540 ;
        RECT 54.940 8.570 55.110 9.520 ;
        RECT 54.510 7.310 54.680 8.370 ;
        RECT 54.940 7.310 55.115 8.570 ;
        RECT 55.370 8.450 55.540 10.050 ;
        RECT 63.630 9.940 63.800 10.110 ;
        RECT 64.585 10.090 64.760 10.600 ;
        RECT 65.015 10.050 65.190 10.600 ;
        RECT 69.245 10.110 69.420 10.600 ;
        RECT 69.770 10.320 69.940 10.600 ;
        RECT 69.770 10.150 70.000 10.320 ;
        RECT 63.630 9.610 64.040 9.940 ;
        RECT 55.910 9.430 56.140 9.580 ;
        RECT 55.910 9.260 56.830 9.430 ;
        RECT 57.350 9.260 57.820 9.430 ;
        RECT 56.360 8.570 56.530 9.260 ;
        RECT 56.730 8.780 56.900 8.890 ;
        RECT 57.350 8.780 57.520 9.260 ;
        RECT 63.630 9.100 63.800 9.610 ;
        RECT 56.730 8.610 57.520 8.780 ;
        RECT 55.370 7.310 55.545 8.450 ;
        RECT 56.730 7.310 56.905 8.610 ;
        RECT 57.350 8.570 57.520 8.610 ;
        RECT 57.720 8.455 57.890 8.890 ;
        RECT 63.630 8.770 64.040 9.100 ;
        RECT 63.630 8.570 63.800 8.770 ;
        RECT 64.585 8.570 64.755 9.520 ;
        RECT 57.720 7.310 57.895 8.455 ;
        RECT 63.630 7.310 63.805 8.570 ;
        RECT 64.585 7.310 64.760 8.570 ;
        RECT 65.015 8.450 65.185 10.050 ;
        RECT 69.245 9.940 69.415 10.110 ;
        RECT 69.245 9.610 69.655 9.940 ;
        RECT 69.245 9.100 69.415 9.610 ;
        RECT 69.245 8.770 69.655 9.100 ;
        RECT 69.245 8.570 69.415 8.770 ;
        RECT 65.015 7.310 65.190 8.450 ;
        RECT 69.245 7.310 69.420 8.570 ;
        RECT 69.830 8.540 70.000 10.150 ;
        RECT 70.200 10.090 70.375 10.600 ;
        RECT 70.630 10.050 70.805 10.600 ;
        RECT 71.995 10.090 72.165 10.600 ;
        RECT 72.985 10.090 73.155 10.600 ;
        RECT 78.890 10.110 79.065 10.600 ;
        RECT 69.770 8.370 70.000 8.540 ;
        RECT 70.200 8.570 70.370 9.520 ;
        RECT 69.770 7.310 69.940 8.370 ;
        RECT 70.200 7.310 70.375 8.570 ;
        RECT 70.630 8.450 70.800 10.050 ;
        RECT 78.890 9.940 79.060 10.110 ;
        RECT 79.845 10.090 80.020 10.600 ;
        RECT 80.275 10.050 80.450 10.600 ;
        RECT 84.505 10.110 84.680 10.600 ;
        RECT 85.030 10.320 85.200 10.600 ;
        RECT 85.030 10.150 85.260 10.320 ;
        RECT 78.890 9.610 79.300 9.940 ;
        RECT 71.170 9.430 71.400 9.580 ;
        RECT 71.170 9.260 72.090 9.430 ;
        RECT 72.610 9.260 73.080 9.430 ;
        RECT 71.620 8.570 71.790 9.260 ;
        RECT 71.990 8.780 72.160 8.890 ;
        RECT 72.610 8.780 72.780 9.260 ;
        RECT 78.890 9.100 79.060 9.610 ;
        RECT 71.990 8.610 72.780 8.780 ;
        RECT 70.630 7.310 70.805 8.450 ;
        RECT 71.990 7.310 72.165 8.610 ;
        RECT 72.610 8.570 72.780 8.610 ;
        RECT 72.980 8.455 73.150 8.890 ;
        RECT 78.890 8.770 79.300 9.100 ;
        RECT 78.890 8.570 79.060 8.770 ;
        RECT 79.845 8.570 80.015 9.520 ;
        RECT 72.980 7.310 73.155 8.455 ;
        RECT 78.890 7.310 79.065 8.570 ;
        RECT 79.845 7.310 80.020 8.570 ;
        RECT 80.275 8.450 80.445 10.050 ;
        RECT 84.505 9.940 84.675 10.110 ;
        RECT 84.505 9.610 84.915 9.940 ;
        RECT 84.505 9.100 84.675 9.610 ;
        RECT 84.505 8.770 84.915 9.100 ;
        RECT 84.505 8.570 84.675 8.770 ;
        RECT 80.275 7.310 80.450 8.450 ;
        RECT 84.505 7.310 84.680 8.570 ;
        RECT 85.090 8.540 85.260 10.150 ;
        RECT 85.460 10.090 85.635 10.600 ;
        RECT 85.890 10.050 86.065 10.600 ;
        RECT 87.255 10.090 87.425 10.600 ;
        RECT 88.245 10.090 88.415 10.600 ;
        RECT 94.150 10.110 94.325 10.600 ;
        RECT 85.030 8.370 85.260 8.540 ;
        RECT 85.460 8.570 85.630 9.520 ;
        RECT 85.030 7.310 85.200 8.370 ;
        RECT 85.460 7.310 85.635 8.570 ;
        RECT 85.890 8.450 86.060 10.050 ;
        RECT 94.150 9.940 94.320 10.110 ;
        RECT 95.105 10.090 95.280 10.600 ;
        RECT 95.535 10.050 95.710 10.600 ;
        RECT 99.765 10.110 99.940 10.600 ;
        RECT 100.290 10.320 100.460 10.600 ;
        RECT 100.290 10.150 100.520 10.320 ;
        RECT 94.150 9.610 94.560 9.940 ;
        RECT 86.430 9.430 86.660 9.580 ;
        RECT 86.430 9.260 87.350 9.430 ;
        RECT 87.870 9.260 88.340 9.430 ;
        RECT 86.880 8.570 87.050 9.260 ;
        RECT 87.250 8.780 87.420 8.890 ;
        RECT 87.870 8.780 88.040 9.260 ;
        RECT 94.150 9.100 94.320 9.610 ;
        RECT 87.250 8.610 88.040 8.780 ;
        RECT 85.890 7.310 86.065 8.450 ;
        RECT 87.250 7.310 87.425 8.610 ;
        RECT 87.870 8.570 88.040 8.610 ;
        RECT 88.240 8.455 88.410 8.890 ;
        RECT 94.150 8.770 94.560 9.100 ;
        RECT 94.150 8.570 94.320 8.770 ;
        RECT 95.105 8.570 95.275 9.520 ;
        RECT 88.240 7.310 88.415 8.455 ;
        RECT 94.150 7.310 94.325 8.570 ;
        RECT 95.105 7.310 95.280 8.570 ;
        RECT 95.535 8.450 95.705 10.050 ;
        RECT 99.765 9.940 99.935 10.110 ;
        RECT 99.765 9.610 100.175 9.940 ;
        RECT 99.765 9.100 99.935 9.610 ;
        RECT 99.765 8.770 100.175 9.100 ;
        RECT 99.765 8.570 99.935 8.770 ;
        RECT 95.535 7.310 95.710 8.450 ;
        RECT 99.765 7.310 99.940 8.570 ;
        RECT 100.350 8.540 100.520 10.150 ;
        RECT 100.720 10.090 100.895 10.600 ;
        RECT 101.150 10.050 101.325 10.600 ;
        RECT 102.515 10.090 102.685 10.600 ;
        RECT 103.505 10.090 103.675 10.600 ;
        RECT 100.290 8.370 100.520 8.540 ;
        RECT 100.720 8.570 100.890 9.520 ;
        RECT 100.290 7.310 100.460 8.370 ;
        RECT 100.720 7.310 100.895 8.570 ;
        RECT 101.150 8.450 101.320 10.050 ;
        RECT 101.690 9.430 101.920 9.580 ;
        RECT 101.690 9.260 102.610 9.430 ;
        RECT 103.130 9.260 103.600 9.430 ;
        RECT 102.140 8.570 102.310 9.260 ;
        RECT 102.510 8.780 102.680 8.890 ;
        RECT 103.130 8.780 103.300 9.260 ;
        RECT 102.510 8.610 103.300 8.780 ;
        RECT 101.150 7.310 101.325 8.450 ;
        RECT 102.510 7.310 102.685 8.610 ;
        RECT 103.130 8.570 103.300 8.610 ;
        RECT 103.500 8.455 103.670 8.890 ;
        RECT 103.500 7.310 103.675 8.455 ;
        RECT 28.825 4.435 28.995 4.795 ;
        RECT 29.765 4.435 29.935 4.795 ;
        RECT 30.245 4.345 30.415 4.765 ;
        RECT 30.605 4.515 30.895 5.075 ;
        RECT 31.685 4.775 31.855 5.105 ;
        RECT 32.165 4.685 32.335 5.075 ;
        RECT 34.060 4.775 34.235 5.105 ;
        RECT 36.005 4.905 36.515 5.075 ;
        RECT 34.585 4.685 34.765 4.795 ;
        RECT 36.345 4.765 36.515 4.905 ;
        RECT 32.055 4.515 32.390 4.685 ;
        RECT 32.885 4.515 33.375 4.685 ;
        RECT 34.585 4.515 35.935 4.685 ;
        RECT 36.345 4.515 36.630 4.765 ;
        RECT 30.725 4.435 30.895 4.515 ;
        RECT 29.525 3.785 29.695 4.235 ;
        RECT 30.005 3.785 30.175 4.115 ;
        RECT 30.965 3.785 31.135 4.115 ;
        RECT 31.445 3.785 31.615 4.515 ;
        RECT 32.885 4.345 33.055 4.515 ;
        RECT 34.585 4.435 34.765 4.515 ;
        RECT 35.765 4.345 35.935 4.515 ;
        RECT 36.455 4.435 36.630 4.515 ;
        RECT 31.925 3.785 32.095 4.235 ;
        RECT 32.405 3.785 32.575 4.115 ;
        RECT 32.885 3.785 33.055 4.115 ;
        RECT 33.365 3.785 33.535 4.235 ;
        RECT 34.325 4.135 34.495 4.235 ;
        RECT 33.845 4.035 34.495 4.135 ;
        RECT 33.765 3.865 34.575 4.035 ;
        RECT 34.805 3.785 34.975 4.115 ;
        RECT 35.285 3.785 35.455 4.235 ;
        RECT 35.765 3.785 35.935 4.115 ;
        RECT 36.245 4.035 36.515 4.235 ;
        RECT 36.125 3.825 36.515 4.035 ;
        RECT 38.725 3.895 38.900 5.155 ;
        RECT 39.250 4.095 39.420 5.155 ;
        RECT 39.250 3.925 39.480 4.095 ;
        RECT 38.725 3.695 38.895 3.895 ;
        RECT 33.845 3.615 34.015 3.655 ;
        RECT 33.485 3.445 34.015 3.615 ;
        RECT 28.825 3.045 28.995 3.395 ;
        RECT 30.725 3.045 30.895 3.395 ;
        RECT 32.125 3.375 32.295 3.395 ;
        RECT 32.125 3.345 32.335 3.375 ;
        RECT 32.025 3.125 32.335 3.345 ;
        RECT 32.165 3.045 32.335 3.125 ;
        RECT 33.125 3.275 33.295 3.395 ;
        RECT 33.125 3.105 34.365 3.275 ;
        RECT 35.045 3.045 35.215 3.395 ;
        RECT 36.005 3.045 36.175 3.395 ;
        RECT 38.725 3.365 39.135 3.695 ;
        RECT 38.725 2.855 38.895 3.365 ;
        RECT 38.725 2.525 39.135 2.855 ;
        RECT 38.725 2.355 38.895 2.525 ;
        RECT 38.725 1.865 38.900 2.355 ;
        RECT 39.310 2.315 39.480 3.925 ;
        RECT 39.680 3.895 39.855 5.155 ;
        RECT 40.110 4.015 40.285 5.155 ;
        RECT 39.680 2.945 39.850 3.895 ;
        RECT 40.110 2.415 40.280 4.015 ;
        RECT 41.470 4.010 41.645 5.155 ;
        RECT 44.085 4.435 44.255 4.795 ;
        RECT 45.025 4.435 45.195 4.795 ;
        RECT 45.505 4.345 45.675 4.765 ;
        RECT 45.865 4.515 46.155 5.075 ;
        RECT 46.945 4.775 47.115 5.105 ;
        RECT 47.425 4.685 47.595 5.075 ;
        RECT 49.320 4.775 49.495 5.105 ;
        RECT 51.265 4.905 51.775 5.075 ;
        RECT 49.845 4.685 50.025 4.795 ;
        RECT 51.605 4.765 51.775 4.905 ;
        RECT 47.315 4.515 47.650 4.685 ;
        RECT 48.145 4.515 48.635 4.685 ;
        RECT 49.845 4.515 51.195 4.685 ;
        RECT 51.605 4.515 51.890 4.765 ;
        RECT 45.985 4.435 46.155 4.515 ;
        RECT 41.100 3.205 41.270 3.895 ;
        RECT 41.470 3.795 41.640 4.010 ;
        RECT 42.085 3.795 42.255 3.895 ;
        RECT 41.470 3.625 42.255 3.795 ;
        RECT 44.785 3.785 44.955 4.235 ;
        RECT 45.265 3.785 45.435 4.115 ;
        RECT 46.225 3.785 46.395 4.115 ;
        RECT 46.705 3.785 46.875 4.515 ;
        RECT 48.145 4.345 48.315 4.515 ;
        RECT 49.845 4.435 50.025 4.515 ;
        RECT 51.025 4.345 51.195 4.515 ;
        RECT 51.715 4.435 51.890 4.515 ;
        RECT 47.185 3.785 47.355 4.235 ;
        RECT 47.665 3.785 47.835 4.115 ;
        RECT 48.145 3.785 48.315 4.115 ;
        RECT 48.625 3.785 48.795 4.235 ;
        RECT 49.585 4.135 49.755 4.235 ;
        RECT 49.105 4.035 49.755 4.135 ;
        RECT 49.025 3.865 49.835 4.035 ;
        RECT 50.065 3.785 50.235 4.115 ;
        RECT 50.545 3.785 50.715 4.235 ;
        RECT 51.025 3.785 51.195 4.115 ;
        RECT 51.505 4.035 51.775 4.235 ;
        RECT 51.385 3.825 51.775 4.035 ;
        RECT 53.985 3.895 54.160 5.155 ;
        RECT 54.510 4.095 54.680 5.155 ;
        RECT 54.510 3.925 54.740 4.095 ;
        RECT 53.985 3.695 54.155 3.895 ;
        RECT 41.470 3.575 41.640 3.625 ;
        RECT 42.085 3.205 42.255 3.625 ;
        RECT 49.105 3.615 49.275 3.655 ;
        RECT 48.745 3.445 49.275 3.615 ;
        RECT 40.650 3.035 41.570 3.205 ;
        RECT 42.085 3.035 42.555 3.205 ;
        RECT 44.085 3.045 44.255 3.395 ;
        RECT 45.985 3.045 46.155 3.395 ;
        RECT 47.385 3.375 47.555 3.395 ;
        RECT 47.385 3.345 47.595 3.375 ;
        RECT 47.285 3.125 47.595 3.345 ;
        RECT 47.425 3.045 47.595 3.125 ;
        RECT 48.385 3.275 48.555 3.395 ;
        RECT 48.385 3.105 49.625 3.275 ;
        RECT 50.305 3.045 50.475 3.395 ;
        RECT 51.265 3.045 51.435 3.395 ;
        RECT 53.985 3.365 54.395 3.695 ;
        RECT 40.650 2.885 40.880 3.035 ;
        RECT 53.985 2.855 54.155 3.365 ;
        RECT 53.985 2.525 54.395 2.855 ;
        RECT 39.250 2.145 39.480 2.315 ;
        RECT 39.250 1.865 39.420 2.145 ;
        RECT 39.680 1.865 39.855 2.375 ;
        RECT 40.110 1.865 40.285 2.415 ;
        RECT 41.475 1.865 41.645 2.375 ;
        RECT 53.985 2.355 54.155 2.525 ;
        RECT 53.985 1.865 54.160 2.355 ;
        RECT 54.570 2.315 54.740 3.925 ;
        RECT 54.940 3.895 55.115 5.155 ;
        RECT 55.370 4.015 55.545 5.155 ;
        RECT 54.940 2.945 55.110 3.895 ;
        RECT 55.370 2.415 55.540 4.015 ;
        RECT 56.730 4.010 56.905 5.155 ;
        RECT 59.345 4.435 59.515 4.795 ;
        RECT 60.285 4.435 60.455 4.795 ;
        RECT 60.765 4.345 60.935 4.765 ;
        RECT 61.125 4.515 61.415 5.075 ;
        RECT 62.205 4.775 62.375 5.105 ;
        RECT 62.685 4.685 62.855 5.075 ;
        RECT 64.580 4.775 64.755 5.105 ;
        RECT 66.525 4.905 67.035 5.075 ;
        RECT 65.105 4.685 65.285 4.795 ;
        RECT 66.865 4.765 67.035 4.905 ;
        RECT 62.575 4.515 62.910 4.685 ;
        RECT 63.405 4.515 63.895 4.685 ;
        RECT 65.105 4.515 66.455 4.685 ;
        RECT 66.865 4.515 67.150 4.765 ;
        RECT 61.245 4.435 61.415 4.515 ;
        RECT 56.360 3.205 56.530 3.895 ;
        RECT 56.730 3.795 56.900 4.010 ;
        RECT 57.345 3.795 57.515 3.895 ;
        RECT 56.730 3.625 57.515 3.795 ;
        RECT 60.045 3.785 60.215 4.235 ;
        RECT 60.525 3.785 60.695 4.115 ;
        RECT 61.485 3.785 61.655 4.115 ;
        RECT 61.965 3.785 62.135 4.515 ;
        RECT 63.405 4.345 63.575 4.515 ;
        RECT 65.105 4.435 65.285 4.515 ;
        RECT 66.285 4.345 66.455 4.515 ;
        RECT 66.975 4.435 67.150 4.515 ;
        RECT 62.445 3.785 62.615 4.235 ;
        RECT 62.925 3.785 63.095 4.115 ;
        RECT 63.405 3.785 63.575 4.115 ;
        RECT 63.885 3.785 64.055 4.235 ;
        RECT 64.845 4.135 65.015 4.235 ;
        RECT 64.365 4.035 65.015 4.135 ;
        RECT 64.285 3.865 65.095 4.035 ;
        RECT 65.325 3.785 65.495 4.115 ;
        RECT 65.805 3.785 65.975 4.235 ;
        RECT 66.285 3.785 66.455 4.115 ;
        RECT 66.765 4.035 67.035 4.235 ;
        RECT 66.645 3.825 67.035 4.035 ;
        RECT 69.245 3.895 69.420 5.155 ;
        RECT 69.770 4.095 69.940 5.155 ;
        RECT 69.770 3.925 70.000 4.095 ;
        RECT 69.245 3.695 69.415 3.895 ;
        RECT 56.730 3.575 56.900 3.625 ;
        RECT 57.345 3.205 57.515 3.625 ;
        RECT 64.365 3.615 64.535 3.655 ;
        RECT 64.005 3.445 64.535 3.615 ;
        RECT 55.910 3.035 56.830 3.205 ;
        RECT 57.345 3.035 57.815 3.205 ;
        RECT 59.345 3.045 59.515 3.395 ;
        RECT 61.245 3.045 61.415 3.395 ;
        RECT 62.645 3.375 62.815 3.395 ;
        RECT 62.645 3.345 62.855 3.375 ;
        RECT 62.545 3.125 62.855 3.345 ;
        RECT 62.685 3.045 62.855 3.125 ;
        RECT 63.645 3.275 63.815 3.395 ;
        RECT 63.645 3.105 64.885 3.275 ;
        RECT 65.565 3.045 65.735 3.395 ;
        RECT 66.525 3.045 66.695 3.395 ;
        RECT 69.245 3.365 69.655 3.695 ;
        RECT 55.910 2.885 56.140 3.035 ;
        RECT 69.245 2.855 69.415 3.365 ;
        RECT 69.245 2.525 69.655 2.855 ;
        RECT 54.510 2.145 54.740 2.315 ;
        RECT 54.510 1.865 54.680 2.145 ;
        RECT 54.940 1.865 55.115 2.375 ;
        RECT 55.370 1.865 55.545 2.415 ;
        RECT 56.735 1.865 56.905 2.375 ;
        RECT 69.245 2.355 69.415 2.525 ;
        RECT 69.245 1.865 69.420 2.355 ;
        RECT 69.830 2.315 70.000 3.925 ;
        RECT 70.200 3.895 70.375 5.155 ;
        RECT 70.630 4.015 70.805 5.155 ;
        RECT 70.200 2.945 70.370 3.895 ;
        RECT 70.630 2.415 70.800 4.015 ;
        RECT 71.990 4.010 72.165 5.155 ;
        RECT 74.605 4.435 74.775 4.795 ;
        RECT 75.545 4.435 75.715 4.795 ;
        RECT 76.025 4.345 76.195 4.765 ;
        RECT 76.385 4.515 76.675 5.075 ;
        RECT 77.465 4.775 77.635 5.105 ;
        RECT 77.945 4.685 78.115 5.075 ;
        RECT 79.840 4.775 80.015 5.105 ;
        RECT 81.785 4.905 82.295 5.075 ;
        RECT 80.365 4.685 80.545 4.795 ;
        RECT 82.125 4.765 82.295 4.905 ;
        RECT 77.835 4.515 78.170 4.685 ;
        RECT 78.665 4.515 79.155 4.685 ;
        RECT 80.365 4.515 81.715 4.685 ;
        RECT 82.125 4.515 82.410 4.765 ;
        RECT 76.505 4.435 76.675 4.515 ;
        RECT 71.620 3.205 71.790 3.895 ;
        RECT 71.990 3.795 72.160 4.010 ;
        RECT 72.605 3.795 72.775 3.895 ;
        RECT 71.990 3.625 72.775 3.795 ;
        RECT 75.305 3.785 75.475 4.235 ;
        RECT 75.785 3.785 75.955 4.115 ;
        RECT 76.745 3.785 76.915 4.115 ;
        RECT 77.225 3.785 77.395 4.515 ;
        RECT 78.665 4.345 78.835 4.515 ;
        RECT 80.365 4.435 80.545 4.515 ;
        RECT 81.545 4.345 81.715 4.515 ;
        RECT 82.235 4.435 82.410 4.515 ;
        RECT 77.705 3.785 77.875 4.235 ;
        RECT 78.185 3.785 78.355 4.115 ;
        RECT 78.665 3.785 78.835 4.115 ;
        RECT 79.145 3.785 79.315 4.235 ;
        RECT 80.105 4.135 80.275 4.235 ;
        RECT 79.625 4.035 80.275 4.135 ;
        RECT 79.545 3.865 80.355 4.035 ;
        RECT 80.585 3.785 80.755 4.115 ;
        RECT 81.065 3.785 81.235 4.235 ;
        RECT 81.545 3.785 81.715 4.115 ;
        RECT 82.025 4.035 82.295 4.235 ;
        RECT 81.905 3.825 82.295 4.035 ;
        RECT 84.505 3.895 84.680 5.155 ;
        RECT 85.030 4.095 85.200 5.155 ;
        RECT 85.030 3.925 85.260 4.095 ;
        RECT 84.505 3.695 84.675 3.895 ;
        RECT 71.990 3.575 72.160 3.625 ;
        RECT 72.605 3.205 72.775 3.625 ;
        RECT 79.625 3.615 79.795 3.655 ;
        RECT 79.265 3.445 79.795 3.615 ;
        RECT 71.170 3.035 72.090 3.205 ;
        RECT 72.605 3.035 73.075 3.205 ;
        RECT 74.605 3.045 74.775 3.395 ;
        RECT 76.505 3.045 76.675 3.395 ;
        RECT 77.905 3.375 78.075 3.395 ;
        RECT 77.905 3.345 78.115 3.375 ;
        RECT 77.805 3.125 78.115 3.345 ;
        RECT 77.945 3.045 78.115 3.125 ;
        RECT 78.905 3.275 79.075 3.395 ;
        RECT 78.905 3.105 80.145 3.275 ;
        RECT 80.825 3.045 80.995 3.395 ;
        RECT 81.785 3.045 81.955 3.395 ;
        RECT 84.505 3.365 84.915 3.695 ;
        RECT 71.170 2.885 71.400 3.035 ;
        RECT 84.505 2.855 84.675 3.365 ;
        RECT 84.505 2.525 84.915 2.855 ;
        RECT 69.770 2.145 70.000 2.315 ;
        RECT 69.770 1.865 69.940 2.145 ;
        RECT 70.200 1.865 70.375 2.375 ;
        RECT 70.630 1.865 70.805 2.415 ;
        RECT 71.995 1.865 72.165 2.375 ;
        RECT 84.505 2.355 84.675 2.525 ;
        RECT 84.505 1.865 84.680 2.355 ;
        RECT 85.090 2.315 85.260 3.925 ;
        RECT 85.460 3.895 85.635 5.155 ;
        RECT 85.890 4.015 86.065 5.155 ;
        RECT 85.460 2.945 85.630 3.895 ;
        RECT 85.890 2.415 86.060 4.015 ;
        RECT 87.250 4.010 87.425 5.155 ;
        RECT 89.865 4.435 90.035 4.795 ;
        RECT 90.805 4.435 90.975 4.795 ;
        RECT 91.285 4.345 91.455 4.765 ;
        RECT 91.645 4.515 91.935 5.075 ;
        RECT 92.725 4.775 92.895 5.105 ;
        RECT 93.205 4.685 93.375 5.075 ;
        RECT 95.100 4.775 95.275 5.105 ;
        RECT 97.045 4.905 97.555 5.075 ;
        RECT 95.625 4.685 95.805 4.795 ;
        RECT 97.385 4.765 97.555 4.905 ;
        RECT 93.095 4.515 93.430 4.685 ;
        RECT 93.925 4.515 94.415 4.685 ;
        RECT 95.625 4.515 96.975 4.685 ;
        RECT 97.385 4.515 97.670 4.765 ;
        RECT 91.765 4.435 91.935 4.515 ;
        RECT 86.880 3.205 87.050 3.895 ;
        RECT 87.250 3.795 87.420 4.010 ;
        RECT 87.865 3.795 88.035 3.895 ;
        RECT 87.250 3.625 88.035 3.795 ;
        RECT 90.565 3.785 90.735 4.235 ;
        RECT 91.045 3.785 91.215 4.115 ;
        RECT 92.005 3.785 92.175 4.115 ;
        RECT 92.485 3.785 92.655 4.515 ;
        RECT 93.925 4.345 94.095 4.515 ;
        RECT 95.625 4.435 95.805 4.515 ;
        RECT 96.805 4.345 96.975 4.515 ;
        RECT 97.495 4.435 97.670 4.515 ;
        RECT 92.965 3.785 93.135 4.235 ;
        RECT 93.445 3.785 93.615 4.115 ;
        RECT 93.925 3.785 94.095 4.115 ;
        RECT 94.405 3.785 94.575 4.235 ;
        RECT 95.365 4.135 95.535 4.235 ;
        RECT 94.885 4.035 95.535 4.135 ;
        RECT 94.805 3.865 95.615 4.035 ;
        RECT 95.845 3.785 96.015 4.115 ;
        RECT 96.325 3.785 96.495 4.235 ;
        RECT 96.805 3.785 96.975 4.115 ;
        RECT 97.285 4.035 97.555 4.235 ;
        RECT 97.165 3.825 97.555 4.035 ;
        RECT 99.765 3.895 99.940 5.155 ;
        RECT 100.290 4.095 100.460 5.155 ;
        RECT 100.290 3.925 100.520 4.095 ;
        RECT 99.765 3.695 99.935 3.895 ;
        RECT 87.250 3.575 87.420 3.625 ;
        RECT 87.865 3.205 88.035 3.625 ;
        RECT 94.885 3.615 95.055 3.655 ;
        RECT 94.525 3.445 95.055 3.615 ;
        RECT 86.430 3.035 87.350 3.205 ;
        RECT 87.865 3.035 88.335 3.205 ;
        RECT 89.865 3.045 90.035 3.395 ;
        RECT 91.765 3.045 91.935 3.395 ;
        RECT 93.165 3.375 93.335 3.395 ;
        RECT 93.165 3.345 93.375 3.375 ;
        RECT 93.065 3.125 93.375 3.345 ;
        RECT 93.205 3.045 93.375 3.125 ;
        RECT 94.165 3.275 94.335 3.395 ;
        RECT 94.165 3.105 95.405 3.275 ;
        RECT 96.085 3.045 96.255 3.395 ;
        RECT 97.045 3.045 97.215 3.395 ;
        RECT 99.765 3.365 100.175 3.695 ;
        RECT 86.430 2.885 86.660 3.035 ;
        RECT 99.765 2.855 99.935 3.365 ;
        RECT 99.765 2.525 100.175 2.855 ;
        RECT 85.030 2.145 85.260 2.315 ;
        RECT 85.030 1.865 85.200 2.145 ;
        RECT 85.460 1.865 85.635 2.375 ;
        RECT 85.890 1.865 86.065 2.415 ;
        RECT 87.255 1.865 87.425 2.375 ;
        RECT 99.765 2.355 99.935 2.525 ;
        RECT 99.765 1.865 99.940 2.355 ;
        RECT 100.350 2.315 100.520 3.925 ;
        RECT 100.720 3.895 100.895 5.155 ;
        RECT 101.150 4.015 101.325 5.155 ;
        RECT 100.720 2.945 100.890 3.895 ;
        RECT 101.150 2.415 101.320 4.015 ;
        RECT 102.510 4.010 102.685 5.155 ;
        RECT 102.140 3.205 102.310 3.895 ;
        RECT 102.510 3.795 102.680 4.010 ;
        RECT 103.125 3.795 103.295 3.895 ;
        RECT 102.510 3.625 103.295 3.795 ;
        RECT 102.510 3.575 102.680 3.625 ;
        RECT 103.125 3.205 103.295 3.625 ;
        RECT 101.690 3.035 102.610 3.205 ;
        RECT 103.125 3.035 103.595 3.205 ;
        RECT 101.690 2.885 101.920 3.035 ;
        RECT 100.290 2.145 100.520 2.315 ;
        RECT 100.290 1.865 100.460 2.145 ;
        RECT 100.720 1.865 100.895 2.375 ;
        RECT 101.150 1.865 101.325 2.415 ;
        RECT 102.515 1.865 102.685 2.375 ;
      LAYER met1 ;
        RECT 26.490 10.060 26.780 10.290 ;
        RECT 34.005 10.060 34.295 10.290 ;
        RECT 39.620 10.060 39.910 10.290 ;
        RECT 26.550 9.610 26.720 10.060 ;
        RECT 34.065 9.715 34.235 10.060 ;
        RECT 26.460 9.320 26.810 9.610 ;
        RECT 33.965 9.345 34.335 9.715 ;
        RECT 39.680 9.580 39.850 10.060 ;
        RECT 41.410 10.030 41.705 10.290 ;
        RECT 42.400 10.030 42.695 10.290 ;
        RECT 49.265 10.060 49.555 10.290 ;
        RECT 54.880 10.060 55.170 10.290 ;
        RECT 40.590 9.580 40.940 9.610 ;
        RECT 39.680 9.550 40.940 9.580 ;
        RECT 39.620 9.410 40.940 9.550 ;
        RECT 34.005 9.320 34.295 9.345 ;
        RECT 39.620 9.320 39.910 9.410 ;
        RECT 40.590 9.320 40.940 9.410 ;
        RECT 34.635 9.180 34.985 9.245 ;
        RECT 40.075 9.180 40.400 9.270 ;
        RECT 34.435 9.150 34.985 9.180 ;
        RECT 40.050 9.150 40.400 9.180 ;
        RECT 34.265 9.145 34.985 9.150 ;
        RECT 39.880 9.145 40.400 9.150 ;
        RECT 34.265 8.980 40.400 9.145 ;
        RECT 34.325 8.975 40.400 8.980 ;
        RECT 34.435 8.950 34.985 8.975 ;
        RECT 40.050 8.950 40.400 8.975 ;
        RECT 34.635 8.895 34.985 8.950 ;
        RECT 40.075 8.945 40.400 8.950 ;
        RECT 41.470 8.930 41.640 10.030 ;
        RECT 42.460 9.300 42.630 10.030 ;
        RECT 49.325 9.715 49.495 10.060 ;
        RECT 49.225 9.345 49.595 9.715 ;
        RECT 54.940 9.580 55.110 10.060 ;
        RECT 56.670 10.030 56.965 10.290 ;
        RECT 57.660 10.030 57.955 10.290 ;
        RECT 64.525 10.060 64.815 10.290 ;
        RECT 70.140 10.060 70.430 10.290 ;
        RECT 55.850 9.580 56.200 9.610 ;
        RECT 54.940 9.550 56.200 9.580 ;
        RECT 54.880 9.410 56.200 9.550 ;
        RECT 49.265 9.320 49.555 9.345 ;
        RECT 54.880 9.320 55.170 9.410 ;
        RECT 55.850 9.320 56.200 9.410 ;
        RECT 42.455 8.950 42.805 9.300 ;
        RECT 49.895 9.180 50.245 9.255 ;
        RECT 55.335 9.180 55.660 9.270 ;
        RECT 49.695 9.150 50.245 9.180 ;
        RECT 55.310 9.150 55.660 9.180 ;
        RECT 49.525 9.145 50.245 9.150 ;
        RECT 55.140 9.145 55.660 9.150 ;
        RECT 49.525 8.980 55.660 9.145 ;
        RECT 49.585 8.975 55.660 8.980 ;
        RECT 49.695 8.950 50.245 8.975 ;
        RECT 55.310 8.950 55.660 8.975 ;
        RECT 42.455 8.930 42.750 8.950 ;
        RECT 41.410 8.925 41.640 8.930 ;
        RECT 26.085 8.790 26.435 8.865 ;
        RECT 39.275 8.820 39.595 8.835 ;
        RECT 39.250 8.790 39.595 8.820 ;
        RECT 25.945 8.620 26.435 8.790 ;
        RECT 39.075 8.620 39.595 8.790 ;
        RECT 41.410 8.690 41.700 8.925 ;
        RECT 42.400 8.865 42.750 8.930 ;
        RECT 49.895 8.905 50.245 8.950 ;
        RECT 55.335 8.945 55.660 8.950 ;
        RECT 56.730 8.930 56.900 10.030 ;
        RECT 57.720 9.305 57.890 10.030 ;
        RECT 64.585 9.715 64.755 10.060 ;
        RECT 64.485 9.345 64.855 9.715 ;
        RECT 70.200 9.580 70.370 10.060 ;
        RECT 71.930 10.030 72.225 10.290 ;
        RECT 72.920 10.030 73.215 10.290 ;
        RECT 79.785 10.060 80.075 10.290 ;
        RECT 85.400 10.060 85.690 10.290 ;
        RECT 71.110 9.580 71.460 9.610 ;
        RECT 70.200 9.550 71.460 9.580 ;
        RECT 70.140 9.410 71.460 9.550 ;
        RECT 64.525 9.320 64.815 9.345 ;
        RECT 70.140 9.320 70.430 9.410 ;
        RECT 71.110 9.320 71.460 9.410 ;
        RECT 57.710 8.950 58.065 9.305 ;
        RECT 65.155 9.180 65.505 9.255 ;
        RECT 70.595 9.180 70.920 9.270 ;
        RECT 64.955 9.150 65.505 9.180 ;
        RECT 70.570 9.150 70.920 9.180 ;
        RECT 64.785 9.145 65.505 9.150 ;
        RECT 70.400 9.145 70.920 9.150 ;
        RECT 64.785 8.980 70.920 9.145 ;
        RECT 64.845 8.975 70.920 8.980 ;
        RECT 64.955 8.950 65.505 8.975 ;
        RECT 70.570 8.950 70.920 8.975 ;
        RECT 57.710 8.930 58.010 8.950 ;
        RECT 56.670 8.925 56.900 8.930 ;
        RECT 42.400 8.690 42.690 8.865 ;
        RECT 54.535 8.820 54.855 8.835 ;
        RECT 54.510 8.790 54.855 8.820 ;
        RECT 54.335 8.620 54.855 8.790 ;
        RECT 56.670 8.690 56.960 8.925 ;
        RECT 57.660 8.860 58.010 8.930 ;
        RECT 65.155 8.905 65.505 8.950 ;
        RECT 70.595 8.945 70.920 8.950 ;
        RECT 71.990 8.930 72.160 10.030 ;
        RECT 72.980 9.300 73.150 10.030 ;
        RECT 79.845 9.715 80.015 10.060 ;
        RECT 79.745 9.345 80.115 9.715 ;
        RECT 85.460 9.580 85.630 10.060 ;
        RECT 87.190 10.030 87.485 10.290 ;
        RECT 88.180 10.030 88.475 10.290 ;
        RECT 95.045 10.060 95.335 10.290 ;
        RECT 100.660 10.060 100.950 10.290 ;
        RECT 86.370 9.580 86.720 9.610 ;
        RECT 85.460 9.550 86.720 9.580 ;
        RECT 85.400 9.410 86.720 9.550 ;
        RECT 79.785 9.320 80.075 9.345 ;
        RECT 85.400 9.320 85.690 9.410 ;
        RECT 86.370 9.320 86.720 9.410 ;
        RECT 72.930 8.950 73.280 9.300 ;
        RECT 80.420 9.180 80.770 9.255 ;
        RECT 85.855 9.180 86.180 9.270 ;
        RECT 80.215 9.150 80.770 9.180 ;
        RECT 85.830 9.150 86.180 9.180 ;
        RECT 80.045 9.145 80.770 9.150 ;
        RECT 85.660 9.145 86.180 9.150 ;
        RECT 80.045 8.980 86.180 9.145 ;
        RECT 80.105 8.975 86.180 8.980 ;
        RECT 80.215 8.950 80.770 8.975 ;
        RECT 85.830 8.950 86.180 8.975 ;
        RECT 72.930 8.930 73.270 8.950 ;
        RECT 71.930 8.925 72.160 8.930 ;
        RECT 57.660 8.690 57.950 8.860 ;
        RECT 69.795 8.820 70.115 8.835 ;
        RECT 69.770 8.790 70.115 8.820 ;
        RECT 69.595 8.620 70.115 8.790 ;
        RECT 71.930 8.690 72.220 8.925 ;
        RECT 72.920 8.860 73.270 8.930 ;
        RECT 80.420 8.905 80.770 8.950 ;
        RECT 85.855 8.945 86.180 8.950 ;
        RECT 87.250 8.930 87.420 10.030 ;
        RECT 88.240 9.300 88.410 10.030 ;
        RECT 95.105 9.715 95.275 10.060 ;
        RECT 95.005 9.345 95.375 9.715 ;
        RECT 100.720 9.580 100.890 10.060 ;
        RECT 102.450 10.030 102.745 10.290 ;
        RECT 103.440 10.030 103.735 10.290 ;
        RECT 101.630 9.580 101.980 9.610 ;
        RECT 100.720 9.550 101.980 9.580 ;
        RECT 100.660 9.410 101.980 9.550 ;
        RECT 95.045 9.320 95.335 9.345 ;
        RECT 100.660 9.320 100.950 9.410 ;
        RECT 101.630 9.320 101.980 9.410 ;
        RECT 88.190 8.950 88.540 9.300 ;
        RECT 95.675 9.180 96.025 9.255 ;
        RECT 101.115 9.180 101.440 9.270 ;
        RECT 95.475 9.150 96.025 9.180 ;
        RECT 101.090 9.150 101.440 9.180 ;
        RECT 95.305 9.145 96.025 9.150 ;
        RECT 100.920 9.145 101.440 9.150 ;
        RECT 95.305 8.980 101.440 9.145 ;
        RECT 95.365 8.975 101.440 8.980 ;
        RECT 95.475 8.950 96.025 8.975 ;
        RECT 101.090 8.950 101.440 8.975 ;
        RECT 88.190 8.930 88.530 8.950 ;
        RECT 87.190 8.925 87.420 8.930 ;
        RECT 72.920 8.690 73.210 8.860 ;
        RECT 85.055 8.820 85.375 8.835 ;
        RECT 85.030 8.790 85.375 8.820 ;
        RECT 84.855 8.620 85.375 8.790 ;
        RECT 87.190 8.690 87.480 8.925 ;
        RECT 88.180 8.860 88.530 8.930 ;
        RECT 95.675 8.905 96.025 8.950 ;
        RECT 101.115 8.945 101.440 8.950 ;
        RECT 102.510 8.930 102.680 10.030 ;
        RECT 103.475 9.995 103.735 10.030 ;
        RECT 103.475 9.915 103.795 9.995 ;
        RECT 103.475 9.565 103.825 9.915 ;
        RECT 103.500 8.930 103.670 9.565 ;
        RECT 102.450 8.925 102.680 8.930 ;
        RECT 103.440 8.925 103.670 8.930 ;
        RECT 88.180 8.690 88.470 8.860 ;
        RECT 100.315 8.820 100.635 8.835 ;
        RECT 100.290 8.790 100.635 8.820 ;
        RECT 100.115 8.620 100.635 8.790 ;
        RECT 102.450 8.690 102.740 8.925 ;
        RECT 103.440 8.690 103.730 8.925 ;
        RECT 26.085 8.575 26.435 8.620 ;
        RECT 39.250 8.590 39.595 8.620 ;
        RECT 54.510 8.590 54.855 8.620 ;
        RECT 69.770 8.590 70.115 8.620 ;
        RECT 85.030 8.590 85.375 8.620 ;
        RECT 100.290 8.590 100.635 8.620 ;
        RECT 39.275 8.545 39.595 8.590 ;
        RECT 54.535 8.545 54.855 8.590 ;
        RECT 69.795 8.545 70.115 8.590 ;
        RECT 85.055 8.545 85.375 8.590 ;
        RECT 100.315 8.545 100.635 8.590 ;
        RECT 30.665 4.895 30.955 5.105 ;
        RECT 29.775 4.875 30.955 4.895 ;
        RECT 28.755 4.585 29.075 4.845 ;
        RECT 29.775 4.825 30.875 4.875 ;
        RECT 31.605 4.865 31.925 5.125 ;
        RECT 32.205 5.105 32.525 5.125 ;
        RECT 32.105 4.875 32.525 5.105 ;
        RECT 32.205 4.865 32.525 4.875 ;
        RECT 33.765 5.105 34.100 5.125 ;
        RECT 33.765 4.875 34.290 5.105 ;
        RECT 35.945 5.065 36.235 5.105 ;
        RECT 36.375 5.065 36.695 5.125 ;
        RECT 35.945 4.925 36.695 5.065 ;
        RECT 35.945 4.875 36.235 4.925 ;
        RECT 33.765 4.865 34.100 4.875 ;
        RECT 36.375 4.865 36.695 4.925 ;
        RECT 45.925 4.895 46.215 5.105 ;
        RECT 45.035 4.875 46.215 4.895 ;
        RECT 29.705 4.755 30.875 4.825 ;
        RECT 29.705 4.595 29.995 4.755 ;
        RECT 32.135 4.585 32.305 4.685 ;
        RECT 34.515 4.585 34.835 4.845 ;
        RECT 44.015 4.585 44.335 4.845 ;
        RECT 45.035 4.825 46.135 4.875 ;
        RECT 46.865 4.865 47.185 5.125 ;
        RECT 47.465 5.105 47.785 5.125 ;
        RECT 47.365 4.875 47.785 5.105 ;
        RECT 47.465 4.865 47.785 4.875 ;
        RECT 49.025 5.105 49.360 5.125 ;
        RECT 49.025 4.875 49.550 5.105 ;
        RECT 51.205 5.065 51.495 5.105 ;
        RECT 51.635 5.065 51.955 5.125 ;
        RECT 51.205 4.925 51.955 5.065 ;
        RECT 51.205 4.875 51.495 4.925 ;
        RECT 49.025 4.865 49.360 4.875 ;
        RECT 51.635 4.865 51.955 4.925 ;
        RECT 61.185 4.895 61.475 5.105 ;
        RECT 60.295 4.875 61.475 4.895 ;
        RECT 44.965 4.755 46.135 4.825 ;
        RECT 44.965 4.595 45.255 4.755 ;
        RECT 47.395 4.585 47.565 4.685 ;
        RECT 49.775 4.585 50.095 4.845 ;
        RECT 59.275 4.585 59.595 4.845 ;
        RECT 60.295 4.825 61.395 4.875 ;
        RECT 62.125 4.865 62.445 5.125 ;
        RECT 62.725 5.105 63.045 5.125 ;
        RECT 62.625 4.875 63.045 5.105 ;
        RECT 62.725 4.865 63.045 4.875 ;
        RECT 64.285 5.105 64.620 5.125 ;
        RECT 64.285 4.875 64.810 5.105 ;
        RECT 66.465 5.065 66.755 5.105 ;
        RECT 66.895 5.065 67.215 5.125 ;
        RECT 66.465 4.925 67.215 5.065 ;
        RECT 66.465 4.875 66.755 4.925 ;
        RECT 64.285 4.865 64.620 4.875 ;
        RECT 66.895 4.865 67.215 4.925 ;
        RECT 76.445 4.895 76.735 5.105 ;
        RECT 75.555 4.875 76.735 4.895 ;
        RECT 60.225 4.755 61.395 4.825 ;
        RECT 60.225 4.595 60.515 4.755 ;
        RECT 62.655 4.585 62.825 4.685 ;
        RECT 65.035 4.585 65.355 4.845 ;
        RECT 74.535 4.585 74.855 4.845 ;
        RECT 75.555 4.825 76.655 4.875 ;
        RECT 77.385 4.865 77.705 5.125 ;
        RECT 77.985 5.105 78.305 5.125 ;
        RECT 77.885 4.875 78.305 5.105 ;
        RECT 77.985 4.865 78.305 4.875 ;
        RECT 79.545 5.105 79.880 5.125 ;
        RECT 79.545 4.875 80.070 5.105 ;
        RECT 81.725 5.065 82.015 5.105 ;
        RECT 82.155 5.065 82.475 5.125 ;
        RECT 81.725 4.925 82.475 5.065 ;
        RECT 81.725 4.875 82.015 4.925 ;
        RECT 79.545 4.865 79.880 4.875 ;
        RECT 82.155 4.865 82.475 4.925 ;
        RECT 91.705 4.895 91.995 5.105 ;
        RECT 90.815 4.875 91.995 4.895 ;
        RECT 75.485 4.755 76.655 4.825 ;
        RECT 75.485 4.595 75.775 4.755 ;
        RECT 77.915 4.585 78.085 4.685 ;
        RECT 80.295 4.585 80.615 4.845 ;
        RECT 89.795 4.585 90.115 4.845 ;
        RECT 90.815 4.825 91.915 4.875 ;
        RECT 92.645 4.865 92.965 5.125 ;
        RECT 93.245 5.105 93.565 5.125 ;
        RECT 93.145 4.875 93.565 5.105 ;
        RECT 93.245 4.865 93.565 4.875 ;
        RECT 94.805 5.105 95.140 5.125 ;
        RECT 94.805 4.875 95.330 5.105 ;
        RECT 96.985 5.065 97.275 5.105 ;
        RECT 97.415 5.065 97.735 5.125 ;
        RECT 96.985 4.925 97.735 5.065 ;
        RECT 96.985 4.875 97.275 4.925 ;
        RECT 94.805 4.865 95.140 4.875 ;
        RECT 97.415 4.865 97.735 4.925 ;
        RECT 90.745 4.755 91.915 4.825 ;
        RECT 90.745 4.595 91.035 4.755 ;
        RECT 93.175 4.585 93.345 4.685 ;
        RECT 95.555 4.585 95.875 4.845 ;
        RECT 31.125 4.545 31.445 4.565 ;
        RECT 30.185 4.505 30.475 4.545 ;
        RECT 30.185 4.315 30.635 4.505 ;
        RECT 29.445 4.025 29.765 4.285 ;
        RECT 29.925 3.745 30.245 4.005 ;
        RECT 30.495 3.985 30.635 4.315 ;
        RECT 31.125 4.315 31.675 4.545 ;
        RECT 31.815 4.445 33.995 4.585 ;
        RECT 46.385 4.545 46.705 4.565 ;
        RECT 31.815 4.365 33.115 4.445 ;
        RECT 31.125 4.305 31.445 4.315 ;
        RECT 31.815 4.085 32.155 4.365 ;
        RECT 32.825 4.315 33.115 4.365 ;
        RECT 31.865 4.035 32.155 4.085 ;
        RECT 33.285 4.025 33.605 4.285 ;
        RECT 30.495 3.845 30.755 3.985 ;
        RECT 28.755 3.185 29.075 3.445 ;
        RECT 30.615 3.425 30.755 3.845 ;
        RECT 30.905 3.945 31.195 3.985 ;
        RECT 31.365 3.945 31.685 4.005 ;
        RECT 30.905 3.805 31.685 3.945 ;
        RECT 30.905 3.755 31.195 3.805 ;
        RECT 31.365 3.745 31.685 3.805 ;
        RECT 32.345 3.755 32.635 3.985 ;
        RECT 32.495 3.505 32.635 3.755 ;
        RECT 32.805 3.745 33.125 4.005 ;
        RECT 33.855 3.805 33.995 4.445 ;
        RECT 35.705 4.505 35.995 4.545 ;
        RECT 45.445 4.505 45.735 4.545 ;
        RECT 35.705 4.365 36.275 4.505 ;
        RECT 34.335 4.285 35.435 4.365 ;
        RECT 35.705 4.315 35.995 4.365 ;
        RECT 34.145 4.265 35.435 4.285 ;
        RECT 36.135 4.265 36.395 4.365 ;
        RECT 34.145 4.225 35.515 4.265 ;
        RECT 36.135 4.225 36.475 4.265 ;
        RECT 34.145 4.035 34.555 4.225 ;
        RECT 35.225 4.035 35.515 4.225 ;
        RECT 36.185 4.035 36.475 4.225 ;
        RECT 34.145 4.025 34.465 4.035 ;
        RECT 34.745 3.805 35.035 3.985 ;
        RECT 33.855 3.755 35.035 3.805 ;
        RECT 33.855 3.705 34.955 3.755 ;
        RECT 35.685 3.745 36.005 4.005 ;
        RECT 37.670 3.995 38.010 4.345 ;
        RECT 45.445 4.315 45.895 4.505 ;
        RECT 44.705 4.025 45.025 4.285 ;
        RECT 33.785 3.665 34.955 3.705 ;
        RECT 32.495 3.445 32.795 3.505 ;
        RECT 33.785 3.455 34.075 3.665 ;
        RECT 37.760 3.490 37.930 3.995 ;
        RECT 39.275 3.875 39.595 3.980 ;
        RECT 39.250 3.860 39.595 3.875 ;
        RECT 39.240 3.845 39.595 3.860 ;
        RECT 39.075 3.675 39.595 3.845 ;
        RECT 39.250 3.660 39.595 3.675 ;
        RECT 39.250 3.645 39.540 3.660 ;
        RECT 40.050 3.490 40.400 3.610 ;
        RECT 41.410 3.540 41.700 3.775 ;
        RECT 45.185 3.745 45.505 4.005 ;
        RECT 45.755 3.985 45.895 4.315 ;
        RECT 46.385 4.315 46.935 4.545 ;
        RECT 47.075 4.445 49.255 4.585 ;
        RECT 61.645 4.545 61.965 4.565 ;
        RECT 47.075 4.365 48.375 4.445 ;
        RECT 46.385 4.305 46.705 4.315 ;
        RECT 47.075 4.085 47.415 4.365 ;
        RECT 48.085 4.315 48.375 4.365 ;
        RECT 47.125 4.035 47.415 4.085 ;
        RECT 48.545 4.025 48.865 4.285 ;
        RECT 45.755 3.845 46.015 3.985 ;
        RECT 41.410 3.535 41.640 3.540 ;
        RECT 30.615 3.385 30.955 3.425 ;
        RECT 31.485 3.385 31.805 3.445 ;
        RECT 30.615 3.245 31.805 3.385 ;
        RECT 30.665 3.195 30.955 3.245 ;
        RECT 31.485 3.185 31.805 3.245 ;
        RECT 31.955 3.185 32.355 3.445 ;
        RECT 32.495 3.385 32.885 3.445 ;
        RECT 33.285 3.425 33.605 3.445 ;
        RECT 33.065 3.385 33.605 3.425 ;
        RECT 32.495 3.365 33.605 3.385 ;
        RECT 32.565 3.245 33.605 3.365 ;
        RECT 32.565 3.185 32.885 3.245 ;
        RECT 33.065 3.195 33.605 3.245 ;
        RECT 33.285 3.185 33.605 3.195 ;
        RECT 34.515 3.385 34.835 3.445 ;
        RECT 34.985 3.385 35.275 3.425 ;
        RECT 34.515 3.245 35.275 3.385 ;
        RECT 34.515 3.185 34.835 3.245 ;
        RECT 34.985 3.195 35.275 3.245 ;
        RECT 35.945 3.385 36.235 3.425 ;
        RECT 36.375 3.385 36.695 3.445 ;
        RECT 35.945 3.245 36.695 3.385 ;
        RECT 37.760 3.320 40.400 3.490 ;
        RECT 39.880 3.315 40.400 3.320 ;
        RECT 40.050 3.260 40.400 3.315 ;
        RECT 35.945 3.195 36.235 3.245 ;
        RECT 36.375 3.185 36.695 3.245 ;
        RECT 39.620 3.120 39.910 3.145 ;
        RECT 40.590 3.120 40.940 3.145 ;
        RECT 39.620 2.950 40.940 3.120 ;
        RECT 39.620 2.915 39.910 2.950 ;
        RECT 39.680 2.405 39.850 2.915 ;
        RECT 40.590 2.855 40.940 2.950 ;
        RECT 41.470 2.435 41.640 3.535 ;
        RECT 44.015 3.185 44.335 3.445 ;
        RECT 45.875 3.425 46.015 3.845 ;
        RECT 46.165 3.945 46.455 3.985 ;
        RECT 46.625 3.945 46.945 4.005 ;
        RECT 46.165 3.805 46.945 3.945 ;
        RECT 46.165 3.755 46.455 3.805 ;
        RECT 46.625 3.745 46.945 3.805 ;
        RECT 47.605 3.755 47.895 3.985 ;
        RECT 47.755 3.505 47.895 3.755 ;
        RECT 48.065 3.745 48.385 4.005 ;
        RECT 49.115 3.805 49.255 4.445 ;
        RECT 50.965 4.505 51.255 4.545 ;
        RECT 60.705 4.505 60.995 4.545 ;
        RECT 50.965 4.365 51.535 4.505 ;
        RECT 49.595 4.285 50.695 4.365 ;
        RECT 50.965 4.315 51.255 4.365 ;
        RECT 49.405 4.265 50.695 4.285 ;
        RECT 51.395 4.265 51.655 4.365 ;
        RECT 49.405 4.225 50.775 4.265 ;
        RECT 51.395 4.225 51.735 4.265 ;
        RECT 49.405 4.035 49.815 4.225 ;
        RECT 50.485 4.035 50.775 4.225 ;
        RECT 51.445 4.035 51.735 4.225 ;
        RECT 49.405 4.025 49.725 4.035 ;
        RECT 50.005 3.805 50.295 3.985 ;
        RECT 49.115 3.755 50.295 3.805 ;
        RECT 49.115 3.705 50.215 3.755 ;
        RECT 50.945 3.745 51.265 4.005 ;
        RECT 52.930 3.995 53.270 4.345 ;
        RECT 60.705 4.315 61.155 4.505 ;
        RECT 59.965 4.025 60.285 4.285 ;
        RECT 49.045 3.665 50.215 3.705 ;
        RECT 47.755 3.445 48.055 3.505 ;
        RECT 49.045 3.455 49.335 3.665 ;
        RECT 53.020 3.490 53.190 3.995 ;
        RECT 54.535 3.875 54.855 3.980 ;
        RECT 54.510 3.860 54.855 3.875 ;
        RECT 54.500 3.845 54.855 3.860 ;
        RECT 54.335 3.675 54.855 3.845 ;
        RECT 54.510 3.660 54.855 3.675 ;
        RECT 54.510 3.645 54.800 3.660 ;
        RECT 55.310 3.490 55.660 3.610 ;
        RECT 56.670 3.540 56.960 3.775 ;
        RECT 60.445 3.745 60.765 4.005 ;
        RECT 61.015 3.985 61.155 4.315 ;
        RECT 61.645 4.315 62.195 4.545 ;
        RECT 62.335 4.445 64.515 4.585 ;
        RECT 76.905 4.545 77.225 4.565 ;
        RECT 62.335 4.365 63.635 4.445 ;
        RECT 61.645 4.305 61.965 4.315 ;
        RECT 62.335 4.085 62.675 4.365 ;
        RECT 63.345 4.315 63.635 4.365 ;
        RECT 62.385 4.035 62.675 4.085 ;
        RECT 63.805 4.025 64.125 4.285 ;
        RECT 61.015 3.845 61.275 3.985 ;
        RECT 56.670 3.535 56.900 3.540 ;
        RECT 45.875 3.385 46.215 3.425 ;
        RECT 46.745 3.385 47.065 3.445 ;
        RECT 45.875 3.245 47.065 3.385 ;
        RECT 45.925 3.195 46.215 3.245 ;
        RECT 46.745 3.185 47.065 3.245 ;
        RECT 47.215 3.185 47.615 3.445 ;
        RECT 47.755 3.385 48.145 3.445 ;
        RECT 48.545 3.425 48.865 3.445 ;
        RECT 48.325 3.385 48.865 3.425 ;
        RECT 47.755 3.365 48.865 3.385 ;
        RECT 47.825 3.245 48.865 3.365 ;
        RECT 47.825 3.185 48.145 3.245 ;
        RECT 48.325 3.195 48.865 3.245 ;
        RECT 48.545 3.185 48.865 3.195 ;
        RECT 49.775 3.385 50.095 3.445 ;
        RECT 50.245 3.385 50.535 3.425 ;
        RECT 49.775 3.245 50.535 3.385 ;
        RECT 49.775 3.185 50.095 3.245 ;
        RECT 50.245 3.195 50.535 3.245 ;
        RECT 51.205 3.385 51.495 3.425 ;
        RECT 51.635 3.385 51.955 3.445 ;
        RECT 51.205 3.245 51.955 3.385 ;
        RECT 53.020 3.320 55.660 3.490 ;
        RECT 55.140 3.315 55.660 3.320 ;
        RECT 55.310 3.260 55.660 3.315 ;
        RECT 51.205 3.195 51.495 3.245 ;
        RECT 51.635 3.185 51.955 3.245 ;
        RECT 54.880 3.120 55.170 3.145 ;
        RECT 55.850 3.120 56.200 3.145 ;
        RECT 54.880 2.950 56.200 3.120 ;
        RECT 54.880 2.915 55.170 2.950 ;
        RECT 39.620 2.175 39.910 2.405 ;
        RECT 41.410 2.175 41.705 2.435 ;
        RECT 54.940 2.405 55.110 2.915 ;
        RECT 55.850 2.855 56.200 2.950 ;
        RECT 56.730 2.435 56.900 3.535 ;
        RECT 59.275 3.185 59.595 3.445 ;
        RECT 61.135 3.425 61.275 3.845 ;
        RECT 61.425 3.945 61.715 3.985 ;
        RECT 61.885 3.945 62.205 4.005 ;
        RECT 61.425 3.805 62.205 3.945 ;
        RECT 61.425 3.755 61.715 3.805 ;
        RECT 61.885 3.745 62.205 3.805 ;
        RECT 62.865 3.755 63.155 3.985 ;
        RECT 63.015 3.505 63.155 3.755 ;
        RECT 63.325 3.745 63.645 4.005 ;
        RECT 64.375 3.805 64.515 4.445 ;
        RECT 66.225 4.505 66.515 4.545 ;
        RECT 75.965 4.505 76.255 4.545 ;
        RECT 66.225 4.365 66.795 4.505 ;
        RECT 64.855 4.285 65.955 4.365 ;
        RECT 66.225 4.315 66.515 4.365 ;
        RECT 64.665 4.265 65.955 4.285 ;
        RECT 66.655 4.265 66.915 4.365 ;
        RECT 64.665 4.225 66.035 4.265 ;
        RECT 66.655 4.225 66.995 4.265 ;
        RECT 64.665 4.035 65.075 4.225 ;
        RECT 65.745 4.035 66.035 4.225 ;
        RECT 66.705 4.035 66.995 4.225 ;
        RECT 64.665 4.025 64.985 4.035 ;
        RECT 65.265 3.805 65.555 3.985 ;
        RECT 64.375 3.755 65.555 3.805 ;
        RECT 64.375 3.705 65.475 3.755 ;
        RECT 66.205 3.745 66.525 4.005 ;
        RECT 68.190 3.995 68.530 4.345 ;
        RECT 75.965 4.315 76.415 4.505 ;
        RECT 75.225 4.025 75.545 4.285 ;
        RECT 64.305 3.665 65.475 3.705 ;
        RECT 63.015 3.445 63.315 3.505 ;
        RECT 64.305 3.455 64.595 3.665 ;
        RECT 68.280 3.490 68.450 3.995 ;
        RECT 69.795 3.875 70.115 3.980 ;
        RECT 69.770 3.860 70.115 3.875 ;
        RECT 69.760 3.845 70.115 3.860 ;
        RECT 69.595 3.675 70.115 3.845 ;
        RECT 69.770 3.660 70.115 3.675 ;
        RECT 69.770 3.645 70.060 3.660 ;
        RECT 70.570 3.490 70.920 3.610 ;
        RECT 71.930 3.540 72.220 3.775 ;
        RECT 75.705 3.745 76.025 4.005 ;
        RECT 76.275 3.985 76.415 4.315 ;
        RECT 76.905 4.315 77.455 4.545 ;
        RECT 77.595 4.445 79.775 4.585 ;
        RECT 92.165 4.545 92.485 4.565 ;
        RECT 77.595 4.365 78.895 4.445 ;
        RECT 76.905 4.305 77.225 4.315 ;
        RECT 77.595 4.085 77.935 4.365 ;
        RECT 78.605 4.315 78.895 4.365 ;
        RECT 77.645 4.035 77.935 4.085 ;
        RECT 79.065 4.025 79.385 4.285 ;
        RECT 76.275 3.845 76.535 3.985 ;
        RECT 71.930 3.535 72.160 3.540 ;
        RECT 61.135 3.385 61.475 3.425 ;
        RECT 62.005 3.385 62.325 3.445 ;
        RECT 61.135 3.245 62.325 3.385 ;
        RECT 61.185 3.195 61.475 3.245 ;
        RECT 62.005 3.185 62.325 3.245 ;
        RECT 62.475 3.185 62.875 3.445 ;
        RECT 63.015 3.385 63.405 3.445 ;
        RECT 63.805 3.425 64.125 3.445 ;
        RECT 63.585 3.385 64.125 3.425 ;
        RECT 63.015 3.365 64.125 3.385 ;
        RECT 63.085 3.245 64.125 3.365 ;
        RECT 63.085 3.185 63.405 3.245 ;
        RECT 63.585 3.195 64.125 3.245 ;
        RECT 63.805 3.185 64.125 3.195 ;
        RECT 65.035 3.385 65.355 3.445 ;
        RECT 65.505 3.385 65.795 3.425 ;
        RECT 65.035 3.245 65.795 3.385 ;
        RECT 65.035 3.185 65.355 3.245 ;
        RECT 65.505 3.195 65.795 3.245 ;
        RECT 66.465 3.385 66.755 3.425 ;
        RECT 66.895 3.385 67.215 3.445 ;
        RECT 66.465 3.245 67.215 3.385 ;
        RECT 68.280 3.320 70.920 3.490 ;
        RECT 70.400 3.315 70.920 3.320 ;
        RECT 70.570 3.260 70.920 3.315 ;
        RECT 66.465 3.195 66.755 3.245 ;
        RECT 66.895 3.185 67.215 3.245 ;
        RECT 70.140 3.120 70.430 3.145 ;
        RECT 71.110 3.120 71.460 3.145 ;
        RECT 70.140 2.950 71.460 3.120 ;
        RECT 70.140 2.915 70.430 2.950 ;
        RECT 54.880 2.175 55.170 2.405 ;
        RECT 56.670 2.175 56.965 2.435 ;
        RECT 70.200 2.405 70.370 2.915 ;
        RECT 71.110 2.855 71.460 2.950 ;
        RECT 71.990 2.435 72.160 3.535 ;
        RECT 74.535 3.185 74.855 3.445 ;
        RECT 76.395 3.425 76.535 3.845 ;
        RECT 76.685 3.945 76.975 3.985 ;
        RECT 77.145 3.945 77.465 4.005 ;
        RECT 76.685 3.805 77.465 3.945 ;
        RECT 76.685 3.755 76.975 3.805 ;
        RECT 77.145 3.745 77.465 3.805 ;
        RECT 78.125 3.755 78.415 3.985 ;
        RECT 78.275 3.505 78.415 3.755 ;
        RECT 78.585 3.745 78.905 4.005 ;
        RECT 79.635 3.805 79.775 4.445 ;
        RECT 81.485 4.505 81.775 4.545 ;
        RECT 91.225 4.505 91.515 4.545 ;
        RECT 81.485 4.365 82.055 4.505 ;
        RECT 80.115 4.285 81.215 4.365 ;
        RECT 81.485 4.315 81.775 4.365 ;
        RECT 79.925 4.265 81.215 4.285 ;
        RECT 81.915 4.265 82.175 4.365 ;
        RECT 79.925 4.225 81.295 4.265 ;
        RECT 81.915 4.225 82.255 4.265 ;
        RECT 79.925 4.035 80.335 4.225 ;
        RECT 81.005 4.035 81.295 4.225 ;
        RECT 81.965 4.035 82.255 4.225 ;
        RECT 79.925 4.025 80.245 4.035 ;
        RECT 80.525 3.805 80.815 3.985 ;
        RECT 79.635 3.755 80.815 3.805 ;
        RECT 79.635 3.705 80.735 3.755 ;
        RECT 81.465 3.745 81.785 4.005 ;
        RECT 83.450 3.995 83.790 4.345 ;
        RECT 91.225 4.315 91.675 4.505 ;
        RECT 90.485 4.025 90.805 4.285 ;
        RECT 79.565 3.665 80.735 3.705 ;
        RECT 78.275 3.445 78.575 3.505 ;
        RECT 79.565 3.455 79.855 3.665 ;
        RECT 83.540 3.490 83.710 3.995 ;
        RECT 85.055 3.875 85.375 3.980 ;
        RECT 85.030 3.860 85.375 3.875 ;
        RECT 85.020 3.845 85.375 3.860 ;
        RECT 84.855 3.675 85.375 3.845 ;
        RECT 85.030 3.660 85.375 3.675 ;
        RECT 85.030 3.645 85.320 3.660 ;
        RECT 85.830 3.490 86.180 3.610 ;
        RECT 87.190 3.540 87.480 3.775 ;
        RECT 90.965 3.745 91.285 4.005 ;
        RECT 91.535 3.985 91.675 4.315 ;
        RECT 92.165 4.315 92.715 4.545 ;
        RECT 92.855 4.445 95.035 4.585 ;
        RECT 92.855 4.365 94.155 4.445 ;
        RECT 92.165 4.305 92.485 4.315 ;
        RECT 92.855 4.085 93.195 4.365 ;
        RECT 93.865 4.315 94.155 4.365 ;
        RECT 92.905 4.035 93.195 4.085 ;
        RECT 94.325 4.025 94.645 4.285 ;
        RECT 91.535 3.845 91.795 3.985 ;
        RECT 87.190 3.535 87.420 3.540 ;
        RECT 76.395 3.385 76.735 3.425 ;
        RECT 77.265 3.385 77.585 3.445 ;
        RECT 76.395 3.245 77.585 3.385 ;
        RECT 76.445 3.195 76.735 3.245 ;
        RECT 77.265 3.185 77.585 3.245 ;
        RECT 77.735 3.185 78.135 3.445 ;
        RECT 78.275 3.385 78.665 3.445 ;
        RECT 79.065 3.425 79.385 3.445 ;
        RECT 78.845 3.385 79.385 3.425 ;
        RECT 78.275 3.365 79.385 3.385 ;
        RECT 78.345 3.245 79.385 3.365 ;
        RECT 78.345 3.185 78.665 3.245 ;
        RECT 78.845 3.195 79.385 3.245 ;
        RECT 79.065 3.185 79.385 3.195 ;
        RECT 80.295 3.385 80.615 3.445 ;
        RECT 80.765 3.385 81.055 3.425 ;
        RECT 80.295 3.245 81.055 3.385 ;
        RECT 80.295 3.185 80.615 3.245 ;
        RECT 80.765 3.195 81.055 3.245 ;
        RECT 81.725 3.385 82.015 3.425 ;
        RECT 82.155 3.385 82.475 3.445 ;
        RECT 81.725 3.245 82.475 3.385 ;
        RECT 83.540 3.320 86.180 3.490 ;
        RECT 85.660 3.315 86.180 3.320 ;
        RECT 85.830 3.260 86.180 3.315 ;
        RECT 81.725 3.195 82.015 3.245 ;
        RECT 82.155 3.185 82.475 3.245 ;
        RECT 85.400 3.120 85.690 3.145 ;
        RECT 86.370 3.120 86.720 3.145 ;
        RECT 85.400 2.950 86.720 3.120 ;
        RECT 85.400 2.915 85.690 2.950 ;
        RECT 70.140 2.175 70.430 2.405 ;
        RECT 71.930 2.175 72.225 2.435 ;
        RECT 85.460 2.405 85.630 2.915 ;
        RECT 86.370 2.855 86.720 2.950 ;
        RECT 87.250 2.435 87.420 3.535 ;
        RECT 89.795 3.185 90.115 3.445 ;
        RECT 91.655 3.425 91.795 3.845 ;
        RECT 91.945 3.945 92.235 3.985 ;
        RECT 92.405 3.945 92.725 4.005 ;
        RECT 91.945 3.805 92.725 3.945 ;
        RECT 91.945 3.755 92.235 3.805 ;
        RECT 92.405 3.745 92.725 3.805 ;
        RECT 93.385 3.755 93.675 3.985 ;
        RECT 93.535 3.505 93.675 3.755 ;
        RECT 93.845 3.745 94.165 4.005 ;
        RECT 94.895 3.805 95.035 4.445 ;
        RECT 96.745 4.505 97.035 4.545 ;
        RECT 96.745 4.365 97.315 4.505 ;
        RECT 95.375 4.285 96.475 4.365 ;
        RECT 96.745 4.315 97.035 4.365 ;
        RECT 95.185 4.265 96.475 4.285 ;
        RECT 97.175 4.265 97.435 4.365 ;
        RECT 95.185 4.225 96.555 4.265 ;
        RECT 97.175 4.225 97.515 4.265 ;
        RECT 95.185 4.035 95.595 4.225 ;
        RECT 96.265 4.035 96.555 4.225 ;
        RECT 97.225 4.035 97.515 4.225 ;
        RECT 95.185 4.025 95.505 4.035 ;
        RECT 95.785 3.805 96.075 3.985 ;
        RECT 94.895 3.755 96.075 3.805 ;
        RECT 94.895 3.705 95.995 3.755 ;
        RECT 96.725 3.745 97.045 4.005 ;
        RECT 98.710 3.995 99.050 4.345 ;
        RECT 94.825 3.665 95.995 3.705 ;
        RECT 93.535 3.445 93.835 3.505 ;
        RECT 94.825 3.455 95.115 3.665 ;
        RECT 98.800 3.490 98.970 3.995 ;
        RECT 100.315 3.875 100.635 3.980 ;
        RECT 100.290 3.860 100.635 3.875 ;
        RECT 100.280 3.845 100.635 3.860 ;
        RECT 100.115 3.675 100.635 3.845 ;
        RECT 100.290 3.660 100.635 3.675 ;
        RECT 100.290 3.645 100.580 3.660 ;
        RECT 101.090 3.490 101.440 3.610 ;
        RECT 102.450 3.540 102.740 3.775 ;
        RECT 102.450 3.535 102.680 3.540 ;
        RECT 91.655 3.385 91.995 3.425 ;
        RECT 92.525 3.385 92.845 3.445 ;
        RECT 91.655 3.245 92.845 3.385 ;
        RECT 91.705 3.195 91.995 3.245 ;
        RECT 92.525 3.185 92.845 3.245 ;
        RECT 92.995 3.185 93.395 3.445 ;
        RECT 93.535 3.385 93.925 3.445 ;
        RECT 94.325 3.425 94.645 3.445 ;
        RECT 94.105 3.385 94.645 3.425 ;
        RECT 93.535 3.365 94.645 3.385 ;
        RECT 93.605 3.245 94.645 3.365 ;
        RECT 93.605 3.185 93.925 3.245 ;
        RECT 94.105 3.195 94.645 3.245 ;
        RECT 94.325 3.185 94.645 3.195 ;
        RECT 95.555 3.385 95.875 3.445 ;
        RECT 96.025 3.385 96.315 3.425 ;
        RECT 95.555 3.245 96.315 3.385 ;
        RECT 95.555 3.185 95.875 3.245 ;
        RECT 96.025 3.195 96.315 3.245 ;
        RECT 96.985 3.385 97.275 3.425 ;
        RECT 97.415 3.385 97.735 3.445 ;
        RECT 96.985 3.245 97.735 3.385 ;
        RECT 98.800 3.320 101.440 3.490 ;
        RECT 100.920 3.315 101.440 3.320 ;
        RECT 101.090 3.260 101.440 3.315 ;
        RECT 96.985 3.195 97.275 3.245 ;
        RECT 97.415 3.185 97.735 3.245 ;
        RECT 100.660 3.120 100.950 3.145 ;
        RECT 101.630 3.120 101.980 3.145 ;
        RECT 100.660 2.950 101.980 3.120 ;
        RECT 100.660 2.915 100.950 2.950 ;
        RECT 85.400 2.175 85.690 2.405 ;
        RECT 87.190 2.175 87.485 2.435 ;
        RECT 100.720 2.405 100.890 2.915 ;
        RECT 101.630 2.855 101.980 2.950 ;
        RECT 102.510 2.435 102.680 3.535 ;
        RECT 100.660 2.175 100.950 2.405 ;
        RECT 102.450 2.175 102.745 2.435 ;
      LAYER met2 ;
        RECT 26.175 10.690 103.675 10.860 ;
        RECT 26.175 8.895 26.345 10.690 ;
        RECT 103.505 9.915 103.675 10.690 ;
        RECT 26.490 9.530 26.780 9.640 ;
        RECT 26.490 9.525 26.810 9.530 ;
        RECT 26.490 9.355 27.710 9.525 ;
        RECT 26.490 9.290 26.780 9.355 ;
        RECT 27.540 9.145 27.710 9.355 ;
        RECT 33.965 9.345 34.335 9.715 ;
        RECT 49.225 9.345 49.595 9.715 ;
        RECT 64.485 9.345 64.855 9.715 ;
        RECT 79.745 9.345 80.115 9.715 ;
        RECT 95.005 9.345 95.375 9.715 ;
        RECT 103.475 9.565 103.825 9.915 ;
        RECT 34.635 9.145 34.985 9.245 ;
        RECT 40.075 9.205 40.400 9.270 ;
        RECT 27.540 8.975 34.985 9.145 ;
        RECT 34.635 8.895 34.985 8.975 ;
        RECT 38.960 9.035 40.400 9.205 ;
        RECT 26.115 8.545 26.405 8.895 ;
        RECT 31.935 5.305 34.375 5.445 ;
        RECT 31.935 5.155 32.075 5.305 ;
        RECT 31.635 5.065 32.075 5.155 ;
        RECT 29.295 4.925 32.075 5.065 ;
        RECT 28.785 4.785 29.045 4.875 ;
        RECT 29.295 4.785 29.435 4.925 ;
        RECT 31.635 4.835 31.895 4.925 ;
        RECT 32.235 4.835 32.495 5.155 ;
        RECT 32.235 4.785 32.435 4.835 ;
        RECT 28.785 4.645 29.435 4.785 ;
        RECT 32.045 4.645 32.435 4.785 ;
        RECT 33.305 4.775 33.585 5.155 ;
        RECT 33.795 4.835 34.070 5.155 ;
        RECT 28.785 4.555 29.045 4.645 ;
        RECT 28.845 3.475 28.985 4.555 ;
        RECT 29.705 4.505 29.985 4.620 ;
        RECT 31.155 4.505 31.415 4.595 ;
        RECT 29.535 4.365 31.415 4.505 ;
        RECT 29.535 4.315 29.985 4.365 ;
        RECT 29.475 4.245 29.985 4.315 ;
        RECT 31.155 4.275 31.415 4.365 ;
        RECT 29.475 4.055 29.735 4.245 ;
        RECT 30.650 4.055 30.955 4.060 ;
        RECT 29.465 3.685 29.745 4.055 ;
        RECT 29.955 3.945 30.215 4.035 ;
        RECT 30.545 3.945 30.955 4.055 ;
        RECT 29.955 3.805 30.955 3.945 ;
        RECT 29.955 3.715 30.215 3.805 ;
        RECT 30.545 3.685 30.955 3.805 ;
        RECT 31.385 3.685 31.665 4.060 ;
        RECT 32.045 3.525 32.185 4.645 ;
        RECT 33.375 4.315 33.515 4.775 ;
        RECT 32.825 3.685 33.105 4.155 ;
        RECT 33.315 4.055 33.575 4.315 ;
        RECT 33.305 3.685 33.585 4.055 ;
        RECT 32.045 3.475 32.355 3.525 ;
        RECT 33.855 3.515 33.995 4.835 ;
        RECT 34.235 4.315 34.375 5.305 ;
        RECT 34.545 4.555 34.805 4.875 ;
        RECT 36.405 4.835 36.665 5.155 ;
        RECT 34.175 3.995 34.435 4.315 ;
        RECT 34.605 3.515 34.745 4.555 ;
        RECT 36.465 4.055 36.605 4.835 ;
        RECT 37.670 4.265 38.010 4.345 ;
        RECT 35.715 3.945 35.975 4.035 ;
        RECT 35.055 3.805 35.975 3.945 ;
        RECT 33.515 3.495 33.995 3.515 ;
        RECT 28.785 3.155 29.045 3.475 ;
        RECT 31.515 3.385 31.775 3.475 ;
        RECT 31.985 3.445 32.355 3.475 ;
        RECT 31.515 3.155 31.835 3.385 ;
        RECT 31.695 3.005 31.835 3.155 ;
        RECT 31.985 3.150 32.395 3.445 ;
        RECT 32.585 3.155 32.865 3.495 ;
        RECT 33.315 3.245 33.995 3.495 ;
        RECT 34.535 3.445 34.815 3.515 ;
        RECT 33.315 3.145 33.795 3.245 ;
        RECT 34.485 3.185 34.860 3.445 ;
        RECT 34.535 3.145 34.815 3.185 ;
        RECT 35.055 3.005 35.195 3.805 ;
        RECT 35.715 3.715 35.975 3.805 ;
        RECT 36.295 3.685 36.605 4.055 ;
        RECT 36.365 3.500 36.605 3.685 ;
        RECT 37.045 4.065 38.010 4.265 ;
        RECT 36.365 3.435 36.675 3.500 ;
        RECT 37.045 3.435 37.245 4.065 ;
        RECT 37.670 3.995 38.010 4.065 ;
        RECT 37.760 3.990 37.930 3.995 ;
        RECT 38.960 3.860 39.120 9.035 ;
        RECT 40.075 8.945 40.400 9.035 ;
        RECT 42.455 9.180 42.805 9.300 ;
        RECT 49.895 9.180 50.245 9.255 ;
        RECT 55.335 9.205 55.660 9.270 ;
        RECT 42.455 8.980 50.245 9.180 ;
        RECT 42.455 8.950 42.805 8.980 ;
        RECT 49.895 8.905 50.245 8.980 ;
        RECT 54.220 9.035 55.660 9.205 ;
        RECT 39.275 8.510 39.595 8.835 ;
        RECT 39.305 8.335 39.475 8.510 ;
        RECT 39.305 8.160 39.480 8.335 ;
        RECT 39.305 7.985 40.280 8.160 ;
        RECT 39.275 3.860 39.595 3.980 ;
        RECT 38.960 3.690 39.595 3.860 ;
        RECT 39.275 3.660 39.595 3.690 ;
        RECT 40.105 3.610 40.280 7.985 ;
        RECT 47.195 5.305 49.635 5.445 ;
        RECT 47.195 5.155 47.335 5.305 ;
        RECT 46.895 5.065 47.335 5.155 ;
        RECT 44.555 4.925 47.335 5.065 ;
        RECT 44.045 4.785 44.305 4.875 ;
        RECT 44.555 4.785 44.695 4.925 ;
        RECT 46.895 4.835 47.155 4.925 ;
        RECT 47.495 4.835 47.755 5.155 ;
        RECT 47.495 4.785 47.695 4.835 ;
        RECT 44.045 4.645 44.695 4.785 ;
        RECT 47.305 4.645 47.695 4.785 ;
        RECT 48.565 4.775 48.845 5.155 ;
        RECT 49.055 4.835 49.330 5.155 ;
        RECT 44.045 4.555 44.305 4.645 ;
        RECT 36.365 3.245 37.245 3.435 ;
        RECT 40.050 3.260 40.400 3.610 ;
        RECT 44.105 3.475 44.245 4.555 ;
        RECT 44.965 4.505 45.245 4.620 ;
        RECT 46.415 4.505 46.675 4.595 ;
        RECT 44.795 4.365 46.675 4.505 ;
        RECT 44.795 4.315 45.245 4.365 ;
        RECT 44.735 4.245 45.245 4.315 ;
        RECT 46.415 4.275 46.675 4.365 ;
        RECT 44.735 4.055 44.995 4.245 ;
        RECT 45.910 4.055 46.215 4.060 ;
        RECT 44.725 3.685 45.005 4.055 ;
        RECT 45.215 3.945 45.475 4.035 ;
        RECT 45.805 3.945 46.215 4.055 ;
        RECT 45.215 3.805 46.215 3.945 ;
        RECT 45.215 3.715 45.475 3.805 ;
        RECT 45.805 3.685 46.215 3.805 ;
        RECT 46.645 3.685 46.925 4.060 ;
        RECT 47.305 3.525 47.445 4.645 ;
        RECT 48.635 4.315 48.775 4.775 ;
        RECT 48.085 3.685 48.365 4.155 ;
        RECT 48.575 4.055 48.835 4.315 ;
        RECT 48.565 3.685 48.845 4.055 ;
        RECT 47.305 3.475 47.615 3.525 ;
        RECT 49.115 3.515 49.255 4.835 ;
        RECT 49.495 4.315 49.635 5.305 ;
        RECT 49.805 4.555 50.065 4.875 ;
        RECT 51.665 4.835 51.925 5.155 ;
        RECT 49.435 3.995 49.695 4.315 ;
        RECT 49.865 3.515 50.005 4.555 ;
        RECT 51.725 4.055 51.865 4.835 ;
        RECT 52.930 4.265 53.270 4.345 ;
        RECT 50.975 3.945 51.235 4.035 ;
        RECT 50.315 3.805 51.235 3.945 ;
        RECT 48.775 3.495 49.255 3.515 ;
        RECT 36.395 3.235 37.245 3.245 ;
        RECT 36.395 3.125 36.675 3.235 ;
        RECT 44.045 3.155 44.305 3.475 ;
        RECT 46.775 3.385 47.035 3.475 ;
        RECT 47.245 3.445 47.615 3.475 ;
        RECT 46.775 3.155 47.095 3.385 ;
        RECT 31.695 2.865 35.195 3.005 ;
        RECT 46.955 3.005 47.095 3.155 ;
        RECT 47.245 3.150 47.655 3.445 ;
        RECT 47.845 3.155 48.125 3.495 ;
        RECT 48.575 3.245 49.255 3.495 ;
        RECT 49.795 3.445 50.075 3.515 ;
        RECT 48.575 3.145 49.055 3.245 ;
        RECT 49.745 3.185 50.120 3.445 ;
        RECT 49.795 3.145 50.075 3.185 ;
        RECT 50.315 3.005 50.455 3.805 ;
        RECT 50.975 3.715 51.235 3.805 ;
        RECT 51.555 3.685 51.865 4.055 ;
        RECT 51.625 3.500 51.865 3.685 ;
        RECT 52.305 4.065 53.270 4.265 ;
        RECT 51.625 3.435 51.935 3.500 ;
        RECT 52.305 3.435 52.505 4.065 ;
        RECT 52.930 3.995 53.270 4.065 ;
        RECT 53.020 3.990 53.190 3.995 ;
        RECT 54.220 3.860 54.380 9.035 ;
        RECT 55.335 8.945 55.660 9.035 ;
        RECT 57.715 9.180 58.065 9.300 ;
        RECT 65.155 9.180 65.505 9.255 ;
        RECT 70.595 9.205 70.920 9.270 ;
        RECT 57.715 8.980 65.505 9.180 ;
        RECT 57.715 8.950 58.065 8.980 ;
        RECT 65.155 8.905 65.505 8.980 ;
        RECT 69.480 9.035 70.920 9.205 ;
        RECT 54.535 8.510 54.855 8.835 ;
        RECT 54.565 8.335 54.735 8.510 ;
        RECT 54.565 8.160 54.740 8.335 ;
        RECT 54.565 7.985 55.540 8.160 ;
        RECT 54.535 3.860 54.855 3.980 ;
        RECT 54.220 3.690 54.855 3.860 ;
        RECT 54.535 3.660 54.855 3.690 ;
        RECT 55.365 3.610 55.540 7.985 ;
        RECT 62.455 5.305 64.895 5.445 ;
        RECT 62.455 5.155 62.595 5.305 ;
        RECT 62.155 5.065 62.595 5.155 ;
        RECT 59.815 4.925 62.595 5.065 ;
        RECT 59.305 4.785 59.565 4.875 ;
        RECT 59.815 4.785 59.955 4.925 ;
        RECT 62.155 4.835 62.415 4.925 ;
        RECT 62.755 4.835 63.015 5.155 ;
        RECT 62.755 4.785 62.955 4.835 ;
        RECT 59.305 4.645 59.955 4.785 ;
        RECT 62.565 4.645 62.955 4.785 ;
        RECT 63.825 4.775 64.105 5.155 ;
        RECT 64.315 4.835 64.590 5.155 ;
        RECT 59.305 4.555 59.565 4.645 ;
        RECT 51.625 3.245 52.505 3.435 ;
        RECT 55.310 3.260 55.660 3.610 ;
        RECT 59.365 3.475 59.505 4.555 ;
        RECT 60.225 4.505 60.505 4.620 ;
        RECT 61.675 4.505 61.935 4.595 ;
        RECT 60.055 4.365 61.935 4.505 ;
        RECT 60.055 4.315 60.505 4.365 ;
        RECT 59.995 4.245 60.505 4.315 ;
        RECT 61.675 4.275 61.935 4.365 ;
        RECT 59.995 4.055 60.255 4.245 ;
        RECT 61.170 4.055 61.475 4.060 ;
        RECT 59.985 3.685 60.265 4.055 ;
        RECT 60.475 3.945 60.735 4.035 ;
        RECT 61.065 3.945 61.475 4.055 ;
        RECT 60.475 3.805 61.475 3.945 ;
        RECT 60.475 3.715 60.735 3.805 ;
        RECT 61.065 3.685 61.475 3.805 ;
        RECT 61.905 3.685 62.185 4.060 ;
        RECT 62.565 3.525 62.705 4.645 ;
        RECT 63.895 4.315 64.035 4.775 ;
        RECT 63.345 3.685 63.625 4.155 ;
        RECT 63.835 4.055 64.095 4.315 ;
        RECT 63.825 3.685 64.105 4.055 ;
        RECT 62.565 3.475 62.875 3.525 ;
        RECT 64.375 3.515 64.515 4.835 ;
        RECT 64.755 4.315 64.895 5.305 ;
        RECT 65.065 4.555 65.325 4.875 ;
        RECT 66.925 4.835 67.185 5.155 ;
        RECT 64.695 3.995 64.955 4.315 ;
        RECT 65.125 3.515 65.265 4.555 ;
        RECT 66.985 4.055 67.125 4.835 ;
        RECT 68.190 4.265 68.530 4.345 ;
        RECT 66.235 3.945 66.495 4.035 ;
        RECT 65.575 3.805 66.495 3.945 ;
        RECT 64.035 3.495 64.515 3.515 ;
        RECT 51.655 3.235 52.505 3.245 ;
        RECT 51.655 3.125 51.935 3.235 ;
        RECT 59.305 3.155 59.565 3.475 ;
        RECT 62.035 3.385 62.295 3.475 ;
        RECT 62.505 3.445 62.875 3.475 ;
        RECT 62.035 3.155 62.355 3.385 ;
        RECT 46.955 2.865 50.455 3.005 ;
        RECT 62.215 3.005 62.355 3.155 ;
        RECT 62.505 3.150 62.915 3.445 ;
        RECT 63.105 3.155 63.385 3.495 ;
        RECT 63.835 3.245 64.515 3.495 ;
        RECT 65.055 3.445 65.335 3.515 ;
        RECT 63.835 3.145 64.315 3.245 ;
        RECT 65.005 3.185 65.380 3.445 ;
        RECT 65.055 3.145 65.335 3.185 ;
        RECT 65.575 3.005 65.715 3.805 ;
        RECT 66.235 3.715 66.495 3.805 ;
        RECT 66.815 3.685 67.125 4.055 ;
        RECT 66.885 3.500 67.125 3.685 ;
        RECT 67.565 4.065 68.530 4.265 ;
        RECT 66.885 3.435 67.195 3.500 ;
        RECT 67.565 3.435 67.765 4.065 ;
        RECT 68.190 3.995 68.530 4.065 ;
        RECT 68.280 3.990 68.450 3.995 ;
        RECT 69.480 3.860 69.640 9.035 ;
        RECT 70.595 8.945 70.920 9.035 ;
        RECT 72.930 9.180 73.280 9.300 ;
        RECT 80.420 9.180 80.770 9.255 ;
        RECT 85.855 9.205 86.180 9.270 ;
        RECT 72.930 8.980 80.770 9.180 ;
        RECT 72.930 8.950 73.280 8.980 ;
        RECT 80.420 8.905 80.770 8.980 ;
        RECT 84.740 9.035 86.180 9.205 ;
        RECT 69.795 8.510 70.115 8.835 ;
        RECT 69.825 8.335 69.995 8.510 ;
        RECT 69.825 8.160 70.000 8.335 ;
        RECT 69.825 7.985 70.800 8.160 ;
        RECT 69.795 3.860 70.115 3.980 ;
        RECT 69.480 3.690 70.115 3.860 ;
        RECT 69.795 3.660 70.115 3.690 ;
        RECT 70.625 3.610 70.800 7.985 ;
        RECT 77.715 5.305 80.155 5.445 ;
        RECT 77.715 5.155 77.855 5.305 ;
        RECT 77.415 5.065 77.855 5.155 ;
        RECT 75.075 4.925 77.855 5.065 ;
        RECT 74.565 4.785 74.825 4.875 ;
        RECT 75.075 4.785 75.215 4.925 ;
        RECT 77.415 4.835 77.675 4.925 ;
        RECT 78.015 4.835 78.275 5.155 ;
        RECT 78.015 4.785 78.215 4.835 ;
        RECT 74.565 4.645 75.215 4.785 ;
        RECT 77.825 4.645 78.215 4.785 ;
        RECT 79.085 4.775 79.365 5.155 ;
        RECT 79.575 4.835 79.850 5.155 ;
        RECT 74.565 4.555 74.825 4.645 ;
        RECT 66.885 3.245 67.765 3.435 ;
        RECT 70.570 3.260 70.920 3.610 ;
        RECT 74.625 3.475 74.765 4.555 ;
        RECT 75.485 4.505 75.765 4.620 ;
        RECT 76.935 4.505 77.195 4.595 ;
        RECT 75.315 4.365 77.195 4.505 ;
        RECT 75.315 4.315 75.765 4.365 ;
        RECT 75.255 4.245 75.765 4.315 ;
        RECT 76.935 4.275 77.195 4.365 ;
        RECT 75.255 4.055 75.515 4.245 ;
        RECT 76.430 4.055 76.735 4.060 ;
        RECT 75.245 3.685 75.525 4.055 ;
        RECT 75.735 3.945 75.995 4.035 ;
        RECT 76.325 3.945 76.735 4.055 ;
        RECT 75.735 3.805 76.735 3.945 ;
        RECT 75.735 3.715 75.995 3.805 ;
        RECT 76.325 3.685 76.735 3.805 ;
        RECT 77.165 3.685 77.445 4.060 ;
        RECT 77.825 3.525 77.965 4.645 ;
        RECT 79.155 4.315 79.295 4.775 ;
        RECT 78.605 3.685 78.885 4.155 ;
        RECT 79.095 4.055 79.355 4.315 ;
        RECT 79.085 3.685 79.365 4.055 ;
        RECT 77.825 3.475 78.135 3.525 ;
        RECT 79.635 3.515 79.775 4.835 ;
        RECT 80.015 4.315 80.155 5.305 ;
        RECT 80.325 4.555 80.585 4.875 ;
        RECT 82.185 4.835 82.445 5.155 ;
        RECT 79.955 3.995 80.215 4.315 ;
        RECT 80.385 3.515 80.525 4.555 ;
        RECT 82.245 4.055 82.385 4.835 ;
        RECT 83.450 4.265 83.790 4.345 ;
        RECT 81.495 3.945 81.755 4.035 ;
        RECT 80.835 3.805 81.755 3.945 ;
        RECT 79.295 3.495 79.775 3.515 ;
        RECT 66.915 3.235 67.765 3.245 ;
        RECT 66.915 3.125 67.195 3.235 ;
        RECT 74.565 3.155 74.825 3.475 ;
        RECT 77.295 3.385 77.555 3.475 ;
        RECT 77.765 3.445 78.135 3.475 ;
        RECT 77.295 3.155 77.615 3.385 ;
        RECT 62.215 2.865 65.715 3.005 ;
        RECT 77.475 3.005 77.615 3.155 ;
        RECT 77.765 3.150 78.175 3.445 ;
        RECT 78.365 3.155 78.645 3.495 ;
        RECT 79.095 3.245 79.775 3.495 ;
        RECT 80.315 3.445 80.595 3.515 ;
        RECT 79.095 3.145 79.575 3.245 ;
        RECT 80.265 3.185 80.640 3.445 ;
        RECT 80.315 3.145 80.595 3.185 ;
        RECT 80.835 3.005 80.975 3.805 ;
        RECT 81.495 3.715 81.755 3.805 ;
        RECT 82.075 3.685 82.385 4.055 ;
        RECT 82.145 3.500 82.385 3.685 ;
        RECT 82.825 4.065 83.790 4.265 ;
        RECT 82.145 3.435 82.455 3.500 ;
        RECT 82.825 3.435 83.025 4.065 ;
        RECT 83.450 3.995 83.790 4.065 ;
        RECT 83.540 3.990 83.710 3.995 ;
        RECT 84.740 3.860 84.900 9.035 ;
        RECT 85.855 8.945 86.180 9.035 ;
        RECT 88.190 9.180 88.540 9.300 ;
        RECT 95.675 9.180 96.025 9.255 ;
        RECT 101.115 9.205 101.440 9.270 ;
        RECT 88.190 8.980 96.025 9.180 ;
        RECT 88.190 8.950 88.540 8.980 ;
        RECT 95.675 8.905 96.025 8.980 ;
        RECT 100.000 9.035 101.440 9.205 ;
        RECT 85.055 8.510 85.375 8.835 ;
        RECT 85.085 8.335 85.255 8.510 ;
        RECT 85.085 8.160 85.260 8.335 ;
        RECT 85.085 7.985 86.060 8.160 ;
        RECT 85.055 3.860 85.375 3.980 ;
        RECT 84.740 3.690 85.375 3.860 ;
        RECT 85.055 3.660 85.375 3.690 ;
        RECT 85.885 3.610 86.060 7.985 ;
        RECT 92.975 5.305 95.415 5.445 ;
        RECT 92.975 5.155 93.115 5.305 ;
        RECT 92.675 5.065 93.115 5.155 ;
        RECT 90.335 4.925 93.115 5.065 ;
        RECT 89.825 4.785 90.085 4.875 ;
        RECT 90.335 4.785 90.475 4.925 ;
        RECT 92.675 4.835 92.935 4.925 ;
        RECT 93.275 4.835 93.535 5.155 ;
        RECT 93.275 4.785 93.475 4.835 ;
        RECT 89.825 4.645 90.475 4.785 ;
        RECT 93.085 4.645 93.475 4.785 ;
        RECT 94.345 4.775 94.625 5.155 ;
        RECT 94.835 4.835 95.110 5.155 ;
        RECT 89.825 4.555 90.085 4.645 ;
        RECT 82.145 3.245 83.025 3.435 ;
        RECT 85.830 3.260 86.180 3.610 ;
        RECT 89.885 3.475 90.025 4.555 ;
        RECT 90.745 4.505 91.025 4.620 ;
        RECT 92.195 4.505 92.455 4.595 ;
        RECT 90.575 4.365 92.455 4.505 ;
        RECT 90.575 4.315 91.025 4.365 ;
        RECT 90.515 4.245 91.025 4.315 ;
        RECT 92.195 4.275 92.455 4.365 ;
        RECT 90.515 4.055 90.775 4.245 ;
        RECT 91.690 4.055 91.995 4.060 ;
        RECT 90.505 3.685 90.785 4.055 ;
        RECT 90.995 3.945 91.255 4.035 ;
        RECT 91.585 3.945 91.995 4.055 ;
        RECT 90.995 3.805 91.995 3.945 ;
        RECT 90.995 3.715 91.255 3.805 ;
        RECT 91.585 3.685 91.995 3.805 ;
        RECT 92.425 3.685 92.705 4.060 ;
        RECT 93.085 3.525 93.225 4.645 ;
        RECT 94.415 4.315 94.555 4.775 ;
        RECT 93.865 3.685 94.145 4.155 ;
        RECT 94.355 4.055 94.615 4.315 ;
        RECT 94.345 3.685 94.625 4.055 ;
        RECT 93.085 3.475 93.395 3.525 ;
        RECT 94.895 3.515 95.035 4.835 ;
        RECT 95.275 4.315 95.415 5.305 ;
        RECT 95.585 4.555 95.845 4.875 ;
        RECT 97.445 4.835 97.705 5.155 ;
        RECT 95.215 3.995 95.475 4.315 ;
        RECT 95.645 3.515 95.785 4.555 ;
        RECT 97.505 4.055 97.645 4.835 ;
        RECT 98.710 4.265 99.050 4.345 ;
        RECT 96.755 3.945 97.015 4.035 ;
        RECT 96.095 3.805 97.015 3.945 ;
        RECT 94.555 3.495 95.035 3.515 ;
        RECT 82.175 3.235 83.025 3.245 ;
        RECT 82.175 3.125 82.455 3.235 ;
        RECT 89.825 3.155 90.085 3.475 ;
        RECT 92.555 3.385 92.815 3.475 ;
        RECT 93.025 3.445 93.395 3.475 ;
        RECT 92.555 3.155 92.875 3.385 ;
        RECT 77.475 2.865 80.975 3.005 ;
        RECT 92.735 3.005 92.875 3.155 ;
        RECT 93.025 3.150 93.435 3.445 ;
        RECT 93.625 3.155 93.905 3.495 ;
        RECT 94.355 3.245 95.035 3.495 ;
        RECT 95.575 3.445 95.855 3.515 ;
        RECT 94.355 3.145 94.835 3.245 ;
        RECT 95.525 3.185 95.900 3.445 ;
        RECT 95.575 3.145 95.855 3.185 ;
        RECT 96.095 3.005 96.235 3.805 ;
        RECT 96.755 3.715 97.015 3.805 ;
        RECT 97.335 3.685 97.645 4.055 ;
        RECT 97.405 3.500 97.645 3.685 ;
        RECT 98.085 4.065 99.050 4.265 ;
        RECT 97.405 3.435 97.715 3.500 ;
        RECT 98.085 3.435 98.285 4.065 ;
        RECT 98.710 3.995 99.050 4.065 ;
        RECT 98.800 3.990 98.970 3.995 ;
        RECT 100.000 3.860 100.160 9.035 ;
        RECT 101.115 8.945 101.440 9.035 ;
        RECT 100.315 8.510 100.635 8.835 ;
        RECT 100.345 8.335 100.515 8.510 ;
        RECT 100.345 8.160 100.520 8.335 ;
        RECT 100.345 7.985 101.320 8.160 ;
        RECT 100.315 3.860 100.635 3.980 ;
        RECT 100.000 3.690 100.635 3.860 ;
        RECT 100.315 3.660 100.635 3.690 ;
        RECT 101.145 3.610 101.320 7.985 ;
        RECT 97.405 3.245 98.285 3.435 ;
        RECT 101.090 3.260 101.440 3.610 ;
        RECT 97.435 3.235 98.285 3.245 ;
        RECT 97.435 3.125 97.715 3.235 ;
        RECT 92.735 2.865 96.235 3.005 ;
      LAYER met3 ;
        RECT 33.965 9.345 34.335 9.715 ;
        RECT 49.225 9.345 49.595 9.715 ;
        RECT 64.485 9.345 64.855 9.715 ;
        RECT 79.745 9.345 80.115 9.715 ;
        RECT 95.005 9.345 95.375 9.715 ;
        RECT 34.000 6.530 34.300 9.345 ;
        RECT 49.260 6.530 49.560 9.345 ;
        RECT 64.520 6.530 64.820 9.345 ;
        RECT 79.780 6.530 80.080 9.345 ;
        RECT 95.040 6.530 95.340 9.345 ;
        RECT 33.995 6.175 34.300 6.530 ;
        RECT 49.255 6.175 49.560 6.530 ;
        RECT 64.515 6.175 64.820 6.530 ;
        RECT 79.775 6.175 80.080 6.530 ;
        RECT 95.035 6.175 95.340 6.530 ;
        RECT 33.995 5.770 34.295 6.175 ;
        RECT 49.255 5.770 49.555 6.175 ;
        RECT 64.515 5.770 64.815 6.175 ;
        RECT 79.775 5.770 80.075 6.175 ;
        RECT 95.035 5.770 95.335 6.175 ;
        RECT 29.765 5.470 34.295 5.770 ;
        RECT 45.025 5.470 49.555 5.770 ;
        RECT 60.285 5.470 64.815 5.770 ;
        RECT 75.545 5.470 80.075 5.770 ;
        RECT 90.805 5.470 95.335 5.770 ;
        RECT 29.765 4.600 30.065 5.470 ;
        RECT 32.560 5.145 32.860 5.470 ;
        RECT 33.285 5.145 33.615 5.155 ;
        RECT 31.375 4.845 33.615 5.145 ;
        RECT 29.685 4.595 30.065 4.600 ;
        RECT 29.455 4.265 30.185 4.595 ;
        RECT 30.645 4.245 30.965 4.625 ;
        RECT 30.645 4.055 30.975 4.245 ;
        RECT 31.375 4.055 31.675 4.845 ;
        RECT 32.560 4.155 32.860 4.845 ;
        RECT 33.275 4.795 33.615 4.845 ;
        RECT 45.025 4.600 45.325 5.470 ;
        RECT 47.820 5.145 48.120 5.470 ;
        RECT 48.545 5.145 48.875 5.155 ;
        RECT 46.635 4.845 48.875 5.145 ;
        RECT 44.945 4.595 45.325 4.600 ;
        RECT 44.715 4.265 45.445 4.595 ;
        RECT 45.905 4.245 46.225 4.625 ;
        RECT 30.645 3.705 30.980 4.055 ;
        RECT 31.355 4.040 31.675 4.055 ;
        RECT 31.355 3.705 31.695 4.040 ;
        RECT 32.355 3.815 33.135 4.155 ;
        RECT 32.560 3.810 33.135 3.815 ;
        RECT 32.795 3.805 33.135 3.810 ;
        RECT 32.805 3.775 33.135 3.805 ;
        RECT 45.905 4.055 46.235 4.245 ;
        RECT 46.635 4.055 46.935 4.845 ;
        RECT 47.820 4.155 48.120 4.845 ;
        RECT 48.535 4.795 48.875 4.845 ;
        RECT 60.285 4.600 60.585 5.470 ;
        RECT 63.080 5.145 63.380 5.470 ;
        RECT 63.805 5.145 64.135 5.155 ;
        RECT 61.895 4.845 64.135 5.145 ;
        RECT 60.205 4.595 60.585 4.600 ;
        RECT 59.975 4.265 60.705 4.595 ;
        RECT 61.165 4.245 61.485 4.625 ;
        RECT 45.905 3.705 46.240 4.055 ;
        RECT 46.615 4.040 46.935 4.055 ;
        RECT 46.615 3.705 46.955 4.040 ;
        RECT 47.615 3.815 48.395 4.155 ;
        RECT 47.820 3.810 48.395 3.815 ;
        RECT 48.055 3.805 48.395 3.810 ;
        RECT 48.065 3.775 48.395 3.805 ;
        RECT 61.165 4.055 61.495 4.245 ;
        RECT 61.895 4.055 62.195 4.845 ;
        RECT 63.080 4.155 63.380 4.845 ;
        RECT 63.795 4.795 64.135 4.845 ;
        RECT 75.545 4.600 75.845 5.470 ;
        RECT 78.340 5.145 78.640 5.470 ;
        RECT 79.065 5.145 79.395 5.155 ;
        RECT 77.155 4.845 79.395 5.145 ;
        RECT 75.465 4.595 75.845 4.600 ;
        RECT 75.235 4.265 75.965 4.595 ;
        RECT 76.425 4.245 76.745 4.625 ;
        RECT 61.165 3.705 61.500 4.055 ;
        RECT 61.875 4.040 62.195 4.055 ;
        RECT 61.875 3.705 62.215 4.040 ;
        RECT 62.875 3.815 63.655 4.155 ;
        RECT 63.080 3.810 63.655 3.815 ;
        RECT 63.315 3.805 63.655 3.810 ;
        RECT 63.325 3.775 63.655 3.805 ;
        RECT 76.425 4.055 76.755 4.245 ;
        RECT 77.155 4.055 77.455 4.845 ;
        RECT 78.340 4.155 78.640 4.845 ;
        RECT 79.055 4.795 79.395 4.845 ;
        RECT 90.805 4.600 91.105 5.470 ;
        RECT 93.600 5.145 93.900 5.470 ;
        RECT 94.325 5.145 94.655 5.155 ;
        RECT 92.415 4.845 94.655 5.145 ;
        RECT 90.725 4.595 91.105 4.600 ;
        RECT 90.495 4.265 91.225 4.595 ;
        RECT 91.685 4.245 92.005 4.625 ;
        RECT 76.425 3.705 76.760 4.055 ;
        RECT 77.135 4.040 77.455 4.055 ;
        RECT 77.135 3.705 77.475 4.040 ;
        RECT 78.135 3.815 78.915 4.155 ;
        RECT 78.340 3.810 78.915 3.815 ;
        RECT 78.575 3.805 78.915 3.810 ;
        RECT 78.585 3.775 78.915 3.805 ;
        RECT 91.685 4.055 92.015 4.245 ;
        RECT 92.415 4.055 92.715 4.845 ;
        RECT 93.600 4.155 93.900 4.845 ;
        RECT 94.315 4.795 94.655 4.845 ;
        RECT 91.685 3.705 92.020 4.055 ;
        RECT 92.395 4.040 92.715 4.055 ;
        RECT 92.395 3.705 92.735 4.040 ;
        RECT 93.395 3.815 94.175 4.155 ;
        RECT 93.600 3.810 94.175 3.815 ;
        RECT 93.835 3.805 94.175 3.810 ;
        RECT 93.845 3.775 94.175 3.805 ;
        RECT 31.925 3.175 32.655 3.505 ;
        RECT 33.470 3.495 33.820 3.500 ;
        RECT 31.925 3.165 32.405 3.175 ;
        RECT 33.470 3.145 34.205 3.495 ;
        RECT 34.505 3.165 35.245 3.495 ;
        RECT 36.365 3.475 36.725 3.480 ;
        RECT 34.505 3.155 34.835 3.165 ;
        RECT 36.205 3.145 36.935 3.475 ;
        RECT 47.185 3.175 47.915 3.505 ;
        RECT 48.730 3.495 49.080 3.500 ;
        RECT 47.185 3.165 47.665 3.175 ;
        RECT 48.730 3.145 49.465 3.495 ;
        RECT 49.765 3.165 50.505 3.495 ;
        RECT 51.625 3.475 51.985 3.480 ;
        RECT 49.765 3.155 50.095 3.165 ;
        RECT 51.465 3.145 52.195 3.475 ;
        RECT 62.445 3.175 63.175 3.505 ;
        RECT 63.990 3.495 64.340 3.500 ;
        RECT 62.445 3.165 62.925 3.175 ;
        RECT 63.990 3.145 64.725 3.495 ;
        RECT 65.025 3.165 65.765 3.495 ;
        RECT 66.885 3.475 67.245 3.480 ;
        RECT 65.025 3.155 65.355 3.165 ;
        RECT 66.725 3.145 67.455 3.475 ;
        RECT 77.705 3.175 78.435 3.505 ;
        RECT 79.250 3.495 79.600 3.500 ;
        RECT 77.705 3.165 78.185 3.175 ;
        RECT 79.250 3.145 79.985 3.495 ;
        RECT 80.285 3.165 81.025 3.495 ;
        RECT 82.145 3.475 82.505 3.480 ;
        RECT 80.285 3.155 80.615 3.165 ;
        RECT 81.985 3.145 82.715 3.475 ;
        RECT 92.965 3.175 93.695 3.505 ;
        RECT 94.510 3.495 94.860 3.500 ;
        RECT 92.965 3.165 93.445 3.175 ;
        RECT 94.510 3.145 95.245 3.495 ;
        RECT 95.545 3.165 96.285 3.495 ;
        RECT 97.405 3.475 97.765 3.480 ;
        RECT 95.545 3.155 95.875 3.165 ;
        RECT 97.245 3.145 97.975 3.475 ;
        RECT 33.470 3.140 33.820 3.145 ;
        RECT 36.365 3.140 36.725 3.145 ;
        RECT 48.730 3.140 49.080 3.145 ;
        RECT 51.625 3.140 51.985 3.145 ;
        RECT 63.990 3.140 64.340 3.145 ;
        RECT 66.885 3.140 67.245 3.145 ;
        RECT 79.250 3.140 79.600 3.145 ;
        RECT 82.145 3.140 82.505 3.145 ;
        RECT 94.510 3.140 94.860 3.145 ;
        RECT 97.405 3.140 97.765 3.145 ;
      LAYER met4 ;
        RECT 30.635 4.265 30.975 4.600 ;
        RECT 45.895 4.265 46.235 4.600 ;
        RECT 61.155 4.265 61.495 4.600 ;
        RECT 76.415 4.265 76.755 4.600 ;
        RECT 91.675 4.265 92.015 4.600 ;
        RECT 30.655 4.095 30.975 4.265 ;
        RECT 32.795 4.095 33.135 4.135 ;
        RECT 30.655 3.795 33.135 4.095 ;
        RECT 45.915 4.095 46.235 4.265 ;
        RECT 48.055 4.095 48.395 4.135 ;
        RECT 45.915 3.795 48.395 4.095 ;
        RECT 61.175 4.095 61.495 4.265 ;
        RECT 63.315 4.095 63.655 4.135 ;
        RECT 61.175 3.795 63.655 4.095 ;
        RECT 76.435 4.095 76.755 4.265 ;
        RECT 78.575 4.095 78.915 4.135 ;
        RECT 76.435 3.795 78.915 4.095 ;
        RECT 91.695 4.095 92.015 4.265 ;
        RECT 93.835 4.095 94.175 4.135 ;
        RECT 91.695 3.795 94.175 4.095 ;
        RECT 32.805 3.775 33.135 3.795 ;
        RECT 48.065 3.775 48.395 3.795 ;
        RECT 63.325 3.775 63.655 3.795 ;
        RECT 78.585 3.775 78.915 3.795 ;
        RECT 93.845 3.775 94.175 3.795 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r1
MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r2
  CLASS BLOCK ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ct_8_b0r2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 103.915 BY 12.465 ;
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 18.635 8.235 18.805 9.505 ;
        RECT 30.320 8.465 30.490 9.505 ;
        RECT 30.315 8.225 30.495 8.465 ;
        RECT 30.320 2.955 30.490 4.225 ;
      LAYER met1 ;
        RECT 18.545 8.405 18.885 8.490 ;
        RECT 18.545 8.375 19.035 8.405 ;
        RECT 20.860 8.375 21.200 8.455 ;
        RECT 18.545 8.200 21.200 8.375 ;
        RECT 18.545 8.150 18.885 8.200 ;
        RECT 20.860 8.175 21.200 8.200 ;
        RECT 30.245 8.405 30.570 8.465 ;
        RECT 30.245 8.235 30.720 8.405 ;
        RECT 30.245 8.140 30.570 8.235 ;
        RECT 30.245 4.790 30.570 5.115 ;
        RECT 30.325 4.255 30.495 4.790 ;
        RECT 30.260 4.225 30.550 4.255 ;
        RECT 30.260 4.055 30.720 4.225 ;
        RECT 30.260 4.025 30.550 4.055 ;
      LAYER met2 ;
        RECT 20.945 9.240 30.495 9.410 ;
        RECT 18.525 8.135 18.900 8.505 ;
        RECT 20.945 8.485 21.115 9.240 ;
        RECT 20.890 8.145 21.170 8.485 ;
        RECT 30.325 8.465 30.495 9.240 ;
        RECT 30.245 8.140 30.570 8.465 ;
        RECT 30.315 5.115 30.485 8.140 ;
        RECT 30.245 4.790 30.570 5.115 ;
      LAYER met3 ;
        RECT 18.545 8.505 18.880 12.385 ;
        RECT 18.525 8.135 18.900 8.505 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 35.855 8.235 36.025 9.505 ;
        RECT 47.540 8.465 47.710 9.505 ;
        RECT 47.535 8.225 47.715 8.465 ;
        RECT 47.540 2.955 47.710 4.225 ;
      LAYER met1 ;
        RECT 35.765 8.405 36.105 8.490 ;
        RECT 35.765 8.375 36.255 8.405 ;
        RECT 38.080 8.375 38.420 8.455 ;
        RECT 35.765 8.200 38.420 8.375 ;
        RECT 35.765 8.150 36.105 8.200 ;
        RECT 38.080 8.175 38.420 8.200 ;
        RECT 47.465 8.405 47.790 8.465 ;
        RECT 47.465 8.235 47.940 8.405 ;
        RECT 47.465 8.140 47.790 8.235 ;
        RECT 47.465 4.790 47.790 5.115 ;
        RECT 47.545 4.255 47.715 4.790 ;
        RECT 47.480 4.225 47.770 4.255 ;
        RECT 47.480 4.055 47.940 4.225 ;
        RECT 47.480 4.025 47.770 4.055 ;
      LAYER met2 ;
        RECT 38.165 9.240 47.715 9.410 ;
        RECT 35.745 8.135 36.120 8.505 ;
        RECT 38.165 8.485 38.335 9.240 ;
        RECT 38.110 8.145 38.390 8.485 ;
        RECT 47.545 8.465 47.715 9.240 ;
        RECT 47.465 8.140 47.790 8.465 ;
        RECT 47.535 5.115 47.705 8.140 ;
        RECT 47.465 4.790 47.790 5.115 ;
      LAYER met3 ;
        RECT 35.765 8.505 36.100 12.385 ;
        RECT 35.745 8.135 36.120 8.505 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 53.075 8.240 53.245 9.510 ;
        RECT 64.760 8.470 64.930 9.510 ;
        RECT 64.755 8.230 64.935 8.470 ;
        RECT 64.760 2.960 64.930 4.230 ;
      LAYER met1 ;
        RECT 52.985 8.410 53.325 8.495 ;
        RECT 52.985 8.380 53.475 8.410 ;
        RECT 55.300 8.380 55.640 8.460 ;
        RECT 52.985 8.205 55.640 8.380 ;
        RECT 52.985 8.155 53.325 8.205 ;
        RECT 55.300 8.180 55.640 8.205 ;
        RECT 64.685 8.410 65.010 8.470 ;
        RECT 64.685 8.240 65.160 8.410 ;
        RECT 64.685 8.145 65.010 8.240 ;
        RECT 64.685 4.795 65.010 5.120 ;
        RECT 64.765 4.260 64.935 4.795 ;
        RECT 64.700 4.230 64.990 4.260 ;
        RECT 64.700 4.060 65.160 4.230 ;
        RECT 64.700 4.030 64.990 4.060 ;
      LAYER met2 ;
        RECT 55.385 9.245 64.935 9.415 ;
        RECT 52.965 8.140 53.340 8.510 ;
        RECT 55.385 8.490 55.555 9.245 ;
        RECT 55.330 8.150 55.610 8.490 ;
        RECT 64.765 8.470 64.935 9.245 ;
        RECT 64.685 8.145 65.010 8.470 ;
        RECT 64.755 5.120 64.925 8.145 ;
        RECT 64.685 4.795 65.010 5.120 ;
      LAYER met3 ;
        RECT 52.985 8.510 53.320 12.390 ;
        RECT 52.965 8.140 53.340 8.510 ;
    END
  END s3
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 103.350 4.010 103.525 5.155 ;
        RECT 103.350 3.575 103.520 4.010 ;
        RECT 103.355 1.865 103.525 2.375 ;
      LAYER met1 ;
        RECT 103.290 3.540 103.580 3.775 ;
        RECT 103.290 3.535 103.520 3.540 ;
        RECT 103.350 2.435 103.520 3.535 ;
        RECT 103.290 2.175 103.585 2.435 ;
    END
  END X5_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 68.910 4.015 69.085 5.160 ;
        RECT 68.910 3.580 69.080 4.015 ;
        RECT 68.915 1.870 69.085 2.380 ;
      LAYER met1 ;
        RECT 68.850 3.545 69.140 3.780 ;
        RECT 68.850 3.540 69.080 3.545 ;
        RECT 68.910 2.440 69.080 3.540 ;
        RECT 68.850 2.180 69.145 2.440 ;
    END
  END X3_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 51.690 4.010 51.865 5.155 ;
        RECT 51.690 3.575 51.860 4.010 ;
        RECT 51.695 1.865 51.865 2.375 ;
      LAYER met1 ;
        RECT 51.630 3.540 51.920 3.775 ;
        RECT 51.630 3.535 51.860 3.540 ;
        RECT 51.690 2.435 51.860 3.535 ;
        RECT 51.630 2.175 51.925 2.435 ;
    END
  END X2_Y1
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 34.470 4.010 34.645 5.155 ;
        RECT 34.470 3.575 34.640 4.010 ;
        RECT 34.475 1.865 34.645 2.375 ;
      LAYER met1 ;
        RECT 34.410 3.540 34.700 3.775 ;
        RECT 34.410 3.535 34.640 3.540 ;
        RECT 34.470 2.435 34.640 3.535 ;
        RECT 34.410 2.175 34.705 2.435 ;
    END
  END X1_Y1
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 87.515 8.235 87.685 9.505 ;
        RECT 99.200 8.465 99.370 9.505 ;
        RECT 99.195 8.225 99.375 8.465 ;
        RECT 99.200 2.955 99.370 4.225 ;
      LAYER met1 ;
        RECT 87.425 8.405 87.765 8.490 ;
        RECT 87.425 8.375 87.915 8.405 ;
        RECT 89.740 8.375 90.080 8.455 ;
        RECT 87.425 8.200 90.080 8.375 ;
        RECT 87.425 8.150 87.765 8.200 ;
        RECT 89.740 8.175 90.080 8.200 ;
        RECT 99.125 8.405 99.450 8.465 ;
        RECT 99.125 8.235 99.600 8.405 ;
        RECT 99.125 8.140 99.450 8.235 ;
        RECT 99.125 4.790 99.450 5.115 ;
        RECT 99.205 4.255 99.375 4.790 ;
        RECT 99.140 4.225 99.430 4.255 ;
        RECT 99.140 4.055 99.600 4.225 ;
        RECT 99.140 4.025 99.430 4.055 ;
      LAYER met2 ;
        RECT 89.825 9.240 99.375 9.410 ;
        RECT 87.405 8.135 87.780 8.505 ;
        RECT 89.825 8.485 89.995 9.240 ;
        RECT 89.770 8.145 90.050 8.485 ;
        RECT 99.205 8.465 99.375 9.240 ;
        RECT 99.125 8.140 99.450 8.465 ;
        RECT 99.195 5.115 99.365 8.140 ;
        RECT 99.125 4.790 99.450 5.115 ;
      LAYER met3 ;
        RECT 87.425 8.505 87.760 12.385 ;
        RECT 87.405 8.135 87.780 8.505 ;
    END
  END s5
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 70.295 8.235 70.465 9.505 ;
        RECT 81.980 8.465 82.150 9.505 ;
        RECT 81.975 8.225 82.155 8.465 ;
        RECT 81.980 2.955 82.150 4.225 ;
      LAYER met1 ;
        RECT 70.205 8.405 70.545 8.490 ;
        RECT 70.205 8.375 70.695 8.405 ;
        RECT 72.520 8.375 72.860 8.455 ;
        RECT 70.205 8.200 72.860 8.375 ;
        RECT 70.205 8.150 70.545 8.200 ;
        RECT 72.520 8.175 72.860 8.200 ;
        RECT 81.905 8.405 82.230 8.465 ;
        RECT 81.905 8.235 82.380 8.405 ;
        RECT 81.905 8.140 82.230 8.235 ;
        RECT 81.905 4.790 82.230 5.115 ;
        RECT 81.985 4.255 82.155 4.790 ;
        RECT 81.920 4.225 82.210 4.255 ;
        RECT 81.920 4.055 82.380 4.225 ;
        RECT 81.920 4.025 82.210 4.055 ;
      LAYER met2 ;
        RECT 72.605 9.240 82.155 9.410 ;
        RECT 70.185 8.135 70.560 8.505 ;
        RECT 72.605 8.485 72.775 9.240 ;
        RECT 72.550 8.145 72.830 8.485 ;
        RECT 81.985 8.465 82.155 9.240 ;
        RECT 81.905 8.140 82.230 8.465 ;
        RECT 81.975 5.115 82.145 8.140 ;
        RECT 81.905 4.790 82.230 5.115 ;
      LAYER met3 ;
        RECT 70.205 8.505 70.540 12.385 ;
        RECT 70.185 8.135 70.560 8.505 ;
    END
  END s4
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 15.225 8.235 15.395 9.505 ;
      LAYER met1 ;
        RECT 15.165 8.430 15.455 8.435 ;
        RECT 15.165 8.405 15.460 8.430 ;
        RECT 15.165 8.235 15.625 8.405 ;
        RECT 15.165 8.205 15.460 8.235 ;
        RECT 15.170 8.200 15.460 8.205 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 52.845 8.745 55.655 8.750 ;
        RECT 64.530 8.745 69.310 8.750 ;
        RECT 14.995 8.740 21.215 8.745 ;
        RECT 30.090 8.740 38.435 8.745 ;
        RECT 47.310 8.740 55.800 8.745 ;
        RECT 14.995 7.140 21.385 8.740 ;
        RECT 29.325 8.130 38.580 8.740 ;
        RECT 46.545 8.130 55.800 8.740 ;
        RECT 63.765 8.740 72.875 8.745 ;
        RECT 81.750 8.740 90.095 8.745 ;
        RECT 98.970 8.740 103.750 8.745 ;
        RECT 63.765 8.135 73.020 8.740 ;
        RECT 29.130 7.140 38.580 8.130 ;
        RECT 46.350 7.145 55.800 8.130 ;
        RECT 63.570 7.145 73.020 8.135 ;
        RECT 80.985 8.130 90.240 8.740 ;
        RECT 98.205 8.130 103.900 8.740 ;
        RECT 46.350 7.140 73.020 7.145 ;
        RECT 80.790 7.140 90.240 8.130 ;
        RECT 98.010 7.140 103.900 8.130 ;
        RECT 14.995 6.655 103.900 7.140 ;
        RECT 15.000 4.775 103.900 6.655 ;
        RECT 14.995 4.315 103.900 4.775 ;
        RECT 14.995 4.310 55.825 4.315 ;
        RECT 14.995 3.710 21.385 4.310 ;
        RECT 29.325 3.720 38.605 4.310 ;
        RECT 46.545 3.720 55.825 4.310 ;
        RECT 63.765 4.310 103.900 4.315 ;
        RECT 63.765 3.725 73.045 4.310 ;
        RECT 64.530 3.720 73.045 3.725 ;
        RECT 80.985 3.720 90.265 4.310 ;
        RECT 98.205 3.720 103.900 4.310 ;
        RECT 30.090 3.715 38.605 3.720 ;
        RECT 47.310 3.715 55.825 3.720 ;
        RECT 35.010 3.710 38.605 3.715 ;
        RECT 69.300 3.710 73.045 3.720 ;
        RECT 81.750 3.715 90.265 3.720 ;
        RECT 98.970 3.715 103.745 3.720 ;
        RECT 86.525 3.710 90.265 3.715 ;
      LAYER li1 ;
        RECT 17.030 10.045 17.205 10.595 ;
        RECT 17.030 8.445 17.200 10.045 ;
        RECT 15.215 7.035 15.385 7.765 ;
        RECT 17.030 7.305 17.205 8.445 ;
        RECT 17.030 7.035 17.200 7.305 ;
        RECT 18.625 7.035 18.795 7.765 ;
        RECT 30.310 7.035 30.480 7.765 ;
        RECT 33.055 7.035 33.225 7.765 ;
        RECT 34.045 7.035 34.215 7.765 ;
        RECT 35.845 7.035 36.015 7.765 ;
        RECT 47.530 7.035 47.700 7.765 ;
        RECT 50.275 7.035 50.445 7.765 ;
        RECT 51.265 7.035 51.435 7.765 ;
        RECT 53.065 7.040 53.235 7.770 ;
        RECT 64.750 7.040 64.920 7.770 ;
        RECT 67.495 7.040 67.665 7.770 ;
        RECT 68.485 7.040 68.655 7.770 ;
        RECT 15.045 7.025 17.795 7.035 ;
        RECT 18.455 7.025 21.205 7.035 ;
        RECT 30.140 7.030 34.865 7.035 ;
        RECT 35.675 7.030 38.425 7.035 ;
        RECT 47.360 7.030 52.085 7.035 ;
        RECT 52.895 7.030 55.645 7.040 ;
        RECT 64.580 7.035 69.305 7.040 ;
        RECT 70.285 7.035 70.455 7.765 ;
        RECT 81.970 7.035 82.140 7.765 ;
        RECT 84.715 7.035 84.885 7.765 ;
        RECT 85.705 7.035 85.875 7.765 ;
        RECT 87.505 7.035 87.675 7.765 ;
        RECT 99.190 7.035 99.360 7.765 ;
        RECT 101.935 7.035 102.105 7.765 ;
        RECT 102.925 7.035 103.095 7.765 ;
        RECT 63.475 7.030 69.460 7.035 ;
        RECT 70.115 7.030 72.865 7.035 ;
        RECT 81.800 7.030 86.525 7.035 ;
        RECT 87.335 7.030 90.085 7.035 ;
        RECT 99.020 7.030 103.745 7.035 ;
        RECT 0.000 7.000 21.470 7.025 ;
        RECT 29.035 7.005 38.580 7.030 ;
        RECT 0.000 6.800 21.940 7.000 ;
        RECT 0.000 5.810 21.945 6.800 ;
        RECT 22.130 5.810 22.410 6.950 ;
        RECT 23.080 5.810 23.340 6.950 ;
        RECT 24.430 5.810 24.710 6.950 ;
        RECT 25.380 5.810 25.640 6.950 ;
        RECT 25.810 5.810 26.070 6.950 ;
        RECT 26.740 5.810 27.020 6.950 ;
        RECT 27.190 5.810 27.450 6.950 ;
        RECT 28.120 5.810 28.400 6.950 ;
        RECT 29.035 6.800 38.585 7.005 ;
        RECT 28.935 5.810 39.165 6.800 ;
        RECT 39.350 5.810 39.630 6.950 ;
        RECT 40.300 5.810 40.560 6.950 ;
        RECT 41.650 5.810 41.930 6.950 ;
        RECT 42.600 5.810 42.860 6.950 ;
        RECT 43.030 5.810 43.290 6.950 ;
        RECT 43.960 5.810 44.240 6.950 ;
        RECT 44.410 5.810 44.670 6.950 ;
        RECT 45.340 5.810 45.620 6.950 ;
        RECT 46.255 6.805 55.805 7.030 ;
        RECT 46.255 6.800 56.385 6.805 ;
        RECT 46.155 5.815 56.385 6.800 ;
        RECT 56.570 5.815 56.850 6.955 ;
        RECT 57.520 5.815 57.780 6.955 ;
        RECT 58.870 5.815 59.150 6.955 ;
        RECT 59.820 5.815 60.080 6.955 ;
        RECT 60.250 5.815 60.510 6.955 ;
        RECT 61.180 5.815 61.460 6.955 ;
        RECT 61.630 5.815 61.890 6.955 ;
        RECT 62.560 5.815 62.840 6.955 ;
        RECT 63.475 6.805 73.025 7.030 ;
        RECT 63.375 6.800 73.025 6.805 ;
        RECT 63.375 5.815 73.605 6.800 ;
        RECT 46.155 5.810 73.605 5.815 ;
        RECT 73.790 5.810 74.070 6.950 ;
        RECT 74.740 5.810 75.000 6.950 ;
        RECT 76.090 5.810 76.370 6.950 ;
        RECT 77.040 5.810 77.300 6.950 ;
        RECT 77.470 5.810 77.730 6.950 ;
        RECT 78.400 5.810 78.680 6.950 ;
        RECT 78.850 5.810 79.110 6.950 ;
        RECT 79.780 5.810 80.060 6.950 ;
        RECT 80.695 6.800 90.245 7.030 ;
        RECT 80.595 5.810 90.825 6.800 ;
        RECT 91.010 5.810 91.290 6.950 ;
        RECT 91.960 5.810 92.220 6.950 ;
        RECT 93.310 5.810 93.590 6.950 ;
        RECT 94.260 5.810 94.520 6.950 ;
        RECT 94.690 5.810 94.950 6.950 ;
        RECT 95.620 5.810 95.900 6.950 ;
        RECT 96.070 5.810 96.330 6.950 ;
        RECT 97.000 5.810 97.280 6.950 ;
        RECT 97.915 6.800 103.900 7.030 ;
        RECT 97.815 5.810 103.900 6.800 ;
        RECT 0.000 5.645 103.900 5.810 ;
        RECT 0.000 5.640 56.380 5.645 ;
        RECT 0.000 5.425 21.940 5.640 ;
        RECT 21.730 4.500 21.940 5.425 ;
        RECT 22.610 4.500 22.840 5.640 ;
        RECT 23.060 4.500 23.390 5.640 ;
        RECT 25.300 4.500 25.630 5.640 ;
        RECT 26.880 5.130 27.050 5.640 ;
        RECT 27.720 4.790 27.890 5.640 ;
        RECT 29.030 5.430 39.160 5.640 ;
        RECT 30.140 5.425 39.160 5.430 ;
        RECT 30.310 4.695 30.480 5.425 ;
        RECT 33.055 4.695 33.225 5.425 ;
        RECT 34.040 4.695 34.210 5.425 ;
        RECT 38.950 4.500 39.160 5.425 ;
        RECT 39.830 4.500 40.060 5.640 ;
        RECT 40.280 4.500 40.610 5.640 ;
        RECT 42.520 4.500 42.850 5.640 ;
        RECT 44.100 5.130 44.270 5.640 ;
        RECT 44.940 4.790 45.110 5.640 ;
        RECT 46.250 5.430 56.380 5.640 ;
        RECT 47.360 5.425 52.080 5.430 ;
        RECT 47.530 4.695 47.700 5.425 ;
        RECT 50.275 4.695 50.445 5.425 ;
        RECT 51.260 4.695 51.430 5.425 ;
        RECT 56.170 4.505 56.380 5.430 ;
        RECT 57.050 4.505 57.280 5.645 ;
        RECT 57.500 4.505 57.830 5.645 ;
        RECT 59.740 4.505 60.070 5.645 ;
        RECT 61.320 5.135 61.490 5.645 ;
        RECT 62.160 4.795 62.330 5.645 ;
        RECT 63.470 5.640 103.900 5.645 ;
        RECT 63.470 5.435 73.600 5.640 ;
        RECT 63.475 5.430 73.600 5.435 ;
        RECT 64.750 4.700 64.920 5.430 ;
        RECT 67.495 4.700 67.665 5.430 ;
        RECT 68.480 4.700 68.650 5.430 ;
        RECT 69.455 5.425 73.600 5.430 ;
        RECT 73.390 4.500 73.600 5.425 ;
        RECT 74.270 4.500 74.500 5.640 ;
        RECT 74.720 4.500 75.050 5.640 ;
        RECT 76.960 4.500 77.290 5.640 ;
        RECT 78.540 5.130 78.710 5.640 ;
        RECT 79.380 4.790 79.550 5.640 ;
        RECT 80.690 5.430 90.820 5.640 ;
        RECT 81.800 5.425 90.820 5.430 ;
        RECT 81.970 4.695 82.140 5.425 ;
        RECT 84.715 4.695 84.885 5.425 ;
        RECT 85.700 4.695 85.870 5.425 ;
        RECT 90.610 4.500 90.820 5.425 ;
        RECT 91.490 4.500 91.720 5.640 ;
        RECT 91.940 4.500 92.270 5.640 ;
        RECT 94.180 4.500 94.510 5.640 ;
        RECT 95.760 5.130 95.930 5.640 ;
        RECT 96.600 4.790 96.770 5.640 ;
        RECT 97.910 5.430 103.900 5.640 ;
        RECT 99.020 5.425 103.740 5.430 ;
        RECT 99.190 4.695 99.360 5.425 ;
        RECT 101.935 4.695 102.105 5.425 ;
        RECT 102.920 4.695 103.090 5.425 ;
      LAYER met1 ;
        RECT 16.970 9.145 17.260 9.175 ;
        RECT 16.800 8.975 17.260 9.145 ;
        RECT 16.970 8.945 17.260 8.975 ;
        RECT 15.045 7.025 17.795 7.035 ;
        RECT 18.455 7.025 21.205 7.035 ;
        RECT 30.140 7.030 34.865 7.035 ;
        RECT 35.675 7.030 38.425 7.035 ;
        RECT 47.360 7.030 52.085 7.035 ;
        RECT 52.895 7.030 55.645 7.040 ;
        RECT 64.580 7.035 69.305 7.040 ;
        RECT 63.475 7.030 69.460 7.035 ;
        RECT 70.115 7.030 72.865 7.035 ;
        RECT 81.800 7.030 86.525 7.035 ;
        RECT 87.335 7.030 90.085 7.035 ;
        RECT 99.020 7.030 103.745 7.035 ;
        RECT 0.000 7.000 21.470 7.025 ;
        RECT 29.035 7.005 38.580 7.030 ;
        RECT 0.000 6.800 21.940 7.000 ;
        RECT 29.035 6.955 38.585 7.005 ;
        RECT 46.255 6.955 55.805 7.030 ;
        RECT 63.475 6.960 73.025 7.030 ;
        RECT 28.945 6.800 38.585 6.955 ;
        RECT 46.165 6.805 55.805 6.955 ;
        RECT 63.385 6.805 73.025 6.960 ;
        RECT 80.695 6.955 90.245 7.030 ;
        RECT 97.915 6.955 103.900 7.030 ;
        RECT 46.165 6.800 56.385 6.805 ;
        RECT 0.000 5.965 21.945 6.800 ;
        RECT 28.935 5.965 39.165 6.800 ;
        RECT 46.155 5.970 56.385 6.800 ;
        RECT 63.375 6.800 73.025 6.805 ;
        RECT 80.605 6.800 90.245 6.955 ;
        RECT 97.825 6.800 103.900 6.955 ;
        RECT 63.375 5.970 73.605 6.800 ;
        RECT 46.155 5.965 73.605 5.970 ;
        RECT 80.595 5.965 90.825 6.800 ;
        RECT 97.815 5.965 103.900 6.800 ;
        RECT 0.000 5.490 103.900 5.965 ;
        RECT 0.000 5.485 56.380 5.490 ;
        RECT 0.000 5.425 21.940 5.485 ;
        RECT 29.030 5.430 39.160 5.485 ;
        RECT 46.250 5.430 56.380 5.485 ;
        RECT 63.470 5.485 103.900 5.490 ;
        RECT 63.470 5.435 73.600 5.485 ;
        RECT 63.475 5.430 73.600 5.435 ;
        RECT 80.690 5.430 90.820 5.485 ;
        RECT 97.910 5.430 103.900 5.485 ;
        RECT 30.140 5.425 39.160 5.430 ;
        RECT 47.360 5.425 52.080 5.430 ;
        RECT 69.455 5.425 73.600 5.430 ;
        RECT 81.800 5.425 90.820 5.430 ;
        RECT 99.020 5.425 103.740 5.430 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 52.235 12.460 69.475 12.465 ;
        RECT 0.045 10.860 103.915 12.460 ;
        RECT 15.215 10.235 15.385 10.860 ;
        RECT 18.625 10.235 18.795 10.860 ;
        RECT 19.580 10.315 19.750 10.595 ;
        RECT 19.580 10.145 19.810 10.315 ;
        RECT 19.640 8.535 19.810 10.145 ;
        RECT 19.580 8.365 19.810 8.535 ;
        RECT 21.585 8.530 21.910 10.860 ;
        RECT 22.235 8.530 22.560 10.860 ;
        RECT 22.885 8.530 23.210 10.860 ;
        RECT 23.535 8.530 23.860 10.860 ;
        RECT 24.185 8.530 24.510 10.860 ;
        RECT 24.835 8.530 25.160 10.860 ;
        RECT 25.485 8.530 25.810 10.860 ;
        RECT 26.135 8.530 26.460 10.860 ;
        RECT 26.785 8.530 27.110 10.860 ;
        RECT 27.435 8.530 27.760 10.860 ;
        RECT 28.085 8.530 28.410 10.860 ;
        RECT 28.735 8.530 28.945 10.860 ;
        RECT 30.310 10.235 30.480 10.860 ;
        RECT 33.055 10.235 33.225 10.860 ;
        RECT 34.045 10.235 34.215 10.860 ;
        RECT 35.845 10.235 36.015 10.860 ;
        RECT 36.800 10.315 36.970 10.595 ;
        RECT 36.800 10.145 37.030 10.315 ;
        RECT 36.860 8.535 37.030 10.145 ;
        RECT 19.580 7.305 19.750 8.365 ;
        RECT 21.585 8.360 28.945 8.530 ;
        RECT 36.800 8.365 37.030 8.535 ;
        RECT 38.805 8.530 39.130 10.860 ;
        RECT 39.455 8.530 39.780 10.860 ;
        RECT 40.105 8.530 40.430 10.860 ;
        RECT 40.755 8.530 41.080 10.860 ;
        RECT 41.405 8.530 41.730 10.860 ;
        RECT 42.055 8.530 42.380 10.860 ;
        RECT 42.705 8.530 43.030 10.860 ;
        RECT 43.355 8.530 43.680 10.860 ;
        RECT 44.005 8.530 44.330 10.860 ;
        RECT 44.655 8.530 44.980 10.860 ;
        RECT 45.305 8.530 45.630 10.860 ;
        RECT 45.955 8.530 46.165 10.860 ;
        RECT 47.530 10.235 47.700 10.860 ;
        RECT 50.275 10.235 50.445 10.860 ;
        RECT 51.265 10.235 51.435 10.860 ;
        RECT 53.065 10.240 53.235 10.860 ;
        RECT 54.020 10.320 54.190 10.600 ;
        RECT 54.020 10.150 54.250 10.320 ;
        RECT 54.080 8.540 54.250 10.150 ;
        RECT 22.130 7.560 22.440 8.360 ;
        RECT 22.140 7.340 22.475 7.390 ;
        RECT 24.060 7.340 24.230 8.360 ;
        RECT 24.430 7.560 24.740 8.360 ;
        RECT 26.710 7.560 27.020 8.360 ;
        RECT 28.090 7.560 28.400 8.360 ;
        RECT 24.440 7.340 24.775 7.390 ;
        RECT 21.670 7.170 22.475 7.340 ;
        RECT 24.050 7.170 24.775 7.340 ;
        RECT 36.800 7.305 36.970 8.365 ;
        RECT 38.805 8.360 46.165 8.530 ;
        RECT 54.020 8.370 54.250 8.540 ;
        RECT 56.025 8.535 56.350 10.860 ;
        RECT 56.675 8.535 57.000 10.860 ;
        RECT 57.325 8.535 57.650 10.860 ;
        RECT 57.975 8.535 58.300 10.860 ;
        RECT 58.625 8.535 58.950 10.860 ;
        RECT 59.275 8.535 59.600 10.860 ;
        RECT 59.925 8.535 60.250 10.860 ;
        RECT 60.575 8.535 60.900 10.860 ;
        RECT 61.225 8.535 61.550 10.860 ;
        RECT 61.875 8.535 62.200 10.860 ;
        RECT 62.525 8.535 62.850 10.860 ;
        RECT 63.175 8.535 63.385 10.860 ;
        RECT 64.750 10.240 64.920 10.860 ;
        RECT 67.495 10.240 67.665 10.860 ;
        RECT 68.485 10.240 68.655 10.860 ;
        RECT 70.285 10.235 70.455 10.860 ;
        RECT 71.240 10.315 71.410 10.595 ;
        RECT 71.240 10.145 71.470 10.315 ;
        RECT 71.300 8.535 71.470 10.145 ;
        RECT 39.350 7.560 39.660 8.360 ;
        RECT 39.360 7.340 39.695 7.390 ;
        RECT 41.280 7.340 41.450 8.360 ;
        RECT 41.650 7.560 41.960 8.360 ;
        RECT 43.930 7.560 44.240 8.360 ;
        RECT 45.310 7.560 45.620 8.360 ;
        RECT 41.660 7.340 41.995 7.390 ;
        RECT 38.890 7.170 39.695 7.340 ;
        RECT 41.270 7.170 41.995 7.340 ;
        RECT 54.020 7.310 54.190 8.370 ;
        RECT 56.025 8.365 63.385 8.535 ;
        RECT 71.240 8.365 71.470 8.535 ;
        RECT 73.245 8.530 73.570 10.860 ;
        RECT 73.895 8.530 74.220 10.860 ;
        RECT 74.545 8.530 74.870 10.860 ;
        RECT 75.195 8.530 75.520 10.860 ;
        RECT 75.845 8.530 76.170 10.860 ;
        RECT 76.495 8.530 76.820 10.860 ;
        RECT 77.145 8.530 77.470 10.860 ;
        RECT 77.795 8.530 78.120 10.860 ;
        RECT 78.445 8.530 78.770 10.860 ;
        RECT 79.095 8.530 79.420 10.860 ;
        RECT 79.745 8.530 80.070 10.860 ;
        RECT 80.395 8.530 80.605 10.860 ;
        RECT 81.970 10.235 82.140 10.860 ;
        RECT 84.715 10.235 84.885 10.860 ;
        RECT 85.705 10.235 85.875 10.860 ;
        RECT 87.505 10.235 87.675 10.860 ;
        RECT 88.460 10.315 88.630 10.595 ;
        RECT 88.460 10.145 88.690 10.315 ;
        RECT 88.520 8.535 88.690 10.145 ;
        RECT 56.570 7.565 56.880 8.365 ;
        RECT 56.580 7.345 56.915 7.395 ;
        RECT 58.500 7.345 58.670 8.365 ;
        RECT 58.870 7.565 59.180 8.365 ;
        RECT 61.150 7.565 61.460 8.365 ;
        RECT 62.530 7.565 62.840 8.365 ;
        RECT 58.880 7.345 59.215 7.395 ;
        RECT 56.110 7.175 56.915 7.345 ;
        RECT 58.490 7.175 59.215 7.345 ;
        RECT 71.240 7.305 71.410 8.365 ;
        RECT 73.245 8.360 80.605 8.530 ;
        RECT 88.460 8.365 88.690 8.535 ;
        RECT 90.465 8.530 90.790 10.860 ;
        RECT 91.115 8.530 91.440 10.860 ;
        RECT 91.765 8.530 92.090 10.860 ;
        RECT 92.415 8.530 92.740 10.860 ;
        RECT 93.065 8.530 93.390 10.860 ;
        RECT 93.715 8.530 94.040 10.860 ;
        RECT 94.365 8.530 94.690 10.860 ;
        RECT 95.015 8.530 95.340 10.860 ;
        RECT 95.665 8.530 95.990 10.860 ;
        RECT 96.315 8.530 96.640 10.860 ;
        RECT 96.965 8.530 97.290 10.860 ;
        RECT 97.615 8.530 97.825 10.860 ;
        RECT 99.190 10.235 99.360 10.860 ;
        RECT 101.935 10.235 102.105 10.860 ;
        RECT 102.925 10.235 103.095 10.860 ;
        RECT 73.790 7.560 74.100 8.360 ;
        RECT 73.800 7.340 74.135 7.390 ;
        RECT 75.720 7.340 75.890 8.360 ;
        RECT 76.090 7.560 76.400 8.360 ;
        RECT 78.370 7.560 78.680 8.360 ;
        RECT 79.750 7.560 80.060 8.360 ;
        RECT 76.100 7.340 76.435 7.390 ;
        RECT 22.140 7.120 22.475 7.170 ;
        RECT 24.440 7.120 24.775 7.170 ;
        RECT 39.360 7.120 39.695 7.170 ;
        RECT 41.660 7.120 41.995 7.170 ;
        RECT 56.580 7.125 56.915 7.175 ;
        RECT 58.880 7.125 59.215 7.175 ;
        RECT 73.330 7.170 74.135 7.340 ;
        RECT 75.710 7.170 76.435 7.340 ;
        RECT 88.460 7.305 88.630 8.365 ;
        RECT 90.465 8.360 97.825 8.530 ;
        RECT 91.010 7.560 91.320 8.360 ;
        RECT 91.020 7.340 91.355 7.390 ;
        RECT 92.940 7.340 93.110 8.360 ;
        RECT 93.310 7.560 93.620 8.360 ;
        RECT 95.590 7.560 95.900 8.360 ;
        RECT 96.970 7.560 97.280 8.360 ;
        RECT 93.320 7.340 93.655 7.390 ;
        RECT 90.550 7.170 91.355 7.340 ;
        RECT 92.930 7.170 93.655 7.340 ;
        RECT 73.800 7.120 74.135 7.170 ;
        RECT 76.100 7.120 76.435 7.170 ;
        RECT 91.020 7.120 91.355 7.170 ;
        RECT 93.320 7.120 93.655 7.170 ;
      LAYER met1 ;
        RECT 52.235 12.460 69.475 12.465 ;
        RECT 0.045 10.860 103.915 12.460 ;
        RECT 19.175 8.785 19.345 10.860 ;
        RECT 19.580 8.785 19.870 8.815 ;
        RECT 19.175 8.600 19.870 8.785 ;
        RECT 19.580 8.585 19.870 8.600 ;
        RECT 21.585 8.685 21.910 10.860 ;
        RECT 22.235 8.685 22.560 10.860 ;
        RECT 22.885 8.685 23.210 10.860 ;
        RECT 23.535 8.685 23.860 10.860 ;
        RECT 24.185 8.685 24.510 10.860 ;
        RECT 24.835 8.685 25.160 10.860 ;
        RECT 25.485 8.685 25.810 10.860 ;
        RECT 26.135 8.685 26.460 10.860 ;
        RECT 26.785 8.685 27.110 10.860 ;
        RECT 27.435 8.685 27.760 10.860 ;
        RECT 28.085 8.685 28.410 10.860 ;
        RECT 28.735 8.685 28.945 10.860 ;
        RECT 21.585 8.330 28.945 8.685 ;
        RECT 36.395 8.785 36.565 10.860 ;
        RECT 36.800 8.785 37.090 8.815 ;
        RECT 36.395 8.600 37.090 8.785 ;
        RECT 36.800 8.585 37.090 8.600 ;
        RECT 38.805 8.685 39.130 10.860 ;
        RECT 39.455 8.685 39.780 10.860 ;
        RECT 40.105 8.685 40.430 10.860 ;
        RECT 40.755 8.685 41.080 10.860 ;
        RECT 41.405 8.685 41.730 10.860 ;
        RECT 42.055 8.685 42.380 10.860 ;
        RECT 42.705 8.685 43.030 10.860 ;
        RECT 43.355 8.685 43.680 10.860 ;
        RECT 44.005 8.685 44.330 10.860 ;
        RECT 44.655 8.685 44.980 10.860 ;
        RECT 45.305 8.685 45.630 10.860 ;
        RECT 45.955 8.685 46.165 10.860 ;
        RECT 38.805 8.330 46.165 8.685 ;
        RECT 53.615 8.790 53.785 10.860 ;
        RECT 54.020 8.790 54.310 8.820 ;
        RECT 53.615 8.605 54.310 8.790 ;
        RECT 54.020 8.590 54.310 8.605 ;
        RECT 56.025 8.690 56.350 10.860 ;
        RECT 56.675 8.690 57.000 10.860 ;
        RECT 57.325 8.690 57.650 10.860 ;
        RECT 57.975 8.690 58.300 10.860 ;
        RECT 58.625 8.690 58.950 10.860 ;
        RECT 59.275 8.690 59.600 10.860 ;
        RECT 59.925 8.690 60.250 10.860 ;
        RECT 60.575 8.690 60.900 10.860 ;
        RECT 61.225 8.690 61.550 10.860 ;
        RECT 61.875 8.690 62.200 10.860 ;
        RECT 62.525 8.690 62.850 10.860 ;
        RECT 63.175 8.690 63.385 10.860 ;
        RECT 56.025 8.335 63.385 8.690 ;
        RECT 70.835 8.785 71.005 10.860 ;
        RECT 71.240 8.785 71.530 8.815 ;
        RECT 70.835 8.600 71.530 8.785 ;
        RECT 71.240 8.585 71.530 8.600 ;
        RECT 73.245 8.685 73.570 10.860 ;
        RECT 73.895 8.685 74.220 10.860 ;
        RECT 74.545 8.685 74.870 10.860 ;
        RECT 75.195 8.685 75.520 10.860 ;
        RECT 75.845 8.685 76.170 10.860 ;
        RECT 76.495 8.685 76.820 10.860 ;
        RECT 77.145 8.685 77.470 10.860 ;
        RECT 77.795 8.685 78.120 10.860 ;
        RECT 78.445 8.685 78.770 10.860 ;
        RECT 79.095 8.685 79.420 10.860 ;
        RECT 79.745 8.685 80.070 10.860 ;
        RECT 80.395 8.685 80.605 10.860 ;
        RECT 73.245 8.330 80.605 8.685 ;
        RECT 88.055 8.785 88.225 10.860 ;
        RECT 88.460 8.785 88.750 8.815 ;
        RECT 88.055 8.600 88.750 8.785 ;
        RECT 88.460 8.585 88.750 8.600 ;
        RECT 90.465 8.685 90.790 10.860 ;
        RECT 91.115 8.685 91.440 10.860 ;
        RECT 91.765 8.685 92.090 10.860 ;
        RECT 92.415 8.685 92.740 10.860 ;
        RECT 93.065 8.685 93.390 10.860 ;
        RECT 93.715 8.685 94.040 10.860 ;
        RECT 94.365 8.685 94.690 10.860 ;
        RECT 95.015 8.685 95.340 10.860 ;
        RECT 95.665 8.685 95.990 10.860 ;
        RECT 96.315 8.685 96.640 10.860 ;
        RECT 96.965 8.685 97.290 10.860 ;
        RECT 97.615 8.685 97.825 10.860 ;
        RECT 90.465 8.330 97.825 8.685 ;
        RECT 21.610 7.325 21.900 7.370 ;
        RECT 23.975 7.325 24.295 7.385 ;
        RECT 21.610 7.185 24.295 7.325 ;
        RECT 21.610 7.140 21.900 7.185 ;
        RECT 23.975 7.125 24.295 7.185 ;
        RECT 38.830 7.325 39.120 7.370 ;
        RECT 41.195 7.325 41.515 7.385 ;
        RECT 38.830 7.185 41.515 7.325 ;
        RECT 38.830 7.140 39.120 7.185 ;
        RECT 41.195 7.125 41.515 7.185 ;
        RECT 56.050 7.330 56.340 7.375 ;
        RECT 58.415 7.330 58.735 7.390 ;
        RECT 56.050 7.190 58.735 7.330 ;
        RECT 56.050 7.145 56.340 7.190 ;
        RECT 58.415 7.130 58.735 7.190 ;
        RECT 73.270 7.325 73.560 7.370 ;
        RECT 75.635 7.325 75.955 7.385 ;
        RECT 73.270 7.185 75.955 7.325 ;
        RECT 73.270 7.140 73.560 7.185 ;
        RECT 75.635 7.125 75.955 7.185 ;
        RECT 90.490 7.325 90.780 7.370 ;
        RECT 92.855 7.325 93.175 7.385 ;
        RECT 90.490 7.185 93.175 7.325 ;
        RECT 90.490 7.140 90.780 7.185 ;
        RECT 92.855 7.125 93.175 7.185 ;
      LAYER met2 ;
        RECT 23.995 7.065 24.275 7.435 ;
        RECT 41.215 7.065 41.495 7.435 ;
        RECT 58.435 7.070 58.715 7.440 ;
        RECT 75.655 7.065 75.935 7.435 ;
        RECT 92.875 7.065 93.155 7.435 ;
      LAYER met3 ;
        RECT 23.970 7.400 24.300 7.415 ;
        RECT 41.190 7.400 41.520 7.415 ;
        RECT 58.410 7.405 58.740 7.420 ;
        RECT 23.500 7.100 24.300 7.400 ;
        RECT 40.720 7.100 41.520 7.400 ;
        RECT 57.940 7.105 58.740 7.405 ;
        RECT 75.630 7.400 75.960 7.415 ;
        RECT 92.850 7.400 93.180 7.415 ;
        RECT 23.970 7.085 24.300 7.100 ;
        RECT 41.190 7.085 41.520 7.100 ;
        RECT 58.410 7.090 58.740 7.105 ;
        RECT 75.160 7.100 75.960 7.400 ;
        RECT 92.380 7.100 93.180 7.400 ;
        RECT 75.630 7.085 75.960 7.100 ;
        RECT 92.850 7.085 93.180 7.100 ;
    END
    PORT
      LAYER li1 ;
        RECT 21.730 3.090 21.940 3.910 ;
        RECT 22.610 3.090 22.840 3.910 ;
        RECT 23.060 3.090 23.330 3.900 ;
        RECT 24.000 3.090 24.240 3.900 ;
        RECT 24.450 3.090 24.690 3.900 ;
        RECT 25.360 3.090 25.630 3.900 ;
        RECT 25.810 3.090 26.100 3.925 ;
        RECT 27.640 3.090 27.970 3.480 ;
        RECT 28.480 3.090 28.810 3.480 ;
        RECT 38.950 3.090 39.160 3.910 ;
        RECT 39.830 3.090 40.060 3.910 ;
        RECT 40.280 3.090 40.550 3.900 ;
        RECT 41.220 3.090 41.460 3.900 ;
        RECT 41.670 3.090 41.910 3.900 ;
        RECT 42.580 3.090 42.850 3.900 ;
        RECT 43.030 3.090 43.320 3.925 ;
        RECT 44.860 3.090 45.190 3.480 ;
        RECT 45.700 3.090 46.030 3.480 ;
        RECT 56.170 3.095 56.380 3.915 ;
        RECT 57.050 3.095 57.280 3.915 ;
        RECT 57.500 3.095 57.770 3.905 ;
        RECT 58.440 3.095 58.680 3.905 ;
        RECT 58.890 3.095 59.130 3.905 ;
        RECT 59.800 3.095 60.070 3.905 ;
        RECT 60.250 3.095 60.540 3.930 ;
        RECT 62.080 3.095 62.410 3.485 ;
        RECT 62.920 3.095 63.250 3.485 ;
        RECT 21.580 2.920 29.325 3.090 ;
        RECT 21.580 1.600 21.925 2.920 ;
        RECT 22.270 1.600 22.600 2.920 ;
        RECT 22.945 1.605 23.290 2.920 ;
        RECT 23.635 1.605 23.980 2.920 ;
        RECT 24.325 1.605 24.670 2.920 ;
        RECT 25.015 1.605 25.360 2.920 ;
        RECT 25.705 1.605 26.050 2.920 ;
        RECT 26.395 1.605 26.740 2.920 ;
        RECT 27.085 1.605 27.430 2.920 ;
        RECT 27.775 1.605 28.120 2.920 ;
        RECT 28.465 1.605 28.810 2.920 ;
        RECT 29.155 1.605 29.325 2.920 ;
        RECT 38.800 2.920 46.545 3.090 ;
        RECT 22.945 1.600 29.325 1.605 ;
        RECT 30.310 1.600 30.480 2.225 ;
        RECT 33.055 1.600 33.225 2.225 ;
        RECT 34.040 1.600 34.210 2.225 ;
        RECT 38.800 1.600 39.145 2.920 ;
        RECT 39.490 1.600 39.820 2.920 ;
        RECT 40.165 1.605 40.510 2.920 ;
        RECT 40.855 1.605 41.200 2.920 ;
        RECT 41.545 1.605 41.890 2.920 ;
        RECT 42.235 1.605 42.580 2.920 ;
        RECT 42.925 1.605 43.270 2.920 ;
        RECT 43.615 1.605 43.960 2.920 ;
        RECT 44.305 1.605 44.650 2.920 ;
        RECT 44.995 1.605 45.340 2.920 ;
        RECT 45.685 1.605 46.030 2.920 ;
        RECT 46.375 1.605 46.545 2.920 ;
        RECT 56.020 2.925 63.765 3.095 ;
        RECT 73.390 3.090 73.600 3.910 ;
        RECT 74.270 3.090 74.500 3.910 ;
        RECT 74.720 3.090 74.990 3.900 ;
        RECT 75.660 3.090 75.900 3.900 ;
        RECT 76.110 3.090 76.350 3.900 ;
        RECT 77.020 3.090 77.290 3.900 ;
        RECT 77.470 3.090 77.760 3.925 ;
        RECT 79.300 3.090 79.630 3.480 ;
        RECT 80.140 3.090 80.470 3.480 ;
        RECT 90.610 3.090 90.820 3.910 ;
        RECT 91.490 3.090 91.720 3.910 ;
        RECT 91.940 3.090 92.210 3.900 ;
        RECT 92.880 3.090 93.120 3.900 ;
        RECT 93.330 3.090 93.570 3.900 ;
        RECT 94.240 3.090 94.510 3.900 ;
        RECT 94.690 3.090 94.980 3.925 ;
        RECT 96.520 3.090 96.850 3.480 ;
        RECT 97.360 3.090 97.690 3.480 ;
        RECT 40.165 1.600 46.545 1.605 ;
        RECT 47.530 1.600 47.700 2.225 ;
        RECT 50.275 1.600 50.445 2.225 ;
        RECT 51.260 1.600 51.430 2.225 ;
        RECT 56.020 1.605 56.365 2.925 ;
        RECT 56.710 1.605 57.040 2.925 ;
        RECT 57.385 1.610 57.730 2.925 ;
        RECT 58.075 1.610 58.420 2.925 ;
        RECT 58.765 1.610 59.110 2.925 ;
        RECT 59.455 1.610 59.800 2.925 ;
        RECT 60.145 1.610 60.490 2.925 ;
        RECT 60.835 1.610 61.180 2.925 ;
        RECT 61.525 1.610 61.870 2.925 ;
        RECT 62.215 1.610 62.560 2.925 ;
        RECT 62.905 1.610 63.250 2.925 ;
        RECT 63.595 1.610 63.765 2.925 ;
        RECT 73.240 2.920 80.985 3.090 ;
        RECT 57.385 1.605 63.765 1.610 ;
        RECT 64.750 1.605 64.920 2.230 ;
        RECT 67.495 1.605 67.665 2.230 ;
        RECT 68.480 1.605 68.650 2.230 ;
        RECT 52.235 1.600 69.475 1.605 ;
        RECT 73.240 1.600 73.585 2.920 ;
        RECT 73.930 1.600 74.260 2.920 ;
        RECT 74.605 1.605 74.950 2.920 ;
        RECT 75.295 1.605 75.640 2.920 ;
        RECT 75.985 1.605 76.330 2.920 ;
        RECT 76.675 1.605 77.020 2.920 ;
        RECT 77.365 1.605 77.710 2.920 ;
        RECT 78.055 1.605 78.400 2.920 ;
        RECT 78.745 1.605 79.090 2.920 ;
        RECT 79.435 1.605 79.780 2.920 ;
        RECT 80.125 1.605 80.470 2.920 ;
        RECT 80.815 1.605 80.985 2.920 ;
        RECT 90.460 2.920 98.205 3.090 ;
        RECT 74.605 1.600 80.985 1.605 ;
        RECT 81.970 1.600 82.140 2.225 ;
        RECT 84.715 1.600 84.885 2.225 ;
        RECT 85.700 1.600 85.870 2.225 ;
        RECT 90.460 1.600 90.805 2.920 ;
        RECT 91.150 1.600 91.480 2.920 ;
        RECT 91.825 1.605 92.170 2.920 ;
        RECT 92.515 1.605 92.860 2.920 ;
        RECT 93.205 1.605 93.550 2.920 ;
        RECT 93.895 1.605 94.240 2.920 ;
        RECT 94.585 1.605 94.930 2.920 ;
        RECT 95.275 1.605 95.620 2.920 ;
        RECT 95.965 1.605 96.310 2.920 ;
        RECT 96.655 1.605 97.000 2.920 ;
        RECT 97.345 1.605 97.690 2.920 ;
        RECT 98.035 1.605 98.205 2.920 ;
        RECT 91.825 1.600 98.205 1.605 ;
        RECT 99.190 1.600 99.360 2.225 ;
        RECT 101.935 1.600 102.105 2.225 ;
        RECT 102.920 1.600 103.090 2.225 ;
        RECT 0.045 0.000 103.915 1.600 ;
      LAYER met1 ;
        RECT 21.580 2.765 29.325 3.120 ;
        RECT 21.580 1.600 21.925 2.765 ;
        RECT 22.270 1.600 22.600 2.765 ;
        RECT 22.945 1.605 23.290 2.765 ;
        RECT 23.635 1.605 23.980 2.765 ;
        RECT 24.325 1.605 24.670 2.765 ;
        RECT 25.015 1.605 25.360 2.765 ;
        RECT 25.705 1.605 26.050 2.765 ;
        RECT 26.395 1.605 26.740 2.765 ;
        RECT 27.085 1.605 27.430 2.765 ;
        RECT 27.775 1.605 28.120 2.765 ;
        RECT 28.465 1.605 28.810 2.765 ;
        RECT 29.155 1.605 29.325 2.765 ;
        RECT 22.945 1.600 29.325 1.605 ;
        RECT 38.800 2.765 46.545 3.120 ;
        RECT 38.800 1.600 39.145 2.765 ;
        RECT 39.490 1.600 39.820 2.765 ;
        RECT 40.165 1.605 40.510 2.765 ;
        RECT 40.855 1.605 41.200 2.765 ;
        RECT 41.545 1.605 41.890 2.765 ;
        RECT 42.235 1.605 42.580 2.765 ;
        RECT 42.925 1.605 43.270 2.765 ;
        RECT 43.615 1.605 43.960 2.765 ;
        RECT 44.305 1.605 44.650 2.765 ;
        RECT 44.995 1.605 45.340 2.765 ;
        RECT 45.685 1.605 46.030 2.765 ;
        RECT 46.375 1.605 46.545 2.765 ;
        RECT 56.020 2.770 63.765 3.125 ;
        RECT 56.020 1.605 56.365 2.770 ;
        RECT 56.710 1.605 57.040 2.770 ;
        RECT 57.385 1.610 57.730 2.770 ;
        RECT 58.075 1.610 58.420 2.770 ;
        RECT 58.765 1.610 59.110 2.770 ;
        RECT 59.455 1.610 59.800 2.770 ;
        RECT 60.145 1.610 60.490 2.770 ;
        RECT 60.835 1.610 61.180 2.770 ;
        RECT 61.525 1.610 61.870 2.770 ;
        RECT 62.215 1.610 62.560 2.770 ;
        RECT 62.905 1.610 63.250 2.770 ;
        RECT 63.595 1.610 63.765 2.770 ;
        RECT 57.385 1.605 63.765 1.610 ;
        RECT 73.240 2.765 80.985 3.120 ;
        RECT 40.165 1.600 46.545 1.605 ;
        RECT 52.235 1.600 69.475 1.605 ;
        RECT 73.240 1.600 73.585 2.765 ;
        RECT 73.930 1.600 74.260 2.765 ;
        RECT 74.605 1.605 74.950 2.765 ;
        RECT 75.295 1.605 75.640 2.765 ;
        RECT 75.985 1.605 76.330 2.765 ;
        RECT 76.675 1.605 77.020 2.765 ;
        RECT 77.365 1.605 77.710 2.765 ;
        RECT 78.055 1.605 78.400 2.765 ;
        RECT 78.745 1.605 79.090 2.765 ;
        RECT 79.435 1.605 79.780 2.765 ;
        RECT 80.125 1.605 80.470 2.765 ;
        RECT 80.815 1.605 80.985 2.765 ;
        RECT 74.605 1.600 80.985 1.605 ;
        RECT 90.460 2.765 98.205 3.120 ;
        RECT 90.460 1.600 90.805 2.765 ;
        RECT 91.150 1.600 91.480 2.765 ;
        RECT 91.825 1.605 92.170 2.765 ;
        RECT 92.515 1.605 92.860 2.765 ;
        RECT 93.205 1.605 93.550 2.765 ;
        RECT 93.895 1.605 94.240 2.765 ;
        RECT 94.585 1.605 94.930 2.765 ;
        RECT 95.275 1.605 95.620 2.765 ;
        RECT 95.965 1.605 96.310 2.765 ;
        RECT 96.655 1.605 97.000 2.765 ;
        RECT 97.345 1.605 97.690 2.765 ;
        RECT 98.035 1.605 98.205 2.765 ;
        RECT 91.825 1.600 98.205 1.605 ;
        RECT 0.045 0.000 103.915 1.600 ;
    END
  END vssd1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 86.130 4.010 86.305 5.155 ;
        RECT 86.130 3.575 86.300 4.010 ;
        RECT 86.135 1.865 86.305 2.375 ;
      LAYER met1 ;
        RECT 86.070 3.540 86.360 3.775 ;
        RECT 86.070 3.535 86.300 3.540 ;
        RECT 86.130 3.370 86.300 3.535 ;
        RECT 86.130 3.200 86.310 3.370 ;
        RECT 86.130 2.435 86.300 3.200 ;
        RECT 86.070 2.175 86.365 2.435 ;
    END
  END X4_Y1
  OBS
      LAYER pwell ;
        RECT 21.460 8.530 22.060 8.745 ;
        RECT 38.680 8.530 39.280 8.745 ;
        RECT 55.900 8.535 56.500 8.750 ;
        RECT 21.460 8.340 22.355 8.530 ;
        RECT 24.485 8.495 24.655 8.530 ;
        RECT 23.580 8.385 24.655 8.495 ;
        RECT 24.370 8.340 24.655 8.385 ;
        RECT 26.795 8.340 26.965 8.530 ;
        RECT 28.175 8.500 28.345 8.530 ;
        RECT 28.175 8.390 28.745 8.500 ;
        RECT 28.175 8.340 28.460 8.390 ;
        RECT 21.460 8.145 23.420 8.340 ;
        RECT 22.070 7.430 23.420 8.145 ;
        RECT 24.370 7.430 28.460 8.340 ;
        RECT 38.680 8.340 39.575 8.530 ;
        RECT 41.705 8.495 41.875 8.530 ;
        RECT 40.800 8.385 41.875 8.495 ;
        RECT 41.590 8.340 41.875 8.385 ;
        RECT 44.015 8.340 44.185 8.530 ;
        RECT 45.395 8.500 45.565 8.530 ;
        RECT 45.395 8.390 45.965 8.500 ;
        RECT 45.395 8.340 45.680 8.390 ;
        RECT 38.680 8.145 40.640 8.340 ;
        RECT 39.290 7.430 40.640 8.145 ;
        RECT 41.590 7.430 45.680 8.340 ;
        RECT 55.900 8.345 56.795 8.535 ;
        RECT 58.925 8.500 59.095 8.535 ;
        RECT 58.020 8.390 59.095 8.500 ;
        RECT 58.810 8.345 59.095 8.390 ;
        RECT 61.235 8.345 61.405 8.535 ;
        RECT 62.615 8.505 62.785 8.535 ;
        RECT 73.120 8.530 73.720 8.745 ;
        RECT 90.340 8.530 90.940 8.745 ;
        RECT 62.615 8.395 63.185 8.505 ;
        RECT 62.615 8.345 62.900 8.395 ;
        RECT 55.900 8.150 57.860 8.345 ;
        RECT 56.510 7.435 57.860 8.150 ;
        RECT 58.810 7.435 62.900 8.345 ;
        RECT 73.120 8.340 74.015 8.530 ;
        RECT 76.145 8.495 76.315 8.530 ;
        RECT 75.240 8.385 76.315 8.495 ;
        RECT 76.030 8.340 76.315 8.385 ;
        RECT 78.455 8.340 78.625 8.530 ;
        RECT 79.835 8.500 80.005 8.530 ;
        RECT 79.835 8.390 80.405 8.500 ;
        RECT 79.835 8.340 80.120 8.390 ;
        RECT 73.120 8.145 75.080 8.340 ;
        RECT 73.730 7.430 75.080 8.145 ;
        RECT 76.030 7.430 80.120 8.340 ;
        RECT 90.340 8.340 91.235 8.530 ;
        RECT 93.365 8.495 93.535 8.530 ;
        RECT 92.460 8.385 93.535 8.495 ;
        RECT 93.250 8.340 93.535 8.385 ;
        RECT 95.675 8.340 95.845 8.530 ;
        RECT 97.055 8.500 97.225 8.530 ;
        RECT 97.055 8.390 97.625 8.500 ;
        RECT 97.055 8.340 97.340 8.390 ;
        RECT 90.340 8.145 92.300 8.340 ;
        RECT 90.950 7.430 92.300 8.145 ;
        RECT 93.250 7.430 97.340 8.340 ;
        RECT 21.600 3.305 28.900 4.020 ;
        RECT 38.820 3.305 46.120 4.020 ;
        RECT 56.040 3.310 63.340 4.025 ;
        RECT 21.460 3.110 28.900 3.305 ;
        RECT 38.680 3.110 46.120 3.305 ;
        RECT 55.900 3.115 63.340 3.310 ;
        RECT 73.260 3.305 80.560 4.020 ;
        RECT 90.480 3.305 97.780 4.020 ;
        RECT 21.460 2.920 22.820 3.110 ;
        RECT 24.025 2.920 24.665 3.110 ;
        RECT 28.630 2.920 28.800 3.110 ;
        RECT 38.680 2.920 40.040 3.110 ;
        RECT 41.245 2.920 41.885 3.110 ;
        RECT 45.850 2.920 46.020 3.110 ;
        RECT 55.900 2.925 57.260 3.115 ;
        RECT 58.465 2.925 59.105 3.115 ;
        RECT 63.070 2.925 63.240 3.115 ;
        RECT 73.120 3.110 80.560 3.305 ;
        RECT 90.340 3.110 97.780 3.305 ;
        RECT 21.460 2.705 22.060 2.920 ;
        RECT 38.680 2.705 39.280 2.920 ;
        RECT 55.900 2.710 56.500 2.925 ;
        RECT 73.120 2.920 74.480 3.110 ;
        RECT 75.685 2.920 76.325 3.110 ;
        RECT 80.290 2.920 80.460 3.110 ;
        RECT 90.340 2.920 91.700 3.110 ;
        RECT 92.905 2.920 93.545 3.110 ;
        RECT 97.510 2.920 97.680 3.110 ;
        RECT 73.120 2.705 73.720 2.920 ;
        RECT 90.340 2.705 90.940 2.920 ;
      LAYER li1 ;
        RECT 15.645 10.105 15.820 10.595 ;
        RECT 16.170 10.315 16.340 10.595 ;
        RECT 16.170 10.145 16.400 10.315 ;
        RECT 15.645 9.935 15.815 10.105 ;
        RECT 15.645 9.605 16.055 9.935 ;
        RECT 15.645 9.095 15.815 9.605 ;
        RECT 15.645 8.765 16.055 9.095 ;
        RECT 15.645 8.565 15.815 8.765 ;
        RECT 15.645 7.305 15.820 8.565 ;
        RECT 16.230 8.535 16.400 10.145 ;
        RECT 16.600 10.085 16.775 10.595 ;
        RECT 19.055 10.105 19.230 10.595 ;
        RECT 19.055 9.935 19.225 10.105 ;
        RECT 20.010 10.085 20.185 10.595 ;
        RECT 20.440 10.045 20.615 10.595 ;
        RECT 30.740 10.105 30.915 10.595 ;
        RECT 31.265 10.315 31.435 10.595 ;
        RECT 31.265 10.145 31.495 10.315 ;
        RECT 19.055 9.605 19.465 9.935 ;
        RECT 16.170 8.365 16.400 8.535 ;
        RECT 16.600 8.565 16.770 9.515 ;
        RECT 19.055 9.095 19.225 9.605 ;
        RECT 19.055 8.765 19.465 9.095 ;
        RECT 19.055 8.565 19.225 8.765 ;
        RECT 20.010 8.565 20.180 9.515 ;
        RECT 16.170 7.305 16.340 8.365 ;
        RECT 16.600 7.305 16.775 8.565 ;
        RECT 19.055 7.305 19.230 8.565 ;
        RECT 20.010 7.305 20.185 8.565 ;
        RECT 20.440 8.445 20.610 10.045 ;
        RECT 30.740 9.935 30.910 10.105 ;
        RECT 30.740 9.605 31.150 9.935 ;
        RECT 30.740 9.095 30.910 9.605 ;
        RECT 30.740 8.765 31.150 9.095 ;
        RECT 30.740 8.565 30.910 8.765 ;
        RECT 20.440 7.305 20.615 8.445 ;
        RECT 22.645 7.560 23.340 8.190 ;
        RECT 22.645 6.960 22.815 7.560 ;
        RECT 22.985 7.340 23.320 7.370 ;
        RECT 23.710 7.340 23.880 8.020 ;
        RECT 22.985 7.170 23.880 7.340 ;
        RECT 24.945 7.560 25.640 8.190 ;
        RECT 25.810 7.560 26.505 8.190 ;
        RECT 27.190 7.560 27.885 8.190 ;
        RECT 22.985 7.120 23.320 7.170 ;
        RECT 24.945 6.960 25.115 7.560 ;
        RECT 25.285 7.340 25.620 7.370 ;
        RECT 25.830 7.340 26.165 7.370 ;
        RECT 25.285 7.170 26.165 7.340 ;
        RECT 25.285 7.120 25.620 7.170 ;
        RECT 25.830 7.120 26.165 7.170 ;
        RECT 26.335 6.960 26.505 7.560 ;
        RECT 26.675 7.120 27.010 7.390 ;
        RECT 27.210 7.120 27.545 7.370 ;
        RECT 27.715 6.960 27.885 7.560 ;
        RECT 28.055 7.120 28.390 7.390 ;
        RECT 30.740 7.305 30.915 8.565 ;
        RECT 31.325 8.535 31.495 10.145 ;
        RECT 31.695 10.085 31.870 10.595 ;
        RECT 32.125 10.045 32.300 10.595 ;
        RECT 33.490 10.085 33.660 10.595 ;
        RECT 34.480 10.085 34.650 10.595 ;
        RECT 36.275 10.105 36.450 10.595 ;
        RECT 31.265 8.365 31.495 8.535 ;
        RECT 31.695 8.565 31.865 9.515 ;
        RECT 31.265 7.305 31.435 8.365 ;
        RECT 31.695 7.305 31.870 8.565 ;
        RECT 32.125 8.445 32.295 10.045 ;
        RECT 36.275 9.935 36.445 10.105 ;
        RECT 37.230 10.085 37.405 10.595 ;
        RECT 37.660 10.045 37.835 10.595 ;
        RECT 47.960 10.105 48.135 10.595 ;
        RECT 48.485 10.315 48.655 10.595 ;
        RECT 48.485 10.145 48.715 10.315 ;
        RECT 33.055 9.425 33.285 9.615 ;
        RECT 36.275 9.605 36.685 9.935 ;
        RECT 33.055 9.385 33.585 9.425 ;
        RECT 33.115 9.255 33.585 9.385 ;
        RECT 34.105 9.255 34.575 9.425 ;
        RECT 33.115 8.565 33.285 9.255 ;
        RECT 33.485 8.780 33.655 8.885 ;
        RECT 34.105 8.780 34.275 9.255 ;
        RECT 36.275 9.095 36.445 9.605 ;
        RECT 33.485 8.605 34.275 8.780 ;
        RECT 32.125 7.305 32.300 8.445 ;
        RECT 33.485 7.305 33.660 8.605 ;
        RECT 34.105 8.565 34.275 8.605 ;
        RECT 34.475 8.450 34.645 8.885 ;
        RECT 36.275 8.765 36.685 9.095 ;
        RECT 36.275 8.565 36.445 8.765 ;
        RECT 37.230 8.565 37.400 9.515 ;
        RECT 34.475 7.305 34.650 8.450 ;
        RECT 36.275 7.305 36.450 8.565 ;
        RECT 37.230 7.305 37.405 8.565 ;
        RECT 37.660 8.445 37.830 10.045 ;
        RECT 47.960 9.935 48.130 10.105 ;
        RECT 47.960 9.605 48.370 9.935 ;
        RECT 47.960 9.095 48.130 9.605 ;
        RECT 47.960 8.765 48.370 9.095 ;
        RECT 47.960 8.565 48.130 8.765 ;
        RECT 37.660 7.305 37.835 8.445 ;
        RECT 39.865 7.560 40.560 8.190 ;
        RECT 39.865 6.960 40.035 7.560 ;
        RECT 40.205 7.340 40.540 7.370 ;
        RECT 40.930 7.340 41.100 8.020 ;
        RECT 40.205 7.170 41.100 7.340 ;
        RECT 42.165 7.560 42.860 8.190 ;
        RECT 43.030 7.560 43.725 8.190 ;
        RECT 44.410 7.560 45.105 8.190 ;
        RECT 40.205 7.120 40.540 7.170 ;
        RECT 42.165 6.960 42.335 7.560 ;
        RECT 42.505 7.340 42.840 7.370 ;
        RECT 43.050 7.340 43.385 7.370 ;
        RECT 42.505 7.170 43.385 7.340 ;
        RECT 42.505 7.120 42.840 7.170 ;
        RECT 43.050 7.120 43.385 7.170 ;
        RECT 43.555 6.960 43.725 7.560 ;
        RECT 43.895 7.120 44.230 7.390 ;
        RECT 44.430 7.120 44.765 7.370 ;
        RECT 44.935 6.960 45.105 7.560 ;
        RECT 45.275 7.120 45.610 7.390 ;
        RECT 47.960 7.305 48.135 8.565 ;
        RECT 48.545 8.535 48.715 10.145 ;
        RECT 48.915 10.085 49.090 10.595 ;
        RECT 49.345 10.045 49.520 10.595 ;
        RECT 50.710 10.085 50.880 10.595 ;
        RECT 51.700 10.085 51.870 10.595 ;
        RECT 53.495 10.110 53.670 10.600 ;
        RECT 48.485 8.365 48.715 8.535 ;
        RECT 48.915 8.565 49.085 9.515 ;
        RECT 48.485 7.305 48.655 8.365 ;
        RECT 48.915 7.305 49.090 8.565 ;
        RECT 49.345 8.445 49.515 10.045 ;
        RECT 53.495 9.940 53.665 10.110 ;
        RECT 54.450 10.090 54.625 10.600 ;
        RECT 54.880 10.050 55.055 10.600 ;
        RECT 65.180 10.110 65.355 10.600 ;
        RECT 65.705 10.320 65.875 10.600 ;
        RECT 65.705 10.150 65.935 10.320 ;
        RECT 50.275 9.425 50.505 9.615 ;
        RECT 53.495 9.610 53.905 9.940 ;
        RECT 50.275 9.385 50.805 9.425 ;
        RECT 50.335 9.255 50.805 9.385 ;
        RECT 51.325 9.255 51.795 9.425 ;
        RECT 50.335 8.565 50.505 9.255 ;
        RECT 50.705 8.780 50.875 8.885 ;
        RECT 51.325 8.780 51.495 9.255 ;
        RECT 53.495 9.100 53.665 9.610 ;
        RECT 50.705 8.605 51.495 8.780 ;
        RECT 49.345 7.305 49.520 8.445 ;
        RECT 50.705 7.305 50.880 8.605 ;
        RECT 51.325 8.565 51.495 8.605 ;
        RECT 51.695 8.450 51.865 8.885 ;
        RECT 53.495 8.770 53.905 9.100 ;
        RECT 53.495 8.570 53.665 8.770 ;
        RECT 54.450 8.570 54.620 9.520 ;
        RECT 51.695 7.305 51.870 8.450 ;
        RECT 53.495 7.310 53.670 8.570 ;
        RECT 54.450 7.310 54.625 8.570 ;
        RECT 54.880 8.450 55.050 10.050 ;
        RECT 65.180 9.940 65.350 10.110 ;
        RECT 65.180 9.610 65.590 9.940 ;
        RECT 65.180 9.100 65.350 9.610 ;
        RECT 65.180 8.770 65.590 9.100 ;
        RECT 65.180 8.570 65.350 8.770 ;
        RECT 54.880 7.310 55.055 8.450 ;
        RECT 57.085 7.565 57.780 8.195 ;
        RECT 57.085 6.965 57.255 7.565 ;
        RECT 57.425 7.345 57.760 7.375 ;
        RECT 58.150 7.345 58.320 8.025 ;
        RECT 57.425 7.175 58.320 7.345 ;
        RECT 59.385 7.565 60.080 8.195 ;
        RECT 60.250 7.565 60.945 8.195 ;
        RECT 61.630 7.565 62.325 8.195 ;
        RECT 57.425 7.125 57.760 7.175 ;
        RECT 59.385 6.965 59.555 7.565 ;
        RECT 59.725 7.345 60.060 7.375 ;
        RECT 60.270 7.345 60.605 7.375 ;
        RECT 59.725 7.175 60.605 7.345 ;
        RECT 59.725 7.125 60.060 7.175 ;
        RECT 60.270 7.125 60.605 7.175 ;
        RECT 60.775 6.965 60.945 7.565 ;
        RECT 61.115 7.125 61.450 7.395 ;
        RECT 61.650 7.125 61.985 7.375 ;
        RECT 62.155 6.965 62.325 7.565 ;
        RECT 62.495 7.125 62.830 7.395 ;
        RECT 65.180 7.310 65.355 8.570 ;
        RECT 65.765 8.540 65.935 10.150 ;
        RECT 66.135 10.090 66.310 10.600 ;
        RECT 66.565 10.050 66.740 10.600 ;
        RECT 67.930 10.090 68.100 10.600 ;
        RECT 68.920 10.090 69.090 10.600 ;
        RECT 70.715 10.105 70.890 10.595 ;
        RECT 65.705 8.370 65.935 8.540 ;
        RECT 66.135 8.570 66.305 9.520 ;
        RECT 65.705 7.310 65.875 8.370 ;
        RECT 66.135 7.310 66.310 8.570 ;
        RECT 66.565 8.450 66.735 10.050 ;
        RECT 70.715 9.935 70.885 10.105 ;
        RECT 71.670 10.085 71.845 10.595 ;
        RECT 72.100 10.045 72.275 10.595 ;
        RECT 82.400 10.105 82.575 10.595 ;
        RECT 82.925 10.315 83.095 10.595 ;
        RECT 82.925 10.145 83.155 10.315 ;
        RECT 67.495 9.430 67.725 9.620 ;
        RECT 70.715 9.605 71.125 9.935 ;
        RECT 67.495 9.390 68.025 9.430 ;
        RECT 67.555 9.260 68.025 9.390 ;
        RECT 68.545 9.260 69.015 9.430 ;
        RECT 67.555 8.570 67.725 9.260 ;
        RECT 67.925 8.785 68.095 8.890 ;
        RECT 68.545 8.785 68.715 9.260 ;
        RECT 70.715 9.095 70.885 9.605 ;
        RECT 67.925 8.610 68.715 8.785 ;
        RECT 66.565 7.310 66.740 8.450 ;
        RECT 67.925 7.310 68.100 8.610 ;
        RECT 68.545 8.570 68.715 8.610 ;
        RECT 68.915 8.455 69.085 8.890 ;
        RECT 70.715 8.765 71.125 9.095 ;
        RECT 70.715 8.565 70.885 8.765 ;
        RECT 71.670 8.565 71.840 9.515 ;
        RECT 68.915 7.310 69.090 8.455 ;
        RECT 70.715 7.305 70.890 8.565 ;
        RECT 71.670 7.305 71.845 8.565 ;
        RECT 72.100 8.445 72.270 10.045 ;
        RECT 82.400 9.935 82.570 10.105 ;
        RECT 82.400 9.605 82.810 9.935 ;
        RECT 82.400 9.095 82.570 9.605 ;
        RECT 82.400 8.765 82.810 9.095 ;
        RECT 82.400 8.565 82.570 8.765 ;
        RECT 72.100 7.305 72.275 8.445 ;
        RECT 74.305 7.560 75.000 8.190 ;
        RECT 22.580 5.980 22.910 6.960 ;
        RECT 24.880 5.980 25.210 6.960 ;
        RECT 26.240 5.980 26.570 6.960 ;
        RECT 27.620 5.980 27.950 6.960 ;
        RECT 39.800 5.980 40.130 6.960 ;
        RECT 42.100 5.980 42.430 6.960 ;
        RECT 43.460 5.980 43.790 6.960 ;
        RECT 44.840 5.980 45.170 6.960 ;
        RECT 57.020 5.985 57.350 6.965 ;
        RECT 59.320 5.985 59.650 6.965 ;
        RECT 60.680 5.985 61.010 6.965 ;
        RECT 62.060 5.985 62.390 6.965 ;
        RECT 74.305 6.960 74.475 7.560 ;
        RECT 74.645 7.340 74.980 7.370 ;
        RECT 75.370 7.340 75.540 8.020 ;
        RECT 74.645 7.170 75.540 7.340 ;
        RECT 76.605 7.560 77.300 8.190 ;
        RECT 77.470 7.560 78.165 8.190 ;
        RECT 78.850 7.560 79.545 8.190 ;
        RECT 74.645 7.120 74.980 7.170 ;
        RECT 76.605 6.960 76.775 7.560 ;
        RECT 76.945 7.340 77.280 7.370 ;
        RECT 77.490 7.340 77.825 7.370 ;
        RECT 76.945 7.170 77.825 7.340 ;
        RECT 76.945 7.120 77.280 7.170 ;
        RECT 77.490 7.120 77.825 7.170 ;
        RECT 77.995 6.960 78.165 7.560 ;
        RECT 78.335 7.120 78.670 7.390 ;
        RECT 78.870 7.120 79.205 7.370 ;
        RECT 79.375 6.960 79.545 7.560 ;
        RECT 79.715 7.120 80.050 7.390 ;
        RECT 82.400 7.305 82.575 8.565 ;
        RECT 82.985 8.535 83.155 10.145 ;
        RECT 83.355 10.085 83.530 10.595 ;
        RECT 83.785 10.045 83.960 10.595 ;
        RECT 85.150 10.085 85.320 10.595 ;
        RECT 86.140 10.085 86.310 10.595 ;
        RECT 87.935 10.105 88.110 10.595 ;
        RECT 82.925 8.365 83.155 8.535 ;
        RECT 83.355 8.565 83.525 9.515 ;
        RECT 82.925 7.305 83.095 8.365 ;
        RECT 83.355 7.305 83.530 8.565 ;
        RECT 83.785 8.445 83.955 10.045 ;
        RECT 87.935 9.935 88.105 10.105 ;
        RECT 88.890 10.085 89.065 10.595 ;
        RECT 89.320 10.045 89.495 10.595 ;
        RECT 99.620 10.105 99.795 10.595 ;
        RECT 100.145 10.315 100.315 10.595 ;
        RECT 100.145 10.145 100.375 10.315 ;
        RECT 84.715 9.425 84.945 9.615 ;
        RECT 87.935 9.605 88.345 9.935 ;
        RECT 84.715 9.385 85.245 9.425 ;
        RECT 84.775 9.255 85.245 9.385 ;
        RECT 85.765 9.255 86.235 9.425 ;
        RECT 84.775 8.565 84.945 9.255 ;
        RECT 85.145 8.780 85.315 8.885 ;
        RECT 85.765 8.780 85.935 9.255 ;
        RECT 87.935 9.095 88.105 9.605 ;
        RECT 85.145 8.605 85.935 8.780 ;
        RECT 83.785 7.305 83.960 8.445 ;
        RECT 85.145 7.305 85.320 8.605 ;
        RECT 85.765 8.565 85.935 8.605 ;
        RECT 86.135 8.450 86.305 8.885 ;
        RECT 87.935 8.765 88.345 9.095 ;
        RECT 87.935 8.565 88.105 8.765 ;
        RECT 88.890 8.565 89.060 9.515 ;
        RECT 86.135 7.305 86.310 8.450 ;
        RECT 87.935 7.305 88.110 8.565 ;
        RECT 88.890 7.305 89.065 8.565 ;
        RECT 89.320 8.445 89.490 10.045 ;
        RECT 99.620 9.935 99.790 10.105 ;
        RECT 99.620 9.605 100.030 9.935 ;
        RECT 99.620 9.095 99.790 9.605 ;
        RECT 99.620 8.765 100.030 9.095 ;
        RECT 99.620 8.565 99.790 8.765 ;
        RECT 89.320 7.305 89.495 8.445 ;
        RECT 91.525 7.560 92.220 8.190 ;
        RECT 91.525 6.960 91.695 7.560 ;
        RECT 91.865 7.340 92.200 7.370 ;
        RECT 92.590 7.340 92.760 8.020 ;
        RECT 91.865 7.170 92.760 7.340 ;
        RECT 93.825 7.560 94.520 8.190 ;
        RECT 94.690 7.560 95.385 8.190 ;
        RECT 96.070 7.560 96.765 8.190 ;
        RECT 91.865 7.120 92.200 7.170 ;
        RECT 93.825 6.960 93.995 7.560 ;
        RECT 94.165 7.340 94.500 7.370 ;
        RECT 94.710 7.340 95.045 7.370 ;
        RECT 94.165 7.170 95.045 7.340 ;
        RECT 94.165 7.120 94.500 7.170 ;
        RECT 94.710 7.120 95.045 7.170 ;
        RECT 95.215 6.960 95.385 7.560 ;
        RECT 95.555 7.120 95.890 7.390 ;
        RECT 96.090 7.120 96.425 7.370 ;
        RECT 96.595 6.960 96.765 7.560 ;
        RECT 96.935 7.120 97.270 7.390 ;
        RECT 99.620 7.305 99.795 8.565 ;
        RECT 100.205 8.535 100.375 10.145 ;
        RECT 100.575 10.085 100.750 10.595 ;
        RECT 101.005 10.045 101.180 10.595 ;
        RECT 102.370 10.085 102.540 10.595 ;
        RECT 103.360 10.085 103.530 10.595 ;
        RECT 100.145 8.365 100.375 8.535 ;
        RECT 100.575 8.565 100.745 9.515 ;
        RECT 100.145 7.305 100.315 8.365 ;
        RECT 100.575 7.305 100.750 8.565 ;
        RECT 101.005 8.445 101.175 10.045 ;
        RECT 101.935 9.425 102.165 9.615 ;
        RECT 101.935 9.385 102.465 9.425 ;
        RECT 101.995 9.255 102.465 9.385 ;
        RECT 102.985 9.255 103.455 9.425 ;
        RECT 101.995 8.565 102.165 9.255 ;
        RECT 102.365 8.780 102.535 8.885 ;
        RECT 102.985 8.780 103.155 9.255 ;
        RECT 102.365 8.605 103.155 8.780 ;
        RECT 101.005 7.305 101.180 8.445 ;
        RECT 102.365 7.305 102.540 8.605 ;
        RECT 102.985 8.565 103.155 8.605 ;
        RECT 103.355 8.450 103.525 8.885 ;
        RECT 103.355 7.305 103.530 8.450 ;
        RECT 74.240 5.980 74.570 6.960 ;
        RECT 76.540 5.980 76.870 6.960 ;
        RECT 77.900 5.980 78.230 6.960 ;
        RECT 79.280 5.980 79.610 6.960 ;
        RECT 91.460 5.980 91.790 6.960 ;
        RECT 93.760 5.980 94.090 6.960 ;
        RECT 95.120 5.980 95.450 6.960 ;
        RECT 96.500 5.980 96.830 6.960 ;
        RECT 22.110 4.490 22.440 5.470 ;
        RECT 23.920 4.670 24.250 5.455 ;
        RECT 23.570 4.500 24.250 4.670 ;
        RECT 24.440 4.670 24.770 5.455 ;
        RECT 24.440 4.500 25.120 4.670 ;
        RECT 22.110 3.890 22.360 4.490 ;
        RECT 22.530 4.280 22.860 4.330 ;
        RECT 23.050 4.280 23.400 4.330 ;
        RECT 22.530 4.110 23.400 4.280 ;
        RECT 22.530 4.080 22.860 4.110 ;
        RECT 23.050 4.080 23.400 4.110 ;
        RECT 23.570 3.900 23.740 4.500 ;
        RECT 23.910 4.080 24.260 4.330 ;
        RECT 24.430 4.080 24.780 4.330 ;
        RECT 24.950 3.900 25.120 4.500 ;
        RECT 25.810 4.620 26.130 5.470 ;
        RECT 26.310 4.960 26.710 5.470 ;
        RECT 27.220 4.960 27.550 5.470 ;
        RECT 26.310 4.790 27.550 4.960 ;
        RECT 28.130 4.620 28.300 5.300 ;
        RECT 28.480 4.790 28.860 5.470 ;
        RECT 25.810 4.540 26.260 4.620 ;
        RECT 25.810 4.370 26.440 4.540 ;
        RECT 25.290 4.080 25.640 4.330 ;
        RECT 22.110 3.260 22.440 3.890 ;
        RECT 23.500 3.260 23.830 3.900 ;
        RECT 24.860 3.260 25.190 3.900 ;
        RECT 26.270 3.490 26.440 4.370 ;
        RECT 27.215 4.450 28.520 4.620 ;
        RECT 26.610 3.830 26.840 4.330 ;
        RECT 27.215 4.250 27.385 4.450 ;
        RECT 27.010 4.080 27.385 4.250 ;
        RECT 27.555 4.080 28.105 4.280 ;
        RECT 28.275 4.000 28.520 4.450 ;
        RECT 28.690 3.830 28.860 4.790 ;
        RECT 26.610 3.660 28.860 3.830 ;
        RECT 30.740 3.895 30.915 5.155 ;
        RECT 31.265 4.095 31.435 5.155 ;
        RECT 31.265 3.925 31.495 4.095 ;
        RECT 30.740 3.695 30.910 3.895 ;
        RECT 26.270 3.320 27.225 3.490 ;
        RECT 28.140 3.340 28.310 3.660 ;
        RECT 30.740 3.365 31.150 3.695 ;
        RECT 30.740 2.855 30.910 3.365 ;
        RECT 30.740 2.525 31.150 2.855 ;
        RECT 30.740 2.355 30.910 2.525 ;
        RECT 30.740 1.865 30.915 2.355 ;
        RECT 31.325 2.315 31.495 3.925 ;
        RECT 31.695 3.895 31.870 5.155 ;
        RECT 32.125 4.015 32.300 5.155 ;
        RECT 31.695 2.945 31.865 3.895 ;
        RECT 32.125 2.415 32.295 4.015 ;
        RECT 33.485 4.010 33.660 5.155 ;
        RECT 39.330 4.490 39.660 5.470 ;
        RECT 41.140 4.670 41.470 5.455 ;
        RECT 40.790 4.500 41.470 4.670 ;
        RECT 41.660 4.670 41.990 5.455 ;
        RECT 41.660 4.500 42.340 4.670 ;
        RECT 33.115 3.205 33.285 3.895 ;
        RECT 33.485 3.805 33.655 4.010 ;
        RECT 34.100 3.805 34.270 3.895 ;
        RECT 33.485 3.625 34.270 3.805 ;
        RECT 33.485 3.575 33.655 3.625 ;
        RECT 34.100 3.205 34.270 3.625 ;
        RECT 39.330 3.890 39.580 4.490 ;
        RECT 39.750 4.280 40.080 4.330 ;
        RECT 40.270 4.280 40.620 4.330 ;
        RECT 39.750 4.110 40.620 4.280 ;
        RECT 39.750 4.080 40.080 4.110 ;
        RECT 40.270 4.080 40.620 4.110 ;
        RECT 40.790 3.900 40.960 4.500 ;
        RECT 41.130 4.080 41.480 4.330 ;
        RECT 41.650 4.080 42.000 4.330 ;
        RECT 42.170 3.900 42.340 4.500 ;
        RECT 43.030 4.620 43.350 5.470 ;
        RECT 43.530 4.960 43.930 5.470 ;
        RECT 44.440 4.960 44.770 5.470 ;
        RECT 43.530 4.790 44.770 4.960 ;
        RECT 45.350 4.620 45.520 5.300 ;
        RECT 45.700 4.790 46.080 5.470 ;
        RECT 43.030 4.540 43.480 4.620 ;
        RECT 43.030 4.370 43.660 4.540 ;
        RECT 42.510 4.080 42.860 4.330 ;
        RECT 39.330 3.260 39.660 3.890 ;
        RECT 40.720 3.260 41.050 3.900 ;
        RECT 42.080 3.260 42.410 3.900 ;
        RECT 43.490 3.490 43.660 4.370 ;
        RECT 44.435 4.450 45.740 4.620 ;
        RECT 43.830 3.830 44.060 4.330 ;
        RECT 44.435 4.250 44.605 4.450 ;
        RECT 44.230 4.080 44.605 4.250 ;
        RECT 44.775 4.080 45.325 4.280 ;
        RECT 45.495 4.000 45.740 4.450 ;
        RECT 45.910 3.830 46.080 4.790 ;
        RECT 43.830 3.660 46.080 3.830 ;
        RECT 47.960 3.895 48.135 5.155 ;
        RECT 48.485 4.095 48.655 5.155 ;
        RECT 48.485 3.925 48.715 4.095 ;
        RECT 47.960 3.695 48.130 3.895 ;
        RECT 43.490 3.320 44.445 3.490 ;
        RECT 45.360 3.340 45.530 3.660 ;
        RECT 47.960 3.365 48.370 3.695 ;
        RECT 33.115 3.175 33.585 3.205 ;
        RECT 33.030 3.035 33.585 3.175 ;
        RECT 34.100 3.035 34.570 3.205 ;
        RECT 33.030 2.945 33.260 3.035 ;
        RECT 47.960 2.855 48.130 3.365 ;
        RECT 47.960 2.525 48.370 2.855 ;
        RECT 31.265 2.145 31.495 2.315 ;
        RECT 31.265 1.865 31.435 2.145 ;
        RECT 31.695 1.865 31.870 2.375 ;
        RECT 32.125 1.865 32.300 2.415 ;
        RECT 33.490 1.865 33.660 2.375 ;
        RECT 47.960 2.355 48.130 2.525 ;
        RECT 47.960 1.865 48.135 2.355 ;
        RECT 48.545 2.315 48.715 3.925 ;
        RECT 48.915 3.895 49.090 5.155 ;
        RECT 49.345 4.015 49.520 5.155 ;
        RECT 48.915 2.945 49.085 3.895 ;
        RECT 49.345 2.415 49.515 4.015 ;
        RECT 50.705 4.010 50.880 5.155 ;
        RECT 56.550 4.495 56.880 5.475 ;
        RECT 58.360 4.675 58.690 5.460 ;
        RECT 58.010 4.505 58.690 4.675 ;
        RECT 58.880 4.675 59.210 5.460 ;
        RECT 58.880 4.505 59.560 4.675 ;
        RECT 50.335 3.205 50.505 3.895 ;
        RECT 50.705 3.805 50.875 4.010 ;
        RECT 56.550 3.895 56.800 4.495 ;
        RECT 56.970 4.285 57.300 4.335 ;
        RECT 57.490 4.285 57.840 4.335 ;
        RECT 56.970 4.115 57.840 4.285 ;
        RECT 56.970 4.085 57.300 4.115 ;
        RECT 57.490 4.085 57.840 4.115 ;
        RECT 58.010 3.905 58.180 4.505 ;
        RECT 58.350 4.085 58.700 4.335 ;
        RECT 58.870 4.085 59.220 4.335 ;
        RECT 59.390 3.905 59.560 4.505 ;
        RECT 60.250 4.625 60.570 5.475 ;
        RECT 60.750 4.965 61.150 5.475 ;
        RECT 61.660 4.965 61.990 5.475 ;
        RECT 60.750 4.795 61.990 4.965 ;
        RECT 62.570 4.625 62.740 5.305 ;
        RECT 62.920 4.795 63.300 5.475 ;
        RECT 60.250 4.545 60.700 4.625 ;
        RECT 60.250 4.375 60.880 4.545 ;
        RECT 59.730 4.085 60.080 4.335 ;
        RECT 51.320 3.805 51.490 3.895 ;
        RECT 50.705 3.625 51.490 3.805 ;
        RECT 50.705 3.575 50.875 3.625 ;
        RECT 51.320 3.205 51.490 3.625 ;
        RECT 56.550 3.265 56.880 3.895 ;
        RECT 57.940 3.265 58.270 3.905 ;
        RECT 59.300 3.265 59.630 3.905 ;
        RECT 60.710 3.495 60.880 4.375 ;
        RECT 61.655 4.455 62.960 4.625 ;
        RECT 61.050 3.835 61.280 4.335 ;
        RECT 61.655 4.255 61.825 4.455 ;
        RECT 61.450 4.085 61.825 4.255 ;
        RECT 61.995 4.085 62.545 4.285 ;
        RECT 62.715 4.005 62.960 4.455 ;
        RECT 63.130 3.835 63.300 4.795 ;
        RECT 61.050 3.665 63.300 3.835 ;
        RECT 65.180 3.900 65.355 5.160 ;
        RECT 65.705 4.100 65.875 5.160 ;
        RECT 65.705 3.930 65.935 4.100 ;
        RECT 65.180 3.700 65.350 3.900 ;
        RECT 60.710 3.325 61.665 3.495 ;
        RECT 62.580 3.345 62.750 3.665 ;
        RECT 65.180 3.370 65.590 3.700 ;
        RECT 50.335 3.175 50.805 3.205 ;
        RECT 50.250 3.035 50.805 3.175 ;
        RECT 51.320 3.035 51.790 3.205 ;
        RECT 50.250 2.945 50.480 3.035 ;
        RECT 65.180 2.860 65.350 3.370 ;
        RECT 65.180 2.530 65.590 2.860 ;
        RECT 48.485 2.145 48.715 2.315 ;
        RECT 48.485 1.865 48.655 2.145 ;
        RECT 48.915 1.865 49.090 2.375 ;
        RECT 49.345 1.865 49.520 2.415 ;
        RECT 50.710 1.865 50.880 2.375 ;
        RECT 65.180 2.360 65.350 2.530 ;
        RECT 65.180 1.870 65.355 2.360 ;
        RECT 65.765 2.320 65.935 3.930 ;
        RECT 66.135 3.900 66.310 5.160 ;
        RECT 66.565 4.020 66.740 5.160 ;
        RECT 66.135 2.950 66.305 3.900 ;
        RECT 66.565 2.420 66.735 4.020 ;
        RECT 67.925 4.015 68.100 5.160 ;
        RECT 73.770 4.490 74.100 5.470 ;
        RECT 75.580 4.670 75.910 5.455 ;
        RECT 75.230 4.500 75.910 4.670 ;
        RECT 76.100 4.670 76.430 5.455 ;
        RECT 76.100 4.500 76.780 4.670 ;
        RECT 67.555 3.210 67.725 3.900 ;
        RECT 67.925 3.810 68.095 4.015 ;
        RECT 68.540 3.810 68.710 3.900 ;
        RECT 67.925 3.630 68.710 3.810 ;
        RECT 67.925 3.580 68.095 3.630 ;
        RECT 68.540 3.210 68.710 3.630 ;
        RECT 73.770 3.890 74.020 4.490 ;
        RECT 74.190 4.280 74.520 4.330 ;
        RECT 74.710 4.280 75.060 4.330 ;
        RECT 74.190 4.110 75.060 4.280 ;
        RECT 74.190 4.080 74.520 4.110 ;
        RECT 74.710 4.080 75.060 4.110 ;
        RECT 75.230 3.900 75.400 4.500 ;
        RECT 75.570 4.080 75.920 4.330 ;
        RECT 76.090 4.080 76.440 4.330 ;
        RECT 76.610 3.900 76.780 4.500 ;
        RECT 77.470 4.620 77.790 5.470 ;
        RECT 77.970 4.960 78.370 5.470 ;
        RECT 78.880 4.960 79.210 5.470 ;
        RECT 77.970 4.790 79.210 4.960 ;
        RECT 79.790 4.620 79.960 5.300 ;
        RECT 80.140 4.790 80.520 5.470 ;
        RECT 77.470 4.540 77.920 4.620 ;
        RECT 77.470 4.370 78.100 4.540 ;
        RECT 76.950 4.080 77.300 4.330 ;
        RECT 73.770 3.260 74.100 3.890 ;
        RECT 75.160 3.260 75.490 3.900 ;
        RECT 76.520 3.260 76.850 3.900 ;
        RECT 77.930 3.490 78.100 4.370 ;
        RECT 78.875 4.450 80.180 4.620 ;
        RECT 78.270 3.830 78.500 4.330 ;
        RECT 78.875 4.250 79.045 4.450 ;
        RECT 78.670 4.080 79.045 4.250 ;
        RECT 79.215 4.080 79.765 4.280 ;
        RECT 79.935 4.000 80.180 4.450 ;
        RECT 80.350 3.830 80.520 4.790 ;
        RECT 78.270 3.660 80.520 3.830 ;
        RECT 82.400 3.895 82.575 5.155 ;
        RECT 82.925 4.095 83.095 5.155 ;
        RECT 82.925 3.925 83.155 4.095 ;
        RECT 82.400 3.695 82.570 3.895 ;
        RECT 77.930 3.320 78.885 3.490 ;
        RECT 79.800 3.340 79.970 3.660 ;
        RECT 82.400 3.365 82.810 3.695 ;
        RECT 67.555 3.180 68.025 3.210 ;
        RECT 67.470 3.040 68.025 3.180 ;
        RECT 68.540 3.040 69.010 3.210 ;
        RECT 67.470 2.950 67.700 3.040 ;
        RECT 82.400 2.855 82.570 3.365 ;
        RECT 82.400 2.525 82.810 2.855 ;
        RECT 65.705 2.150 65.935 2.320 ;
        RECT 65.705 1.870 65.875 2.150 ;
        RECT 66.135 1.870 66.310 2.380 ;
        RECT 66.565 1.870 66.740 2.420 ;
        RECT 67.930 1.870 68.100 2.380 ;
        RECT 82.400 2.355 82.570 2.525 ;
        RECT 82.400 1.865 82.575 2.355 ;
        RECT 82.985 2.315 83.155 3.925 ;
        RECT 83.355 3.895 83.530 5.155 ;
        RECT 83.785 4.015 83.960 5.155 ;
        RECT 83.355 2.945 83.525 3.895 ;
        RECT 83.785 2.415 83.955 4.015 ;
        RECT 85.145 4.010 85.320 5.155 ;
        RECT 90.990 4.490 91.320 5.470 ;
        RECT 92.800 4.670 93.130 5.455 ;
        RECT 92.450 4.500 93.130 4.670 ;
        RECT 93.320 4.670 93.650 5.455 ;
        RECT 93.320 4.500 94.000 4.670 ;
        RECT 84.775 3.205 84.945 3.895 ;
        RECT 85.145 3.805 85.315 4.010 ;
        RECT 85.760 3.805 85.930 3.895 ;
        RECT 85.145 3.625 85.930 3.805 ;
        RECT 85.145 3.575 85.315 3.625 ;
        RECT 85.760 3.205 85.930 3.625 ;
        RECT 90.990 3.890 91.240 4.490 ;
        RECT 91.410 4.280 91.740 4.330 ;
        RECT 91.930 4.280 92.280 4.330 ;
        RECT 91.410 4.110 92.280 4.280 ;
        RECT 91.410 4.080 91.740 4.110 ;
        RECT 91.930 4.080 92.280 4.110 ;
        RECT 92.450 3.900 92.620 4.500 ;
        RECT 92.790 4.080 93.140 4.330 ;
        RECT 93.310 4.080 93.660 4.330 ;
        RECT 93.830 3.900 94.000 4.500 ;
        RECT 94.690 4.620 95.010 5.470 ;
        RECT 95.190 4.960 95.590 5.470 ;
        RECT 96.100 4.960 96.430 5.470 ;
        RECT 95.190 4.790 96.430 4.960 ;
        RECT 97.010 4.620 97.180 5.300 ;
        RECT 97.360 4.790 97.740 5.470 ;
        RECT 94.690 4.540 95.140 4.620 ;
        RECT 94.690 4.370 95.320 4.540 ;
        RECT 94.170 4.080 94.520 4.330 ;
        RECT 90.990 3.260 91.320 3.890 ;
        RECT 92.380 3.260 92.710 3.900 ;
        RECT 93.740 3.260 94.070 3.900 ;
        RECT 95.150 3.490 95.320 4.370 ;
        RECT 96.095 4.450 97.400 4.620 ;
        RECT 95.490 3.830 95.720 4.330 ;
        RECT 96.095 4.250 96.265 4.450 ;
        RECT 95.890 4.080 96.265 4.250 ;
        RECT 96.435 4.080 96.985 4.280 ;
        RECT 97.155 4.000 97.400 4.450 ;
        RECT 97.570 3.830 97.740 4.790 ;
        RECT 95.490 3.660 97.740 3.830 ;
        RECT 99.620 3.895 99.795 5.155 ;
        RECT 100.145 4.095 100.315 5.155 ;
        RECT 100.145 3.925 100.375 4.095 ;
        RECT 99.620 3.695 99.790 3.895 ;
        RECT 95.150 3.320 96.105 3.490 ;
        RECT 97.020 3.340 97.190 3.660 ;
        RECT 99.620 3.365 100.030 3.695 ;
        RECT 84.775 3.175 85.245 3.205 ;
        RECT 84.690 3.035 85.245 3.175 ;
        RECT 85.760 3.035 86.230 3.205 ;
        RECT 84.690 2.945 84.920 3.035 ;
        RECT 99.620 2.855 99.790 3.365 ;
        RECT 99.620 2.525 100.030 2.855 ;
        RECT 82.925 2.145 83.155 2.315 ;
        RECT 82.925 1.865 83.095 2.145 ;
        RECT 83.355 1.865 83.530 2.375 ;
        RECT 83.785 1.865 83.960 2.415 ;
        RECT 85.150 1.865 85.320 2.375 ;
        RECT 99.620 2.355 99.790 2.525 ;
        RECT 99.620 1.865 99.795 2.355 ;
        RECT 100.205 2.315 100.375 3.925 ;
        RECT 100.575 3.895 100.750 5.155 ;
        RECT 101.005 4.015 101.180 5.155 ;
        RECT 100.575 2.945 100.745 3.895 ;
        RECT 101.005 2.415 101.175 4.015 ;
        RECT 102.365 4.010 102.540 5.155 ;
        RECT 101.995 3.205 102.165 3.895 ;
        RECT 102.365 3.805 102.535 4.010 ;
        RECT 102.980 3.805 103.150 3.895 ;
        RECT 102.365 3.625 103.150 3.805 ;
        RECT 102.365 3.575 102.535 3.625 ;
        RECT 102.980 3.205 103.150 3.625 ;
        RECT 101.995 3.175 102.465 3.205 ;
        RECT 101.910 3.035 102.465 3.175 ;
        RECT 102.980 3.035 103.450 3.205 ;
        RECT 101.910 2.945 102.140 3.035 ;
        RECT 100.145 2.145 100.375 2.315 ;
        RECT 100.145 1.865 100.315 2.145 ;
        RECT 100.575 1.865 100.750 2.375 ;
        RECT 101.005 1.865 101.180 2.415 ;
        RECT 102.370 1.865 102.540 2.375 ;
      LAYER met1 ;
        RECT 16.540 10.055 16.830 10.285 ;
        RECT 19.950 10.055 20.240 10.285 ;
        RECT 31.635 10.055 31.925 10.285 ;
        RECT 16.600 9.590 16.770 10.055 ;
        RECT 20.010 9.690 20.180 10.055 ;
        RECT 16.510 9.310 16.850 9.590 ;
        RECT 19.915 9.320 20.285 9.690 ;
        RECT 31.695 9.575 31.865 10.055 ;
        RECT 33.425 10.025 33.720 10.285 ;
        RECT 34.415 10.025 34.710 10.285 ;
        RECT 37.170 10.055 37.460 10.285 ;
        RECT 48.855 10.055 49.145 10.285 ;
        RECT 33.055 9.650 33.285 9.675 ;
        RECT 33.025 9.575 33.315 9.650 ;
        RECT 31.695 9.545 33.315 9.575 ;
        RECT 31.635 9.405 33.315 9.545 ;
        RECT 19.950 9.315 20.240 9.320 ;
        RECT 31.635 9.315 31.925 9.405 ;
        RECT 33.025 9.355 33.315 9.405 ;
        RECT 33.055 9.325 33.285 9.355 ;
        RECT 32.090 9.175 32.415 9.265 ;
        RECT 20.380 9.145 20.670 9.175 ;
        RECT 32.065 9.145 32.415 9.175 ;
        RECT 20.210 9.140 20.670 9.145 ;
        RECT 20.210 8.975 20.700 9.140 ;
        RECT 31.895 8.975 32.415 9.145 ;
        RECT 20.360 8.860 20.700 8.975 ;
        RECT 32.065 8.945 32.415 8.975 ;
        RECT 32.090 8.940 32.415 8.945 ;
        RECT 33.485 8.925 33.655 10.025 ;
        RECT 34.475 9.270 34.645 10.025 ;
        RECT 37.230 9.690 37.400 10.055 ;
        RECT 37.135 9.320 37.505 9.690 ;
        RECT 48.915 9.575 49.085 10.055 ;
        RECT 50.645 10.025 50.940 10.285 ;
        RECT 51.635 10.025 51.930 10.285 ;
        RECT 54.390 10.060 54.680 10.290 ;
        RECT 66.075 10.060 66.365 10.290 ;
        RECT 50.275 9.650 50.505 9.675 ;
        RECT 50.245 9.575 50.535 9.650 ;
        RECT 48.915 9.545 50.535 9.575 ;
        RECT 48.855 9.405 50.535 9.545 ;
        RECT 37.170 9.315 37.460 9.320 ;
        RECT 48.855 9.315 49.145 9.405 ;
        RECT 50.245 9.355 50.535 9.405 ;
        RECT 50.275 9.325 50.505 9.355 ;
        RECT 34.475 8.945 34.805 9.270 ;
        RECT 49.310 9.175 49.635 9.265 ;
        RECT 37.600 9.145 37.890 9.175 ;
        RECT 49.285 9.145 49.635 9.175 ;
        RECT 37.430 9.140 37.890 9.145 ;
        RECT 37.430 8.975 37.920 9.140 ;
        RECT 49.115 8.975 49.635 9.145 ;
        RECT 34.475 8.925 34.765 8.945 ;
        RECT 33.425 8.920 33.655 8.925 ;
        RECT 16.135 8.785 16.475 8.850 ;
        RECT 31.290 8.815 31.610 8.890 ;
        RECT 31.265 8.785 31.610 8.815 ;
        RECT 15.995 8.615 16.475 8.785 ;
        RECT 31.090 8.615 31.610 8.785 ;
        RECT 33.425 8.685 33.715 8.920 ;
        RECT 34.415 8.855 34.765 8.925 ;
        RECT 37.580 8.860 37.920 8.975 ;
        RECT 49.285 8.945 49.635 8.975 ;
        RECT 49.310 8.940 49.635 8.945 ;
        RECT 50.705 8.925 50.875 10.025 ;
        RECT 51.695 9.270 51.865 10.025 ;
        RECT 54.450 9.695 54.620 10.060 ;
        RECT 54.355 9.325 54.725 9.695 ;
        RECT 66.135 9.580 66.305 10.060 ;
        RECT 67.865 10.030 68.160 10.290 ;
        RECT 68.855 10.030 69.150 10.290 ;
        RECT 71.610 10.055 71.900 10.285 ;
        RECT 83.295 10.055 83.585 10.285 ;
        RECT 67.495 9.655 67.725 9.680 ;
        RECT 67.465 9.580 67.755 9.655 ;
        RECT 66.135 9.550 67.755 9.580 ;
        RECT 66.075 9.410 67.755 9.550 ;
        RECT 54.390 9.320 54.680 9.325 ;
        RECT 66.075 9.320 66.365 9.410 ;
        RECT 67.465 9.360 67.755 9.410 ;
        RECT 67.495 9.330 67.725 9.360 ;
        RECT 51.695 8.945 52.025 9.270 ;
        RECT 66.530 9.180 66.855 9.270 ;
        RECT 54.820 9.150 55.110 9.180 ;
        RECT 66.505 9.150 66.855 9.180 ;
        RECT 54.650 9.145 55.110 9.150 ;
        RECT 54.650 8.980 55.140 9.145 ;
        RECT 66.335 8.980 66.855 9.150 ;
        RECT 51.695 8.925 51.985 8.945 ;
        RECT 50.645 8.920 50.875 8.925 ;
        RECT 34.415 8.685 34.705 8.855 ;
        RECT 48.510 8.815 48.830 8.890 ;
        RECT 48.485 8.785 48.830 8.815 ;
        RECT 48.310 8.615 48.830 8.785 ;
        RECT 50.645 8.685 50.935 8.920 ;
        RECT 51.635 8.855 51.985 8.925 ;
        RECT 54.800 8.865 55.140 8.980 ;
        RECT 66.505 8.950 66.855 8.980 ;
        RECT 66.530 8.945 66.855 8.950 ;
        RECT 67.925 8.930 68.095 10.030 ;
        RECT 68.915 9.275 69.085 10.030 ;
        RECT 71.670 9.690 71.840 10.055 ;
        RECT 71.575 9.320 71.945 9.690 ;
        RECT 83.355 9.575 83.525 10.055 ;
        RECT 85.085 10.025 85.380 10.285 ;
        RECT 86.075 10.025 86.370 10.285 ;
        RECT 88.830 10.055 89.120 10.285 ;
        RECT 100.515 10.055 100.805 10.285 ;
        RECT 84.715 9.650 84.945 9.675 ;
        RECT 84.685 9.575 84.975 9.650 ;
        RECT 83.355 9.545 84.975 9.575 ;
        RECT 83.295 9.405 84.975 9.545 ;
        RECT 71.610 9.315 71.900 9.320 ;
        RECT 83.295 9.315 83.585 9.405 ;
        RECT 84.685 9.355 84.975 9.405 ;
        RECT 84.715 9.325 84.945 9.355 ;
        RECT 68.915 8.950 69.245 9.275 ;
        RECT 83.750 9.175 84.075 9.265 ;
        RECT 72.040 9.145 72.330 9.175 ;
        RECT 83.725 9.145 84.075 9.175 ;
        RECT 71.870 9.140 72.330 9.145 ;
        RECT 71.870 8.975 72.360 9.140 ;
        RECT 83.555 8.975 84.075 9.145 ;
        RECT 68.915 8.930 69.205 8.950 ;
        RECT 67.865 8.925 68.095 8.930 ;
        RECT 51.635 8.685 51.925 8.855 ;
        RECT 65.730 8.820 66.050 8.895 ;
        RECT 65.705 8.790 66.050 8.820 ;
        RECT 65.530 8.620 66.050 8.790 ;
        RECT 67.865 8.690 68.155 8.925 ;
        RECT 68.855 8.860 69.205 8.930 ;
        RECT 72.020 8.860 72.360 8.975 ;
        RECT 83.725 8.945 84.075 8.975 ;
        RECT 83.750 8.940 84.075 8.945 ;
        RECT 85.145 8.925 85.315 10.025 ;
        RECT 86.135 9.270 86.305 10.025 ;
        RECT 88.890 9.690 89.060 10.055 ;
        RECT 88.795 9.320 89.165 9.690 ;
        RECT 100.575 9.575 100.745 10.055 ;
        RECT 102.305 10.025 102.600 10.285 ;
        RECT 103.295 10.025 103.590 10.285 ;
        RECT 101.935 9.650 102.165 9.675 ;
        RECT 101.905 9.575 102.195 9.650 ;
        RECT 100.575 9.545 102.195 9.575 ;
        RECT 100.515 9.405 102.195 9.545 ;
        RECT 88.830 9.315 89.120 9.320 ;
        RECT 100.515 9.315 100.805 9.405 ;
        RECT 101.905 9.355 102.195 9.405 ;
        RECT 101.935 9.325 102.165 9.355 ;
        RECT 86.135 8.945 86.465 9.270 ;
        RECT 100.970 9.175 101.295 9.265 ;
        RECT 89.260 9.145 89.550 9.175 ;
        RECT 100.945 9.145 101.295 9.175 ;
        RECT 89.090 9.140 89.550 9.145 ;
        RECT 89.090 8.975 89.580 9.140 ;
        RECT 100.775 8.975 101.295 9.145 ;
        RECT 86.135 8.925 86.425 8.945 ;
        RECT 85.085 8.920 85.315 8.925 ;
        RECT 68.855 8.690 69.145 8.860 ;
        RECT 82.950 8.815 83.270 8.890 ;
        RECT 82.925 8.785 83.270 8.815 ;
        RECT 16.135 8.570 16.475 8.615 ;
        RECT 31.265 8.585 31.610 8.615 ;
        RECT 48.485 8.585 48.830 8.615 ;
        RECT 65.705 8.590 66.050 8.620 ;
        RECT 82.750 8.615 83.270 8.785 ;
        RECT 85.085 8.685 85.375 8.920 ;
        RECT 86.075 8.850 86.425 8.925 ;
        RECT 89.240 8.860 89.580 8.975 ;
        RECT 100.945 8.945 101.295 8.975 ;
        RECT 100.970 8.940 101.295 8.945 ;
        RECT 102.365 8.925 102.535 10.025 ;
        RECT 103.325 10.000 103.590 10.025 ;
        RECT 103.325 9.585 103.650 10.000 ;
        RECT 103.355 8.925 103.525 9.585 ;
        RECT 102.305 8.920 102.535 8.925 ;
        RECT 103.295 8.920 103.525 8.925 ;
        RECT 86.075 8.685 86.365 8.850 ;
        RECT 100.170 8.815 100.490 8.890 ;
        RECT 100.145 8.785 100.490 8.815 ;
        RECT 99.970 8.615 100.490 8.785 ;
        RECT 102.305 8.685 102.595 8.920 ;
        RECT 103.295 8.685 103.585 8.920 ;
        RECT 31.290 8.565 31.610 8.585 ;
        RECT 48.510 8.565 48.830 8.585 ;
        RECT 65.730 8.570 66.050 8.590 ;
        RECT 82.925 8.585 83.270 8.615 ;
        RECT 100.145 8.585 100.490 8.615 ;
        RECT 82.950 8.565 83.270 8.585 ;
        RECT 100.170 8.565 100.490 8.585 ;
        RECT 23.650 8.005 23.940 8.050 ;
        RECT 24.655 8.005 24.975 8.035 ;
        RECT 26.015 8.005 26.335 8.050 ;
        RECT 23.650 7.865 25.565 8.005 ;
        RECT 23.650 7.820 23.940 7.865 ;
        RECT 24.650 7.835 24.980 7.865 ;
        RECT 24.655 7.775 24.975 7.835 ;
        RECT 25.425 7.650 25.565 7.865 ;
        RECT 26.015 7.865 26.610 8.005 ;
        RECT 26.015 7.790 26.335 7.865 ;
        RECT 27.390 7.805 28.035 8.050 ;
        RECT 40.870 8.005 41.160 8.050 ;
        RECT 41.875 8.005 42.195 8.035 ;
        RECT 43.235 8.005 43.555 8.050 ;
        RECT 40.870 7.865 42.785 8.005 ;
        RECT 40.870 7.820 41.160 7.865 ;
        RECT 41.870 7.835 42.200 7.865 ;
        RECT 27.715 7.775 28.035 7.805 ;
        RECT 41.875 7.775 42.195 7.835 ;
        RECT 42.645 7.650 42.785 7.865 ;
        RECT 43.235 7.865 43.830 8.005 ;
        RECT 43.235 7.790 43.555 7.865 ;
        RECT 44.610 7.805 45.255 8.050 ;
        RECT 58.090 8.010 58.380 8.055 ;
        RECT 59.095 8.010 59.415 8.040 ;
        RECT 60.455 8.010 60.775 8.055 ;
        RECT 58.090 7.870 60.005 8.010 ;
        RECT 58.090 7.825 58.380 7.870 ;
        RECT 59.090 7.840 59.420 7.870 ;
        RECT 44.935 7.775 45.255 7.805 ;
        RECT 59.095 7.780 59.415 7.840 ;
        RECT 59.865 7.655 60.005 7.870 ;
        RECT 60.455 7.870 61.050 8.010 ;
        RECT 60.455 7.795 60.775 7.870 ;
        RECT 61.830 7.810 62.475 8.055 ;
        RECT 75.310 8.005 75.600 8.050 ;
        RECT 76.315 8.005 76.635 8.035 ;
        RECT 77.675 8.005 77.995 8.050 ;
        RECT 75.310 7.865 77.225 8.005 ;
        RECT 75.310 7.820 75.600 7.865 ;
        RECT 76.310 7.835 76.640 7.865 ;
        RECT 62.155 7.780 62.475 7.810 ;
        RECT 76.315 7.775 76.635 7.835 ;
        RECT 25.425 7.510 27.435 7.650 ;
        RECT 42.645 7.510 44.655 7.650 ;
        RECT 59.865 7.515 61.875 7.655 ;
        RECT 27.295 7.370 27.435 7.510 ;
        RECT 44.515 7.370 44.655 7.510 ;
        RECT 61.735 7.375 61.875 7.515 ;
        RECT 77.085 7.650 77.225 7.865 ;
        RECT 77.675 7.865 78.270 8.005 ;
        RECT 77.675 7.790 77.995 7.865 ;
        RECT 79.050 7.805 79.695 8.050 ;
        RECT 92.530 8.005 92.820 8.050 ;
        RECT 93.535 8.005 93.855 8.035 ;
        RECT 94.895 8.005 95.215 8.050 ;
        RECT 92.530 7.865 94.445 8.005 ;
        RECT 92.530 7.820 92.820 7.865 ;
        RECT 93.530 7.835 93.860 7.865 ;
        RECT 79.375 7.775 79.695 7.805 ;
        RECT 93.535 7.775 93.855 7.835 ;
        RECT 94.305 7.650 94.445 7.865 ;
        RECT 94.895 7.865 95.490 8.005 ;
        RECT 94.895 7.790 95.215 7.865 ;
        RECT 96.270 7.805 96.915 8.050 ;
        RECT 96.595 7.775 96.915 7.805 ;
        RECT 77.085 7.510 79.095 7.650 ;
        RECT 94.305 7.510 96.315 7.650 ;
        RECT 25.340 7.125 25.985 7.370 ;
        RECT 25.665 7.110 25.985 7.125 ;
        RECT 26.695 7.110 27.015 7.370 ;
        RECT 27.220 7.140 27.510 7.370 ;
        RECT 28.070 7.140 28.360 7.370 ;
        RECT 26.785 6.970 26.925 7.110 ;
        RECT 28.145 6.970 28.285 7.140 ;
        RECT 42.560 7.125 43.205 7.370 ;
        RECT 42.885 7.110 43.205 7.125 ;
        RECT 43.915 7.110 44.235 7.370 ;
        RECT 44.440 7.140 44.730 7.370 ;
        RECT 45.290 7.140 45.580 7.370 ;
        RECT 26.785 6.830 28.285 6.970 ;
        RECT 44.005 6.970 44.145 7.110 ;
        RECT 45.365 6.970 45.505 7.140 ;
        RECT 59.780 7.130 60.425 7.375 ;
        RECT 60.105 7.115 60.425 7.130 ;
        RECT 61.135 7.115 61.455 7.375 ;
        RECT 61.660 7.145 61.950 7.375 ;
        RECT 62.510 7.145 62.800 7.375 ;
        RECT 78.955 7.370 79.095 7.510 ;
        RECT 96.175 7.370 96.315 7.510 ;
        RECT 44.005 6.830 45.505 6.970 ;
        RECT 61.225 6.975 61.365 7.115 ;
        RECT 62.585 6.975 62.725 7.145 ;
        RECT 77.000 7.125 77.645 7.370 ;
        RECT 77.325 7.110 77.645 7.125 ;
        RECT 78.355 7.110 78.675 7.370 ;
        RECT 78.880 7.140 79.170 7.370 ;
        RECT 79.730 7.140 80.020 7.370 ;
        RECT 61.225 6.835 62.725 6.975 ;
        RECT 78.445 6.970 78.585 7.110 ;
        RECT 79.805 6.970 79.945 7.140 ;
        RECT 94.220 7.125 94.865 7.370 ;
        RECT 94.545 7.110 94.865 7.125 ;
        RECT 95.575 7.110 95.895 7.370 ;
        RECT 96.100 7.140 96.390 7.370 ;
        RECT 96.950 7.140 97.240 7.370 ;
        RECT 78.445 6.830 79.945 6.970 ;
        RECT 95.665 6.970 95.805 7.110 ;
        RECT 97.025 6.970 97.165 7.140 ;
        RECT 95.665 6.830 97.165 6.970 ;
        RECT 22.615 6.305 22.935 6.365 ;
        RECT 22.340 6.165 22.935 6.305 ;
        RECT 22.615 6.105 22.935 6.165 ;
        RECT 24.890 6.305 25.180 6.350 ;
        RECT 27.035 6.305 27.355 6.365 ;
        RECT 39.835 6.305 40.155 6.365 ;
        RECT 24.890 6.165 27.355 6.305 ;
        RECT 39.560 6.165 40.155 6.305 ;
        RECT 24.890 6.120 25.180 6.165 ;
        RECT 27.035 6.105 27.355 6.165 ;
        RECT 39.835 6.105 40.155 6.165 ;
        RECT 42.110 6.305 42.400 6.350 ;
        RECT 44.255 6.305 44.575 6.365 ;
        RECT 57.055 6.310 57.375 6.370 ;
        RECT 42.110 6.165 44.575 6.305 ;
        RECT 56.780 6.170 57.375 6.310 ;
        RECT 42.110 6.120 42.400 6.165 ;
        RECT 44.255 6.105 44.575 6.165 ;
        RECT 57.055 6.110 57.375 6.170 ;
        RECT 59.330 6.310 59.620 6.355 ;
        RECT 61.475 6.310 61.795 6.370 ;
        RECT 59.330 6.170 61.795 6.310 ;
        RECT 74.275 6.305 74.595 6.365 ;
        RECT 59.330 6.125 59.620 6.170 ;
        RECT 61.475 6.110 61.795 6.170 ;
        RECT 74.000 6.165 74.595 6.305 ;
        RECT 74.275 6.105 74.595 6.165 ;
        RECT 76.550 6.305 76.840 6.350 ;
        RECT 78.695 6.305 79.015 6.365 ;
        RECT 91.495 6.305 91.815 6.365 ;
        RECT 76.550 6.165 79.015 6.305 ;
        RECT 91.220 6.165 91.815 6.305 ;
        RECT 76.550 6.120 76.840 6.165 ;
        RECT 78.695 6.105 79.015 6.165 ;
        RECT 91.495 6.105 91.815 6.165 ;
        RECT 93.770 6.305 94.060 6.350 ;
        RECT 95.915 6.305 96.235 6.365 ;
        RECT 93.770 6.165 96.235 6.305 ;
        RECT 93.770 6.120 94.060 6.165 ;
        RECT 95.915 6.105 96.235 6.165 ;
        RECT 23.990 5.285 24.280 5.330 ;
        RECT 26.355 5.285 26.675 5.345 ;
        RECT 23.990 5.145 26.675 5.285 ;
        RECT 23.990 5.100 24.280 5.145 ;
        RECT 26.355 5.085 26.675 5.145 ;
        RECT 27.035 5.285 27.355 5.345 ;
        RECT 28.070 5.285 28.360 5.330 ;
        RECT 27.035 5.145 28.360 5.285 ;
        RECT 27.035 5.085 27.355 5.145 ;
        RECT 28.070 5.100 28.360 5.145 ;
        RECT 41.210 5.285 41.500 5.330 ;
        RECT 43.575 5.285 43.895 5.345 ;
        RECT 41.210 5.145 43.895 5.285 ;
        RECT 41.210 5.100 41.500 5.145 ;
        RECT 43.575 5.085 43.895 5.145 ;
        RECT 44.255 5.285 44.575 5.345 ;
        RECT 45.290 5.285 45.580 5.330 ;
        RECT 44.255 5.145 45.580 5.285 ;
        RECT 44.255 5.085 44.575 5.145 ;
        RECT 45.290 5.100 45.580 5.145 ;
        RECT 58.430 5.290 58.720 5.335 ;
        RECT 60.795 5.290 61.115 5.350 ;
        RECT 58.430 5.150 61.115 5.290 ;
        RECT 58.430 5.105 58.720 5.150 ;
        RECT 60.795 5.090 61.115 5.150 ;
        RECT 61.475 5.290 61.795 5.350 ;
        RECT 62.510 5.290 62.800 5.335 ;
        RECT 61.475 5.150 62.800 5.290 ;
        RECT 61.475 5.090 61.795 5.150 ;
        RECT 62.510 5.105 62.800 5.150 ;
        RECT 75.650 5.285 75.940 5.330 ;
        RECT 78.015 5.285 78.335 5.345 ;
        RECT 75.650 5.145 78.335 5.285 ;
        RECT 75.650 5.100 75.940 5.145 ;
        RECT 78.015 5.085 78.335 5.145 ;
        RECT 78.695 5.285 79.015 5.345 ;
        RECT 79.730 5.285 80.020 5.330 ;
        RECT 78.695 5.145 80.020 5.285 ;
        RECT 78.695 5.085 79.015 5.145 ;
        RECT 79.730 5.100 80.020 5.145 ;
        RECT 92.870 5.285 93.160 5.330 ;
        RECT 95.235 5.285 95.555 5.345 ;
        RECT 92.870 5.145 95.555 5.285 ;
        RECT 92.870 5.100 93.160 5.145 ;
        RECT 95.235 5.085 95.555 5.145 ;
        RECT 95.915 5.285 96.235 5.345 ;
        RECT 96.950 5.285 97.240 5.330 ;
        RECT 95.915 5.145 97.240 5.285 ;
        RECT 95.915 5.085 96.235 5.145 ;
        RECT 96.950 5.100 97.240 5.145 ;
        RECT 22.120 4.945 22.410 4.990 ;
        RECT 24.995 4.945 25.315 5.005 ;
        RECT 22.120 4.805 25.315 4.945 ;
        RECT 22.120 4.760 22.410 4.805 ;
        RECT 22.615 4.265 22.935 4.325 ;
        RECT 24.575 4.315 24.715 4.805 ;
        RECT 24.995 4.745 25.315 4.805 ;
        RECT 39.340 4.945 39.630 4.990 ;
        RECT 42.215 4.945 42.535 5.005 ;
        RECT 39.340 4.805 42.535 4.945 ;
        RECT 39.340 4.760 39.630 4.805 ;
        RECT 26.015 4.605 26.335 4.665 ;
        RECT 25.740 4.465 26.335 4.605 ;
        RECT 26.015 4.405 26.335 4.465 ;
        RECT 23.990 4.270 24.280 4.315 ;
        RECT 22.340 4.125 22.935 4.265 ;
        RECT 22.615 4.065 22.935 4.125 ;
        RECT 23.385 4.130 24.280 4.270 ;
        RECT 23.385 3.985 23.525 4.130 ;
        RECT 23.990 4.085 24.280 4.130 ;
        RECT 24.500 4.085 24.790 4.315 ;
        RECT 25.335 4.265 25.655 4.325 ;
        RECT 27.715 4.265 28.035 4.325 ;
        RECT 39.835 4.265 40.155 4.325 ;
        RECT 41.795 4.315 41.935 4.805 ;
        RECT 42.215 4.745 42.535 4.805 ;
        RECT 56.560 4.950 56.850 4.995 ;
        RECT 59.435 4.950 59.755 5.010 ;
        RECT 56.560 4.810 59.755 4.950 ;
        RECT 56.560 4.765 56.850 4.810 ;
        RECT 43.235 4.605 43.555 4.665 ;
        RECT 42.960 4.465 43.555 4.605 ;
        RECT 43.235 4.405 43.555 4.465 ;
        RECT 41.210 4.270 41.500 4.315 ;
        RECT 25.060 4.125 25.655 4.265 ;
        RECT 27.440 4.125 28.035 4.265 ;
        RECT 39.560 4.125 40.155 4.265 ;
        RECT 25.335 4.065 25.655 4.125 ;
        RECT 27.715 4.065 28.035 4.125 ;
        RECT 39.835 4.065 40.155 4.125 ;
        RECT 40.605 4.130 41.500 4.270 ;
        RECT 40.605 3.985 40.745 4.130 ;
        RECT 41.210 4.085 41.500 4.130 ;
        RECT 41.720 4.085 42.010 4.315 ;
        RECT 42.555 4.265 42.875 4.325 ;
        RECT 44.935 4.265 45.255 4.325 ;
        RECT 57.055 4.270 57.375 4.330 ;
        RECT 59.015 4.320 59.155 4.810 ;
        RECT 59.435 4.750 59.755 4.810 ;
        RECT 73.780 4.945 74.070 4.990 ;
        RECT 76.655 4.945 76.975 5.005 ;
        RECT 73.780 4.805 76.975 4.945 ;
        RECT 73.780 4.760 74.070 4.805 ;
        RECT 60.455 4.610 60.775 4.670 ;
        RECT 60.180 4.470 60.775 4.610 ;
        RECT 60.455 4.410 60.775 4.470 ;
        RECT 58.430 4.275 58.720 4.320 ;
        RECT 42.280 4.125 42.875 4.265 ;
        RECT 44.660 4.125 45.255 4.265 ;
        RECT 56.780 4.130 57.375 4.270 ;
        RECT 42.555 4.065 42.875 4.125 ;
        RECT 44.935 4.065 45.255 4.125 ;
        RECT 57.055 4.070 57.375 4.130 ;
        RECT 57.825 4.135 58.720 4.275 ;
        RECT 57.825 3.990 57.965 4.135 ;
        RECT 58.430 4.090 58.720 4.135 ;
        RECT 58.940 4.090 59.230 4.320 ;
        RECT 59.775 4.270 60.095 4.330 ;
        RECT 62.155 4.270 62.475 4.330 ;
        RECT 59.500 4.130 60.095 4.270 ;
        RECT 61.880 4.130 62.475 4.270 ;
        RECT 74.275 4.265 74.595 4.325 ;
        RECT 76.235 4.315 76.375 4.805 ;
        RECT 76.655 4.745 76.975 4.805 ;
        RECT 91.000 4.945 91.290 4.990 ;
        RECT 93.875 4.945 94.195 5.005 ;
        RECT 91.000 4.805 94.195 4.945 ;
        RECT 91.000 4.760 91.290 4.805 ;
        RECT 77.675 4.605 77.995 4.665 ;
        RECT 77.400 4.465 77.995 4.605 ;
        RECT 77.675 4.405 77.995 4.465 ;
        RECT 75.650 4.270 75.940 4.315 ;
        RECT 59.775 4.070 60.095 4.130 ;
        RECT 62.155 4.070 62.475 4.130 ;
        RECT 74.000 4.125 74.595 4.265 ;
        RECT 74.275 4.065 74.595 4.125 ;
        RECT 75.045 4.130 75.940 4.270 ;
        RECT 23.295 3.725 23.615 3.985 ;
        RECT 31.290 3.875 31.610 3.980 ;
        RECT 31.265 3.860 31.610 3.875 ;
        RECT 24.655 3.800 24.975 3.815 ;
        RECT 24.655 3.755 25.160 3.800 ;
        RECT 24.565 3.615 25.160 3.755 ;
        RECT 30.975 3.690 31.610 3.860 ;
        RECT 31.090 3.675 31.610 3.690 ;
        RECT 31.265 3.660 31.610 3.675 ;
        RECT 31.265 3.645 31.555 3.660 ;
        RECT 24.655 3.570 25.160 3.615 ;
        RECT 24.655 3.555 24.975 3.570 ;
        RECT 29.620 3.290 29.945 3.615 ;
        RECT 32.065 3.485 32.415 3.610 ;
        RECT 33.425 3.540 33.715 3.775 ;
        RECT 40.515 3.725 40.835 3.985 ;
        RECT 48.510 3.875 48.830 3.980 ;
        RECT 48.485 3.860 48.830 3.875 ;
        RECT 41.875 3.800 42.195 3.815 ;
        RECT 41.875 3.755 42.380 3.800 ;
        RECT 41.785 3.615 42.380 3.755 ;
        RECT 48.195 3.690 48.830 3.860 ;
        RECT 48.310 3.675 48.830 3.690 ;
        RECT 48.485 3.660 48.830 3.675 ;
        RECT 48.485 3.645 48.775 3.660 ;
        RECT 41.875 3.570 42.380 3.615 ;
        RECT 41.875 3.555 42.195 3.570 ;
        RECT 33.425 3.535 33.655 3.540 ;
        RECT 31.895 3.315 32.415 3.485 ;
        RECT 32.065 3.260 32.415 3.315 ;
        RECT 33.030 3.205 33.260 3.235 ;
        RECT 31.635 3.120 31.925 3.145 ;
        RECT 33.000 3.120 33.290 3.205 ;
        RECT 31.635 2.950 33.290 3.120 ;
        RECT 31.635 2.915 31.925 2.950 ;
        RECT 31.695 2.405 31.865 2.915 ;
        RECT 33.000 2.910 33.290 2.950 ;
        RECT 33.030 2.885 33.260 2.910 ;
        RECT 33.485 2.435 33.655 3.535 ;
        RECT 46.840 3.290 47.165 3.615 ;
        RECT 49.285 3.485 49.635 3.610 ;
        RECT 50.645 3.540 50.935 3.775 ;
        RECT 57.735 3.730 58.055 3.990 ;
        RECT 75.045 3.985 75.185 4.130 ;
        RECT 75.650 4.085 75.940 4.130 ;
        RECT 76.160 4.085 76.450 4.315 ;
        RECT 76.995 4.265 77.315 4.325 ;
        RECT 79.375 4.265 79.695 4.325 ;
        RECT 91.495 4.265 91.815 4.325 ;
        RECT 93.455 4.315 93.595 4.805 ;
        RECT 93.875 4.745 94.195 4.805 ;
        RECT 94.895 4.605 95.215 4.665 ;
        RECT 94.620 4.465 95.215 4.605 ;
        RECT 94.895 4.405 95.215 4.465 ;
        RECT 92.870 4.270 93.160 4.315 ;
        RECT 76.720 4.125 77.315 4.265 ;
        RECT 79.100 4.125 79.695 4.265 ;
        RECT 91.220 4.125 91.815 4.265 ;
        RECT 76.995 4.065 77.315 4.125 ;
        RECT 79.375 4.065 79.695 4.125 ;
        RECT 91.495 4.065 91.815 4.125 ;
        RECT 92.265 4.130 93.160 4.270 ;
        RECT 92.265 3.985 92.405 4.130 ;
        RECT 92.870 4.085 93.160 4.130 ;
        RECT 93.380 4.085 93.670 4.315 ;
        RECT 94.215 4.265 94.535 4.325 ;
        RECT 96.595 4.265 96.915 4.325 ;
        RECT 93.940 4.125 94.535 4.265 ;
        RECT 96.320 4.125 96.915 4.265 ;
        RECT 94.215 4.065 94.535 4.125 ;
        RECT 96.595 4.065 96.915 4.125 ;
        RECT 65.730 3.880 66.050 3.985 ;
        RECT 65.705 3.865 66.050 3.880 ;
        RECT 59.095 3.805 59.415 3.820 ;
        RECT 59.095 3.760 59.600 3.805 ;
        RECT 59.005 3.620 59.600 3.760 ;
        RECT 65.415 3.695 66.050 3.865 ;
        RECT 65.530 3.680 66.050 3.695 ;
        RECT 65.705 3.665 66.050 3.680 ;
        RECT 65.705 3.650 65.995 3.665 ;
        RECT 59.095 3.575 59.600 3.620 ;
        RECT 59.095 3.560 59.415 3.575 ;
        RECT 50.645 3.535 50.875 3.540 ;
        RECT 49.115 3.315 49.635 3.485 ;
        RECT 49.285 3.260 49.635 3.315 ;
        RECT 50.250 3.205 50.480 3.235 ;
        RECT 48.855 3.120 49.145 3.145 ;
        RECT 50.220 3.120 50.510 3.205 ;
        RECT 48.855 2.950 50.510 3.120 ;
        RECT 48.855 2.915 49.145 2.950 ;
        RECT 31.635 2.175 31.925 2.405 ;
        RECT 33.425 2.175 33.720 2.435 ;
        RECT 48.915 2.405 49.085 2.915 ;
        RECT 50.220 2.910 50.510 2.950 ;
        RECT 50.250 2.885 50.480 2.910 ;
        RECT 50.705 2.435 50.875 3.535 ;
        RECT 64.060 3.295 64.385 3.620 ;
        RECT 66.505 3.490 66.855 3.615 ;
        RECT 67.865 3.545 68.155 3.780 ;
        RECT 74.955 3.725 75.275 3.985 ;
        RECT 82.950 3.875 83.270 3.980 ;
        RECT 82.925 3.860 83.270 3.875 ;
        RECT 76.315 3.800 76.635 3.815 ;
        RECT 76.315 3.755 76.820 3.800 ;
        RECT 76.225 3.615 76.820 3.755 ;
        RECT 82.635 3.690 83.270 3.860 ;
        RECT 82.750 3.675 83.270 3.690 ;
        RECT 82.925 3.660 83.270 3.675 ;
        RECT 82.925 3.645 83.215 3.660 ;
        RECT 76.315 3.570 76.820 3.615 ;
        RECT 76.315 3.555 76.635 3.570 ;
        RECT 67.865 3.540 68.095 3.545 ;
        RECT 66.335 3.320 66.855 3.490 ;
        RECT 66.505 3.265 66.855 3.320 ;
        RECT 67.470 3.210 67.700 3.240 ;
        RECT 66.075 3.125 66.365 3.150 ;
        RECT 67.440 3.125 67.730 3.210 ;
        RECT 66.075 2.955 67.730 3.125 ;
        RECT 66.075 2.920 66.365 2.955 ;
        RECT 48.855 2.175 49.145 2.405 ;
        RECT 50.645 2.175 50.940 2.435 ;
        RECT 66.135 2.410 66.305 2.920 ;
        RECT 67.440 2.915 67.730 2.955 ;
        RECT 67.470 2.890 67.700 2.915 ;
        RECT 67.925 2.440 68.095 3.540 ;
        RECT 81.280 3.290 81.605 3.615 ;
        RECT 83.725 3.485 84.075 3.610 ;
        RECT 85.085 3.540 85.375 3.775 ;
        RECT 92.175 3.725 92.495 3.985 ;
        RECT 100.170 3.875 100.490 3.980 ;
        RECT 100.145 3.860 100.490 3.875 ;
        RECT 93.535 3.800 93.855 3.815 ;
        RECT 93.535 3.755 94.040 3.800 ;
        RECT 93.445 3.615 94.040 3.755 ;
        RECT 99.855 3.690 100.490 3.860 ;
        RECT 99.970 3.675 100.490 3.690 ;
        RECT 100.145 3.660 100.490 3.675 ;
        RECT 100.145 3.645 100.435 3.660 ;
        RECT 93.535 3.570 94.040 3.615 ;
        RECT 93.535 3.555 93.855 3.570 ;
        RECT 85.085 3.535 85.315 3.540 ;
        RECT 83.555 3.315 84.075 3.485 ;
        RECT 83.725 3.260 84.075 3.315 ;
        RECT 84.690 3.205 84.920 3.235 ;
        RECT 83.295 3.120 83.585 3.145 ;
        RECT 84.660 3.120 84.950 3.205 ;
        RECT 83.295 2.950 84.950 3.120 ;
        RECT 83.295 2.915 83.585 2.950 ;
        RECT 66.075 2.180 66.365 2.410 ;
        RECT 67.865 2.180 68.160 2.440 ;
        RECT 83.355 2.405 83.525 2.915 ;
        RECT 84.660 2.910 84.950 2.950 ;
        RECT 84.690 2.885 84.920 2.910 ;
        RECT 85.145 2.435 85.315 3.535 ;
        RECT 98.500 3.290 98.825 3.615 ;
        RECT 100.945 3.485 101.295 3.610 ;
        RECT 102.305 3.540 102.595 3.775 ;
        RECT 102.305 3.535 102.535 3.540 ;
        RECT 100.775 3.315 101.295 3.485 ;
        RECT 100.945 3.260 101.295 3.315 ;
        RECT 101.910 3.205 102.140 3.235 ;
        RECT 100.515 3.120 100.805 3.145 ;
        RECT 101.880 3.120 102.170 3.205 ;
        RECT 100.515 2.950 102.170 3.120 ;
        RECT 100.515 2.915 100.805 2.950 ;
        RECT 83.295 2.175 83.585 2.405 ;
        RECT 85.085 2.175 85.380 2.435 ;
        RECT 100.575 2.405 100.745 2.915 ;
        RECT 101.880 2.910 102.170 2.950 ;
        RECT 101.910 2.885 102.140 2.910 ;
        RECT 102.365 2.435 102.535 3.535 ;
        RECT 100.515 2.175 100.805 2.405 ;
        RECT 102.305 2.175 102.600 2.435 ;
      LAYER met2 ;
        RECT 16.210 10.055 103.530 10.225 ;
        RECT 16.210 8.880 16.380 10.055 ;
        RECT 103.360 9.910 103.530 10.055 ;
        RECT 16.540 9.515 16.820 9.620 ;
        RECT 16.540 9.345 17.745 9.515 ;
        RECT 16.540 9.280 16.820 9.345 ;
        RECT 17.575 9.140 17.745 9.345 ;
        RECT 19.915 9.320 20.285 9.690 ;
        RECT 20.440 9.550 31.135 9.720 ;
        RECT 20.440 9.170 20.610 9.550 ;
        RECT 30.975 9.200 31.135 9.550 ;
        RECT 37.135 9.320 37.505 9.690 ;
        RECT 37.660 9.550 48.355 9.720 ;
        RECT 32.090 9.200 32.415 9.265 ;
        RECT 20.390 9.140 20.670 9.170 ;
        RECT 17.575 8.970 20.670 9.140 ;
        RECT 16.165 8.540 16.445 8.880 ;
        RECT 20.390 8.830 20.670 8.970 ;
        RECT 30.975 9.030 32.415 9.200 ;
        RECT 24.675 7.725 24.955 8.095 ;
        RECT 26.045 8.050 26.305 8.095 ;
        RECT 26.015 7.805 26.335 8.050 ;
        RECT 26.045 7.760 26.305 7.805 ;
        RECT 27.745 7.760 28.005 8.095 ;
        RECT 25.685 7.065 25.965 7.435 ;
        RECT 26.105 6.645 26.245 7.760 ;
        RECT 26.725 7.065 27.005 7.435 ;
        RECT 25.425 6.505 26.245 6.645 ;
        RECT 22.645 6.075 22.905 6.395 ;
        RECT 22.705 4.355 22.845 6.075 ;
        RECT 25.425 5.800 25.565 6.505 ;
        RECT 27.065 6.075 27.325 6.395 ;
        RECT 23.315 5.430 23.595 5.800 ;
        RECT 25.355 5.430 25.635 5.800 ;
        RECT 22.645 4.035 22.905 4.355 ;
        RECT 23.385 4.015 23.525 5.430 ;
        RECT 25.005 4.690 25.285 5.060 ;
        RECT 25.425 4.355 25.565 5.430 ;
        RECT 26.375 5.030 26.655 5.400 ;
        RECT 27.125 5.375 27.265 6.075 ;
        RECT 27.065 5.055 27.325 5.375 ;
        RECT 25.365 4.035 25.625 4.355 ;
        RECT 26.035 4.350 26.315 4.720 ;
        RECT 27.805 4.355 27.945 7.760 ;
        RECT 27.745 4.035 28.005 4.355 ;
        RECT 23.325 3.695 23.585 4.015 ;
        RECT 24.675 3.815 24.955 3.870 ;
        RECT 30.975 3.860 31.135 9.030 ;
        RECT 32.090 8.940 32.415 9.030 ;
        RECT 34.480 9.145 34.805 9.270 ;
        RECT 37.660 9.170 37.830 9.550 ;
        RECT 48.195 9.200 48.355 9.550 ;
        RECT 54.355 9.325 54.725 9.695 ;
        RECT 54.880 9.555 65.575 9.725 ;
        RECT 49.310 9.200 49.635 9.265 ;
        RECT 34.480 9.140 35.715 9.145 ;
        RECT 37.610 9.140 37.890 9.170 ;
        RECT 34.480 8.975 37.890 9.140 ;
        RECT 34.480 8.945 34.805 8.975 ;
        RECT 35.715 8.970 37.890 8.975 ;
        RECT 31.290 8.565 31.610 8.890 ;
        RECT 37.610 8.830 37.890 8.970 ;
        RECT 48.195 9.030 49.635 9.200 ;
        RECT 31.320 8.330 31.490 8.565 ;
        RECT 31.320 8.155 31.495 8.330 ;
        RECT 31.320 7.980 32.295 8.155 ;
        RECT 31.290 3.860 31.610 3.980 ;
        RECT 24.675 3.640 29.325 3.815 ;
        RECT 30.975 3.690 31.610 3.860 ;
        RECT 31.290 3.660 31.610 3.690 ;
        RECT 24.675 3.500 24.955 3.640 ;
        RECT 29.150 3.490 29.325 3.640 ;
        RECT 29.620 3.490 29.945 3.615 ;
        RECT 32.120 3.610 32.295 7.980 ;
        RECT 41.895 7.725 42.175 8.095 ;
        RECT 43.265 8.050 43.525 8.095 ;
        RECT 43.235 7.805 43.555 8.050 ;
        RECT 43.265 7.760 43.525 7.805 ;
        RECT 44.965 7.760 45.225 8.095 ;
        RECT 42.905 7.065 43.185 7.435 ;
        RECT 43.325 6.645 43.465 7.760 ;
        RECT 43.945 7.065 44.225 7.435 ;
        RECT 42.645 6.505 43.465 6.645 ;
        RECT 39.865 6.075 40.125 6.395 ;
        RECT 39.925 4.355 40.065 6.075 ;
        RECT 42.645 5.800 42.785 6.505 ;
        RECT 44.285 6.075 44.545 6.395 ;
        RECT 40.535 5.430 40.815 5.800 ;
        RECT 42.575 5.430 42.855 5.800 ;
        RECT 39.865 4.035 40.125 4.355 ;
        RECT 40.605 4.015 40.745 5.430 ;
        RECT 42.225 4.690 42.505 5.060 ;
        RECT 42.645 4.355 42.785 5.430 ;
        RECT 43.595 5.030 43.875 5.400 ;
        RECT 44.345 5.375 44.485 6.075 ;
        RECT 44.285 5.055 44.545 5.375 ;
        RECT 42.585 4.035 42.845 4.355 ;
        RECT 43.255 4.350 43.535 4.720 ;
        RECT 45.025 4.355 45.165 7.760 ;
        RECT 44.965 4.035 45.225 4.355 ;
        RECT 40.545 3.695 40.805 4.015 ;
        RECT 41.895 3.815 42.175 3.870 ;
        RECT 48.195 3.860 48.355 9.030 ;
        RECT 49.310 8.940 49.635 9.030 ;
        RECT 51.700 9.145 52.025 9.270 ;
        RECT 54.880 9.175 55.050 9.555 ;
        RECT 65.415 9.205 65.575 9.555 ;
        RECT 71.575 9.320 71.945 9.690 ;
        RECT 72.100 9.550 82.795 9.720 ;
        RECT 66.530 9.205 66.855 9.270 ;
        RECT 51.700 9.140 52.885 9.145 ;
        RECT 54.830 9.140 55.110 9.175 ;
        RECT 51.700 8.975 55.120 9.140 ;
        RECT 51.700 8.945 52.025 8.975 ;
        RECT 52.885 8.970 55.120 8.975 ;
        RECT 65.415 9.035 66.855 9.205 ;
        RECT 48.510 8.565 48.830 8.890 ;
        RECT 54.830 8.835 55.110 8.970 ;
        RECT 48.540 8.330 48.710 8.565 ;
        RECT 48.540 8.155 48.715 8.330 ;
        RECT 48.540 7.980 49.515 8.155 ;
        RECT 48.510 3.860 48.830 3.980 ;
        RECT 41.895 3.640 46.545 3.815 ;
        RECT 48.195 3.690 48.830 3.860 ;
        RECT 48.510 3.660 48.830 3.690 ;
        RECT 32.065 3.490 32.415 3.610 ;
        RECT 41.895 3.500 42.175 3.640 ;
        RECT 29.150 3.320 32.415 3.490 ;
        RECT 46.370 3.490 46.545 3.640 ;
        RECT 46.840 3.490 47.165 3.615 ;
        RECT 49.340 3.610 49.515 7.980 ;
        RECT 59.115 7.730 59.395 8.100 ;
        RECT 60.485 8.055 60.745 8.100 ;
        RECT 60.455 7.810 60.775 8.055 ;
        RECT 60.485 7.765 60.745 7.810 ;
        RECT 62.185 7.765 62.445 8.100 ;
        RECT 60.125 7.070 60.405 7.440 ;
        RECT 60.545 6.650 60.685 7.765 ;
        RECT 61.165 7.070 61.445 7.440 ;
        RECT 59.865 6.510 60.685 6.650 ;
        RECT 57.085 6.080 57.345 6.400 ;
        RECT 57.145 4.360 57.285 6.080 ;
        RECT 59.865 5.805 60.005 6.510 ;
        RECT 61.505 6.080 61.765 6.400 ;
        RECT 57.755 5.435 58.035 5.805 ;
        RECT 59.795 5.435 60.075 5.805 ;
        RECT 57.085 4.040 57.345 4.360 ;
        RECT 57.825 4.020 57.965 5.435 ;
        RECT 59.445 4.695 59.725 5.065 ;
        RECT 59.865 4.360 60.005 5.435 ;
        RECT 60.815 5.035 61.095 5.405 ;
        RECT 61.565 5.380 61.705 6.080 ;
        RECT 61.505 5.060 61.765 5.380 ;
        RECT 59.805 4.040 60.065 4.360 ;
        RECT 60.475 4.355 60.755 4.725 ;
        RECT 62.245 4.360 62.385 7.765 ;
        RECT 62.185 4.040 62.445 4.360 ;
        RECT 57.765 3.700 58.025 4.020 ;
        RECT 59.115 3.820 59.395 3.875 ;
        RECT 65.415 3.865 65.575 9.035 ;
        RECT 66.530 8.945 66.855 9.035 ;
        RECT 68.920 9.150 69.245 9.275 ;
        RECT 72.100 9.170 72.270 9.550 ;
        RECT 82.635 9.200 82.795 9.550 ;
        RECT 88.795 9.320 89.165 9.690 ;
        RECT 89.320 9.550 100.015 9.720 ;
        RECT 103.325 9.585 103.650 9.910 ;
        RECT 83.750 9.200 84.075 9.265 ;
        RECT 68.920 9.145 69.970 9.150 ;
        RECT 68.920 9.140 70.045 9.145 ;
        RECT 72.050 9.140 72.330 9.170 ;
        RECT 68.920 8.980 72.330 9.140 ;
        RECT 68.920 8.950 69.245 8.980 ;
        RECT 69.970 8.975 72.330 8.980 ;
        RECT 70.045 8.970 72.330 8.975 ;
        RECT 65.730 8.570 66.050 8.895 ;
        RECT 72.050 8.830 72.330 8.970 ;
        RECT 82.635 9.030 84.075 9.200 ;
        RECT 65.760 8.335 65.930 8.570 ;
        RECT 65.760 8.160 65.935 8.335 ;
        RECT 65.760 7.985 66.735 8.160 ;
        RECT 65.730 3.865 66.050 3.985 ;
        RECT 59.115 3.645 63.765 3.820 ;
        RECT 65.415 3.695 66.050 3.865 ;
        RECT 65.730 3.665 66.050 3.695 ;
        RECT 49.285 3.490 49.635 3.610 ;
        RECT 59.115 3.505 59.395 3.645 ;
        RECT 46.370 3.320 49.635 3.490 ;
        RECT 63.590 3.495 63.765 3.645 ;
        RECT 64.060 3.495 64.385 3.620 ;
        RECT 66.560 3.615 66.735 7.985 ;
        RECT 76.335 7.725 76.615 8.095 ;
        RECT 77.705 8.050 77.965 8.095 ;
        RECT 77.675 7.805 77.995 8.050 ;
        RECT 77.705 7.760 77.965 7.805 ;
        RECT 79.405 7.760 79.665 8.095 ;
        RECT 77.345 7.065 77.625 7.435 ;
        RECT 77.765 6.645 77.905 7.760 ;
        RECT 78.385 7.065 78.665 7.435 ;
        RECT 77.085 6.505 77.905 6.645 ;
        RECT 74.305 6.075 74.565 6.395 ;
        RECT 74.365 4.355 74.505 6.075 ;
        RECT 77.085 5.800 77.225 6.505 ;
        RECT 78.725 6.075 78.985 6.395 ;
        RECT 74.975 5.430 75.255 5.800 ;
        RECT 77.015 5.430 77.295 5.800 ;
        RECT 74.305 4.035 74.565 4.355 ;
        RECT 75.045 4.015 75.185 5.430 ;
        RECT 76.665 4.690 76.945 5.060 ;
        RECT 77.085 4.355 77.225 5.430 ;
        RECT 78.035 5.030 78.315 5.400 ;
        RECT 78.785 5.375 78.925 6.075 ;
        RECT 78.725 5.055 78.985 5.375 ;
        RECT 77.025 4.035 77.285 4.355 ;
        RECT 77.695 4.350 77.975 4.720 ;
        RECT 79.465 4.355 79.605 7.760 ;
        RECT 79.405 4.035 79.665 4.355 ;
        RECT 74.985 3.695 75.245 4.015 ;
        RECT 76.335 3.815 76.615 3.870 ;
        RECT 82.635 3.860 82.795 9.030 ;
        RECT 83.750 8.940 84.075 9.030 ;
        RECT 86.140 9.145 86.465 9.270 ;
        RECT 89.320 9.170 89.490 9.550 ;
        RECT 99.855 9.200 100.015 9.550 ;
        RECT 100.970 9.200 101.295 9.265 ;
        RECT 86.140 9.140 86.925 9.145 ;
        RECT 89.270 9.140 89.550 9.170 ;
        RECT 86.140 8.975 89.550 9.140 ;
        RECT 86.140 8.945 86.465 8.975 ;
        RECT 86.925 8.970 89.550 8.975 ;
        RECT 82.950 8.565 83.270 8.890 ;
        RECT 89.270 8.830 89.550 8.970 ;
        RECT 99.855 9.030 101.295 9.200 ;
        RECT 82.980 8.330 83.150 8.565 ;
        RECT 82.980 8.155 83.155 8.330 ;
        RECT 82.980 7.980 83.955 8.155 ;
        RECT 82.950 3.860 83.270 3.980 ;
        RECT 76.335 3.640 80.985 3.815 ;
        RECT 82.635 3.690 83.270 3.860 ;
        RECT 82.950 3.660 83.270 3.690 ;
        RECT 66.505 3.495 66.855 3.615 ;
        RECT 76.335 3.500 76.615 3.640 ;
        RECT 63.590 3.325 66.855 3.495 ;
        RECT 29.620 3.290 29.945 3.320 ;
        RECT 32.065 3.260 32.415 3.320 ;
        RECT 46.840 3.290 47.165 3.320 ;
        RECT 49.285 3.260 49.635 3.320 ;
        RECT 64.060 3.295 64.385 3.325 ;
        RECT 66.505 3.265 66.855 3.325 ;
        RECT 80.810 3.490 80.985 3.640 ;
        RECT 81.280 3.490 81.605 3.615 ;
        RECT 83.780 3.610 83.955 7.980 ;
        RECT 93.555 7.725 93.835 8.095 ;
        RECT 94.925 8.050 95.185 8.095 ;
        RECT 94.895 7.805 95.215 8.050 ;
        RECT 94.925 7.760 95.185 7.805 ;
        RECT 96.625 7.760 96.885 8.095 ;
        RECT 94.565 7.065 94.845 7.435 ;
        RECT 94.985 6.645 95.125 7.760 ;
        RECT 95.605 7.065 95.885 7.435 ;
        RECT 94.305 6.505 95.125 6.645 ;
        RECT 91.525 6.075 91.785 6.395 ;
        RECT 91.585 4.355 91.725 6.075 ;
        RECT 94.305 5.800 94.445 6.505 ;
        RECT 95.945 6.075 96.205 6.395 ;
        RECT 92.195 5.430 92.475 5.800 ;
        RECT 94.235 5.430 94.515 5.800 ;
        RECT 91.525 4.035 91.785 4.355 ;
        RECT 92.265 4.015 92.405 5.430 ;
        RECT 93.885 4.690 94.165 5.060 ;
        RECT 94.305 4.355 94.445 5.430 ;
        RECT 95.255 5.030 95.535 5.400 ;
        RECT 96.005 5.375 96.145 6.075 ;
        RECT 95.945 5.055 96.205 5.375 ;
        RECT 94.245 4.035 94.505 4.355 ;
        RECT 94.915 4.350 95.195 4.720 ;
        RECT 96.685 4.355 96.825 7.760 ;
        RECT 96.625 4.035 96.885 4.355 ;
        RECT 92.205 3.695 92.465 4.015 ;
        RECT 93.555 3.815 93.835 3.870 ;
        RECT 99.855 3.860 100.015 9.030 ;
        RECT 100.970 8.940 101.295 9.030 ;
        RECT 100.170 8.565 100.490 8.890 ;
        RECT 100.200 8.330 100.370 8.565 ;
        RECT 100.200 8.155 100.375 8.330 ;
        RECT 100.200 7.980 101.175 8.155 ;
        RECT 100.170 3.860 100.490 3.980 ;
        RECT 93.555 3.640 98.205 3.815 ;
        RECT 99.855 3.690 100.490 3.860 ;
        RECT 100.170 3.660 100.490 3.690 ;
        RECT 83.725 3.490 84.075 3.610 ;
        RECT 93.555 3.500 93.835 3.640 ;
        RECT 80.810 3.320 84.075 3.490 ;
        RECT 98.030 3.490 98.205 3.640 ;
        RECT 98.500 3.490 98.825 3.615 ;
        RECT 101.000 3.610 101.175 7.980 ;
        RECT 100.945 3.490 101.295 3.610 ;
        RECT 98.030 3.320 101.295 3.490 ;
        RECT 81.280 3.290 81.605 3.320 ;
        RECT 83.725 3.260 84.075 3.320 ;
        RECT 98.500 3.290 98.825 3.320 ;
        RECT 100.945 3.260 101.295 3.320 ;
      LAYER met3 ;
        RECT 19.915 9.620 20.285 9.690 ;
        RECT 37.135 9.620 37.505 9.690 ;
        RECT 54.355 9.625 54.725 9.695 ;
        RECT 19.915 9.320 27.065 9.620 ;
        RECT 37.135 9.320 44.285 9.620 ;
        RECT 54.355 9.325 61.505 9.625 ;
        RECT 24.680 8.090 24.980 9.320 ;
        RECT 24.180 7.790 24.980 8.090 ;
        RECT 24.560 7.745 24.980 7.790 ;
        RECT 25.710 8.100 26.015 9.320 ;
        RECT 24.560 7.720 24.860 7.745 ;
        RECT 25.710 7.430 26.010 8.100 ;
        RECT 26.765 7.465 27.065 9.320 ;
        RECT 41.900 8.090 42.200 9.320 ;
        RECT 41.400 7.790 42.200 8.090 ;
        RECT 41.780 7.745 42.200 7.790 ;
        RECT 42.930 8.100 43.235 9.320 ;
        RECT 41.780 7.720 42.080 7.745 ;
        RECT 25.670 7.415 26.010 7.430 ;
        RECT 25.660 7.400 26.010 7.415 ;
        RECT 25.190 7.100 26.010 7.400 ;
        RECT 26.690 7.400 27.065 7.465 ;
        RECT 42.930 7.430 43.230 8.100 ;
        RECT 43.985 7.465 44.285 9.320 ;
        RECT 59.120 8.095 59.420 9.325 ;
        RECT 58.620 7.795 59.420 8.095 ;
        RECT 59.000 7.750 59.420 7.795 ;
        RECT 60.150 8.105 60.455 9.325 ;
        RECT 59.000 7.725 59.300 7.750 ;
        RECT 42.890 7.415 43.230 7.430 ;
        RECT 42.880 7.400 43.230 7.415 ;
        RECT 26.690 7.100 27.500 7.400 ;
        RECT 42.410 7.100 43.230 7.400 ;
        RECT 43.910 7.400 44.285 7.465 ;
        RECT 60.150 7.435 60.450 8.105 ;
        RECT 61.205 7.470 61.505 9.325 ;
        RECT 71.575 9.620 71.945 9.690 ;
        RECT 88.795 9.620 89.165 9.690 ;
        RECT 71.575 9.320 78.725 9.620 ;
        RECT 88.795 9.320 95.945 9.620 ;
        RECT 76.340 8.090 76.640 9.320 ;
        RECT 75.840 7.790 76.640 8.090 ;
        RECT 76.220 7.745 76.640 7.790 ;
        RECT 77.370 8.100 77.675 9.320 ;
        RECT 76.220 7.720 76.520 7.745 ;
        RECT 60.110 7.420 60.450 7.435 ;
        RECT 60.100 7.405 60.450 7.420 ;
        RECT 43.910 7.100 44.720 7.400 ;
        RECT 59.630 7.105 60.450 7.405 ;
        RECT 61.130 7.405 61.505 7.470 ;
        RECT 77.370 7.430 77.670 8.100 ;
        RECT 78.425 7.465 78.725 9.320 ;
        RECT 93.560 8.090 93.860 9.320 ;
        RECT 93.060 7.790 93.860 8.090 ;
        RECT 93.440 7.745 93.860 7.790 ;
        RECT 94.590 8.100 94.895 9.320 ;
        RECT 93.440 7.720 93.740 7.745 ;
        RECT 77.330 7.415 77.670 7.430 ;
        RECT 61.130 7.105 61.940 7.405 ;
        RECT 77.320 7.400 77.670 7.415 ;
        RECT 25.660 7.085 26.010 7.100 ;
        RECT 26.700 7.085 27.055 7.100 ;
        RECT 42.880 7.085 43.230 7.100 ;
        RECT 43.920 7.085 44.275 7.100 ;
        RECT 60.100 7.090 60.450 7.105 ;
        RECT 61.140 7.090 61.495 7.105 ;
        RECT 76.850 7.100 77.670 7.400 ;
        RECT 78.350 7.400 78.725 7.465 ;
        RECT 94.590 7.430 94.890 8.100 ;
        RECT 95.645 7.465 95.945 9.320 ;
        RECT 94.550 7.415 94.890 7.430 ;
        RECT 94.540 7.400 94.890 7.415 ;
        RECT 78.350 7.100 79.160 7.400 ;
        RECT 94.070 7.100 94.890 7.400 ;
        RECT 95.570 7.400 95.945 7.465 ;
        RECT 95.570 7.100 96.380 7.400 ;
        RECT 60.110 7.085 60.450 7.090 ;
        RECT 25.670 7.080 26.010 7.085 ;
        RECT 25.685 7.040 25.985 7.080 ;
        RECT 26.755 7.060 27.055 7.085 ;
        RECT 42.890 7.080 43.230 7.085 ;
        RECT 42.905 7.040 43.205 7.080 ;
        RECT 43.975 7.060 44.275 7.085 ;
        RECT 60.125 7.045 60.425 7.085 ;
        RECT 61.195 7.065 61.495 7.090 ;
        RECT 77.320 7.085 77.670 7.100 ;
        RECT 78.360 7.085 78.715 7.100 ;
        RECT 94.540 7.085 94.890 7.100 ;
        RECT 95.580 7.085 95.935 7.100 ;
        RECT 77.330 7.080 77.670 7.085 ;
        RECT 77.345 7.040 77.645 7.080 ;
        RECT 78.415 7.060 78.715 7.085 ;
        RECT 94.550 7.080 94.890 7.085 ;
        RECT 94.565 7.040 94.865 7.080 ;
        RECT 95.635 7.060 95.935 7.085 ;
        RECT 23.290 5.765 23.620 5.780 ;
        RECT 25.330 5.765 25.660 5.780 ;
        RECT 23.290 5.465 25.660 5.765 ;
        RECT 23.290 5.450 23.620 5.465 ;
        RECT 25.330 5.450 25.660 5.465 ;
        RECT 40.510 5.765 40.840 5.780 ;
        RECT 42.550 5.765 42.880 5.780 ;
        RECT 40.510 5.465 42.880 5.765 ;
        RECT 40.510 5.450 40.840 5.465 ;
        RECT 42.550 5.450 42.880 5.465 ;
        RECT 57.730 5.770 58.060 5.785 ;
        RECT 59.770 5.770 60.100 5.785 ;
        RECT 57.730 5.470 60.100 5.770 ;
        RECT 57.730 5.455 58.060 5.470 ;
        RECT 59.770 5.455 60.100 5.470 ;
        RECT 74.950 5.765 75.280 5.780 ;
        RECT 76.990 5.765 77.320 5.780 ;
        RECT 74.950 5.465 77.320 5.765 ;
        RECT 74.950 5.450 75.280 5.465 ;
        RECT 76.990 5.450 77.320 5.465 ;
        RECT 92.170 5.765 92.500 5.780 ;
        RECT 94.210 5.765 94.540 5.780 ;
        RECT 92.170 5.465 94.540 5.765 ;
        RECT 92.170 5.450 92.500 5.465 ;
        RECT 94.210 5.450 94.540 5.465 ;
        RECT 26.350 5.365 26.680 5.380 ;
        RECT 43.570 5.365 43.900 5.380 ;
        RECT 60.790 5.370 61.120 5.385 ;
        RECT 26.350 5.065 27.150 5.365 ;
        RECT 43.570 5.065 44.370 5.365 ;
        RECT 60.790 5.070 61.590 5.370 ;
        RECT 78.010 5.365 78.340 5.380 ;
        RECT 95.230 5.365 95.560 5.380 ;
        RECT 26.350 5.050 26.680 5.065 ;
        RECT 43.570 5.050 43.900 5.065 ;
        RECT 60.790 5.055 61.120 5.070 ;
        RECT 78.010 5.065 78.810 5.365 ;
        RECT 95.230 5.065 96.030 5.365 ;
        RECT 24.980 5.025 25.310 5.040 ;
        RECT 24.520 4.725 25.320 5.025 ;
        RECT 26.365 5.020 26.665 5.050 ;
        RECT 42.200 5.025 42.530 5.040 ;
        RECT 41.740 4.725 42.540 5.025 ;
        RECT 43.585 5.020 43.885 5.050 ;
        RECT 59.420 5.030 59.750 5.045 ;
        RECT 58.960 4.730 59.760 5.030 ;
        RECT 60.805 5.025 61.105 5.055 ;
        RECT 78.010 5.050 78.340 5.065 ;
        RECT 95.230 5.050 95.560 5.065 ;
        RECT 76.640 5.025 76.970 5.040 ;
        RECT 24.980 4.710 25.310 4.725 ;
        RECT 42.200 4.710 42.530 4.725 ;
        RECT 59.420 4.715 59.750 4.730 ;
        RECT 76.180 4.725 76.980 5.025 ;
        RECT 78.025 5.020 78.325 5.050 ;
        RECT 93.860 5.025 94.190 5.040 ;
        RECT 93.400 4.725 94.200 5.025 ;
        RECT 95.245 5.020 95.545 5.050 ;
        RECT 76.640 4.710 76.970 4.725 ;
        RECT 93.860 4.710 94.190 4.725 ;
        RECT 26.010 4.685 26.340 4.700 ;
        RECT 43.230 4.685 43.560 4.700 ;
        RECT 60.450 4.690 60.780 4.705 ;
        RECT 26.010 4.385 26.810 4.685 ;
        RECT 43.230 4.385 44.030 4.685 ;
        RECT 60.450 4.390 61.250 4.690 ;
        RECT 77.670 4.685 78.000 4.700 ;
        RECT 94.890 4.685 95.220 4.700 ;
        RECT 26.010 4.370 26.395 4.385 ;
        RECT 43.230 4.370 43.615 4.385 ;
        RECT 60.450 4.375 60.835 4.390 ;
        RECT 26.095 4.360 26.395 4.370 ;
        RECT 43.315 4.360 43.615 4.370 ;
        RECT 60.535 4.365 60.835 4.375 ;
        RECT 77.670 4.385 78.470 4.685 ;
        RECT 94.890 4.385 95.690 4.685 ;
        RECT 77.670 4.370 78.055 4.385 ;
        RECT 94.890 4.370 95.275 4.385 ;
        RECT 77.755 4.360 78.055 4.370 ;
        RECT 94.975 4.360 95.275 4.370 ;
        RECT 24.650 3.835 24.980 3.850 ;
        RECT 41.870 3.835 42.200 3.850 ;
        RECT 59.090 3.840 59.420 3.855 ;
        RECT 24.180 3.535 24.980 3.835 ;
        RECT 41.400 3.535 42.200 3.835 ;
        RECT 58.620 3.540 59.420 3.840 ;
        RECT 76.310 3.835 76.640 3.850 ;
        RECT 93.530 3.835 93.860 3.850 ;
        RECT 59.080 3.535 59.420 3.540 ;
        RECT 75.840 3.535 76.640 3.835 ;
        RECT 93.060 3.535 93.860 3.835 ;
        RECT 24.640 3.530 24.980 3.535 ;
        RECT 41.860 3.530 42.200 3.535 ;
        RECT 24.650 3.520 24.980 3.530 ;
        RECT 41.870 3.520 42.200 3.530 ;
        RECT 59.090 3.525 59.420 3.535 ;
        RECT 76.300 3.530 76.640 3.535 ;
        RECT 93.520 3.530 93.860 3.535 ;
        RECT 76.310 3.520 76.640 3.530 ;
        RECT 93.530 3.520 93.860 3.530 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r2
MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r2
  CLASS BLOCK ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ea_8_b0r2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 99.425 BY 12.460 ;
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 23.805 8.235 23.975 9.505 ;
        RECT 29.420 8.235 29.590 9.505 ;
        RECT 29.420 2.955 29.590 4.225 ;
      LAYER met1 ;
        RECT 23.720 8.405 24.070 8.465 ;
        RECT 29.340 8.405 29.680 8.475 ;
        RECT 23.720 8.375 24.205 8.405 ;
        RECT 29.340 8.400 29.820 8.405 ;
        RECT 29.325 8.375 29.820 8.400 ;
        RECT 23.720 8.235 29.820 8.375 ;
        RECT 23.720 8.205 29.680 8.235 ;
        RECT 23.720 8.175 24.070 8.205 ;
        RECT 29.340 8.125 29.680 8.205 ;
        RECT 29.350 4.225 29.690 4.350 ;
        RECT 29.350 4.055 29.820 4.225 ;
        RECT 29.350 4.000 29.690 4.055 ;
      LAYER met2 ;
        RECT 23.750 8.130 24.040 8.510 ;
        RECT 29.340 8.125 29.680 8.475 ;
        RECT 29.425 4.350 29.595 8.125 ;
        RECT 29.350 4.000 29.690 4.350 ;
      LAYER met3 ;
        RECT 23.715 8.465 24.065 12.460 ;
        RECT 23.720 8.130 24.070 8.465 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 40.130 8.235 40.300 9.505 ;
        RECT 45.745 8.235 45.915 9.505 ;
        RECT 45.745 2.955 45.915 4.225 ;
      LAYER met1 ;
        RECT 40.045 8.405 40.395 8.465 ;
        RECT 45.665 8.405 46.005 8.475 ;
        RECT 40.045 8.375 40.530 8.405 ;
        RECT 45.665 8.400 46.145 8.405 ;
        RECT 45.650 8.375 46.145 8.400 ;
        RECT 40.045 8.235 46.145 8.375 ;
        RECT 40.045 8.205 46.005 8.235 ;
        RECT 40.045 8.175 40.395 8.205 ;
        RECT 45.665 8.125 46.005 8.205 ;
        RECT 45.675 4.225 46.015 4.350 ;
        RECT 45.675 4.055 46.145 4.225 ;
        RECT 45.675 4.000 46.015 4.055 ;
      LAYER met2 ;
        RECT 40.075 8.130 40.365 8.510 ;
        RECT 45.665 8.125 46.005 8.475 ;
        RECT 45.750 4.350 45.920 8.125 ;
        RECT 45.675 4.000 46.015 4.350 ;
      LAYER met3 ;
        RECT 40.040 8.465 40.390 12.460 ;
        RECT 40.045 8.130 40.395 8.465 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 56.455 8.235 56.625 9.505 ;
        RECT 62.070 8.235 62.240 9.505 ;
        RECT 62.070 2.955 62.240 4.225 ;
      LAYER met1 ;
        RECT 56.370 8.405 56.720 8.465 ;
        RECT 61.990 8.405 62.330 8.475 ;
        RECT 56.370 8.375 56.855 8.405 ;
        RECT 61.990 8.400 62.470 8.405 ;
        RECT 61.975 8.375 62.470 8.400 ;
        RECT 56.370 8.235 62.470 8.375 ;
        RECT 56.370 8.205 62.330 8.235 ;
        RECT 56.370 8.175 56.720 8.205 ;
        RECT 61.990 8.125 62.330 8.205 ;
        RECT 62.000 4.225 62.340 4.350 ;
        RECT 62.000 4.055 62.470 4.225 ;
        RECT 62.000 4.000 62.340 4.055 ;
      LAYER met2 ;
        RECT 56.400 8.130 56.690 8.510 ;
        RECT 61.990 8.125 62.330 8.475 ;
        RECT 62.075 4.350 62.245 8.125 ;
        RECT 62.000 4.000 62.340 4.350 ;
      LAYER met3 ;
        RECT 56.365 8.465 56.715 12.460 ;
        RECT 56.370 8.130 56.720 8.465 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 72.780 8.235 72.950 9.505 ;
        RECT 78.395 8.235 78.565 9.505 ;
        RECT 78.395 2.955 78.565 4.225 ;
      LAYER met1 ;
        RECT 72.695 8.405 73.045 8.465 ;
        RECT 78.315 8.405 78.655 8.475 ;
        RECT 72.695 8.375 73.180 8.405 ;
        RECT 78.315 8.400 78.795 8.405 ;
        RECT 78.300 8.375 78.795 8.400 ;
        RECT 72.695 8.235 78.795 8.375 ;
        RECT 72.695 8.205 78.655 8.235 ;
        RECT 72.695 8.175 73.045 8.205 ;
        RECT 78.315 8.125 78.655 8.205 ;
        RECT 78.325 4.225 78.665 4.350 ;
        RECT 78.325 4.055 78.795 4.225 ;
        RECT 78.325 4.000 78.665 4.055 ;
      LAYER met2 ;
        RECT 72.725 8.130 73.015 8.510 ;
        RECT 78.315 8.125 78.655 8.475 ;
        RECT 78.400 4.350 78.570 8.125 ;
        RECT 78.325 4.000 78.665 4.350 ;
      LAYER met3 ;
        RECT 72.690 8.465 73.040 12.460 ;
        RECT 72.695 8.130 73.045 8.465 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 89.105 8.235 89.275 9.505 ;
        RECT 94.720 8.235 94.890 9.505 ;
        RECT 94.720 2.955 94.890 4.225 ;
      LAYER met1 ;
        RECT 89.020 8.405 89.370 8.465 ;
        RECT 94.640 8.405 94.980 8.475 ;
        RECT 89.020 8.375 89.505 8.405 ;
        RECT 94.640 8.400 95.120 8.405 ;
        RECT 94.625 8.375 95.120 8.400 ;
        RECT 89.020 8.235 95.120 8.375 ;
        RECT 89.020 8.205 94.980 8.235 ;
        RECT 89.020 8.175 89.370 8.205 ;
        RECT 94.640 8.125 94.980 8.205 ;
        RECT 94.650 4.225 94.990 4.350 ;
        RECT 94.650 4.055 95.120 4.225 ;
        RECT 94.650 4.000 94.990 4.055 ;
      LAYER met2 ;
        RECT 89.050 8.130 89.340 8.510 ;
        RECT 94.640 8.125 94.980 8.475 ;
        RECT 94.725 4.350 94.895 8.125 ;
        RECT 94.650 4.000 94.990 4.350 ;
      LAYER met3 ;
        RECT 89.015 8.465 89.365 12.460 ;
        RECT 89.020 8.130 89.370 8.465 ;
    END
  END s5
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 33.575 5.100 33.750 5.160 ;
        RECT 33.570 4.755 33.750 5.100 ;
        RECT 33.575 4.015 33.750 4.755 ;
        RECT 33.575 3.580 33.745 4.015 ;
        RECT 33.580 1.870 33.750 2.380 ;
      LAYER met1 ;
        RECT 33.515 3.545 33.805 3.780 ;
        RECT 33.515 3.540 33.745 3.545 ;
        RECT 33.575 2.440 33.745 3.540 ;
        RECT 33.515 2.180 33.810 2.440 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 49.900 5.100 50.075 5.160 ;
        RECT 49.895 4.755 50.075 5.100 ;
        RECT 49.900 4.015 50.075 4.755 ;
        RECT 49.900 3.580 50.070 4.015 ;
        RECT 49.905 1.870 50.075 2.380 ;
      LAYER met1 ;
        RECT 49.840 3.545 50.130 3.780 ;
        RECT 49.840 3.540 50.070 3.545 ;
        RECT 49.900 2.440 50.070 3.540 ;
        RECT 49.840 2.180 50.135 2.440 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 66.225 5.100 66.400 5.160 ;
        RECT 66.220 4.755 66.400 5.100 ;
        RECT 66.225 4.015 66.400 4.755 ;
        RECT 66.225 3.580 66.395 4.015 ;
        RECT 66.230 1.870 66.400 2.380 ;
      LAYER met1 ;
        RECT 66.165 3.545 66.455 3.780 ;
        RECT 66.165 3.540 66.395 3.545 ;
        RECT 66.225 2.440 66.395 3.540 ;
        RECT 66.165 2.180 66.460 2.440 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 82.550 5.100 82.725 5.160 ;
        RECT 82.545 4.755 82.725 5.100 ;
        RECT 82.550 4.015 82.725 4.755 ;
        RECT 82.550 3.580 82.720 4.015 ;
        RECT 82.555 1.870 82.725 2.380 ;
      LAYER met1 ;
        RECT 82.490 3.545 82.780 3.780 ;
        RECT 82.490 3.540 82.720 3.545 ;
        RECT 82.550 2.440 82.720 3.540 ;
        RECT 82.490 2.180 82.785 2.440 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 98.875 5.100 99.050 5.160 ;
        RECT 98.870 4.755 99.050 5.100 ;
        RECT 98.875 4.015 99.050 4.755 ;
        RECT 98.875 3.580 99.045 4.015 ;
        RECT 98.880 1.870 99.050 2.380 ;
      LAYER met1 ;
        RECT 98.815 3.545 99.105 3.780 ;
        RECT 98.815 3.540 99.045 3.545 ;
        RECT 98.875 2.440 99.045 3.540 ;
        RECT 98.815 2.180 99.110 2.440 ;
    END
  END X5_Y1
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 15.225 8.235 15.395 9.505 ;
      LAYER met1 ;
        RECT 15.165 8.430 15.455 8.435 ;
        RECT 15.165 8.405 15.460 8.430 ;
        RECT 15.165 8.235 15.625 8.405 ;
        RECT 15.165 8.205 15.460 8.235 ;
        RECT 15.170 8.200 15.460 8.205 ;
    END
  END start
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 25.665 3.925 25.835 4.125 ;
        RECT 27.625 3.925 27.795 4.125 ;
        RECT 41.990 3.925 42.160 4.125 ;
        RECT 43.950 3.925 44.120 4.125 ;
        RECT 58.315 3.925 58.485 4.125 ;
        RECT 60.275 3.925 60.445 4.125 ;
        RECT 74.640 3.925 74.810 4.125 ;
        RECT 76.600 3.925 76.770 4.125 ;
        RECT 90.965 3.925 91.135 4.125 ;
        RECT 92.925 3.925 93.095 4.125 ;
        RECT 25.345 3.755 25.835 3.925 ;
        RECT 27.305 3.755 27.795 3.925 ;
        RECT 41.670 3.755 42.160 3.925 ;
        RECT 43.630 3.755 44.120 3.925 ;
        RECT 57.995 3.755 58.485 3.925 ;
        RECT 59.955 3.755 60.445 3.925 ;
        RECT 74.320 3.755 74.810 3.925 ;
        RECT 76.280 3.755 76.770 3.925 ;
        RECT 90.645 3.755 91.135 3.925 ;
        RECT 92.605 3.755 93.095 3.925 ;
        RECT 18.865 2.765 19.035 3.265 ;
        RECT 19.825 2.765 19.995 3.265 ;
        RECT 20.785 2.765 20.955 3.265 ;
        RECT 21.305 2.765 21.475 3.265 ;
        RECT 22.265 2.765 22.435 3.265 ;
        RECT 24.705 2.765 24.875 3.265 ;
        RECT 26.665 2.780 26.835 3.265 ;
        RECT 26.485 2.765 26.835 2.780 ;
        RECT 35.190 2.765 35.360 3.265 ;
        RECT 36.150 2.765 36.320 3.265 ;
        RECT 37.110 2.765 37.280 3.265 ;
        RECT 37.630 2.765 37.800 3.265 ;
        RECT 38.590 2.765 38.760 3.265 ;
        RECT 41.030 2.765 41.200 3.265 ;
        RECT 42.990 2.780 43.160 3.265 ;
        RECT 42.810 2.765 43.160 2.780 ;
        RECT 51.515 2.765 51.685 3.265 ;
        RECT 52.475 2.765 52.645 3.265 ;
        RECT 53.435 2.765 53.605 3.265 ;
        RECT 53.955 2.765 54.125 3.265 ;
        RECT 54.915 2.765 55.085 3.265 ;
        RECT 57.355 2.765 57.525 3.265 ;
        RECT 59.315 2.780 59.485 3.265 ;
        RECT 59.135 2.765 59.485 2.780 ;
        RECT 67.840 2.765 68.010 3.265 ;
        RECT 68.800 2.765 68.970 3.265 ;
        RECT 69.760 2.765 69.930 3.265 ;
        RECT 70.280 2.765 70.450 3.265 ;
        RECT 71.240 2.765 71.410 3.265 ;
        RECT 73.680 2.765 73.850 3.265 ;
        RECT 75.640 2.780 75.810 3.265 ;
        RECT 75.460 2.765 75.810 2.780 ;
        RECT 84.165 2.765 84.335 3.265 ;
        RECT 85.125 2.765 85.295 3.265 ;
        RECT 86.085 2.765 86.255 3.265 ;
        RECT 86.605 2.765 86.775 3.265 ;
        RECT 87.565 2.765 87.735 3.265 ;
        RECT 90.005 2.765 90.175 3.265 ;
        RECT 91.965 2.780 92.135 3.265 ;
        RECT 91.785 2.765 92.135 2.780 ;
        RECT 18.535 1.600 28.350 2.765 ;
        RECT 29.410 1.600 29.580 2.225 ;
        RECT 32.155 1.600 32.325 2.225 ;
        RECT 33.145 1.600 33.315 2.230 ;
        RECT 34.860 1.600 44.675 2.765 ;
        RECT 45.735 1.600 45.905 2.225 ;
        RECT 48.480 1.600 48.650 2.225 ;
        RECT 49.470 1.600 49.640 2.230 ;
        RECT 51.185 1.600 61.000 2.765 ;
        RECT 62.060 1.600 62.230 2.225 ;
        RECT 64.805 1.600 64.975 2.225 ;
        RECT 65.795 1.600 65.965 2.230 ;
        RECT 67.510 1.600 77.325 2.765 ;
        RECT 78.385 1.600 78.555 2.225 ;
        RECT 81.130 1.600 81.300 2.225 ;
        RECT 82.120 1.600 82.290 2.230 ;
        RECT 83.835 1.600 93.650 2.765 ;
        RECT 94.710 1.600 94.880 2.225 ;
        RECT 97.455 1.600 97.625 2.225 ;
        RECT 98.445 1.600 98.615 2.230 ;
        RECT 0.000 0.000 99.420 1.600 ;
      LAYER met1 ;
        RECT 27.465 4.255 27.705 4.350 ;
        RECT 43.790 4.255 44.030 4.350 ;
        RECT 60.115 4.255 60.355 4.350 ;
        RECT 76.440 4.255 76.680 4.350 ;
        RECT 92.765 4.255 93.005 4.350 ;
        RECT 25.935 4.240 27.705 4.255 ;
        RECT 42.260 4.240 44.030 4.255 ;
        RECT 58.585 4.240 60.355 4.255 ;
        RECT 74.910 4.240 76.680 4.255 ;
        RECT 91.235 4.240 93.005 4.255 ;
        RECT 25.935 4.155 28.350 4.240 ;
        RECT 42.260 4.155 44.675 4.240 ;
        RECT 58.585 4.155 61.000 4.240 ;
        RECT 74.910 4.155 77.325 4.240 ;
        RECT 91.235 4.155 93.650 4.240 ;
        RECT 25.605 4.115 28.350 4.155 ;
        RECT 25.605 3.975 26.075 4.115 ;
        RECT 27.395 4.055 28.350 4.115 ;
        RECT 27.395 3.975 27.855 4.055 ;
        RECT 25.605 3.925 25.895 3.975 ;
        RECT 27.425 3.925 27.855 3.975 ;
        RECT 27.425 3.915 27.745 3.925 ;
        RECT 28.165 2.880 28.350 4.055 ;
        RECT 41.930 4.115 44.675 4.155 ;
        RECT 41.930 3.975 42.400 4.115 ;
        RECT 43.720 4.055 44.675 4.115 ;
        RECT 43.720 3.975 44.180 4.055 ;
        RECT 41.930 3.925 42.220 3.975 ;
        RECT 43.750 3.925 44.180 3.975 ;
        RECT 43.750 3.915 44.070 3.925 ;
        RECT 44.490 2.880 44.675 4.055 ;
        RECT 58.255 4.115 61.000 4.155 ;
        RECT 58.255 3.975 58.725 4.115 ;
        RECT 60.045 4.055 61.000 4.115 ;
        RECT 60.045 3.975 60.505 4.055 ;
        RECT 58.255 3.925 58.545 3.975 ;
        RECT 60.075 3.925 60.505 3.975 ;
        RECT 60.075 3.915 60.395 3.925 ;
        RECT 60.815 2.880 61.000 4.055 ;
        RECT 74.580 4.115 77.325 4.155 ;
        RECT 74.580 3.975 75.050 4.115 ;
        RECT 76.370 4.055 77.325 4.115 ;
        RECT 76.370 3.975 76.830 4.055 ;
        RECT 74.580 3.925 74.870 3.975 ;
        RECT 76.400 3.925 76.830 3.975 ;
        RECT 76.400 3.915 76.720 3.925 ;
        RECT 77.140 2.880 77.325 4.055 ;
        RECT 90.905 4.115 93.650 4.155 ;
        RECT 90.905 3.975 91.375 4.115 ;
        RECT 92.695 4.055 93.650 4.115 ;
        RECT 92.695 3.975 93.155 4.055 ;
        RECT 90.905 3.925 91.195 3.975 ;
        RECT 92.725 3.925 93.155 3.975 ;
        RECT 92.725 3.915 93.045 3.925 ;
        RECT 93.465 2.880 93.650 4.055 ;
        RECT 28.160 2.860 28.350 2.880 ;
        RECT 44.485 2.860 44.675 2.880 ;
        RECT 60.810 2.860 61.000 2.880 ;
        RECT 77.135 2.860 77.325 2.880 ;
        RECT 93.460 2.860 93.650 2.880 ;
        RECT 28.155 2.795 28.350 2.860 ;
        RECT 44.480 2.795 44.675 2.860 ;
        RECT 60.805 2.795 61.000 2.860 ;
        RECT 77.130 2.795 77.325 2.860 ;
        RECT 93.455 2.795 93.650 2.860 ;
        RECT 18.535 1.600 28.350 2.795 ;
        RECT 34.860 1.600 44.675 2.795 ;
        RECT 51.185 1.600 61.000 2.795 ;
        RECT 67.510 1.600 77.325 2.795 ;
        RECT 83.835 1.600 93.650 2.795 ;
        RECT 0.000 0.000 99.420 1.600 ;
      LAYER met2 ;
        RECT 27.445 4.135 27.725 4.510 ;
        RECT 43.770 4.135 44.050 4.510 ;
        RECT 60.095 4.135 60.375 4.510 ;
        RECT 76.420 4.135 76.700 4.510 ;
        RECT 92.745 4.135 93.025 4.510 ;
        RECT 27.455 3.885 27.715 4.135 ;
        RECT 43.780 3.885 44.040 4.135 ;
        RECT 60.105 3.885 60.365 4.135 ;
        RECT 76.430 3.885 76.690 4.135 ;
        RECT 92.755 3.885 93.015 4.135 ;
      LAYER met3 ;
        RECT 27.425 4.485 27.755 4.885 ;
        RECT 43.750 4.485 44.080 4.885 ;
        RECT 60.075 4.485 60.405 4.885 ;
        RECT 76.400 4.485 76.730 4.885 ;
        RECT 92.725 4.485 93.055 4.885 ;
        RECT 27.420 4.155 27.755 4.485 ;
        RECT 43.745 4.155 44.080 4.485 ;
        RECT 60.070 4.155 60.405 4.485 ;
        RECT 76.395 4.155 76.730 4.485 ;
        RECT 92.720 4.155 93.055 4.485 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 10.860 99.425 12.460 ;
        RECT 15.215 10.235 15.385 10.860 ;
        RECT 23.795 10.235 23.965 10.860 ;
        RECT 24.750 10.315 24.920 10.595 ;
        RECT 24.750 10.145 24.980 10.315 ;
        RECT 29.410 10.235 29.580 10.860 ;
        RECT 32.155 10.235 32.325 10.860 ;
        RECT 33.150 10.230 33.320 10.860 ;
        RECT 40.120 10.235 40.290 10.860 ;
        RECT 41.075 10.315 41.245 10.595 ;
        RECT 41.075 10.145 41.305 10.315 ;
        RECT 45.735 10.235 45.905 10.860 ;
        RECT 48.480 10.235 48.650 10.860 ;
        RECT 49.475 10.230 49.645 10.860 ;
        RECT 56.445 10.235 56.615 10.860 ;
        RECT 57.400 10.315 57.570 10.595 ;
        RECT 57.400 10.145 57.630 10.315 ;
        RECT 62.060 10.235 62.230 10.860 ;
        RECT 64.805 10.235 64.975 10.860 ;
        RECT 65.800 10.230 65.970 10.860 ;
        RECT 72.770 10.235 72.940 10.860 ;
        RECT 73.725 10.315 73.895 10.595 ;
        RECT 73.725 10.145 73.955 10.315 ;
        RECT 78.385 10.235 78.555 10.860 ;
        RECT 81.130 10.235 81.300 10.860 ;
        RECT 82.125 10.230 82.295 10.860 ;
        RECT 89.095 10.235 89.265 10.860 ;
        RECT 90.050 10.315 90.220 10.595 ;
        RECT 90.050 10.145 90.280 10.315 ;
        RECT 94.710 10.235 94.880 10.860 ;
        RECT 97.455 10.235 97.625 10.860 ;
        RECT 98.450 10.230 98.620 10.860 ;
        RECT 24.810 8.535 24.980 10.145 ;
        RECT 41.135 8.535 41.305 10.145 ;
        RECT 57.460 8.535 57.630 10.145 ;
        RECT 73.785 8.535 73.955 10.145 ;
        RECT 90.110 8.535 90.280 10.145 ;
        RECT 24.750 8.365 24.980 8.535 ;
        RECT 41.075 8.365 41.305 8.535 ;
        RECT 57.400 8.365 57.630 8.535 ;
        RECT 73.725 8.365 73.955 8.535 ;
        RECT 90.050 8.365 90.280 8.535 ;
        RECT 24.750 7.305 24.920 8.365 ;
        RECT 41.075 7.305 41.245 8.365 ;
        RECT 57.400 7.305 57.570 8.365 ;
        RECT 73.725 7.305 73.895 8.365 ;
        RECT 90.050 7.305 90.220 8.365 ;
      LAYER met1 ;
        RECT 0.000 10.860 99.425 12.460 ;
        RECT 24.370 8.785 24.545 10.860 ;
        RECT 24.750 8.785 25.040 8.815 ;
        RECT 24.370 8.600 25.040 8.785 ;
        RECT 40.695 8.785 40.870 10.860 ;
        RECT 41.075 8.785 41.365 8.815 ;
        RECT 40.695 8.600 41.365 8.785 ;
        RECT 57.020 8.785 57.195 10.860 ;
        RECT 57.400 8.785 57.690 8.815 ;
        RECT 57.020 8.600 57.690 8.785 ;
        RECT 73.345 8.785 73.520 10.860 ;
        RECT 73.725 8.785 74.015 8.815 ;
        RECT 73.345 8.600 74.015 8.785 ;
        RECT 89.670 8.785 89.845 10.860 ;
        RECT 90.050 8.785 90.340 8.815 ;
        RECT 89.670 8.600 90.340 8.785 ;
        RECT 24.750 8.585 25.040 8.600 ;
        RECT 41.075 8.585 41.365 8.600 ;
        RECT 57.400 8.585 57.690 8.600 ;
        RECT 73.725 8.585 74.015 8.600 ;
        RECT 90.050 8.585 90.340 8.600 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 14.995 8.740 17.805 8.745 ;
        RECT 23.575 8.740 26.385 8.745 ;
        RECT 29.190 8.740 32.980 8.745 ;
        RECT 39.900 8.740 42.710 8.745 ;
        RECT 45.515 8.740 49.305 8.745 ;
        RECT 56.225 8.740 59.035 8.745 ;
        RECT 61.840 8.740 65.630 8.745 ;
        RECT 72.550 8.740 75.360 8.745 ;
        RECT 78.165 8.740 81.955 8.745 ;
        RECT 88.875 8.740 91.685 8.745 ;
        RECT 94.490 8.740 98.280 8.745 ;
        RECT 14.995 6.655 99.420 8.740 ;
        RECT 15.000 4.000 99.420 6.655 ;
        RECT 17.785 3.985 99.420 4.000 ;
        RECT 28.175 3.720 34.120 3.985 ;
        RECT 44.500 3.720 50.445 3.985 ;
        RECT 60.825 3.720 66.770 3.985 ;
        RECT 77.150 3.720 83.095 3.985 ;
        RECT 93.475 3.720 99.420 3.985 ;
        RECT 29.190 3.715 32.980 3.720 ;
        RECT 45.515 3.715 49.305 3.720 ;
        RECT 61.840 3.715 65.630 3.720 ;
        RECT 78.165 3.715 81.955 3.720 ;
        RECT 94.490 3.715 98.280 3.720 ;
      LAYER li1 ;
        RECT 17.030 10.045 17.205 10.595 ;
        RECT 17.030 8.445 17.200 10.045 ;
        RECT 15.215 7.035 15.385 7.765 ;
        RECT 17.030 7.305 17.205 8.445 ;
        RECT 17.030 7.035 17.200 7.305 ;
        RECT 23.795 7.035 23.965 7.765 ;
        RECT 29.410 7.035 29.580 7.765 ;
        RECT 32.155 7.035 32.325 7.765 ;
        RECT 33.150 7.035 33.320 7.760 ;
        RECT 40.120 7.035 40.290 7.765 ;
        RECT 45.735 7.035 45.905 7.765 ;
        RECT 48.480 7.035 48.650 7.765 ;
        RECT 49.475 7.035 49.645 7.760 ;
        RECT 56.445 7.035 56.615 7.765 ;
        RECT 62.060 7.035 62.230 7.765 ;
        RECT 64.805 7.035 64.975 7.765 ;
        RECT 65.800 7.035 65.970 7.760 ;
        RECT 72.770 7.035 72.940 7.765 ;
        RECT 78.385 7.035 78.555 7.765 ;
        RECT 81.130 7.035 81.300 7.765 ;
        RECT 82.125 7.035 82.295 7.760 ;
        RECT 89.095 7.035 89.265 7.765 ;
        RECT 94.710 7.035 94.880 7.765 ;
        RECT 97.455 7.035 97.625 7.765 ;
        RECT 98.450 7.035 98.620 7.760 ;
        RECT 0.000 5.435 99.420 7.035 ;
        RECT 17.790 5.430 99.420 5.435 ;
        RECT 18.535 5.315 28.195 5.430 ;
        RECT 29.240 5.425 32.975 5.430 ;
        RECT 19.825 4.815 19.995 5.315 ;
        RECT 22.265 4.815 22.435 5.315 ;
        RECT 23.225 4.815 23.395 5.315 ;
        RECT 24.225 4.815 24.395 5.315 ;
        RECT 26.665 4.815 26.835 5.315 ;
        RECT 27.625 4.815 27.795 5.315 ;
        RECT 29.410 4.695 29.580 5.425 ;
        RECT 32.155 4.695 32.325 5.425 ;
        RECT 33.145 4.700 33.315 5.430 ;
        RECT 34.860 5.315 44.520 5.430 ;
        RECT 45.565 5.425 49.300 5.430 ;
        RECT 36.150 4.815 36.320 5.315 ;
        RECT 38.590 4.815 38.760 5.315 ;
        RECT 39.550 4.815 39.720 5.315 ;
        RECT 40.550 4.815 40.720 5.315 ;
        RECT 42.990 4.815 43.160 5.315 ;
        RECT 43.950 4.815 44.120 5.315 ;
        RECT 45.735 4.695 45.905 5.425 ;
        RECT 48.480 4.695 48.650 5.425 ;
        RECT 49.470 4.700 49.640 5.430 ;
        RECT 51.185 5.315 60.845 5.430 ;
        RECT 61.890 5.425 65.625 5.430 ;
        RECT 52.475 4.815 52.645 5.315 ;
        RECT 54.915 4.815 55.085 5.315 ;
        RECT 55.875 4.815 56.045 5.315 ;
        RECT 56.875 4.815 57.045 5.315 ;
        RECT 59.315 4.815 59.485 5.315 ;
        RECT 60.275 4.815 60.445 5.315 ;
        RECT 62.060 4.695 62.230 5.425 ;
        RECT 64.805 4.695 64.975 5.425 ;
        RECT 65.795 4.700 65.965 5.430 ;
        RECT 67.510 5.315 77.170 5.430 ;
        RECT 78.215 5.425 81.950 5.430 ;
        RECT 68.800 4.815 68.970 5.315 ;
        RECT 71.240 4.815 71.410 5.315 ;
        RECT 72.200 4.815 72.370 5.315 ;
        RECT 73.200 4.815 73.370 5.315 ;
        RECT 75.640 4.815 75.810 5.315 ;
        RECT 76.600 4.815 76.770 5.315 ;
        RECT 78.385 4.695 78.555 5.425 ;
        RECT 81.130 4.695 81.300 5.425 ;
        RECT 82.120 4.700 82.290 5.430 ;
        RECT 83.835 5.315 93.495 5.430 ;
        RECT 94.540 5.425 98.275 5.430 ;
        RECT 85.125 4.815 85.295 5.315 ;
        RECT 87.565 4.815 87.735 5.315 ;
        RECT 88.525 4.815 88.695 5.315 ;
        RECT 89.525 4.815 89.695 5.315 ;
        RECT 91.965 4.815 92.135 5.315 ;
        RECT 92.925 4.815 93.095 5.315 ;
        RECT 94.710 4.695 94.880 5.425 ;
        RECT 97.455 4.695 97.625 5.425 ;
        RECT 98.445 4.700 98.615 5.430 ;
      LAYER met1 ;
        RECT 16.970 9.145 17.260 9.175 ;
        RECT 16.800 8.975 17.260 9.145 ;
        RECT 16.970 8.945 17.260 8.975 ;
        RECT 0.000 5.435 99.420 7.035 ;
        RECT 17.790 5.430 99.420 5.435 ;
        RECT 18.535 5.285 28.195 5.430 ;
        RECT 29.240 5.425 32.975 5.430 ;
        RECT 34.860 5.285 44.520 5.430 ;
        RECT 45.565 5.425 49.300 5.430 ;
        RECT 51.185 5.285 60.845 5.430 ;
        RECT 61.890 5.425 65.625 5.430 ;
        RECT 67.510 5.285 77.170 5.430 ;
        RECT 78.215 5.425 81.950 5.430 ;
        RECT 83.835 5.285 93.495 5.430 ;
        RECT 94.540 5.425 98.275 5.430 ;
    END
  END vccd1
  OBS
      LAYER pwell ;
        RECT 18.695 2.625 18.865 2.765 ;
        RECT 18.675 2.605 18.865 2.625 ;
        RECT 21.135 2.605 21.305 2.765 ;
        RECT 23.575 2.605 23.745 2.765 ;
        RECT 26.015 2.625 26.185 2.765 ;
        RECT 35.020 2.625 35.190 2.765 ;
        RECT 26.015 2.605 26.205 2.625 ;
        RECT 18.675 2.595 18.845 2.605 ;
        RECT 26.035 2.595 26.205 2.605 ;
        RECT 35.000 2.605 35.190 2.625 ;
        RECT 37.460 2.605 37.630 2.765 ;
        RECT 39.900 2.605 40.070 2.765 ;
        RECT 42.340 2.625 42.510 2.765 ;
        RECT 51.345 2.625 51.515 2.765 ;
        RECT 42.340 2.605 42.530 2.625 ;
        RECT 35.000 2.595 35.170 2.605 ;
        RECT 42.360 2.595 42.530 2.605 ;
        RECT 51.325 2.605 51.515 2.625 ;
        RECT 53.785 2.605 53.955 2.765 ;
        RECT 56.225 2.605 56.395 2.765 ;
        RECT 58.665 2.625 58.835 2.765 ;
        RECT 67.670 2.625 67.840 2.765 ;
        RECT 58.665 2.605 58.855 2.625 ;
        RECT 51.325 2.595 51.495 2.605 ;
        RECT 58.685 2.595 58.855 2.605 ;
        RECT 67.650 2.605 67.840 2.625 ;
        RECT 70.110 2.605 70.280 2.765 ;
        RECT 72.550 2.605 72.720 2.765 ;
        RECT 74.990 2.625 75.160 2.765 ;
        RECT 83.995 2.625 84.165 2.765 ;
        RECT 74.990 2.605 75.180 2.625 ;
        RECT 67.650 2.595 67.820 2.605 ;
        RECT 75.010 2.595 75.180 2.605 ;
        RECT 83.975 2.605 84.165 2.625 ;
        RECT 86.435 2.605 86.605 2.765 ;
        RECT 88.875 2.605 89.045 2.765 ;
        RECT 91.315 2.625 91.485 2.765 ;
        RECT 91.315 2.605 91.505 2.625 ;
        RECT 83.975 2.595 84.145 2.605 ;
        RECT 91.335 2.595 91.505 2.605 ;
      LAYER li1 ;
        RECT 15.645 10.105 15.820 10.595 ;
        RECT 16.170 10.315 16.340 10.595 ;
        RECT 16.170 10.145 16.400 10.315 ;
        RECT 15.645 9.935 15.815 10.105 ;
        RECT 15.645 9.605 16.055 9.935 ;
        RECT 15.645 9.095 15.815 9.605 ;
        RECT 15.645 8.765 16.055 9.095 ;
        RECT 15.645 8.565 15.815 8.765 ;
        RECT 15.645 7.305 15.820 8.565 ;
        RECT 16.230 8.535 16.400 10.145 ;
        RECT 16.600 10.085 16.775 10.595 ;
        RECT 24.225 10.105 24.400 10.595 ;
        RECT 24.225 9.935 24.395 10.105 ;
        RECT 25.180 10.085 25.355 10.595 ;
        RECT 25.610 10.045 25.785 10.595 ;
        RECT 29.840 10.105 30.015 10.595 ;
        RECT 30.365 10.315 30.535 10.595 ;
        RECT 30.365 10.145 30.595 10.315 ;
        RECT 24.225 9.605 24.635 9.935 ;
        RECT 16.170 8.365 16.400 8.535 ;
        RECT 16.600 8.565 16.770 9.515 ;
        RECT 24.225 9.095 24.395 9.605 ;
        RECT 24.225 8.765 24.635 9.095 ;
        RECT 24.225 8.565 24.395 8.765 ;
        RECT 25.180 8.565 25.350 9.515 ;
        RECT 16.170 7.305 16.340 8.365 ;
        RECT 16.600 7.305 16.775 8.565 ;
        RECT 24.225 7.305 24.400 8.565 ;
        RECT 25.180 7.305 25.355 8.565 ;
        RECT 25.610 8.445 25.780 10.045 ;
        RECT 29.840 9.935 30.010 10.105 ;
        RECT 29.840 9.605 30.250 9.935 ;
        RECT 29.840 9.095 30.010 9.605 ;
        RECT 29.840 8.765 30.250 9.095 ;
        RECT 29.840 8.565 30.010 8.765 ;
        RECT 25.610 7.305 25.785 8.445 ;
        RECT 29.840 7.305 30.015 8.565 ;
        RECT 30.425 8.535 30.595 10.145 ;
        RECT 30.795 10.085 30.970 10.595 ;
        RECT 31.225 10.045 31.400 10.595 ;
        RECT 32.590 10.085 32.760 10.595 ;
        RECT 33.585 10.080 33.755 10.590 ;
        RECT 40.550 10.105 40.725 10.595 ;
        RECT 30.365 8.365 30.595 8.535 ;
        RECT 30.795 8.565 30.965 9.515 ;
        RECT 30.365 7.305 30.535 8.365 ;
        RECT 30.795 7.305 30.970 8.565 ;
        RECT 31.225 8.445 31.395 10.045 ;
        RECT 40.550 9.935 40.720 10.105 ;
        RECT 41.505 10.085 41.680 10.595 ;
        RECT 41.935 10.045 42.110 10.595 ;
        RECT 46.165 10.105 46.340 10.595 ;
        RECT 46.690 10.315 46.860 10.595 ;
        RECT 46.690 10.145 46.920 10.315 ;
        RECT 40.550 9.605 40.960 9.935 ;
        RECT 31.765 9.425 31.995 9.575 ;
        RECT 31.765 9.255 32.685 9.425 ;
        RECT 32.215 8.565 32.385 9.255 ;
        RECT 33.210 9.250 33.680 9.420 ;
        RECT 32.585 8.775 32.755 8.885 ;
        RECT 33.210 8.775 33.380 9.250 ;
        RECT 40.550 9.095 40.720 9.605 ;
        RECT 32.585 8.605 33.380 8.775 ;
        RECT 31.225 7.305 31.400 8.445 ;
        RECT 32.585 7.305 32.760 8.605 ;
        RECT 33.210 8.560 33.380 8.605 ;
        RECT 33.580 8.445 33.750 8.880 ;
        RECT 40.550 8.765 40.960 9.095 ;
        RECT 40.550 8.565 40.720 8.765 ;
        RECT 41.505 8.565 41.675 9.515 ;
        RECT 33.580 7.300 33.755 8.445 ;
        RECT 40.550 7.305 40.725 8.565 ;
        RECT 41.505 7.305 41.680 8.565 ;
        RECT 41.935 8.445 42.105 10.045 ;
        RECT 46.165 9.935 46.335 10.105 ;
        RECT 46.165 9.605 46.575 9.935 ;
        RECT 46.165 9.095 46.335 9.605 ;
        RECT 46.165 8.765 46.575 9.095 ;
        RECT 46.165 8.565 46.335 8.765 ;
        RECT 41.935 7.305 42.110 8.445 ;
        RECT 46.165 7.305 46.340 8.565 ;
        RECT 46.750 8.535 46.920 10.145 ;
        RECT 47.120 10.085 47.295 10.595 ;
        RECT 47.550 10.045 47.725 10.595 ;
        RECT 48.915 10.085 49.085 10.595 ;
        RECT 49.910 10.080 50.080 10.590 ;
        RECT 56.875 10.105 57.050 10.595 ;
        RECT 46.690 8.365 46.920 8.535 ;
        RECT 47.120 8.565 47.290 9.515 ;
        RECT 46.690 7.305 46.860 8.365 ;
        RECT 47.120 7.305 47.295 8.565 ;
        RECT 47.550 8.445 47.720 10.045 ;
        RECT 56.875 9.935 57.045 10.105 ;
        RECT 57.830 10.085 58.005 10.595 ;
        RECT 58.260 10.045 58.435 10.595 ;
        RECT 62.490 10.105 62.665 10.595 ;
        RECT 63.015 10.315 63.185 10.595 ;
        RECT 63.015 10.145 63.245 10.315 ;
        RECT 56.875 9.605 57.285 9.935 ;
        RECT 48.090 9.425 48.320 9.575 ;
        RECT 48.090 9.255 49.010 9.425 ;
        RECT 48.540 8.565 48.710 9.255 ;
        RECT 49.535 9.250 50.005 9.420 ;
        RECT 48.910 8.775 49.080 8.885 ;
        RECT 49.535 8.775 49.705 9.250 ;
        RECT 56.875 9.095 57.045 9.605 ;
        RECT 48.910 8.605 49.705 8.775 ;
        RECT 47.550 7.305 47.725 8.445 ;
        RECT 48.910 7.305 49.085 8.605 ;
        RECT 49.535 8.560 49.705 8.605 ;
        RECT 49.905 8.445 50.075 8.880 ;
        RECT 56.875 8.765 57.285 9.095 ;
        RECT 56.875 8.565 57.045 8.765 ;
        RECT 57.830 8.565 58.000 9.515 ;
        RECT 49.905 7.300 50.080 8.445 ;
        RECT 56.875 7.305 57.050 8.565 ;
        RECT 57.830 7.305 58.005 8.565 ;
        RECT 58.260 8.445 58.430 10.045 ;
        RECT 62.490 9.935 62.660 10.105 ;
        RECT 62.490 9.605 62.900 9.935 ;
        RECT 62.490 9.095 62.660 9.605 ;
        RECT 62.490 8.765 62.900 9.095 ;
        RECT 62.490 8.565 62.660 8.765 ;
        RECT 58.260 7.305 58.435 8.445 ;
        RECT 62.490 7.305 62.665 8.565 ;
        RECT 63.075 8.535 63.245 10.145 ;
        RECT 63.445 10.085 63.620 10.595 ;
        RECT 63.875 10.045 64.050 10.595 ;
        RECT 65.240 10.085 65.410 10.595 ;
        RECT 66.235 10.080 66.405 10.590 ;
        RECT 73.200 10.105 73.375 10.595 ;
        RECT 63.015 8.365 63.245 8.535 ;
        RECT 63.445 8.565 63.615 9.515 ;
        RECT 63.015 7.305 63.185 8.365 ;
        RECT 63.445 7.305 63.620 8.565 ;
        RECT 63.875 8.445 64.045 10.045 ;
        RECT 73.200 9.935 73.370 10.105 ;
        RECT 74.155 10.085 74.330 10.595 ;
        RECT 74.585 10.045 74.760 10.595 ;
        RECT 78.815 10.105 78.990 10.595 ;
        RECT 79.340 10.315 79.510 10.595 ;
        RECT 79.340 10.145 79.570 10.315 ;
        RECT 73.200 9.605 73.610 9.935 ;
        RECT 64.415 9.425 64.645 9.575 ;
        RECT 64.415 9.255 65.335 9.425 ;
        RECT 64.865 8.565 65.035 9.255 ;
        RECT 65.860 9.250 66.330 9.420 ;
        RECT 65.235 8.775 65.405 8.885 ;
        RECT 65.860 8.775 66.030 9.250 ;
        RECT 73.200 9.095 73.370 9.605 ;
        RECT 65.235 8.605 66.030 8.775 ;
        RECT 63.875 7.305 64.050 8.445 ;
        RECT 65.235 7.305 65.410 8.605 ;
        RECT 65.860 8.560 66.030 8.605 ;
        RECT 66.230 8.445 66.400 8.880 ;
        RECT 73.200 8.765 73.610 9.095 ;
        RECT 73.200 8.565 73.370 8.765 ;
        RECT 74.155 8.565 74.325 9.515 ;
        RECT 66.230 7.300 66.405 8.445 ;
        RECT 73.200 7.305 73.375 8.565 ;
        RECT 74.155 7.305 74.330 8.565 ;
        RECT 74.585 8.445 74.755 10.045 ;
        RECT 78.815 9.935 78.985 10.105 ;
        RECT 78.815 9.605 79.225 9.935 ;
        RECT 78.815 9.095 78.985 9.605 ;
        RECT 78.815 8.765 79.225 9.095 ;
        RECT 78.815 8.565 78.985 8.765 ;
        RECT 74.585 7.305 74.760 8.445 ;
        RECT 78.815 7.305 78.990 8.565 ;
        RECT 79.400 8.535 79.570 10.145 ;
        RECT 79.770 10.085 79.945 10.595 ;
        RECT 80.200 10.045 80.375 10.595 ;
        RECT 81.565 10.085 81.735 10.595 ;
        RECT 82.560 10.080 82.730 10.590 ;
        RECT 89.525 10.105 89.700 10.595 ;
        RECT 79.340 8.365 79.570 8.535 ;
        RECT 79.770 8.565 79.940 9.515 ;
        RECT 79.340 7.305 79.510 8.365 ;
        RECT 79.770 7.305 79.945 8.565 ;
        RECT 80.200 8.445 80.370 10.045 ;
        RECT 89.525 9.935 89.695 10.105 ;
        RECT 90.480 10.085 90.655 10.595 ;
        RECT 90.910 10.045 91.085 10.595 ;
        RECT 95.140 10.105 95.315 10.595 ;
        RECT 95.665 10.315 95.835 10.595 ;
        RECT 95.665 10.145 95.895 10.315 ;
        RECT 89.525 9.605 89.935 9.935 ;
        RECT 80.740 9.425 80.970 9.575 ;
        RECT 80.740 9.255 81.660 9.425 ;
        RECT 81.190 8.565 81.360 9.255 ;
        RECT 82.185 9.250 82.655 9.420 ;
        RECT 81.560 8.775 81.730 8.885 ;
        RECT 82.185 8.775 82.355 9.250 ;
        RECT 89.525 9.095 89.695 9.605 ;
        RECT 81.560 8.605 82.355 8.775 ;
        RECT 80.200 7.305 80.375 8.445 ;
        RECT 81.560 7.305 81.735 8.605 ;
        RECT 82.185 8.560 82.355 8.605 ;
        RECT 82.555 8.445 82.725 8.880 ;
        RECT 89.525 8.765 89.935 9.095 ;
        RECT 89.525 8.565 89.695 8.765 ;
        RECT 90.480 8.565 90.650 9.515 ;
        RECT 82.555 7.300 82.730 8.445 ;
        RECT 89.525 7.305 89.700 8.565 ;
        RECT 90.480 7.305 90.655 8.565 ;
        RECT 90.910 8.445 91.080 10.045 ;
        RECT 95.140 9.935 95.310 10.105 ;
        RECT 95.140 9.605 95.550 9.935 ;
        RECT 95.140 9.095 95.310 9.605 ;
        RECT 95.140 8.765 95.550 9.095 ;
        RECT 95.140 8.565 95.310 8.765 ;
        RECT 90.910 7.305 91.085 8.445 ;
        RECT 95.140 7.305 95.315 8.565 ;
        RECT 95.725 8.535 95.895 10.145 ;
        RECT 96.095 10.085 96.270 10.595 ;
        RECT 96.525 10.045 96.700 10.595 ;
        RECT 97.890 10.085 98.060 10.595 ;
        RECT 98.885 10.080 99.055 10.590 ;
        RECT 95.665 8.365 95.895 8.535 ;
        RECT 96.095 8.565 96.265 9.515 ;
        RECT 95.665 7.305 95.835 8.365 ;
        RECT 96.095 7.305 96.270 8.565 ;
        RECT 96.525 8.445 96.695 10.045 ;
        RECT 97.065 9.425 97.295 9.575 ;
        RECT 97.065 9.255 97.985 9.425 ;
        RECT 97.515 8.565 97.685 9.255 ;
        RECT 98.510 9.250 98.980 9.420 ;
        RECT 97.885 8.775 98.055 8.885 ;
        RECT 98.510 8.775 98.680 9.250 ;
        RECT 97.885 8.605 98.680 8.775 ;
        RECT 96.525 7.305 96.700 8.445 ;
        RECT 97.885 7.305 98.060 8.605 ;
        RECT 98.510 8.560 98.680 8.605 ;
        RECT 98.880 8.445 99.050 8.880 ;
        RECT 98.880 7.300 99.055 8.445 ;
        RECT 19.225 4.795 19.515 4.965 ;
        RECT 18.865 4.235 19.035 4.655 ;
        RECT 19.225 3.925 19.395 4.795 ;
        RECT 20.545 4.515 20.955 4.685 ;
        RECT 19.025 3.755 19.395 3.925 ;
        RECT 19.585 4.235 20.235 4.405 ;
        RECT 20.785 4.325 20.955 4.515 ;
        RECT 21.305 4.235 21.475 4.655 ;
        RECT 21.665 4.515 21.955 4.685 ;
        RECT 19.585 3.675 19.755 4.235 ;
        RECT 20.065 3.675 20.235 4.005 ;
        RECT 21.665 3.925 21.835 4.515 ;
        RECT 22.745 4.325 22.915 4.685 ;
        RECT 25.185 4.665 25.355 4.995 ;
        RECT 26.185 4.665 26.355 4.995 ;
        RECT 23.665 4.495 24.955 4.575 ;
        RECT 25.585 4.495 25.915 4.575 ;
        RECT 23.665 4.405 25.915 4.495 ;
        RECT 27.065 4.405 27.395 4.575 ;
        RECT 24.705 4.325 25.835 4.405 ;
        RECT 26.305 4.235 27.315 4.405 ;
        RECT 20.465 3.755 20.955 3.925 ;
        RECT 21.465 3.755 21.835 3.925 ;
        RECT 20.785 3.675 20.955 3.755 ;
        RECT 22.025 3.675 22.195 4.005 ;
        RECT 22.505 3.675 22.675 4.125 ;
        RECT 22.905 3.755 24.235 3.925 ;
        RECT 23.985 3.675 24.155 3.755 ;
        RECT 24.465 3.675 24.635 4.005 ;
        RECT 24.945 3.675 25.115 4.125 ;
        RECT 26.305 4.005 26.475 4.235 ;
        RECT 26.305 3.755 26.595 4.005 ;
        RECT 26.425 3.675 26.595 3.755 ;
        RECT 26.905 3.675 27.075 4.005 ;
        RECT 29.840 3.895 30.015 5.155 ;
        RECT 30.365 4.095 30.535 5.155 ;
        RECT 30.365 3.925 30.595 4.095 ;
        RECT 29.840 3.695 30.010 3.895 ;
        RECT 22.985 3.525 23.155 3.565 ;
        RECT 22.985 3.355 23.475 3.525 ;
        RECT 25.425 3.395 25.835 3.565 ;
        RECT 19.345 2.935 19.515 3.285 ;
        RECT 20.305 2.935 20.475 3.285 ;
        RECT 21.785 2.935 21.955 3.285 ;
        RECT 23.745 2.935 23.915 3.285 ;
        RECT 25.665 2.935 25.835 3.395 ;
        RECT 29.840 3.365 30.250 3.695 ;
        RECT 26.185 2.935 26.355 3.285 ;
        RECT 27.145 3.185 27.315 3.285 ;
        RECT 27.145 3.015 27.875 3.185 ;
        RECT 29.840 2.855 30.010 3.365 ;
        RECT 29.840 2.525 30.250 2.855 ;
        RECT 29.840 2.355 30.010 2.525 ;
        RECT 29.840 1.865 30.015 2.355 ;
        RECT 30.425 2.315 30.595 3.925 ;
        RECT 30.795 3.895 30.970 5.155 ;
        RECT 31.225 4.015 31.400 5.155 ;
        RECT 30.795 2.945 30.965 3.895 ;
        RECT 31.225 2.415 31.395 4.015 ;
        RECT 32.585 4.010 32.760 5.155 ;
        RECT 35.550 4.795 35.840 4.965 ;
        RECT 35.190 4.235 35.360 4.655 ;
        RECT 32.215 3.205 32.385 3.895 ;
        RECT 32.585 3.795 32.755 4.010 ;
        RECT 35.550 3.925 35.720 4.795 ;
        RECT 36.870 4.515 37.280 4.685 ;
        RECT 33.205 3.795 33.375 3.900 ;
        RECT 32.585 3.625 33.375 3.795 ;
        RECT 35.350 3.755 35.720 3.925 ;
        RECT 35.910 4.235 36.560 4.405 ;
        RECT 37.110 4.325 37.280 4.515 ;
        RECT 37.630 4.235 37.800 4.655 ;
        RECT 37.990 4.515 38.280 4.685 ;
        RECT 35.910 3.675 36.080 4.235 ;
        RECT 36.390 3.675 36.560 4.005 ;
        RECT 37.990 3.925 38.160 4.515 ;
        RECT 39.070 4.325 39.240 4.685 ;
        RECT 41.510 4.665 41.680 4.995 ;
        RECT 42.510 4.665 42.680 4.995 ;
        RECT 39.990 4.495 41.280 4.575 ;
        RECT 41.910 4.495 42.240 4.575 ;
        RECT 39.990 4.405 42.240 4.495 ;
        RECT 43.390 4.405 43.720 4.575 ;
        RECT 41.030 4.325 42.160 4.405 ;
        RECT 42.630 4.235 43.640 4.405 ;
        RECT 36.790 3.755 37.280 3.925 ;
        RECT 37.790 3.755 38.160 3.925 ;
        RECT 37.110 3.675 37.280 3.755 ;
        RECT 38.350 3.675 38.520 4.005 ;
        RECT 38.830 3.675 39.000 4.125 ;
        RECT 39.230 3.755 40.560 3.925 ;
        RECT 40.310 3.675 40.480 3.755 ;
        RECT 40.790 3.675 40.960 4.005 ;
        RECT 41.270 3.675 41.440 4.125 ;
        RECT 42.630 4.005 42.800 4.235 ;
        RECT 42.630 3.755 42.920 4.005 ;
        RECT 42.750 3.675 42.920 3.755 ;
        RECT 43.230 3.675 43.400 4.005 ;
        RECT 46.165 3.895 46.340 5.155 ;
        RECT 46.690 4.095 46.860 5.155 ;
        RECT 46.690 3.925 46.920 4.095 ;
        RECT 46.165 3.695 46.335 3.895 ;
        RECT 32.585 3.575 32.755 3.625 ;
        RECT 33.205 3.210 33.375 3.625 ;
        RECT 39.310 3.525 39.480 3.565 ;
        RECT 39.310 3.355 39.800 3.525 ;
        RECT 41.750 3.395 42.160 3.565 ;
        RECT 31.765 3.035 32.685 3.205 ;
        RECT 33.205 3.040 33.675 3.210 ;
        RECT 31.765 2.885 31.995 3.035 ;
        RECT 35.670 2.935 35.840 3.285 ;
        RECT 36.630 2.935 36.800 3.285 ;
        RECT 38.110 2.935 38.280 3.285 ;
        RECT 40.070 2.935 40.240 3.285 ;
        RECT 41.990 2.935 42.160 3.395 ;
        RECT 46.165 3.365 46.575 3.695 ;
        RECT 42.510 2.935 42.680 3.285 ;
        RECT 43.470 3.185 43.640 3.285 ;
        RECT 43.470 3.015 44.200 3.185 ;
        RECT 46.165 2.855 46.335 3.365 ;
        RECT 46.165 2.525 46.575 2.855 ;
        RECT 30.365 2.145 30.595 2.315 ;
        RECT 30.365 1.865 30.535 2.145 ;
        RECT 30.795 1.865 30.970 2.375 ;
        RECT 31.225 1.865 31.400 2.415 ;
        RECT 32.590 1.865 32.760 2.375 ;
        RECT 46.165 2.355 46.335 2.525 ;
        RECT 46.165 1.865 46.340 2.355 ;
        RECT 46.750 2.315 46.920 3.925 ;
        RECT 47.120 3.895 47.295 5.155 ;
        RECT 47.550 4.015 47.725 5.155 ;
        RECT 47.120 2.945 47.290 3.895 ;
        RECT 47.550 2.415 47.720 4.015 ;
        RECT 48.910 4.010 49.085 5.155 ;
        RECT 51.875 4.795 52.165 4.965 ;
        RECT 51.515 4.235 51.685 4.655 ;
        RECT 48.540 3.205 48.710 3.895 ;
        RECT 48.910 3.795 49.080 4.010 ;
        RECT 51.875 3.925 52.045 4.795 ;
        RECT 53.195 4.515 53.605 4.685 ;
        RECT 49.530 3.795 49.700 3.900 ;
        RECT 48.910 3.625 49.700 3.795 ;
        RECT 51.675 3.755 52.045 3.925 ;
        RECT 52.235 4.235 52.885 4.405 ;
        RECT 53.435 4.325 53.605 4.515 ;
        RECT 53.955 4.235 54.125 4.655 ;
        RECT 54.315 4.515 54.605 4.685 ;
        RECT 52.235 3.675 52.405 4.235 ;
        RECT 52.715 3.675 52.885 4.005 ;
        RECT 54.315 3.925 54.485 4.515 ;
        RECT 55.395 4.325 55.565 4.685 ;
        RECT 57.835 4.665 58.005 4.995 ;
        RECT 58.835 4.665 59.005 4.995 ;
        RECT 56.315 4.495 57.605 4.575 ;
        RECT 58.235 4.495 58.565 4.575 ;
        RECT 56.315 4.405 58.565 4.495 ;
        RECT 59.715 4.405 60.045 4.575 ;
        RECT 57.355 4.325 58.485 4.405 ;
        RECT 58.955 4.235 59.965 4.405 ;
        RECT 53.115 3.755 53.605 3.925 ;
        RECT 54.115 3.755 54.485 3.925 ;
        RECT 53.435 3.675 53.605 3.755 ;
        RECT 54.675 3.675 54.845 4.005 ;
        RECT 55.155 3.675 55.325 4.125 ;
        RECT 55.555 3.755 56.885 3.925 ;
        RECT 56.635 3.675 56.805 3.755 ;
        RECT 57.115 3.675 57.285 4.005 ;
        RECT 57.595 3.675 57.765 4.125 ;
        RECT 58.955 4.005 59.125 4.235 ;
        RECT 58.955 3.755 59.245 4.005 ;
        RECT 59.075 3.675 59.245 3.755 ;
        RECT 59.555 3.675 59.725 4.005 ;
        RECT 62.490 3.895 62.665 5.155 ;
        RECT 63.015 4.095 63.185 5.155 ;
        RECT 63.015 3.925 63.245 4.095 ;
        RECT 62.490 3.695 62.660 3.895 ;
        RECT 48.910 3.575 49.080 3.625 ;
        RECT 49.530 3.210 49.700 3.625 ;
        RECT 55.635 3.525 55.805 3.565 ;
        RECT 55.635 3.355 56.125 3.525 ;
        RECT 58.075 3.395 58.485 3.565 ;
        RECT 48.090 3.035 49.010 3.205 ;
        RECT 49.530 3.040 50.000 3.210 ;
        RECT 48.090 2.885 48.320 3.035 ;
        RECT 51.995 2.935 52.165 3.285 ;
        RECT 52.955 2.935 53.125 3.285 ;
        RECT 54.435 2.935 54.605 3.285 ;
        RECT 56.395 2.935 56.565 3.285 ;
        RECT 58.315 2.935 58.485 3.395 ;
        RECT 62.490 3.365 62.900 3.695 ;
        RECT 58.835 2.935 59.005 3.285 ;
        RECT 59.795 3.185 59.965 3.285 ;
        RECT 59.795 3.015 60.525 3.185 ;
        RECT 62.490 2.855 62.660 3.365 ;
        RECT 62.490 2.525 62.900 2.855 ;
        RECT 46.690 2.145 46.920 2.315 ;
        RECT 46.690 1.865 46.860 2.145 ;
        RECT 47.120 1.865 47.295 2.375 ;
        RECT 47.550 1.865 47.725 2.415 ;
        RECT 48.915 1.865 49.085 2.375 ;
        RECT 62.490 2.355 62.660 2.525 ;
        RECT 62.490 1.865 62.665 2.355 ;
        RECT 63.075 2.315 63.245 3.925 ;
        RECT 63.445 3.895 63.620 5.155 ;
        RECT 63.875 4.015 64.050 5.155 ;
        RECT 63.445 2.945 63.615 3.895 ;
        RECT 63.875 2.415 64.045 4.015 ;
        RECT 65.235 4.010 65.410 5.155 ;
        RECT 68.200 4.795 68.490 4.965 ;
        RECT 67.840 4.235 68.010 4.655 ;
        RECT 64.865 3.205 65.035 3.895 ;
        RECT 65.235 3.795 65.405 4.010 ;
        RECT 68.200 3.925 68.370 4.795 ;
        RECT 69.520 4.515 69.930 4.685 ;
        RECT 65.855 3.795 66.025 3.900 ;
        RECT 65.235 3.625 66.025 3.795 ;
        RECT 68.000 3.755 68.370 3.925 ;
        RECT 68.560 4.235 69.210 4.405 ;
        RECT 69.760 4.325 69.930 4.515 ;
        RECT 70.280 4.235 70.450 4.655 ;
        RECT 70.640 4.515 70.930 4.685 ;
        RECT 68.560 3.675 68.730 4.235 ;
        RECT 69.040 3.675 69.210 4.005 ;
        RECT 70.640 3.925 70.810 4.515 ;
        RECT 71.720 4.325 71.890 4.685 ;
        RECT 74.160 4.665 74.330 4.995 ;
        RECT 75.160 4.665 75.330 4.995 ;
        RECT 72.640 4.495 73.930 4.575 ;
        RECT 74.560 4.495 74.890 4.575 ;
        RECT 72.640 4.405 74.890 4.495 ;
        RECT 76.040 4.405 76.370 4.575 ;
        RECT 73.680 4.325 74.810 4.405 ;
        RECT 75.280 4.235 76.290 4.405 ;
        RECT 69.440 3.755 69.930 3.925 ;
        RECT 70.440 3.755 70.810 3.925 ;
        RECT 69.760 3.675 69.930 3.755 ;
        RECT 71.000 3.675 71.170 4.005 ;
        RECT 71.480 3.675 71.650 4.125 ;
        RECT 71.880 3.755 73.210 3.925 ;
        RECT 72.960 3.675 73.130 3.755 ;
        RECT 73.440 3.675 73.610 4.005 ;
        RECT 73.920 3.675 74.090 4.125 ;
        RECT 75.280 4.005 75.450 4.235 ;
        RECT 75.280 3.755 75.570 4.005 ;
        RECT 75.400 3.675 75.570 3.755 ;
        RECT 75.880 3.675 76.050 4.005 ;
        RECT 78.815 3.895 78.990 5.155 ;
        RECT 79.340 4.095 79.510 5.155 ;
        RECT 79.340 3.925 79.570 4.095 ;
        RECT 78.815 3.695 78.985 3.895 ;
        RECT 65.235 3.575 65.405 3.625 ;
        RECT 65.855 3.210 66.025 3.625 ;
        RECT 71.960 3.525 72.130 3.565 ;
        RECT 71.960 3.355 72.450 3.525 ;
        RECT 74.400 3.395 74.810 3.565 ;
        RECT 64.415 3.035 65.335 3.205 ;
        RECT 65.855 3.040 66.325 3.210 ;
        RECT 64.415 2.885 64.645 3.035 ;
        RECT 68.320 2.935 68.490 3.285 ;
        RECT 69.280 2.935 69.450 3.285 ;
        RECT 70.760 2.935 70.930 3.285 ;
        RECT 72.720 2.935 72.890 3.285 ;
        RECT 74.640 2.935 74.810 3.395 ;
        RECT 78.815 3.365 79.225 3.695 ;
        RECT 75.160 2.935 75.330 3.285 ;
        RECT 76.120 3.185 76.290 3.285 ;
        RECT 76.120 3.015 76.850 3.185 ;
        RECT 78.815 2.855 78.985 3.365 ;
        RECT 78.815 2.525 79.225 2.855 ;
        RECT 63.015 2.145 63.245 2.315 ;
        RECT 63.015 1.865 63.185 2.145 ;
        RECT 63.445 1.865 63.620 2.375 ;
        RECT 63.875 1.865 64.050 2.415 ;
        RECT 65.240 1.865 65.410 2.375 ;
        RECT 78.815 2.355 78.985 2.525 ;
        RECT 78.815 1.865 78.990 2.355 ;
        RECT 79.400 2.315 79.570 3.925 ;
        RECT 79.770 3.895 79.945 5.155 ;
        RECT 80.200 4.015 80.375 5.155 ;
        RECT 79.770 2.945 79.940 3.895 ;
        RECT 80.200 2.415 80.370 4.015 ;
        RECT 81.560 4.010 81.735 5.155 ;
        RECT 84.525 4.795 84.815 4.965 ;
        RECT 84.165 4.235 84.335 4.655 ;
        RECT 81.190 3.205 81.360 3.895 ;
        RECT 81.560 3.795 81.730 4.010 ;
        RECT 84.525 3.925 84.695 4.795 ;
        RECT 85.845 4.515 86.255 4.685 ;
        RECT 82.180 3.795 82.350 3.900 ;
        RECT 81.560 3.625 82.350 3.795 ;
        RECT 84.325 3.755 84.695 3.925 ;
        RECT 84.885 4.235 85.535 4.405 ;
        RECT 86.085 4.325 86.255 4.515 ;
        RECT 86.605 4.235 86.775 4.655 ;
        RECT 86.965 4.515 87.255 4.685 ;
        RECT 84.885 3.675 85.055 4.235 ;
        RECT 85.365 3.675 85.535 4.005 ;
        RECT 86.965 3.925 87.135 4.515 ;
        RECT 88.045 4.325 88.215 4.685 ;
        RECT 90.485 4.665 90.655 4.995 ;
        RECT 91.485 4.665 91.655 4.995 ;
        RECT 88.965 4.495 90.255 4.575 ;
        RECT 90.885 4.495 91.215 4.575 ;
        RECT 88.965 4.405 91.215 4.495 ;
        RECT 92.365 4.405 92.695 4.575 ;
        RECT 90.005 4.325 91.135 4.405 ;
        RECT 91.605 4.235 92.615 4.405 ;
        RECT 85.765 3.755 86.255 3.925 ;
        RECT 86.765 3.755 87.135 3.925 ;
        RECT 86.085 3.675 86.255 3.755 ;
        RECT 87.325 3.675 87.495 4.005 ;
        RECT 87.805 3.675 87.975 4.125 ;
        RECT 88.205 3.755 89.535 3.925 ;
        RECT 89.285 3.675 89.455 3.755 ;
        RECT 89.765 3.675 89.935 4.005 ;
        RECT 90.245 3.675 90.415 4.125 ;
        RECT 91.605 4.005 91.775 4.235 ;
        RECT 91.605 3.755 91.895 4.005 ;
        RECT 91.725 3.675 91.895 3.755 ;
        RECT 92.205 3.675 92.375 4.005 ;
        RECT 95.140 3.895 95.315 5.155 ;
        RECT 95.665 4.095 95.835 5.155 ;
        RECT 95.665 3.925 95.895 4.095 ;
        RECT 95.140 3.695 95.310 3.895 ;
        RECT 81.560 3.575 81.730 3.625 ;
        RECT 82.180 3.210 82.350 3.625 ;
        RECT 88.285 3.525 88.455 3.565 ;
        RECT 88.285 3.355 88.775 3.525 ;
        RECT 90.725 3.395 91.135 3.565 ;
        RECT 80.740 3.035 81.660 3.205 ;
        RECT 82.180 3.040 82.650 3.210 ;
        RECT 80.740 2.885 80.970 3.035 ;
        RECT 84.645 2.935 84.815 3.285 ;
        RECT 85.605 2.935 85.775 3.285 ;
        RECT 87.085 2.935 87.255 3.285 ;
        RECT 89.045 2.935 89.215 3.285 ;
        RECT 90.965 2.935 91.135 3.395 ;
        RECT 95.140 3.365 95.550 3.695 ;
        RECT 91.485 2.935 91.655 3.285 ;
        RECT 92.445 3.185 92.615 3.285 ;
        RECT 92.445 3.015 93.175 3.185 ;
        RECT 95.140 2.855 95.310 3.365 ;
        RECT 95.140 2.525 95.550 2.855 ;
        RECT 79.340 2.145 79.570 2.315 ;
        RECT 79.340 1.865 79.510 2.145 ;
        RECT 79.770 1.865 79.945 2.375 ;
        RECT 80.200 1.865 80.375 2.415 ;
        RECT 81.565 1.865 81.735 2.375 ;
        RECT 95.140 2.355 95.310 2.525 ;
        RECT 95.140 1.865 95.315 2.355 ;
        RECT 95.725 2.315 95.895 3.925 ;
        RECT 96.095 3.895 96.270 5.155 ;
        RECT 96.525 4.015 96.700 5.155 ;
        RECT 96.095 2.945 96.265 3.895 ;
        RECT 96.525 2.415 96.695 4.015 ;
        RECT 97.885 4.010 98.060 5.155 ;
        RECT 97.515 3.205 97.685 3.895 ;
        RECT 97.885 3.795 98.055 4.010 ;
        RECT 98.505 3.795 98.675 3.900 ;
        RECT 97.885 3.625 98.675 3.795 ;
        RECT 97.885 3.575 98.055 3.625 ;
        RECT 98.505 3.210 98.675 3.625 ;
        RECT 97.065 3.035 97.985 3.205 ;
        RECT 98.505 3.040 98.975 3.210 ;
        RECT 97.065 2.885 97.295 3.035 ;
        RECT 95.665 2.145 95.895 2.315 ;
        RECT 95.665 1.865 95.835 2.145 ;
        RECT 96.095 1.865 96.270 2.375 ;
        RECT 96.525 1.865 96.700 2.415 ;
        RECT 97.890 1.865 98.060 2.375 ;
      LAYER met1 ;
        RECT 16.540 10.055 16.830 10.285 ;
        RECT 25.120 10.055 25.410 10.285 ;
        RECT 30.735 10.055 31.025 10.285 ;
        RECT 16.600 9.605 16.770 10.055 ;
        RECT 25.180 9.710 25.350 10.055 ;
        RECT 16.510 9.315 16.860 9.605 ;
        RECT 25.100 9.360 25.470 9.710 ;
        RECT 30.795 9.575 30.965 10.055 ;
        RECT 32.525 10.025 32.820 10.285 ;
        RECT 31.705 9.575 32.055 9.605 ;
        RECT 30.795 9.545 32.055 9.575 ;
        RECT 30.735 9.405 32.055 9.545 ;
        RECT 25.100 9.340 25.410 9.360 ;
        RECT 25.120 9.315 25.410 9.340 ;
        RECT 30.735 9.315 31.025 9.405 ;
        RECT 31.705 9.315 32.055 9.405 ;
        RECT 25.550 9.145 25.840 9.175 ;
        RECT 25.380 9.140 25.840 9.145 ;
        RECT 26.585 9.140 26.935 9.240 ;
        RECT 31.190 9.175 31.515 9.265 ;
        RECT 31.165 9.145 31.515 9.175 ;
        RECT 30.995 9.140 31.515 9.145 ;
        RECT 25.380 8.975 31.515 9.140 ;
        RECT 25.550 8.970 31.515 8.975 ;
        RECT 25.550 8.945 25.840 8.970 ;
        RECT 26.585 8.890 26.935 8.970 ;
        RECT 31.165 8.945 31.515 8.970 ;
        RECT 31.190 8.940 31.515 8.945 ;
        RECT 32.585 8.925 32.755 10.025 ;
        RECT 33.520 10.020 33.815 10.280 ;
        RECT 41.445 10.055 41.735 10.285 ;
        RECT 47.060 10.055 47.350 10.285 ;
        RECT 33.580 9.290 33.750 10.020 ;
        RECT 41.505 9.710 41.675 10.055 ;
        RECT 41.425 9.360 41.795 9.710 ;
        RECT 47.120 9.575 47.290 10.055 ;
        RECT 48.850 10.025 49.145 10.285 ;
        RECT 48.030 9.575 48.380 9.605 ;
        RECT 47.120 9.545 48.380 9.575 ;
        RECT 47.060 9.405 48.380 9.545 ;
        RECT 41.425 9.340 41.735 9.360 ;
        RECT 41.445 9.315 41.735 9.340 ;
        RECT 47.060 9.315 47.350 9.405 ;
        RECT 48.030 9.315 48.380 9.405 ;
        RECT 32.525 8.920 32.755 8.925 ;
        RECT 33.570 8.940 33.920 9.290 ;
        RECT 42.075 9.175 42.425 9.245 ;
        RECT 47.515 9.175 47.840 9.265 ;
        RECT 41.875 9.145 42.425 9.175 ;
        RECT 47.490 9.145 47.840 9.175 ;
        RECT 41.705 9.140 42.425 9.145 ;
        RECT 47.320 9.140 47.840 9.145 ;
        RECT 41.705 8.975 47.840 9.140 ;
        RECT 41.875 8.970 47.840 8.975 ;
        RECT 41.875 8.945 42.425 8.970 ;
        RECT 47.490 8.945 47.840 8.970 ;
        RECT 33.570 8.920 33.870 8.940 ;
        RECT 16.135 8.785 16.485 8.860 ;
        RECT 30.390 8.815 30.710 8.830 ;
        RECT 30.365 8.785 30.710 8.815 ;
        RECT 15.995 8.615 16.485 8.785 ;
        RECT 30.190 8.615 30.710 8.785 ;
        RECT 32.525 8.685 32.815 8.920 ;
        RECT 33.520 8.850 33.870 8.920 ;
        RECT 42.075 8.895 42.425 8.945 ;
        RECT 47.515 8.940 47.840 8.945 ;
        RECT 48.910 8.925 49.080 10.025 ;
        RECT 49.845 10.020 50.140 10.280 ;
        RECT 57.770 10.055 58.060 10.285 ;
        RECT 63.385 10.055 63.675 10.285 ;
        RECT 49.905 9.300 50.075 10.020 ;
        RECT 57.830 9.710 58.000 10.055 ;
        RECT 57.750 9.360 58.120 9.710 ;
        RECT 63.445 9.575 63.615 10.055 ;
        RECT 65.175 10.025 65.470 10.285 ;
        RECT 64.355 9.575 64.705 9.605 ;
        RECT 63.445 9.545 64.705 9.575 ;
        RECT 63.385 9.405 64.705 9.545 ;
        RECT 57.750 9.340 58.060 9.360 ;
        RECT 57.770 9.315 58.060 9.340 ;
        RECT 63.385 9.315 63.675 9.405 ;
        RECT 64.355 9.315 64.705 9.405 ;
        RECT 48.850 8.920 49.080 8.925 ;
        RECT 49.890 8.945 50.245 9.300 ;
        RECT 58.400 9.175 58.750 9.250 ;
        RECT 63.840 9.175 64.165 9.265 ;
        RECT 58.200 9.145 58.750 9.175 ;
        RECT 63.815 9.145 64.165 9.175 ;
        RECT 58.030 9.140 58.750 9.145 ;
        RECT 63.645 9.140 64.165 9.145 ;
        RECT 58.030 8.975 64.165 9.140 ;
        RECT 58.200 8.970 64.165 8.975 ;
        RECT 58.200 8.945 58.750 8.970 ;
        RECT 63.815 8.945 64.165 8.970 ;
        RECT 49.890 8.920 50.195 8.945 ;
        RECT 33.520 8.680 33.810 8.850 ;
        RECT 46.715 8.815 47.035 8.830 ;
        RECT 46.690 8.785 47.035 8.815 ;
        RECT 46.515 8.615 47.035 8.785 ;
        RECT 48.850 8.685 49.140 8.920 ;
        RECT 49.845 8.850 50.195 8.920 ;
        RECT 58.400 8.900 58.750 8.945 ;
        RECT 63.840 8.940 64.165 8.945 ;
        RECT 65.235 8.925 65.405 10.025 ;
        RECT 66.170 10.020 66.465 10.280 ;
        RECT 74.095 10.055 74.385 10.285 ;
        RECT 79.710 10.055 80.000 10.285 ;
        RECT 66.230 9.290 66.400 10.020 ;
        RECT 74.155 9.710 74.325 10.055 ;
        RECT 74.075 9.360 74.445 9.710 ;
        RECT 79.770 9.575 79.940 10.055 ;
        RECT 81.500 10.025 81.795 10.285 ;
        RECT 80.680 9.575 81.030 9.605 ;
        RECT 79.770 9.545 81.030 9.575 ;
        RECT 79.710 9.405 81.030 9.545 ;
        RECT 74.075 9.340 74.385 9.360 ;
        RECT 74.095 9.315 74.385 9.340 ;
        RECT 79.710 9.315 80.000 9.405 ;
        RECT 80.680 9.315 81.030 9.405 ;
        RECT 65.175 8.920 65.405 8.925 ;
        RECT 66.175 8.940 66.525 9.290 ;
        RECT 74.725 9.175 75.075 9.245 ;
        RECT 80.165 9.175 80.490 9.265 ;
        RECT 74.525 9.145 75.075 9.175 ;
        RECT 80.140 9.145 80.490 9.175 ;
        RECT 74.355 9.140 75.075 9.145 ;
        RECT 79.970 9.140 80.490 9.145 ;
        RECT 74.355 8.975 80.490 9.140 ;
        RECT 74.525 8.970 80.490 8.975 ;
        RECT 74.525 8.945 75.075 8.970 ;
        RECT 80.140 8.945 80.490 8.970 ;
        RECT 66.175 8.920 66.520 8.940 ;
        RECT 49.845 8.680 50.135 8.850 ;
        RECT 63.040 8.815 63.360 8.830 ;
        RECT 63.015 8.785 63.360 8.815 ;
        RECT 62.840 8.615 63.360 8.785 ;
        RECT 65.175 8.685 65.465 8.920 ;
        RECT 66.170 8.845 66.520 8.920 ;
        RECT 74.725 8.895 75.075 8.945 ;
        RECT 80.165 8.940 80.490 8.945 ;
        RECT 81.560 8.925 81.730 10.025 ;
        RECT 82.495 10.020 82.790 10.280 ;
        RECT 90.420 10.055 90.710 10.285 ;
        RECT 96.035 10.055 96.325 10.285 ;
        RECT 82.555 9.290 82.725 10.020 ;
        RECT 90.480 9.710 90.650 10.055 ;
        RECT 90.400 9.360 90.770 9.710 ;
        RECT 96.095 9.575 96.265 10.055 ;
        RECT 97.825 10.025 98.120 10.285 ;
        RECT 97.005 9.575 97.355 9.605 ;
        RECT 96.095 9.545 97.355 9.575 ;
        RECT 96.035 9.405 97.355 9.545 ;
        RECT 90.400 9.340 90.710 9.360 ;
        RECT 90.420 9.315 90.710 9.340 ;
        RECT 96.035 9.315 96.325 9.405 ;
        RECT 97.005 9.315 97.355 9.405 ;
        RECT 81.500 8.920 81.730 8.925 ;
        RECT 82.500 8.940 82.850 9.290 ;
        RECT 91.055 9.175 91.405 9.245 ;
        RECT 96.490 9.175 96.815 9.265 ;
        RECT 90.850 9.145 91.405 9.175 ;
        RECT 96.465 9.145 96.815 9.175 ;
        RECT 90.680 9.140 91.405 9.145 ;
        RECT 96.295 9.140 96.815 9.145 ;
        RECT 90.680 8.975 96.815 9.140 ;
        RECT 90.850 8.970 96.815 8.975 ;
        RECT 90.850 8.945 91.405 8.970 ;
        RECT 96.465 8.945 96.815 8.970 ;
        RECT 82.500 8.920 82.845 8.940 ;
        RECT 66.170 8.680 66.460 8.845 ;
        RECT 79.365 8.815 79.685 8.830 ;
        RECT 79.340 8.785 79.685 8.815 ;
        RECT 79.165 8.615 79.685 8.785 ;
        RECT 81.500 8.685 81.790 8.920 ;
        RECT 82.495 8.845 82.845 8.920 ;
        RECT 91.055 8.895 91.405 8.945 ;
        RECT 96.490 8.940 96.815 8.945 ;
        RECT 97.885 8.925 98.055 10.025 ;
        RECT 98.820 10.020 99.115 10.280 ;
        RECT 98.850 9.980 99.115 10.020 ;
        RECT 98.850 9.910 99.175 9.980 ;
        RECT 98.850 9.560 99.200 9.910 ;
        RECT 97.825 8.920 98.055 8.925 ;
        RECT 98.880 8.920 99.050 9.560 ;
        RECT 82.495 8.680 82.785 8.845 ;
        RECT 95.690 8.815 96.010 8.830 ;
        RECT 95.665 8.785 96.010 8.815 ;
        RECT 95.490 8.615 96.010 8.785 ;
        RECT 97.825 8.685 98.115 8.920 ;
        RECT 98.820 8.915 99.050 8.920 ;
        RECT 98.820 8.680 99.110 8.915 ;
        RECT 16.135 8.570 16.485 8.615 ;
        RECT 30.365 8.585 30.710 8.615 ;
        RECT 46.690 8.585 47.035 8.615 ;
        RECT 63.015 8.585 63.360 8.615 ;
        RECT 79.340 8.585 79.685 8.615 ;
        RECT 95.665 8.585 96.010 8.615 ;
        RECT 30.390 8.540 30.710 8.585 ;
        RECT 46.715 8.540 47.035 8.585 ;
        RECT 63.040 8.540 63.360 8.585 ;
        RECT 79.365 8.540 79.685 8.585 ;
        RECT 95.690 8.540 96.010 8.585 ;
        RECT 19.285 4.955 19.575 4.995 ;
        RECT 19.985 4.955 20.305 5.015 ;
        RECT 19.285 4.815 20.305 4.955 ;
        RECT 19.285 4.765 19.615 4.815 ;
        RECT 19.985 4.755 20.305 4.815 ;
        RECT 25.125 4.955 25.415 4.995 ;
        RECT 25.125 4.765 25.455 4.955 ;
        RECT 20.485 4.675 20.775 4.715 ;
        RECT 21.705 4.675 22.025 4.735 ;
        RECT 22.545 4.715 22.865 4.735 ;
        RECT 22.545 4.675 22.975 4.715 ;
        RECT 20.485 4.485 20.935 4.675 ;
        RECT 18.785 4.195 19.105 4.455 ;
        RECT 19.745 4.435 20.065 4.455 ;
        RECT 19.745 4.205 20.295 4.435 ;
        RECT 20.795 4.255 20.935 4.485 ;
        RECT 21.705 4.535 22.975 4.675 ;
        RECT 21.705 4.475 22.025 4.535 ;
        RECT 22.545 4.485 22.975 4.535 ;
        RECT 22.545 4.475 22.865 4.485 ;
        RECT 19.745 4.195 20.065 4.205 ;
        RECT 18.875 3.275 19.015 4.195 ;
        RECT 20.435 4.115 20.935 4.255 ;
        RECT 21.245 4.205 21.535 4.435 ;
        RECT 19.745 3.875 20.065 3.895 ;
        RECT 19.745 3.645 20.295 3.875 ;
        RECT 19.745 3.635 20.065 3.645 ;
        RECT 20.435 3.335 20.575 4.115 ;
        RECT 21.315 3.895 21.455 4.205 ;
        RECT 22.515 4.155 25.095 4.255 ;
        RECT 22.445 4.115 25.175 4.155 ;
        RECT 22.445 3.925 23.105 4.115 ;
        RECT 24.885 3.925 25.175 4.115 ;
        RECT 22.785 3.915 23.105 3.925 ;
        RECT 20.965 3.875 21.455 3.895 ;
        RECT 20.725 3.645 21.455 3.875 ;
        RECT 20.965 3.635 21.455 3.645 ;
        RECT 21.945 3.635 22.265 3.895 ;
        RECT 23.785 3.875 24.105 3.895 ;
        RECT 23.785 3.645 24.215 3.875 ;
        RECT 23.785 3.635 24.105 3.645 ;
        RECT 24.385 3.635 24.705 3.895 ;
        RECT 19.285 3.275 19.575 3.315 ;
        RECT 18.875 3.135 19.575 3.275 ;
        RECT 19.285 3.085 19.575 3.135 ;
        RECT 20.225 3.135 20.575 3.335 ;
        RECT 21.315 3.275 21.455 3.635 ;
        RECT 22.425 3.555 22.745 3.615 ;
        RECT 25.315 3.595 25.455 4.765 ;
        RECT 26.125 4.735 26.415 4.995 ;
        RECT 35.610 4.955 35.900 4.995 ;
        RECT 36.310 4.955 36.630 5.015 ;
        RECT 35.610 4.815 36.630 4.955 ;
        RECT 35.610 4.765 35.940 4.815 ;
        RECT 36.310 4.755 36.630 4.815 ;
        RECT 41.450 4.955 41.740 4.995 ;
        RECT 41.450 4.765 41.780 4.955 ;
        RECT 26.105 4.475 26.425 4.735 ;
        RECT 36.810 4.675 37.100 4.715 ;
        RECT 38.030 4.675 38.350 4.735 ;
        RECT 38.870 4.715 39.190 4.735 ;
        RECT 38.870 4.675 39.300 4.715 ;
        RECT 36.810 4.485 37.260 4.675 ;
        RECT 35.110 4.195 35.430 4.455 ;
        RECT 36.070 4.435 36.390 4.455 ;
        RECT 36.070 4.205 36.620 4.435 ;
        RECT 37.120 4.255 37.260 4.485 ;
        RECT 38.030 4.535 39.300 4.675 ;
        RECT 38.030 4.475 38.350 4.535 ;
        RECT 38.870 4.485 39.300 4.535 ;
        RECT 38.870 4.475 39.190 4.485 ;
        RECT 36.070 4.195 36.390 4.205 ;
        RECT 26.225 3.875 26.545 3.895 ;
        RECT 30.390 3.875 30.710 3.980 ;
        RECT 26.225 3.635 26.695 3.875 ;
        RECT 26.845 3.835 27.135 3.875 ;
        RECT 30.365 3.860 30.710 3.875 ;
        RECT 30.360 3.845 30.710 3.860 ;
        RECT 26.845 3.695 27.295 3.835 ;
        RECT 26.845 3.645 27.775 3.695 ;
        RECT 30.190 3.675 30.710 3.845 ;
        RECT 30.365 3.660 30.710 3.675 ;
        RECT 30.365 3.645 30.655 3.660 ;
        RECT 22.925 3.555 23.215 3.595 ;
        RECT 25.315 3.555 25.655 3.595 ;
        RECT 22.425 3.415 23.215 3.555 ;
        RECT 22.425 3.355 22.745 3.415 ;
        RECT 22.925 3.365 23.215 3.415 ;
        RECT 24.955 3.415 25.655 3.555 ;
        RECT 24.955 3.395 25.095 3.415 ;
        RECT 23.495 3.335 25.095 3.395 ;
        RECT 25.365 3.365 25.655 3.415 ;
        RECT 26.555 3.395 26.695 3.635 ;
        RECT 27.155 3.615 27.775 3.645 ;
        RECT 27.155 3.555 27.865 3.615 ;
        RECT 21.725 3.275 22.015 3.315 ;
        RECT 21.315 3.135 22.015 3.275 ;
        RECT 20.225 3.075 20.545 3.135 ;
        RECT 21.725 3.085 22.015 3.135 ;
        RECT 23.405 3.255 25.095 3.335 ;
        RECT 25.845 3.315 26.165 3.335 ;
        RECT 23.405 3.085 23.975 3.255 ;
        RECT 25.845 3.085 26.415 3.315 ;
        RECT 26.555 3.275 26.815 3.395 ;
        RECT 27.545 3.355 27.865 3.555 ;
        RECT 31.165 3.490 31.515 3.610 ;
        RECT 32.525 3.540 32.815 3.775 ;
        RECT 32.525 3.535 32.755 3.540 ;
        RECT 28.860 3.320 31.515 3.490 ;
        RECT 27.085 3.275 27.375 3.315 ;
        RECT 26.555 3.255 27.375 3.275 ;
        RECT 26.675 3.135 27.375 3.255 ;
        RECT 27.085 3.085 27.375 3.135 ;
        RECT 28.860 3.105 29.030 3.320 ;
        RECT 30.995 3.315 31.515 3.320 ;
        RECT 31.165 3.260 31.515 3.315 ;
        RECT 30.735 3.120 31.025 3.145 ;
        RECT 31.705 3.120 32.055 3.145 ;
        RECT 23.405 3.075 23.725 3.085 ;
        RECT 25.845 3.075 26.165 3.085 ;
        RECT 28.770 2.755 29.110 3.105 ;
        RECT 30.735 2.950 32.055 3.120 ;
        RECT 30.735 2.915 31.025 2.950 ;
        RECT 30.795 2.405 30.965 2.915 ;
        RECT 31.705 2.855 32.055 2.950 ;
        RECT 32.585 2.435 32.755 3.535 ;
        RECT 35.200 3.275 35.340 4.195 ;
        RECT 36.760 4.115 37.260 4.255 ;
        RECT 37.570 4.205 37.860 4.435 ;
        RECT 36.070 3.875 36.390 3.895 ;
        RECT 36.070 3.645 36.620 3.875 ;
        RECT 36.070 3.635 36.390 3.645 ;
        RECT 36.760 3.335 36.900 4.115 ;
        RECT 37.640 3.895 37.780 4.205 ;
        RECT 38.840 4.155 41.420 4.255 ;
        RECT 38.770 4.115 41.500 4.155 ;
        RECT 38.770 3.925 39.430 4.115 ;
        RECT 41.210 3.925 41.500 4.115 ;
        RECT 39.110 3.915 39.430 3.925 ;
        RECT 37.290 3.875 37.780 3.895 ;
        RECT 37.050 3.645 37.780 3.875 ;
        RECT 37.290 3.635 37.780 3.645 ;
        RECT 38.270 3.635 38.590 3.895 ;
        RECT 40.110 3.875 40.430 3.895 ;
        RECT 40.110 3.645 40.540 3.875 ;
        RECT 40.110 3.635 40.430 3.645 ;
        RECT 40.710 3.635 41.030 3.895 ;
        RECT 35.610 3.275 35.900 3.315 ;
        RECT 35.200 3.135 35.900 3.275 ;
        RECT 35.610 3.085 35.900 3.135 ;
        RECT 36.550 3.135 36.900 3.335 ;
        RECT 37.640 3.275 37.780 3.635 ;
        RECT 38.750 3.555 39.070 3.615 ;
        RECT 41.640 3.595 41.780 4.765 ;
        RECT 42.450 4.735 42.740 4.995 ;
        RECT 51.935 4.955 52.225 4.995 ;
        RECT 52.635 4.955 52.955 5.015 ;
        RECT 51.935 4.815 52.955 4.955 ;
        RECT 51.935 4.765 52.265 4.815 ;
        RECT 52.635 4.755 52.955 4.815 ;
        RECT 57.775 4.955 58.065 4.995 ;
        RECT 57.775 4.765 58.105 4.955 ;
        RECT 42.430 4.475 42.750 4.735 ;
        RECT 53.135 4.675 53.425 4.715 ;
        RECT 54.355 4.675 54.675 4.735 ;
        RECT 55.195 4.715 55.515 4.735 ;
        RECT 55.195 4.675 55.625 4.715 ;
        RECT 53.135 4.485 53.585 4.675 ;
        RECT 51.435 4.195 51.755 4.455 ;
        RECT 52.395 4.435 52.715 4.455 ;
        RECT 52.395 4.205 52.945 4.435 ;
        RECT 53.445 4.255 53.585 4.485 ;
        RECT 54.355 4.535 55.625 4.675 ;
        RECT 54.355 4.475 54.675 4.535 ;
        RECT 55.195 4.485 55.625 4.535 ;
        RECT 55.195 4.475 55.515 4.485 ;
        RECT 52.395 4.195 52.715 4.205 ;
        RECT 42.550 3.875 42.870 3.895 ;
        RECT 46.715 3.875 47.035 3.980 ;
        RECT 42.550 3.635 43.020 3.875 ;
        RECT 43.170 3.835 43.460 3.875 ;
        RECT 46.690 3.860 47.035 3.875 ;
        RECT 46.685 3.845 47.035 3.860 ;
        RECT 43.170 3.695 43.620 3.835 ;
        RECT 43.170 3.645 44.100 3.695 ;
        RECT 46.515 3.675 47.035 3.845 ;
        RECT 46.690 3.660 47.035 3.675 ;
        RECT 46.690 3.645 46.980 3.660 ;
        RECT 39.250 3.555 39.540 3.595 ;
        RECT 41.640 3.555 41.980 3.595 ;
        RECT 38.750 3.415 39.540 3.555 ;
        RECT 38.750 3.355 39.070 3.415 ;
        RECT 39.250 3.365 39.540 3.415 ;
        RECT 41.280 3.415 41.980 3.555 ;
        RECT 41.280 3.395 41.420 3.415 ;
        RECT 39.820 3.335 41.420 3.395 ;
        RECT 41.690 3.365 41.980 3.415 ;
        RECT 42.880 3.395 43.020 3.635 ;
        RECT 43.480 3.615 44.100 3.645 ;
        RECT 43.480 3.555 44.190 3.615 ;
        RECT 38.050 3.275 38.340 3.315 ;
        RECT 37.640 3.135 38.340 3.275 ;
        RECT 36.550 3.075 36.870 3.135 ;
        RECT 38.050 3.085 38.340 3.135 ;
        RECT 39.730 3.255 41.420 3.335 ;
        RECT 42.170 3.315 42.490 3.335 ;
        RECT 39.730 3.085 40.300 3.255 ;
        RECT 42.170 3.085 42.740 3.315 ;
        RECT 42.880 3.275 43.140 3.395 ;
        RECT 43.870 3.355 44.190 3.555 ;
        RECT 47.490 3.490 47.840 3.610 ;
        RECT 48.850 3.540 49.140 3.775 ;
        RECT 48.850 3.535 49.080 3.540 ;
        RECT 45.185 3.320 47.840 3.490 ;
        RECT 43.410 3.275 43.700 3.315 ;
        RECT 42.880 3.255 43.700 3.275 ;
        RECT 43.000 3.135 43.700 3.255 ;
        RECT 43.410 3.085 43.700 3.135 ;
        RECT 45.185 3.105 45.355 3.320 ;
        RECT 47.320 3.315 47.840 3.320 ;
        RECT 47.490 3.260 47.840 3.315 ;
        RECT 47.060 3.120 47.350 3.145 ;
        RECT 48.030 3.120 48.380 3.145 ;
        RECT 39.730 3.075 40.050 3.085 ;
        RECT 42.170 3.075 42.490 3.085 ;
        RECT 45.095 2.755 45.435 3.105 ;
        RECT 47.060 2.950 48.380 3.120 ;
        RECT 47.060 2.915 47.350 2.950 ;
        RECT 30.735 2.175 31.025 2.405 ;
        RECT 32.525 2.175 32.820 2.435 ;
        RECT 47.120 2.405 47.290 2.915 ;
        RECT 48.030 2.855 48.380 2.950 ;
        RECT 48.910 2.435 49.080 3.535 ;
        RECT 51.525 3.275 51.665 4.195 ;
        RECT 53.085 4.115 53.585 4.255 ;
        RECT 53.895 4.205 54.185 4.435 ;
        RECT 52.395 3.875 52.715 3.895 ;
        RECT 52.395 3.645 52.945 3.875 ;
        RECT 52.395 3.635 52.715 3.645 ;
        RECT 53.085 3.335 53.225 4.115 ;
        RECT 53.965 3.895 54.105 4.205 ;
        RECT 55.165 4.155 57.745 4.255 ;
        RECT 55.095 4.115 57.825 4.155 ;
        RECT 55.095 3.925 55.755 4.115 ;
        RECT 57.535 3.925 57.825 4.115 ;
        RECT 55.435 3.915 55.755 3.925 ;
        RECT 53.615 3.875 54.105 3.895 ;
        RECT 53.375 3.645 54.105 3.875 ;
        RECT 53.615 3.635 54.105 3.645 ;
        RECT 54.595 3.635 54.915 3.895 ;
        RECT 56.435 3.875 56.755 3.895 ;
        RECT 56.435 3.645 56.865 3.875 ;
        RECT 56.435 3.635 56.755 3.645 ;
        RECT 57.035 3.635 57.355 3.895 ;
        RECT 51.935 3.275 52.225 3.315 ;
        RECT 51.525 3.135 52.225 3.275 ;
        RECT 51.935 3.085 52.225 3.135 ;
        RECT 52.875 3.135 53.225 3.335 ;
        RECT 53.965 3.275 54.105 3.635 ;
        RECT 55.075 3.555 55.395 3.615 ;
        RECT 57.965 3.595 58.105 4.765 ;
        RECT 58.775 4.735 59.065 4.995 ;
        RECT 68.260 4.955 68.550 4.995 ;
        RECT 68.960 4.955 69.280 5.015 ;
        RECT 68.260 4.815 69.280 4.955 ;
        RECT 68.260 4.765 68.590 4.815 ;
        RECT 68.960 4.755 69.280 4.815 ;
        RECT 74.100 4.955 74.390 4.995 ;
        RECT 74.100 4.765 74.430 4.955 ;
        RECT 58.755 4.475 59.075 4.735 ;
        RECT 69.460 4.675 69.750 4.715 ;
        RECT 70.680 4.675 71.000 4.735 ;
        RECT 71.520 4.715 71.840 4.735 ;
        RECT 71.520 4.675 71.950 4.715 ;
        RECT 69.460 4.485 69.910 4.675 ;
        RECT 67.760 4.195 68.080 4.455 ;
        RECT 68.720 4.435 69.040 4.455 ;
        RECT 68.720 4.205 69.270 4.435 ;
        RECT 69.770 4.255 69.910 4.485 ;
        RECT 70.680 4.535 71.950 4.675 ;
        RECT 70.680 4.475 71.000 4.535 ;
        RECT 71.520 4.485 71.950 4.535 ;
        RECT 71.520 4.475 71.840 4.485 ;
        RECT 68.720 4.195 69.040 4.205 ;
        RECT 58.875 3.875 59.195 3.895 ;
        RECT 63.040 3.875 63.360 3.980 ;
        RECT 58.875 3.635 59.345 3.875 ;
        RECT 59.495 3.835 59.785 3.875 ;
        RECT 63.015 3.860 63.360 3.875 ;
        RECT 63.010 3.845 63.360 3.860 ;
        RECT 59.495 3.695 59.945 3.835 ;
        RECT 59.495 3.645 60.425 3.695 ;
        RECT 62.840 3.675 63.360 3.845 ;
        RECT 63.015 3.660 63.360 3.675 ;
        RECT 63.015 3.645 63.305 3.660 ;
        RECT 55.575 3.555 55.865 3.595 ;
        RECT 57.965 3.555 58.305 3.595 ;
        RECT 55.075 3.415 55.865 3.555 ;
        RECT 55.075 3.355 55.395 3.415 ;
        RECT 55.575 3.365 55.865 3.415 ;
        RECT 57.605 3.415 58.305 3.555 ;
        RECT 57.605 3.395 57.745 3.415 ;
        RECT 56.145 3.335 57.745 3.395 ;
        RECT 58.015 3.365 58.305 3.415 ;
        RECT 59.205 3.395 59.345 3.635 ;
        RECT 59.805 3.615 60.425 3.645 ;
        RECT 59.805 3.555 60.515 3.615 ;
        RECT 54.375 3.275 54.665 3.315 ;
        RECT 53.965 3.135 54.665 3.275 ;
        RECT 52.875 3.075 53.195 3.135 ;
        RECT 54.375 3.085 54.665 3.135 ;
        RECT 56.055 3.255 57.745 3.335 ;
        RECT 58.495 3.315 58.815 3.335 ;
        RECT 56.055 3.085 56.625 3.255 ;
        RECT 58.495 3.085 59.065 3.315 ;
        RECT 59.205 3.275 59.465 3.395 ;
        RECT 60.195 3.355 60.515 3.555 ;
        RECT 63.815 3.490 64.165 3.610 ;
        RECT 65.175 3.540 65.465 3.775 ;
        RECT 65.175 3.535 65.405 3.540 ;
        RECT 61.510 3.320 64.165 3.490 ;
        RECT 59.735 3.275 60.025 3.315 ;
        RECT 59.205 3.255 60.025 3.275 ;
        RECT 59.325 3.135 60.025 3.255 ;
        RECT 59.735 3.085 60.025 3.135 ;
        RECT 61.510 3.105 61.680 3.320 ;
        RECT 63.645 3.315 64.165 3.320 ;
        RECT 63.815 3.260 64.165 3.315 ;
        RECT 63.385 3.120 63.675 3.145 ;
        RECT 64.355 3.120 64.705 3.145 ;
        RECT 56.055 3.075 56.375 3.085 ;
        RECT 58.495 3.075 58.815 3.085 ;
        RECT 61.420 2.755 61.760 3.105 ;
        RECT 63.385 2.950 64.705 3.120 ;
        RECT 63.385 2.915 63.675 2.950 ;
        RECT 47.060 2.175 47.350 2.405 ;
        RECT 48.850 2.175 49.145 2.435 ;
        RECT 63.445 2.405 63.615 2.915 ;
        RECT 64.355 2.855 64.705 2.950 ;
        RECT 65.235 2.435 65.405 3.535 ;
        RECT 67.850 3.275 67.990 4.195 ;
        RECT 69.410 4.115 69.910 4.255 ;
        RECT 70.220 4.205 70.510 4.435 ;
        RECT 68.720 3.875 69.040 3.895 ;
        RECT 68.720 3.645 69.270 3.875 ;
        RECT 68.720 3.635 69.040 3.645 ;
        RECT 69.410 3.335 69.550 4.115 ;
        RECT 70.290 3.895 70.430 4.205 ;
        RECT 71.490 4.155 74.070 4.255 ;
        RECT 71.420 4.115 74.150 4.155 ;
        RECT 71.420 3.925 72.080 4.115 ;
        RECT 73.860 3.925 74.150 4.115 ;
        RECT 71.760 3.915 72.080 3.925 ;
        RECT 69.940 3.875 70.430 3.895 ;
        RECT 69.700 3.645 70.430 3.875 ;
        RECT 69.940 3.635 70.430 3.645 ;
        RECT 70.920 3.635 71.240 3.895 ;
        RECT 72.760 3.875 73.080 3.895 ;
        RECT 72.760 3.645 73.190 3.875 ;
        RECT 72.760 3.635 73.080 3.645 ;
        RECT 73.360 3.635 73.680 3.895 ;
        RECT 68.260 3.275 68.550 3.315 ;
        RECT 67.850 3.135 68.550 3.275 ;
        RECT 68.260 3.085 68.550 3.135 ;
        RECT 69.200 3.135 69.550 3.335 ;
        RECT 70.290 3.275 70.430 3.635 ;
        RECT 71.400 3.555 71.720 3.615 ;
        RECT 74.290 3.595 74.430 4.765 ;
        RECT 75.100 4.735 75.390 4.995 ;
        RECT 84.585 4.955 84.875 4.995 ;
        RECT 85.285 4.955 85.605 5.015 ;
        RECT 84.585 4.815 85.605 4.955 ;
        RECT 84.585 4.765 84.915 4.815 ;
        RECT 85.285 4.755 85.605 4.815 ;
        RECT 90.425 4.955 90.715 4.995 ;
        RECT 90.425 4.765 90.755 4.955 ;
        RECT 75.080 4.475 75.400 4.735 ;
        RECT 85.785 4.675 86.075 4.715 ;
        RECT 87.005 4.675 87.325 4.735 ;
        RECT 87.845 4.715 88.165 4.735 ;
        RECT 87.845 4.675 88.275 4.715 ;
        RECT 85.785 4.485 86.235 4.675 ;
        RECT 84.085 4.195 84.405 4.455 ;
        RECT 85.045 4.435 85.365 4.455 ;
        RECT 85.045 4.205 85.595 4.435 ;
        RECT 86.095 4.255 86.235 4.485 ;
        RECT 87.005 4.535 88.275 4.675 ;
        RECT 87.005 4.475 87.325 4.535 ;
        RECT 87.845 4.485 88.275 4.535 ;
        RECT 87.845 4.475 88.165 4.485 ;
        RECT 85.045 4.195 85.365 4.205 ;
        RECT 75.200 3.875 75.520 3.895 ;
        RECT 79.365 3.875 79.685 3.980 ;
        RECT 75.200 3.635 75.670 3.875 ;
        RECT 75.820 3.835 76.110 3.875 ;
        RECT 79.340 3.860 79.685 3.875 ;
        RECT 79.335 3.845 79.685 3.860 ;
        RECT 75.820 3.695 76.270 3.835 ;
        RECT 75.820 3.645 76.750 3.695 ;
        RECT 79.165 3.675 79.685 3.845 ;
        RECT 79.340 3.660 79.685 3.675 ;
        RECT 79.340 3.645 79.630 3.660 ;
        RECT 71.900 3.555 72.190 3.595 ;
        RECT 74.290 3.555 74.630 3.595 ;
        RECT 71.400 3.415 72.190 3.555 ;
        RECT 71.400 3.355 71.720 3.415 ;
        RECT 71.900 3.365 72.190 3.415 ;
        RECT 73.930 3.415 74.630 3.555 ;
        RECT 73.930 3.395 74.070 3.415 ;
        RECT 72.470 3.335 74.070 3.395 ;
        RECT 74.340 3.365 74.630 3.415 ;
        RECT 75.530 3.395 75.670 3.635 ;
        RECT 76.130 3.615 76.750 3.645 ;
        RECT 76.130 3.555 76.840 3.615 ;
        RECT 70.700 3.275 70.990 3.315 ;
        RECT 70.290 3.135 70.990 3.275 ;
        RECT 69.200 3.075 69.520 3.135 ;
        RECT 70.700 3.085 70.990 3.135 ;
        RECT 72.380 3.255 74.070 3.335 ;
        RECT 74.820 3.315 75.140 3.335 ;
        RECT 72.380 3.085 72.950 3.255 ;
        RECT 74.820 3.085 75.390 3.315 ;
        RECT 75.530 3.275 75.790 3.395 ;
        RECT 76.520 3.355 76.840 3.555 ;
        RECT 80.140 3.490 80.490 3.610 ;
        RECT 81.500 3.540 81.790 3.775 ;
        RECT 81.500 3.535 81.730 3.540 ;
        RECT 77.835 3.320 80.490 3.490 ;
        RECT 76.060 3.275 76.350 3.315 ;
        RECT 75.530 3.255 76.350 3.275 ;
        RECT 75.650 3.135 76.350 3.255 ;
        RECT 76.060 3.085 76.350 3.135 ;
        RECT 77.835 3.105 78.005 3.320 ;
        RECT 79.970 3.315 80.490 3.320 ;
        RECT 80.140 3.260 80.490 3.315 ;
        RECT 79.710 3.120 80.000 3.145 ;
        RECT 80.680 3.120 81.030 3.145 ;
        RECT 72.380 3.075 72.700 3.085 ;
        RECT 74.820 3.075 75.140 3.085 ;
        RECT 77.745 2.755 78.085 3.105 ;
        RECT 79.710 2.950 81.030 3.120 ;
        RECT 79.710 2.915 80.000 2.950 ;
        RECT 63.385 2.175 63.675 2.405 ;
        RECT 65.175 2.175 65.470 2.435 ;
        RECT 79.770 2.405 79.940 2.915 ;
        RECT 80.680 2.855 81.030 2.950 ;
        RECT 81.560 2.435 81.730 3.535 ;
        RECT 84.175 3.275 84.315 4.195 ;
        RECT 85.735 4.115 86.235 4.255 ;
        RECT 86.545 4.205 86.835 4.435 ;
        RECT 85.045 3.875 85.365 3.895 ;
        RECT 85.045 3.645 85.595 3.875 ;
        RECT 85.045 3.635 85.365 3.645 ;
        RECT 85.735 3.335 85.875 4.115 ;
        RECT 86.615 3.895 86.755 4.205 ;
        RECT 87.815 4.155 90.395 4.255 ;
        RECT 87.745 4.115 90.475 4.155 ;
        RECT 87.745 3.925 88.405 4.115 ;
        RECT 90.185 3.925 90.475 4.115 ;
        RECT 88.085 3.915 88.405 3.925 ;
        RECT 86.265 3.875 86.755 3.895 ;
        RECT 86.025 3.645 86.755 3.875 ;
        RECT 86.265 3.635 86.755 3.645 ;
        RECT 87.245 3.635 87.565 3.895 ;
        RECT 89.085 3.875 89.405 3.895 ;
        RECT 89.085 3.645 89.515 3.875 ;
        RECT 89.085 3.635 89.405 3.645 ;
        RECT 89.685 3.635 90.005 3.895 ;
        RECT 84.585 3.275 84.875 3.315 ;
        RECT 84.175 3.135 84.875 3.275 ;
        RECT 84.585 3.085 84.875 3.135 ;
        RECT 85.525 3.135 85.875 3.335 ;
        RECT 86.615 3.275 86.755 3.635 ;
        RECT 87.725 3.555 88.045 3.615 ;
        RECT 90.615 3.595 90.755 4.765 ;
        RECT 91.425 4.735 91.715 4.995 ;
        RECT 91.405 4.475 91.725 4.735 ;
        RECT 91.525 3.875 91.845 3.895 ;
        RECT 95.690 3.875 96.010 3.980 ;
        RECT 91.525 3.635 91.995 3.875 ;
        RECT 92.145 3.835 92.435 3.875 ;
        RECT 95.665 3.860 96.010 3.875 ;
        RECT 95.660 3.845 96.010 3.860 ;
        RECT 92.145 3.695 92.595 3.835 ;
        RECT 92.145 3.645 93.075 3.695 ;
        RECT 95.490 3.675 96.010 3.845 ;
        RECT 95.665 3.660 96.010 3.675 ;
        RECT 95.665 3.645 95.955 3.660 ;
        RECT 88.225 3.555 88.515 3.595 ;
        RECT 90.615 3.555 90.955 3.595 ;
        RECT 87.725 3.415 88.515 3.555 ;
        RECT 87.725 3.355 88.045 3.415 ;
        RECT 88.225 3.365 88.515 3.415 ;
        RECT 90.255 3.415 90.955 3.555 ;
        RECT 90.255 3.395 90.395 3.415 ;
        RECT 88.795 3.335 90.395 3.395 ;
        RECT 90.665 3.365 90.955 3.415 ;
        RECT 91.855 3.395 91.995 3.635 ;
        RECT 92.455 3.615 93.075 3.645 ;
        RECT 92.455 3.555 93.165 3.615 ;
        RECT 87.025 3.275 87.315 3.315 ;
        RECT 86.615 3.135 87.315 3.275 ;
        RECT 85.525 3.075 85.845 3.135 ;
        RECT 87.025 3.085 87.315 3.135 ;
        RECT 88.705 3.255 90.395 3.335 ;
        RECT 91.145 3.315 91.465 3.335 ;
        RECT 88.705 3.085 89.275 3.255 ;
        RECT 91.145 3.085 91.715 3.315 ;
        RECT 91.855 3.275 92.115 3.395 ;
        RECT 92.845 3.355 93.165 3.555 ;
        RECT 96.465 3.490 96.815 3.610 ;
        RECT 97.825 3.540 98.115 3.775 ;
        RECT 97.825 3.535 98.055 3.540 ;
        RECT 94.160 3.320 96.815 3.490 ;
        RECT 92.385 3.275 92.675 3.315 ;
        RECT 91.855 3.255 92.675 3.275 ;
        RECT 91.975 3.135 92.675 3.255 ;
        RECT 92.385 3.085 92.675 3.135 ;
        RECT 94.160 3.105 94.330 3.320 ;
        RECT 96.295 3.315 96.815 3.320 ;
        RECT 96.465 3.260 96.815 3.315 ;
        RECT 96.035 3.120 96.325 3.145 ;
        RECT 97.005 3.120 97.355 3.145 ;
        RECT 88.705 3.075 89.025 3.085 ;
        RECT 91.145 3.075 91.465 3.085 ;
        RECT 94.070 2.755 94.410 3.105 ;
        RECT 96.035 2.950 97.355 3.120 ;
        RECT 96.035 2.915 96.325 2.950 ;
        RECT 79.710 2.175 80.000 2.405 ;
        RECT 81.500 2.175 81.795 2.435 ;
        RECT 96.095 2.405 96.265 2.915 ;
        RECT 97.005 2.855 97.355 2.950 ;
        RECT 97.885 2.435 98.055 3.535 ;
        RECT 96.035 2.175 96.325 2.405 ;
        RECT 97.825 2.175 98.120 2.435 ;
      LAYER met2 ;
        RECT 16.225 10.685 99.050 10.855 ;
        RECT 16.225 8.890 16.395 10.685 ;
        RECT 98.880 9.910 99.050 10.685 ;
        RECT 16.540 9.510 16.830 9.635 ;
        RECT 16.540 9.505 16.860 9.510 ;
        RECT 16.540 9.335 17.880 9.505 ;
        RECT 25.100 9.340 25.470 9.710 ;
        RECT 41.425 9.340 41.795 9.710 ;
        RECT 57.750 9.340 58.120 9.710 ;
        RECT 74.075 9.340 74.445 9.710 ;
        RECT 90.400 9.340 90.770 9.710 ;
        RECT 98.850 9.560 99.200 9.910 ;
        RECT 16.540 9.285 16.830 9.335 ;
        RECT 17.710 9.140 17.880 9.335 ;
        RECT 26.585 9.140 26.935 9.240 ;
        RECT 31.190 9.200 31.515 9.265 ;
        RECT 17.710 8.970 26.935 9.140 ;
        RECT 26.585 8.890 26.935 8.970 ;
        RECT 30.075 9.030 31.515 9.200 ;
        RECT 16.165 8.540 16.455 8.890 ;
        RECT 19.595 5.185 23.255 5.325 ;
        RECT 18.805 4.135 19.085 4.510 ;
        RECT 19.595 4.505 19.735 5.185 ;
        RECT 20.015 4.955 20.275 5.045 ;
        RECT 20.015 4.815 21.695 4.955 ;
        RECT 20.015 4.725 20.275 4.815 ;
        RECT 21.555 4.765 21.695 4.815 ;
        RECT 21.555 4.535 21.995 4.765 ;
        RECT 19.595 4.255 20.045 4.505 ;
        RECT 21.735 4.445 21.995 4.535 ;
        RECT 22.515 4.445 22.835 4.765 ;
        RECT 23.115 4.505 23.255 5.185 ;
        RECT 23.425 4.955 23.705 5.070 ;
        RECT 24.505 4.955 26.685 5.065 ;
        RECT 23.425 4.905 26.685 4.955 ;
        RECT 23.425 4.815 24.645 4.905 ;
        RECT 23.425 4.695 23.705 4.815 ;
        RECT 25.345 4.505 25.645 4.510 ;
        RECT 19.765 4.135 20.045 4.255 ;
        RECT 18.865 2.515 19.035 4.135 ;
        RECT 21.055 3.950 21.455 4.115 ;
        RECT 21.055 3.925 21.525 3.950 ;
        RECT 19.775 3.835 20.035 3.925 ;
        RECT 19.775 3.695 20.815 3.835 ;
        RECT 19.775 3.605 20.035 3.695 ;
        RECT 20.245 3.015 20.525 3.390 ;
        RECT 20.675 3.045 20.815 3.695 ;
        RECT 20.995 3.605 21.525 3.925 ;
        RECT 21.245 3.575 21.525 3.605 ;
        RECT 21.965 3.575 22.245 3.950 ;
        RECT 22.515 3.645 22.655 4.445 ;
        RECT 23.115 4.395 25.645 4.505 ;
        RECT 26.135 4.445 26.395 4.765 ;
        RECT 26.135 4.395 26.335 4.445 ;
        RECT 23.115 4.365 26.335 4.395 ;
        RECT 25.365 4.255 26.335 4.365 ;
        RECT 22.815 4.115 23.075 4.205 ;
        RECT 25.365 4.135 25.645 4.255 ;
        RECT 22.815 3.950 23.135 4.115 ;
        RECT 22.815 3.885 23.205 3.950 ;
        RECT 22.455 3.325 22.715 3.645 ;
        RECT 22.925 3.575 23.205 3.885 ;
        RECT 23.805 3.575 24.085 3.950 ;
        RECT 24.415 3.605 24.675 3.925 ;
        RECT 23.435 3.045 23.695 3.365 ;
        RECT 20.675 2.905 23.635 3.045 ;
        RECT 24.475 2.905 24.615 3.605 ;
        RECT 25.485 3.575 25.765 3.945 ;
        RECT 25.555 2.905 25.695 3.575 ;
        RECT 25.935 3.365 26.075 4.255 ;
        RECT 26.535 3.925 26.685 4.905 ;
        RECT 26.255 3.785 26.685 3.925 ;
        RECT 30.075 3.860 30.235 9.030 ;
        RECT 31.190 8.940 31.515 9.030 ;
        RECT 33.570 9.170 33.920 9.290 ;
        RECT 42.075 9.170 42.425 9.245 ;
        RECT 47.515 9.200 47.840 9.265 ;
        RECT 33.570 8.970 42.425 9.170 ;
        RECT 33.570 8.940 33.920 8.970 ;
        RECT 42.075 8.895 42.425 8.970 ;
        RECT 46.400 9.030 47.840 9.200 ;
        RECT 30.390 8.505 30.710 8.830 ;
        RECT 30.420 8.330 30.590 8.505 ;
        RECT 30.420 8.155 30.595 8.330 ;
        RECT 30.420 7.980 31.395 8.155 ;
        RECT 30.390 3.860 30.710 3.980 ;
        RECT 26.255 3.605 26.515 3.785 ;
        RECT 26.965 3.555 27.245 3.785 ;
        RECT 30.075 3.690 30.710 3.860 ;
        RECT 30.390 3.660 30.710 3.690 ;
        RECT 27.575 3.555 27.835 3.645 ;
        RECT 31.220 3.610 31.395 7.980 ;
        RECT 35.920 5.185 39.580 5.325 ;
        RECT 35.130 4.135 35.410 4.510 ;
        RECT 35.920 4.505 36.060 5.185 ;
        RECT 36.340 4.955 36.600 5.045 ;
        RECT 36.340 4.815 38.020 4.955 ;
        RECT 36.340 4.725 36.600 4.815 ;
        RECT 37.880 4.765 38.020 4.815 ;
        RECT 37.880 4.535 38.320 4.765 ;
        RECT 35.920 4.255 36.370 4.505 ;
        RECT 38.060 4.445 38.320 4.535 ;
        RECT 38.840 4.445 39.160 4.765 ;
        RECT 39.440 4.505 39.580 5.185 ;
        RECT 39.750 4.955 40.030 5.070 ;
        RECT 40.830 4.955 43.010 5.065 ;
        RECT 39.750 4.905 43.010 4.955 ;
        RECT 39.750 4.815 40.970 4.905 ;
        RECT 39.750 4.695 40.030 4.815 ;
        RECT 41.670 4.505 41.970 4.510 ;
        RECT 36.090 4.135 36.370 4.255 ;
        RECT 26.675 3.415 27.835 3.555 ;
        RECT 25.875 3.045 26.135 3.365 ;
        RECT 26.675 2.905 26.815 3.415 ;
        RECT 27.575 3.325 27.835 3.415 ;
        RECT 31.165 3.260 31.515 3.610 ;
        RECT 28.860 3.105 29.030 3.110 ;
        RECT 24.475 2.765 26.815 2.905 ;
        RECT 28.770 2.755 29.110 3.105 ;
        RECT 28.770 2.515 29.030 2.755 ;
        RECT 18.865 2.355 29.030 2.515 ;
        RECT 35.190 2.515 35.360 4.135 ;
        RECT 37.380 3.950 37.780 4.115 ;
        RECT 37.380 3.925 37.850 3.950 ;
        RECT 36.100 3.835 36.360 3.925 ;
        RECT 36.100 3.695 37.140 3.835 ;
        RECT 36.100 3.605 36.360 3.695 ;
        RECT 36.570 3.015 36.850 3.390 ;
        RECT 37.000 3.045 37.140 3.695 ;
        RECT 37.320 3.605 37.850 3.925 ;
        RECT 37.570 3.575 37.850 3.605 ;
        RECT 38.290 3.575 38.570 3.950 ;
        RECT 38.840 3.645 38.980 4.445 ;
        RECT 39.440 4.395 41.970 4.505 ;
        RECT 42.460 4.445 42.720 4.765 ;
        RECT 42.460 4.395 42.660 4.445 ;
        RECT 39.440 4.365 42.660 4.395 ;
        RECT 41.690 4.255 42.660 4.365 ;
        RECT 39.140 4.115 39.400 4.205 ;
        RECT 41.690 4.135 41.970 4.255 ;
        RECT 39.140 3.950 39.460 4.115 ;
        RECT 39.140 3.885 39.530 3.950 ;
        RECT 38.780 3.325 39.040 3.645 ;
        RECT 39.250 3.575 39.530 3.885 ;
        RECT 40.130 3.575 40.410 3.950 ;
        RECT 40.740 3.605 41.000 3.925 ;
        RECT 39.760 3.045 40.020 3.365 ;
        RECT 37.000 2.905 39.960 3.045 ;
        RECT 40.800 2.905 40.940 3.605 ;
        RECT 41.810 3.575 42.090 3.945 ;
        RECT 41.880 2.905 42.020 3.575 ;
        RECT 42.260 3.365 42.400 4.255 ;
        RECT 42.860 3.925 43.010 4.905 ;
        RECT 42.580 3.785 43.010 3.925 ;
        RECT 46.400 3.860 46.560 9.030 ;
        RECT 47.515 8.940 47.840 9.030 ;
        RECT 49.895 9.175 50.245 9.295 ;
        RECT 58.400 9.175 58.750 9.250 ;
        RECT 63.840 9.200 64.165 9.265 ;
        RECT 49.895 8.975 58.750 9.175 ;
        RECT 49.895 8.945 50.245 8.975 ;
        RECT 58.400 8.900 58.750 8.975 ;
        RECT 62.725 9.030 64.165 9.200 ;
        RECT 46.715 8.505 47.035 8.830 ;
        RECT 46.745 8.330 46.915 8.505 ;
        RECT 46.745 8.155 46.920 8.330 ;
        RECT 46.745 7.980 47.720 8.155 ;
        RECT 46.715 3.860 47.035 3.980 ;
        RECT 42.580 3.605 42.840 3.785 ;
        RECT 43.290 3.555 43.570 3.785 ;
        RECT 46.400 3.690 47.035 3.860 ;
        RECT 46.715 3.660 47.035 3.690 ;
        RECT 43.900 3.555 44.160 3.645 ;
        RECT 47.545 3.610 47.720 7.980 ;
        RECT 52.245 5.185 55.905 5.325 ;
        RECT 51.455 4.135 51.735 4.510 ;
        RECT 52.245 4.505 52.385 5.185 ;
        RECT 52.665 4.955 52.925 5.045 ;
        RECT 52.665 4.815 54.345 4.955 ;
        RECT 52.665 4.725 52.925 4.815 ;
        RECT 54.205 4.765 54.345 4.815 ;
        RECT 54.205 4.535 54.645 4.765 ;
        RECT 52.245 4.255 52.695 4.505 ;
        RECT 54.385 4.445 54.645 4.535 ;
        RECT 55.165 4.445 55.485 4.765 ;
        RECT 55.765 4.505 55.905 5.185 ;
        RECT 56.075 4.955 56.355 5.070 ;
        RECT 57.155 4.955 59.335 5.065 ;
        RECT 56.075 4.905 59.335 4.955 ;
        RECT 56.075 4.815 57.295 4.905 ;
        RECT 56.075 4.695 56.355 4.815 ;
        RECT 57.995 4.505 58.295 4.510 ;
        RECT 52.415 4.135 52.695 4.255 ;
        RECT 43.000 3.415 44.160 3.555 ;
        RECT 42.200 3.045 42.460 3.365 ;
        RECT 43.000 2.905 43.140 3.415 ;
        RECT 43.900 3.325 44.160 3.415 ;
        RECT 47.490 3.260 47.840 3.610 ;
        RECT 45.185 3.105 45.355 3.110 ;
        RECT 40.800 2.765 43.140 2.905 ;
        RECT 45.095 2.755 45.435 3.105 ;
        RECT 45.095 2.515 45.355 2.755 ;
        RECT 35.190 2.355 45.355 2.515 ;
        RECT 51.515 2.515 51.685 4.135 ;
        RECT 53.705 3.950 54.105 4.115 ;
        RECT 53.705 3.925 54.175 3.950 ;
        RECT 52.425 3.835 52.685 3.925 ;
        RECT 52.425 3.695 53.465 3.835 ;
        RECT 52.425 3.605 52.685 3.695 ;
        RECT 52.895 3.015 53.175 3.390 ;
        RECT 53.325 3.045 53.465 3.695 ;
        RECT 53.645 3.605 54.175 3.925 ;
        RECT 53.895 3.575 54.175 3.605 ;
        RECT 54.615 3.575 54.895 3.950 ;
        RECT 55.165 3.645 55.305 4.445 ;
        RECT 55.765 4.395 58.295 4.505 ;
        RECT 58.785 4.445 59.045 4.765 ;
        RECT 58.785 4.395 58.985 4.445 ;
        RECT 55.765 4.365 58.985 4.395 ;
        RECT 58.015 4.255 58.985 4.365 ;
        RECT 55.465 4.115 55.725 4.205 ;
        RECT 58.015 4.135 58.295 4.255 ;
        RECT 55.465 3.950 55.785 4.115 ;
        RECT 55.465 3.885 55.855 3.950 ;
        RECT 55.105 3.325 55.365 3.645 ;
        RECT 55.575 3.575 55.855 3.885 ;
        RECT 56.455 3.575 56.735 3.950 ;
        RECT 57.065 3.605 57.325 3.925 ;
        RECT 56.085 3.045 56.345 3.365 ;
        RECT 53.325 2.905 56.285 3.045 ;
        RECT 57.125 2.905 57.265 3.605 ;
        RECT 58.135 3.575 58.415 3.945 ;
        RECT 58.205 2.905 58.345 3.575 ;
        RECT 58.585 3.365 58.725 4.255 ;
        RECT 59.185 3.925 59.335 4.905 ;
        RECT 58.905 3.785 59.335 3.925 ;
        RECT 62.725 3.860 62.885 9.030 ;
        RECT 63.840 8.940 64.165 9.030 ;
        RECT 66.175 9.170 66.525 9.290 ;
        RECT 74.725 9.170 75.075 9.245 ;
        RECT 80.165 9.200 80.490 9.265 ;
        RECT 66.175 8.970 75.075 9.170 ;
        RECT 66.175 8.940 66.525 8.970 ;
        RECT 74.725 8.895 75.075 8.970 ;
        RECT 79.050 9.030 80.490 9.200 ;
        RECT 63.040 8.505 63.360 8.830 ;
        RECT 63.070 8.330 63.240 8.505 ;
        RECT 63.070 8.155 63.245 8.330 ;
        RECT 63.070 7.980 64.045 8.155 ;
        RECT 63.040 3.860 63.360 3.980 ;
        RECT 58.905 3.605 59.165 3.785 ;
        RECT 59.615 3.555 59.895 3.785 ;
        RECT 62.725 3.690 63.360 3.860 ;
        RECT 63.040 3.660 63.360 3.690 ;
        RECT 60.225 3.555 60.485 3.645 ;
        RECT 63.870 3.610 64.045 7.980 ;
        RECT 68.570 5.185 72.230 5.325 ;
        RECT 67.780 4.135 68.060 4.510 ;
        RECT 68.570 4.505 68.710 5.185 ;
        RECT 68.990 4.955 69.250 5.045 ;
        RECT 68.990 4.815 70.670 4.955 ;
        RECT 68.990 4.725 69.250 4.815 ;
        RECT 70.530 4.765 70.670 4.815 ;
        RECT 70.530 4.535 70.970 4.765 ;
        RECT 68.570 4.255 69.020 4.505 ;
        RECT 70.710 4.445 70.970 4.535 ;
        RECT 71.490 4.445 71.810 4.765 ;
        RECT 72.090 4.505 72.230 5.185 ;
        RECT 72.400 4.955 72.680 5.070 ;
        RECT 73.480 4.955 75.660 5.065 ;
        RECT 72.400 4.905 75.660 4.955 ;
        RECT 72.400 4.815 73.620 4.905 ;
        RECT 72.400 4.695 72.680 4.815 ;
        RECT 74.320 4.505 74.620 4.510 ;
        RECT 68.740 4.135 69.020 4.255 ;
        RECT 59.325 3.415 60.485 3.555 ;
        RECT 58.525 3.045 58.785 3.365 ;
        RECT 59.325 2.905 59.465 3.415 ;
        RECT 60.225 3.325 60.485 3.415 ;
        RECT 63.815 3.260 64.165 3.610 ;
        RECT 61.510 3.105 61.680 3.110 ;
        RECT 57.125 2.765 59.465 2.905 ;
        RECT 61.420 2.755 61.760 3.105 ;
        RECT 61.420 2.515 61.680 2.755 ;
        RECT 51.515 2.355 61.680 2.515 ;
        RECT 67.840 2.515 68.010 4.135 ;
        RECT 70.030 3.950 70.430 4.115 ;
        RECT 70.030 3.925 70.500 3.950 ;
        RECT 68.750 3.835 69.010 3.925 ;
        RECT 68.750 3.695 69.790 3.835 ;
        RECT 68.750 3.605 69.010 3.695 ;
        RECT 69.220 3.015 69.500 3.390 ;
        RECT 69.650 3.045 69.790 3.695 ;
        RECT 69.970 3.605 70.500 3.925 ;
        RECT 70.220 3.575 70.500 3.605 ;
        RECT 70.940 3.575 71.220 3.950 ;
        RECT 71.490 3.645 71.630 4.445 ;
        RECT 72.090 4.395 74.620 4.505 ;
        RECT 75.110 4.445 75.370 4.765 ;
        RECT 75.110 4.395 75.310 4.445 ;
        RECT 72.090 4.365 75.310 4.395 ;
        RECT 74.340 4.255 75.310 4.365 ;
        RECT 71.790 4.115 72.050 4.205 ;
        RECT 74.340 4.135 74.620 4.255 ;
        RECT 71.790 3.950 72.110 4.115 ;
        RECT 71.790 3.885 72.180 3.950 ;
        RECT 71.430 3.325 71.690 3.645 ;
        RECT 71.900 3.575 72.180 3.885 ;
        RECT 72.780 3.575 73.060 3.950 ;
        RECT 73.390 3.605 73.650 3.925 ;
        RECT 72.410 3.045 72.670 3.365 ;
        RECT 69.650 2.905 72.610 3.045 ;
        RECT 73.450 2.905 73.590 3.605 ;
        RECT 74.460 3.575 74.740 3.945 ;
        RECT 74.530 2.905 74.670 3.575 ;
        RECT 74.910 3.365 75.050 4.255 ;
        RECT 75.510 3.925 75.660 4.905 ;
        RECT 75.230 3.785 75.660 3.925 ;
        RECT 79.050 3.860 79.210 9.030 ;
        RECT 80.165 8.940 80.490 9.030 ;
        RECT 82.500 9.170 82.850 9.290 ;
        RECT 91.055 9.170 91.405 9.245 ;
        RECT 96.490 9.200 96.815 9.265 ;
        RECT 82.500 8.970 91.405 9.170 ;
        RECT 82.500 8.940 82.850 8.970 ;
        RECT 91.055 8.895 91.405 8.970 ;
        RECT 95.375 9.030 96.815 9.200 ;
        RECT 79.365 8.505 79.685 8.830 ;
        RECT 79.395 8.330 79.565 8.505 ;
        RECT 79.395 8.155 79.570 8.330 ;
        RECT 79.395 7.980 80.370 8.155 ;
        RECT 79.365 3.860 79.685 3.980 ;
        RECT 75.230 3.605 75.490 3.785 ;
        RECT 75.940 3.555 76.220 3.785 ;
        RECT 79.050 3.690 79.685 3.860 ;
        RECT 79.365 3.660 79.685 3.690 ;
        RECT 76.550 3.555 76.810 3.645 ;
        RECT 80.195 3.610 80.370 7.980 ;
        RECT 84.895 5.185 88.555 5.325 ;
        RECT 84.105 4.135 84.385 4.510 ;
        RECT 84.895 4.505 85.035 5.185 ;
        RECT 85.315 4.955 85.575 5.045 ;
        RECT 85.315 4.815 86.995 4.955 ;
        RECT 85.315 4.725 85.575 4.815 ;
        RECT 86.855 4.765 86.995 4.815 ;
        RECT 86.855 4.535 87.295 4.765 ;
        RECT 84.895 4.255 85.345 4.505 ;
        RECT 87.035 4.445 87.295 4.535 ;
        RECT 87.815 4.445 88.135 4.765 ;
        RECT 88.415 4.505 88.555 5.185 ;
        RECT 88.725 4.955 89.005 5.070 ;
        RECT 89.805 4.955 91.985 5.065 ;
        RECT 88.725 4.905 91.985 4.955 ;
        RECT 88.725 4.815 89.945 4.905 ;
        RECT 88.725 4.695 89.005 4.815 ;
        RECT 90.645 4.505 90.945 4.510 ;
        RECT 85.065 4.135 85.345 4.255 ;
        RECT 75.650 3.415 76.810 3.555 ;
        RECT 74.850 3.045 75.110 3.365 ;
        RECT 75.650 2.905 75.790 3.415 ;
        RECT 76.550 3.325 76.810 3.415 ;
        RECT 80.140 3.260 80.490 3.610 ;
        RECT 77.835 3.105 78.005 3.110 ;
        RECT 73.450 2.765 75.790 2.905 ;
        RECT 77.745 2.755 78.085 3.105 ;
        RECT 77.745 2.515 78.005 2.755 ;
        RECT 67.840 2.355 78.005 2.515 ;
        RECT 84.165 2.515 84.335 4.135 ;
        RECT 86.355 3.950 86.755 4.115 ;
        RECT 86.355 3.925 86.825 3.950 ;
        RECT 85.075 3.835 85.335 3.925 ;
        RECT 85.075 3.695 86.115 3.835 ;
        RECT 85.075 3.605 85.335 3.695 ;
        RECT 85.545 3.015 85.825 3.390 ;
        RECT 85.975 3.045 86.115 3.695 ;
        RECT 86.295 3.605 86.825 3.925 ;
        RECT 86.545 3.575 86.825 3.605 ;
        RECT 87.265 3.575 87.545 3.950 ;
        RECT 87.815 3.645 87.955 4.445 ;
        RECT 88.415 4.395 90.945 4.505 ;
        RECT 91.435 4.445 91.695 4.765 ;
        RECT 91.435 4.395 91.635 4.445 ;
        RECT 88.415 4.365 91.635 4.395 ;
        RECT 90.665 4.255 91.635 4.365 ;
        RECT 88.115 4.115 88.375 4.205 ;
        RECT 90.665 4.135 90.945 4.255 ;
        RECT 88.115 3.950 88.435 4.115 ;
        RECT 88.115 3.885 88.505 3.950 ;
        RECT 87.755 3.325 88.015 3.645 ;
        RECT 88.225 3.575 88.505 3.885 ;
        RECT 89.105 3.575 89.385 3.950 ;
        RECT 89.715 3.605 89.975 3.925 ;
        RECT 88.735 3.045 88.995 3.365 ;
        RECT 85.975 2.905 88.935 3.045 ;
        RECT 89.775 2.905 89.915 3.605 ;
        RECT 90.785 3.575 91.065 3.945 ;
        RECT 90.855 2.905 90.995 3.575 ;
        RECT 91.235 3.365 91.375 4.255 ;
        RECT 91.835 3.925 91.985 4.905 ;
        RECT 91.555 3.785 91.985 3.925 ;
        RECT 95.375 3.860 95.535 9.030 ;
        RECT 96.490 8.940 96.815 9.030 ;
        RECT 95.690 8.505 96.010 8.830 ;
        RECT 95.720 8.330 95.890 8.505 ;
        RECT 95.720 8.155 95.895 8.330 ;
        RECT 95.720 7.980 96.695 8.155 ;
        RECT 95.690 3.860 96.010 3.980 ;
        RECT 91.555 3.605 91.815 3.785 ;
        RECT 92.265 3.555 92.545 3.785 ;
        RECT 95.375 3.690 96.010 3.860 ;
        RECT 95.690 3.660 96.010 3.690 ;
        RECT 92.875 3.555 93.135 3.645 ;
        RECT 96.520 3.610 96.695 7.980 ;
        RECT 91.975 3.415 93.135 3.555 ;
        RECT 91.175 3.045 91.435 3.365 ;
        RECT 91.975 2.905 92.115 3.415 ;
        RECT 92.875 3.325 93.135 3.415 ;
        RECT 96.465 3.260 96.815 3.610 ;
        RECT 94.160 3.105 94.330 3.110 ;
        RECT 89.775 2.765 92.115 2.905 ;
        RECT 94.070 2.755 94.410 3.105 ;
        RECT 94.070 2.515 94.330 2.755 ;
        RECT 84.165 2.355 94.330 2.515 ;
        RECT 28.805 2.350 29.030 2.355 ;
        RECT 45.130 2.350 45.355 2.355 ;
        RECT 61.455 2.350 61.680 2.355 ;
        RECT 77.780 2.350 78.005 2.355 ;
        RECT 94.105 2.350 94.330 2.355 ;
      LAYER met3 ;
        RECT 25.100 9.675 25.470 9.710 ;
        RECT 41.425 9.675 41.795 9.710 ;
        RECT 57.750 9.675 58.120 9.710 ;
        RECT 74.075 9.675 74.445 9.710 ;
        RECT 90.400 9.675 90.770 9.710 ;
        RECT 25.100 9.375 27.085 9.675 ;
        RECT 25.100 9.340 25.470 9.375 ;
        RECT 23.400 5.035 23.735 5.055 ;
        RECT 22.195 4.735 23.735 5.035 ;
        RECT 18.780 3.755 19.115 4.490 ;
        RECT 21.225 3.930 21.555 4.325 ;
        RECT 22.195 3.930 22.495 4.735 ;
        RECT 23.400 4.715 23.735 4.735 ;
        RECT 25.340 4.165 25.675 4.490 ;
        RECT 20.225 3.360 20.555 3.765 ;
        RECT 21.220 3.595 21.555 3.930 ;
        RECT 21.940 3.615 22.495 3.930 ;
        RECT 22.900 3.875 23.235 3.930 ;
        RECT 23.780 3.875 24.115 3.930 ;
        RECT 21.940 3.595 22.275 3.615 ;
        RECT 22.900 3.600 25.045 3.875 ;
        RECT 25.345 3.755 25.675 4.165 ;
        RECT 26.785 3.875 27.085 9.375 ;
        RECT 41.425 9.375 43.410 9.675 ;
        RECT 41.425 9.340 41.795 9.375 ;
        RECT 39.725 5.035 40.060 5.055 ;
        RECT 38.520 4.735 40.060 5.035 ;
        RECT 20.220 3.035 20.555 3.360 ;
        RECT 22.905 3.575 25.045 3.600 ;
        RECT 22.905 3.195 23.235 3.575 ;
        RECT 23.785 3.195 24.115 3.575 ;
        RECT 24.745 3.455 25.045 3.575 ;
        RECT 25.985 3.575 27.275 3.875 ;
        RECT 35.105 3.755 35.440 4.490 ;
        RECT 37.550 3.930 37.880 4.325 ;
        RECT 38.520 3.930 38.820 4.735 ;
        RECT 39.725 4.715 40.060 4.735 ;
        RECT 41.665 4.165 42.000 4.490 ;
        RECT 25.985 3.455 26.290 3.575 ;
        RECT 24.745 3.155 26.290 3.455 ;
        RECT 26.940 3.415 27.275 3.575 ;
        RECT 26.945 3.035 27.275 3.415 ;
        RECT 36.550 3.360 36.880 3.765 ;
        RECT 37.545 3.595 37.880 3.930 ;
        RECT 38.265 3.615 38.820 3.930 ;
        RECT 39.225 3.875 39.560 3.930 ;
        RECT 40.105 3.875 40.440 3.930 ;
        RECT 38.265 3.595 38.600 3.615 ;
        RECT 39.225 3.600 41.370 3.875 ;
        RECT 41.670 3.755 42.000 4.165 ;
        RECT 43.110 3.875 43.410 9.375 ;
        RECT 57.750 9.375 59.735 9.675 ;
        RECT 57.750 9.340 58.120 9.375 ;
        RECT 56.050 5.035 56.385 5.055 ;
        RECT 54.845 4.735 56.385 5.035 ;
        RECT 36.545 3.035 36.880 3.360 ;
        RECT 39.230 3.575 41.370 3.600 ;
        RECT 39.230 3.195 39.560 3.575 ;
        RECT 40.110 3.195 40.440 3.575 ;
        RECT 41.070 3.455 41.370 3.575 ;
        RECT 42.310 3.575 43.600 3.875 ;
        RECT 51.430 3.755 51.765 4.490 ;
        RECT 53.875 3.930 54.205 4.325 ;
        RECT 54.845 3.930 55.145 4.735 ;
        RECT 56.050 4.715 56.385 4.735 ;
        RECT 57.990 4.165 58.325 4.490 ;
        RECT 42.310 3.455 42.615 3.575 ;
        RECT 41.070 3.155 42.615 3.455 ;
        RECT 43.265 3.415 43.600 3.575 ;
        RECT 43.270 3.035 43.600 3.415 ;
        RECT 52.875 3.360 53.205 3.765 ;
        RECT 53.870 3.595 54.205 3.930 ;
        RECT 54.590 3.615 55.145 3.930 ;
        RECT 55.550 3.875 55.885 3.930 ;
        RECT 56.430 3.875 56.765 3.930 ;
        RECT 54.590 3.595 54.925 3.615 ;
        RECT 55.550 3.600 57.695 3.875 ;
        RECT 57.995 3.755 58.325 4.165 ;
        RECT 59.435 3.875 59.735 9.375 ;
        RECT 74.075 9.375 76.060 9.675 ;
        RECT 74.075 9.340 74.445 9.375 ;
        RECT 72.375 5.035 72.710 5.055 ;
        RECT 71.170 4.735 72.710 5.035 ;
        RECT 52.870 3.035 53.205 3.360 ;
        RECT 55.555 3.575 57.695 3.600 ;
        RECT 55.555 3.195 55.885 3.575 ;
        RECT 56.435 3.195 56.765 3.575 ;
        RECT 57.395 3.455 57.695 3.575 ;
        RECT 58.635 3.575 59.925 3.875 ;
        RECT 67.755 3.755 68.090 4.490 ;
        RECT 70.200 3.930 70.530 4.325 ;
        RECT 71.170 3.930 71.470 4.735 ;
        RECT 72.375 4.715 72.710 4.735 ;
        RECT 74.315 4.165 74.650 4.490 ;
        RECT 58.635 3.455 58.940 3.575 ;
        RECT 57.395 3.155 58.940 3.455 ;
        RECT 59.590 3.415 59.925 3.575 ;
        RECT 59.595 3.035 59.925 3.415 ;
        RECT 69.200 3.360 69.530 3.765 ;
        RECT 70.195 3.595 70.530 3.930 ;
        RECT 70.915 3.615 71.470 3.930 ;
        RECT 71.875 3.875 72.210 3.930 ;
        RECT 72.755 3.875 73.090 3.930 ;
        RECT 70.915 3.595 71.250 3.615 ;
        RECT 71.875 3.600 74.020 3.875 ;
        RECT 74.320 3.755 74.650 4.165 ;
        RECT 75.760 3.875 76.060 9.375 ;
        RECT 90.400 9.375 92.385 9.675 ;
        RECT 90.400 9.340 90.770 9.375 ;
        RECT 88.700 5.035 89.035 5.055 ;
        RECT 87.495 4.735 89.035 5.035 ;
        RECT 69.195 3.035 69.530 3.360 ;
        RECT 71.880 3.575 74.020 3.600 ;
        RECT 71.880 3.195 72.210 3.575 ;
        RECT 72.760 3.195 73.090 3.575 ;
        RECT 73.720 3.455 74.020 3.575 ;
        RECT 74.960 3.575 76.250 3.875 ;
        RECT 84.080 3.755 84.415 4.490 ;
        RECT 86.525 3.930 86.855 4.325 ;
        RECT 87.495 3.930 87.795 4.735 ;
        RECT 88.700 4.715 89.035 4.735 ;
        RECT 90.640 4.165 90.975 4.490 ;
        RECT 74.960 3.455 75.265 3.575 ;
        RECT 73.720 3.155 75.265 3.455 ;
        RECT 75.915 3.415 76.250 3.575 ;
        RECT 75.920 3.035 76.250 3.415 ;
        RECT 85.525 3.360 85.855 3.765 ;
        RECT 86.520 3.595 86.855 3.930 ;
        RECT 87.240 3.615 87.795 3.930 ;
        RECT 88.200 3.875 88.535 3.930 ;
        RECT 89.080 3.875 89.415 3.930 ;
        RECT 87.240 3.595 87.575 3.615 ;
        RECT 88.200 3.600 90.345 3.875 ;
        RECT 90.645 3.755 90.975 4.165 ;
        RECT 92.085 3.875 92.385 9.375 ;
        RECT 85.520 3.035 85.855 3.360 ;
        RECT 88.205 3.575 90.345 3.600 ;
        RECT 88.205 3.195 88.535 3.575 ;
        RECT 89.085 3.195 89.415 3.575 ;
        RECT 90.045 3.455 90.345 3.575 ;
        RECT 91.285 3.575 92.575 3.875 ;
        RECT 91.285 3.455 91.590 3.575 ;
        RECT 90.045 3.155 91.590 3.455 ;
        RECT 92.240 3.415 92.575 3.575 ;
        RECT 92.245 3.035 92.575 3.415 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r2
MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r2
  CLASS BLOCK ;
  FOREIGN sky130_osu_ring_oscillator_mpr2et_8_b0r2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.600 BY 12.465 ;
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 26.040 8.240 26.210 9.510 ;
        RECT 31.655 8.240 31.825 9.510 ;
        RECT 31.655 2.955 31.825 4.225 ;
      LAYER met1 ;
        RECT 25.950 8.410 26.300 8.495 ;
        RECT 31.575 8.410 31.915 8.485 ;
        RECT 25.950 8.380 26.440 8.410 ;
        RECT 31.575 8.405 32.055 8.410 ;
        RECT 31.560 8.380 32.060 8.405 ;
        RECT 25.950 8.235 32.060 8.380 ;
        RECT 25.950 8.210 31.915 8.235 ;
        RECT 25.950 8.145 26.300 8.210 ;
        RECT 31.575 8.135 31.915 8.210 ;
        RECT 31.585 4.225 31.925 4.350 ;
        RECT 31.585 4.055 32.055 4.225 ;
        RECT 31.585 4.000 31.925 4.055 ;
      LAYER met2 ;
        RECT 31.575 8.135 31.915 8.485 ;
        RECT 31.660 4.350 31.830 8.135 ;
        RECT 31.585 4.000 31.925 4.350 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 44.600 8.240 44.770 9.510 ;
        RECT 50.215 8.240 50.385 9.510 ;
        RECT 50.215 2.955 50.385 4.225 ;
      LAYER met1 ;
        RECT 44.510 8.410 44.860 8.495 ;
        RECT 50.135 8.410 50.475 8.485 ;
        RECT 44.510 8.380 45.000 8.410 ;
        RECT 50.135 8.405 50.615 8.410 ;
        RECT 50.120 8.380 50.620 8.405 ;
        RECT 44.510 8.235 50.620 8.380 ;
        RECT 44.510 8.210 50.475 8.235 ;
        RECT 44.510 8.145 44.860 8.210 ;
        RECT 50.135 8.135 50.475 8.210 ;
        RECT 50.145 4.225 50.485 4.350 ;
        RECT 50.145 4.055 50.615 4.225 ;
        RECT 50.145 4.000 50.485 4.055 ;
      LAYER met2 ;
        RECT 50.135 8.135 50.475 8.485 ;
        RECT 50.220 4.350 50.390 8.135 ;
        RECT 50.145 4.000 50.485 4.350 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 63.160 8.240 63.330 9.510 ;
        RECT 68.775 8.240 68.945 9.510 ;
        RECT 68.775 2.955 68.945 4.225 ;
      LAYER met1 ;
        RECT 63.070 8.410 63.420 8.495 ;
        RECT 68.695 8.410 69.035 8.485 ;
        RECT 63.070 8.380 63.560 8.410 ;
        RECT 68.695 8.405 69.175 8.410 ;
        RECT 68.680 8.380 69.180 8.405 ;
        RECT 63.070 8.235 69.180 8.380 ;
        RECT 63.070 8.210 69.035 8.235 ;
        RECT 63.070 8.145 63.420 8.210 ;
        RECT 68.695 8.135 69.035 8.210 ;
        RECT 68.705 4.225 69.045 4.350 ;
        RECT 68.705 4.055 69.175 4.225 ;
        RECT 68.705 4.000 69.045 4.055 ;
      LAYER met2 ;
        RECT 68.695 8.135 69.035 8.485 ;
        RECT 68.780 4.350 68.950 8.135 ;
        RECT 68.705 4.000 69.045 4.350 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 81.720 8.240 81.890 9.510 ;
        RECT 87.335 8.240 87.505 9.510 ;
        RECT 87.335 2.955 87.505 4.225 ;
      LAYER met1 ;
        RECT 81.630 8.410 81.980 8.495 ;
        RECT 87.255 8.410 87.595 8.485 ;
        RECT 81.630 8.380 82.120 8.410 ;
        RECT 87.255 8.405 87.735 8.410 ;
        RECT 87.240 8.380 87.740 8.405 ;
        RECT 81.630 8.235 87.740 8.380 ;
        RECT 81.630 8.210 87.595 8.235 ;
        RECT 81.630 8.145 81.980 8.210 ;
        RECT 87.255 8.135 87.595 8.210 ;
        RECT 87.265 4.225 87.605 4.350 ;
        RECT 87.265 4.055 87.735 4.225 ;
        RECT 87.265 4.000 87.605 4.055 ;
      LAYER met2 ;
        RECT 87.255 8.135 87.595 8.485 ;
        RECT 87.340 4.350 87.510 8.135 ;
        RECT 87.265 4.000 87.605 4.350 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 100.280 8.240 100.450 9.510 ;
        RECT 105.895 8.240 106.065 9.510 ;
        RECT 105.895 2.955 106.065 4.225 ;
      LAYER met1 ;
        RECT 100.190 8.410 100.540 8.495 ;
        RECT 105.815 8.410 106.155 8.485 ;
        RECT 100.190 8.380 100.680 8.410 ;
        RECT 105.815 8.405 106.295 8.410 ;
        RECT 105.800 8.380 106.300 8.405 ;
        RECT 100.190 8.235 106.300 8.380 ;
        RECT 100.190 8.210 106.155 8.235 ;
        RECT 100.190 8.145 100.540 8.210 ;
        RECT 105.815 8.135 106.155 8.210 ;
        RECT 105.825 4.225 106.165 4.350 ;
        RECT 105.825 4.055 106.295 4.225 ;
        RECT 105.825 4.000 106.165 4.055 ;
      LAYER met2 ;
        RECT 105.815 8.135 106.155 8.485 ;
        RECT 105.900 4.350 106.070 8.135 ;
        RECT 105.825 4.000 106.165 4.350 ;
    END
  END s5
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 35.810 4.015 35.985 5.160 ;
        RECT 35.810 3.580 35.980 4.015 ;
        RECT 35.815 1.870 35.985 2.380 ;
      LAYER met1 ;
        RECT 35.750 3.545 36.040 3.780 ;
        RECT 35.750 3.540 35.980 3.545 ;
        RECT 35.810 2.440 35.980 3.540 ;
        RECT 35.750 2.180 36.045 2.440 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 54.370 4.015 54.545 5.160 ;
        RECT 54.370 3.580 54.540 4.015 ;
        RECT 54.375 1.870 54.545 2.380 ;
      LAYER met1 ;
        RECT 54.310 3.545 54.600 3.780 ;
        RECT 54.310 3.540 54.540 3.545 ;
        RECT 54.370 2.440 54.540 3.540 ;
        RECT 54.310 2.180 54.605 2.440 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 72.930 4.015 73.105 5.160 ;
        RECT 72.930 3.580 73.100 4.015 ;
        RECT 72.935 1.870 73.105 2.380 ;
      LAYER met1 ;
        RECT 72.870 3.545 73.160 3.780 ;
        RECT 72.870 3.540 73.100 3.545 ;
        RECT 72.930 2.440 73.100 3.540 ;
        RECT 72.870 2.180 73.165 2.440 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 91.490 4.015 91.665 5.160 ;
        RECT 91.490 3.580 91.660 4.015 ;
        RECT 91.495 1.870 91.665 2.380 ;
      LAYER met1 ;
        RECT 91.430 3.545 91.720 3.780 ;
        RECT 91.430 3.540 91.660 3.545 ;
        RECT 91.490 2.440 91.660 3.540 ;
        RECT 91.430 2.180 91.725 2.440 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 110.050 4.015 110.225 5.160 ;
        RECT 110.050 3.580 110.220 4.015 ;
        RECT 110.055 1.870 110.225 2.380 ;
      LAYER met1 ;
        RECT 109.990 3.545 110.280 3.780 ;
        RECT 109.990 3.540 110.220 3.545 ;
        RECT 110.050 2.440 110.220 3.540 ;
        RECT 109.990 2.180 110.285 2.440 ;
    END
  END X5_Y1
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 15.225 8.240 15.395 9.510 ;
      LAYER met1 ;
        RECT 15.140 8.410 15.480 8.455 ;
        RECT 15.140 8.240 15.625 8.410 ;
        RECT 15.140 8.195 15.480 8.240 ;
    END
  END start
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 10.865 110.600 12.465 ;
        RECT 15.215 10.240 15.385 10.865 ;
        RECT 26.030 10.240 26.200 10.865 ;
        RECT 26.985 10.320 27.155 10.600 ;
        RECT 26.985 10.150 27.215 10.320 ;
        RECT 31.645 10.240 31.815 10.865 ;
        RECT 34.390 10.240 34.560 10.865 ;
        RECT 35.385 10.235 35.555 10.865 ;
        RECT 44.590 10.240 44.760 10.865 ;
        RECT 45.545 10.320 45.715 10.600 ;
        RECT 45.545 10.150 45.775 10.320 ;
        RECT 50.205 10.240 50.375 10.865 ;
        RECT 52.950 10.240 53.120 10.865 ;
        RECT 53.945 10.235 54.115 10.865 ;
        RECT 63.150 10.240 63.320 10.865 ;
        RECT 64.105 10.320 64.275 10.600 ;
        RECT 64.105 10.150 64.335 10.320 ;
        RECT 68.765 10.240 68.935 10.865 ;
        RECT 71.510 10.240 71.680 10.865 ;
        RECT 72.505 10.235 72.675 10.865 ;
        RECT 81.710 10.240 81.880 10.865 ;
        RECT 82.665 10.320 82.835 10.600 ;
        RECT 82.665 10.150 82.895 10.320 ;
        RECT 87.325 10.240 87.495 10.865 ;
        RECT 90.070 10.240 90.240 10.865 ;
        RECT 91.065 10.235 91.235 10.865 ;
        RECT 100.270 10.240 100.440 10.865 ;
        RECT 101.225 10.320 101.395 10.600 ;
        RECT 101.225 10.150 101.455 10.320 ;
        RECT 105.885 10.240 106.055 10.865 ;
        RECT 108.630 10.240 108.800 10.865 ;
        RECT 109.625 10.235 109.795 10.865 ;
        RECT 27.045 8.540 27.215 10.150 ;
        RECT 45.605 8.540 45.775 10.150 ;
        RECT 64.165 8.540 64.335 10.150 ;
        RECT 82.725 8.540 82.895 10.150 ;
        RECT 101.285 8.540 101.455 10.150 ;
        RECT 26.985 8.370 27.215 8.540 ;
        RECT 45.545 8.370 45.775 8.540 ;
        RECT 64.105 8.370 64.335 8.540 ;
        RECT 82.665 8.370 82.895 8.540 ;
        RECT 101.225 8.370 101.455 8.540 ;
        RECT 26.985 7.310 27.155 8.370 ;
        RECT 45.545 7.310 45.715 8.370 ;
        RECT 64.105 7.310 64.275 8.370 ;
        RECT 82.665 7.310 82.835 8.370 ;
        RECT 101.225 7.310 101.395 8.370 ;
      LAYER met1 ;
        RECT 0.000 10.865 110.600 12.465 ;
        RECT 26.545 8.790 26.715 10.865 ;
        RECT 26.985 8.790 27.275 8.820 ;
        RECT 26.545 8.605 27.275 8.790 ;
        RECT 45.105 8.790 45.275 10.865 ;
        RECT 45.545 8.790 45.835 8.820 ;
        RECT 45.105 8.605 45.835 8.790 ;
        RECT 63.665 8.790 63.835 10.865 ;
        RECT 64.105 8.790 64.395 8.820 ;
        RECT 63.665 8.605 64.395 8.790 ;
        RECT 82.225 8.790 82.395 10.865 ;
        RECT 82.665 8.790 82.955 8.820 ;
        RECT 82.225 8.605 82.955 8.790 ;
        RECT 100.785 8.790 100.955 10.865 ;
        RECT 101.225 8.790 101.515 8.820 ;
        RECT 100.785 8.605 101.515 8.790 ;
        RECT 26.985 8.590 27.275 8.605 ;
        RECT 45.545 8.590 45.835 8.605 ;
        RECT 64.105 8.590 64.395 8.605 ;
        RECT 82.665 8.590 82.955 8.605 ;
        RECT 101.225 8.590 101.515 8.605 ;
    END
    PORT
      LAYER li1 ;
        RECT 20.190 4.345 20.480 4.515 ;
        RECT 38.750 4.345 39.040 4.515 ;
        RECT 57.310 4.345 57.600 4.515 ;
        RECT 75.870 4.345 76.160 4.515 ;
        RECT 94.430 4.345 94.720 4.515 ;
        RECT 20.190 4.035 20.360 4.345 ;
        RECT 19.990 3.865 20.360 4.035 ;
        RECT 22.030 3.785 22.200 4.115 ;
        RECT 38.750 4.035 38.920 4.345 ;
        RECT 38.550 3.865 38.920 4.035 ;
        RECT 40.590 3.785 40.760 4.115 ;
        RECT 57.310 4.035 57.480 4.345 ;
        RECT 57.110 3.865 57.480 4.035 ;
        RECT 59.150 3.785 59.320 4.115 ;
        RECT 75.870 4.035 76.040 4.345 ;
        RECT 75.670 3.865 76.040 4.035 ;
        RECT 77.710 3.785 77.880 4.115 ;
        RECT 94.430 4.035 94.600 4.345 ;
        RECT 94.230 3.865 94.600 4.035 ;
        RECT 96.270 3.785 96.440 4.115 ;
        RECT 19.350 2.875 19.520 3.375 ;
        RECT 20.830 2.890 21.000 3.375 ;
        RECT 20.830 2.875 21.090 2.890 ;
        RECT 22.750 2.875 22.920 3.375 ;
        RECT 23.195 2.875 23.390 2.890 ;
        RECT 24.230 2.875 24.400 3.375 ;
        RECT 25.190 2.875 25.360 3.375 ;
        RECT 26.190 2.875 26.360 3.375 ;
        RECT 27.150 2.875 27.320 3.375 ;
        RECT 27.670 2.875 27.840 3.375 ;
        RECT 28.630 2.875 28.800 3.375 ;
        RECT 29.590 2.875 29.760 3.375 ;
        RECT 30.395 2.875 30.585 2.880 ;
        RECT 37.910 2.875 38.080 3.375 ;
        RECT 39.390 2.890 39.560 3.375 ;
        RECT 39.390 2.875 39.650 2.890 ;
        RECT 41.310 2.875 41.480 3.375 ;
        RECT 41.755 2.875 41.950 2.890 ;
        RECT 42.790 2.875 42.960 3.375 ;
        RECT 43.750 2.875 43.920 3.375 ;
        RECT 44.750 2.875 44.920 3.375 ;
        RECT 45.710 2.875 45.880 3.375 ;
        RECT 46.230 2.875 46.400 3.375 ;
        RECT 47.190 2.875 47.360 3.375 ;
        RECT 48.150 2.875 48.320 3.375 ;
        RECT 48.955 2.875 49.145 2.880 ;
        RECT 56.470 2.875 56.640 3.375 ;
        RECT 57.950 2.890 58.120 3.375 ;
        RECT 57.950 2.875 58.210 2.890 ;
        RECT 59.870 2.875 60.040 3.375 ;
        RECT 60.315 2.875 60.510 2.890 ;
        RECT 61.350 2.875 61.520 3.375 ;
        RECT 62.310 2.875 62.480 3.375 ;
        RECT 63.310 2.875 63.480 3.375 ;
        RECT 64.270 2.875 64.440 3.375 ;
        RECT 64.790 2.875 64.960 3.375 ;
        RECT 65.750 2.875 65.920 3.375 ;
        RECT 66.710 2.875 66.880 3.375 ;
        RECT 67.515 2.875 67.705 2.880 ;
        RECT 75.030 2.875 75.200 3.375 ;
        RECT 76.510 2.890 76.680 3.375 ;
        RECT 76.510 2.875 76.770 2.890 ;
        RECT 78.430 2.875 78.600 3.375 ;
        RECT 78.875 2.875 79.070 2.890 ;
        RECT 79.910 2.875 80.080 3.375 ;
        RECT 80.870 2.875 81.040 3.375 ;
        RECT 81.870 2.875 82.040 3.375 ;
        RECT 82.830 2.875 83.000 3.375 ;
        RECT 83.350 2.875 83.520 3.375 ;
        RECT 84.310 2.875 84.480 3.375 ;
        RECT 85.270 2.875 85.440 3.375 ;
        RECT 86.075 2.875 86.265 2.880 ;
        RECT 93.590 2.875 93.760 3.375 ;
        RECT 95.070 2.890 95.240 3.375 ;
        RECT 95.070 2.875 95.330 2.890 ;
        RECT 96.990 2.875 97.160 3.375 ;
        RECT 97.435 2.875 97.630 2.890 ;
        RECT 98.470 2.875 98.640 3.375 ;
        RECT 99.430 2.875 99.600 3.375 ;
        RECT 100.430 2.875 100.600 3.375 ;
        RECT 101.390 2.875 101.560 3.375 ;
        RECT 101.910 2.875 102.080 3.375 ;
        RECT 102.870 2.875 103.040 3.375 ;
        RECT 103.830 2.875 104.000 3.375 ;
        RECT 104.635 2.875 104.825 2.880 ;
        RECT 18.540 1.600 30.585 2.875 ;
        RECT 31.645 1.600 31.815 2.225 ;
        RECT 34.390 1.600 34.560 2.225 ;
        RECT 35.380 1.600 35.550 2.230 ;
        RECT 37.100 1.600 49.145 2.875 ;
        RECT 50.205 1.600 50.375 2.225 ;
        RECT 52.950 1.600 53.120 2.225 ;
        RECT 53.940 1.600 54.110 2.230 ;
        RECT 55.660 1.600 67.705 2.875 ;
        RECT 68.765 1.600 68.935 2.225 ;
        RECT 71.510 1.600 71.680 2.225 ;
        RECT 72.500 1.600 72.670 2.230 ;
        RECT 74.220 1.600 86.265 2.875 ;
        RECT 87.325 1.600 87.495 2.225 ;
        RECT 90.070 1.600 90.240 2.225 ;
        RECT 91.060 1.600 91.230 2.230 ;
        RECT 92.780 1.600 104.825 2.875 ;
        RECT 105.885 1.600 106.055 2.225 ;
        RECT 108.630 1.600 108.800 2.225 ;
        RECT 109.620 1.600 109.790 2.230 ;
        RECT 0.000 0.000 110.595 1.600 ;
      LAYER met1 ;
        RECT 20.230 4.305 20.550 4.565 ;
        RECT 38.790 4.305 39.110 4.565 ;
        RECT 57.350 4.305 57.670 4.565 ;
        RECT 75.910 4.305 76.230 4.565 ;
        RECT 94.470 4.305 94.790 4.565 ;
        RECT 21.970 3.805 22.260 4.035 ;
        RECT 40.530 3.805 40.820 4.035 ;
        RECT 59.090 3.805 59.380 4.035 ;
        RECT 77.650 3.805 77.940 4.035 ;
        RECT 96.210 3.805 96.500 4.035 ;
        RECT 21.200 3.665 22.260 3.805 ;
        RECT 39.760 3.665 40.820 3.805 ;
        RECT 58.320 3.665 59.380 3.805 ;
        RECT 76.880 3.665 77.940 3.805 ;
        RECT 95.440 3.665 96.500 3.805 ;
        RECT 18.540 2.880 30.500 2.905 ;
        RECT 37.100 2.880 49.060 2.905 ;
        RECT 55.660 2.880 67.620 2.905 ;
        RECT 74.220 2.880 86.180 2.905 ;
        RECT 92.780 2.880 104.740 2.905 ;
        RECT 18.540 1.600 30.585 2.880 ;
        RECT 37.100 1.600 49.145 2.880 ;
        RECT 55.660 1.600 67.705 2.880 ;
        RECT 74.220 1.600 86.265 2.880 ;
        RECT 92.780 1.600 104.825 2.880 ;
        RECT 0.000 0.000 110.595 1.600 ;
      LAYER met2 ;
        RECT 20.260 4.505 20.520 4.595 ;
        RECT 38.820 4.505 39.080 4.595 ;
        RECT 57.380 4.505 57.640 4.595 ;
        RECT 75.940 4.505 76.200 4.595 ;
        RECT 94.500 4.505 94.760 4.595 ;
        RECT 20.200 4.275 20.520 4.505 ;
        RECT 38.760 4.275 39.080 4.505 ;
        RECT 57.320 4.275 57.640 4.505 ;
        RECT 75.880 4.275 76.200 4.505 ;
        RECT 94.440 4.275 94.760 4.505 ;
        RECT 20.200 3.945 20.340 4.275 ;
        RECT 20.510 3.945 20.790 4.060 ;
        RECT 21.980 3.945 22.240 4.035 ;
        RECT 20.200 3.805 22.240 3.945 ;
        RECT 38.760 3.945 38.900 4.275 ;
        RECT 39.070 3.945 39.350 4.060 ;
        RECT 40.540 3.945 40.800 4.035 ;
        RECT 38.760 3.805 40.800 3.945 ;
        RECT 57.320 3.945 57.460 4.275 ;
        RECT 57.630 3.945 57.910 4.060 ;
        RECT 59.100 3.945 59.360 4.035 ;
        RECT 57.320 3.805 59.360 3.945 ;
        RECT 75.880 3.945 76.020 4.275 ;
        RECT 76.190 3.945 76.470 4.060 ;
        RECT 77.660 3.945 77.920 4.035 ;
        RECT 75.880 3.805 77.920 3.945 ;
        RECT 94.440 3.945 94.580 4.275 ;
        RECT 94.750 3.945 95.030 4.060 ;
        RECT 96.220 3.945 96.480 4.035 ;
        RECT 94.440 3.805 96.480 3.945 ;
        RECT 20.510 3.685 20.790 3.805 ;
        RECT 21.980 3.715 22.240 3.805 ;
        RECT 39.070 3.685 39.350 3.805 ;
        RECT 40.540 3.715 40.800 3.805 ;
        RECT 57.630 3.685 57.910 3.805 ;
        RECT 59.100 3.715 59.360 3.805 ;
        RECT 76.190 3.685 76.470 3.805 ;
        RECT 77.660 3.715 77.920 3.805 ;
        RECT 94.750 3.685 95.030 3.805 ;
        RECT 96.220 3.715 96.480 3.805 ;
        RECT 20.610 2.635 20.780 3.685 ;
        RECT 39.170 2.635 39.340 3.685 ;
        RECT 57.730 2.635 57.900 3.685 ;
        RECT 76.290 2.635 76.460 3.685 ;
        RECT 94.850 2.635 95.020 3.685 ;
        RECT 20.585 2.295 20.925 2.635 ;
        RECT 39.145 2.295 39.485 2.635 ;
        RECT 57.705 2.295 58.045 2.635 ;
        RECT 76.265 2.295 76.605 2.635 ;
        RECT 94.825 2.295 95.165 2.635 ;
      LAYER met3 ;
        RECT 20.490 4.035 20.815 4.040 ;
        RECT 39.050 4.035 39.375 4.040 ;
        RECT 57.610 4.035 57.935 4.040 ;
        RECT 76.170 4.035 76.495 4.040 ;
        RECT 94.730 4.035 95.055 4.040 ;
        RECT 20.150 3.705 20.880 4.035 ;
        RECT 38.710 3.705 39.440 4.035 ;
        RECT 57.270 3.705 58.000 4.035 ;
        RECT 75.830 3.705 76.560 4.035 ;
        RECT 94.390 3.705 95.120 4.035 ;
        RECT 20.490 3.700 20.815 3.705 ;
        RECT 39.050 3.700 39.375 3.705 ;
        RECT 57.610 3.700 57.935 3.705 ;
        RECT 76.170 3.700 76.495 3.705 ;
        RECT 94.730 3.700 95.055 3.705 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 34.545 8.750 36.580 8.755 ;
        RECT 14.995 8.745 20.160 8.750 ;
        RECT 25.810 8.745 28.620 8.750 ;
        RECT 31.425 8.745 38.720 8.750 ;
        RECT 44.370 8.745 47.180 8.750 ;
        RECT 49.985 8.745 57.280 8.750 ;
        RECT 62.930 8.745 65.740 8.750 ;
        RECT 68.545 8.745 75.840 8.750 ;
        RECT 81.490 8.745 84.300 8.750 ;
        RECT 87.105 8.745 94.400 8.750 ;
        RECT 100.050 8.745 102.860 8.750 ;
        RECT 105.665 8.745 109.455 8.750 ;
        RECT 14.995 6.660 110.595 8.745 ;
        RECT 15.000 4.100 110.595 6.660 ;
        RECT 18.300 4.095 110.595 4.100 ;
        RECT 30.405 3.720 36.355 4.095 ;
        RECT 48.965 3.720 54.915 4.095 ;
        RECT 67.525 3.720 73.475 4.095 ;
        RECT 86.085 3.720 92.035 4.095 ;
        RECT 104.645 3.720 110.595 4.095 ;
        RECT 31.425 3.715 35.215 3.720 ;
        RECT 49.985 3.715 53.775 3.720 ;
        RECT 68.545 3.715 72.335 3.720 ;
        RECT 87.105 3.715 90.895 3.720 ;
        RECT 105.665 3.715 109.455 3.720 ;
      LAYER li1 ;
        RECT 17.030 10.050 17.205 10.600 ;
        RECT 17.030 8.450 17.200 10.050 ;
        RECT 15.215 7.040 15.385 7.770 ;
        RECT 17.030 7.310 17.205 8.450 ;
        RECT 17.030 7.040 17.200 7.310 ;
        RECT 26.030 7.040 26.200 7.770 ;
        RECT 31.645 7.040 31.815 7.770 ;
        RECT 34.390 7.040 34.560 7.770 ;
        RECT 35.385 7.040 35.555 7.765 ;
        RECT 44.590 7.040 44.760 7.770 ;
        RECT 50.205 7.040 50.375 7.770 ;
        RECT 52.950 7.040 53.120 7.770 ;
        RECT 53.945 7.040 54.115 7.765 ;
        RECT 63.150 7.040 63.320 7.770 ;
        RECT 68.765 7.040 68.935 7.770 ;
        RECT 71.510 7.040 71.680 7.770 ;
        RECT 72.505 7.040 72.675 7.765 ;
        RECT 81.710 7.040 81.880 7.770 ;
        RECT 87.325 7.040 87.495 7.770 ;
        RECT 90.070 7.040 90.240 7.770 ;
        RECT 91.065 7.040 91.235 7.765 ;
        RECT 100.270 7.040 100.440 7.770 ;
        RECT 105.885 7.040 106.055 7.770 ;
        RECT 108.630 7.040 108.800 7.770 ;
        RECT 109.625 7.040 109.795 7.765 ;
        RECT 0.000 7.035 110.495 7.040 ;
        RECT 0.000 5.440 110.595 7.035 ;
        RECT 18.540 5.430 36.355 5.440 ;
        RECT 37.100 5.430 54.915 5.440 ;
        RECT 55.660 5.430 73.475 5.440 ;
        RECT 74.220 5.430 92.035 5.440 ;
        RECT 92.780 5.430 110.595 5.440 ;
        RECT 18.540 5.425 30.500 5.430 ;
        RECT 31.475 5.425 35.210 5.430 ;
        RECT 19.350 4.925 19.520 5.425 ;
        RECT 20.310 4.925 20.480 5.425 ;
        RECT 21.310 4.925 21.480 5.425 ;
        RECT 23.270 4.925 23.440 5.425 ;
        RECT 24.230 4.925 24.400 5.425 ;
        RECT 26.190 4.925 26.360 5.425 ;
        RECT 28.630 4.925 28.800 5.425 ;
        RECT 31.645 4.695 31.815 5.425 ;
        RECT 34.390 4.695 34.560 5.425 ;
        RECT 35.380 4.700 35.550 5.430 ;
        RECT 37.100 5.425 49.060 5.430 ;
        RECT 50.035 5.425 53.770 5.430 ;
        RECT 37.910 4.925 38.080 5.425 ;
        RECT 38.870 4.925 39.040 5.425 ;
        RECT 39.870 4.925 40.040 5.425 ;
        RECT 41.830 4.925 42.000 5.425 ;
        RECT 42.790 4.925 42.960 5.425 ;
        RECT 44.750 4.925 44.920 5.425 ;
        RECT 47.190 4.925 47.360 5.425 ;
        RECT 50.205 4.695 50.375 5.425 ;
        RECT 52.950 4.695 53.120 5.425 ;
        RECT 53.940 4.700 54.110 5.430 ;
        RECT 55.660 5.425 67.620 5.430 ;
        RECT 68.595 5.425 72.330 5.430 ;
        RECT 56.470 4.925 56.640 5.425 ;
        RECT 57.430 4.925 57.600 5.425 ;
        RECT 58.430 4.925 58.600 5.425 ;
        RECT 60.390 4.925 60.560 5.425 ;
        RECT 61.350 4.925 61.520 5.425 ;
        RECT 63.310 4.925 63.480 5.425 ;
        RECT 65.750 4.925 65.920 5.425 ;
        RECT 68.765 4.695 68.935 5.425 ;
        RECT 71.510 4.695 71.680 5.425 ;
        RECT 72.500 4.700 72.670 5.430 ;
        RECT 74.220 5.425 86.180 5.430 ;
        RECT 87.155 5.425 90.890 5.430 ;
        RECT 75.030 4.925 75.200 5.425 ;
        RECT 75.990 4.925 76.160 5.425 ;
        RECT 76.990 4.925 77.160 5.425 ;
        RECT 78.950 4.925 79.120 5.425 ;
        RECT 79.910 4.925 80.080 5.425 ;
        RECT 81.870 4.925 82.040 5.425 ;
        RECT 84.310 4.925 84.480 5.425 ;
        RECT 87.325 4.695 87.495 5.425 ;
        RECT 90.070 4.695 90.240 5.425 ;
        RECT 91.060 4.700 91.230 5.430 ;
        RECT 92.780 5.425 104.740 5.430 ;
        RECT 105.715 5.425 109.450 5.430 ;
        RECT 93.590 4.925 93.760 5.425 ;
        RECT 94.550 4.925 94.720 5.425 ;
        RECT 95.550 4.925 95.720 5.425 ;
        RECT 97.510 4.925 97.680 5.425 ;
        RECT 98.470 4.925 98.640 5.425 ;
        RECT 100.430 4.925 100.600 5.425 ;
        RECT 102.870 4.925 103.040 5.425 ;
        RECT 105.885 4.695 106.055 5.425 ;
        RECT 108.630 4.695 108.800 5.425 ;
        RECT 109.620 4.700 109.790 5.430 ;
      LAYER met1 ;
        RECT 16.970 9.150 17.260 9.180 ;
        RECT 16.800 8.980 17.260 9.150 ;
        RECT 16.970 8.950 17.260 8.980 ;
        RECT 0.000 7.035 110.495 7.040 ;
        RECT 0.000 5.440 110.595 7.035 ;
        RECT 18.540 5.430 36.355 5.440 ;
        RECT 37.100 5.430 54.915 5.440 ;
        RECT 55.660 5.430 73.475 5.440 ;
        RECT 74.220 5.430 92.035 5.440 ;
        RECT 92.780 5.430 110.595 5.440 ;
        RECT 18.540 5.395 30.500 5.430 ;
        RECT 31.475 5.425 35.210 5.430 ;
        RECT 37.100 5.395 49.060 5.430 ;
        RECT 50.035 5.425 53.770 5.430 ;
        RECT 55.660 5.395 67.620 5.430 ;
        RECT 68.595 5.425 72.330 5.430 ;
        RECT 74.220 5.395 86.180 5.430 ;
        RECT 87.155 5.425 90.890 5.430 ;
        RECT 92.780 5.395 104.740 5.430 ;
        RECT 105.715 5.425 109.450 5.430 ;
    END
  END vccd1
  OBS
      LAYER pwell ;
        RECT 18.700 2.735 18.870 2.875 ;
        RECT 18.680 2.715 18.870 2.735 ;
        RECT 18.680 2.705 18.850 2.715 ;
        RECT 20.660 2.705 20.830 2.875 ;
        RECT 23.100 2.705 23.270 2.875 ;
        RECT 25.540 2.705 25.710 2.875 ;
        RECT 27.500 2.705 27.670 2.875 ;
        RECT 37.260 2.735 37.430 2.875 ;
        RECT 37.240 2.715 37.430 2.735 ;
        RECT 37.240 2.705 37.410 2.715 ;
        RECT 39.220 2.705 39.390 2.875 ;
        RECT 41.660 2.705 41.830 2.875 ;
        RECT 44.100 2.705 44.270 2.875 ;
        RECT 46.060 2.705 46.230 2.875 ;
        RECT 55.820 2.735 55.990 2.875 ;
        RECT 55.800 2.715 55.990 2.735 ;
        RECT 55.800 2.705 55.970 2.715 ;
        RECT 57.780 2.705 57.950 2.875 ;
        RECT 60.220 2.705 60.390 2.875 ;
        RECT 62.660 2.705 62.830 2.875 ;
        RECT 64.620 2.705 64.790 2.875 ;
        RECT 74.380 2.735 74.550 2.875 ;
        RECT 74.360 2.715 74.550 2.735 ;
        RECT 74.360 2.705 74.530 2.715 ;
        RECT 76.340 2.705 76.510 2.875 ;
        RECT 78.780 2.705 78.950 2.875 ;
        RECT 81.220 2.705 81.390 2.875 ;
        RECT 83.180 2.705 83.350 2.875 ;
        RECT 92.940 2.735 93.110 2.875 ;
        RECT 92.920 2.715 93.110 2.735 ;
        RECT 92.920 2.705 93.090 2.715 ;
        RECT 94.900 2.705 95.070 2.875 ;
        RECT 97.340 2.705 97.510 2.875 ;
        RECT 99.780 2.705 99.950 2.875 ;
        RECT 101.740 2.705 101.910 2.875 ;
      LAYER li1 ;
        RECT 15.645 10.110 15.820 10.600 ;
        RECT 16.170 10.320 16.340 10.600 ;
        RECT 16.170 10.150 16.400 10.320 ;
        RECT 15.645 9.940 15.815 10.110 ;
        RECT 15.645 9.610 16.055 9.940 ;
        RECT 15.645 9.100 15.815 9.610 ;
        RECT 15.645 8.770 16.055 9.100 ;
        RECT 15.645 8.570 15.815 8.770 ;
        RECT 15.645 7.310 15.820 8.570 ;
        RECT 16.230 8.540 16.400 10.150 ;
        RECT 16.600 10.090 16.775 10.600 ;
        RECT 26.460 10.110 26.635 10.600 ;
        RECT 26.460 9.940 26.630 10.110 ;
        RECT 27.415 10.090 27.590 10.600 ;
        RECT 27.845 10.050 28.020 10.600 ;
        RECT 32.075 10.110 32.250 10.600 ;
        RECT 32.600 10.320 32.770 10.600 ;
        RECT 32.600 10.150 32.830 10.320 ;
        RECT 26.460 9.610 26.870 9.940 ;
        RECT 16.170 8.370 16.400 8.540 ;
        RECT 16.600 8.570 16.770 9.520 ;
        RECT 26.460 9.100 26.630 9.610 ;
        RECT 26.460 8.770 26.870 9.100 ;
        RECT 26.460 8.570 26.630 8.770 ;
        RECT 27.415 8.570 27.585 9.520 ;
        RECT 16.170 7.310 16.340 8.370 ;
        RECT 16.600 7.310 16.775 8.570 ;
        RECT 26.460 7.310 26.635 8.570 ;
        RECT 27.415 7.310 27.590 8.570 ;
        RECT 27.845 8.450 28.015 10.050 ;
        RECT 32.075 9.940 32.245 10.110 ;
        RECT 32.075 9.610 32.485 9.940 ;
        RECT 32.075 9.100 32.245 9.610 ;
        RECT 32.075 8.770 32.485 9.100 ;
        RECT 32.075 8.570 32.245 8.770 ;
        RECT 27.845 7.310 28.020 8.450 ;
        RECT 32.075 7.310 32.250 8.570 ;
        RECT 32.660 8.540 32.830 10.150 ;
        RECT 33.030 10.090 33.205 10.600 ;
        RECT 33.460 10.050 33.635 10.600 ;
        RECT 34.825 10.090 34.995 10.600 ;
        RECT 35.820 10.085 35.990 10.595 ;
        RECT 45.020 10.110 45.195 10.600 ;
        RECT 32.600 8.370 32.830 8.540 ;
        RECT 33.030 8.570 33.200 9.520 ;
        RECT 32.600 7.310 32.770 8.370 ;
        RECT 33.030 7.310 33.205 8.570 ;
        RECT 33.460 8.450 33.630 10.050 ;
        RECT 45.020 9.940 45.190 10.110 ;
        RECT 45.975 10.090 46.150 10.600 ;
        RECT 46.405 10.050 46.580 10.600 ;
        RECT 50.635 10.110 50.810 10.600 ;
        RECT 51.160 10.320 51.330 10.600 ;
        RECT 51.160 10.150 51.390 10.320 ;
        RECT 45.020 9.610 45.430 9.940 ;
        RECT 34.390 9.430 34.620 9.600 ;
        RECT 34.390 9.370 34.920 9.430 ;
        RECT 34.450 9.260 34.920 9.370 ;
        RECT 34.450 8.570 34.620 9.260 ;
        RECT 35.445 9.255 35.915 9.425 ;
        RECT 34.820 8.810 34.990 8.890 ;
        RECT 35.445 8.810 35.615 9.255 ;
        RECT 45.020 9.100 45.190 9.610 ;
        RECT 34.820 8.610 35.615 8.810 ;
        RECT 33.460 7.310 33.635 8.450 ;
        RECT 34.820 7.310 34.995 8.610 ;
        RECT 35.445 8.565 35.615 8.610 ;
        RECT 35.815 8.450 35.985 8.885 ;
        RECT 45.020 8.770 45.430 9.100 ;
        RECT 45.020 8.570 45.190 8.770 ;
        RECT 45.975 8.570 46.145 9.520 ;
        RECT 35.815 7.305 35.990 8.450 ;
        RECT 45.020 7.310 45.195 8.570 ;
        RECT 45.975 7.310 46.150 8.570 ;
        RECT 46.405 8.450 46.575 10.050 ;
        RECT 50.635 9.940 50.805 10.110 ;
        RECT 50.635 9.610 51.045 9.940 ;
        RECT 50.635 9.100 50.805 9.610 ;
        RECT 50.635 8.770 51.045 9.100 ;
        RECT 50.635 8.570 50.805 8.770 ;
        RECT 46.405 7.310 46.580 8.450 ;
        RECT 50.635 7.310 50.810 8.570 ;
        RECT 51.220 8.540 51.390 10.150 ;
        RECT 51.590 10.090 51.765 10.600 ;
        RECT 52.020 10.050 52.195 10.600 ;
        RECT 53.385 10.090 53.555 10.600 ;
        RECT 54.380 10.085 54.550 10.595 ;
        RECT 63.580 10.110 63.755 10.600 ;
        RECT 51.160 8.370 51.390 8.540 ;
        RECT 51.590 8.570 51.760 9.520 ;
        RECT 51.160 7.310 51.330 8.370 ;
        RECT 51.590 7.310 51.765 8.570 ;
        RECT 52.020 8.450 52.190 10.050 ;
        RECT 63.580 9.940 63.750 10.110 ;
        RECT 64.535 10.090 64.710 10.600 ;
        RECT 64.965 10.050 65.140 10.600 ;
        RECT 69.195 10.110 69.370 10.600 ;
        RECT 69.720 10.320 69.890 10.600 ;
        RECT 69.720 10.150 69.950 10.320 ;
        RECT 63.580 9.610 63.990 9.940 ;
        RECT 52.950 9.430 53.180 9.600 ;
        RECT 52.950 9.370 53.480 9.430 ;
        RECT 53.010 9.260 53.480 9.370 ;
        RECT 53.010 8.570 53.180 9.260 ;
        RECT 54.005 9.255 54.475 9.425 ;
        RECT 53.380 8.810 53.550 8.890 ;
        RECT 54.005 8.810 54.175 9.255 ;
        RECT 63.580 9.100 63.750 9.610 ;
        RECT 53.380 8.610 54.175 8.810 ;
        RECT 52.020 7.310 52.195 8.450 ;
        RECT 53.380 7.310 53.555 8.610 ;
        RECT 54.005 8.565 54.175 8.610 ;
        RECT 54.375 8.450 54.545 8.885 ;
        RECT 63.580 8.770 63.990 9.100 ;
        RECT 63.580 8.570 63.750 8.770 ;
        RECT 64.535 8.570 64.705 9.520 ;
        RECT 54.375 7.305 54.550 8.450 ;
        RECT 63.580 7.310 63.755 8.570 ;
        RECT 64.535 7.310 64.710 8.570 ;
        RECT 64.965 8.450 65.135 10.050 ;
        RECT 69.195 9.940 69.365 10.110 ;
        RECT 69.195 9.610 69.605 9.940 ;
        RECT 69.195 9.100 69.365 9.610 ;
        RECT 69.195 8.770 69.605 9.100 ;
        RECT 69.195 8.570 69.365 8.770 ;
        RECT 64.965 7.310 65.140 8.450 ;
        RECT 69.195 7.310 69.370 8.570 ;
        RECT 69.780 8.540 69.950 10.150 ;
        RECT 70.150 10.090 70.325 10.600 ;
        RECT 70.580 10.050 70.755 10.600 ;
        RECT 71.945 10.090 72.115 10.600 ;
        RECT 72.940 10.085 73.110 10.595 ;
        RECT 82.140 10.110 82.315 10.600 ;
        RECT 69.720 8.370 69.950 8.540 ;
        RECT 70.150 8.570 70.320 9.520 ;
        RECT 69.720 7.310 69.890 8.370 ;
        RECT 70.150 7.310 70.325 8.570 ;
        RECT 70.580 8.450 70.750 10.050 ;
        RECT 82.140 9.940 82.310 10.110 ;
        RECT 83.095 10.090 83.270 10.600 ;
        RECT 83.525 10.050 83.700 10.600 ;
        RECT 87.755 10.110 87.930 10.600 ;
        RECT 88.280 10.320 88.450 10.600 ;
        RECT 88.280 10.150 88.510 10.320 ;
        RECT 82.140 9.610 82.550 9.940 ;
        RECT 71.510 9.430 71.740 9.600 ;
        RECT 71.510 9.370 72.040 9.430 ;
        RECT 71.570 9.260 72.040 9.370 ;
        RECT 71.570 8.570 71.740 9.260 ;
        RECT 72.565 9.255 73.035 9.425 ;
        RECT 71.940 8.810 72.110 8.890 ;
        RECT 72.565 8.810 72.735 9.255 ;
        RECT 82.140 9.100 82.310 9.610 ;
        RECT 71.940 8.610 72.735 8.810 ;
        RECT 70.580 7.310 70.755 8.450 ;
        RECT 71.940 7.310 72.115 8.610 ;
        RECT 72.565 8.565 72.735 8.610 ;
        RECT 72.935 8.450 73.105 8.885 ;
        RECT 82.140 8.770 82.550 9.100 ;
        RECT 82.140 8.570 82.310 8.770 ;
        RECT 83.095 8.570 83.265 9.520 ;
        RECT 72.935 7.305 73.110 8.450 ;
        RECT 82.140 7.310 82.315 8.570 ;
        RECT 83.095 7.310 83.270 8.570 ;
        RECT 83.525 8.450 83.695 10.050 ;
        RECT 87.755 9.940 87.925 10.110 ;
        RECT 87.755 9.610 88.165 9.940 ;
        RECT 87.755 9.100 87.925 9.610 ;
        RECT 87.755 8.770 88.165 9.100 ;
        RECT 87.755 8.570 87.925 8.770 ;
        RECT 83.525 7.310 83.700 8.450 ;
        RECT 87.755 7.310 87.930 8.570 ;
        RECT 88.340 8.540 88.510 10.150 ;
        RECT 88.710 10.090 88.885 10.600 ;
        RECT 89.140 10.050 89.315 10.600 ;
        RECT 90.505 10.090 90.675 10.600 ;
        RECT 91.500 10.085 91.670 10.595 ;
        RECT 100.700 10.110 100.875 10.600 ;
        RECT 88.280 8.370 88.510 8.540 ;
        RECT 88.710 8.570 88.880 9.520 ;
        RECT 88.280 7.310 88.450 8.370 ;
        RECT 88.710 7.310 88.885 8.570 ;
        RECT 89.140 8.450 89.310 10.050 ;
        RECT 100.700 9.940 100.870 10.110 ;
        RECT 101.655 10.090 101.830 10.600 ;
        RECT 102.085 10.050 102.260 10.600 ;
        RECT 106.315 10.110 106.490 10.600 ;
        RECT 106.840 10.320 107.010 10.600 ;
        RECT 106.840 10.150 107.070 10.320 ;
        RECT 100.700 9.610 101.110 9.940 ;
        RECT 90.070 9.430 90.300 9.600 ;
        RECT 90.070 9.370 90.600 9.430 ;
        RECT 90.130 9.260 90.600 9.370 ;
        RECT 90.130 8.570 90.300 9.260 ;
        RECT 91.125 9.255 91.595 9.425 ;
        RECT 90.500 8.810 90.670 8.890 ;
        RECT 91.125 8.810 91.295 9.255 ;
        RECT 100.700 9.100 100.870 9.610 ;
        RECT 90.500 8.610 91.295 8.810 ;
        RECT 89.140 7.310 89.315 8.450 ;
        RECT 90.500 7.310 90.675 8.610 ;
        RECT 91.125 8.565 91.295 8.610 ;
        RECT 91.495 8.450 91.665 8.885 ;
        RECT 100.700 8.770 101.110 9.100 ;
        RECT 100.700 8.570 100.870 8.770 ;
        RECT 101.655 8.570 101.825 9.520 ;
        RECT 91.495 7.305 91.670 8.450 ;
        RECT 100.700 7.310 100.875 8.570 ;
        RECT 101.655 7.310 101.830 8.570 ;
        RECT 102.085 8.450 102.255 10.050 ;
        RECT 106.315 9.940 106.485 10.110 ;
        RECT 106.315 9.610 106.725 9.940 ;
        RECT 106.315 9.100 106.485 9.610 ;
        RECT 106.315 8.770 106.725 9.100 ;
        RECT 106.315 8.570 106.485 8.770 ;
        RECT 102.085 7.310 102.260 8.450 ;
        RECT 106.315 7.310 106.490 8.570 ;
        RECT 106.900 8.540 107.070 10.150 ;
        RECT 107.270 10.090 107.445 10.600 ;
        RECT 107.700 10.050 107.875 10.600 ;
        RECT 109.065 10.090 109.235 10.600 ;
        RECT 110.060 10.085 110.230 10.595 ;
        RECT 106.840 8.370 107.070 8.540 ;
        RECT 107.270 8.570 107.440 9.520 ;
        RECT 106.840 7.310 107.010 8.370 ;
        RECT 107.270 7.310 107.445 8.570 ;
        RECT 107.700 8.450 107.870 10.050 ;
        RECT 108.630 9.430 108.860 9.600 ;
        RECT 108.630 9.370 109.160 9.430 ;
        RECT 108.690 9.260 109.160 9.370 ;
        RECT 108.690 8.570 108.860 9.260 ;
        RECT 109.685 9.255 110.155 9.425 ;
        RECT 109.060 8.810 109.230 8.890 ;
        RECT 109.685 8.810 109.855 9.255 ;
        RECT 109.060 8.610 109.855 8.810 ;
        RECT 107.700 7.310 107.875 8.450 ;
        RECT 109.060 7.310 109.235 8.610 ;
        RECT 109.685 8.565 109.855 8.610 ;
        RECT 110.055 8.450 110.225 8.885 ;
        RECT 110.055 7.305 110.230 8.450 ;
        RECT 18.870 4.575 19.040 4.935 ;
        RECT 19.830 4.605 20.000 4.765 ;
        RECT 21.790 4.685 21.960 4.795 ;
        RECT 19.210 4.435 20.000 4.605 ;
        RECT 20.750 4.515 22.040 4.685 ;
        RECT 19.210 4.375 19.380 4.435 ;
        RECT 19.110 4.205 19.380 4.375 ;
        RECT 19.830 4.345 20.000 4.435 ;
        RECT 22.270 4.345 22.440 4.765 ;
        RECT 22.750 4.435 22.920 4.795 ;
        RECT 23.670 4.515 24.160 4.685 ;
        RECT 19.110 4.135 19.280 4.205 ;
        RECT 18.870 3.865 19.280 4.135 ;
        RECT 19.110 3.785 19.280 3.865 ;
        RECT 19.590 3.785 19.760 4.115 ;
        RECT 20.740 3.865 21.320 4.035 ;
        RECT 20.740 3.785 20.910 3.865 ;
        RECT 21.550 3.785 21.720 4.235 ;
        RECT 23.270 4.035 23.440 4.515 ;
        RECT 23.990 4.345 25.000 4.515 ;
        RECT 25.190 4.435 25.360 5.075 ;
        RECT 25.710 4.775 25.880 5.105 ;
        RECT 26.670 4.905 27.320 5.075 ;
        RECT 27.030 4.515 27.320 4.905 ;
        RECT 28.030 4.905 28.320 5.075 ;
        RECT 24.830 4.115 25.000 4.345 ;
        RECT 25.710 4.375 25.880 4.515 ;
        RECT 27.150 4.435 27.320 4.515 ;
        RECT 25.710 4.205 26.600 4.375 ;
        RECT 27.670 4.345 27.840 4.765 ;
        RECT 28.030 4.515 28.200 4.905 ;
        RECT 28.870 4.515 29.840 4.685 ;
        RECT 28.030 4.345 28.320 4.515 ;
        RECT 28.870 4.345 29.040 4.515 ;
        RECT 22.430 3.865 22.920 4.035 ;
        RECT 23.270 3.865 23.760 4.035 ;
        RECT 22.750 3.785 22.920 3.865 ;
        RECT 23.990 3.785 24.160 4.115 ;
        RECT 24.470 3.785 24.640 4.115 ;
        RECT 24.830 3.865 25.120 4.115 ;
        RECT 24.950 3.785 25.120 3.865 ;
        RECT 25.710 3.865 26.200 4.035 ;
        RECT 25.710 3.785 25.880 3.865 ;
        RECT 26.430 3.785 26.600 4.205 ;
        RECT 27.150 4.135 27.320 4.235 ;
        RECT 26.910 4.035 27.320 4.135 ;
        RECT 28.030 4.035 28.200 4.345 ;
        RECT 26.830 3.965 27.320 4.035 ;
        RECT 26.830 3.865 27.160 3.965 ;
        RECT 27.830 3.865 28.200 4.035 ;
        RECT 28.390 4.035 28.560 4.115 ;
        RECT 28.390 3.865 29.120 4.035 ;
        RECT 28.390 3.785 28.560 3.865 ;
        RECT 29.350 3.785 29.520 4.235 ;
        RECT 32.075 3.895 32.250 5.155 ;
        RECT 32.600 4.095 32.770 5.155 ;
        RECT 32.600 3.925 32.830 4.095 ;
        RECT 32.075 3.695 32.245 3.895 ;
        RECT 18.870 3.045 19.040 3.395 ;
        RECT 19.830 3.295 20.000 3.395 ;
        RECT 22.270 3.295 22.440 3.395 ;
        RECT 23.750 3.295 23.920 3.395 ;
        RECT 19.830 3.125 20.560 3.295 ;
        RECT 21.710 3.125 22.440 3.295 ;
        RECT 23.190 3.125 23.920 3.295 ;
        RECT 24.710 3.045 24.880 3.395 ;
        RECT 25.710 3.045 25.880 3.395 ;
        RECT 26.670 3.045 26.840 3.395 ;
        RECT 28.150 3.045 28.320 3.395 ;
        RECT 29.110 3.045 29.280 3.395 ;
        RECT 32.075 3.365 32.485 3.695 ;
        RECT 32.075 2.855 32.245 3.365 ;
        RECT 32.075 2.525 32.485 2.855 ;
        RECT 32.075 2.355 32.245 2.525 ;
        RECT 32.075 1.865 32.250 2.355 ;
        RECT 32.660 2.315 32.830 3.925 ;
        RECT 33.030 3.895 33.205 5.155 ;
        RECT 33.460 4.015 33.635 5.155 ;
        RECT 33.030 2.945 33.200 3.895 ;
        RECT 33.460 2.415 33.630 4.015 ;
        RECT 34.820 4.010 34.995 5.155 ;
        RECT 37.430 4.575 37.600 4.935 ;
        RECT 38.390 4.605 38.560 4.765 ;
        RECT 40.350 4.685 40.520 4.795 ;
        RECT 37.770 4.435 38.560 4.605 ;
        RECT 39.310 4.515 40.600 4.685 ;
        RECT 37.770 4.375 37.940 4.435 ;
        RECT 37.670 4.205 37.940 4.375 ;
        RECT 38.390 4.345 38.560 4.435 ;
        RECT 40.830 4.345 41.000 4.765 ;
        RECT 41.310 4.435 41.480 4.795 ;
        RECT 42.230 4.515 42.720 4.685 ;
        RECT 37.670 4.135 37.840 4.205 ;
        RECT 34.450 3.205 34.620 3.895 ;
        RECT 34.820 3.805 34.990 4.010 ;
        RECT 35.440 3.805 35.610 3.900 ;
        RECT 37.430 3.865 37.840 4.135 ;
        RECT 34.820 3.625 35.610 3.805 ;
        RECT 37.670 3.785 37.840 3.865 ;
        RECT 38.150 3.785 38.320 4.115 ;
        RECT 39.300 3.865 39.880 4.035 ;
        RECT 39.300 3.785 39.470 3.865 ;
        RECT 40.110 3.785 40.280 4.235 ;
        RECT 41.830 4.035 42.000 4.515 ;
        RECT 42.550 4.345 43.560 4.515 ;
        RECT 43.750 4.435 43.920 5.075 ;
        RECT 44.270 4.775 44.440 5.105 ;
        RECT 45.230 4.905 45.880 5.075 ;
        RECT 45.590 4.515 45.880 4.905 ;
        RECT 46.590 4.905 46.880 5.075 ;
        RECT 43.390 4.115 43.560 4.345 ;
        RECT 44.270 4.375 44.440 4.515 ;
        RECT 45.710 4.435 45.880 4.515 ;
        RECT 44.270 4.205 45.160 4.375 ;
        RECT 46.230 4.345 46.400 4.765 ;
        RECT 46.590 4.515 46.760 4.905 ;
        RECT 47.430 4.515 48.400 4.685 ;
        RECT 46.590 4.345 46.880 4.515 ;
        RECT 47.430 4.345 47.600 4.515 ;
        RECT 40.990 3.865 41.480 4.035 ;
        RECT 41.830 3.865 42.320 4.035 ;
        RECT 41.310 3.785 41.480 3.865 ;
        RECT 42.550 3.785 42.720 4.115 ;
        RECT 43.030 3.785 43.200 4.115 ;
        RECT 43.390 3.865 43.680 4.115 ;
        RECT 43.510 3.785 43.680 3.865 ;
        RECT 44.270 3.865 44.760 4.035 ;
        RECT 44.270 3.785 44.440 3.865 ;
        RECT 44.990 3.785 45.160 4.205 ;
        RECT 45.710 4.135 45.880 4.235 ;
        RECT 45.470 4.035 45.880 4.135 ;
        RECT 46.590 4.035 46.760 4.345 ;
        RECT 45.390 3.965 45.880 4.035 ;
        RECT 45.390 3.865 45.720 3.965 ;
        RECT 46.390 3.865 46.760 4.035 ;
        RECT 46.950 4.035 47.120 4.115 ;
        RECT 46.950 3.865 47.680 4.035 ;
        RECT 46.950 3.785 47.120 3.865 ;
        RECT 47.910 3.785 48.080 4.235 ;
        RECT 50.635 3.895 50.810 5.155 ;
        RECT 51.160 4.095 51.330 5.155 ;
        RECT 51.160 3.925 51.390 4.095 ;
        RECT 34.820 3.575 34.990 3.625 ;
        RECT 35.440 3.210 35.610 3.625 ;
        RECT 50.635 3.695 50.805 3.895 ;
        RECT 34.450 3.175 34.920 3.205 ;
        RECT 34.390 3.035 34.920 3.175 ;
        RECT 35.440 3.040 35.910 3.210 ;
        RECT 37.430 3.045 37.600 3.395 ;
        RECT 38.390 3.295 38.560 3.395 ;
        RECT 40.830 3.295 41.000 3.395 ;
        RECT 42.310 3.295 42.480 3.395 ;
        RECT 38.390 3.125 39.120 3.295 ;
        RECT 40.270 3.125 41.000 3.295 ;
        RECT 41.750 3.125 42.480 3.295 ;
        RECT 43.270 3.045 43.440 3.395 ;
        RECT 44.270 3.045 44.440 3.395 ;
        RECT 45.230 3.045 45.400 3.395 ;
        RECT 46.710 3.045 46.880 3.395 ;
        RECT 47.670 3.045 47.840 3.395 ;
        RECT 50.635 3.365 51.045 3.695 ;
        RECT 34.390 2.945 34.620 3.035 ;
        RECT 50.635 2.855 50.805 3.365 ;
        RECT 50.635 2.525 51.045 2.855 ;
        RECT 32.600 2.145 32.830 2.315 ;
        RECT 32.600 1.865 32.770 2.145 ;
        RECT 33.030 1.865 33.205 2.375 ;
        RECT 33.460 1.865 33.635 2.415 ;
        RECT 34.825 1.865 34.995 2.375 ;
        RECT 50.635 2.355 50.805 2.525 ;
        RECT 50.635 1.865 50.810 2.355 ;
        RECT 51.220 2.315 51.390 3.925 ;
        RECT 51.590 3.895 51.765 5.155 ;
        RECT 52.020 4.015 52.195 5.155 ;
        RECT 51.590 2.945 51.760 3.895 ;
        RECT 52.020 2.415 52.190 4.015 ;
        RECT 53.380 4.010 53.555 5.155 ;
        RECT 55.990 4.575 56.160 4.935 ;
        RECT 56.950 4.605 57.120 4.765 ;
        RECT 58.910 4.685 59.080 4.795 ;
        RECT 56.330 4.435 57.120 4.605 ;
        RECT 57.870 4.515 59.160 4.685 ;
        RECT 56.330 4.375 56.500 4.435 ;
        RECT 56.230 4.205 56.500 4.375 ;
        RECT 56.950 4.345 57.120 4.435 ;
        RECT 59.390 4.345 59.560 4.765 ;
        RECT 59.870 4.435 60.040 4.795 ;
        RECT 60.790 4.515 61.280 4.685 ;
        RECT 56.230 4.135 56.400 4.205 ;
        RECT 53.010 3.205 53.180 3.895 ;
        RECT 53.380 3.805 53.550 4.010 ;
        RECT 54.000 3.805 54.170 3.900 ;
        RECT 55.990 3.865 56.400 4.135 ;
        RECT 53.380 3.625 54.170 3.805 ;
        RECT 56.230 3.785 56.400 3.865 ;
        RECT 56.710 3.785 56.880 4.115 ;
        RECT 57.860 3.865 58.440 4.035 ;
        RECT 57.860 3.785 58.030 3.865 ;
        RECT 58.670 3.785 58.840 4.235 ;
        RECT 60.390 4.035 60.560 4.515 ;
        RECT 61.110 4.345 62.120 4.515 ;
        RECT 62.310 4.435 62.480 5.075 ;
        RECT 62.830 4.775 63.000 5.105 ;
        RECT 63.790 4.905 64.440 5.075 ;
        RECT 64.150 4.515 64.440 4.905 ;
        RECT 65.150 4.905 65.440 5.075 ;
        RECT 61.950 4.115 62.120 4.345 ;
        RECT 62.830 4.375 63.000 4.515 ;
        RECT 64.270 4.435 64.440 4.515 ;
        RECT 62.830 4.205 63.720 4.375 ;
        RECT 64.790 4.345 64.960 4.765 ;
        RECT 65.150 4.515 65.320 4.905 ;
        RECT 65.990 4.515 66.960 4.685 ;
        RECT 65.150 4.345 65.440 4.515 ;
        RECT 65.990 4.345 66.160 4.515 ;
        RECT 59.550 3.865 60.040 4.035 ;
        RECT 60.390 3.865 60.880 4.035 ;
        RECT 59.870 3.785 60.040 3.865 ;
        RECT 61.110 3.785 61.280 4.115 ;
        RECT 61.590 3.785 61.760 4.115 ;
        RECT 61.950 3.865 62.240 4.115 ;
        RECT 62.070 3.785 62.240 3.865 ;
        RECT 62.830 3.865 63.320 4.035 ;
        RECT 62.830 3.785 63.000 3.865 ;
        RECT 63.550 3.785 63.720 4.205 ;
        RECT 64.270 4.135 64.440 4.235 ;
        RECT 64.030 4.035 64.440 4.135 ;
        RECT 65.150 4.035 65.320 4.345 ;
        RECT 63.950 3.965 64.440 4.035 ;
        RECT 63.950 3.865 64.280 3.965 ;
        RECT 64.950 3.865 65.320 4.035 ;
        RECT 65.510 4.035 65.680 4.115 ;
        RECT 65.510 3.865 66.240 4.035 ;
        RECT 65.510 3.785 65.680 3.865 ;
        RECT 66.470 3.785 66.640 4.235 ;
        RECT 69.195 3.895 69.370 5.155 ;
        RECT 69.720 4.095 69.890 5.155 ;
        RECT 69.720 3.925 69.950 4.095 ;
        RECT 53.380 3.575 53.550 3.625 ;
        RECT 54.000 3.210 54.170 3.625 ;
        RECT 69.195 3.695 69.365 3.895 ;
        RECT 53.010 3.175 53.480 3.205 ;
        RECT 52.950 3.035 53.480 3.175 ;
        RECT 54.000 3.040 54.470 3.210 ;
        RECT 55.990 3.045 56.160 3.395 ;
        RECT 56.950 3.295 57.120 3.395 ;
        RECT 59.390 3.295 59.560 3.395 ;
        RECT 60.870 3.295 61.040 3.395 ;
        RECT 56.950 3.125 57.680 3.295 ;
        RECT 58.830 3.125 59.560 3.295 ;
        RECT 60.310 3.125 61.040 3.295 ;
        RECT 61.830 3.045 62.000 3.395 ;
        RECT 62.830 3.045 63.000 3.395 ;
        RECT 63.790 3.045 63.960 3.395 ;
        RECT 65.270 3.045 65.440 3.395 ;
        RECT 66.230 3.045 66.400 3.395 ;
        RECT 69.195 3.365 69.605 3.695 ;
        RECT 52.950 2.945 53.180 3.035 ;
        RECT 69.195 2.855 69.365 3.365 ;
        RECT 69.195 2.525 69.605 2.855 ;
        RECT 51.160 2.145 51.390 2.315 ;
        RECT 51.160 1.865 51.330 2.145 ;
        RECT 51.590 1.865 51.765 2.375 ;
        RECT 52.020 1.865 52.195 2.415 ;
        RECT 53.385 1.865 53.555 2.375 ;
        RECT 69.195 2.355 69.365 2.525 ;
        RECT 69.195 1.865 69.370 2.355 ;
        RECT 69.780 2.315 69.950 3.925 ;
        RECT 70.150 3.895 70.325 5.155 ;
        RECT 70.580 4.015 70.755 5.155 ;
        RECT 70.150 2.945 70.320 3.895 ;
        RECT 70.580 2.415 70.750 4.015 ;
        RECT 71.940 4.010 72.115 5.155 ;
        RECT 74.550 4.575 74.720 4.935 ;
        RECT 75.510 4.605 75.680 4.765 ;
        RECT 77.470 4.685 77.640 4.795 ;
        RECT 74.890 4.435 75.680 4.605 ;
        RECT 76.430 4.515 77.720 4.685 ;
        RECT 74.890 4.375 75.060 4.435 ;
        RECT 74.790 4.205 75.060 4.375 ;
        RECT 75.510 4.345 75.680 4.435 ;
        RECT 77.950 4.345 78.120 4.765 ;
        RECT 78.430 4.435 78.600 4.795 ;
        RECT 79.350 4.515 79.840 4.685 ;
        RECT 74.790 4.135 74.960 4.205 ;
        RECT 71.570 3.205 71.740 3.895 ;
        RECT 71.940 3.805 72.110 4.010 ;
        RECT 72.560 3.805 72.730 3.900 ;
        RECT 74.550 3.865 74.960 4.135 ;
        RECT 71.940 3.625 72.730 3.805 ;
        RECT 74.790 3.785 74.960 3.865 ;
        RECT 75.270 3.785 75.440 4.115 ;
        RECT 76.420 3.865 77.000 4.035 ;
        RECT 76.420 3.785 76.590 3.865 ;
        RECT 77.230 3.785 77.400 4.235 ;
        RECT 78.950 4.035 79.120 4.515 ;
        RECT 79.670 4.345 80.680 4.515 ;
        RECT 80.870 4.435 81.040 5.075 ;
        RECT 81.390 4.775 81.560 5.105 ;
        RECT 82.350 4.905 83.000 5.075 ;
        RECT 82.710 4.515 83.000 4.905 ;
        RECT 83.710 4.905 84.000 5.075 ;
        RECT 80.510 4.115 80.680 4.345 ;
        RECT 81.390 4.375 81.560 4.515 ;
        RECT 82.830 4.435 83.000 4.515 ;
        RECT 81.390 4.205 82.280 4.375 ;
        RECT 83.350 4.345 83.520 4.765 ;
        RECT 83.710 4.515 83.880 4.905 ;
        RECT 84.550 4.515 85.520 4.685 ;
        RECT 83.710 4.345 84.000 4.515 ;
        RECT 84.550 4.345 84.720 4.515 ;
        RECT 78.110 3.865 78.600 4.035 ;
        RECT 78.950 3.865 79.440 4.035 ;
        RECT 78.430 3.785 78.600 3.865 ;
        RECT 79.670 3.785 79.840 4.115 ;
        RECT 80.150 3.785 80.320 4.115 ;
        RECT 80.510 3.865 80.800 4.115 ;
        RECT 80.630 3.785 80.800 3.865 ;
        RECT 81.390 3.865 81.880 4.035 ;
        RECT 81.390 3.785 81.560 3.865 ;
        RECT 82.110 3.785 82.280 4.205 ;
        RECT 82.830 4.135 83.000 4.235 ;
        RECT 82.590 4.035 83.000 4.135 ;
        RECT 83.710 4.035 83.880 4.345 ;
        RECT 82.510 3.965 83.000 4.035 ;
        RECT 82.510 3.865 82.840 3.965 ;
        RECT 83.510 3.865 83.880 4.035 ;
        RECT 84.070 4.035 84.240 4.115 ;
        RECT 84.070 3.865 84.800 4.035 ;
        RECT 84.070 3.785 84.240 3.865 ;
        RECT 85.030 3.785 85.200 4.235 ;
        RECT 87.755 3.895 87.930 5.155 ;
        RECT 88.280 4.095 88.450 5.155 ;
        RECT 88.280 3.925 88.510 4.095 ;
        RECT 71.940 3.575 72.110 3.625 ;
        RECT 72.560 3.210 72.730 3.625 ;
        RECT 87.755 3.695 87.925 3.895 ;
        RECT 71.570 3.175 72.040 3.205 ;
        RECT 71.510 3.035 72.040 3.175 ;
        RECT 72.560 3.040 73.030 3.210 ;
        RECT 74.550 3.045 74.720 3.395 ;
        RECT 75.510 3.295 75.680 3.395 ;
        RECT 77.950 3.295 78.120 3.395 ;
        RECT 79.430 3.295 79.600 3.395 ;
        RECT 75.510 3.125 76.240 3.295 ;
        RECT 77.390 3.125 78.120 3.295 ;
        RECT 78.870 3.125 79.600 3.295 ;
        RECT 80.390 3.045 80.560 3.395 ;
        RECT 81.390 3.045 81.560 3.395 ;
        RECT 82.350 3.045 82.520 3.395 ;
        RECT 83.830 3.045 84.000 3.395 ;
        RECT 84.790 3.045 84.960 3.395 ;
        RECT 87.755 3.365 88.165 3.695 ;
        RECT 71.510 2.945 71.740 3.035 ;
        RECT 87.755 2.855 87.925 3.365 ;
        RECT 87.755 2.525 88.165 2.855 ;
        RECT 69.720 2.145 69.950 2.315 ;
        RECT 69.720 1.865 69.890 2.145 ;
        RECT 70.150 1.865 70.325 2.375 ;
        RECT 70.580 1.865 70.755 2.415 ;
        RECT 71.945 1.865 72.115 2.375 ;
        RECT 87.755 2.355 87.925 2.525 ;
        RECT 87.755 1.865 87.930 2.355 ;
        RECT 88.340 2.315 88.510 3.925 ;
        RECT 88.710 3.895 88.885 5.155 ;
        RECT 89.140 4.015 89.315 5.155 ;
        RECT 88.710 2.945 88.880 3.895 ;
        RECT 89.140 2.415 89.310 4.015 ;
        RECT 90.500 4.010 90.675 5.155 ;
        RECT 93.110 4.575 93.280 4.935 ;
        RECT 94.070 4.605 94.240 4.765 ;
        RECT 96.030 4.685 96.200 4.795 ;
        RECT 93.450 4.435 94.240 4.605 ;
        RECT 94.990 4.515 96.280 4.685 ;
        RECT 93.450 4.375 93.620 4.435 ;
        RECT 93.350 4.205 93.620 4.375 ;
        RECT 94.070 4.345 94.240 4.435 ;
        RECT 96.510 4.345 96.680 4.765 ;
        RECT 96.990 4.435 97.160 4.795 ;
        RECT 97.910 4.515 98.400 4.685 ;
        RECT 93.350 4.135 93.520 4.205 ;
        RECT 90.130 3.205 90.300 3.895 ;
        RECT 90.500 3.805 90.670 4.010 ;
        RECT 91.120 3.805 91.290 3.900 ;
        RECT 93.110 3.865 93.520 4.135 ;
        RECT 90.500 3.625 91.290 3.805 ;
        RECT 93.350 3.785 93.520 3.865 ;
        RECT 93.830 3.785 94.000 4.115 ;
        RECT 94.980 3.865 95.560 4.035 ;
        RECT 94.980 3.785 95.150 3.865 ;
        RECT 95.790 3.785 95.960 4.235 ;
        RECT 97.510 4.035 97.680 4.515 ;
        RECT 98.230 4.345 99.240 4.515 ;
        RECT 99.430 4.435 99.600 5.075 ;
        RECT 99.950 4.775 100.120 5.105 ;
        RECT 100.910 4.905 101.560 5.075 ;
        RECT 101.270 4.515 101.560 4.905 ;
        RECT 102.270 4.905 102.560 5.075 ;
        RECT 99.070 4.115 99.240 4.345 ;
        RECT 99.950 4.375 100.120 4.515 ;
        RECT 101.390 4.435 101.560 4.515 ;
        RECT 99.950 4.205 100.840 4.375 ;
        RECT 101.910 4.345 102.080 4.765 ;
        RECT 102.270 4.515 102.440 4.905 ;
        RECT 103.110 4.515 104.080 4.685 ;
        RECT 102.270 4.345 102.560 4.515 ;
        RECT 103.110 4.345 103.280 4.515 ;
        RECT 96.670 3.865 97.160 4.035 ;
        RECT 97.510 3.865 98.000 4.035 ;
        RECT 96.990 3.785 97.160 3.865 ;
        RECT 98.230 3.785 98.400 4.115 ;
        RECT 98.710 3.785 98.880 4.115 ;
        RECT 99.070 3.865 99.360 4.115 ;
        RECT 99.190 3.785 99.360 3.865 ;
        RECT 99.950 3.865 100.440 4.035 ;
        RECT 99.950 3.785 100.120 3.865 ;
        RECT 100.670 3.785 100.840 4.205 ;
        RECT 101.390 4.135 101.560 4.235 ;
        RECT 101.150 4.035 101.560 4.135 ;
        RECT 102.270 4.035 102.440 4.345 ;
        RECT 101.070 3.965 101.560 4.035 ;
        RECT 101.070 3.865 101.400 3.965 ;
        RECT 102.070 3.865 102.440 4.035 ;
        RECT 102.630 4.035 102.800 4.115 ;
        RECT 102.630 3.865 103.360 4.035 ;
        RECT 102.630 3.785 102.800 3.865 ;
        RECT 103.590 3.785 103.760 4.235 ;
        RECT 106.315 3.895 106.490 5.155 ;
        RECT 106.840 4.095 107.010 5.155 ;
        RECT 106.840 3.925 107.070 4.095 ;
        RECT 90.500 3.575 90.670 3.625 ;
        RECT 91.120 3.210 91.290 3.625 ;
        RECT 106.315 3.695 106.485 3.895 ;
        RECT 90.130 3.175 90.600 3.205 ;
        RECT 90.070 3.035 90.600 3.175 ;
        RECT 91.120 3.040 91.590 3.210 ;
        RECT 93.110 3.045 93.280 3.395 ;
        RECT 94.070 3.295 94.240 3.395 ;
        RECT 96.510 3.295 96.680 3.395 ;
        RECT 97.990 3.295 98.160 3.395 ;
        RECT 94.070 3.125 94.800 3.295 ;
        RECT 95.950 3.125 96.680 3.295 ;
        RECT 97.430 3.125 98.160 3.295 ;
        RECT 98.950 3.045 99.120 3.395 ;
        RECT 99.950 3.045 100.120 3.395 ;
        RECT 100.910 3.045 101.080 3.395 ;
        RECT 102.390 3.045 102.560 3.395 ;
        RECT 103.350 3.045 103.520 3.395 ;
        RECT 106.315 3.365 106.725 3.695 ;
        RECT 90.070 2.945 90.300 3.035 ;
        RECT 106.315 2.855 106.485 3.365 ;
        RECT 106.315 2.525 106.725 2.855 ;
        RECT 88.280 2.145 88.510 2.315 ;
        RECT 88.280 1.865 88.450 2.145 ;
        RECT 88.710 1.865 88.885 2.375 ;
        RECT 89.140 1.865 89.315 2.415 ;
        RECT 90.505 1.865 90.675 2.375 ;
        RECT 106.315 2.355 106.485 2.525 ;
        RECT 106.315 1.865 106.490 2.355 ;
        RECT 106.900 2.315 107.070 3.925 ;
        RECT 107.270 3.895 107.445 5.155 ;
        RECT 107.700 4.015 107.875 5.155 ;
        RECT 107.270 2.945 107.440 3.895 ;
        RECT 107.700 2.415 107.870 4.015 ;
        RECT 109.060 4.010 109.235 5.155 ;
        RECT 108.690 3.205 108.860 3.895 ;
        RECT 109.060 3.805 109.230 4.010 ;
        RECT 109.680 3.805 109.850 3.900 ;
        RECT 109.060 3.625 109.850 3.805 ;
        RECT 109.060 3.575 109.230 3.625 ;
        RECT 109.680 3.210 109.850 3.625 ;
        RECT 108.690 3.175 109.160 3.205 ;
        RECT 108.630 3.035 109.160 3.175 ;
        RECT 109.680 3.040 110.150 3.210 ;
        RECT 108.630 2.945 108.860 3.035 ;
        RECT 106.840 2.145 107.070 2.315 ;
        RECT 106.840 1.865 107.010 2.145 ;
        RECT 107.270 1.865 107.445 2.375 ;
        RECT 107.700 1.865 107.875 2.415 ;
        RECT 109.065 1.865 109.235 2.375 ;
      LAYER met1 ;
        RECT 16.540 10.060 16.830 10.290 ;
        RECT 27.355 10.060 27.645 10.290 ;
        RECT 32.970 10.060 33.260 10.290 ;
        RECT 16.600 9.610 16.770 10.060 ;
        RECT 27.415 9.715 27.585 10.060 ;
        RECT 16.510 9.320 16.860 9.610 ;
        RECT 27.315 9.345 27.695 9.715 ;
        RECT 33.030 9.580 33.200 10.060 ;
        RECT 34.760 10.030 35.055 10.290 ;
        RECT 34.390 9.635 34.620 9.660 ;
        RECT 34.360 9.580 34.650 9.635 ;
        RECT 33.030 9.550 34.650 9.580 ;
        RECT 32.970 9.410 34.650 9.550 ;
        RECT 27.355 9.320 27.645 9.345 ;
        RECT 32.970 9.320 33.260 9.410 ;
        RECT 34.360 9.335 34.650 9.410 ;
        RECT 34.390 9.310 34.620 9.335 ;
        RECT 27.990 9.180 28.340 9.245 ;
        RECT 33.425 9.180 33.750 9.270 ;
        RECT 27.785 9.150 28.340 9.180 ;
        RECT 33.400 9.150 33.750 9.180 ;
        RECT 27.615 9.145 28.340 9.150 ;
        RECT 33.230 9.145 33.750 9.150 ;
        RECT 27.615 8.975 33.750 9.145 ;
        RECT 27.785 8.950 28.340 8.975 ;
        RECT 33.400 8.950 33.750 8.975 ;
        RECT 27.990 8.895 28.340 8.950 ;
        RECT 33.425 8.945 33.750 8.950 ;
        RECT 34.820 8.930 34.990 10.030 ;
        RECT 35.755 10.025 36.050 10.285 ;
        RECT 45.915 10.060 46.205 10.290 ;
        RECT 51.530 10.060 51.820 10.290 ;
        RECT 35.815 9.295 35.985 10.025 ;
        RECT 45.975 9.715 46.145 10.060 ;
        RECT 45.875 9.345 46.255 9.715 ;
        RECT 51.590 9.580 51.760 10.060 ;
        RECT 53.320 10.030 53.615 10.290 ;
        RECT 52.950 9.635 53.180 9.660 ;
        RECT 52.920 9.580 53.210 9.635 ;
        RECT 51.590 9.550 53.210 9.580 ;
        RECT 51.530 9.410 53.210 9.550 ;
        RECT 45.915 9.320 46.205 9.345 ;
        RECT 51.530 9.320 51.820 9.410 ;
        RECT 52.920 9.335 53.210 9.410 ;
        RECT 52.950 9.310 53.180 9.335 ;
        RECT 34.760 8.925 34.990 8.930 ;
        RECT 35.805 8.945 36.155 9.295 ;
        RECT 46.550 9.180 46.900 9.250 ;
        RECT 51.985 9.180 52.310 9.270 ;
        RECT 46.345 9.150 46.900 9.180 ;
        RECT 51.960 9.150 52.310 9.180 ;
        RECT 46.175 9.145 46.900 9.150 ;
        RECT 51.790 9.145 52.310 9.150 ;
        RECT 46.175 8.975 52.310 9.145 ;
        RECT 46.345 8.950 46.900 8.975 ;
        RECT 51.960 8.950 52.310 8.975 ;
        RECT 35.805 8.925 36.105 8.945 ;
        RECT 16.135 8.790 16.485 8.865 ;
        RECT 32.625 8.820 32.945 8.835 ;
        RECT 32.600 8.790 32.945 8.820 ;
        RECT 15.995 8.620 16.485 8.790 ;
        RECT 32.425 8.620 32.945 8.790 ;
        RECT 34.760 8.690 35.050 8.925 ;
        RECT 35.755 8.855 36.105 8.925 ;
        RECT 46.550 8.900 46.900 8.950 ;
        RECT 51.985 8.945 52.310 8.950 ;
        RECT 53.380 8.930 53.550 10.030 ;
        RECT 54.315 10.025 54.610 10.285 ;
        RECT 64.475 10.060 64.765 10.290 ;
        RECT 70.090 10.060 70.380 10.290 ;
        RECT 54.375 9.305 54.545 10.025 ;
        RECT 64.535 9.715 64.705 10.060 ;
        RECT 64.435 9.345 64.815 9.715 ;
        RECT 70.150 9.580 70.320 10.060 ;
        RECT 71.880 10.030 72.175 10.290 ;
        RECT 71.510 9.635 71.740 9.660 ;
        RECT 71.480 9.580 71.770 9.635 ;
        RECT 70.150 9.550 71.770 9.580 ;
        RECT 70.090 9.410 71.770 9.550 ;
        RECT 64.475 9.320 64.765 9.345 ;
        RECT 70.090 9.320 70.380 9.410 ;
        RECT 71.480 9.335 71.770 9.410 ;
        RECT 71.510 9.310 71.740 9.335 ;
        RECT 53.320 8.925 53.550 8.930 ;
        RECT 54.360 8.950 54.715 9.305 ;
        RECT 65.105 9.180 65.455 9.255 ;
        RECT 70.545 9.180 70.870 9.270 ;
        RECT 64.905 9.150 65.455 9.180 ;
        RECT 70.520 9.150 70.870 9.180 ;
        RECT 64.735 9.145 65.455 9.150 ;
        RECT 70.350 9.145 70.870 9.150 ;
        RECT 64.735 8.975 70.870 9.145 ;
        RECT 64.905 8.950 65.455 8.975 ;
        RECT 70.520 8.950 70.870 8.975 ;
        RECT 54.360 8.925 54.665 8.950 ;
        RECT 35.755 8.685 36.045 8.855 ;
        RECT 51.185 8.820 51.505 8.835 ;
        RECT 51.160 8.790 51.505 8.820 ;
        RECT 50.985 8.620 51.505 8.790 ;
        RECT 53.320 8.690 53.610 8.925 ;
        RECT 54.315 8.850 54.665 8.925 ;
        RECT 65.105 8.905 65.455 8.950 ;
        RECT 70.545 8.945 70.870 8.950 ;
        RECT 71.940 8.930 72.110 10.030 ;
        RECT 72.875 10.025 73.170 10.285 ;
        RECT 83.035 10.060 83.325 10.290 ;
        RECT 88.650 10.060 88.940 10.290 ;
        RECT 72.935 9.295 73.105 10.025 ;
        RECT 83.095 9.715 83.265 10.060 ;
        RECT 82.995 9.345 83.375 9.715 ;
        RECT 88.710 9.580 88.880 10.060 ;
        RECT 90.440 10.030 90.735 10.290 ;
        RECT 90.070 9.635 90.300 9.660 ;
        RECT 90.040 9.580 90.330 9.635 ;
        RECT 88.710 9.550 90.330 9.580 ;
        RECT 88.650 9.410 90.330 9.550 ;
        RECT 83.035 9.320 83.325 9.345 ;
        RECT 88.650 9.320 88.940 9.410 ;
        RECT 90.040 9.335 90.330 9.410 ;
        RECT 90.070 9.310 90.300 9.335 ;
        RECT 71.880 8.925 72.110 8.930 ;
        RECT 72.880 8.945 73.230 9.295 ;
        RECT 83.665 9.180 84.015 9.250 ;
        RECT 89.105 9.180 89.430 9.270 ;
        RECT 83.465 9.150 84.015 9.180 ;
        RECT 89.080 9.150 89.430 9.180 ;
        RECT 83.295 9.145 84.015 9.150 ;
        RECT 88.910 9.145 89.430 9.150 ;
        RECT 83.295 8.975 89.430 9.145 ;
        RECT 83.465 8.950 84.015 8.975 ;
        RECT 89.080 8.950 89.430 8.975 ;
        RECT 72.880 8.925 73.225 8.945 ;
        RECT 54.315 8.685 54.605 8.850 ;
        RECT 69.745 8.820 70.065 8.835 ;
        RECT 69.720 8.790 70.065 8.820 ;
        RECT 69.545 8.620 70.065 8.790 ;
        RECT 71.880 8.690 72.170 8.925 ;
        RECT 72.875 8.855 73.225 8.925 ;
        RECT 83.665 8.900 84.015 8.950 ;
        RECT 89.105 8.945 89.430 8.950 ;
        RECT 90.500 8.930 90.670 10.030 ;
        RECT 91.435 10.025 91.730 10.285 ;
        RECT 101.595 10.060 101.885 10.290 ;
        RECT 107.210 10.060 107.500 10.290 ;
        RECT 91.495 9.295 91.665 10.025 ;
        RECT 101.655 9.715 101.825 10.060 ;
        RECT 101.555 9.345 101.935 9.715 ;
        RECT 107.270 9.580 107.440 10.060 ;
        RECT 109.000 10.030 109.295 10.290 ;
        RECT 108.630 9.635 108.860 9.660 ;
        RECT 108.600 9.580 108.890 9.635 ;
        RECT 107.270 9.550 108.890 9.580 ;
        RECT 107.210 9.410 108.890 9.550 ;
        RECT 101.595 9.320 101.885 9.345 ;
        RECT 107.210 9.320 107.500 9.410 ;
        RECT 108.600 9.335 108.890 9.410 ;
        RECT 108.630 9.310 108.860 9.335 ;
        RECT 90.440 8.925 90.670 8.930 ;
        RECT 91.440 8.945 91.790 9.295 ;
        RECT 102.225 9.180 102.575 9.250 ;
        RECT 107.665 9.180 107.990 9.270 ;
        RECT 102.025 9.150 102.575 9.180 ;
        RECT 107.640 9.150 107.990 9.180 ;
        RECT 101.855 9.145 102.575 9.150 ;
        RECT 107.470 9.145 107.990 9.150 ;
        RECT 101.855 8.975 107.990 9.145 ;
        RECT 102.025 8.950 102.575 8.975 ;
        RECT 107.640 8.950 107.990 8.975 ;
        RECT 91.440 8.925 91.785 8.945 ;
        RECT 72.875 8.685 73.165 8.855 ;
        RECT 88.305 8.820 88.625 8.835 ;
        RECT 88.280 8.790 88.625 8.820 ;
        RECT 88.105 8.620 88.625 8.790 ;
        RECT 90.440 8.690 90.730 8.925 ;
        RECT 91.435 8.855 91.785 8.925 ;
        RECT 102.225 8.900 102.575 8.950 ;
        RECT 107.665 8.945 107.990 8.950 ;
        RECT 109.060 8.930 109.230 10.030 ;
        RECT 109.995 10.025 110.290 10.285 ;
        RECT 110.025 10.000 110.290 10.025 ;
        RECT 110.025 9.915 110.350 10.000 ;
        RECT 110.025 9.565 110.375 9.915 ;
        RECT 109.000 8.925 109.230 8.930 ;
        RECT 110.055 8.925 110.225 9.565 ;
        RECT 91.435 8.685 91.725 8.855 ;
        RECT 106.865 8.820 107.185 8.835 ;
        RECT 106.840 8.790 107.185 8.820 ;
        RECT 106.665 8.620 107.185 8.790 ;
        RECT 109.000 8.690 109.290 8.925 ;
        RECT 109.995 8.920 110.225 8.925 ;
        RECT 109.995 8.685 110.285 8.920 ;
        RECT 16.135 8.575 16.485 8.620 ;
        RECT 32.600 8.590 32.945 8.620 ;
        RECT 51.160 8.590 51.505 8.620 ;
        RECT 69.720 8.590 70.065 8.620 ;
        RECT 88.280 8.590 88.625 8.620 ;
        RECT 106.840 8.590 107.185 8.620 ;
        RECT 32.625 8.545 32.945 8.590 ;
        RECT 51.185 8.545 51.505 8.590 ;
        RECT 69.745 8.545 70.065 8.590 ;
        RECT 88.305 8.545 88.625 8.590 ;
        RECT 106.865 8.545 107.185 8.590 ;
        RECT 23.550 5.065 23.870 5.125 ;
        RECT 18.790 4.555 19.110 4.965 ;
        RECT 23.550 4.925 24.620 5.065 ;
        RECT 21.800 4.825 22.900 4.895 ;
        RECT 23.550 4.865 23.870 4.925 ;
        RECT 21.730 4.755 22.980 4.825 ;
        RECT 21.730 4.595 22.020 4.755 ;
        RECT 22.690 4.595 22.980 4.755 ;
        RECT 18.870 3.425 19.030 4.555 ;
        RECT 19.750 4.305 20.070 4.565 ;
        RECT 20.870 4.445 21.190 4.565 ;
        RECT 22.210 4.505 22.500 4.545 ;
        RECT 20.870 4.305 21.700 4.445 ;
        RECT 22.210 4.315 22.540 4.505 ;
        RECT 21.490 4.265 21.700 4.305 ;
        RECT 21.490 4.035 21.780 4.265 ;
        RECT 19.270 3.985 19.590 4.005 ;
        RECT 19.270 3.845 20.220 3.985 ;
        RECT 20.680 3.945 20.970 3.985 ;
        RECT 19.270 3.755 19.820 3.845 ;
        RECT 20.080 3.805 20.220 3.845 ;
        RECT 20.580 3.805 20.970 3.945 ;
        RECT 20.080 3.755 20.970 3.805 ;
        RECT 19.270 3.745 19.590 3.755 ;
        RECT 20.080 3.665 20.720 3.755 ;
        RECT 18.810 3.195 19.100 3.425 ;
        RECT 19.750 3.385 20.070 3.445 ;
        RECT 21.710 3.385 22.030 3.445 ;
        RECT 22.400 3.425 22.540 4.315 ;
        RECT 23.190 4.305 23.510 4.565 ;
        RECT 23.910 4.305 24.230 4.565 ;
        RECT 24.480 4.505 24.620 4.925 ;
        RECT 25.110 4.865 25.430 5.125 ;
        RECT 25.650 5.065 25.940 5.105 ;
        RECT 26.110 5.065 26.430 5.125 ;
        RECT 25.650 4.925 26.430 5.065 ;
        RECT 25.650 4.875 25.940 4.925 ;
        RECT 26.110 4.865 26.430 4.925 ;
        RECT 26.590 4.865 26.910 5.125 ;
        RECT 27.070 4.865 27.390 5.125 ;
        RECT 28.070 4.895 28.390 5.125 ;
        RECT 42.110 5.065 42.430 5.125 ;
        RECT 28.070 4.865 29.500 4.895 ;
        RECT 28.160 4.755 29.500 4.865 ;
        RECT 25.650 4.505 25.940 4.545 ;
        RECT 24.480 4.365 25.940 4.505 ;
        RECT 25.650 4.315 25.940 4.365 ;
        RECT 27.590 4.305 27.910 4.565 ;
        RECT 28.160 4.545 28.300 4.755 ;
        RECT 28.090 4.315 28.380 4.545 ;
        RECT 28.810 4.505 29.100 4.545 ;
        RECT 28.810 4.315 29.140 4.505 ;
        RECT 27.090 4.225 27.380 4.265 ;
        RECT 27.590 4.225 27.820 4.305 ;
        RECT 27.090 4.085 27.820 4.225 ;
        RECT 27.090 4.035 27.380 4.085 ;
        RECT 22.930 3.985 23.250 4.005 ;
        RECT 22.690 3.945 23.250 3.985 ;
        RECT 23.930 3.945 24.220 3.985 ;
        RECT 22.690 3.805 24.220 3.945 ;
        RECT 22.690 3.755 23.250 3.805 ;
        RECT 23.930 3.755 24.220 3.805 ;
        RECT 24.410 3.945 24.700 3.985 ;
        RECT 24.410 3.805 25.340 3.945 ;
        RECT 24.410 3.755 24.700 3.805 ;
        RECT 22.930 3.745 23.250 3.755 ;
        RECT 19.750 3.245 22.030 3.385 ;
        RECT 19.750 3.185 20.070 3.245 ;
        RECT 21.710 3.185 22.030 3.245 ;
        RECT 22.210 3.385 22.540 3.425 ;
        RECT 23.190 3.385 23.510 3.445 ;
        RECT 23.910 3.425 24.230 3.445 ;
        RECT 22.210 3.245 23.510 3.385 ;
        RECT 22.210 3.195 22.500 3.245 ;
        RECT 23.190 3.185 23.510 3.245 ;
        RECT 23.690 3.195 24.230 3.425 ;
        RECT 23.910 3.185 24.230 3.195 ;
        RECT 24.630 3.185 24.950 3.445 ;
        RECT 25.200 3.385 25.340 3.805 ;
        RECT 25.630 3.805 25.950 4.005 ;
        RECT 28.330 3.805 28.620 3.985 ;
        RECT 25.630 3.755 28.620 3.805 ;
        RECT 25.630 3.745 28.540 3.755 ;
        RECT 25.720 3.665 28.540 3.745 ;
        RECT 29.000 3.445 29.140 4.315 ;
        RECT 29.360 4.265 29.500 4.755 ;
        RECT 31.020 4.445 31.360 4.795 ;
        RECT 37.350 4.555 37.670 4.965 ;
        RECT 42.110 4.925 43.180 5.065 ;
        RECT 40.360 4.825 41.460 4.895 ;
        RECT 42.110 4.865 42.430 4.925 ;
        RECT 40.290 4.755 41.540 4.825 ;
        RECT 40.290 4.595 40.580 4.755 ;
        RECT 41.250 4.595 41.540 4.755 ;
        RECT 29.290 4.035 29.580 4.265 ;
        RECT 31.110 3.490 31.280 4.445 ;
        RECT 32.625 3.875 32.945 3.980 ;
        RECT 32.600 3.860 32.945 3.875 ;
        RECT 32.595 3.845 32.945 3.860 ;
        RECT 32.425 3.675 32.945 3.845 ;
        RECT 32.600 3.660 32.945 3.675 ;
        RECT 32.600 3.645 32.890 3.660 ;
        RECT 33.400 3.490 33.750 3.610 ;
        RECT 34.760 3.540 35.050 3.775 ;
        RECT 34.760 3.535 34.990 3.540 ;
        RECT 25.870 3.425 26.190 3.445 ;
        RECT 25.650 3.385 26.190 3.425 ;
        RECT 25.200 3.245 26.190 3.385 ;
        RECT 25.650 3.195 26.190 3.245 ;
        RECT 25.870 3.185 26.190 3.195 ;
        RECT 26.470 3.185 27.150 3.445 ;
        RECT 27.590 3.385 27.910 3.445 ;
        RECT 28.090 3.385 28.380 3.425 ;
        RECT 27.590 3.245 28.380 3.385 ;
        RECT 29.000 3.245 29.350 3.445 ;
        RECT 31.110 3.320 33.750 3.490 ;
        RECT 33.230 3.315 33.750 3.320 ;
        RECT 33.400 3.260 33.750 3.315 ;
        RECT 27.590 3.185 27.910 3.245 ;
        RECT 28.090 3.195 28.380 3.245 ;
        RECT 29.030 3.185 29.350 3.245 ;
        RECT 34.390 3.220 34.620 3.235 ;
        RECT 32.970 3.120 33.260 3.145 ;
        RECT 34.360 3.120 34.655 3.220 ;
        RECT 32.970 2.950 34.655 3.120 ;
        RECT 32.970 2.915 33.260 2.950 ;
        RECT 33.030 2.405 33.200 2.915 ;
        RECT 34.360 2.900 34.655 2.950 ;
        RECT 34.390 2.885 34.620 2.900 ;
        RECT 34.820 2.435 34.990 3.535 ;
        RECT 37.430 3.425 37.590 4.555 ;
        RECT 38.310 4.305 38.630 4.565 ;
        RECT 39.430 4.445 39.750 4.565 ;
        RECT 40.770 4.505 41.060 4.545 ;
        RECT 39.430 4.305 40.260 4.445 ;
        RECT 40.770 4.315 41.100 4.505 ;
        RECT 40.050 4.265 40.260 4.305 ;
        RECT 40.050 4.035 40.340 4.265 ;
        RECT 37.830 3.985 38.150 4.005 ;
        RECT 37.830 3.845 38.780 3.985 ;
        RECT 39.240 3.945 39.530 3.985 ;
        RECT 37.830 3.755 38.380 3.845 ;
        RECT 38.640 3.805 38.780 3.845 ;
        RECT 39.140 3.805 39.530 3.945 ;
        RECT 38.640 3.755 39.530 3.805 ;
        RECT 37.830 3.745 38.150 3.755 ;
        RECT 38.640 3.665 39.280 3.755 ;
        RECT 37.370 3.195 37.660 3.425 ;
        RECT 38.310 3.385 38.630 3.445 ;
        RECT 40.270 3.385 40.590 3.445 ;
        RECT 40.960 3.425 41.100 4.315 ;
        RECT 41.750 4.305 42.070 4.565 ;
        RECT 42.470 4.305 42.790 4.565 ;
        RECT 43.040 4.505 43.180 4.925 ;
        RECT 43.670 4.865 43.990 5.125 ;
        RECT 44.210 5.065 44.500 5.105 ;
        RECT 44.670 5.065 44.990 5.125 ;
        RECT 44.210 4.925 44.990 5.065 ;
        RECT 44.210 4.875 44.500 4.925 ;
        RECT 44.670 4.865 44.990 4.925 ;
        RECT 45.150 4.865 45.470 5.125 ;
        RECT 45.630 4.865 45.950 5.125 ;
        RECT 46.630 4.895 46.950 5.125 ;
        RECT 60.670 5.065 60.990 5.125 ;
        RECT 46.630 4.865 48.060 4.895 ;
        RECT 46.720 4.755 48.060 4.865 ;
        RECT 44.210 4.505 44.500 4.545 ;
        RECT 43.040 4.365 44.500 4.505 ;
        RECT 44.210 4.315 44.500 4.365 ;
        RECT 46.150 4.305 46.470 4.565 ;
        RECT 46.720 4.545 46.860 4.755 ;
        RECT 46.650 4.315 46.940 4.545 ;
        RECT 47.370 4.505 47.660 4.545 ;
        RECT 47.370 4.315 47.700 4.505 ;
        RECT 45.650 4.225 45.940 4.265 ;
        RECT 46.150 4.225 46.380 4.305 ;
        RECT 45.650 4.085 46.380 4.225 ;
        RECT 45.650 4.035 45.940 4.085 ;
        RECT 41.490 3.985 41.810 4.005 ;
        RECT 41.250 3.945 41.810 3.985 ;
        RECT 42.490 3.945 42.780 3.985 ;
        RECT 41.250 3.805 42.780 3.945 ;
        RECT 41.250 3.755 41.810 3.805 ;
        RECT 42.490 3.755 42.780 3.805 ;
        RECT 42.970 3.945 43.260 3.985 ;
        RECT 42.970 3.805 43.900 3.945 ;
        RECT 42.970 3.755 43.260 3.805 ;
        RECT 41.490 3.745 41.810 3.755 ;
        RECT 38.310 3.245 40.590 3.385 ;
        RECT 38.310 3.185 38.630 3.245 ;
        RECT 40.270 3.185 40.590 3.245 ;
        RECT 40.770 3.385 41.100 3.425 ;
        RECT 41.750 3.385 42.070 3.445 ;
        RECT 42.470 3.425 42.790 3.445 ;
        RECT 40.770 3.245 42.070 3.385 ;
        RECT 40.770 3.195 41.060 3.245 ;
        RECT 41.750 3.185 42.070 3.245 ;
        RECT 42.250 3.195 42.790 3.425 ;
        RECT 42.470 3.185 42.790 3.195 ;
        RECT 43.190 3.185 43.510 3.445 ;
        RECT 43.760 3.385 43.900 3.805 ;
        RECT 44.190 3.805 44.510 4.005 ;
        RECT 46.890 3.805 47.180 3.985 ;
        RECT 44.190 3.755 47.180 3.805 ;
        RECT 44.190 3.745 47.100 3.755 ;
        RECT 44.280 3.665 47.100 3.745 ;
        RECT 47.560 3.445 47.700 4.315 ;
        RECT 47.920 4.265 48.060 4.755 ;
        RECT 49.580 4.445 49.920 4.795 ;
        RECT 55.910 4.555 56.230 4.965 ;
        RECT 60.670 4.925 61.740 5.065 ;
        RECT 58.920 4.825 60.020 4.895 ;
        RECT 60.670 4.865 60.990 4.925 ;
        RECT 58.850 4.755 60.100 4.825 ;
        RECT 58.850 4.595 59.140 4.755 ;
        RECT 59.810 4.595 60.100 4.755 ;
        RECT 47.850 4.035 48.140 4.265 ;
        RECT 49.670 3.490 49.840 4.445 ;
        RECT 51.185 3.875 51.505 3.980 ;
        RECT 51.160 3.860 51.505 3.875 ;
        RECT 51.155 3.845 51.505 3.860 ;
        RECT 50.985 3.675 51.505 3.845 ;
        RECT 51.160 3.660 51.505 3.675 ;
        RECT 51.160 3.645 51.450 3.660 ;
        RECT 51.960 3.490 52.310 3.610 ;
        RECT 53.320 3.540 53.610 3.775 ;
        RECT 53.320 3.535 53.550 3.540 ;
        RECT 44.430 3.425 44.750 3.445 ;
        RECT 44.210 3.385 44.750 3.425 ;
        RECT 43.760 3.245 44.750 3.385 ;
        RECT 44.210 3.195 44.750 3.245 ;
        RECT 44.430 3.185 44.750 3.195 ;
        RECT 45.030 3.185 45.710 3.445 ;
        RECT 46.150 3.385 46.470 3.445 ;
        RECT 46.650 3.385 46.940 3.425 ;
        RECT 46.150 3.245 46.940 3.385 ;
        RECT 47.560 3.245 47.910 3.445 ;
        RECT 49.670 3.320 52.310 3.490 ;
        RECT 51.790 3.315 52.310 3.320 ;
        RECT 51.960 3.260 52.310 3.315 ;
        RECT 46.150 3.185 46.470 3.245 ;
        RECT 46.650 3.195 46.940 3.245 ;
        RECT 47.590 3.185 47.910 3.245 ;
        RECT 52.950 3.220 53.180 3.235 ;
        RECT 51.530 3.120 51.820 3.145 ;
        RECT 52.920 3.120 53.215 3.220 ;
        RECT 51.530 2.950 53.215 3.120 ;
        RECT 51.530 2.915 51.820 2.950 ;
        RECT 32.970 2.175 33.260 2.405 ;
        RECT 34.760 2.175 35.055 2.435 ;
        RECT 51.590 2.405 51.760 2.915 ;
        RECT 52.920 2.900 53.215 2.950 ;
        RECT 52.950 2.885 53.180 2.900 ;
        RECT 53.380 2.435 53.550 3.535 ;
        RECT 55.990 3.425 56.150 4.555 ;
        RECT 56.870 4.305 57.190 4.565 ;
        RECT 57.990 4.445 58.310 4.565 ;
        RECT 59.330 4.505 59.620 4.545 ;
        RECT 57.990 4.305 58.820 4.445 ;
        RECT 59.330 4.315 59.660 4.505 ;
        RECT 58.610 4.265 58.820 4.305 ;
        RECT 58.610 4.035 58.900 4.265 ;
        RECT 56.390 3.985 56.710 4.005 ;
        RECT 56.390 3.845 57.340 3.985 ;
        RECT 57.800 3.945 58.090 3.985 ;
        RECT 56.390 3.755 56.940 3.845 ;
        RECT 57.200 3.805 57.340 3.845 ;
        RECT 57.700 3.805 58.090 3.945 ;
        RECT 57.200 3.755 58.090 3.805 ;
        RECT 56.390 3.745 56.710 3.755 ;
        RECT 57.200 3.665 57.840 3.755 ;
        RECT 55.930 3.195 56.220 3.425 ;
        RECT 56.870 3.385 57.190 3.445 ;
        RECT 58.830 3.385 59.150 3.445 ;
        RECT 59.520 3.425 59.660 4.315 ;
        RECT 60.310 4.305 60.630 4.565 ;
        RECT 61.030 4.305 61.350 4.565 ;
        RECT 61.600 4.505 61.740 4.925 ;
        RECT 62.230 4.865 62.550 5.125 ;
        RECT 62.770 5.065 63.060 5.105 ;
        RECT 63.230 5.065 63.550 5.125 ;
        RECT 62.770 4.925 63.550 5.065 ;
        RECT 62.770 4.875 63.060 4.925 ;
        RECT 63.230 4.865 63.550 4.925 ;
        RECT 63.710 4.865 64.030 5.125 ;
        RECT 64.190 4.865 64.510 5.125 ;
        RECT 65.190 4.895 65.510 5.125 ;
        RECT 79.230 5.065 79.550 5.125 ;
        RECT 65.190 4.865 66.620 4.895 ;
        RECT 65.280 4.755 66.620 4.865 ;
        RECT 62.770 4.505 63.060 4.545 ;
        RECT 61.600 4.365 63.060 4.505 ;
        RECT 62.770 4.315 63.060 4.365 ;
        RECT 64.710 4.305 65.030 4.565 ;
        RECT 65.280 4.545 65.420 4.755 ;
        RECT 65.210 4.315 65.500 4.545 ;
        RECT 65.930 4.505 66.220 4.545 ;
        RECT 65.930 4.315 66.260 4.505 ;
        RECT 64.210 4.225 64.500 4.265 ;
        RECT 64.710 4.225 64.940 4.305 ;
        RECT 64.210 4.085 64.940 4.225 ;
        RECT 64.210 4.035 64.500 4.085 ;
        RECT 60.050 3.985 60.370 4.005 ;
        RECT 59.810 3.945 60.370 3.985 ;
        RECT 61.050 3.945 61.340 3.985 ;
        RECT 59.810 3.805 61.340 3.945 ;
        RECT 59.810 3.755 60.370 3.805 ;
        RECT 61.050 3.755 61.340 3.805 ;
        RECT 61.530 3.945 61.820 3.985 ;
        RECT 61.530 3.805 62.460 3.945 ;
        RECT 61.530 3.755 61.820 3.805 ;
        RECT 60.050 3.745 60.370 3.755 ;
        RECT 56.870 3.245 59.150 3.385 ;
        RECT 56.870 3.185 57.190 3.245 ;
        RECT 58.830 3.185 59.150 3.245 ;
        RECT 59.330 3.385 59.660 3.425 ;
        RECT 60.310 3.385 60.630 3.445 ;
        RECT 61.030 3.425 61.350 3.445 ;
        RECT 59.330 3.245 60.630 3.385 ;
        RECT 59.330 3.195 59.620 3.245 ;
        RECT 60.310 3.185 60.630 3.245 ;
        RECT 60.810 3.195 61.350 3.425 ;
        RECT 61.030 3.185 61.350 3.195 ;
        RECT 61.750 3.185 62.070 3.445 ;
        RECT 62.320 3.385 62.460 3.805 ;
        RECT 62.750 3.805 63.070 4.005 ;
        RECT 65.450 3.805 65.740 3.985 ;
        RECT 62.750 3.755 65.740 3.805 ;
        RECT 62.750 3.745 65.660 3.755 ;
        RECT 62.840 3.665 65.660 3.745 ;
        RECT 66.120 3.445 66.260 4.315 ;
        RECT 66.480 4.265 66.620 4.755 ;
        RECT 68.140 4.445 68.480 4.795 ;
        RECT 74.470 4.555 74.790 4.965 ;
        RECT 79.230 4.925 80.300 5.065 ;
        RECT 77.480 4.825 78.580 4.895 ;
        RECT 79.230 4.865 79.550 4.925 ;
        RECT 77.410 4.755 78.660 4.825 ;
        RECT 77.410 4.595 77.700 4.755 ;
        RECT 78.370 4.595 78.660 4.755 ;
        RECT 66.410 4.035 66.700 4.265 ;
        RECT 68.230 3.490 68.400 4.445 ;
        RECT 69.745 3.875 70.065 3.980 ;
        RECT 69.720 3.860 70.065 3.875 ;
        RECT 69.715 3.845 70.065 3.860 ;
        RECT 69.545 3.675 70.065 3.845 ;
        RECT 69.720 3.660 70.065 3.675 ;
        RECT 69.720 3.645 70.010 3.660 ;
        RECT 70.520 3.490 70.870 3.610 ;
        RECT 71.880 3.540 72.170 3.775 ;
        RECT 71.880 3.535 72.110 3.540 ;
        RECT 62.990 3.425 63.310 3.445 ;
        RECT 62.770 3.385 63.310 3.425 ;
        RECT 62.320 3.245 63.310 3.385 ;
        RECT 62.770 3.195 63.310 3.245 ;
        RECT 62.990 3.185 63.310 3.195 ;
        RECT 63.590 3.185 64.270 3.445 ;
        RECT 64.710 3.385 65.030 3.445 ;
        RECT 65.210 3.385 65.500 3.425 ;
        RECT 64.710 3.245 65.500 3.385 ;
        RECT 66.120 3.245 66.470 3.445 ;
        RECT 68.230 3.320 70.870 3.490 ;
        RECT 70.350 3.315 70.870 3.320 ;
        RECT 70.520 3.260 70.870 3.315 ;
        RECT 64.710 3.185 65.030 3.245 ;
        RECT 65.210 3.195 65.500 3.245 ;
        RECT 66.150 3.185 66.470 3.245 ;
        RECT 71.510 3.220 71.740 3.235 ;
        RECT 70.090 3.120 70.380 3.145 ;
        RECT 71.480 3.120 71.775 3.220 ;
        RECT 70.090 2.950 71.775 3.120 ;
        RECT 70.090 2.915 70.380 2.950 ;
        RECT 51.530 2.175 51.820 2.405 ;
        RECT 53.320 2.175 53.615 2.435 ;
        RECT 70.150 2.405 70.320 2.915 ;
        RECT 71.480 2.900 71.775 2.950 ;
        RECT 71.510 2.885 71.740 2.900 ;
        RECT 71.940 2.435 72.110 3.535 ;
        RECT 74.550 3.425 74.710 4.555 ;
        RECT 75.430 4.305 75.750 4.565 ;
        RECT 76.550 4.445 76.870 4.565 ;
        RECT 77.890 4.505 78.180 4.545 ;
        RECT 76.550 4.305 77.380 4.445 ;
        RECT 77.890 4.315 78.220 4.505 ;
        RECT 77.170 4.265 77.380 4.305 ;
        RECT 77.170 4.035 77.460 4.265 ;
        RECT 74.950 3.985 75.270 4.005 ;
        RECT 74.950 3.845 75.900 3.985 ;
        RECT 76.360 3.945 76.650 3.985 ;
        RECT 74.950 3.755 75.500 3.845 ;
        RECT 75.760 3.805 75.900 3.845 ;
        RECT 76.260 3.805 76.650 3.945 ;
        RECT 75.760 3.755 76.650 3.805 ;
        RECT 74.950 3.745 75.270 3.755 ;
        RECT 75.760 3.665 76.400 3.755 ;
        RECT 74.490 3.195 74.780 3.425 ;
        RECT 75.430 3.385 75.750 3.445 ;
        RECT 77.390 3.385 77.710 3.445 ;
        RECT 78.080 3.425 78.220 4.315 ;
        RECT 78.870 4.305 79.190 4.565 ;
        RECT 79.590 4.305 79.910 4.565 ;
        RECT 80.160 4.505 80.300 4.925 ;
        RECT 80.790 4.865 81.110 5.125 ;
        RECT 81.330 5.065 81.620 5.105 ;
        RECT 81.790 5.065 82.110 5.125 ;
        RECT 81.330 4.925 82.110 5.065 ;
        RECT 81.330 4.875 81.620 4.925 ;
        RECT 81.790 4.865 82.110 4.925 ;
        RECT 82.270 4.865 82.590 5.125 ;
        RECT 82.750 4.865 83.070 5.125 ;
        RECT 83.750 4.895 84.070 5.125 ;
        RECT 97.790 5.065 98.110 5.125 ;
        RECT 83.750 4.865 85.180 4.895 ;
        RECT 83.840 4.755 85.180 4.865 ;
        RECT 81.330 4.505 81.620 4.545 ;
        RECT 80.160 4.365 81.620 4.505 ;
        RECT 81.330 4.315 81.620 4.365 ;
        RECT 83.270 4.305 83.590 4.565 ;
        RECT 83.840 4.545 83.980 4.755 ;
        RECT 83.770 4.315 84.060 4.545 ;
        RECT 84.490 4.505 84.780 4.545 ;
        RECT 84.490 4.315 84.820 4.505 ;
        RECT 82.770 4.225 83.060 4.265 ;
        RECT 83.270 4.225 83.500 4.305 ;
        RECT 82.770 4.085 83.500 4.225 ;
        RECT 82.770 4.035 83.060 4.085 ;
        RECT 78.610 3.985 78.930 4.005 ;
        RECT 78.370 3.945 78.930 3.985 ;
        RECT 79.610 3.945 79.900 3.985 ;
        RECT 78.370 3.805 79.900 3.945 ;
        RECT 78.370 3.755 78.930 3.805 ;
        RECT 79.610 3.755 79.900 3.805 ;
        RECT 80.090 3.945 80.380 3.985 ;
        RECT 80.090 3.805 81.020 3.945 ;
        RECT 80.090 3.755 80.380 3.805 ;
        RECT 78.610 3.745 78.930 3.755 ;
        RECT 75.430 3.245 77.710 3.385 ;
        RECT 75.430 3.185 75.750 3.245 ;
        RECT 77.390 3.185 77.710 3.245 ;
        RECT 77.890 3.385 78.220 3.425 ;
        RECT 78.870 3.385 79.190 3.445 ;
        RECT 79.590 3.425 79.910 3.445 ;
        RECT 77.890 3.245 79.190 3.385 ;
        RECT 77.890 3.195 78.180 3.245 ;
        RECT 78.870 3.185 79.190 3.245 ;
        RECT 79.370 3.195 79.910 3.425 ;
        RECT 79.590 3.185 79.910 3.195 ;
        RECT 80.310 3.185 80.630 3.445 ;
        RECT 80.880 3.385 81.020 3.805 ;
        RECT 81.310 3.805 81.630 4.005 ;
        RECT 84.010 3.805 84.300 3.985 ;
        RECT 81.310 3.755 84.300 3.805 ;
        RECT 81.310 3.745 84.220 3.755 ;
        RECT 81.400 3.665 84.220 3.745 ;
        RECT 84.680 3.445 84.820 4.315 ;
        RECT 85.040 4.265 85.180 4.755 ;
        RECT 86.700 4.445 87.040 4.795 ;
        RECT 93.030 4.555 93.350 4.965 ;
        RECT 97.790 4.925 98.860 5.065 ;
        RECT 96.040 4.825 97.140 4.895 ;
        RECT 97.790 4.865 98.110 4.925 ;
        RECT 95.970 4.755 97.220 4.825 ;
        RECT 95.970 4.595 96.260 4.755 ;
        RECT 96.930 4.595 97.220 4.755 ;
        RECT 84.970 4.035 85.260 4.265 ;
        RECT 86.790 3.490 86.960 4.445 ;
        RECT 88.305 3.875 88.625 3.980 ;
        RECT 88.280 3.860 88.625 3.875 ;
        RECT 88.275 3.845 88.625 3.860 ;
        RECT 88.105 3.675 88.625 3.845 ;
        RECT 88.280 3.660 88.625 3.675 ;
        RECT 88.280 3.645 88.570 3.660 ;
        RECT 89.080 3.490 89.430 3.610 ;
        RECT 90.440 3.540 90.730 3.775 ;
        RECT 90.440 3.535 90.670 3.540 ;
        RECT 81.550 3.425 81.870 3.445 ;
        RECT 81.330 3.385 81.870 3.425 ;
        RECT 80.880 3.245 81.870 3.385 ;
        RECT 81.330 3.195 81.870 3.245 ;
        RECT 81.550 3.185 81.870 3.195 ;
        RECT 82.150 3.185 82.830 3.445 ;
        RECT 83.270 3.385 83.590 3.445 ;
        RECT 83.770 3.385 84.060 3.425 ;
        RECT 83.270 3.245 84.060 3.385 ;
        RECT 84.680 3.245 85.030 3.445 ;
        RECT 86.790 3.320 89.430 3.490 ;
        RECT 88.910 3.315 89.430 3.320 ;
        RECT 89.080 3.260 89.430 3.315 ;
        RECT 83.270 3.185 83.590 3.245 ;
        RECT 83.770 3.195 84.060 3.245 ;
        RECT 84.710 3.185 85.030 3.245 ;
        RECT 90.070 3.220 90.300 3.235 ;
        RECT 88.650 3.120 88.940 3.145 ;
        RECT 90.040 3.120 90.335 3.220 ;
        RECT 88.650 2.950 90.335 3.120 ;
        RECT 88.650 2.915 88.940 2.950 ;
        RECT 70.090 2.175 70.380 2.405 ;
        RECT 71.880 2.175 72.175 2.435 ;
        RECT 88.710 2.405 88.880 2.915 ;
        RECT 90.040 2.900 90.335 2.950 ;
        RECT 90.070 2.885 90.300 2.900 ;
        RECT 90.500 2.435 90.670 3.535 ;
        RECT 93.110 3.425 93.270 4.555 ;
        RECT 93.990 4.305 94.310 4.565 ;
        RECT 95.110 4.445 95.430 4.565 ;
        RECT 96.450 4.505 96.740 4.545 ;
        RECT 95.110 4.305 95.940 4.445 ;
        RECT 96.450 4.315 96.780 4.505 ;
        RECT 95.730 4.265 95.940 4.305 ;
        RECT 95.730 4.035 96.020 4.265 ;
        RECT 93.510 3.985 93.830 4.005 ;
        RECT 93.510 3.845 94.460 3.985 ;
        RECT 94.920 3.945 95.210 3.985 ;
        RECT 93.510 3.755 94.060 3.845 ;
        RECT 94.320 3.805 94.460 3.845 ;
        RECT 94.820 3.805 95.210 3.945 ;
        RECT 94.320 3.755 95.210 3.805 ;
        RECT 93.510 3.745 93.830 3.755 ;
        RECT 94.320 3.665 94.960 3.755 ;
        RECT 93.050 3.195 93.340 3.425 ;
        RECT 93.990 3.385 94.310 3.445 ;
        RECT 95.950 3.385 96.270 3.445 ;
        RECT 96.640 3.425 96.780 4.315 ;
        RECT 97.430 4.305 97.750 4.565 ;
        RECT 98.150 4.305 98.470 4.565 ;
        RECT 98.720 4.505 98.860 4.925 ;
        RECT 99.350 4.865 99.670 5.125 ;
        RECT 99.890 5.065 100.180 5.105 ;
        RECT 100.350 5.065 100.670 5.125 ;
        RECT 99.890 4.925 100.670 5.065 ;
        RECT 99.890 4.875 100.180 4.925 ;
        RECT 100.350 4.865 100.670 4.925 ;
        RECT 100.830 4.865 101.150 5.125 ;
        RECT 101.310 4.865 101.630 5.125 ;
        RECT 102.310 4.895 102.630 5.125 ;
        RECT 102.310 4.865 103.740 4.895 ;
        RECT 102.400 4.755 103.740 4.865 ;
        RECT 99.890 4.505 100.180 4.545 ;
        RECT 98.720 4.365 100.180 4.505 ;
        RECT 99.890 4.315 100.180 4.365 ;
        RECT 101.830 4.305 102.150 4.565 ;
        RECT 102.400 4.545 102.540 4.755 ;
        RECT 102.330 4.315 102.620 4.545 ;
        RECT 103.050 4.505 103.340 4.545 ;
        RECT 103.050 4.315 103.380 4.505 ;
        RECT 101.330 4.225 101.620 4.265 ;
        RECT 101.830 4.225 102.060 4.305 ;
        RECT 101.330 4.085 102.060 4.225 ;
        RECT 101.330 4.035 101.620 4.085 ;
        RECT 97.170 3.985 97.490 4.005 ;
        RECT 96.930 3.945 97.490 3.985 ;
        RECT 98.170 3.945 98.460 3.985 ;
        RECT 96.930 3.805 98.460 3.945 ;
        RECT 96.930 3.755 97.490 3.805 ;
        RECT 98.170 3.755 98.460 3.805 ;
        RECT 98.650 3.945 98.940 3.985 ;
        RECT 98.650 3.805 99.580 3.945 ;
        RECT 98.650 3.755 98.940 3.805 ;
        RECT 97.170 3.745 97.490 3.755 ;
        RECT 93.990 3.245 96.270 3.385 ;
        RECT 93.990 3.185 94.310 3.245 ;
        RECT 95.950 3.185 96.270 3.245 ;
        RECT 96.450 3.385 96.780 3.425 ;
        RECT 97.430 3.385 97.750 3.445 ;
        RECT 98.150 3.425 98.470 3.445 ;
        RECT 96.450 3.245 97.750 3.385 ;
        RECT 96.450 3.195 96.740 3.245 ;
        RECT 97.430 3.185 97.750 3.245 ;
        RECT 97.930 3.195 98.470 3.425 ;
        RECT 98.150 3.185 98.470 3.195 ;
        RECT 98.870 3.185 99.190 3.445 ;
        RECT 99.440 3.385 99.580 3.805 ;
        RECT 99.870 3.805 100.190 4.005 ;
        RECT 102.570 3.805 102.860 3.985 ;
        RECT 99.870 3.755 102.860 3.805 ;
        RECT 99.870 3.745 102.780 3.755 ;
        RECT 99.960 3.665 102.780 3.745 ;
        RECT 103.240 3.445 103.380 4.315 ;
        RECT 103.600 4.265 103.740 4.755 ;
        RECT 105.260 4.445 105.600 4.795 ;
        RECT 103.530 4.035 103.820 4.265 ;
        RECT 105.350 3.490 105.520 4.445 ;
        RECT 106.865 3.875 107.185 3.980 ;
        RECT 106.840 3.860 107.185 3.875 ;
        RECT 106.835 3.845 107.185 3.860 ;
        RECT 106.665 3.675 107.185 3.845 ;
        RECT 106.840 3.660 107.185 3.675 ;
        RECT 106.840 3.645 107.130 3.660 ;
        RECT 107.640 3.490 107.990 3.610 ;
        RECT 109.000 3.540 109.290 3.775 ;
        RECT 109.000 3.535 109.230 3.540 ;
        RECT 100.110 3.425 100.430 3.445 ;
        RECT 99.890 3.385 100.430 3.425 ;
        RECT 99.440 3.245 100.430 3.385 ;
        RECT 99.890 3.195 100.430 3.245 ;
        RECT 100.110 3.185 100.430 3.195 ;
        RECT 100.710 3.185 101.390 3.445 ;
        RECT 101.830 3.385 102.150 3.445 ;
        RECT 102.330 3.385 102.620 3.425 ;
        RECT 101.830 3.245 102.620 3.385 ;
        RECT 103.240 3.245 103.590 3.445 ;
        RECT 105.350 3.320 107.990 3.490 ;
        RECT 107.470 3.315 107.990 3.320 ;
        RECT 107.640 3.260 107.990 3.315 ;
        RECT 101.830 3.185 102.150 3.245 ;
        RECT 102.330 3.195 102.620 3.245 ;
        RECT 103.270 3.185 103.590 3.245 ;
        RECT 108.630 3.220 108.860 3.235 ;
        RECT 107.210 3.120 107.500 3.145 ;
        RECT 108.600 3.120 108.895 3.220 ;
        RECT 107.210 2.950 108.895 3.120 ;
        RECT 107.210 2.915 107.500 2.950 ;
        RECT 88.650 2.175 88.940 2.405 ;
        RECT 90.440 2.175 90.735 2.435 ;
        RECT 107.270 2.405 107.440 2.915 ;
        RECT 108.600 2.900 108.895 2.950 ;
        RECT 108.630 2.885 108.860 2.900 ;
        RECT 109.060 2.435 109.230 3.535 ;
        RECT 107.210 2.175 107.500 2.405 ;
        RECT 109.000 2.175 109.295 2.435 ;
      LAYER met2 ;
        RECT 16.225 10.690 110.225 10.860 ;
        RECT 16.225 8.895 16.395 10.690 ;
        RECT 110.055 9.915 110.225 10.690 ;
        RECT 16.540 9.520 16.830 9.640 ;
        RECT 16.540 9.515 16.860 9.520 ;
        RECT 16.540 9.345 17.730 9.515 ;
        RECT 27.315 9.345 27.690 9.715 ;
        RECT 45.875 9.345 46.250 9.715 ;
        RECT 64.435 9.345 64.810 9.715 ;
        RECT 82.995 9.345 83.370 9.715 ;
        RECT 101.555 9.345 101.930 9.715 ;
        RECT 110.025 9.565 110.375 9.915 ;
        RECT 16.540 9.290 16.830 9.345 ;
        RECT 17.560 9.145 17.730 9.345 ;
        RECT 27.990 9.145 28.340 9.245 ;
        RECT 33.425 9.205 33.750 9.270 ;
        RECT 17.560 8.975 28.340 9.145 ;
        RECT 27.990 8.895 28.340 8.975 ;
        RECT 32.310 9.035 33.750 9.205 ;
        RECT 16.165 8.545 16.455 8.895 ;
        RECT 25.190 5.430 31.280 5.620 ;
        RECT 25.190 5.180 25.360 5.430 ;
        RECT 18.810 4.805 19.090 5.180 ;
        RECT 23.580 4.835 23.840 5.155 ;
        RECT 18.820 4.555 19.080 4.805 ;
        RECT 21.250 4.595 21.530 4.620 ;
        RECT 19.780 4.275 20.040 4.595 ;
        RECT 20.900 4.505 21.530 4.595 ;
        RECT 23.220 4.505 23.480 4.595 ;
        RECT 20.900 4.365 23.480 4.505 ;
        RECT 20.900 4.275 21.530 4.365 ;
        RECT 23.220 4.275 23.480 4.365 ;
        RECT 19.290 3.685 19.570 4.060 ;
        RECT 19.840 3.475 19.980 4.275 ;
        RECT 21.250 4.245 21.530 4.275 ;
        RECT 22.690 4.035 22.970 4.060 ;
        RECT 22.690 3.715 23.220 4.035 ;
        RECT 22.690 3.685 22.970 3.715 ;
        RECT 19.780 3.155 20.040 3.475 ;
        RECT 21.740 3.385 22.000 3.475 ;
        RECT 23.220 3.385 23.480 3.475 ;
        RECT 23.640 3.385 23.780 4.835 ;
        RECT 25.130 4.805 25.410 5.180 ;
        RECT 26.140 4.835 26.400 5.155 ;
        RECT 26.620 4.835 26.880 5.155 ;
        RECT 23.930 4.245 24.210 4.620 ;
        RECT 25.200 4.615 25.340 4.805 ;
        RECT 25.010 4.505 25.340 4.615 ;
        RECT 24.720 4.365 25.340 4.505 ;
        RECT 24.000 3.475 24.140 4.245 ;
        RECT 24.720 3.475 24.860 4.365 ;
        RECT 25.010 4.245 25.290 4.365 ;
        RECT 25.660 3.945 25.920 4.035 ;
        RECT 25.080 3.805 25.920 3.945 ;
        RECT 21.740 3.245 22.780 3.385 ;
        RECT 21.740 3.155 22.000 3.245 ;
        RECT 22.640 3.005 22.780 3.245 ;
        RECT 23.220 3.245 23.780 3.385 ;
        RECT 23.220 3.155 23.480 3.245 ;
        RECT 23.940 3.155 24.200 3.475 ;
        RECT 24.660 3.155 24.920 3.475 ;
        RECT 25.080 3.005 25.220 3.805 ;
        RECT 25.660 3.715 25.920 3.805 ;
        RECT 26.200 3.475 26.340 4.835 ;
        RECT 26.620 4.785 26.820 4.835 ;
        RECT 27.090 4.805 27.370 5.180 ;
        RECT 28.090 4.805 28.370 5.180 ;
        RECT 31.090 4.795 31.280 5.430 ;
        RECT 26.560 4.615 26.820 4.785 ;
        RECT 26.560 4.245 27.060 4.615 ;
        RECT 27.620 4.275 27.880 4.595 ;
        RECT 31.020 4.445 31.360 4.795 ;
        RECT 31.110 4.440 31.280 4.445 ;
        RECT 26.560 3.475 26.700 4.245 ;
        RECT 27.680 3.475 27.820 4.275 ;
        RECT 32.310 3.860 32.470 9.035 ;
        RECT 33.425 8.945 33.750 9.035 ;
        RECT 35.805 9.175 36.155 9.295 ;
        RECT 46.550 9.175 46.900 9.250 ;
        RECT 51.985 9.205 52.310 9.270 ;
        RECT 35.805 8.975 46.900 9.175 ;
        RECT 35.805 8.945 36.155 8.975 ;
        RECT 46.550 8.900 46.900 8.975 ;
        RECT 50.870 9.035 52.310 9.205 ;
        RECT 32.625 8.510 32.945 8.835 ;
        RECT 32.655 8.335 32.825 8.510 ;
        RECT 32.655 8.160 32.830 8.335 ;
        RECT 32.655 7.985 33.630 8.160 ;
        RECT 32.625 3.860 32.945 3.980 ;
        RECT 32.310 3.690 32.945 3.860 ;
        RECT 32.625 3.660 32.945 3.690 ;
        RECT 33.455 3.610 33.630 7.985 ;
        RECT 43.750 5.430 49.840 5.620 ;
        RECT 43.750 5.180 43.920 5.430 ;
        RECT 37.370 4.805 37.650 5.180 ;
        RECT 42.140 4.835 42.400 5.155 ;
        RECT 37.380 4.555 37.640 4.805 ;
        RECT 39.810 4.595 40.090 4.620 ;
        RECT 38.340 4.275 38.600 4.595 ;
        RECT 39.460 4.505 40.090 4.595 ;
        RECT 41.780 4.505 42.040 4.595 ;
        RECT 39.460 4.365 42.040 4.505 ;
        RECT 39.460 4.275 40.090 4.365 ;
        RECT 41.780 4.275 42.040 4.365 ;
        RECT 37.850 3.685 38.130 4.060 ;
        RECT 25.900 3.245 26.340 3.475 ;
        RECT 25.900 3.155 26.160 3.245 ;
        RECT 26.500 3.155 26.760 3.475 ;
        RECT 27.620 3.155 27.880 3.475 ;
        RECT 29.050 3.125 29.330 3.500 ;
        RECT 33.400 3.260 33.750 3.610 ;
        RECT 38.400 3.475 38.540 4.275 ;
        RECT 39.810 4.245 40.090 4.275 ;
        RECT 41.250 4.035 41.530 4.060 ;
        RECT 41.250 3.715 41.780 4.035 ;
        RECT 41.250 3.685 41.530 3.715 ;
        RECT 38.340 3.155 38.600 3.475 ;
        RECT 40.300 3.385 40.560 3.475 ;
        RECT 41.780 3.385 42.040 3.475 ;
        RECT 42.200 3.385 42.340 4.835 ;
        RECT 43.690 4.805 43.970 5.180 ;
        RECT 44.700 4.835 44.960 5.155 ;
        RECT 45.180 4.835 45.440 5.155 ;
        RECT 42.490 4.245 42.770 4.620 ;
        RECT 43.760 4.615 43.900 4.805 ;
        RECT 43.570 4.505 43.900 4.615 ;
        RECT 43.280 4.365 43.900 4.505 ;
        RECT 42.560 3.475 42.700 4.245 ;
        RECT 43.280 3.475 43.420 4.365 ;
        RECT 43.570 4.245 43.850 4.365 ;
        RECT 44.220 3.945 44.480 4.035 ;
        RECT 43.640 3.805 44.480 3.945 ;
        RECT 40.300 3.245 41.340 3.385 ;
        RECT 40.300 3.155 40.560 3.245 ;
        RECT 22.640 2.865 25.220 3.005 ;
        RECT 41.200 3.005 41.340 3.245 ;
        RECT 41.780 3.245 42.340 3.385 ;
        RECT 41.780 3.155 42.040 3.245 ;
        RECT 42.500 3.155 42.760 3.475 ;
        RECT 43.220 3.155 43.480 3.475 ;
        RECT 43.640 3.005 43.780 3.805 ;
        RECT 44.220 3.715 44.480 3.805 ;
        RECT 44.760 3.475 44.900 4.835 ;
        RECT 45.180 4.785 45.380 4.835 ;
        RECT 45.650 4.805 45.930 5.180 ;
        RECT 46.650 4.805 46.930 5.180 ;
        RECT 49.650 4.795 49.840 5.430 ;
        RECT 45.120 4.615 45.380 4.785 ;
        RECT 45.120 4.245 45.620 4.615 ;
        RECT 46.180 4.275 46.440 4.595 ;
        RECT 49.580 4.445 49.920 4.795 ;
        RECT 49.670 4.440 49.840 4.445 ;
        RECT 45.120 3.475 45.260 4.245 ;
        RECT 46.240 3.475 46.380 4.275 ;
        RECT 50.870 3.860 51.030 9.035 ;
        RECT 51.985 8.945 52.310 9.035 ;
        RECT 54.365 9.180 54.715 9.300 ;
        RECT 65.105 9.180 65.455 9.255 ;
        RECT 70.545 9.205 70.870 9.270 ;
        RECT 54.365 8.980 65.455 9.180 ;
        RECT 54.365 8.950 54.715 8.980 ;
        RECT 65.105 8.905 65.455 8.980 ;
        RECT 69.430 9.035 70.870 9.205 ;
        RECT 51.185 8.510 51.505 8.835 ;
        RECT 51.215 8.335 51.385 8.510 ;
        RECT 51.215 8.160 51.390 8.335 ;
        RECT 51.215 7.985 52.190 8.160 ;
        RECT 51.185 3.860 51.505 3.980 ;
        RECT 50.870 3.690 51.505 3.860 ;
        RECT 51.185 3.660 51.505 3.690 ;
        RECT 52.015 3.610 52.190 7.985 ;
        RECT 62.310 5.430 68.400 5.620 ;
        RECT 62.310 5.180 62.480 5.430 ;
        RECT 55.930 4.805 56.210 5.180 ;
        RECT 60.700 4.835 60.960 5.155 ;
        RECT 55.940 4.555 56.200 4.805 ;
        RECT 58.370 4.595 58.650 4.620 ;
        RECT 56.900 4.275 57.160 4.595 ;
        RECT 58.020 4.505 58.650 4.595 ;
        RECT 60.340 4.505 60.600 4.595 ;
        RECT 58.020 4.365 60.600 4.505 ;
        RECT 58.020 4.275 58.650 4.365 ;
        RECT 60.340 4.275 60.600 4.365 ;
        RECT 56.410 3.685 56.690 4.060 ;
        RECT 44.460 3.245 44.900 3.475 ;
        RECT 44.460 3.155 44.720 3.245 ;
        RECT 45.060 3.155 45.320 3.475 ;
        RECT 46.180 3.155 46.440 3.475 ;
        RECT 47.610 3.125 47.890 3.500 ;
        RECT 51.960 3.260 52.310 3.610 ;
        RECT 56.960 3.475 57.100 4.275 ;
        RECT 58.370 4.245 58.650 4.275 ;
        RECT 59.810 4.035 60.090 4.060 ;
        RECT 59.810 3.715 60.340 4.035 ;
        RECT 59.810 3.685 60.090 3.715 ;
        RECT 56.900 3.155 57.160 3.475 ;
        RECT 58.860 3.385 59.120 3.475 ;
        RECT 60.340 3.385 60.600 3.475 ;
        RECT 60.760 3.385 60.900 4.835 ;
        RECT 62.250 4.805 62.530 5.180 ;
        RECT 63.260 4.835 63.520 5.155 ;
        RECT 63.740 4.835 64.000 5.155 ;
        RECT 61.050 4.245 61.330 4.620 ;
        RECT 62.320 4.615 62.460 4.805 ;
        RECT 62.130 4.505 62.460 4.615 ;
        RECT 61.840 4.365 62.460 4.505 ;
        RECT 61.120 3.475 61.260 4.245 ;
        RECT 61.840 3.475 61.980 4.365 ;
        RECT 62.130 4.245 62.410 4.365 ;
        RECT 62.780 3.945 63.040 4.035 ;
        RECT 62.200 3.805 63.040 3.945 ;
        RECT 58.860 3.245 59.900 3.385 ;
        RECT 58.860 3.155 59.120 3.245 ;
        RECT 41.200 2.865 43.780 3.005 ;
        RECT 59.760 3.005 59.900 3.245 ;
        RECT 60.340 3.245 60.900 3.385 ;
        RECT 60.340 3.155 60.600 3.245 ;
        RECT 61.060 3.155 61.320 3.475 ;
        RECT 61.780 3.155 62.040 3.475 ;
        RECT 62.200 3.005 62.340 3.805 ;
        RECT 62.780 3.715 63.040 3.805 ;
        RECT 63.320 3.475 63.460 4.835 ;
        RECT 63.740 4.785 63.940 4.835 ;
        RECT 64.210 4.805 64.490 5.180 ;
        RECT 65.210 4.805 65.490 5.180 ;
        RECT 68.210 4.795 68.400 5.430 ;
        RECT 63.680 4.615 63.940 4.785 ;
        RECT 63.680 4.245 64.180 4.615 ;
        RECT 64.740 4.275 65.000 4.595 ;
        RECT 68.140 4.445 68.480 4.795 ;
        RECT 68.230 4.440 68.400 4.445 ;
        RECT 63.680 3.475 63.820 4.245 ;
        RECT 64.800 3.475 64.940 4.275 ;
        RECT 69.430 3.860 69.590 9.035 ;
        RECT 70.545 8.945 70.870 9.035 ;
        RECT 72.880 9.175 73.230 9.295 ;
        RECT 83.665 9.175 84.015 9.250 ;
        RECT 89.105 9.205 89.430 9.270 ;
        RECT 72.880 8.975 84.015 9.175 ;
        RECT 72.880 8.945 73.230 8.975 ;
        RECT 83.665 8.900 84.015 8.975 ;
        RECT 87.990 9.035 89.430 9.205 ;
        RECT 69.745 8.510 70.065 8.835 ;
        RECT 69.775 8.335 69.945 8.510 ;
        RECT 69.775 8.160 69.950 8.335 ;
        RECT 69.775 7.985 70.750 8.160 ;
        RECT 69.745 3.860 70.065 3.980 ;
        RECT 69.430 3.690 70.065 3.860 ;
        RECT 69.745 3.660 70.065 3.690 ;
        RECT 70.575 3.610 70.750 7.985 ;
        RECT 80.870 5.430 86.960 5.620 ;
        RECT 80.870 5.180 81.040 5.430 ;
        RECT 74.490 4.805 74.770 5.180 ;
        RECT 79.260 4.835 79.520 5.155 ;
        RECT 74.500 4.555 74.760 4.805 ;
        RECT 76.930 4.595 77.210 4.620 ;
        RECT 75.460 4.275 75.720 4.595 ;
        RECT 76.580 4.505 77.210 4.595 ;
        RECT 78.900 4.505 79.160 4.595 ;
        RECT 76.580 4.365 79.160 4.505 ;
        RECT 76.580 4.275 77.210 4.365 ;
        RECT 78.900 4.275 79.160 4.365 ;
        RECT 74.970 3.685 75.250 4.060 ;
        RECT 63.020 3.245 63.460 3.475 ;
        RECT 63.020 3.155 63.280 3.245 ;
        RECT 63.620 3.155 63.880 3.475 ;
        RECT 64.740 3.155 65.000 3.475 ;
        RECT 66.170 3.125 66.450 3.500 ;
        RECT 70.520 3.260 70.870 3.610 ;
        RECT 75.520 3.475 75.660 4.275 ;
        RECT 76.930 4.245 77.210 4.275 ;
        RECT 78.370 4.035 78.650 4.060 ;
        RECT 78.370 3.715 78.900 4.035 ;
        RECT 78.370 3.685 78.650 3.715 ;
        RECT 75.460 3.155 75.720 3.475 ;
        RECT 77.420 3.385 77.680 3.475 ;
        RECT 78.900 3.385 79.160 3.475 ;
        RECT 79.320 3.385 79.460 4.835 ;
        RECT 80.810 4.805 81.090 5.180 ;
        RECT 81.820 4.835 82.080 5.155 ;
        RECT 82.300 4.835 82.560 5.155 ;
        RECT 79.610 4.245 79.890 4.620 ;
        RECT 80.880 4.615 81.020 4.805 ;
        RECT 80.690 4.505 81.020 4.615 ;
        RECT 80.400 4.365 81.020 4.505 ;
        RECT 79.680 3.475 79.820 4.245 ;
        RECT 80.400 3.475 80.540 4.365 ;
        RECT 80.690 4.245 80.970 4.365 ;
        RECT 81.340 3.945 81.600 4.035 ;
        RECT 80.760 3.805 81.600 3.945 ;
        RECT 77.420 3.245 78.460 3.385 ;
        RECT 77.420 3.155 77.680 3.245 ;
        RECT 59.760 2.865 62.340 3.005 ;
        RECT 78.320 3.005 78.460 3.245 ;
        RECT 78.900 3.245 79.460 3.385 ;
        RECT 78.900 3.155 79.160 3.245 ;
        RECT 79.620 3.155 79.880 3.475 ;
        RECT 80.340 3.155 80.600 3.475 ;
        RECT 80.760 3.005 80.900 3.805 ;
        RECT 81.340 3.715 81.600 3.805 ;
        RECT 81.880 3.475 82.020 4.835 ;
        RECT 82.300 4.785 82.500 4.835 ;
        RECT 82.770 4.805 83.050 5.180 ;
        RECT 83.770 4.805 84.050 5.180 ;
        RECT 86.770 4.795 86.960 5.430 ;
        RECT 82.240 4.615 82.500 4.785 ;
        RECT 82.240 4.245 82.740 4.615 ;
        RECT 83.300 4.275 83.560 4.595 ;
        RECT 86.700 4.445 87.040 4.795 ;
        RECT 86.790 4.440 86.960 4.445 ;
        RECT 82.240 3.475 82.380 4.245 ;
        RECT 83.360 3.475 83.500 4.275 ;
        RECT 87.990 3.860 88.150 9.035 ;
        RECT 89.105 8.945 89.430 9.035 ;
        RECT 91.440 9.175 91.790 9.295 ;
        RECT 102.225 9.175 102.575 9.250 ;
        RECT 107.665 9.205 107.990 9.270 ;
        RECT 91.440 8.975 102.575 9.175 ;
        RECT 91.440 8.945 91.790 8.975 ;
        RECT 102.225 8.900 102.575 8.975 ;
        RECT 106.550 9.035 107.990 9.205 ;
        RECT 88.305 8.510 88.625 8.835 ;
        RECT 88.335 8.335 88.505 8.510 ;
        RECT 88.335 8.160 88.510 8.335 ;
        RECT 88.335 7.985 89.310 8.160 ;
        RECT 88.305 3.860 88.625 3.980 ;
        RECT 87.990 3.690 88.625 3.860 ;
        RECT 88.305 3.660 88.625 3.690 ;
        RECT 89.135 3.610 89.310 7.985 ;
        RECT 99.430 5.430 105.520 5.620 ;
        RECT 99.430 5.180 99.600 5.430 ;
        RECT 93.050 4.805 93.330 5.180 ;
        RECT 97.820 4.835 98.080 5.155 ;
        RECT 93.060 4.555 93.320 4.805 ;
        RECT 95.490 4.595 95.770 4.620 ;
        RECT 94.020 4.275 94.280 4.595 ;
        RECT 95.140 4.505 95.770 4.595 ;
        RECT 97.460 4.505 97.720 4.595 ;
        RECT 95.140 4.365 97.720 4.505 ;
        RECT 95.140 4.275 95.770 4.365 ;
        RECT 97.460 4.275 97.720 4.365 ;
        RECT 93.530 3.685 93.810 4.060 ;
        RECT 81.580 3.245 82.020 3.475 ;
        RECT 81.580 3.155 81.840 3.245 ;
        RECT 82.180 3.155 82.440 3.475 ;
        RECT 83.300 3.155 83.560 3.475 ;
        RECT 84.730 3.125 85.010 3.500 ;
        RECT 89.080 3.260 89.430 3.610 ;
        RECT 94.080 3.475 94.220 4.275 ;
        RECT 95.490 4.245 95.770 4.275 ;
        RECT 96.930 4.035 97.210 4.060 ;
        RECT 96.930 3.715 97.460 4.035 ;
        RECT 96.930 3.685 97.210 3.715 ;
        RECT 94.020 3.155 94.280 3.475 ;
        RECT 95.980 3.385 96.240 3.475 ;
        RECT 97.460 3.385 97.720 3.475 ;
        RECT 97.880 3.385 98.020 4.835 ;
        RECT 99.370 4.805 99.650 5.180 ;
        RECT 100.380 4.835 100.640 5.155 ;
        RECT 100.860 4.835 101.120 5.155 ;
        RECT 98.170 4.245 98.450 4.620 ;
        RECT 99.440 4.615 99.580 4.805 ;
        RECT 99.250 4.505 99.580 4.615 ;
        RECT 98.960 4.365 99.580 4.505 ;
        RECT 98.240 3.475 98.380 4.245 ;
        RECT 98.960 3.475 99.100 4.365 ;
        RECT 99.250 4.245 99.530 4.365 ;
        RECT 99.900 3.945 100.160 4.035 ;
        RECT 99.320 3.805 100.160 3.945 ;
        RECT 95.980 3.245 97.020 3.385 ;
        RECT 95.980 3.155 96.240 3.245 ;
        RECT 78.320 2.865 80.900 3.005 ;
        RECT 96.880 3.005 97.020 3.245 ;
        RECT 97.460 3.245 98.020 3.385 ;
        RECT 97.460 3.155 97.720 3.245 ;
        RECT 98.180 3.155 98.440 3.475 ;
        RECT 98.900 3.155 99.160 3.475 ;
        RECT 99.320 3.005 99.460 3.805 ;
        RECT 99.900 3.715 100.160 3.805 ;
        RECT 100.440 3.475 100.580 4.835 ;
        RECT 100.860 4.785 101.060 4.835 ;
        RECT 101.330 4.805 101.610 5.180 ;
        RECT 102.330 4.805 102.610 5.180 ;
        RECT 105.330 4.795 105.520 5.430 ;
        RECT 100.800 4.615 101.060 4.785 ;
        RECT 100.800 4.245 101.300 4.615 ;
        RECT 101.860 4.275 102.120 4.595 ;
        RECT 105.260 4.445 105.600 4.795 ;
        RECT 105.350 4.440 105.520 4.445 ;
        RECT 100.800 3.475 100.940 4.245 ;
        RECT 101.920 3.475 102.060 4.275 ;
        RECT 106.550 3.860 106.710 9.035 ;
        RECT 107.665 8.945 107.990 9.035 ;
        RECT 106.865 8.510 107.185 8.835 ;
        RECT 106.895 8.335 107.065 8.510 ;
        RECT 106.895 8.160 107.070 8.335 ;
        RECT 106.895 7.985 107.870 8.160 ;
        RECT 106.865 3.860 107.185 3.980 ;
        RECT 106.550 3.690 107.185 3.860 ;
        RECT 106.865 3.660 107.185 3.690 ;
        RECT 107.695 3.610 107.870 7.985 ;
        RECT 100.140 3.245 100.580 3.475 ;
        RECT 100.140 3.155 100.400 3.245 ;
        RECT 100.740 3.155 101.000 3.475 ;
        RECT 101.860 3.155 102.120 3.475 ;
        RECT 103.290 3.125 103.570 3.500 ;
        RECT 107.640 3.260 107.990 3.610 ;
        RECT 96.880 2.865 99.460 3.005 ;
      LAYER met3 ;
        RECT 27.315 9.685 27.690 9.715 ;
        RECT 45.875 9.685 46.250 9.715 ;
        RECT 64.435 9.685 64.810 9.715 ;
        RECT 82.995 9.685 83.370 9.715 ;
        RECT 101.555 9.685 101.930 9.715 ;
        RECT 27.315 9.385 28.320 9.685 ;
        RECT 27.315 9.345 27.690 9.385 ;
        RECT 28.020 6.995 28.320 9.385 ;
        RECT 45.875 9.385 46.880 9.685 ;
        RECT 45.875 9.345 46.250 9.385 ;
        RECT 46.580 6.995 46.880 9.385 ;
        RECT 64.435 9.385 65.440 9.685 ;
        RECT 64.435 9.345 64.810 9.385 ;
        RECT 65.140 6.995 65.440 9.385 ;
        RECT 82.995 9.385 84.000 9.685 ;
        RECT 82.995 9.345 83.370 9.385 ;
        RECT 83.700 6.995 84.000 9.385 ;
        RECT 101.555 9.385 102.560 9.685 ;
        RECT 101.555 9.345 101.930 9.385 ;
        RECT 102.260 6.995 102.560 9.385 ;
        RECT 18.185 6.695 28.320 6.995 ;
        RECT 36.745 6.695 46.880 6.995 ;
        RECT 55.305 6.695 65.440 6.995 ;
        RECT 73.865 6.695 84.000 6.995 ;
        RECT 92.425 6.695 102.560 6.995 ;
        RECT 18.185 4.015 18.485 6.695 ;
        RECT 18.785 5.155 19.110 5.160 ;
        RECT 18.785 4.825 19.520 5.155 ;
        RECT 18.785 4.820 19.110 4.825 ;
        RECT 21.260 4.600 21.560 6.695 ;
        RECT 21.225 4.595 21.560 4.600 ;
        RECT 21.225 4.265 21.960 4.595 ;
        RECT 21.225 4.260 21.555 4.265 ;
        RECT 22.695 4.040 22.995 6.695 ;
        RECT 25.105 5.155 25.435 5.160 ;
        RECT 27.070 5.155 27.395 5.160 ;
        RECT 28.075 5.155 28.395 5.160 ;
        RECT 25.105 4.825 25.840 5.155 ;
        RECT 26.810 4.825 27.540 5.155 ;
        RECT 27.840 4.825 28.400 5.155 ;
        RECT 25.105 4.820 25.435 4.825 ;
        RECT 27.070 4.820 27.395 4.825 ;
        RECT 23.905 4.595 24.225 4.600 ;
        RECT 23.905 4.260 24.460 4.595 ;
        RECT 19.120 4.035 19.640 4.040 ;
        RECT 22.665 4.035 22.995 4.040 ;
        RECT 19.120 4.015 19.850 4.035 ;
        RECT 18.185 3.715 19.850 4.015 ;
        RECT 19.120 3.705 19.850 3.715 ;
        RECT 22.665 3.705 23.400 4.035 ;
        RECT 22.665 3.700 22.990 3.705 ;
        RECT 24.160 3.465 24.460 4.260 ;
        RECT 27.840 3.465 28.140 4.825 ;
        RECT 36.745 4.015 37.045 6.695 ;
        RECT 37.345 5.155 37.670 5.160 ;
        RECT 37.345 4.825 38.080 5.155 ;
        RECT 37.345 4.820 37.670 4.825 ;
        RECT 39.820 4.600 40.120 6.695 ;
        RECT 39.785 4.595 40.120 4.600 ;
        RECT 39.785 4.265 40.520 4.595 ;
        RECT 39.785 4.260 40.115 4.265 ;
        RECT 41.255 4.040 41.555 6.695 ;
        RECT 43.665 5.155 43.995 5.160 ;
        RECT 45.630 5.155 45.955 5.160 ;
        RECT 46.635 5.155 46.955 5.160 ;
        RECT 43.665 4.825 44.400 5.155 ;
        RECT 45.370 4.825 46.100 5.155 ;
        RECT 46.400 4.825 46.960 5.155 ;
        RECT 43.665 4.820 43.995 4.825 ;
        RECT 45.630 4.820 45.955 4.825 ;
        RECT 42.465 4.595 42.785 4.600 ;
        RECT 42.465 4.260 43.020 4.595 ;
        RECT 37.680 4.035 38.200 4.040 ;
        RECT 41.225 4.035 41.555 4.040 ;
        RECT 37.680 4.015 38.410 4.035 ;
        RECT 36.745 3.715 38.410 4.015 ;
        RECT 37.680 3.705 38.410 3.715 ;
        RECT 41.225 3.705 41.960 4.035 ;
        RECT 41.225 3.700 41.550 3.705 ;
        RECT 24.160 3.165 28.140 3.465 ;
        RECT 29.025 3.475 29.350 3.480 ;
        RECT 29.025 3.145 29.760 3.475 ;
        RECT 42.720 3.465 43.020 4.260 ;
        RECT 46.400 3.465 46.700 4.825 ;
        RECT 55.305 4.015 55.605 6.695 ;
        RECT 55.905 5.155 56.230 5.160 ;
        RECT 55.905 4.825 56.640 5.155 ;
        RECT 55.905 4.820 56.230 4.825 ;
        RECT 58.380 4.600 58.680 6.695 ;
        RECT 58.345 4.595 58.680 4.600 ;
        RECT 58.345 4.265 59.080 4.595 ;
        RECT 58.345 4.260 58.675 4.265 ;
        RECT 59.815 4.040 60.115 6.695 ;
        RECT 62.225 5.155 62.555 5.160 ;
        RECT 64.190 5.155 64.515 5.160 ;
        RECT 65.195 5.155 65.515 5.160 ;
        RECT 62.225 4.825 62.960 5.155 ;
        RECT 63.930 4.825 64.660 5.155 ;
        RECT 64.960 4.825 65.520 5.155 ;
        RECT 62.225 4.820 62.555 4.825 ;
        RECT 64.190 4.820 64.515 4.825 ;
        RECT 61.025 4.595 61.345 4.600 ;
        RECT 61.025 4.260 61.580 4.595 ;
        RECT 56.240 4.035 56.760 4.040 ;
        RECT 59.785 4.035 60.115 4.040 ;
        RECT 56.240 4.015 56.970 4.035 ;
        RECT 55.305 3.715 56.970 4.015 ;
        RECT 56.240 3.705 56.970 3.715 ;
        RECT 59.785 3.705 60.520 4.035 ;
        RECT 59.785 3.700 60.110 3.705 ;
        RECT 42.720 3.165 46.700 3.465 ;
        RECT 47.585 3.475 47.910 3.480 ;
        RECT 47.585 3.145 48.320 3.475 ;
        RECT 61.280 3.465 61.580 4.260 ;
        RECT 64.960 3.465 65.260 4.825 ;
        RECT 73.865 4.015 74.165 6.695 ;
        RECT 74.465 5.155 74.790 5.160 ;
        RECT 74.465 4.825 75.200 5.155 ;
        RECT 74.465 4.820 74.790 4.825 ;
        RECT 76.940 4.600 77.240 6.695 ;
        RECT 76.905 4.595 77.240 4.600 ;
        RECT 76.905 4.265 77.640 4.595 ;
        RECT 76.905 4.260 77.235 4.265 ;
        RECT 78.375 4.040 78.675 6.695 ;
        RECT 80.785 5.155 81.115 5.160 ;
        RECT 82.750 5.155 83.075 5.160 ;
        RECT 83.755 5.155 84.075 5.160 ;
        RECT 80.785 4.825 81.520 5.155 ;
        RECT 82.490 4.825 83.220 5.155 ;
        RECT 83.520 4.825 84.080 5.155 ;
        RECT 80.785 4.820 81.115 4.825 ;
        RECT 82.750 4.820 83.075 4.825 ;
        RECT 79.585 4.595 79.905 4.600 ;
        RECT 79.585 4.260 80.140 4.595 ;
        RECT 74.800 4.035 75.320 4.040 ;
        RECT 78.345 4.035 78.675 4.040 ;
        RECT 74.800 4.015 75.530 4.035 ;
        RECT 73.865 3.715 75.530 4.015 ;
        RECT 74.800 3.705 75.530 3.715 ;
        RECT 78.345 3.705 79.080 4.035 ;
        RECT 78.345 3.700 78.670 3.705 ;
        RECT 61.280 3.165 65.260 3.465 ;
        RECT 66.145 3.475 66.470 3.480 ;
        RECT 66.145 3.145 66.880 3.475 ;
        RECT 79.840 3.465 80.140 4.260 ;
        RECT 83.520 3.465 83.820 4.825 ;
        RECT 92.425 4.015 92.725 6.695 ;
        RECT 93.025 5.155 93.350 5.160 ;
        RECT 93.025 4.825 93.760 5.155 ;
        RECT 93.025 4.820 93.350 4.825 ;
        RECT 95.500 4.600 95.800 6.695 ;
        RECT 95.465 4.595 95.800 4.600 ;
        RECT 95.465 4.265 96.200 4.595 ;
        RECT 95.465 4.260 95.795 4.265 ;
        RECT 96.935 4.040 97.235 6.695 ;
        RECT 99.345 5.155 99.675 5.160 ;
        RECT 101.310 5.155 101.635 5.160 ;
        RECT 102.315 5.155 102.635 5.160 ;
        RECT 99.345 4.825 100.080 5.155 ;
        RECT 101.050 4.825 101.780 5.155 ;
        RECT 102.080 4.825 102.640 5.155 ;
        RECT 99.345 4.820 99.675 4.825 ;
        RECT 101.310 4.820 101.635 4.825 ;
        RECT 98.145 4.595 98.465 4.600 ;
        RECT 98.145 4.260 98.700 4.595 ;
        RECT 93.360 4.035 93.880 4.040 ;
        RECT 96.905 4.035 97.235 4.040 ;
        RECT 93.360 4.015 94.090 4.035 ;
        RECT 92.425 3.715 94.090 4.015 ;
        RECT 93.360 3.705 94.090 3.715 ;
        RECT 96.905 3.705 97.640 4.035 ;
        RECT 96.905 3.700 97.230 3.705 ;
        RECT 79.840 3.165 83.820 3.465 ;
        RECT 84.705 3.475 85.030 3.480 ;
        RECT 84.705 3.145 85.440 3.475 ;
        RECT 98.400 3.465 98.700 4.260 ;
        RECT 102.080 3.465 102.380 4.825 ;
        RECT 98.400 3.165 102.380 3.465 ;
        RECT 103.265 3.475 103.590 3.480 ;
        RECT 103.265 3.145 104.000 3.475 ;
        RECT 29.025 3.140 29.350 3.145 ;
        RECT 47.585 3.140 47.910 3.145 ;
        RECT 66.145 3.140 66.470 3.145 ;
        RECT 84.705 3.140 85.030 3.145 ;
        RECT 103.265 3.140 103.590 3.145 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r2
MACRO mux16x1_project
  CLASS BLOCK ;
  FOREIGN mux16x1_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 110.000 ;
  PIN data_in[0]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 9.685 96.565 10.015 96.935 ;
      LAYER met1 ;
        RECT 5.130 96.800 5.450 96.860 ;
        RECT 9.745 96.800 10.035 96.845 ;
        RECT 5.130 96.660 10.035 96.800 ;
        RECT 5.130 96.600 5.450 96.660 ;
        RECT 9.745 96.615 10.035 96.660 ;
      LAYER met2 ;
        RECT 5.150 104.875 5.430 105.245 ;
        RECT 5.220 96.890 5.360 104.875 ;
        RECT 5.160 96.570 5.420 96.890 ;
      LAYER met3 ;
        RECT 0.000 105.210 4.000 105.360 ;
        RECT 5.125 105.210 5.455 105.225 ;
        RECT 0.000 104.910 5.455 105.210 ;
        RECT 0.000 104.760 4.000 104.910 ;
        RECT 5.125 104.895 5.455 104.910 ;
    END
  END data_in[0]
  PIN data_in[10]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 36.725 7.335 37.095 ;
      LAYER met1 ;
        RECT 4.670 36.960 4.990 37.020 ;
        RECT 6.985 36.960 7.275 37.005 ;
        RECT 4.670 36.820 7.275 36.960 ;
        RECT 4.670 36.760 4.990 36.820 ;
        RECT 6.985 36.775 7.275 36.820 ;
      LAYER met2 ;
        RECT 4.690 36.875 4.970 37.245 ;
        RECT 4.700 36.730 4.960 36.875 ;
      LAYER met3 ;
        RECT 0.000 37.210 4.000 37.360 ;
        RECT 4.665 37.210 4.995 37.225 ;
        RECT 0.000 36.910 4.995 37.210 ;
        RECT 0.000 36.760 4.000 36.910 ;
        RECT 4.665 36.895 4.995 36.910 ;
    END
  END data_in[10]
  PIN data_in[11]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 28.185 7.335 28.555 ;
      LAYER met1 ;
        RECT 4.670 28.460 4.990 28.520 ;
        RECT 6.985 28.460 7.275 28.505 ;
        RECT 4.670 28.320 7.275 28.460 ;
        RECT 4.670 28.260 4.990 28.320 ;
        RECT 6.985 28.275 7.275 28.320 ;
      LAYER met2 ;
        RECT 4.690 30.075 4.970 30.445 ;
        RECT 4.760 28.550 4.900 30.075 ;
        RECT 4.700 28.230 4.960 28.550 ;
      LAYER met3 ;
        RECT 0.000 30.410 4.000 30.560 ;
        RECT 4.665 30.410 4.995 30.425 ;
        RECT 0.000 30.110 4.995 30.410 ;
        RECT 0.000 29.960 4.000 30.110 ;
        RECT 4.665 30.095 4.995 30.110 ;
    END
  END data_in[11]
  PIN data_in[12]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 22.745 7.335 23.115 ;
      LAYER met1 ;
        RECT 4.670 23.020 4.990 23.080 ;
        RECT 6.985 23.020 7.275 23.065 ;
        RECT 4.670 22.880 7.275 23.020 ;
        RECT 4.670 22.820 4.990 22.880 ;
        RECT 6.985 22.835 7.275 22.880 ;
      LAYER met2 ;
        RECT 4.690 23.275 4.970 23.645 ;
        RECT 4.760 23.110 4.900 23.275 ;
        RECT 4.700 22.790 4.960 23.110 ;
      LAYER met3 ;
        RECT 0.000 23.610 4.000 23.760 ;
        RECT 4.665 23.610 4.995 23.625 ;
        RECT 0.000 23.310 4.995 23.610 ;
        RECT 0.000 23.160 4.000 23.310 ;
        RECT 4.665 23.295 4.995 23.310 ;
    END
  END data_in[12]
  PIN data_in[13]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 17.305 7.335 17.675 ;
      LAYER met1 ;
        RECT 4.670 17.580 4.990 17.640 ;
        RECT 6.985 17.580 7.275 17.625 ;
        RECT 4.670 17.440 7.275 17.580 ;
        RECT 4.670 17.380 4.990 17.440 ;
        RECT 6.985 17.395 7.275 17.440 ;
      LAYER met2 ;
        RECT 4.700 17.350 4.960 17.670 ;
        RECT 4.760 16.845 4.900 17.350 ;
        RECT 4.690 16.475 4.970 16.845 ;
      LAYER met3 ;
        RECT 0.000 16.810 4.000 16.960 ;
        RECT 4.665 16.810 4.995 16.825 ;
        RECT 0.000 16.510 4.995 16.810 ;
        RECT 0.000 16.360 4.000 16.510 ;
        RECT 4.665 16.495 4.995 16.510 ;
    END
  END data_in[13]
  PIN data_in[14]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 11.865 7.335 12.235 ;
      LAYER met1 ;
        RECT 4.670 12.140 4.990 12.200 ;
        RECT 6.985 12.140 7.275 12.185 ;
        RECT 4.670 12.000 7.275 12.140 ;
        RECT 4.670 11.940 4.990 12.000 ;
        RECT 6.985 11.955 7.275 12.000 ;
      LAYER met2 ;
        RECT 4.700 11.910 4.960 12.230 ;
        RECT 4.760 10.045 4.900 11.910 ;
        RECT 4.690 9.675 4.970 10.045 ;
      LAYER met3 ;
        RECT 0.000 10.010 4.000 10.160 ;
        RECT 4.665 10.010 4.995 10.025 ;
        RECT 0.000 9.710 4.995 10.010 ;
        RECT 0.000 9.560 4.000 9.710 ;
        RECT 4.665 9.695 4.995 9.710 ;
    END
  END data_in[14]
  PIN data_in[15]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 8.385 11.865 8.715 12.235 ;
      LAYER met1 ;
        RECT 8.350 11.940 8.670 12.200 ;
      LAYER met2 ;
        RECT 8.380 11.910 8.640 12.230 ;
        RECT 8.440 3.925 8.580 11.910 ;
        RECT 8.370 3.555 8.650 3.925 ;
      LAYER met3 ;
        RECT 8.345 3.890 8.675 3.905 ;
        RECT 4.910 3.590 8.675 3.890 ;
        RECT 0.000 3.210 4.000 3.360 ;
        RECT 4.910 3.210 5.210 3.590 ;
        RECT 8.345 3.575 8.675 3.590 ;
        RECT 0.000 2.910 5.210 3.210 ;
        RECT 0.000 2.760 4.000 2.910 ;
    END
  END data_in[15]
  PIN data_in[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 11.065 96.565 11.395 96.935 ;
      LAYER met1 ;
        RECT 5.590 97.480 5.910 97.540 ;
        RECT 5.590 97.340 8.120 97.480 ;
        RECT 5.590 97.280 5.910 97.340 ;
        RECT 7.980 97.140 8.120 97.340 ;
        RECT 7.980 97.000 11.340 97.140 ;
        RECT 11.200 96.845 11.340 97.000 ;
        RECT 11.125 96.615 11.415 96.845 ;
      LAYER met2 ;
        RECT 5.610 98.075 5.890 98.445 ;
        RECT 5.680 97.570 5.820 98.075 ;
        RECT 5.620 97.250 5.880 97.570 ;
      LAYER met3 ;
        RECT 0.000 98.410 4.000 98.560 ;
        RECT 5.585 98.410 5.915 98.425 ;
        RECT 0.000 98.110 5.915 98.410 ;
        RECT 0.000 97.960 4.000 98.110 ;
        RECT 5.585 98.095 5.915 98.110 ;
    END
  END data_in[1]
  PIN data_in[2]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 93.465 7.335 93.835 ;
      LAYER met1 ;
        RECT 4.670 93.740 4.990 93.800 ;
        RECT 6.985 93.740 7.275 93.785 ;
        RECT 4.670 93.600 7.275 93.740 ;
        RECT 4.670 93.540 4.990 93.600 ;
        RECT 6.985 93.555 7.275 93.600 ;
      LAYER met2 ;
        RECT 4.700 93.510 4.960 93.830 ;
        RECT 4.760 91.645 4.900 93.510 ;
        RECT 4.690 91.275 4.970 91.645 ;
      LAYER met3 ;
        RECT 0.000 91.610 4.000 91.760 ;
        RECT 4.665 91.610 4.995 91.625 ;
        RECT 0.000 91.310 4.995 91.610 ;
        RECT 0.000 91.160 4.000 91.310 ;
        RECT 4.665 91.295 4.995 91.310 ;
    END
  END data_in[2]
  PIN data_in[3]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 85.685 7.335 86.055 ;
      LAYER met1 ;
        RECT 4.670 85.920 4.990 85.980 ;
        RECT 6.985 85.920 7.275 85.965 ;
        RECT 4.670 85.780 7.275 85.920 ;
        RECT 4.670 85.720 4.990 85.780 ;
        RECT 6.985 85.735 7.275 85.780 ;
      LAYER met2 ;
        RECT 4.700 85.690 4.960 86.010 ;
        RECT 4.760 84.845 4.900 85.690 ;
        RECT 4.690 84.475 4.970 84.845 ;
      LAYER met3 ;
        RECT 0.000 84.810 4.000 84.960 ;
        RECT 4.665 84.810 4.995 84.825 ;
        RECT 0.000 84.510 4.995 84.810 ;
        RECT 0.000 84.360 4.000 84.510 ;
        RECT 4.665 84.495 4.995 84.510 ;
    END
  END data_in[3]
  PIN data_in[4]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 77.145 7.335 77.515 ;
      LAYER met1 ;
        RECT 4.670 77.420 4.990 77.480 ;
        RECT 6.985 77.420 7.275 77.465 ;
        RECT 4.670 77.280 7.275 77.420 ;
        RECT 4.670 77.220 4.990 77.280 ;
        RECT 6.985 77.235 7.275 77.280 ;
      LAYER met2 ;
        RECT 4.690 77.675 4.970 78.045 ;
        RECT 4.760 77.510 4.900 77.675 ;
        RECT 4.700 77.190 4.960 77.510 ;
      LAYER met3 ;
        RECT 0.000 78.010 4.000 78.160 ;
        RECT 4.665 78.010 4.995 78.025 ;
        RECT 0.000 77.710 4.995 78.010 ;
        RECT 0.000 77.560 4.000 77.710 ;
        RECT 4.665 77.695 4.995 77.710 ;
    END
  END data_in[4]
  PIN data_in[5]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 71.705 7.335 72.075 ;
      LAYER met1 ;
        RECT 4.670 71.980 4.990 72.040 ;
        RECT 6.985 71.980 7.275 72.025 ;
        RECT 4.670 71.840 7.275 71.980 ;
        RECT 4.670 71.780 4.990 71.840 ;
        RECT 6.985 71.795 7.275 71.840 ;
      LAYER met2 ;
        RECT 4.700 71.750 4.960 72.070 ;
        RECT 4.760 71.245 4.900 71.750 ;
        RECT 4.690 70.875 4.970 71.245 ;
      LAYER met3 ;
        RECT 0.000 71.210 4.000 71.360 ;
        RECT 4.665 71.210 4.995 71.225 ;
        RECT 0.000 70.910 4.995 71.210 ;
        RECT 0.000 70.760 4.000 70.910 ;
        RECT 4.665 70.895 4.995 70.910 ;
    END
  END data_in[5]
  PIN data_in[6]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 66.265 7.335 66.635 ;
      LAYER met1 ;
        RECT 4.670 66.540 4.990 66.600 ;
        RECT 6.985 66.540 7.275 66.585 ;
        RECT 4.670 66.400 7.275 66.540 ;
        RECT 4.670 66.340 4.990 66.400 ;
        RECT 6.985 66.355 7.275 66.400 ;
      LAYER met2 ;
        RECT 4.700 66.310 4.960 66.630 ;
        RECT 4.760 64.445 4.900 66.310 ;
        RECT 4.690 64.075 4.970 64.445 ;
      LAYER met3 ;
        RECT 0.000 64.410 4.000 64.560 ;
        RECT 4.665 64.410 4.995 64.425 ;
        RECT 0.000 64.110 4.995 64.410 ;
        RECT 0.000 63.960 4.000 64.110 ;
        RECT 4.665 64.095 4.995 64.110 ;
    END
  END data_in[6]
  PIN data_in[7]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 58.485 7.335 58.855 ;
      LAYER met1 ;
        RECT 4.670 58.720 4.990 58.780 ;
        RECT 6.985 58.720 7.275 58.765 ;
        RECT 4.670 58.580 7.275 58.720 ;
        RECT 4.670 58.520 4.990 58.580 ;
        RECT 6.985 58.535 7.275 58.580 ;
      LAYER met2 ;
        RECT 4.700 58.490 4.960 58.810 ;
        RECT 4.760 57.645 4.900 58.490 ;
        RECT 4.690 57.275 4.970 57.645 ;
      LAYER met3 ;
        RECT 0.000 57.610 4.000 57.760 ;
        RECT 4.665 57.610 4.995 57.625 ;
        RECT 0.000 57.310 4.995 57.610 ;
        RECT 0.000 57.160 4.000 57.310 ;
        RECT 4.665 57.295 4.995 57.310 ;
    END
  END data_in[7]
  PIN data_in[8]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 53.045 7.335 53.415 ;
      LAYER met1 ;
        RECT 4.670 53.280 4.990 53.340 ;
        RECT 6.985 53.280 7.275 53.325 ;
        RECT 4.670 53.140 7.275 53.280 ;
        RECT 4.670 53.080 4.990 53.140 ;
        RECT 6.985 53.095 7.275 53.140 ;
      LAYER met2 ;
        RECT 4.700 53.050 4.960 53.370 ;
        RECT 4.760 50.845 4.900 53.050 ;
        RECT 4.690 50.475 4.970 50.845 ;
      LAYER met3 ;
        RECT 0.000 50.810 4.000 50.960 ;
        RECT 4.665 50.810 4.995 50.825 ;
        RECT 0.000 50.510 4.995 50.810 ;
        RECT 0.000 50.360 4.000 50.510 ;
        RECT 4.665 50.495 4.995 50.510 ;
    END
  END data_in[8]
  PIN data_in[9]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 7.005 44.505 7.335 44.875 ;
      LAYER met1 ;
        RECT 4.670 44.780 4.990 44.840 ;
        RECT 6.985 44.780 7.275 44.825 ;
        RECT 4.670 44.640 7.275 44.780 ;
        RECT 4.670 44.580 4.990 44.640 ;
        RECT 6.985 44.595 7.275 44.640 ;
      LAYER met2 ;
        RECT 4.700 44.550 4.960 44.870 ;
        RECT 4.760 44.045 4.900 44.550 ;
        RECT 4.690 43.675 4.970 44.045 ;
      LAYER met3 ;
        RECT 0.000 44.010 4.000 44.160 ;
        RECT 4.665 44.010 4.995 44.025 ;
        RECT 0.000 43.710 4.995 44.010 ;
        RECT 0.000 43.560 4.000 43.710 ;
        RECT 4.665 43.695 4.995 43.710 ;
    END
  END data_in[9]
  PIN select[0]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 7.325 96.595 7.685 97.175 ;
      LAYER met1 ;
        RECT 6.970 97.140 7.290 97.200 ;
        RECT 7.445 97.140 7.735 97.185 ;
        RECT 6.970 97.000 7.735 97.140 ;
        RECT 6.970 96.940 7.290 97.000 ;
        RECT 7.445 96.955 7.735 97.000 ;
      LAYER met2 ;
        RECT 6.070 106.490 6.350 110.000 ;
        RECT 6.070 106.350 7.200 106.490 ;
        RECT 6.070 106.000 6.350 106.350 ;
        RECT 7.060 97.230 7.200 106.350 ;
        RECT 7.000 96.910 7.260 97.230 ;
    END
  END select[0]
  PIN select[1]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 18.945 96.565 19.300 96.935 ;
      LAYER met1 ;
        RECT 18.470 96.800 18.790 96.860 ;
        RECT 18.945 96.800 19.235 96.845 ;
        RECT 18.470 96.660 19.235 96.800 ;
        RECT 18.470 96.600 18.790 96.660 ;
        RECT 18.945 96.615 19.235 96.660 ;
      LAYER met2 ;
        RECT 18.490 106.000 18.770 110.000 ;
        RECT 18.560 96.890 18.700 106.000 ;
        RECT 18.500 96.570 18.760 96.890 ;
    END
  END select[1]
  PIN select[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 32.795 96.595 33.155 97.175 ;
      LAYER met1 ;
        RECT 30.890 97.140 31.210 97.200 ;
        RECT 32.745 97.140 33.035 97.185 ;
        RECT 30.890 97.000 33.035 97.140 ;
        RECT 30.890 96.940 31.210 97.000 ;
        RECT 32.745 96.955 33.035 97.000 ;
      LAYER met2 ;
        RECT 30.910 106.000 31.190 110.000 ;
        RECT 30.980 97.230 31.120 106.000 ;
        RECT 30.920 96.910 31.180 97.230 ;
    END
  END select[2]
  PIN select[3]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 42.335 96.565 42.675 96.935 ;
      LAYER met1 ;
        RECT 42.850 97.280 43.170 97.540 ;
        RECT 42.405 96.800 42.695 96.845 ;
        RECT 42.940 96.800 43.080 97.280 ;
        RECT 42.405 96.660 43.080 96.800 ;
        RECT 42.405 96.615 42.695 96.660 ;
      LAYER met2 ;
        RECT 43.330 106.490 43.610 110.000 ;
        RECT 42.940 106.350 43.610 106.490 ;
        RECT 42.940 97.570 43.080 106.350 ;
        RECT 43.330 106.000 43.610 106.350 ;
        RECT 42.880 97.250 43.140 97.570 ;
    END
  END select[3]
  PIN vccd1
    ANTENNAGATEAREA 491.182983 ;
    ANTENNADIFFAREA 144.292252 ;
    PORT
      LAYER nwell ;
        RECT 5.330 93.785 44.350 96.615 ;
        RECT 5.330 88.345 44.350 91.175 ;
        RECT 5.330 82.905 44.350 85.735 ;
        RECT 5.330 77.465 44.350 80.295 ;
        RECT 5.330 72.025 44.350 74.855 ;
        RECT 5.330 66.585 44.350 69.415 ;
        RECT 5.330 61.145 44.350 63.975 ;
        RECT 5.330 55.705 44.350 58.535 ;
        RECT 5.330 50.265 44.350 53.095 ;
        RECT 5.330 44.825 44.350 47.655 ;
        RECT 5.330 39.385 44.350 42.215 ;
        RECT 5.330 33.945 44.350 36.775 ;
        RECT 5.330 28.505 44.350 31.335 ;
        RECT 5.330 23.065 44.350 25.895 ;
        RECT 5.330 17.625 44.350 20.455 ;
        RECT 5.330 12.185 44.350 15.015 ;
      LAYER li1 ;
        RECT 6.295 96.375 6.815 96.915 ;
        RECT 5.605 95.285 6.815 96.375 ;
        RECT 7.425 95.285 7.755 96.065 ;
        RECT 8.315 95.285 8.650 95.710 ;
        RECT 9.265 95.285 9.595 96.045 ;
        RECT 10.645 95.285 10.975 96.045 ;
        RECT 14.990 95.720 15.340 96.970 ;
        RECT 17.795 96.375 18.315 96.915 ;
        RECT 11.585 95.285 16.930 95.720 ;
        RECT 17.105 95.285 18.315 96.375 ;
        RECT 18.485 95.285 18.775 96.450 ;
        RECT 19.420 95.285 19.750 96.045 ;
        RECT 20.350 95.285 20.610 96.435 ;
        RECT 24.190 95.720 24.540 96.970 ;
        RECT 28.125 96.375 29.815 96.895 ;
        RECT 30.675 96.375 31.195 96.915 ;
        RECT 20.785 95.285 26.130 95.720 ;
        RECT 26.305 95.285 29.815 96.375 ;
        RECT 29.985 95.285 31.195 96.375 ;
        RECT 31.365 95.285 31.655 96.450 ;
        RECT 31.830 95.285 32.165 95.710 ;
        RECT 32.725 95.285 33.055 96.065 ;
        RECT 37.070 95.720 37.420 96.970 ;
        RECT 40.105 96.375 40.855 96.895 ;
        RECT 33.665 95.285 39.010 95.720 ;
        RECT 39.185 95.285 40.855 96.375 ;
        RECT 42.865 96.375 43.385 96.915 ;
        RECT 41.925 95.285 42.255 96.045 ;
        RECT 42.865 95.285 44.075 96.375 ;
        RECT 5.520 95.115 44.160 95.285 ;
        RECT 5.605 94.025 6.815 95.115 ;
        RECT 7.425 94.355 7.755 95.115 ;
        RECT 8.365 94.680 13.710 95.115 ;
        RECT 6.295 93.485 6.815 94.025 ;
        RECT 11.770 93.430 12.120 94.680 ;
        RECT 13.885 94.025 17.395 95.115 ;
        RECT 15.705 93.505 17.395 94.025 ;
        RECT 18.485 93.950 18.775 95.115 ;
        RECT 18.945 94.680 24.290 95.115 ;
        RECT 24.465 94.680 29.810 95.115 ;
        RECT 29.985 94.680 35.330 95.115 ;
        RECT 35.505 94.680 40.850 95.115 ;
        RECT 22.350 93.430 22.700 94.680 ;
        RECT 27.870 93.430 28.220 94.680 ;
        RECT 33.390 93.430 33.740 94.680 ;
        RECT 38.910 93.430 39.260 94.680 ;
        RECT 41.025 94.025 42.695 95.115 ;
        RECT 41.945 93.505 42.695 94.025 ;
        RECT 42.865 94.025 44.075 95.115 ;
        RECT 42.865 93.485 43.385 94.025 ;
        RECT 6.295 90.935 6.815 91.475 ;
        RECT 5.605 89.845 6.815 90.935 ;
        RECT 10.390 90.280 10.740 91.530 ;
        RECT 15.910 90.280 16.260 91.530 ;
        RECT 21.430 90.280 21.780 91.530 ;
        RECT 26.950 90.280 27.300 91.530 ;
        RECT 29.985 90.935 30.735 91.455 ;
        RECT 6.985 89.845 12.330 90.280 ;
        RECT 12.505 89.845 17.850 90.280 ;
        RECT 18.025 89.845 23.370 90.280 ;
        RECT 23.545 89.845 28.890 90.280 ;
        RECT 29.065 89.845 30.735 90.935 ;
        RECT 31.365 89.845 31.655 91.010 ;
        RECT 35.230 90.280 35.580 91.530 ;
        RECT 40.750 90.280 41.100 91.530 ;
        RECT 42.865 90.935 43.385 91.475 ;
        RECT 31.825 89.845 37.170 90.280 ;
        RECT 37.345 89.845 42.690 90.280 ;
        RECT 42.865 89.845 44.075 90.935 ;
        RECT 5.520 89.675 44.160 89.845 ;
        RECT 5.605 88.585 6.815 89.675 ;
        RECT 6.985 89.240 12.330 89.675 ;
        RECT 12.505 89.240 17.850 89.675 ;
        RECT 6.295 88.045 6.815 88.585 ;
        RECT 10.390 87.990 10.740 89.240 ;
        RECT 15.910 87.990 16.260 89.240 ;
        RECT 18.485 88.510 18.775 89.675 ;
        RECT 18.945 89.240 24.290 89.675 ;
        RECT 24.465 89.240 29.810 89.675 ;
        RECT 29.985 89.240 35.330 89.675 ;
        RECT 35.505 89.240 40.850 89.675 ;
        RECT 22.350 87.990 22.700 89.240 ;
        RECT 27.870 87.990 28.220 89.240 ;
        RECT 33.390 87.990 33.740 89.240 ;
        RECT 38.910 87.990 39.260 89.240 ;
        RECT 41.025 88.585 42.695 89.675 ;
        RECT 41.945 88.065 42.695 88.585 ;
        RECT 42.865 88.585 44.075 89.675 ;
        RECT 42.865 88.045 43.385 88.585 ;
        RECT 6.295 85.495 6.815 86.035 ;
        RECT 5.605 84.405 6.815 85.495 ;
        RECT 7.425 84.405 7.755 85.165 ;
        RECT 11.770 84.840 12.120 86.090 ;
        RECT 17.290 84.840 17.640 86.090 ;
        RECT 22.810 84.840 23.160 86.090 ;
        RECT 28.330 84.840 28.680 86.090 ;
        RECT 8.365 84.405 13.710 84.840 ;
        RECT 13.885 84.405 19.230 84.840 ;
        RECT 19.405 84.405 24.750 84.840 ;
        RECT 24.925 84.405 30.270 84.840 ;
        RECT 31.365 84.405 31.655 85.570 ;
        RECT 35.230 84.840 35.580 86.090 ;
        RECT 40.750 84.840 41.100 86.090 ;
        RECT 42.865 85.495 43.385 86.035 ;
        RECT 31.825 84.405 37.170 84.840 ;
        RECT 37.345 84.405 42.690 84.840 ;
        RECT 42.865 84.405 44.075 85.495 ;
        RECT 5.520 84.235 44.160 84.405 ;
        RECT 5.605 83.145 6.815 84.235 ;
        RECT 6.985 83.800 12.330 84.235 ;
        RECT 12.505 83.800 17.850 84.235 ;
        RECT 6.295 82.605 6.815 83.145 ;
        RECT 10.390 82.550 10.740 83.800 ;
        RECT 15.910 82.550 16.260 83.800 ;
        RECT 18.485 83.070 18.775 84.235 ;
        RECT 18.945 83.800 24.290 84.235 ;
        RECT 24.465 83.800 29.810 84.235 ;
        RECT 29.985 83.800 35.330 84.235 ;
        RECT 35.505 83.800 40.850 84.235 ;
        RECT 22.350 82.550 22.700 83.800 ;
        RECT 27.870 82.550 28.220 83.800 ;
        RECT 33.390 82.550 33.740 83.800 ;
        RECT 38.910 82.550 39.260 83.800 ;
        RECT 41.025 83.145 42.695 84.235 ;
        RECT 41.945 82.625 42.695 83.145 ;
        RECT 42.865 83.145 44.075 84.235 ;
        RECT 42.865 82.605 43.385 83.145 ;
        RECT 6.295 80.055 6.815 80.595 ;
        RECT 5.605 78.965 6.815 80.055 ;
        RECT 20.050 79.400 20.400 80.650 ;
        RECT 25.570 79.400 25.920 80.650 ;
        RECT 29.505 80.055 31.195 80.575 ;
        RECT 7.415 78.965 7.745 79.345 ;
        RECT 10.135 78.965 10.465 79.345 ;
        RECT 11.960 78.965 12.290 79.345 ;
        RECT 12.880 78.965 13.230 79.345 ;
        RECT 15.715 78.965 16.045 79.345 ;
        RECT 16.645 78.965 21.990 79.400 ;
        RECT 22.165 78.965 27.510 79.400 ;
        RECT 27.685 78.965 31.195 80.055 ;
        RECT 31.365 78.965 31.655 80.130 ;
        RECT 35.230 79.400 35.580 80.650 ;
        RECT 40.750 79.400 41.100 80.650 ;
        RECT 42.865 80.055 43.385 80.595 ;
        RECT 31.825 78.965 37.170 79.400 ;
        RECT 37.345 78.965 42.690 79.400 ;
        RECT 42.865 78.965 44.075 80.055 ;
        RECT 5.520 78.795 44.160 78.965 ;
        RECT 5.605 77.705 6.815 78.795 ;
        RECT 7.425 78.035 7.755 78.795 ;
        RECT 8.365 78.360 13.710 78.795 ;
        RECT 6.295 77.165 6.815 77.705 ;
        RECT 11.770 77.110 12.120 78.360 ;
        RECT 13.885 77.705 17.395 78.795 ;
        RECT 15.705 77.185 17.395 77.705 ;
        RECT 18.485 77.630 18.775 78.795 ;
        RECT 18.945 78.360 24.290 78.795 ;
        RECT 24.465 78.360 29.810 78.795 ;
        RECT 29.985 78.360 35.330 78.795 ;
        RECT 35.505 78.360 40.850 78.795 ;
        RECT 22.350 77.110 22.700 78.360 ;
        RECT 27.870 77.110 28.220 78.360 ;
        RECT 33.390 77.110 33.740 78.360 ;
        RECT 38.910 77.110 39.260 78.360 ;
        RECT 41.025 77.705 42.695 78.795 ;
        RECT 41.945 77.185 42.695 77.705 ;
        RECT 42.865 77.705 44.075 78.795 ;
        RECT 42.865 77.165 43.385 77.705 ;
        RECT 6.295 74.615 6.815 75.155 ;
        RECT 5.605 73.525 6.815 74.615 ;
        RECT 20.050 73.960 20.400 75.210 ;
        RECT 25.570 73.960 25.920 75.210 ;
        RECT 29.505 74.615 31.195 75.135 ;
        RECT 7.415 73.525 7.745 73.905 ;
        RECT 10.135 73.525 10.465 73.905 ;
        RECT 11.960 73.525 12.290 73.905 ;
        RECT 12.880 73.525 13.230 73.905 ;
        RECT 15.715 73.525 16.045 73.905 ;
        RECT 16.645 73.525 21.990 73.960 ;
        RECT 22.165 73.525 27.510 73.960 ;
        RECT 27.685 73.525 31.195 74.615 ;
        RECT 31.365 73.525 31.655 74.690 ;
        RECT 35.230 73.960 35.580 75.210 ;
        RECT 40.750 73.960 41.100 75.210 ;
        RECT 42.865 74.615 43.385 75.155 ;
        RECT 31.825 73.525 37.170 73.960 ;
        RECT 37.345 73.525 42.690 73.960 ;
        RECT 42.865 73.525 44.075 74.615 ;
        RECT 5.520 73.355 44.160 73.525 ;
        RECT 5.605 72.265 6.815 73.355 ;
        RECT 7.425 72.595 7.755 73.355 ;
        RECT 8.365 72.265 10.955 73.355 ;
        RECT 6.295 71.725 6.815 72.265 ;
        RECT 9.745 71.745 10.955 72.265 ;
        RECT 12.095 72.215 12.265 73.355 ;
        RECT 14.635 72.595 14.805 73.355 ;
        RECT 15.725 72.265 18.315 73.355 ;
        RECT 17.105 71.745 18.315 72.265 ;
        RECT 18.485 72.190 18.775 73.355 ;
        RECT 18.945 72.920 24.290 73.355 ;
        RECT 24.465 72.920 29.810 73.355 ;
        RECT 29.985 72.920 35.330 73.355 ;
        RECT 35.505 72.920 40.850 73.355 ;
        RECT 22.350 71.670 22.700 72.920 ;
        RECT 27.870 71.670 28.220 72.920 ;
        RECT 33.390 71.670 33.740 72.920 ;
        RECT 38.910 71.670 39.260 72.920 ;
        RECT 41.025 72.265 42.695 73.355 ;
        RECT 41.945 71.745 42.695 72.265 ;
        RECT 42.865 72.265 44.075 73.355 ;
        RECT 42.865 71.725 43.385 72.265 ;
        RECT 6.295 69.175 6.815 69.715 ;
        RECT 5.605 68.085 6.815 69.175 ;
        RECT 10.390 68.520 10.740 69.770 ;
        RECT 15.910 68.520 16.260 69.770 ;
        RECT 21.430 68.520 21.780 69.770 ;
        RECT 26.950 68.520 27.300 69.770 ;
        RECT 29.985 69.175 30.735 69.695 ;
        RECT 6.985 68.085 12.330 68.520 ;
        RECT 12.505 68.085 17.850 68.520 ;
        RECT 18.025 68.085 23.370 68.520 ;
        RECT 23.545 68.085 28.890 68.520 ;
        RECT 29.065 68.085 30.735 69.175 ;
        RECT 31.365 68.085 31.655 69.250 ;
        RECT 35.230 68.520 35.580 69.770 ;
        RECT 40.750 68.520 41.100 69.770 ;
        RECT 42.865 69.175 43.385 69.715 ;
        RECT 31.825 68.085 37.170 68.520 ;
        RECT 37.345 68.085 42.690 68.520 ;
        RECT 42.865 68.085 44.075 69.175 ;
        RECT 5.520 67.915 44.160 68.085 ;
        RECT 5.605 66.825 6.815 67.915 ;
        RECT 7.425 67.155 7.755 67.915 ;
        RECT 8.365 67.480 13.710 67.915 ;
        RECT 6.295 66.285 6.815 66.825 ;
        RECT 11.770 66.230 12.120 67.480 ;
        RECT 13.885 66.825 17.395 67.915 ;
        RECT 15.705 66.305 17.395 66.825 ;
        RECT 18.485 66.750 18.775 67.915 ;
        RECT 18.945 67.480 24.290 67.915 ;
        RECT 24.465 67.480 29.810 67.915 ;
        RECT 29.985 67.480 35.330 67.915 ;
        RECT 35.505 67.480 40.850 67.915 ;
        RECT 22.350 66.230 22.700 67.480 ;
        RECT 27.870 66.230 28.220 67.480 ;
        RECT 33.390 66.230 33.740 67.480 ;
        RECT 38.910 66.230 39.260 67.480 ;
        RECT 41.025 66.825 42.695 67.915 ;
        RECT 41.945 66.305 42.695 66.825 ;
        RECT 42.865 66.825 44.075 67.915 ;
        RECT 42.865 66.285 43.385 66.825 ;
        RECT 6.295 63.735 6.815 64.275 ;
        RECT 5.605 62.645 6.815 63.735 ;
        RECT 10.390 63.080 10.740 64.330 ;
        RECT 15.910 63.080 16.260 64.330 ;
        RECT 21.430 63.080 21.780 64.330 ;
        RECT 26.950 63.080 27.300 64.330 ;
        RECT 29.985 63.735 30.735 64.255 ;
        RECT 6.985 62.645 12.330 63.080 ;
        RECT 12.505 62.645 17.850 63.080 ;
        RECT 18.025 62.645 23.370 63.080 ;
        RECT 23.545 62.645 28.890 63.080 ;
        RECT 29.065 62.645 30.735 63.735 ;
        RECT 31.365 62.645 31.655 63.810 ;
        RECT 35.230 63.080 35.580 64.330 ;
        RECT 40.750 63.080 41.100 64.330 ;
        RECT 42.865 63.735 43.385 64.275 ;
        RECT 31.825 62.645 37.170 63.080 ;
        RECT 37.345 62.645 42.690 63.080 ;
        RECT 42.865 62.645 44.075 63.735 ;
        RECT 5.520 62.475 44.160 62.645 ;
        RECT 5.605 61.385 6.815 62.475 ;
        RECT 6.985 61.385 10.495 62.475 ;
        RECT 6.295 60.845 6.815 61.385 ;
        RECT 8.805 60.865 10.495 61.385 ;
        RECT 12.455 61.335 12.785 62.475 ;
        RECT 12.965 62.040 18.310 62.475 ;
        RECT 16.370 60.790 16.720 62.040 ;
        RECT 18.485 61.310 18.775 62.475 ;
        RECT 18.945 62.040 24.290 62.475 ;
        RECT 24.465 62.040 29.810 62.475 ;
        RECT 29.985 62.040 35.330 62.475 ;
        RECT 35.505 62.040 40.850 62.475 ;
        RECT 22.350 60.790 22.700 62.040 ;
        RECT 27.870 60.790 28.220 62.040 ;
        RECT 33.390 60.790 33.740 62.040 ;
        RECT 38.910 60.790 39.260 62.040 ;
        RECT 41.025 61.385 42.695 62.475 ;
        RECT 41.945 60.865 42.695 61.385 ;
        RECT 42.865 61.385 44.075 62.475 ;
        RECT 42.865 60.845 43.385 61.385 ;
        RECT 6.295 58.295 6.815 58.835 ;
        RECT 10.185 58.295 11.875 58.815 ;
        RECT 5.605 57.205 6.815 58.295 ;
        RECT 7.425 57.205 7.755 57.965 ;
        RECT 8.365 57.205 11.875 58.295 ;
        RECT 13.535 57.205 13.705 57.645 ;
        RECT 18.670 57.640 19.020 58.890 ;
        RECT 24.190 57.640 24.540 58.890 ;
        RECT 28.125 58.295 29.815 58.815 ;
        RECT 30.675 58.295 31.195 58.835 ;
        RECT 14.310 57.205 14.640 57.565 ;
        RECT 15.265 57.205 20.610 57.640 ;
        RECT 20.785 57.205 26.130 57.640 ;
        RECT 26.305 57.205 29.815 58.295 ;
        RECT 29.985 57.205 31.195 58.295 ;
        RECT 31.365 57.205 31.655 58.370 ;
        RECT 35.230 57.640 35.580 58.890 ;
        RECT 40.750 57.640 41.100 58.890 ;
        RECT 42.865 58.295 43.385 58.835 ;
        RECT 31.825 57.205 37.170 57.640 ;
        RECT 37.345 57.205 42.690 57.640 ;
        RECT 42.865 57.205 44.075 58.295 ;
        RECT 5.520 57.035 44.160 57.205 ;
        RECT 5.605 55.945 6.815 57.035 ;
        RECT 6.985 56.600 12.330 57.035 ;
        RECT 12.505 56.600 17.850 57.035 ;
        RECT 6.295 55.405 6.815 55.945 ;
        RECT 10.390 55.350 10.740 56.600 ;
        RECT 15.910 55.350 16.260 56.600 ;
        RECT 18.485 55.870 18.775 57.035 ;
        RECT 18.945 56.600 24.290 57.035 ;
        RECT 24.465 56.600 29.810 57.035 ;
        RECT 29.985 56.600 35.330 57.035 ;
        RECT 22.350 55.350 22.700 56.600 ;
        RECT 27.870 55.350 28.220 56.600 ;
        RECT 33.390 55.350 33.740 56.600 ;
        RECT 35.595 56.235 35.765 57.035 ;
        RECT 36.435 56.235 36.605 57.035 ;
        RECT 37.275 56.235 37.445 57.035 ;
        RECT 38.035 56.235 38.365 57.035 ;
        RECT 38.875 56.235 39.205 57.035 ;
        RECT 39.715 56.235 40.045 57.035 ;
        RECT 40.555 56.235 40.885 57.035 ;
        RECT 41.395 56.235 41.725 57.035 ;
        RECT 42.235 55.885 42.565 57.035 ;
        RECT 42.865 55.945 44.075 57.035 ;
        RECT 42.865 55.405 43.385 55.945 ;
        RECT 6.295 52.855 6.815 53.395 ;
        RECT 5.605 51.765 6.815 52.855 ;
        RECT 7.425 51.765 7.755 52.525 ;
        RECT 11.770 52.200 12.120 53.450 ;
        RECT 17.290 52.200 17.640 53.450 ;
        RECT 22.810 52.200 23.160 53.450 ;
        RECT 28.330 52.200 28.680 53.450 ;
        RECT 8.365 51.765 13.710 52.200 ;
        RECT 13.885 51.765 19.230 52.200 ;
        RECT 19.405 51.765 24.750 52.200 ;
        RECT 24.925 51.765 30.270 52.200 ;
        RECT 31.365 51.765 31.655 52.930 ;
        RECT 35.230 52.200 35.580 53.450 ;
        RECT 40.750 52.200 41.100 53.450 ;
        RECT 42.865 52.855 43.385 53.395 ;
        RECT 31.825 51.765 37.170 52.200 ;
        RECT 37.345 51.765 42.690 52.200 ;
        RECT 42.865 51.765 44.075 52.855 ;
        RECT 5.520 51.595 44.160 51.765 ;
        RECT 5.605 50.505 6.815 51.595 ;
        RECT 6.985 51.160 12.330 51.595 ;
        RECT 12.505 51.160 17.850 51.595 ;
        RECT 6.295 49.965 6.815 50.505 ;
        RECT 10.390 49.910 10.740 51.160 ;
        RECT 15.910 49.910 16.260 51.160 ;
        RECT 18.485 50.430 18.775 51.595 ;
        RECT 18.945 51.160 24.290 51.595 ;
        RECT 24.465 51.160 29.810 51.595 ;
        RECT 29.985 51.160 35.330 51.595 ;
        RECT 35.505 51.160 40.850 51.595 ;
        RECT 22.350 49.910 22.700 51.160 ;
        RECT 27.870 49.910 28.220 51.160 ;
        RECT 33.390 49.910 33.740 51.160 ;
        RECT 38.910 49.910 39.260 51.160 ;
        RECT 41.025 50.505 42.695 51.595 ;
        RECT 41.945 49.985 42.695 50.505 ;
        RECT 42.865 50.505 44.075 51.595 ;
        RECT 42.865 49.965 43.385 50.505 ;
        RECT 6.295 47.415 6.815 47.955 ;
        RECT 5.605 46.325 6.815 47.415 ;
        RECT 7.715 46.325 8.045 46.835 ;
        RECT 13.150 46.760 13.500 48.010 ;
        RECT 18.670 46.760 19.020 48.010 ;
        RECT 24.190 46.760 24.540 48.010 ;
        RECT 28.125 47.415 29.815 47.935 ;
        RECT 30.675 47.415 31.195 47.955 ;
        RECT 9.745 46.325 15.090 46.760 ;
        RECT 15.265 46.325 20.610 46.760 ;
        RECT 20.785 46.325 26.130 46.760 ;
        RECT 26.305 46.325 29.815 47.415 ;
        RECT 29.985 46.325 31.195 47.415 ;
        RECT 31.365 46.325 31.655 47.490 ;
        RECT 35.230 46.760 35.580 48.010 ;
        RECT 40.750 46.760 41.100 48.010 ;
        RECT 42.865 47.415 43.385 47.955 ;
        RECT 31.825 46.325 37.170 46.760 ;
        RECT 37.345 46.325 42.690 46.760 ;
        RECT 42.865 46.325 44.075 47.415 ;
        RECT 5.520 46.155 44.160 46.325 ;
        RECT 5.605 45.065 6.815 46.155 ;
        RECT 7.425 45.395 7.755 46.155 ;
        RECT 8.365 45.720 13.710 46.155 ;
        RECT 6.295 44.525 6.815 45.065 ;
        RECT 11.770 44.470 12.120 45.720 ;
        RECT 13.885 45.065 17.395 46.155 ;
        RECT 15.705 44.545 17.395 45.065 ;
        RECT 18.485 44.990 18.775 46.155 ;
        RECT 18.945 45.720 24.290 46.155 ;
        RECT 24.465 45.720 29.810 46.155 ;
        RECT 29.985 45.720 35.330 46.155 ;
        RECT 35.505 45.720 40.850 46.155 ;
        RECT 22.350 44.470 22.700 45.720 ;
        RECT 27.870 44.470 28.220 45.720 ;
        RECT 33.390 44.470 33.740 45.720 ;
        RECT 38.910 44.470 39.260 45.720 ;
        RECT 41.025 45.065 42.695 46.155 ;
        RECT 41.945 44.545 42.695 45.065 ;
        RECT 42.865 45.065 44.075 46.155 ;
        RECT 42.865 44.525 43.385 45.065 ;
        RECT 6.295 41.975 6.815 42.515 ;
        RECT 5.605 40.885 6.815 41.975 ;
        RECT 7.735 40.885 7.905 41.645 ;
        RECT 10.275 40.885 10.445 42.025 ;
        RECT 11.590 40.885 11.920 41.600 ;
        RECT 18.210 41.320 18.560 42.570 ;
        RECT 23.730 41.320 24.080 42.570 ;
        RECT 29.250 41.320 29.600 42.570 ;
        RECT 14.805 40.885 20.150 41.320 ;
        RECT 20.325 40.885 25.670 41.320 ;
        RECT 25.845 40.885 31.190 41.320 ;
        RECT 31.365 40.885 31.655 42.050 ;
        RECT 35.230 41.320 35.580 42.570 ;
        RECT 40.750 41.320 41.100 42.570 ;
        RECT 42.865 41.975 43.385 42.515 ;
        RECT 31.825 40.885 37.170 41.320 ;
        RECT 37.345 40.885 42.690 41.320 ;
        RECT 42.865 40.885 44.075 41.975 ;
        RECT 5.520 40.715 44.160 40.885 ;
        RECT 5.605 39.625 6.815 40.715 ;
        RECT 6.985 40.205 7.245 40.715 ;
        RECT 7.905 40.210 8.520 40.715 ;
        RECT 8.325 40.035 8.520 40.210 ;
        RECT 9.335 40.170 9.550 40.715 ;
        RECT 10.205 40.280 15.550 40.715 ;
        RECT 8.325 39.845 8.655 40.035 ;
        RECT 6.295 39.085 6.815 39.625 ;
        RECT 13.610 39.030 13.960 40.280 ;
        RECT 15.725 39.625 18.315 40.715 ;
        RECT 17.105 39.105 18.315 39.625 ;
        RECT 18.485 39.550 18.775 40.715 ;
        RECT 18.945 40.280 24.290 40.715 ;
        RECT 24.465 40.280 29.810 40.715 ;
        RECT 29.985 40.280 35.330 40.715 ;
        RECT 35.505 40.280 40.850 40.715 ;
        RECT 22.350 39.030 22.700 40.280 ;
        RECT 27.870 39.030 28.220 40.280 ;
        RECT 33.390 39.030 33.740 40.280 ;
        RECT 38.910 39.030 39.260 40.280 ;
        RECT 41.025 39.625 42.695 40.715 ;
        RECT 41.945 39.105 42.695 39.625 ;
        RECT 42.865 39.625 44.075 40.715 ;
        RECT 42.865 39.085 43.385 39.625 ;
        RECT 6.295 36.535 6.815 37.075 ;
        RECT 5.605 35.445 6.815 36.535 ;
        RECT 7.425 35.445 7.755 36.205 ;
        RECT 11.770 35.880 12.120 37.130 ;
        RECT 17.290 35.880 17.640 37.130 ;
        RECT 22.810 35.880 23.160 37.130 ;
        RECT 28.330 35.880 28.680 37.130 ;
        RECT 8.365 35.445 13.710 35.880 ;
        RECT 13.885 35.445 19.230 35.880 ;
        RECT 19.405 35.445 24.750 35.880 ;
        RECT 24.925 35.445 30.270 35.880 ;
        RECT 31.365 35.445 31.655 36.610 ;
        RECT 35.230 35.880 35.580 37.130 ;
        RECT 40.750 35.880 41.100 37.130 ;
        RECT 42.865 36.535 43.385 37.075 ;
        RECT 31.825 35.445 37.170 35.880 ;
        RECT 37.345 35.445 42.690 35.880 ;
        RECT 42.865 35.445 44.075 36.535 ;
        RECT 5.520 35.275 44.160 35.445 ;
        RECT 5.605 34.185 6.815 35.275 ;
        RECT 6.985 34.185 8.195 35.275 ;
        RECT 8.865 34.815 9.115 35.275 ;
        RECT 9.795 34.815 10.045 35.275 ;
        RECT 11.115 34.815 11.365 35.275 ;
        RECT 12.045 34.840 17.390 35.275 ;
        RECT 6.295 33.645 6.815 34.185 ;
        RECT 7.675 33.645 8.195 34.185 ;
        RECT 15.450 33.590 15.800 34.840 ;
        RECT 18.485 34.110 18.775 35.275 ;
        RECT 18.945 34.840 24.290 35.275 ;
        RECT 24.465 34.840 29.810 35.275 ;
        RECT 29.985 34.840 35.330 35.275 ;
        RECT 35.505 34.840 40.850 35.275 ;
        RECT 22.350 33.590 22.700 34.840 ;
        RECT 27.870 33.590 28.220 34.840 ;
        RECT 33.390 33.590 33.740 34.840 ;
        RECT 38.910 33.590 39.260 34.840 ;
        RECT 41.025 34.185 42.695 35.275 ;
        RECT 41.945 33.665 42.695 34.185 ;
        RECT 42.865 34.185 44.075 35.275 ;
        RECT 42.865 33.645 43.385 34.185 ;
        RECT 6.295 31.095 6.815 31.635 ;
        RECT 5.605 30.005 6.815 31.095 ;
        RECT 7.905 30.005 8.165 31.145 ;
        RECT 10.190 30.005 10.470 30.805 ;
        RECT 11.885 30.005 12.170 30.805 ;
        RECT 12.840 30.005 13.090 31.145 ;
        RECT 17.290 30.440 17.640 31.690 ;
        RECT 22.810 30.440 23.160 31.690 ;
        RECT 28.330 30.440 28.680 31.690 ;
        RECT 13.885 30.005 19.230 30.440 ;
        RECT 19.405 30.005 24.750 30.440 ;
        RECT 24.925 30.005 30.270 30.440 ;
        RECT 31.365 30.005 31.655 31.170 ;
        RECT 35.230 30.440 35.580 31.690 ;
        RECT 40.750 30.440 41.100 31.690 ;
        RECT 42.865 31.095 43.385 31.635 ;
        RECT 31.825 30.005 37.170 30.440 ;
        RECT 37.345 30.005 42.690 30.440 ;
        RECT 42.865 30.005 44.075 31.095 ;
        RECT 5.520 29.835 44.160 30.005 ;
        RECT 5.605 28.745 6.815 29.835 ;
        RECT 7.425 29.075 7.755 29.835 ;
        RECT 6.295 28.205 6.815 28.745 ;
        RECT 8.825 28.695 9.085 29.835 ;
        RECT 9.755 28.695 10.035 29.835 ;
        RECT 10.205 29.400 15.550 29.835 ;
        RECT 13.610 28.150 13.960 29.400 ;
        RECT 15.725 28.745 18.315 29.835 ;
        RECT 17.105 28.225 18.315 28.745 ;
        RECT 18.485 28.670 18.775 29.835 ;
        RECT 18.945 29.400 24.290 29.835 ;
        RECT 24.465 29.400 29.810 29.835 ;
        RECT 29.985 29.400 35.330 29.835 ;
        RECT 35.505 29.400 40.850 29.835 ;
        RECT 22.350 28.150 22.700 29.400 ;
        RECT 27.870 28.150 28.220 29.400 ;
        RECT 33.390 28.150 33.740 29.400 ;
        RECT 38.910 28.150 39.260 29.400 ;
        RECT 41.025 28.745 42.695 29.835 ;
        RECT 41.945 28.225 42.695 28.745 ;
        RECT 42.865 28.745 44.075 29.835 ;
        RECT 42.865 28.205 43.385 28.745 ;
        RECT 6.295 25.655 6.815 26.195 ;
        RECT 5.605 24.565 6.815 25.655 ;
        RECT 7.735 24.565 7.905 25.325 ;
        RECT 10.275 24.565 10.445 25.705 ;
        RECT 14.530 25.000 14.880 26.250 ;
        RECT 20.050 25.000 20.400 26.250 ;
        RECT 25.570 25.000 25.920 26.250 ;
        RECT 29.505 25.655 31.195 26.175 ;
        RECT 11.125 24.565 16.470 25.000 ;
        RECT 16.645 24.565 21.990 25.000 ;
        RECT 22.165 24.565 27.510 25.000 ;
        RECT 27.685 24.565 31.195 25.655 ;
        RECT 31.365 24.565 31.655 25.730 ;
        RECT 35.230 25.000 35.580 26.250 ;
        RECT 40.750 25.000 41.100 26.250 ;
        RECT 42.865 25.655 43.385 26.195 ;
        RECT 31.825 24.565 37.170 25.000 ;
        RECT 37.345 24.565 42.690 25.000 ;
        RECT 42.865 24.565 44.075 25.655 ;
        RECT 5.520 24.395 44.160 24.565 ;
        RECT 5.605 23.305 6.815 24.395 ;
        RECT 7.425 23.635 7.755 24.395 ;
        RECT 8.365 23.960 13.710 24.395 ;
        RECT 6.295 22.765 6.815 23.305 ;
        RECT 11.770 22.710 12.120 23.960 ;
        RECT 13.885 23.305 17.395 24.395 ;
        RECT 15.705 22.785 17.395 23.305 ;
        RECT 18.485 23.230 18.775 24.395 ;
        RECT 18.945 23.960 24.290 24.395 ;
        RECT 24.465 23.960 29.810 24.395 ;
        RECT 29.985 23.960 35.330 24.395 ;
        RECT 35.505 23.960 40.850 24.395 ;
        RECT 22.350 22.710 22.700 23.960 ;
        RECT 27.870 22.710 28.220 23.960 ;
        RECT 33.390 22.710 33.740 23.960 ;
        RECT 38.910 22.710 39.260 23.960 ;
        RECT 41.025 23.305 42.695 24.395 ;
        RECT 41.945 22.785 42.695 23.305 ;
        RECT 42.865 23.305 44.075 24.395 ;
        RECT 42.865 22.765 43.385 23.305 ;
        RECT 6.295 20.215 6.815 20.755 ;
        RECT 5.605 19.125 6.815 20.215 ;
        RECT 10.390 19.560 10.740 20.810 ;
        RECT 15.910 19.560 16.260 20.810 ;
        RECT 21.430 19.560 21.780 20.810 ;
        RECT 26.950 19.560 27.300 20.810 ;
        RECT 29.985 20.215 30.735 20.735 ;
        RECT 6.985 19.125 12.330 19.560 ;
        RECT 12.505 19.125 17.850 19.560 ;
        RECT 18.025 19.125 23.370 19.560 ;
        RECT 23.545 19.125 28.890 19.560 ;
        RECT 29.065 19.125 30.735 20.215 ;
        RECT 31.365 19.125 31.655 20.290 ;
        RECT 35.230 19.560 35.580 20.810 ;
        RECT 40.750 19.560 41.100 20.810 ;
        RECT 42.865 20.215 43.385 20.755 ;
        RECT 31.825 19.125 37.170 19.560 ;
        RECT 37.345 19.125 42.690 19.560 ;
        RECT 42.865 19.125 44.075 20.215 ;
        RECT 5.520 18.955 44.160 19.125 ;
        RECT 5.605 17.865 6.815 18.955 ;
        RECT 7.425 18.195 7.755 18.955 ;
        RECT 8.365 18.520 13.710 18.955 ;
        RECT 6.295 17.325 6.815 17.865 ;
        RECT 11.770 17.270 12.120 18.520 ;
        RECT 13.885 17.865 17.395 18.955 ;
        RECT 15.705 17.345 17.395 17.865 ;
        RECT 18.485 17.790 18.775 18.955 ;
        RECT 18.945 18.520 24.290 18.955 ;
        RECT 24.465 18.520 29.810 18.955 ;
        RECT 29.985 18.520 35.330 18.955 ;
        RECT 35.505 18.520 40.850 18.955 ;
        RECT 22.350 17.270 22.700 18.520 ;
        RECT 27.870 17.270 28.220 18.520 ;
        RECT 33.390 17.270 33.740 18.520 ;
        RECT 38.910 17.270 39.260 18.520 ;
        RECT 41.025 17.865 42.695 18.955 ;
        RECT 41.945 17.345 42.695 17.865 ;
        RECT 42.865 17.865 44.075 18.955 ;
        RECT 42.865 17.325 43.385 17.865 ;
        RECT 6.295 14.775 6.815 15.315 ;
        RECT 5.605 13.685 6.815 14.775 ;
        RECT 10.390 14.120 10.740 15.370 ;
        RECT 15.910 14.120 16.260 15.370 ;
        RECT 21.430 14.120 21.780 15.370 ;
        RECT 26.950 14.120 27.300 15.370 ;
        RECT 29.985 14.775 30.735 15.295 ;
        RECT 6.985 13.685 12.330 14.120 ;
        RECT 12.505 13.685 17.850 14.120 ;
        RECT 18.025 13.685 23.370 14.120 ;
        RECT 23.545 13.685 28.890 14.120 ;
        RECT 29.065 13.685 30.735 14.775 ;
        RECT 31.365 13.685 31.655 14.850 ;
        RECT 35.230 14.120 35.580 15.370 ;
        RECT 40.750 14.120 41.100 15.370 ;
        RECT 42.865 14.775 43.385 15.315 ;
        RECT 31.825 13.685 37.170 14.120 ;
        RECT 37.345 13.685 42.690 14.120 ;
        RECT 42.865 13.685 44.075 14.775 ;
        RECT 5.520 13.515 44.160 13.685 ;
        RECT 5.605 12.425 6.815 13.515 ;
        RECT 7.425 12.755 7.755 13.515 ;
        RECT 8.805 12.755 9.135 13.515 ;
        RECT 9.745 13.080 15.090 13.515 ;
        RECT 6.295 11.885 6.815 12.425 ;
        RECT 13.150 11.830 13.500 13.080 ;
        RECT 15.265 12.425 17.855 13.515 ;
        RECT 16.645 11.905 17.855 12.425 ;
        RECT 18.485 12.350 18.775 13.515 ;
        RECT 18.945 13.080 24.290 13.515 ;
        RECT 24.465 13.080 29.810 13.515 ;
        RECT 22.350 11.830 22.700 13.080 ;
        RECT 27.870 11.830 28.220 13.080 ;
        RECT 29.985 12.425 31.195 13.515 ;
        RECT 30.675 11.885 31.195 12.425 ;
        RECT 31.365 12.350 31.655 13.515 ;
        RECT 31.825 13.080 37.170 13.515 ;
        RECT 37.345 13.080 42.690 13.515 ;
        RECT 35.230 11.830 35.580 13.080 ;
        RECT 40.750 11.830 41.100 13.080 ;
        RECT 42.865 12.425 44.075 13.515 ;
        RECT 42.865 11.885 43.385 12.425 ;
      LAYER met1 ;
        RECT 5.520 94.960 44.160 95.440 ;
        RECT 5.520 89.520 44.160 90.000 ;
        RECT 5.520 84.080 44.160 84.560 ;
        RECT 5.520 78.640 44.160 79.120 ;
        RECT 5.520 73.200 44.160 73.680 ;
        RECT 5.520 67.760 44.160 68.240 ;
        RECT 5.520 62.320 44.160 62.800 ;
        RECT 5.520 56.880 44.160 57.360 ;
        RECT 5.520 51.440 44.160 51.920 ;
        RECT 5.520 46.000 44.160 46.480 ;
        RECT 5.520 40.560 44.160 41.040 ;
        RECT 5.520 35.120 44.160 35.600 ;
        RECT 5.520 29.680 44.160 30.160 ;
        RECT 5.520 24.240 44.160 24.720 ;
        RECT 5.520 18.800 44.160 19.280 ;
        RECT 5.520 13.360 44.160 13.840 ;
      LAYER met2 ;
        RECT 9.580 95.015 11.120 95.385 ;
        RECT 19.240 95.015 20.780 95.385 ;
        RECT 28.900 95.015 30.440 95.385 ;
        RECT 38.560 95.015 40.100 95.385 ;
        RECT 9.580 89.575 11.120 89.945 ;
        RECT 19.240 89.575 20.780 89.945 ;
        RECT 28.900 89.575 30.440 89.945 ;
        RECT 38.560 89.575 40.100 89.945 ;
        RECT 9.580 84.135 11.120 84.505 ;
        RECT 19.240 84.135 20.780 84.505 ;
        RECT 28.900 84.135 30.440 84.505 ;
        RECT 38.560 84.135 40.100 84.505 ;
        RECT 9.580 78.695 11.120 79.065 ;
        RECT 19.240 78.695 20.780 79.065 ;
        RECT 28.900 78.695 30.440 79.065 ;
        RECT 38.560 78.695 40.100 79.065 ;
        RECT 9.580 73.255 11.120 73.625 ;
        RECT 19.240 73.255 20.780 73.625 ;
        RECT 28.900 73.255 30.440 73.625 ;
        RECT 38.560 73.255 40.100 73.625 ;
        RECT 9.580 67.815 11.120 68.185 ;
        RECT 19.240 67.815 20.780 68.185 ;
        RECT 28.900 67.815 30.440 68.185 ;
        RECT 38.560 67.815 40.100 68.185 ;
        RECT 9.580 62.375 11.120 62.745 ;
        RECT 19.240 62.375 20.780 62.745 ;
        RECT 28.900 62.375 30.440 62.745 ;
        RECT 38.560 62.375 40.100 62.745 ;
        RECT 9.580 56.935 11.120 57.305 ;
        RECT 19.240 56.935 20.780 57.305 ;
        RECT 28.900 56.935 30.440 57.305 ;
        RECT 38.560 56.935 40.100 57.305 ;
        RECT 9.580 51.495 11.120 51.865 ;
        RECT 19.240 51.495 20.780 51.865 ;
        RECT 28.900 51.495 30.440 51.865 ;
        RECT 38.560 51.495 40.100 51.865 ;
        RECT 9.580 46.055 11.120 46.425 ;
        RECT 19.240 46.055 20.780 46.425 ;
        RECT 28.900 46.055 30.440 46.425 ;
        RECT 38.560 46.055 40.100 46.425 ;
        RECT 9.580 40.615 11.120 40.985 ;
        RECT 19.240 40.615 20.780 40.985 ;
        RECT 28.900 40.615 30.440 40.985 ;
        RECT 38.560 40.615 40.100 40.985 ;
        RECT 9.580 35.175 11.120 35.545 ;
        RECT 19.240 35.175 20.780 35.545 ;
        RECT 28.900 35.175 30.440 35.545 ;
        RECT 38.560 35.175 40.100 35.545 ;
        RECT 9.580 29.735 11.120 30.105 ;
        RECT 19.240 29.735 20.780 30.105 ;
        RECT 28.900 29.735 30.440 30.105 ;
        RECT 38.560 29.735 40.100 30.105 ;
        RECT 9.580 24.295 11.120 24.665 ;
        RECT 19.240 24.295 20.780 24.665 ;
        RECT 28.900 24.295 30.440 24.665 ;
        RECT 38.560 24.295 40.100 24.665 ;
        RECT 9.580 18.855 11.120 19.225 ;
        RECT 19.240 18.855 20.780 19.225 ;
        RECT 28.900 18.855 30.440 19.225 ;
        RECT 38.560 18.855 40.100 19.225 ;
        RECT 9.580 13.415 11.120 13.785 ;
        RECT 19.240 13.415 20.780 13.785 ;
        RECT 28.900 13.415 30.440 13.785 ;
        RECT 38.560 13.415 40.100 13.785 ;
      LAYER met3 ;
        RECT 9.560 95.035 11.140 95.365 ;
        RECT 19.220 95.035 20.800 95.365 ;
        RECT 28.880 95.035 30.460 95.365 ;
        RECT 38.540 95.035 40.120 95.365 ;
        RECT 9.560 89.595 11.140 89.925 ;
        RECT 19.220 89.595 20.800 89.925 ;
        RECT 28.880 89.595 30.460 89.925 ;
        RECT 38.540 89.595 40.120 89.925 ;
        RECT 9.560 84.155 11.140 84.485 ;
        RECT 19.220 84.155 20.800 84.485 ;
        RECT 28.880 84.155 30.460 84.485 ;
        RECT 38.540 84.155 40.120 84.485 ;
        RECT 9.560 78.715 11.140 79.045 ;
        RECT 19.220 78.715 20.800 79.045 ;
        RECT 28.880 78.715 30.460 79.045 ;
        RECT 38.540 78.715 40.120 79.045 ;
        RECT 9.560 73.275 11.140 73.605 ;
        RECT 19.220 73.275 20.800 73.605 ;
        RECT 28.880 73.275 30.460 73.605 ;
        RECT 38.540 73.275 40.120 73.605 ;
        RECT 9.560 67.835 11.140 68.165 ;
        RECT 19.220 67.835 20.800 68.165 ;
        RECT 28.880 67.835 30.460 68.165 ;
        RECT 38.540 67.835 40.120 68.165 ;
        RECT 9.560 62.395 11.140 62.725 ;
        RECT 19.220 62.395 20.800 62.725 ;
        RECT 28.880 62.395 30.460 62.725 ;
        RECT 38.540 62.395 40.120 62.725 ;
        RECT 9.560 56.955 11.140 57.285 ;
        RECT 19.220 56.955 20.800 57.285 ;
        RECT 28.880 56.955 30.460 57.285 ;
        RECT 38.540 56.955 40.120 57.285 ;
        RECT 9.560 51.515 11.140 51.845 ;
        RECT 19.220 51.515 20.800 51.845 ;
        RECT 28.880 51.515 30.460 51.845 ;
        RECT 38.540 51.515 40.120 51.845 ;
        RECT 9.560 46.075 11.140 46.405 ;
        RECT 19.220 46.075 20.800 46.405 ;
        RECT 28.880 46.075 30.460 46.405 ;
        RECT 38.540 46.075 40.120 46.405 ;
        RECT 9.560 40.635 11.140 40.965 ;
        RECT 19.220 40.635 20.800 40.965 ;
        RECT 28.880 40.635 30.460 40.965 ;
        RECT 38.540 40.635 40.120 40.965 ;
        RECT 9.560 35.195 11.140 35.525 ;
        RECT 19.220 35.195 20.800 35.525 ;
        RECT 28.880 35.195 30.460 35.525 ;
        RECT 38.540 35.195 40.120 35.525 ;
        RECT 9.560 29.755 11.140 30.085 ;
        RECT 19.220 29.755 20.800 30.085 ;
        RECT 28.880 29.755 30.460 30.085 ;
        RECT 38.540 29.755 40.120 30.085 ;
        RECT 9.560 24.315 11.140 24.645 ;
        RECT 19.220 24.315 20.800 24.645 ;
        RECT 28.880 24.315 30.460 24.645 ;
        RECT 38.540 24.315 40.120 24.645 ;
        RECT 9.560 18.875 11.140 19.205 ;
        RECT 19.220 18.875 20.800 19.205 ;
        RECT 28.880 18.875 30.460 19.205 ;
        RECT 38.540 18.875 40.120 19.205 ;
        RECT 9.560 13.435 11.140 13.765 ;
        RECT 19.220 13.435 20.800 13.765 ;
        RECT 28.880 13.435 30.460 13.765 ;
        RECT 38.540 13.435 40.120 13.765 ;
      LAYER met4 ;
        RECT 9.550 10.640 11.150 98.160 ;
        RECT 19.210 10.640 20.810 98.160 ;
        RECT 28.870 10.640 30.470 98.160 ;
        RECT 38.530 10.640 40.130 98.160 ;
    END
  END vccd1
  PIN vssd1
    ANTENNAGATEAREA 776.962158 ;
    ANTENNADIFFAREA 93.163246 ;
    PORT
      LAYER pwell ;
        RECT 18.415 96.945 18.845 97.730 ;
        RECT 31.295 96.945 31.725 97.730 ;
        RECT 18.415 92.670 18.845 93.455 ;
        RECT 31.295 91.505 31.725 92.290 ;
        RECT 18.415 87.230 18.845 88.015 ;
        RECT 31.295 86.065 31.725 86.850 ;
        RECT 18.415 81.790 18.845 82.575 ;
        RECT 31.295 80.625 31.725 81.410 ;
        RECT 18.415 76.350 18.845 77.135 ;
        RECT 31.295 75.185 31.725 75.970 ;
        RECT 18.415 70.910 18.845 71.695 ;
        RECT 31.295 69.745 31.725 70.530 ;
        RECT 18.415 65.470 18.845 66.255 ;
        RECT 31.295 64.305 31.725 65.090 ;
        RECT 18.415 60.030 18.845 60.815 ;
        RECT 31.295 58.865 31.725 59.650 ;
        RECT 18.415 54.590 18.845 55.375 ;
        RECT 31.295 53.425 31.725 54.210 ;
        RECT 18.415 49.150 18.845 49.935 ;
        RECT 31.295 47.985 31.725 48.770 ;
        RECT 18.415 43.710 18.845 44.495 ;
        RECT 31.295 42.545 31.725 43.330 ;
        RECT 18.415 38.270 18.845 39.055 ;
        RECT 31.295 37.105 31.725 37.890 ;
        RECT 18.415 32.830 18.845 33.615 ;
        RECT 31.295 31.665 31.725 32.450 ;
        RECT 18.415 27.390 18.845 28.175 ;
        RECT 31.295 26.225 31.725 27.010 ;
        RECT 18.415 21.950 18.845 22.735 ;
        RECT 31.295 20.785 31.725 21.570 ;
        RECT 18.415 16.510 18.845 17.295 ;
        RECT 31.295 15.345 31.725 16.130 ;
        RECT 18.415 11.070 18.845 11.855 ;
        RECT 31.295 11.070 31.725 11.855 ;
      LAYER li1 ;
        RECT 5.520 97.835 44.160 98.005 ;
        RECT 5.605 97.085 6.815 97.835 ;
        RECT 7.455 97.355 7.730 97.835 ;
        RECT 8.315 97.435 8.650 97.835 ;
        RECT 9.265 97.455 9.595 97.835 ;
        RECT 10.645 97.455 10.975 97.835 ;
        RECT 11.585 97.290 16.930 97.835 ;
        RECT 5.605 96.545 6.125 97.085 ;
        RECT 13.170 96.460 13.510 97.290 ;
        RECT 17.105 97.085 18.315 97.835 ;
        RECT 18.485 97.110 18.775 97.835 ;
        RECT 19.420 97.455 19.750 97.835 ;
        RECT 17.105 96.545 17.625 97.085 ;
        RECT 20.350 96.995 20.610 97.835 ;
        RECT 20.785 97.290 26.130 97.835 ;
        RECT 22.370 96.460 22.710 97.290 ;
        RECT 26.305 97.065 29.815 97.835 ;
        RECT 29.985 97.085 31.195 97.835 ;
        RECT 31.365 97.110 31.655 97.835 ;
        RECT 31.830 97.435 32.165 97.835 ;
        RECT 32.750 97.355 33.025 97.835 ;
        RECT 33.665 97.290 39.010 97.835 ;
        RECT 26.305 96.545 27.955 97.065 ;
        RECT 29.985 96.545 30.505 97.085 ;
        RECT 35.250 96.460 35.590 97.290 ;
        RECT 39.185 97.065 40.855 97.835 ;
        RECT 41.925 97.455 42.255 97.835 ;
        RECT 42.865 97.085 44.075 97.835 ;
        RECT 39.185 96.545 39.935 97.065 ;
        RECT 43.555 96.545 44.075 97.085 ;
        RECT 5.605 93.315 6.125 93.855 ;
        RECT 5.605 92.565 6.815 93.315 ;
        RECT 9.950 93.110 10.290 93.940 ;
        RECT 13.885 93.335 15.535 93.855 ;
        RECT 7.425 92.565 7.755 92.945 ;
        RECT 8.365 92.565 13.710 93.110 ;
        RECT 13.885 92.565 17.395 93.335 ;
        RECT 18.485 92.565 18.775 93.290 ;
        RECT 20.530 93.110 20.870 93.940 ;
        RECT 26.050 93.110 26.390 93.940 ;
        RECT 31.570 93.110 31.910 93.940 ;
        RECT 37.090 93.110 37.430 93.940 ;
        RECT 41.025 93.335 41.775 93.855 ;
        RECT 18.945 92.565 24.290 93.110 ;
        RECT 24.465 92.565 29.810 93.110 ;
        RECT 29.985 92.565 35.330 93.110 ;
        RECT 35.505 92.565 40.850 93.110 ;
        RECT 41.025 92.565 42.695 93.335 ;
        RECT 43.555 93.315 44.075 93.855 ;
        RECT 42.865 92.565 44.075 93.315 ;
        RECT 5.520 92.395 44.160 92.565 ;
        RECT 5.605 91.645 6.815 92.395 ;
        RECT 6.985 91.850 12.330 92.395 ;
        RECT 12.505 91.850 17.850 92.395 ;
        RECT 18.025 91.850 23.370 92.395 ;
        RECT 23.545 91.850 28.890 92.395 ;
        RECT 5.605 91.105 6.125 91.645 ;
        RECT 8.570 91.020 8.910 91.850 ;
        RECT 14.090 91.020 14.430 91.850 ;
        RECT 19.610 91.020 19.950 91.850 ;
        RECT 25.130 91.020 25.470 91.850 ;
        RECT 29.065 91.625 30.735 92.395 ;
        RECT 31.365 91.670 31.655 92.395 ;
        RECT 31.825 91.850 37.170 92.395 ;
        RECT 37.345 91.850 42.690 92.395 ;
        RECT 29.065 91.105 29.815 91.625 ;
        RECT 33.410 91.020 33.750 91.850 ;
        RECT 38.930 91.020 39.270 91.850 ;
        RECT 42.865 91.645 44.075 92.395 ;
        RECT 43.555 91.105 44.075 91.645 ;
        RECT 5.605 87.875 6.125 88.415 ;
        RECT 5.605 87.125 6.815 87.875 ;
        RECT 8.570 87.670 8.910 88.500 ;
        RECT 14.090 87.670 14.430 88.500 ;
        RECT 6.985 87.125 12.330 87.670 ;
        RECT 12.505 87.125 17.850 87.670 ;
        RECT 18.485 87.125 18.775 87.850 ;
        RECT 20.530 87.670 20.870 88.500 ;
        RECT 26.050 87.670 26.390 88.500 ;
        RECT 31.570 87.670 31.910 88.500 ;
        RECT 37.090 87.670 37.430 88.500 ;
        RECT 41.025 87.895 41.775 88.415 ;
        RECT 18.945 87.125 24.290 87.670 ;
        RECT 24.465 87.125 29.810 87.670 ;
        RECT 29.985 87.125 35.330 87.670 ;
        RECT 35.505 87.125 40.850 87.670 ;
        RECT 41.025 87.125 42.695 87.895 ;
        RECT 43.555 87.875 44.075 88.415 ;
        RECT 42.865 87.125 44.075 87.875 ;
        RECT 5.520 86.955 44.160 87.125 ;
        RECT 5.605 86.205 6.815 86.955 ;
        RECT 7.425 86.575 7.755 86.955 ;
        RECT 8.365 86.410 13.710 86.955 ;
        RECT 13.885 86.410 19.230 86.955 ;
        RECT 19.405 86.410 24.750 86.955 ;
        RECT 24.925 86.410 30.270 86.955 ;
        RECT 5.605 85.665 6.125 86.205 ;
        RECT 9.950 85.580 10.290 86.410 ;
        RECT 15.470 85.580 15.810 86.410 ;
        RECT 20.990 85.580 21.330 86.410 ;
        RECT 26.510 85.580 26.850 86.410 ;
        RECT 31.365 86.230 31.655 86.955 ;
        RECT 31.825 86.410 37.170 86.955 ;
        RECT 37.345 86.410 42.690 86.955 ;
        RECT 33.410 85.580 33.750 86.410 ;
        RECT 38.930 85.580 39.270 86.410 ;
        RECT 42.865 86.205 44.075 86.955 ;
        RECT 43.555 85.665 44.075 86.205 ;
        RECT 5.605 82.435 6.125 82.975 ;
        RECT 5.605 81.685 6.815 82.435 ;
        RECT 8.570 82.230 8.910 83.060 ;
        RECT 14.090 82.230 14.430 83.060 ;
        RECT 6.985 81.685 12.330 82.230 ;
        RECT 12.505 81.685 17.850 82.230 ;
        RECT 18.485 81.685 18.775 82.410 ;
        RECT 20.530 82.230 20.870 83.060 ;
        RECT 26.050 82.230 26.390 83.060 ;
        RECT 31.570 82.230 31.910 83.060 ;
        RECT 37.090 82.230 37.430 83.060 ;
        RECT 41.025 82.455 41.775 82.975 ;
        RECT 18.945 81.685 24.290 82.230 ;
        RECT 24.465 81.685 29.810 82.230 ;
        RECT 29.985 81.685 35.330 82.230 ;
        RECT 35.505 81.685 40.850 82.230 ;
        RECT 41.025 81.685 42.695 82.455 ;
        RECT 43.555 82.435 44.075 82.975 ;
        RECT 42.865 81.685 44.075 82.435 ;
        RECT 5.520 81.515 44.160 81.685 ;
        RECT 5.605 80.765 6.815 81.515 ;
        RECT 7.415 81.135 7.745 81.515 ;
        RECT 9.700 80.795 9.990 81.515 ;
        RECT 12.050 81.055 12.220 81.515 ;
        RECT 12.910 81.135 13.240 81.515 ;
        RECT 15.795 81.055 15.965 81.515 ;
        RECT 16.645 80.970 21.990 81.515 ;
        RECT 22.165 80.970 27.510 81.515 ;
        RECT 5.605 80.225 6.125 80.765 ;
        RECT 18.230 80.140 18.570 80.970 ;
        RECT 23.750 80.140 24.090 80.970 ;
        RECT 27.685 80.745 31.195 81.515 ;
        RECT 31.365 80.790 31.655 81.515 ;
        RECT 31.825 80.970 37.170 81.515 ;
        RECT 37.345 80.970 42.690 81.515 ;
        RECT 27.685 80.225 29.335 80.745 ;
        RECT 33.410 80.140 33.750 80.970 ;
        RECT 38.930 80.140 39.270 80.970 ;
        RECT 42.865 80.765 44.075 81.515 ;
        RECT 43.555 80.225 44.075 80.765 ;
        RECT 5.605 76.995 6.125 77.535 ;
        RECT 5.605 76.245 6.815 76.995 ;
        RECT 9.950 76.790 10.290 77.620 ;
        RECT 13.885 77.015 15.535 77.535 ;
        RECT 7.425 76.245 7.755 76.625 ;
        RECT 8.365 76.245 13.710 76.790 ;
        RECT 13.885 76.245 17.395 77.015 ;
        RECT 18.485 76.245 18.775 76.970 ;
        RECT 20.530 76.790 20.870 77.620 ;
        RECT 26.050 76.790 26.390 77.620 ;
        RECT 31.570 76.790 31.910 77.620 ;
        RECT 37.090 76.790 37.430 77.620 ;
        RECT 41.025 77.015 41.775 77.535 ;
        RECT 18.945 76.245 24.290 76.790 ;
        RECT 24.465 76.245 29.810 76.790 ;
        RECT 29.985 76.245 35.330 76.790 ;
        RECT 35.505 76.245 40.850 76.790 ;
        RECT 41.025 76.245 42.695 77.015 ;
        RECT 43.555 76.995 44.075 77.535 ;
        RECT 42.865 76.245 44.075 76.995 ;
        RECT 5.520 76.075 44.160 76.245 ;
        RECT 5.605 75.325 6.815 76.075 ;
        RECT 7.415 75.695 7.745 76.075 ;
        RECT 9.700 75.355 9.990 76.075 ;
        RECT 12.050 75.615 12.220 76.075 ;
        RECT 12.910 75.695 13.240 76.075 ;
        RECT 15.795 75.615 15.965 76.075 ;
        RECT 16.645 75.530 21.990 76.075 ;
        RECT 22.165 75.530 27.510 76.075 ;
        RECT 5.605 74.785 6.125 75.325 ;
        RECT 18.230 74.700 18.570 75.530 ;
        RECT 23.750 74.700 24.090 75.530 ;
        RECT 27.685 75.305 31.195 76.075 ;
        RECT 31.365 75.350 31.655 76.075 ;
        RECT 31.825 75.530 37.170 76.075 ;
        RECT 37.345 75.530 42.690 76.075 ;
        RECT 27.685 74.785 29.335 75.305 ;
        RECT 33.410 74.700 33.750 75.530 ;
        RECT 38.930 74.700 39.270 75.530 ;
        RECT 42.865 75.325 44.075 76.075 ;
        RECT 43.555 74.785 44.075 75.325 ;
        RECT 5.605 71.555 6.125 72.095 ;
        RECT 8.365 71.575 9.575 72.095 ;
        RECT 15.725 71.575 16.935 72.095 ;
        RECT 5.605 70.805 6.815 71.555 ;
        RECT 7.425 70.805 7.755 71.185 ;
        RECT 8.365 70.805 10.955 71.575 ;
        RECT 12.015 70.805 12.345 71.205 ;
        RECT 14.305 70.805 14.815 71.340 ;
        RECT 15.725 70.805 18.315 71.575 ;
        RECT 18.485 70.805 18.775 71.530 ;
        RECT 20.530 71.350 20.870 72.180 ;
        RECT 26.050 71.350 26.390 72.180 ;
        RECT 31.570 71.350 31.910 72.180 ;
        RECT 37.090 71.350 37.430 72.180 ;
        RECT 41.025 71.575 41.775 72.095 ;
        RECT 18.945 70.805 24.290 71.350 ;
        RECT 24.465 70.805 29.810 71.350 ;
        RECT 29.985 70.805 35.330 71.350 ;
        RECT 35.505 70.805 40.850 71.350 ;
        RECT 41.025 70.805 42.695 71.575 ;
        RECT 43.555 71.555 44.075 72.095 ;
        RECT 42.865 70.805 44.075 71.555 ;
        RECT 5.520 70.635 44.160 70.805 ;
        RECT 5.605 69.885 6.815 70.635 ;
        RECT 6.985 70.090 12.330 70.635 ;
        RECT 12.505 70.090 17.850 70.635 ;
        RECT 18.025 70.090 23.370 70.635 ;
        RECT 23.545 70.090 28.890 70.635 ;
        RECT 5.605 69.345 6.125 69.885 ;
        RECT 8.570 69.260 8.910 70.090 ;
        RECT 14.090 69.260 14.430 70.090 ;
        RECT 19.610 69.260 19.950 70.090 ;
        RECT 25.130 69.260 25.470 70.090 ;
        RECT 29.065 69.865 30.735 70.635 ;
        RECT 31.365 69.910 31.655 70.635 ;
        RECT 31.825 70.090 37.170 70.635 ;
        RECT 37.345 70.090 42.690 70.635 ;
        RECT 29.065 69.345 29.815 69.865 ;
        RECT 33.410 69.260 33.750 70.090 ;
        RECT 38.930 69.260 39.270 70.090 ;
        RECT 42.865 69.885 44.075 70.635 ;
        RECT 43.555 69.345 44.075 69.885 ;
        RECT 5.605 66.115 6.125 66.655 ;
        RECT 5.605 65.365 6.815 66.115 ;
        RECT 9.950 65.910 10.290 66.740 ;
        RECT 13.885 66.135 15.535 66.655 ;
        RECT 7.425 65.365 7.755 65.745 ;
        RECT 8.365 65.365 13.710 65.910 ;
        RECT 13.885 65.365 17.395 66.135 ;
        RECT 18.485 65.365 18.775 66.090 ;
        RECT 20.530 65.910 20.870 66.740 ;
        RECT 26.050 65.910 26.390 66.740 ;
        RECT 31.570 65.910 31.910 66.740 ;
        RECT 37.090 65.910 37.430 66.740 ;
        RECT 41.025 66.135 41.775 66.655 ;
        RECT 18.945 65.365 24.290 65.910 ;
        RECT 24.465 65.365 29.810 65.910 ;
        RECT 29.985 65.365 35.330 65.910 ;
        RECT 35.505 65.365 40.850 65.910 ;
        RECT 41.025 65.365 42.695 66.135 ;
        RECT 43.555 66.115 44.075 66.655 ;
        RECT 42.865 65.365 44.075 66.115 ;
        RECT 5.520 65.195 44.160 65.365 ;
        RECT 5.605 64.445 6.815 65.195 ;
        RECT 6.985 64.650 12.330 65.195 ;
        RECT 12.505 64.650 17.850 65.195 ;
        RECT 18.025 64.650 23.370 65.195 ;
        RECT 23.545 64.650 28.890 65.195 ;
        RECT 5.605 63.905 6.125 64.445 ;
        RECT 8.570 63.820 8.910 64.650 ;
        RECT 14.090 63.820 14.430 64.650 ;
        RECT 19.610 63.820 19.950 64.650 ;
        RECT 25.130 63.820 25.470 64.650 ;
        RECT 29.065 64.425 30.735 65.195 ;
        RECT 31.365 64.470 31.655 65.195 ;
        RECT 31.825 64.650 37.170 65.195 ;
        RECT 37.345 64.650 42.690 65.195 ;
        RECT 29.065 63.905 29.815 64.425 ;
        RECT 33.410 63.820 33.750 64.650 ;
        RECT 38.930 63.820 39.270 64.650 ;
        RECT 42.865 64.445 44.075 65.195 ;
        RECT 43.555 63.905 44.075 64.445 ;
        RECT 5.605 60.675 6.125 61.215 ;
        RECT 6.985 60.695 8.635 61.215 ;
        RECT 5.605 59.925 6.815 60.675 ;
        RECT 6.985 59.925 10.495 60.695 ;
        RECT 11.605 59.925 11.845 60.735 ;
        RECT 12.515 59.925 12.785 60.735 ;
        RECT 14.550 60.470 14.890 61.300 ;
        RECT 12.965 59.925 18.310 60.470 ;
        RECT 18.485 59.925 18.775 60.650 ;
        RECT 20.530 60.470 20.870 61.300 ;
        RECT 26.050 60.470 26.390 61.300 ;
        RECT 31.570 60.470 31.910 61.300 ;
        RECT 37.090 60.470 37.430 61.300 ;
        RECT 41.025 60.695 41.775 61.215 ;
        RECT 18.945 59.925 24.290 60.470 ;
        RECT 24.465 59.925 29.810 60.470 ;
        RECT 29.985 59.925 35.330 60.470 ;
        RECT 35.505 59.925 40.850 60.470 ;
        RECT 41.025 59.925 42.695 60.695 ;
        RECT 43.555 60.675 44.075 61.215 ;
        RECT 42.865 59.925 44.075 60.675 ;
        RECT 5.520 59.755 44.160 59.925 ;
        RECT 5.605 59.005 6.815 59.755 ;
        RECT 7.425 59.375 7.755 59.755 ;
        RECT 5.605 58.465 6.125 59.005 ;
        RECT 8.365 58.985 11.875 59.755 ;
        RECT 12.055 59.015 12.385 59.755 ;
        RECT 13.090 59.395 13.420 59.755 ;
        RECT 8.365 58.465 10.015 58.985 ;
        RECT 14.785 58.975 15.080 59.755 ;
        RECT 15.265 59.210 20.610 59.755 ;
        RECT 20.785 59.210 26.130 59.755 ;
        RECT 16.850 58.380 17.190 59.210 ;
        RECT 22.370 58.380 22.710 59.210 ;
        RECT 26.305 58.985 29.815 59.755 ;
        RECT 29.985 59.005 31.195 59.755 ;
        RECT 31.365 59.030 31.655 59.755 ;
        RECT 31.825 59.210 37.170 59.755 ;
        RECT 37.345 59.210 42.690 59.755 ;
        RECT 26.305 58.465 27.955 58.985 ;
        RECT 29.985 58.465 30.505 59.005 ;
        RECT 33.410 58.380 33.750 59.210 ;
        RECT 38.930 58.380 39.270 59.210 ;
        RECT 42.865 59.005 44.075 59.755 ;
        RECT 43.555 58.465 44.075 59.005 ;
        RECT 5.605 55.235 6.125 55.775 ;
        RECT 5.605 54.485 6.815 55.235 ;
        RECT 8.570 55.030 8.910 55.860 ;
        RECT 14.090 55.030 14.430 55.860 ;
        RECT 6.985 54.485 12.330 55.030 ;
        RECT 12.505 54.485 17.850 55.030 ;
        RECT 18.485 54.485 18.775 55.210 ;
        RECT 20.530 55.030 20.870 55.860 ;
        RECT 26.050 55.030 26.390 55.860 ;
        RECT 31.570 55.030 31.910 55.860 ;
        RECT 18.945 54.485 24.290 55.030 ;
        RECT 24.465 54.485 29.810 55.030 ;
        RECT 29.985 54.485 35.330 55.030 ;
        RECT 35.515 54.485 35.845 54.965 ;
        RECT 36.355 54.485 36.685 54.965 ;
        RECT 37.195 54.485 37.525 54.965 ;
        RECT 38.035 54.485 38.365 54.965 ;
        RECT 38.875 54.485 39.205 54.965 ;
        RECT 39.715 54.485 40.045 54.965 ;
        RECT 40.555 54.485 40.885 54.965 ;
        RECT 41.395 54.485 41.725 54.965 ;
        RECT 42.235 54.485 42.565 55.285 ;
        RECT 43.555 55.235 44.075 55.775 ;
        RECT 42.865 54.485 44.075 55.235 ;
        RECT 5.520 54.315 44.160 54.485 ;
        RECT 5.605 53.565 6.815 54.315 ;
        RECT 7.425 53.935 7.755 54.315 ;
        RECT 8.365 53.770 13.710 54.315 ;
        RECT 13.885 53.770 19.230 54.315 ;
        RECT 19.405 53.770 24.750 54.315 ;
        RECT 24.925 53.770 30.270 54.315 ;
        RECT 5.605 53.025 6.125 53.565 ;
        RECT 9.950 52.940 10.290 53.770 ;
        RECT 15.470 52.940 15.810 53.770 ;
        RECT 20.990 52.940 21.330 53.770 ;
        RECT 26.510 52.940 26.850 53.770 ;
        RECT 31.365 53.590 31.655 54.315 ;
        RECT 31.825 53.770 37.170 54.315 ;
        RECT 37.345 53.770 42.690 54.315 ;
        RECT 33.410 52.940 33.750 53.770 ;
        RECT 38.930 52.940 39.270 53.770 ;
        RECT 42.865 53.565 44.075 54.315 ;
        RECT 43.555 53.025 44.075 53.565 ;
        RECT 5.605 49.795 6.125 50.335 ;
        RECT 5.605 49.045 6.815 49.795 ;
        RECT 8.570 49.590 8.910 50.420 ;
        RECT 14.090 49.590 14.430 50.420 ;
        RECT 6.985 49.045 12.330 49.590 ;
        RECT 12.505 49.045 17.850 49.590 ;
        RECT 18.485 49.045 18.775 49.770 ;
        RECT 20.530 49.590 20.870 50.420 ;
        RECT 26.050 49.590 26.390 50.420 ;
        RECT 31.570 49.590 31.910 50.420 ;
        RECT 37.090 49.590 37.430 50.420 ;
        RECT 41.025 49.815 41.775 50.335 ;
        RECT 18.945 49.045 24.290 49.590 ;
        RECT 24.465 49.045 29.810 49.590 ;
        RECT 29.985 49.045 35.330 49.590 ;
        RECT 35.505 49.045 40.850 49.590 ;
        RECT 41.025 49.045 42.695 49.815 ;
        RECT 43.555 49.795 44.075 50.335 ;
        RECT 42.865 49.045 44.075 49.795 ;
        RECT 5.520 48.875 44.160 49.045 ;
        RECT 5.605 48.125 6.815 48.875 ;
        RECT 7.715 48.135 8.045 48.875 ;
        RECT 8.555 48.475 8.885 48.875 ;
        RECT 9.745 48.330 15.090 48.875 ;
        RECT 15.265 48.330 20.610 48.875 ;
        RECT 20.785 48.330 26.130 48.875 ;
        RECT 5.605 47.585 6.125 48.125 ;
        RECT 11.330 47.500 11.670 48.330 ;
        RECT 16.850 47.500 17.190 48.330 ;
        RECT 22.370 47.500 22.710 48.330 ;
        RECT 26.305 48.105 29.815 48.875 ;
        RECT 29.985 48.125 31.195 48.875 ;
        RECT 31.365 48.150 31.655 48.875 ;
        RECT 31.825 48.330 37.170 48.875 ;
        RECT 37.345 48.330 42.690 48.875 ;
        RECT 26.305 47.585 27.955 48.105 ;
        RECT 29.985 47.585 30.505 48.125 ;
        RECT 33.410 47.500 33.750 48.330 ;
        RECT 38.930 47.500 39.270 48.330 ;
        RECT 42.865 48.125 44.075 48.875 ;
        RECT 43.555 47.585 44.075 48.125 ;
        RECT 5.605 44.355 6.125 44.895 ;
        RECT 5.605 43.605 6.815 44.355 ;
        RECT 9.950 44.150 10.290 44.980 ;
        RECT 13.885 44.375 15.535 44.895 ;
        RECT 7.425 43.605 7.755 43.985 ;
        RECT 8.365 43.605 13.710 44.150 ;
        RECT 13.885 43.605 17.395 44.375 ;
        RECT 18.485 43.605 18.775 44.330 ;
        RECT 20.530 44.150 20.870 44.980 ;
        RECT 26.050 44.150 26.390 44.980 ;
        RECT 31.570 44.150 31.910 44.980 ;
        RECT 37.090 44.150 37.430 44.980 ;
        RECT 41.025 44.375 41.775 44.895 ;
        RECT 18.945 43.605 24.290 44.150 ;
        RECT 24.465 43.605 29.810 44.150 ;
        RECT 29.985 43.605 35.330 44.150 ;
        RECT 35.505 43.605 40.850 44.150 ;
        RECT 41.025 43.605 42.695 44.375 ;
        RECT 43.555 44.355 44.075 44.895 ;
        RECT 42.865 43.605 44.075 44.355 ;
        RECT 5.520 43.435 44.160 43.605 ;
        RECT 5.605 42.685 6.815 43.435 ;
        RECT 7.725 42.900 8.235 43.435 ;
        RECT 10.195 43.035 10.525 43.435 ;
        RECT 11.210 42.760 11.450 43.435 ;
        RECT 12.840 42.985 13.170 43.435 ;
        RECT 14.090 42.995 14.405 43.435 ;
        RECT 14.805 42.890 20.150 43.435 ;
        RECT 20.325 42.890 25.670 43.435 ;
        RECT 25.845 42.890 31.190 43.435 ;
        RECT 5.605 42.145 6.125 42.685 ;
        RECT 16.390 42.060 16.730 42.890 ;
        RECT 21.910 42.060 22.250 42.890 ;
        RECT 27.430 42.060 27.770 42.890 ;
        RECT 31.365 42.710 31.655 43.435 ;
        RECT 31.825 42.890 37.170 43.435 ;
        RECT 37.345 42.890 42.690 43.435 ;
        RECT 33.410 42.060 33.750 42.890 ;
        RECT 38.930 42.060 39.270 42.890 ;
        RECT 42.865 42.685 44.075 43.435 ;
        RECT 43.555 42.145 44.075 42.685 ;
        RECT 5.605 38.915 6.125 39.455 ;
        RECT 5.605 38.165 6.815 38.915 ;
        RECT 6.985 38.165 7.245 38.985 ;
        RECT 11.790 38.710 12.130 39.540 ;
        RECT 15.725 38.935 16.935 39.455 ;
        RECT 9.275 38.165 9.605 38.625 ;
        RECT 10.205 38.165 15.550 38.710 ;
        RECT 15.725 38.165 18.315 38.935 ;
        RECT 18.485 38.165 18.775 38.890 ;
        RECT 20.530 38.710 20.870 39.540 ;
        RECT 26.050 38.710 26.390 39.540 ;
        RECT 31.570 38.710 31.910 39.540 ;
        RECT 37.090 38.710 37.430 39.540 ;
        RECT 41.025 38.935 41.775 39.455 ;
        RECT 18.945 38.165 24.290 38.710 ;
        RECT 24.465 38.165 29.810 38.710 ;
        RECT 29.985 38.165 35.330 38.710 ;
        RECT 35.505 38.165 40.850 38.710 ;
        RECT 41.025 38.165 42.695 38.935 ;
        RECT 43.555 38.915 44.075 39.455 ;
        RECT 42.865 38.165 44.075 38.915 ;
        RECT 5.520 37.995 44.160 38.165 ;
        RECT 5.605 37.245 6.815 37.995 ;
        RECT 7.425 37.615 7.755 37.995 ;
        RECT 8.365 37.450 13.710 37.995 ;
        RECT 13.885 37.450 19.230 37.995 ;
        RECT 19.405 37.450 24.750 37.995 ;
        RECT 24.925 37.450 30.270 37.995 ;
        RECT 5.605 36.705 6.125 37.245 ;
        RECT 9.950 36.620 10.290 37.450 ;
        RECT 15.470 36.620 15.810 37.450 ;
        RECT 20.990 36.620 21.330 37.450 ;
        RECT 26.510 36.620 26.850 37.450 ;
        RECT 31.365 37.270 31.655 37.995 ;
        RECT 31.825 37.450 37.170 37.995 ;
        RECT 37.345 37.450 42.690 37.995 ;
        RECT 33.410 36.620 33.750 37.450 ;
        RECT 38.930 36.620 39.270 37.450 ;
        RECT 42.865 37.245 44.075 37.995 ;
        RECT 43.555 36.705 44.075 37.245 ;
        RECT 5.605 33.475 6.125 34.015 ;
        RECT 6.985 33.475 7.505 34.015 ;
        RECT 5.605 32.725 6.815 33.475 ;
        RECT 6.985 32.725 8.195 33.475 ;
        RECT 8.365 32.725 8.705 33.450 ;
        RECT 13.630 33.270 13.970 34.100 ;
        RECT 11.035 32.725 11.365 33.205 ;
        RECT 12.045 32.725 17.390 33.270 ;
        RECT 18.485 32.725 18.775 33.450 ;
        RECT 20.530 33.270 20.870 34.100 ;
        RECT 26.050 33.270 26.390 34.100 ;
        RECT 31.570 33.270 31.910 34.100 ;
        RECT 37.090 33.270 37.430 34.100 ;
        RECT 41.025 33.495 41.775 34.015 ;
        RECT 18.945 32.725 24.290 33.270 ;
        RECT 24.465 32.725 29.810 33.270 ;
        RECT 29.985 32.725 35.330 33.270 ;
        RECT 35.505 32.725 40.850 33.270 ;
        RECT 41.025 32.725 42.695 33.495 ;
        RECT 43.555 33.475 44.075 34.015 ;
        RECT 42.865 32.725 44.075 33.475 ;
        RECT 5.520 32.555 44.160 32.725 ;
        RECT 5.605 31.805 6.815 32.555 ;
        RECT 5.605 31.265 6.125 31.805 ;
        RECT 7.905 31.735 8.165 32.555 ;
        RECT 9.275 32.155 9.605 32.555 ;
        RECT 10.115 32.155 10.490 32.555 ;
        RECT 12.760 32.155 13.090 32.555 ;
        RECT 13.885 32.010 19.230 32.555 ;
        RECT 19.405 32.010 24.750 32.555 ;
        RECT 24.925 32.010 30.270 32.555 ;
        RECT 15.470 31.180 15.810 32.010 ;
        RECT 20.990 31.180 21.330 32.010 ;
        RECT 26.510 31.180 26.850 32.010 ;
        RECT 31.365 31.830 31.655 32.555 ;
        RECT 31.825 32.010 37.170 32.555 ;
        RECT 37.345 32.010 42.690 32.555 ;
        RECT 33.410 31.180 33.750 32.010 ;
        RECT 38.930 31.180 39.270 32.010 ;
        RECT 42.865 31.805 44.075 32.555 ;
        RECT 43.555 31.265 44.075 31.805 ;
        RECT 5.605 28.035 6.125 28.575 ;
        RECT 5.605 27.285 6.815 28.035 ;
        RECT 7.425 27.285 7.755 27.665 ;
        RECT 9.725 27.285 10.035 28.085 ;
        RECT 11.790 27.830 12.130 28.660 ;
        RECT 15.725 28.055 16.935 28.575 ;
        RECT 10.205 27.285 15.550 27.830 ;
        RECT 15.725 27.285 18.315 28.055 ;
        RECT 18.485 27.285 18.775 28.010 ;
        RECT 20.530 27.830 20.870 28.660 ;
        RECT 26.050 27.830 26.390 28.660 ;
        RECT 31.570 27.830 31.910 28.660 ;
        RECT 37.090 27.830 37.430 28.660 ;
        RECT 41.025 28.055 41.775 28.575 ;
        RECT 18.945 27.285 24.290 27.830 ;
        RECT 24.465 27.285 29.810 27.830 ;
        RECT 29.985 27.285 35.330 27.830 ;
        RECT 35.505 27.285 40.850 27.830 ;
        RECT 41.025 27.285 42.695 28.055 ;
        RECT 43.555 28.035 44.075 28.575 ;
        RECT 42.865 27.285 44.075 28.035 ;
        RECT 5.520 27.115 44.160 27.285 ;
        RECT 5.605 26.365 6.815 27.115 ;
        RECT 7.725 26.580 8.235 27.115 ;
        RECT 10.195 26.715 10.525 27.115 ;
        RECT 11.125 26.570 16.470 27.115 ;
        RECT 16.645 26.570 21.990 27.115 ;
        RECT 22.165 26.570 27.510 27.115 ;
        RECT 5.605 25.825 6.125 26.365 ;
        RECT 12.710 25.740 13.050 26.570 ;
        RECT 18.230 25.740 18.570 26.570 ;
        RECT 23.750 25.740 24.090 26.570 ;
        RECT 27.685 26.345 31.195 27.115 ;
        RECT 31.365 26.390 31.655 27.115 ;
        RECT 31.825 26.570 37.170 27.115 ;
        RECT 37.345 26.570 42.690 27.115 ;
        RECT 27.685 25.825 29.335 26.345 ;
        RECT 33.410 25.740 33.750 26.570 ;
        RECT 38.930 25.740 39.270 26.570 ;
        RECT 42.865 26.365 44.075 27.115 ;
        RECT 43.555 25.825 44.075 26.365 ;
        RECT 5.605 22.595 6.125 23.135 ;
        RECT 5.605 21.845 6.815 22.595 ;
        RECT 9.950 22.390 10.290 23.220 ;
        RECT 13.885 22.615 15.535 23.135 ;
        RECT 7.425 21.845 7.755 22.225 ;
        RECT 8.365 21.845 13.710 22.390 ;
        RECT 13.885 21.845 17.395 22.615 ;
        RECT 18.485 21.845 18.775 22.570 ;
        RECT 20.530 22.390 20.870 23.220 ;
        RECT 26.050 22.390 26.390 23.220 ;
        RECT 31.570 22.390 31.910 23.220 ;
        RECT 37.090 22.390 37.430 23.220 ;
        RECT 41.025 22.615 41.775 23.135 ;
        RECT 18.945 21.845 24.290 22.390 ;
        RECT 24.465 21.845 29.810 22.390 ;
        RECT 29.985 21.845 35.330 22.390 ;
        RECT 35.505 21.845 40.850 22.390 ;
        RECT 41.025 21.845 42.695 22.615 ;
        RECT 43.555 22.595 44.075 23.135 ;
        RECT 42.865 21.845 44.075 22.595 ;
        RECT 5.520 21.675 44.160 21.845 ;
        RECT 5.605 20.925 6.815 21.675 ;
        RECT 6.985 21.130 12.330 21.675 ;
        RECT 12.505 21.130 17.850 21.675 ;
        RECT 18.025 21.130 23.370 21.675 ;
        RECT 23.545 21.130 28.890 21.675 ;
        RECT 5.605 20.385 6.125 20.925 ;
        RECT 8.570 20.300 8.910 21.130 ;
        RECT 14.090 20.300 14.430 21.130 ;
        RECT 19.610 20.300 19.950 21.130 ;
        RECT 25.130 20.300 25.470 21.130 ;
        RECT 29.065 20.905 30.735 21.675 ;
        RECT 31.365 20.950 31.655 21.675 ;
        RECT 31.825 21.130 37.170 21.675 ;
        RECT 37.345 21.130 42.690 21.675 ;
        RECT 29.065 20.385 29.815 20.905 ;
        RECT 33.410 20.300 33.750 21.130 ;
        RECT 38.930 20.300 39.270 21.130 ;
        RECT 42.865 20.925 44.075 21.675 ;
        RECT 43.555 20.385 44.075 20.925 ;
        RECT 5.605 17.155 6.125 17.695 ;
        RECT 5.605 16.405 6.815 17.155 ;
        RECT 9.950 16.950 10.290 17.780 ;
        RECT 13.885 17.175 15.535 17.695 ;
        RECT 7.425 16.405 7.755 16.785 ;
        RECT 8.365 16.405 13.710 16.950 ;
        RECT 13.885 16.405 17.395 17.175 ;
        RECT 18.485 16.405 18.775 17.130 ;
        RECT 20.530 16.950 20.870 17.780 ;
        RECT 26.050 16.950 26.390 17.780 ;
        RECT 31.570 16.950 31.910 17.780 ;
        RECT 37.090 16.950 37.430 17.780 ;
        RECT 41.025 17.175 41.775 17.695 ;
        RECT 18.945 16.405 24.290 16.950 ;
        RECT 24.465 16.405 29.810 16.950 ;
        RECT 29.985 16.405 35.330 16.950 ;
        RECT 35.505 16.405 40.850 16.950 ;
        RECT 41.025 16.405 42.695 17.175 ;
        RECT 43.555 17.155 44.075 17.695 ;
        RECT 42.865 16.405 44.075 17.155 ;
        RECT 5.520 16.235 44.160 16.405 ;
        RECT 5.605 15.485 6.815 16.235 ;
        RECT 6.985 15.690 12.330 16.235 ;
        RECT 12.505 15.690 17.850 16.235 ;
        RECT 18.025 15.690 23.370 16.235 ;
        RECT 23.545 15.690 28.890 16.235 ;
        RECT 5.605 14.945 6.125 15.485 ;
        RECT 8.570 14.860 8.910 15.690 ;
        RECT 14.090 14.860 14.430 15.690 ;
        RECT 19.610 14.860 19.950 15.690 ;
        RECT 25.130 14.860 25.470 15.690 ;
        RECT 29.065 15.465 30.735 16.235 ;
        RECT 31.365 15.510 31.655 16.235 ;
        RECT 31.825 15.690 37.170 16.235 ;
        RECT 37.345 15.690 42.690 16.235 ;
        RECT 29.065 14.945 29.815 15.465 ;
        RECT 33.410 14.860 33.750 15.690 ;
        RECT 38.930 14.860 39.270 15.690 ;
        RECT 42.865 15.485 44.075 16.235 ;
        RECT 43.555 14.945 44.075 15.485 ;
        RECT 5.605 11.715 6.125 12.255 ;
        RECT 5.605 10.965 6.815 11.715 ;
        RECT 11.330 11.510 11.670 12.340 ;
        RECT 15.265 11.735 16.475 12.255 ;
        RECT 7.425 10.965 7.755 11.345 ;
        RECT 8.805 10.965 9.135 11.345 ;
        RECT 9.745 10.965 15.090 11.510 ;
        RECT 15.265 10.965 17.855 11.735 ;
        RECT 18.485 10.965 18.775 11.690 ;
        RECT 20.530 11.510 20.870 12.340 ;
        RECT 26.050 11.510 26.390 12.340 ;
        RECT 29.985 11.715 30.505 12.255 ;
        RECT 18.945 10.965 24.290 11.510 ;
        RECT 24.465 10.965 29.810 11.510 ;
        RECT 29.985 10.965 31.195 11.715 ;
        RECT 31.365 10.965 31.655 11.690 ;
        RECT 33.410 11.510 33.750 12.340 ;
        RECT 38.930 11.510 39.270 12.340 ;
        RECT 43.555 11.715 44.075 12.255 ;
        RECT 31.825 10.965 37.170 11.510 ;
        RECT 37.345 10.965 42.690 11.510 ;
        RECT 42.865 10.965 44.075 11.715 ;
        RECT 5.520 10.795 44.160 10.965 ;
      LAYER met1 ;
        RECT 5.520 97.680 44.960 98.160 ;
        RECT 5.520 92.240 44.960 92.720 ;
        RECT 5.520 86.800 44.960 87.280 ;
        RECT 5.520 81.360 44.960 81.840 ;
        RECT 5.520 75.920 44.960 76.400 ;
        RECT 5.520 70.480 44.960 70.960 ;
        RECT 5.520 65.040 44.960 65.520 ;
        RECT 5.520 59.600 44.960 60.080 ;
        RECT 5.520 54.160 44.960 54.640 ;
        RECT 5.520 48.720 44.960 49.200 ;
        RECT 5.520 43.280 44.960 43.760 ;
        RECT 5.520 37.840 44.960 38.320 ;
        RECT 5.520 32.400 44.960 32.880 ;
        RECT 5.520 26.960 44.960 27.440 ;
        RECT 5.520 21.520 44.960 22.000 ;
        RECT 5.520 16.080 44.960 16.560 ;
        RECT 5.520 10.640 44.960 11.120 ;
      LAYER met2 ;
        RECT 14.410 97.735 15.950 98.105 ;
        RECT 24.070 97.735 25.610 98.105 ;
        RECT 33.730 97.735 35.270 98.105 ;
        RECT 43.390 97.735 44.930 98.105 ;
        RECT 14.410 92.295 15.950 92.665 ;
        RECT 24.070 92.295 25.610 92.665 ;
        RECT 33.730 92.295 35.270 92.665 ;
        RECT 43.390 92.295 44.930 92.665 ;
        RECT 14.410 86.855 15.950 87.225 ;
        RECT 24.070 86.855 25.610 87.225 ;
        RECT 33.730 86.855 35.270 87.225 ;
        RECT 43.390 86.855 44.930 87.225 ;
        RECT 14.410 81.415 15.950 81.785 ;
        RECT 24.070 81.415 25.610 81.785 ;
        RECT 33.730 81.415 35.270 81.785 ;
        RECT 43.390 81.415 44.930 81.785 ;
        RECT 14.410 75.975 15.950 76.345 ;
        RECT 24.070 75.975 25.610 76.345 ;
        RECT 33.730 75.975 35.270 76.345 ;
        RECT 43.390 75.975 44.930 76.345 ;
        RECT 14.410 70.535 15.950 70.905 ;
        RECT 24.070 70.535 25.610 70.905 ;
        RECT 33.730 70.535 35.270 70.905 ;
        RECT 43.390 70.535 44.930 70.905 ;
        RECT 14.410 65.095 15.950 65.465 ;
        RECT 24.070 65.095 25.610 65.465 ;
        RECT 33.730 65.095 35.270 65.465 ;
        RECT 43.390 65.095 44.930 65.465 ;
        RECT 14.410 59.655 15.950 60.025 ;
        RECT 24.070 59.655 25.610 60.025 ;
        RECT 33.730 59.655 35.270 60.025 ;
        RECT 43.390 59.655 44.930 60.025 ;
        RECT 14.410 54.215 15.950 54.585 ;
        RECT 24.070 54.215 25.610 54.585 ;
        RECT 33.730 54.215 35.270 54.585 ;
        RECT 43.390 54.215 44.930 54.585 ;
        RECT 14.410 48.775 15.950 49.145 ;
        RECT 24.070 48.775 25.610 49.145 ;
        RECT 33.730 48.775 35.270 49.145 ;
        RECT 43.390 48.775 44.930 49.145 ;
        RECT 14.410 43.335 15.950 43.705 ;
        RECT 24.070 43.335 25.610 43.705 ;
        RECT 33.730 43.335 35.270 43.705 ;
        RECT 43.390 43.335 44.930 43.705 ;
        RECT 14.410 37.895 15.950 38.265 ;
        RECT 24.070 37.895 25.610 38.265 ;
        RECT 33.730 37.895 35.270 38.265 ;
        RECT 43.390 37.895 44.930 38.265 ;
        RECT 14.410 32.455 15.950 32.825 ;
        RECT 24.070 32.455 25.610 32.825 ;
        RECT 33.730 32.455 35.270 32.825 ;
        RECT 43.390 32.455 44.930 32.825 ;
        RECT 14.410 27.015 15.950 27.385 ;
        RECT 24.070 27.015 25.610 27.385 ;
        RECT 33.730 27.015 35.270 27.385 ;
        RECT 43.390 27.015 44.930 27.385 ;
        RECT 14.410 21.575 15.950 21.945 ;
        RECT 24.070 21.575 25.610 21.945 ;
        RECT 33.730 21.575 35.270 21.945 ;
        RECT 43.390 21.575 44.930 21.945 ;
        RECT 14.410 16.135 15.950 16.505 ;
        RECT 24.070 16.135 25.610 16.505 ;
        RECT 33.730 16.135 35.270 16.505 ;
        RECT 43.390 16.135 44.930 16.505 ;
        RECT 14.410 10.695 15.950 11.065 ;
        RECT 24.070 10.695 25.610 11.065 ;
        RECT 33.730 10.695 35.270 11.065 ;
        RECT 43.390 10.695 44.930 11.065 ;
      LAYER met3 ;
        RECT 14.390 97.755 15.970 98.085 ;
        RECT 24.050 97.755 25.630 98.085 ;
        RECT 33.710 97.755 35.290 98.085 ;
        RECT 43.370 97.755 44.950 98.085 ;
        RECT 14.390 92.315 15.970 92.645 ;
        RECT 24.050 92.315 25.630 92.645 ;
        RECT 33.710 92.315 35.290 92.645 ;
        RECT 43.370 92.315 44.950 92.645 ;
        RECT 14.390 86.875 15.970 87.205 ;
        RECT 24.050 86.875 25.630 87.205 ;
        RECT 33.710 86.875 35.290 87.205 ;
        RECT 43.370 86.875 44.950 87.205 ;
        RECT 14.390 81.435 15.970 81.765 ;
        RECT 24.050 81.435 25.630 81.765 ;
        RECT 33.710 81.435 35.290 81.765 ;
        RECT 43.370 81.435 44.950 81.765 ;
        RECT 14.390 75.995 15.970 76.325 ;
        RECT 24.050 75.995 25.630 76.325 ;
        RECT 33.710 75.995 35.290 76.325 ;
        RECT 43.370 75.995 44.950 76.325 ;
        RECT 14.390 70.555 15.970 70.885 ;
        RECT 24.050 70.555 25.630 70.885 ;
        RECT 33.710 70.555 35.290 70.885 ;
        RECT 43.370 70.555 44.950 70.885 ;
        RECT 14.390 65.115 15.970 65.445 ;
        RECT 24.050 65.115 25.630 65.445 ;
        RECT 33.710 65.115 35.290 65.445 ;
        RECT 43.370 65.115 44.950 65.445 ;
        RECT 14.390 59.675 15.970 60.005 ;
        RECT 24.050 59.675 25.630 60.005 ;
        RECT 33.710 59.675 35.290 60.005 ;
        RECT 43.370 59.675 44.950 60.005 ;
        RECT 14.390 54.235 15.970 54.565 ;
        RECT 24.050 54.235 25.630 54.565 ;
        RECT 33.710 54.235 35.290 54.565 ;
        RECT 43.370 54.235 44.950 54.565 ;
        RECT 14.390 48.795 15.970 49.125 ;
        RECT 24.050 48.795 25.630 49.125 ;
        RECT 33.710 48.795 35.290 49.125 ;
        RECT 43.370 48.795 44.950 49.125 ;
        RECT 14.390 43.355 15.970 43.685 ;
        RECT 24.050 43.355 25.630 43.685 ;
        RECT 33.710 43.355 35.290 43.685 ;
        RECT 43.370 43.355 44.950 43.685 ;
        RECT 14.390 37.915 15.970 38.245 ;
        RECT 24.050 37.915 25.630 38.245 ;
        RECT 33.710 37.915 35.290 38.245 ;
        RECT 43.370 37.915 44.950 38.245 ;
        RECT 14.390 32.475 15.970 32.805 ;
        RECT 24.050 32.475 25.630 32.805 ;
        RECT 33.710 32.475 35.290 32.805 ;
        RECT 43.370 32.475 44.950 32.805 ;
        RECT 14.390 27.035 15.970 27.365 ;
        RECT 24.050 27.035 25.630 27.365 ;
        RECT 33.710 27.035 35.290 27.365 ;
        RECT 43.370 27.035 44.950 27.365 ;
        RECT 14.390 21.595 15.970 21.925 ;
        RECT 24.050 21.595 25.630 21.925 ;
        RECT 33.710 21.595 35.290 21.925 ;
        RECT 43.370 21.595 44.950 21.925 ;
        RECT 14.390 16.155 15.970 16.485 ;
        RECT 24.050 16.155 25.630 16.485 ;
        RECT 33.710 16.155 35.290 16.485 ;
        RECT 43.370 16.155 44.950 16.485 ;
        RECT 14.390 10.715 15.970 11.045 ;
        RECT 24.050 10.715 25.630 11.045 ;
        RECT 33.710 10.715 35.290 11.045 ;
        RECT 43.370 10.715 44.950 11.045 ;
      LAYER met4 ;
        RECT 14.380 10.640 15.980 98.160 ;
        RECT 24.040 10.640 25.640 98.160 ;
        RECT 33.700 10.640 35.300 98.160 ;
        RECT 43.360 10.640 44.960 98.160 ;
    END
  END vssd1
  PIN y
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER li1 ;
        RECT 37.695 56.015 37.865 56.865 ;
        RECT 38.535 56.015 38.705 56.865 ;
        RECT 39.375 56.015 39.545 56.865 ;
        RECT 40.215 56.015 40.385 56.865 ;
        RECT 41.055 56.015 41.225 56.865 ;
        RECT 41.895 56.015 42.065 56.865 ;
        RECT 37.695 55.845 42.065 56.015 ;
        RECT 40.130 55.305 42.065 55.845 ;
        RECT 37.695 55.135 42.065 55.305 ;
        RECT 37.695 54.655 37.865 55.135 ;
        RECT 38.535 54.655 38.705 55.135 ;
        RECT 39.375 54.655 39.545 55.135 ;
        RECT 40.215 54.655 40.385 55.135 ;
        RECT 41.055 54.655 41.225 55.135 ;
        RECT 41.895 54.655 42.065 55.135 ;
      LAYER met1 ;
        RECT 41.010 55.120 41.330 55.380 ;
      LAYER met2 ;
        RECT 41.040 55.090 41.300 55.410 ;
        RECT 41.100 53.565 41.240 55.090 ;
        RECT 41.030 53.195 41.310 53.565 ;
      LAYER met3 ;
        RECT 46.000 54.890 50.000 55.040 ;
        RECT 45.390 54.590 50.000 54.890 ;
        RECT 41.005 53.530 41.335 53.545 ;
        RECT 45.390 53.530 45.690 54.590 ;
        RECT 46.000 54.440 50.000 54.590 ;
        RECT 41.005 53.230 45.690 53.530 ;
        RECT 41.005 53.215 41.335 53.230 ;
    END
  END y
  OBS
      LAYER pwell ;
        RECT 5.665 97.815 5.835 98.005 ;
        RECT 7.045 97.815 7.215 98.005 ;
        RECT 9.805 97.815 9.975 98.005 ;
        RECT 11.185 97.815 11.355 98.005 ;
        RECT 11.645 97.815 11.815 98.005 ;
        RECT 17.165 97.815 17.335 98.005 ;
        RECT 19.005 97.815 19.175 98.005 ;
        RECT 20.845 97.815 21.015 98.005 ;
        RECT 26.365 97.815 26.535 98.005 ;
        RECT 30.045 97.815 30.215 98.005 ;
        RECT 33.265 97.815 33.435 98.005 ;
        RECT 33.725 97.815 33.895 98.005 ;
        RECT 39.245 97.815 39.415 98.005 ;
        RECT 41.080 97.865 41.200 97.975 ;
        RECT 42.455 97.815 42.625 98.005 ;
        RECT 43.845 97.815 44.015 98.005 ;
        RECT 5.525 97.005 6.895 97.815 ;
        RECT 6.905 97.135 8.735 97.815 ;
        RECT 8.745 97.035 10.115 97.815 ;
        RECT 10.125 97.035 11.495 97.815 ;
        RECT 11.505 97.005 17.015 97.815 ;
        RECT 17.025 97.005 18.395 97.815 ;
        RECT 18.865 97.135 20.695 97.815 ;
        RECT 19.350 96.905 20.695 97.135 ;
        RECT 20.705 97.005 26.215 97.815 ;
        RECT 26.225 97.005 29.895 97.815 ;
        RECT 29.905 97.005 31.275 97.815 ;
        RECT 31.745 97.135 33.575 97.815 ;
        RECT 33.585 97.005 39.095 97.815 ;
        RECT 39.105 97.005 40.935 97.815 ;
        RECT 41.405 97.035 42.775 97.815 ;
        RECT 42.785 97.005 44.155 97.815 ;
        RECT 5.525 92.585 6.895 93.395 ;
        RECT 6.905 92.585 8.275 93.365 ;
        RECT 8.285 92.585 13.795 93.395 ;
        RECT 13.805 92.585 17.475 93.395 ;
        RECT 18.865 92.585 24.375 93.395 ;
        RECT 24.385 92.585 29.895 93.395 ;
        RECT 29.905 92.585 35.415 93.395 ;
        RECT 35.425 92.585 40.935 93.395 ;
        RECT 40.945 92.585 42.775 93.395 ;
        RECT 42.785 92.585 44.155 93.395 ;
        RECT 5.665 92.375 5.835 92.585 ;
        RECT 7.045 92.375 7.215 92.585 ;
        RECT 8.425 92.395 8.595 92.585 ;
        RECT 12.565 92.375 12.735 92.565 ;
        RECT 13.945 92.395 14.115 92.585 ;
        RECT 17.635 92.430 17.795 92.540 ;
        RECT 18.085 92.375 18.255 92.565 ;
        RECT 19.005 92.395 19.175 92.585 ;
        RECT 23.605 92.375 23.775 92.565 ;
        RECT 24.525 92.395 24.695 92.585 ;
        RECT 29.125 92.375 29.295 92.565 ;
        RECT 30.045 92.395 30.215 92.585 ;
        RECT 30.960 92.425 31.080 92.535 ;
        RECT 31.885 92.375 32.055 92.565 ;
        RECT 35.565 92.395 35.735 92.585 ;
        RECT 37.405 92.375 37.575 92.565 ;
        RECT 41.085 92.395 41.255 92.585 ;
        RECT 43.845 92.375 44.015 92.585 ;
        RECT 5.525 91.565 6.895 92.375 ;
        RECT 6.905 91.565 12.415 92.375 ;
        RECT 12.425 91.565 17.935 92.375 ;
        RECT 17.945 91.565 23.455 92.375 ;
        RECT 23.465 91.565 28.975 92.375 ;
        RECT 28.985 91.565 30.815 92.375 ;
        RECT 31.745 91.565 37.255 92.375 ;
        RECT 37.265 91.565 42.775 92.375 ;
        RECT 42.785 91.565 44.155 92.375 ;
        RECT 5.525 87.145 6.895 87.955 ;
        RECT 6.905 87.145 12.415 87.955 ;
        RECT 12.425 87.145 17.935 87.955 ;
        RECT 18.865 87.145 24.375 87.955 ;
        RECT 24.385 87.145 29.895 87.955 ;
        RECT 29.905 87.145 35.415 87.955 ;
        RECT 35.425 87.145 40.935 87.955 ;
        RECT 40.945 87.145 42.775 87.955 ;
        RECT 42.785 87.145 44.155 87.955 ;
        RECT 5.665 86.935 5.835 87.145 ;
        RECT 7.045 86.935 7.215 87.145 ;
        RECT 8.425 86.935 8.595 87.125 ;
        RECT 12.565 86.955 12.735 87.145 ;
        RECT 13.945 86.935 14.115 87.125 ;
        RECT 18.080 86.985 18.200 87.095 ;
        RECT 19.005 86.955 19.175 87.145 ;
        RECT 19.465 86.935 19.635 87.125 ;
        RECT 24.525 86.955 24.695 87.145 ;
        RECT 24.985 86.935 25.155 87.125 ;
        RECT 30.045 86.955 30.215 87.145 ;
        RECT 30.515 86.980 30.675 87.090 ;
        RECT 31.885 86.935 32.055 87.125 ;
        RECT 35.565 86.955 35.735 87.145 ;
        RECT 37.405 86.935 37.575 87.125 ;
        RECT 41.085 86.955 41.255 87.145 ;
        RECT 43.845 86.935 44.015 87.145 ;
        RECT 5.525 86.125 6.895 86.935 ;
        RECT 6.905 86.155 8.275 86.935 ;
        RECT 8.285 86.125 13.795 86.935 ;
        RECT 13.805 86.125 19.315 86.935 ;
        RECT 19.325 86.125 24.835 86.935 ;
        RECT 24.845 86.125 30.355 86.935 ;
        RECT 31.745 86.125 37.255 86.935 ;
        RECT 37.265 86.125 42.775 86.935 ;
        RECT 42.785 86.125 44.155 86.935 ;
        RECT 5.525 81.705 6.895 82.515 ;
        RECT 6.905 81.705 12.415 82.515 ;
        RECT 12.425 81.705 17.935 82.515 ;
        RECT 18.865 81.705 24.375 82.515 ;
        RECT 24.385 81.705 29.895 82.515 ;
        RECT 29.905 81.705 35.415 82.515 ;
        RECT 35.425 81.705 40.935 82.515 ;
        RECT 40.945 81.705 42.775 82.515 ;
        RECT 42.785 81.705 44.155 82.515 ;
        RECT 5.665 81.495 5.835 81.705 ;
        RECT 7.045 81.495 7.215 81.705 ;
        RECT 12.565 81.515 12.735 81.705 ;
        RECT 16.705 81.495 16.875 81.685 ;
        RECT 18.080 81.545 18.200 81.655 ;
        RECT 19.005 81.515 19.175 81.705 ;
        RECT 22.225 81.495 22.395 81.685 ;
        RECT 24.525 81.515 24.695 81.705 ;
        RECT 27.745 81.495 27.915 81.685 ;
        RECT 30.045 81.515 30.215 81.705 ;
        RECT 31.885 81.495 32.055 81.685 ;
        RECT 35.565 81.515 35.735 81.705 ;
        RECT 37.405 81.495 37.575 81.685 ;
        RECT 41.085 81.515 41.255 81.705 ;
        RECT 43.845 81.495 44.015 81.705 ;
        RECT 5.525 80.685 6.895 81.495 ;
        RECT 6.905 81.325 8.665 81.495 ;
        RECT 6.905 81.280 9.160 81.325 ;
        RECT 6.905 81.245 10.100 81.280 ;
        RECT 11.460 81.245 16.555 81.495 ;
        RECT 6.905 80.815 16.555 81.245 ;
        RECT 8.230 80.645 11.460 80.815 ;
        RECT 9.170 80.600 11.460 80.645 ;
        RECT 10.110 80.565 11.460 80.600 ;
        RECT 14.535 80.585 16.555 80.815 ;
        RECT 16.565 80.685 22.075 81.495 ;
        RECT 22.085 80.685 27.595 81.495 ;
        RECT 27.605 80.685 31.275 81.495 ;
        RECT 31.745 80.685 37.255 81.495 ;
        RECT 37.265 80.685 42.775 81.495 ;
        RECT 42.785 80.685 44.155 81.495 ;
        RECT 14.535 80.565 15.455 80.585 ;
        RECT 5.525 76.265 6.895 77.075 ;
        RECT 6.905 76.265 8.275 77.045 ;
        RECT 8.285 76.265 13.795 77.075 ;
        RECT 13.805 76.265 17.475 77.075 ;
        RECT 18.865 76.265 24.375 77.075 ;
        RECT 24.385 76.265 29.895 77.075 ;
        RECT 29.905 76.265 35.415 77.075 ;
        RECT 35.425 76.265 40.935 77.075 ;
        RECT 40.945 76.265 42.775 77.075 ;
        RECT 42.785 76.265 44.155 77.075 ;
        RECT 5.665 76.055 5.835 76.265 ;
        RECT 7.045 76.055 7.215 76.265 ;
        RECT 8.425 76.075 8.595 76.265 ;
        RECT 13.945 76.075 14.115 76.265 ;
        RECT 16.705 76.055 16.875 76.245 ;
        RECT 17.635 76.110 17.795 76.220 ;
        RECT 19.005 76.075 19.175 76.265 ;
        RECT 22.225 76.055 22.395 76.245 ;
        RECT 24.525 76.075 24.695 76.265 ;
        RECT 27.745 76.055 27.915 76.245 ;
        RECT 30.045 76.075 30.215 76.265 ;
        RECT 31.885 76.055 32.055 76.245 ;
        RECT 35.565 76.075 35.735 76.265 ;
        RECT 37.405 76.055 37.575 76.245 ;
        RECT 41.085 76.075 41.255 76.265 ;
        RECT 43.845 76.055 44.015 76.265 ;
        RECT 5.525 75.245 6.895 76.055 ;
        RECT 6.905 75.885 8.665 76.055 ;
        RECT 6.905 75.840 9.160 75.885 ;
        RECT 6.905 75.805 10.100 75.840 ;
        RECT 11.460 75.805 16.555 76.055 ;
        RECT 6.905 75.375 16.555 75.805 ;
        RECT 8.230 75.205 11.460 75.375 ;
        RECT 9.170 75.160 11.460 75.205 ;
        RECT 10.110 75.125 11.460 75.160 ;
        RECT 14.535 75.145 16.555 75.375 ;
        RECT 16.565 75.245 22.075 76.055 ;
        RECT 22.085 75.245 27.595 76.055 ;
        RECT 27.605 75.245 31.275 76.055 ;
        RECT 31.745 75.245 37.255 76.055 ;
        RECT 37.265 75.245 42.775 76.055 ;
        RECT 42.785 75.245 44.155 76.055 ;
        RECT 14.535 75.125 15.455 75.145 ;
        RECT 5.525 70.825 6.895 71.635 ;
        RECT 6.905 70.825 8.275 71.605 ;
        RECT 8.285 70.825 11.035 71.635 ;
        RECT 11.505 71.505 12.435 71.735 ;
        RECT 11.505 70.825 15.405 71.505 ;
        RECT 15.645 70.825 18.395 71.635 ;
        RECT 18.865 70.825 24.375 71.635 ;
        RECT 24.385 70.825 29.895 71.635 ;
        RECT 29.905 70.825 35.415 71.635 ;
        RECT 35.425 70.825 40.935 71.635 ;
        RECT 40.945 70.825 42.775 71.635 ;
        RECT 42.785 70.825 44.155 71.635 ;
        RECT 5.665 70.615 5.835 70.825 ;
        RECT 7.045 70.615 7.215 70.825 ;
        RECT 8.425 70.635 8.595 70.825 ;
        RECT 11.180 70.665 11.300 70.775 ;
        RECT 11.920 70.635 12.090 70.825 ;
        RECT 12.565 70.615 12.735 70.805 ;
        RECT 15.785 70.635 15.955 70.825 ;
        RECT 18.085 70.615 18.255 70.805 ;
        RECT 19.005 70.635 19.175 70.825 ;
        RECT 23.605 70.615 23.775 70.805 ;
        RECT 24.525 70.635 24.695 70.825 ;
        RECT 29.125 70.615 29.295 70.805 ;
        RECT 30.045 70.635 30.215 70.825 ;
        RECT 30.960 70.665 31.080 70.775 ;
        RECT 31.885 70.615 32.055 70.805 ;
        RECT 35.565 70.635 35.735 70.825 ;
        RECT 37.405 70.615 37.575 70.805 ;
        RECT 41.085 70.635 41.255 70.825 ;
        RECT 43.845 70.615 44.015 70.825 ;
        RECT 5.525 69.805 6.895 70.615 ;
        RECT 6.905 69.805 12.415 70.615 ;
        RECT 12.425 69.805 17.935 70.615 ;
        RECT 17.945 69.805 23.455 70.615 ;
        RECT 23.465 69.805 28.975 70.615 ;
        RECT 28.985 69.805 30.815 70.615 ;
        RECT 31.745 69.805 37.255 70.615 ;
        RECT 37.265 69.805 42.775 70.615 ;
        RECT 42.785 69.805 44.155 70.615 ;
        RECT 5.525 65.385 6.895 66.195 ;
        RECT 6.905 65.385 8.275 66.165 ;
        RECT 8.285 65.385 13.795 66.195 ;
        RECT 13.805 65.385 17.475 66.195 ;
        RECT 18.865 65.385 24.375 66.195 ;
        RECT 24.385 65.385 29.895 66.195 ;
        RECT 29.905 65.385 35.415 66.195 ;
        RECT 35.425 65.385 40.935 66.195 ;
        RECT 40.945 65.385 42.775 66.195 ;
        RECT 42.785 65.385 44.155 66.195 ;
        RECT 5.665 65.175 5.835 65.385 ;
        RECT 7.045 65.175 7.215 65.385 ;
        RECT 8.425 65.195 8.595 65.385 ;
        RECT 12.565 65.175 12.735 65.365 ;
        RECT 13.945 65.195 14.115 65.385 ;
        RECT 17.635 65.230 17.795 65.340 ;
        RECT 18.085 65.175 18.255 65.365 ;
        RECT 19.005 65.195 19.175 65.385 ;
        RECT 23.605 65.175 23.775 65.365 ;
        RECT 24.525 65.195 24.695 65.385 ;
        RECT 29.125 65.175 29.295 65.365 ;
        RECT 30.045 65.195 30.215 65.385 ;
        RECT 30.960 65.225 31.080 65.335 ;
        RECT 31.885 65.175 32.055 65.365 ;
        RECT 35.565 65.195 35.735 65.385 ;
        RECT 37.405 65.175 37.575 65.365 ;
        RECT 41.085 65.195 41.255 65.385 ;
        RECT 43.845 65.175 44.015 65.385 ;
        RECT 5.525 64.365 6.895 65.175 ;
        RECT 6.905 64.365 12.415 65.175 ;
        RECT 12.425 64.365 17.935 65.175 ;
        RECT 17.945 64.365 23.455 65.175 ;
        RECT 23.465 64.365 28.975 65.175 ;
        RECT 28.985 64.365 30.815 65.175 ;
        RECT 31.745 64.365 37.255 65.175 ;
        RECT 37.265 64.365 42.775 65.175 ;
        RECT 42.785 64.365 44.155 65.175 ;
        RECT 5.525 59.945 6.895 60.755 ;
        RECT 6.905 59.945 10.575 60.755 ;
        RECT 11.505 59.945 12.855 60.855 ;
        RECT 12.885 59.945 18.395 60.755 ;
        RECT 18.865 59.945 24.375 60.755 ;
        RECT 24.385 59.945 29.895 60.755 ;
        RECT 29.905 59.945 35.415 60.755 ;
        RECT 35.425 59.945 40.935 60.755 ;
        RECT 40.945 59.945 42.775 60.755 ;
        RECT 42.785 59.945 44.155 60.755 ;
        RECT 5.665 59.735 5.835 59.945 ;
        RECT 7.045 59.735 7.215 59.945 ;
        RECT 8.425 59.735 8.595 59.925 ;
        RECT 10.735 59.790 10.895 59.900 ;
        RECT 11.650 59.755 11.820 59.945 ;
        RECT 13.025 59.755 13.195 59.945 ;
        RECT 14.865 59.735 15.035 59.925 ;
        RECT 15.325 59.735 15.495 59.925 ;
        RECT 19.005 59.755 19.175 59.945 ;
        RECT 20.845 59.735 21.015 59.925 ;
        RECT 24.525 59.755 24.695 59.945 ;
        RECT 26.365 59.735 26.535 59.925 ;
        RECT 30.045 59.735 30.215 59.945 ;
        RECT 31.885 59.735 32.055 59.925 ;
        RECT 35.565 59.755 35.735 59.945 ;
        RECT 37.405 59.735 37.575 59.925 ;
        RECT 41.085 59.755 41.255 59.945 ;
        RECT 43.845 59.735 44.015 59.945 ;
        RECT 5.525 58.925 6.895 59.735 ;
        RECT 6.905 58.955 8.275 59.735 ;
        RECT 8.285 58.925 11.955 59.735 ;
        RECT 11.965 58.825 15.175 59.735 ;
        RECT 15.185 58.925 20.695 59.735 ;
        RECT 20.705 58.925 26.215 59.735 ;
        RECT 26.225 58.925 29.895 59.735 ;
        RECT 29.905 58.925 31.275 59.735 ;
        RECT 31.745 58.925 37.255 59.735 ;
        RECT 37.265 58.925 42.775 59.735 ;
        RECT 42.785 58.925 44.155 59.735 ;
        RECT 5.525 54.505 6.895 55.315 ;
        RECT 6.905 54.505 12.415 55.315 ;
        RECT 12.425 54.505 17.935 55.315 ;
        RECT 18.865 54.505 24.375 55.315 ;
        RECT 24.385 54.505 29.895 55.315 ;
        RECT 29.905 54.505 35.415 55.315 ;
        RECT 35.425 54.505 42.775 55.415 ;
        RECT 42.785 54.505 44.155 55.315 ;
        RECT 5.665 54.295 5.835 54.505 ;
        RECT 7.045 54.295 7.215 54.505 ;
        RECT 8.425 54.295 8.595 54.485 ;
        RECT 12.565 54.315 12.735 54.505 ;
        RECT 13.945 54.295 14.115 54.485 ;
        RECT 18.080 54.345 18.200 54.455 ;
        RECT 19.005 54.315 19.175 54.505 ;
        RECT 19.465 54.295 19.635 54.485 ;
        RECT 24.525 54.315 24.695 54.505 ;
        RECT 24.985 54.295 25.155 54.485 ;
        RECT 30.045 54.315 30.215 54.505 ;
        RECT 30.515 54.340 30.675 54.450 ;
        RECT 31.885 54.295 32.055 54.485 ;
        RECT 35.990 54.315 36.160 54.505 ;
        RECT 37.405 54.295 37.575 54.485 ;
        RECT 43.845 54.295 44.015 54.505 ;
        RECT 5.525 53.485 6.895 54.295 ;
        RECT 6.905 53.515 8.275 54.295 ;
        RECT 8.285 53.485 13.795 54.295 ;
        RECT 13.805 53.485 19.315 54.295 ;
        RECT 19.325 53.485 24.835 54.295 ;
        RECT 24.845 53.485 30.355 54.295 ;
        RECT 31.745 53.485 37.255 54.295 ;
        RECT 37.265 53.485 42.775 54.295 ;
        RECT 42.785 53.485 44.155 54.295 ;
        RECT 5.525 49.065 6.895 49.875 ;
        RECT 6.905 49.065 12.415 49.875 ;
        RECT 12.425 49.065 17.935 49.875 ;
        RECT 18.865 49.065 24.375 49.875 ;
        RECT 24.385 49.065 29.895 49.875 ;
        RECT 29.905 49.065 35.415 49.875 ;
        RECT 35.425 49.065 40.935 49.875 ;
        RECT 40.945 49.065 42.775 49.875 ;
        RECT 42.785 49.065 44.155 49.875 ;
        RECT 5.665 48.855 5.835 49.065 ;
        RECT 7.045 48.875 7.215 49.065 ;
        RECT 9.345 48.875 9.515 49.045 ;
        RECT 9.345 48.855 9.475 48.875 ;
        RECT 9.805 48.855 9.975 49.045 ;
        RECT 12.565 48.875 12.735 49.065 ;
        RECT 15.325 48.855 15.495 49.045 ;
        RECT 18.080 48.905 18.200 49.015 ;
        RECT 19.005 48.875 19.175 49.065 ;
        RECT 20.845 48.855 21.015 49.045 ;
        RECT 24.525 48.875 24.695 49.065 ;
        RECT 26.365 48.855 26.535 49.045 ;
        RECT 30.045 48.855 30.215 49.065 ;
        RECT 31.885 48.855 32.055 49.045 ;
        RECT 35.565 48.875 35.735 49.065 ;
        RECT 37.405 48.855 37.575 49.045 ;
        RECT 41.085 48.875 41.255 49.065 ;
        RECT 43.845 48.855 44.015 49.065 ;
        RECT 5.525 48.045 6.895 48.855 ;
        RECT 7.625 48.625 9.475 48.855 ;
        RECT 7.140 47.945 9.475 48.625 ;
        RECT 9.665 48.045 15.175 48.855 ;
        RECT 15.185 48.045 20.695 48.855 ;
        RECT 20.705 48.045 26.215 48.855 ;
        RECT 26.225 48.045 29.895 48.855 ;
        RECT 29.905 48.045 31.275 48.855 ;
        RECT 31.745 48.045 37.255 48.855 ;
        RECT 37.265 48.045 42.775 48.855 ;
        RECT 42.785 48.045 44.155 48.855 ;
        RECT 5.525 43.625 6.895 44.435 ;
        RECT 6.905 43.625 8.275 44.405 ;
        RECT 8.285 43.625 13.795 44.435 ;
        RECT 13.805 43.625 17.475 44.435 ;
        RECT 18.865 43.625 24.375 44.435 ;
        RECT 24.385 43.625 29.895 44.435 ;
        RECT 29.905 43.625 35.415 44.435 ;
        RECT 35.425 43.625 40.935 44.435 ;
        RECT 40.945 43.625 42.775 44.435 ;
        RECT 42.785 43.625 44.155 44.435 ;
        RECT 5.665 43.415 5.835 43.625 ;
        RECT 7.045 43.435 7.215 43.625 ;
        RECT 8.425 43.435 8.595 43.625 ;
        RECT 10.450 43.415 10.620 43.605 ;
        RECT 12.575 43.415 12.745 43.585 ;
        RECT 13.945 43.435 14.115 43.625 ;
        RECT 14.405 43.415 14.575 43.605 ;
        RECT 14.865 43.415 15.035 43.605 ;
        RECT 17.635 43.470 17.795 43.580 ;
        RECT 19.005 43.435 19.175 43.625 ;
        RECT 20.385 43.415 20.555 43.605 ;
        RECT 24.525 43.435 24.695 43.625 ;
        RECT 25.905 43.415 26.075 43.605 ;
        RECT 30.045 43.435 30.215 43.625 ;
        RECT 31.885 43.415 32.055 43.605 ;
        RECT 35.565 43.435 35.735 43.625 ;
        RECT 37.405 43.415 37.575 43.605 ;
        RECT 41.085 43.435 41.255 43.625 ;
        RECT 43.845 43.415 44.015 43.625 ;
        RECT 5.525 42.605 6.895 43.415 ;
        RECT 7.135 42.735 11.035 43.415 ;
        RECT 10.105 42.505 11.035 42.735 ;
        RECT 11.045 42.505 14.695 43.415 ;
        RECT 14.725 42.605 20.235 43.415 ;
        RECT 20.245 42.605 25.755 43.415 ;
        RECT 25.765 42.605 31.275 43.415 ;
        RECT 31.745 42.605 37.255 43.415 ;
        RECT 37.265 42.605 42.775 43.415 ;
        RECT 42.785 42.605 44.155 43.415 ;
        RECT 5.525 38.185 6.895 38.995 ;
        RECT 6.905 38.895 7.835 39.095 ;
        RECT 9.165 38.895 10.115 39.095 ;
        RECT 6.905 38.415 10.115 38.895 ;
        RECT 7.050 38.215 10.115 38.415 ;
        RECT 5.665 37.975 5.835 38.185 ;
        RECT 7.050 38.165 7.220 38.215 ;
        RECT 9.180 38.185 10.115 38.215 ;
        RECT 10.125 38.185 15.635 38.995 ;
        RECT 15.645 38.185 18.395 38.995 ;
        RECT 18.865 38.185 24.375 38.995 ;
        RECT 24.385 38.185 29.895 38.995 ;
        RECT 29.905 38.185 35.415 38.995 ;
        RECT 35.425 38.185 40.935 38.995 ;
        RECT 40.945 38.185 42.775 38.995 ;
        RECT 42.785 38.185 44.155 38.995 ;
        RECT 7.045 37.995 7.220 38.165 ;
        RECT 7.045 37.975 7.215 37.995 ;
        RECT 8.425 37.975 8.595 38.165 ;
        RECT 10.265 37.995 10.435 38.185 ;
        RECT 13.945 37.975 14.115 38.165 ;
        RECT 15.785 37.995 15.955 38.185 ;
        RECT 19.005 37.995 19.175 38.185 ;
        RECT 19.465 37.975 19.635 38.165 ;
        RECT 24.525 37.995 24.695 38.185 ;
        RECT 24.985 37.975 25.155 38.165 ;
        RECT 30.045 37.995 30.215 38.185 ;
        RECT 30.515 38.020 30.675 38.130 ;
        RECT 31.885 37.975 32.055 38.165 ;
        RECT 35.565 37.995 35.735 38.185 ;
        RECT 37.405 37.975 37.575 38.165 ;
        RECT 41.085 37.995 41.255 38.185 ;
        RECT 43.845 37.975 44.015 38.185 ;
        RECT 5.525 37.165 6.895 37.975 ;
        RECT 6.905 37.195 8.275 37.975 ;
        RECT 8.285 37.165 13.795 37.975 ;
        RECT 13.805 37.165 19.315 37.975 ;
        RECT 19.325 37.165 24.835 37.975 ;
        RECT 24.845 37.165 30.355 37.975 ;
        RECT 31.745 37.165 37.255 37.975 ;
        RECT 37.265 37.165 42.775 37.975 ;
        RECT 42.785 37.165 44.155 37.975 ;
        RECT 5.525 32.745 6.895 33.555 ;
        RECT 6.905 32.745 8.275 33.555 ;
        RECT 8.285 32.745 11.955 33.655 ;
        RECT 11.965 32.745 17.475 33.555 ;
        RECT 18.865 32.745 24.375 33.555 ;
        RECT 24.385 32.745 29.895 33.555 ;
        RECT 29.905 32.745 35.415 33.555 ;
        RECT 35.425 32.745 40.935 33.555 ;
        RECT 40.945 32.745 42.775 33.555 ;
        RECT 42.785 32.745 44.155 33.555 ;
        RECT 5.665 32.535 5.835 32.745 ;
        RECT 7.045 32.555 7.215 32.745 ;
        RECT 5.525 31.725 6.895 32.535 ;
        RECT 7.965 32.505 8.135 32.725 ;
        RECT 11.640 32.555 11.810 32.745 ;
        RECT 12.105 32.555 12.275 32.745 ;
        RECT 13.485 32.535 13.655 32.725 ;
        RECT 13.945 32.535 14.115 32.725 ;
        RECT 17.635 32.590 17.795 32.700 ;
        RECT 19.005 32.555 19.175 32.745 ;
        RECT 19.465 32.535 19.635 32.725 ;
        RECT 24.525 32.555 24.695 32.745 ;
        RECT 24.985 32.535 25.155 32.725 ;
        RECT 30.045 32.555 30.215 32.745 ;
        RECT 30.515 32.580 30.675 32.690 ;
        RECT 31.885 32.535 32.055 32.725 ;
        RECT 35.565 32.555 35.735 32.745 ;
        RECT 37.405 32.535 37.575 32.725 ;
        RECT 41.085 32.555 41.255 32.745 ;
        RECT 43.845 32.535 44.015 32.745 ;
        RECT 10.090 32.505 11.035 32.535 ;
        RECT 7.965 32.305 11.035 32.505 ;
        RECT 7.825 31.825 11.035 32.305 ;
        RECT 7.825 31.625 8.755 31.825 ;
        RECT 10.090 31.625 11.035 31.825 ;
        RECT 11.275 32.305 13.655 32.535 ;
        RECT 11.275 31.625 13.665 32.305 ;
        RECT 13.805 31.725 19.315 32.535 ;
        RECT 19.325 31.725 24.835 32.535 ;
        RECT 24.845 31.725 30.355 32.535 ;
        RECT 31.745 31.725 37.255 32.535 ;
        RECT 37.265 31.725 42.775 32.535 ;
        RECT 42.785 31.725 44.155 32.535 ;
        RECT 5.525 27.305 6.895 28.115 ;
        RECT 6.905 27.305 8.275 28.085 ;
        RECT 8.745 27.305 10.095 28.215 ;
        RECT 10.125 27.305 15.635 28.115 ;
        RECT 15.645 27.305 18.395 28.115 ;
        RECT 18.865 27.305 24.375 28.115 ;
        RECT 24.385 27.305 29.895 28.115 ;
        RECT 29.905 27.305 35.415 28.115 ;
        RECT 35.425 27.305 40.935 28.115 ;
        RECT 40.945 27.305 42.775 28.115 ;
        RECT 42.785 27.305 44.155 28.115 ;
        RECT 5.665 27.095 5.835 27.305 ;
        RECT 7.045 27.115 7.215 27.305 ;
        RECT 8.420 27.145 8.540 27.255 ;
        RECT 9.810 27.115 9.980 27.305 ;
        RECT 10.265 27.115 10.435 27.305 ;
        RECT 10.450 27.095 10.620 27.285 ;
        RECT 11.185 27.095 11.355 27.285 ;
        RECT 15.785 27.115 15.955 27.305 ;
        RECT 16.705 27.095 16.875 27.285 ;
        RECT 19.005 27.115 19.175 27.305 ;
        RECT 22.225 27.095 22.395 27.285 ;
        RECT 24.525 27.115 24.695 27.305 ;
        RECT 27.745 27.095 27.915 27.285 ;
        RECT 30.045 27.115 30.215 27.305 ;
        RECT 31.885 27.095 32.055 27.285 ;
        RECT 35.565 27.115 35.735 27.305 ;
        RECT 37.405 27.095 37.575 27.285 ;
        RECT 41.085 27.115 41.255 27.305 ;
        RECT 43.845 27.095 44.015 27.305 ;
        RECT 5.525 26.285 6.895 27.095 ;
        RECT 7.135 26.415 11.035 27.095 ;
        RECT 10.105 26.185 11.035 26.415 ;
        RECT 11.045 26.285 16.555 27.095 ;
        RECT 16.565 26.285 22.075 27.095 ;
        RECT 22.085 26.285 27.595 27.095 ;
        RECT 27.605 26.285 31.275 27.095 ;
        RECT 31.745 26.285 37.255 27.095 ;
        RECT 37.265 26.285 42.775 27.095 ;
        RECT 42.785 26.285 44.155 27.095 ;
        RECT 5.525 21.865 6.895 22.675 ;
        RECT 6.905 21.865 8.275 22.645 ;
        RECT 8.285 21.865 13.795 22.675 ;
        RECT 13.805 21.865 17.475 22.675 ;
        RECT 18.865 21.865 24.375 22.675 ;
        RECT 24.385 21.865 29.895 22.675 ;
        RECT 29.905 21.865 35.415 22.675 ;
        RECT 35.425 21.865 40.935 22.675 ;
        RECT 40.945 21.865 42.775 22.675 ;
        RECT 42.785 21.865 44.155 22.675 ;
        RECT 5.665 21.655 5.835 21.865 ;
        RECT 7.045 21.655 7.215 21.865 ;
        RECT 8.425 21.675 8.595 21.865 ;
        RECT 12.565 21.655 12.735 21.845 ;
        RECT 13.945 21.675 14.115 21.865 ;
        RECT 17.635 21.710 17.795 21.820 ;
        RECT 18.085 21.655 18.255 21.845 ;
        RECT 19.005 21.675 19.175 21.865 ;
        RECT 23.605 21.655 23.775 21.845 ;
        RECT 24.525 21.675 24.695 21.865 ;
        RECT 29.125 21.655 29.295 21.845 ;
        RECT 30.045 21.675 30.215 21.865 ;
        RECT 30.960 21.705 31.080 21.815 ;
        RECT 31.885 21.655 32.055 21.845 ;
        RECT 35.565 21.675 35.735 21.865 ;
        RECT 37.405 21.655 37.575 21.845 ;
        RECT 41.085 21.675 41.255 21.865 ;
        RECT 43.845 21.655 44.015 21.865 ;
        RECT 5.525 20.845 6.895 21.655 ;
        RECT 6.905 20.845 12.415 21.655 ;
        RECT 12.425 20.845 17.935 21.655 ;
        RECT 17.945 20.845 23.455 21.655 ;
        RECT 23.465 20.845 28.975 21.655 ;
        RECT 28.985 20.845 30.815 21.655 ;
        RECT 31.745 20.845 37.255 21.655 ;
        RECT 37.265 20.845 42.775 21.655 ;
        RECT 42.785 20.845 44.155 21.655 ;
        RECT 5.525 16.425 6.895 17.235 ;
        RECT 6.905 16.425 8.275 17.205 ;
        RECT 8.285 16.425 13.795 17.235 ;
        RECT 13.805 16.425 17.475 17.235 ;
        RECT 18.865 16.425 24.375 17.235 ;
        RECT 24.385 16.425 29.895 17.235 ;
        RECT 29.905 16.425 35.415 17.235 ;
        RECT 35.425 16.425 40.935 17.235 ;
        RECT 40.945 16.425 42.775 17.235 ;
        RECT 42.785 16.425 44.155 17.235 ;
        RECT 5.665 16.215 5.835 16.425 ;
        RECT 7.045 16.215 7.215 16.425 ;
        RECT 8.425 16.235 8.595 16.425 ;
        RECT 12.565 16.215 12.735 16.405 ;
        RECT 13.945 16.235 14.115 16.425 ;
        RECT 17.635 16.270 17.795 16.380 ;
        RECT 18.085 16.215 18.255 16.405 ;
        RECT 19.005 16.235 19.175 16.425 ;
        RECT 23.605 16.215 23.775 16.405 ;
        RECT 24.525 16.235 24.695 16.425 ;
        RECT 29.125 16.215 29.295 16.405 ;
        RECT 30.045 16.235 30.215 16.425 ;
        RECT 30.960 16.265 31.080 16.375 ;
        RECT 31.885 16.215 32.055 16.405 ;
        RECT 35.565 16.235 35.735 16.425 ;
        RECT 37.405 16.215 37.575 16.405 ;
        RECT 41.085 16.235 41.255 16.425 ;
        RECT 43.845 16.215 44.015 16.425 ;
        RECT 5.525 15.405 6.895 16.215 ;
        RECT 6.905 15.405 12.415 16.215 ;
        RECT 12.425 15.405 17.935 16.215 ;
        RECT 17.945 15.405 23.455 16.215 ;
        RECT 23.465 15.405 28.975 16.215 ;
        RECT 28.985 15.405 30.815 16.215 ;
        RECT 31.745 15.405 37.255 16.215 ;
        RECT 37.265 15.405 42.775 16.215 ;
        RECT 42.785 15.405 44.155 16.215 ;
        RECT 5.525 10.985 6.895 11.795 ;
        RECT 6.905 10.985 8.275 11.765 ;
        RECT 8.285 10.985 9.655 11.765 ;
        RECT 9.665 10.985 15.175 11.795 ;
        RECT 15.185 10.985 17.935 11.795 ;
        RECT 18.865 10.985 24.375 11.795 ;
        RECT 24.385 10.985 29.895 11.795 ;
        RECT 29.905 10.985 31.275 11.795 ;
        RECT 31.745 10.985 37.255 11.795 ;
        RECT 37.265 10.985 42.775 11.795 ;
        RECT 42.785 10.985 44.155 11.795 ;
        RECT 5.665 10.795 5.835 10.985 ;
        RECT 7.045 10.795 7.215 10.985 ;
        RECT 8.425 10.795 8.595 10.985 ;
        RECT 9.805 10.795 9.975 10.985 ;
        RECT 15.325 10.795 15.495 10.985 ;
        RECT 18.080 10.825 18.200 10.935 ;
        RECT 19.005 10.795 19.175 10.985 ;
        RECT 24.525 10.795 24.695 10.985 ;
        RECT 30.045 10.795 30.215 10.985 ;
        RECT 31.885 10.795 32.055 10.985 ;
        RECT 37.405 10.795 37.575 10.985 ;
        RECT 43.845 10.795 44.015 10.985 ;
      LAYER li1 ;
        RECT 6.985 97.335 7.245 97.665 ;
        RECT 6.985 96.425 7.155 97.335 ;
        RECT 7.940 97.265 8.145 97.665 ;
        RECT 7.940 97.095 8.625 97.265 ;
        RECT 7.865 96.425 8.115 96.925 ;
        RECT 6.985 96.255 8.115 96.425 ;
        RECT 6.985 95.485 7.255 96.255 ;
        RECT 8.285 96.065 8.625 97.095 ;
        RECT 7.960 95.890 8.625 96.065 ;
        RECT 8.825 97.160 9.085 97.665 ;
        RECT 9.775 97.285 9.945 97.665 ;
        RECT 8.825 96.360 8.995 97.160 ;
        RECT 9.280 97.115 9.945 97.285 ;
        RECT 10.205 97.160 10.465 97.665 ;
        RECT 11.155 97.285 11.325 97.665 ;
        RECT 9.280 96.860 9.450 97.115 ;
        RECT 9.165 96.530 9.450 96.860 ;
        RECT 9.280 96.385 9.450 96.530 ;
        RECT 7.960 95.485 8.145 95.890 ;
        RECT 8.825 95.455 9.095 96.360 ;
        RECT 9.280 96.215 9.945 96.385 ;
        RECT 9.775 95.455 9.945 96.215 ;
        RECT 10.205 96.360 10.375 97.160 ;
        RECT 10.660 97.115 11.325 97.285 ;
        RECT 19.035 97.285 19.205 97.665 ;
        RECT 19.035 97.115 19.750 97.285 ;
        RECT 10.660 96.860 10.830 97.115 ;
        RECT 10.545 96.530 10.830 96.860 ;
        RECT 10.660 96.385 10.830 96.530 ;
        RECT 19.580 96.925 19.750 97.115 ;
        RECT 19.920 97.090 20.175 97.665 ;
        RECT 32.335 97.265 32.540 97.665 ;
        RECT 33.235 97.335 33.495 97.665 ;
        RECT 19.580 96.595 19.835 96.925 ;
        RECT 19.580 96.385 19.750 96.595 ;
        RECT 10.205 95.455 10.475 96.360 ;
        RECT 10.660 96.215 11.325 96.385 ;
        RECT 11.155 95.455 11.325 96.215 ;
        RECT 19.035 96.215 19.750 96.385 ;
        RECT 20.005 96.360 20.175 97.090 ;
        RECT 19.035 95.455 19.205 96.215 ;
        RECT 19.920 95.455 20.175 96.360 ;
        RECT 31.855 97.095 32.540 97.265 ;
        RECT 31.855 96.065 32.195 97.095 ;
        RECT 32.365 96.425 32.615 96.925 ;
        RECT 33.325 96.425 33.495 97.335 ;
        RECT 32.365 96.255 33.495 96.425 ;
        RECT 31.855 95.890 32.520 96.065 ;
        RECT 32.335 95.485 32.520 95.890 ;
        RECT 33.225 95.485 33.495 96.255 ;
        RECT 41.485 97.160 41.745 97.665 ;
        RECT 42.435 97.285 42.605 97.665 ;
        RECT 41.485 96.360 41.665 97.160 ;
        RECT 41.940 97.115 42.605 97.285 ;
        RECT 41.940 96.860 42.110 97.115 ;
        RECT 41.835 96.530 42.110 96.860 ;
        RECT 41.940 96.385 42.110 96.530 ;
        RECT 41.485 95.455 41.755 96.360 ;
        RECT 41.940 96.215 42.615 96.385 ;
        RECT 42.435 95.455 42.615 96.215 ;
        RECT 7.075 94.185 7.245 94.945 ;
        RECT 7.075 94.015 7.740 94.185 ;
        RECT 7.925 94.040 8.195 94.945 ;
        RECT 7.570 93.870 7.740 94.015 ;
        RECT 7.570 93.540 7.855 93.870 ;
        RECT 7.570 93.285 7.740 93.540 ;
        RECT 7.075 93.115 7.740 93.285 ;
        RECT 8.025 93.240 8.195 94.040 ;
        RECT 7.075 92.735 7.245 93.115 ;
        RECT 7.935 92.735 8.195 93.240 ;
        RECT 7.075 86.405 7.245 86.785 ;
        RECT 7.075 86.235 7.740 86.405 ;
        RECT 7.935 86.280 8.195 86.785 ;
        RECT 7.570 85.980 7.740 86.235 ;
        RECT 7.570 85.650 7.855 85.980 ;
        RECT 7.570 85.505 7.740 85.650 ;
        RECT 7.075 85.335 7.740 85.505 ;
        RECT 8.025 85.480 8.195 86.280 ;
        RECT 7.075 84.575 7.245 85.335 ;
        RECT 7.925 84.575 8.195 85.480 ;
        RECT 7.075 80.965 7.245 81.340 ;
        RECT 7.915 81.175 8.990 81.345 ;
        RECT 7.915 80.965 8.085 81.175 ;
        RECT 7.075 80.795 8.085 80.965 ;
        RECT 8.310 80.835 8.650 81.005 ;
        RECT 8.820 80.840 8.990 81.175 ;
        RECT 10.280 81.175 11.880 81.345 ;
        RECT 8.310 80.665 8.600 80.835 ;
        RECT 7.050 80.495 7.395 80.605 ;
        RECT 7.045 80.325 7.395 80.495 ;
        RECT 7.050 79.985 7.395 80.325 ;
        RECT 7.705 79.985 8.140 80.605 ;
        RECT 8.310 80.145 8.480 80.665 ;
        RECT 9.160 80.495 9.520 81.170 ;
        RECT 10.280 80.805 10.450 81.175 ;
        RECT 11.525 81.135 11.880 81.175 ;
        RECT 10.620 80.755 10.950 81.005 ;
        RECT 10.635 80.680 10.950 80.755 ;
        RECT 11.120 80.885 11.290 81.005 ;
        RECT 12.395 80.885 12.640 81.305 ;
        RECT 13.410 80.945 13.585 81.275 ;
        RECT 13.930 81.185 14.100 81.345 ;
        RECT 13.930 81.015 14.460 81.185 ;
        RECT 14.630 81.175 15.625 81.345 ;
        RECT 14.630 81.015 14.800 81.175 ;
        RECT 11.120 80.715 12.640 80.885 ;
        RECT 8.980 80.315 9.520 80.495 ;
        RECT 9.160 80.205 9.520 80.315 ;
        RECT 8.310 79.975 8.945 80.145 ;
        RECT 9.160 79.975 9.965 80.205 ;
        RECT 7.075 79.635 8.605 79.805 ;
        RECT 7.075 79.135 7.245 79.635 ;
        RECT 8.435 79.475 8.605 79.635 ;
        RECT 8.775 79.645 8.945 79.975 ;
        RECT 8.775 79.475 9.105 79.645 ;
        RECT 7.915 79.305 8.085 79.465 ;
        RECT 9.275 79.305 9.445 79.805 ;
        RECT 7.915 79.135 9.445 79.305 ;
        RECT 9.615 79.135 9.965 79.975 ;
        RECT 10.165 79.605 10.465 80.605 ;
        RECT 10.635 80.155 10.805 80.680 ;
        RECT 11.120 80.675 11.290 80.715 ;
        RECT 10.975 80.495 11.305 80.505 ;
        RECT 10.975 80.335 11.360 80.495 ;
        RECT 11.190 80.325 11.360 80.335 ;
        RECT 11.700 80.155 11.945 80.545 ;
        RECT 10.635 79.985 11.395 80.155 ;
        RECT 11.645 79.985 11.945 80.155 ;
        RECT 10.725 79.305 10.895 79.815 ;
        RECT 11.065 79.475 11.395 79.985 ;
        RECT 11.700 79.925 11.945 79.985 ;
        RECT 12.150 79.925 12.480 80.545 ;
        RECT 12.955 79.925 13.245 80.605 ;
        RECT 13.415 80.495 13.585 80.945 ;
        RECT 13.880 80.665 14.120 80.835 ;
        RECT 13.415 80.325 13.705 80.495 ;
        RECT 11.565 79.515 12.630 79.685 ;
        RECT 11.565 79.305 11.735 79.515 ;
        RECT 10.725 79.135 11.735 79.305 ;
        RECT 12.460 79.135 12.630 79.515 ;
        RECT 13.415 79.465 13.585 80.325 ;
        RECT 13.400 79.135 13.585 79.465 ;
        RECT 13.880 79.465 14.050 80.665 ;
        RECT 14.290 79.845 14.460 81.015 ;
        RECT 15.110 80.835 15.285 81.005 ;
        RECT 14.870 80.675 15.285 80.835 ;
        RECT 15.455 80.885 15.625 81.175 ;
        RECT 15.455 80.715 16.025 80.885 ;
        RECT 14.870 80.665 15.280 80.675 ;
        RECT 15.090 80.325 15.545 80.495 ;
        RECT 15.855 79.935 16.025 80.715 ;
        RECT 14.290 79.615 15.075 79.845 ;
        RECT 14.745 79.475 15.075 79.615 ;
        RECT 15.375 79.765 16.025 79.935 ;
        RECT 13.880 79.135 14.090 79.465 ;
        RECT 14.260 79.305 14.590 79.345 ;
        RECT 15.375 79.305 15.545 79.765 ;
        RECT 14.260 79.135 15.545 79.305 ;
        RECT 16.215 79.135 16.475 81.345 ;
        RECT 7.075 77.865 7.245 78.625 ;
        RECT 7.075 77.695 7.740 77.865 ;
        RECT 7.925 77.720 8.195 78.625 ;
        RECT 7.570 77.550 7.740 77.695 ;
        RECT 7.570 77.220 7.855 77.550 ;
        RECT 7.570 76.965 7.740 77.220 ;
        RECT 7.075 76.795 7.740 76.965 ;
        RECT 8.025 76.920 8.195 77.720 ;
        RECT 7.075 76.415 7.245 76.795 ;
        RECT 7.935 76.415 8.195 76.920 ;
        RECT 7.075 75.525 7.245 75.900 ;
        RECT 7.915 75.735 8.990 75.905 ;
        RECT 7.915 75.525 8.085 75.735 ;
        RECT 7.075 75.355 8.085 75.525 ;
        RECT 8.310 75.395 8.650 75.565 ;
        RECT 8.820 75.400 8.990 75.735 ;
        RECT 10.280 75.735 11.880 75.905 ;
        RECT 8.310 75.225 8.600 75.395 ;
        RECT 7.050 75.055 7.395 75.165 ;
        RECT 7.045 74.885 7.395 75.055 ;
        RECT 7.050 74.545 7.395 74.885 ;
        RECT 7.705 74.545 8.140 75.165 ;
        RECT 8.310 74.705 8.480 75.225 ;
        RECT 9.160 75.055 9.520 75.730 ;
        RECT 10.280 75.365 10.450 75.735 ;
        RECT 11.525 75.695 11.880 75.735 ;
        RECT 10.620 75.315 10.950 75.565 ;
        RECT 10.635 75.240 10.950 75.315 ;
        RECT 11.120 75.445 11.290 75.565 ;
        RECT 12.395 75.445 12.640 75.865 ;
        RECT 13.410 75.505 13.585 75.835 ;
        RECT 13.930 75.745 14.100 75.905 ;
        RECT 13.930 75.575 14.460 75.745 ;
        RECT 14.630 75.735 15.625 75.905 ;
        RECT 14.630 75.575 14.800 75.735 ;
        RECT 11.120 75.275 12.640 75.445 ;
        RECT 8.980 74.875 9.520 75.055 ;
        RECT 9.160 74.765 9.520 74.875 ;
        RECT 8.310 74.535 8.945 74.705 ;
        RECT 9.160 74.535 9.965 74.765 ;
        RECT 7.075 74.195 8.605 74.365 ;
        RECT 7.075 73.695 7.245 74.195 ;
        RECT 8.435 74.035 8.605 74.195 ;
        RECT 8.775 74.205 8.945 74.535 ;
        RECT 8.775 74.035 9.105 74.205 ;
        RECT 7.915 73.865 8.085 74.025 ;
        RECT 9.275 73.865 9.445 74.365 ;
        RECT 7.915 73.695 9.445 73.865 ;
        RECT 9.615 73.695 9.965 74.535 ;
        RECT 10.165 74.165 10.465 75.165 ;
        RECT 10.635 74.715 10.805 75.240 ;
        RECT 11.120 75.235 11.290 75.275 ;
        RECT 10.975 75.055 11.305 75.065 ;
        RECT 10.975 74.895 11.360 75.055 ;
        RECT 11.190 74.885 11.360 74.895 ;
        RECT 11.700 74.715 11.945 75.105 ;
        RECT 10.635 74.545 11.395 74.715 ;
        RECT 11.645 74.545 11.945 74.715 ;
        RECT 10.725 73.865 10.895 74.375 ;
        RECT 11.065 74.035 11.395 74.545 ;
        RECT 11.700 74.485 11.945 74.545 ;
        RECT 12.150 74.485 12.480 75.105 ;
        RECT 12.955 74.485 13.245 75.165 ;
        RECT 13.415 75.055 13.585 75.505 ;
        RECT 13.880 75.225 14.120 75.395 ;
        RECT 13.415 74.885 13.705 75.055 ;
        RECT 11.565 74.075 12.630 74.245 ;
        RECT 11.565 73.865 11.735 74.075 ;
        RECT 10.725 73.695 11.735 73.865 ;
        RECT 12.460 73.695 12.630 74.075 ;
        RECT 13.415 74.025 13.585 74.885 ;
        RECT 13.400 73.695 13.585 74.025 ;
        RECT 13.880 74.025 14.050 75.225 ;
        RECT 14.290 74.405 14.460 75.575 ;
        RECT 15.110 75.395 15.285 75.565 ;
        RECT 14.870 75.235 15.285 75.395 ;
        RECT 15.455 75.445 15.625 75.735 ;
        RECT 15.455 75.275 16.025 75.445 ;
        RECT 14.870 75.225 15.280 75.235 ;
        RECT 15.090 74.885 15.545 75.055 ;
        RECT 15.855 74.495 16.025 75.275 ;
        RECT 14.290 74.175 15.075 74.405 ;
        RECT 14.745 74.035 15.075 74.175 ;
        RECT 15.375 74.325 16.025 74.495 ;
        RECT 13.880 73.695 14.090 74.025 ;
        RECT 14.260 73.865 14.590 73.905 ;
        RECT 15.375 73.865 15.545 74.325 ;
        RECT 14.260 73.695 15.545 73.865 ;
        RECT 16.215 73.695 16.475 75.905 ;
        RECT 7.075 72.425 7.245 73.185 ;
        RECT 7.075 72.255 7.740 72.425 ;
        RECT 7.925 72.280 8.195 73.185 ;
        RECT 7.570 72.110 7.740 72.255 ;
        RECT 7.570 71.780 7.855 72.110 ;
        RECT 7.570 71.525 7.740 71.780 ;
        RECT 7.075 71.355 7.740 71.525 ;
        RECT 8.025 71.480 8.195 72.280 ;
        RECT 7.075 70.975 7.245 71.355 ;
        RECT 7.935 70.975 8.195 71.480 ;
        RECT 11.590 72.215 11.925 73.185 ;
        RECT 12.435 73.015 14.465 73.185 ;
        RECT 11.590 71.545 11.760 72.215 ;
        RECT 12.435 72.045 12.605 73.015 ;
        RECT 11.930 71.715 12.185 72.045 ;
        RECT 12.410 71.715 12.605 72.045 ;
        RECT 12.775 72.675 13.900 72.845 ;
        RECT 12.015 71.545 12.185 71.715 ;
        RECT 12.775 71.545 12.945 72.675 ;
        RECT 11.590 70.975 11.845 71.545 ;
        RECT 12.015 71.375 12.945 71.545 ;
        RECT 13.115 72.335 14.125 72.505 ;
        RECT 13.115 71.535 13.285 72.335 ;
        RECT 13.490 71.655 13.765 72.135 ;
        RECT 13.485 71.485 13.765 71.655 ;
        RECT 12.770 71.340 12.945 71.375 ;
        RECT 12.770 70.975 13.300 71.340 ;
        RECT 13.490 70.975 13.765 71.485 ;
        RECT 13.935 70.975 14.125 72.335 ;
        RECT 14.295 72.350 14.465 73.015 ;
        RECT 15.040 72.595 15.555 73.005 ;
        RECT 14.295 72.160 15.045 72.350 ;
        RECT 15.215 71.785 15.555 72.595 ;
        RECT 14.325 71.615 15.555 71.785 ;
        RECT 15.035 71.010 15.280 71.615 ;
        RECT 7.075 66.985 7.245 67.745 ;
        RECT 7.075 66.815 7.740 66.985 ;
        RECT 7.925 66.840 8.195 67.745 ;
        RECT 7.570 66.670 7.740 66.815 ;
        RECT 7.570 66.340 7.855 66.670 ;
        RECT 7.570 66.085 7.740 66.340 ;
        RECT 7.075 65.915 7.740 66.085 ;
        RECT 8.025 66.040 8.195 66.840 ;
        RECT 7.075 65.535 7.245 65.915 ;
        RECT 7.935 65.535 8.195 66.040 ;
        RECT 11.595 61.505 11.925 62.290 ;
        RECT 11.595 61.335 12.275 61.505 ;
        RECT 11.585 60.915 11.935 61.165 ;
        RECT 12.105 60.735 12.275 61.335 ;
        RECT 12.445 60.915 12.795 61.165 ;
        RECT 12.015 60.095 12.345 60.735 ;
        RECT 7.075 59.205 7.245 59.585 ;
        RECT 7.075 59.035 7.740 59.205 ;
        RECT 7.935 59.080 8.195 59.585 ;
        RECT 7.570 58.780 7.740 59.035 ;
        RECT 7.570 58.450 7.855 58.780 ;
        RECT 7.570 58.305 7.740 58.450 ;
        RECT 7.075 58.135 7.740 58.305 ;
        RECT 8.025 58.280 8.195 59.080 ;
        RECT 12.565 59.225 12.885 59.585 ;
        RECT 13.880 59.225 14.225 59.585 ;
        RECT 12.565 59.055 14.225 59.225 ;
        RECT 7.075 57.375 7.245 58.135 ;
        RECT 7.925 57.375 8.195 58.280 ;
        RECT 12.105 58.215 12.380 58.845 ;
        RECT 12.090 57.555 12.395 58.045 ;
        RECT 12.565 57.725 12.865 59.055 ;
        RECT 13.245 58.595 13.575 58.765 ;
        RECT 13.250 58.345 13.575 58.595 ;
        RECT 13.755 58.515 14.365 58.845 ;
        RECT 14.535 58.345 15.035 58.805 ;
        RECT 13.250 58.165 15.035 58.345 ;
        RECT 13.035 57.815 15.070 57.985 ;
        RECT 13.035 57.555 13.365 57.815 ;
        RECT 12.090 57.375 13.365 57.555 ;
        RECT 13.960 57.735 15.070 57.815 ;
        RECT 13.960 57.375 14.130 57.735 ;
        RECT 14.810 57.375 15.070 57.735 ;
        RECT 35.935 56.015 36.265 56.865 ;
        RECT 36.775 56.015 37.105 56.865 ;
        RECT 35.935 55.845 37.435 56.015 ;
        RECT 35.555 55.475 37.080 55.675 ;
        RECT 37.260 55.645 37.435 55.845 ;
        RECT 37.260 55.475 39.885 55.645 ;
        RECT 37.260 55.305 37.435 55.475 ;
        RECT 36.015 55.135 37.435 55.305 ;
        RECT 36.015 54.655 36.185 55.135 ;
        RECT 36.855 54.660 37.025 55.135 ;
        RECT 7.075 53.765 7.245 54.145 ;
        RECT 7.075 53.595 7.740 53.765 ;
        RECT 7.935 53.640 8.195 54.145 ;
        RECT 7.570 53.340 7.740 53.595 ;
        RECT 7.570 53.010 7.855 53.340 ;
        RECT 7.570 52.865 7.740 53.010 ;
        RECT 7.075 52.695 7.740 52.865 ;
        RECT 8.025 52.840 8.195 53.640 ;
        RECT 7.075 51.935 7.245 52.695 ;
        RECT 7.925 51.935 8.195 52.840 ;
        RECT 7.310 48.305 7.480 48.555 ;
        RECT 6.985 48.135 7.480 48.305 ;
        RECT 8.215 48.305 8.385 48.650 ;
        RECT 9.055 48.305 9.575 48.705 ;
        RECT 8.215 48.135 9.575 48.305 ;
        RECT 6.985 47.175 7.155 48.135 ;
        RECT 7.325 47.345 7.675 47.965 ;
        RECT 7.845 47.345 8.185 47.965 ;
        RECT 8.355 47.345 8.595 47.965 ;
        RECT 8.775 47.715 9.235 47.885 ;
        RECT 8.775 47.175 8.945 47.715 ;
        RECT 9.405 47.515 9.575 48.135 ;
        RECT 6.985 47.005 8.945 47.175 ;
        RECT 9.115 46.505 9.575 47.515 ;
        RECT 7.075 45.225 7.245 45.985 ;
        RECT 7.075 45.055 7.740 45.225 ;
        RECT 7.925 45.080 8.195 45.985 ;
        RECT 7.570 44.910 7.740 45.055 ;
        RECT 7.570 44.580 7.855 44.910 ;
        RECT 7.570 44.325 7.740 44.580 ;
        RECT 7.075 44.155 7.740 44.325 ;
        RECT 8.025 44.280 8.195 45.080 ;
        RECT 7.075 43.775 7.245 44.155 ;
        RECT 7.935 43.775 8.195 44.280 ;
        RECT 7.260 42.625 7.505 43.230 ;
        RECT 6.985 42.455 8.215 42.625 ;
        RECT 6.985 41.645 7.325 42.455 ;
        RECT 7.495 41.890 8.245 42.080 ;
        RECT 6.985 41.235 7.500 41.645 ;
        RECT 8.075 41.225 8.245 41.890 ;
        RECT 8.415 41.905 8.605 43.265 ;
        RECT 8.775 43.095 9.050 43.265 ;
        RECT 8.775 42.925 9.055 43.095 ;
        RECT 8.775 42.105 9.050 42.925 ;
        RECT 9.240 42.900 9.770 43.265 ;
        RECT 9.595 42.865 9.770 42.900 ;
        RECT 9.255 41.905 9.425 42.705 ;
        RECT 8.415 41.735 9.425 41.905 ;
        RECT 9.595 42.695 10.525 42.865 ;
        RECT 10.695 42.695 10.950 43.265 ;
        RECT 9.595 41.565 9.765 42.695 ;
        RECT 10.355 42.525 10.525 42.695 ;
        RECT 8.640 41.395 9.765 41.565 ;
        RECT 9.935 42.195 10.130 42.525 ;
        RECT 10.355 42.195 10.610 42.525 ;
        RECT 9.935 41.225 10.105 42.195 ;
        RECT 10.780 42.025 10.950 42.695 ;
        RECT 11.630 42.500 11.815 43.170 ;
        RECT 12.300 42.815 12.630 43.215 ;
        RECT 13.345 42.820 13.675 43.260 ;
        RECT 13.345 42.815 14.575 42.820 ;
        RECT 12.300 42.705 14.575 42.815 ;
        RECT 12.420 42.640 14.575 42.705 ;
        RECT 11.180 42.230 11.815 42.500 ;
        RECT 11.995 42.120 12.280 42.525 ;
        RECT 12.450 42.120 12.780 42.470 ;
        RECT 8.075 41.055 10.105 41.225 ;
        RECT 10.615 41.055 10.950 42.025 ;
        RECT 11.215 41.770 12.325 41.940 ;
        RECT 11.215 41.060 11.410 41.770 ;
        RECT 12.095 41.060 12.325 41.770 ;
        RECT 12.505 41.065 12.780 42.120 ;
        RECT 12.950 41.065 13.285 42.470 ;
        RECT 13.485 41.065 13.935 42.470 ;
        RECT 14.190 41.060 14.575 42.640 ;
        RECT 6.985 39.155 7.325 40.035 ;
        RECT 7.495 39.325 7.665 40.545 ;
        RECT 8.690 40.205 9.165 40.545 ;
        RECT 7.905 39.675 8.155 40.040 ;
        RECT 8.875 39.675 9.590 39.970 ;
        RECT 9.760 39.845 10.035 40.545 ;
        RECT 7.905 39.505 9.695 39.675 ;
        RECT 7.495 39.075 8.290 39.325 ;
        RECT 7.495 38.985 7.745 39.075 ;
        RECT 7.415 38.565 7.745 38.985 ;
        RECT 8.460 38.650 8.715 39.505 ;
        RECT 7.925 38.385 8.715 38.650 ;
        RECT 8.885 38.805 9.295 39.325 ;
        RECT 9.465 39.075 9.695 39.505 ;
        RECT 9.865 38.815 10.035 39.845 ;
        RECT 8.885 38.385 9.085 38.805 ;
        RECT 9.775 38.335 10.035 38.815 ;
        RECT 7.075 37.445 7.245 37.825 ;
        RECT 7.075 37.275 7.740 37.445 ;
        RECT 7.935 37.320 8.195 37.825 ;
        RECT 7.570 37.020 7.740 37.275 ;
        RECT 7.570 36.690 7.855 37.020 ;
        RECT 7.570 36.545 7.740 36.690 ;
        RECT 7.075 36.375 7.740 36.545 ;
        RECT 8.025 36.520 8.195 37.320 ;
        RECT 7.075 35.615 7.245 36.375 ;
        RECT 7.925 35.615 8.195 36.520 ;
        RECT 8.455 34.605 8.625 35.105 ;
        RECT 9.415 34.605 9.585 35.105 ;
        RECT 10.255 34.605 10.425 35.105 ;
        RECT 8.455 34.435 10.425 34.605 ;
        RECT 10.595 34.635 10.925 35.065 ;
        RECT 11.535 34.805 11.875 35.065 ;
        RECT 10.595 34.465 11.445 34.635 ;
        RECT 8.390 33.635 8.645 34.265 ;
        RECT 8.875 33.635 9.255 34.265 ;
        RECT 10.125 34.255 10.425 34.260 ;
        RECT 10.125 34.085 10.435 34.255 ;
        RECT 10.125 33.965 10.425 34.085 ;
        RECT 8.875 33.035 9.080 33.635 ;
        RECT 9.515 33.240 9.735 33.965 ;
        RECT 10.045 33.635 10.425 33.965 ;
        RECT 10.625 33.715 10.955 34.275 ;
        RECT 11.275 33.545 11.445 34.465 ;
        RECT 10.625 33.450 11.445 33.545 ;
        RECT 10.430 33.375 11.445 33.450 ;
        RECT 9.310 33.055 10.260 33.240 ;
        RECT 10.430 32.940 10.845 33.375 ;
        RECT 11.615 33.200 11.875 34.805 ;
        RECT 11.535 32.940 11.875 33.200 ;
        RECT 8.335 31.735 8.665 32.155 ;
        RECT 8.845 31.985 9.105 32.385 ;
        RECT 9.775 31.985 9.945 32.335 ;
        RECT 8.845 31.815 10.510 31.985 ;
        RECT 10.680 31.880 10.955 32.225 ;
        RECT 8.415 31.645 8.665 31.735 ;
        RECT 10.340 31.645 10.510 31.815 ;
        RECT 7.910 31.315 8.245 31.565 ;
        RECT 8.415 31.315 9.130 31.645 ;
        RECT 9.345 31.315 10.170 31.645 ;
        RECT 10.340 31.315 10.615 31.645 ;
        RECT 8.415 30.755 8.585 31.315 ;
        RECT 8.845 30.855 9.175 31.145 ;
        RECT 9.345 31.025 9.590 31.315 ;
        RECT 10.340 31.145 10.510 31.315 ;
        RECT 10.785 31.145 10.955 31.880 ;
        RECT 9.850 30.975 10.510 31.145 ;
        RECT 9.850 30.855 10.020 30.975 ;
        RECT 8.845 30.685 10.020 30.855 ;
        RECT 8.405 30.185 10.020 30.515 ;
        RECT 10.680 30.175 10.955 31.145 ;
        RECT 11.125 32.155 11.715 32.385 ;
        RECT 11.125 31.145 11.415 32.155 ;
        RECT 13.290 31.985 13.715 32.195 ;
        RECT 11.585 31.815 13.715 31.985 ;
        RECT 11.585 31.315 11.755 31.815 ;
        RECT 12.045 31.315 12.375 31.645 ;
        RECT 12.565 31.315 12.835 31.645 ;
        RECT 13.025 31.315 13.375 31.645 ;
        RECT 11.125 30.975 12.670 31.145 ;
        RECT 13.545 31.045 13.715 31.815 ;
        RECT 11.125 30.175 11.715 30.975 ;
        RECT 12.340 30.175 12.670 30.975 ;
        RECT 13.290 30.715 13.715 31.045 ;
        RECT 7.075 28.905 7.245 29.665 ;
        RECT 7.075 28.735 7.740 28.905 ;
        RECT 7.925 28.760 8.195 29.665 ;
        RECT 7.570 28.590 7.740 28.735 ;
        RECT 7.570 28.260 7.855 28.590 ;
        RECT 7.570 28.005 7.740 28.260 ;
        RECT 7.075 27.835 7.740 28.005 ;
        RECT 8.025 27.960 8.195 28.760 ;
        RECT 9.255 28.685 9.585 29.665 ;
        RECT 8.845 28.275 9.180 28.525 ;
        RECT 9.350 28.085 9.520 28.685 ;
        RECT 9.690 28.255 10.025 28.525 ;
        RECT 7.075 27.455 7.245 27.835 ;
        RECT 7.935 27.455 8.195 27.960 ;
        RECT 8.825 27.455 9.520 28.085 ;
        RECT 7.260 26.305 7.505 26.910 ;
        RECT 6.985 26.135 8.215 26.305 ;
        RECT 6.985 25.325 7.325 26.135 ;
        RECT 7.495 25.570 8.245 25.760 ;
        RECT 6.985 24.915 7.500 25.325 ;
        RECT 8.075 24.905 8.245 25.570 ;
        RECT 8.415 25.585 8.605 26.945 ;
        RECT 8.775 26.095 9.050 26.945 ;
        RECT 9.240 26.580 9.770 26.945 ;
        RECT 9.595 26.545 9.770 26.580 ;
        RECT 8.775 25.925 9.055 26.095 ;
        RECT 8.775 25.785 9.050 25.925 ;
        RECT 9.255 25.585 9.425 26.385 ;
        RECT 8.415 25.415 9.425 25.585 ;
        RECT 9.595 26.375 10.525 26.545 ;
        RECT 10.695 26.375 10.950 26.945 ;
        RECT 9.595 25.245 9.765 26.375 ;
        RECT 10.355 26.205 10.525 26.375 ;
        RECT 8.640 25.075 9.765 25.245 ;
        RECT 9.935 25.875 10.130 26.205 ;
        RECT 10.355 25.875 10.610 26.205 ;
        RECT 9.935 24.905 10.105 25.875 ;
        RECT 10.780 25.705 10.950 26.375 ;
        RECT 8.075 24.735 10.105 24.905 ;
        RECT 10.615 24.735 10.950 25.705 ;
        RECT 7.075 23.465 7.245 24.225 ;
        RECT 7.075 23.295 7.740 23.465 ;
        RECT 7.925 23.320 8.195 24.225 ;
        RECT 7.570 23.150 7.740 23.295 ;
        RECT 7.570 22.820 7.855 23.150 ;
        RECT 7.570 22.565 7.740 22.820 ;
        RECT 7.075 22.395 7.740 22.565 ;
        RECT 8.025 22.520 8.195 23.320 ;
        RECT 7.075 22.015 7.245 22.395 ;
        RECT 7.935 22.015 8.195 22.520 ;
        RECT 7.075 18.025 7.245 18.785 ;
        RECT 7.075 17.855 7.740 18.025 ;
        RECT 7.925 17.880 8.195 18.785 ;
        RECT 7.570 17.710 7.740 17.855 ;
        RECT 7.570 17.380 7.855 17.710 ;
        RECT 7.570 17.125 7.740 17.380 ;
        RECT 7.075 16.955 7.740 17.125 ;
        RECT 8.025 17.080 8.195 17.880 ;
        RECT 7.075 16.575 7.245 16.955 ;
        RECT 7.935 16.575 8.195 17.080 ;
        RECT 7.075 12.585 7.245 13.345 ;
        RECT 7.075 12.415 7.740 12.585 ;
        RECT 7.925 12.440 8.195 13.345 ;
        RECT 7.570 12.270 7.740 12.415 ;
        RECT 7.570 11.940 7.855 12.270 ;
        RECT 7.570 11.685 7.740 11.940 ;
        RECT 7.075 11.515 7.740 11.685 ;
        RECT 8.025 11.640 8.195 12.440 ;
        RECT 8.455 12.585 8.625 13.345 ;
        RECT 8.455 12.415 9.120 12.585 ;
        RECT 9.305 12.440 9.575 13.345 ;
        RECT 8.950 12.270 9.120 12.415 ;
        RECT 8.950 11.940 9.235 12.270 ;
        RECT 8.950 11.685 9.120 11.940 ;
        RECT 7.075 11.135 7.245 11.515 ;
        RECT 7.935 11.135 8.195 11.640 ;
        RECT 8.455 11.515 9.120 11.685 ;
        RECT 9.405 11.640 9.575 12.440 ;
        RECT 8.455 11.135 8.625 11.515 ;
        RECT 9.315 11.135 9.575 11.640 ;
      LAYER met1 ;
        RECT 8.810 97.480 9.130 97.540 ;
        RECT 10.205 97.480 10.495 97.525 ;
        RECT 8.810 97.340 10.495 97.480 ;
        RECT 8.810 97.280 9.130 97.340 ;
        RECT 10.205 97.295 10.495 97.340 ;
        RECT 12.490 97.480 12.810 97.540 ;
        RECT 19.865 97.480 20.155 97.525 ;
        RECT 12.490 97.340 20.155 97.480 ;
        RECT 12.490 97.280 12.810 97.340 ;
        RECT 19.865 97.295 20.155 97.340 ;
        RECT 8.365 96.460 8.655 96.505 ;
        RECT 11.570 96.460 11.890 96.520 ;
        RECT 8.365 96.320 11.890 96.460 ;
        RECT 8.365 96.275 8.655 96.320 ;
        RECT 11.570 96.260 11.890 96.320 ;
        RECT 31.810 95.920 32.130 96.180 ;
        RECT 8.350 95.780 8.670 95.840 ;
        RECT 8.825 95.780 9.115 95.825 ;
        RECT 8.350 95.640 9.115 95.780 ;
        RECT 8.350 95.580 8.670 95.640 ;
        RECT 8.825 95.595 9.115 95.640 ;
        RECT 41.470 95.580 41.790 95.840 ;
        RECT 7.890 92.860 8.210 93.120 ;
        RECT 6.970 84.900 7.290 84.960 ;
        RECT 7.905 84.900 8.195 84.945 ;
        RECT 6.970 84.760 8.195 84.900 ;
        RECT 6.970 84.700 7.290 84.760 ;
        RECT 7.905 84.715 8.195 84.760 ;
        RECT 7.430 83.200 7.750 83.260 ;
        RECT 8.350 83.200 8.670 83.260 ;
        RECT 7.430 83.060 8.670 83.200 ;
        RECT 7.430 83.000 7.750 83.060 ;
        RECT 8.350 83.000 8.670 83.060 ;
        RECT 8.370 80.820 8.660 80.865 ;
        RECT 13.890 80.820 14.180 80.865 ;
        RECT 14.810 80.820 15.100 80.865 ;
        RECT 8.370 80.680 15.100 80.820 ;
        RECT 8.370 80.635 8.660 80.680 ;
        RECT 13.890 80.635 14.180 80.680 ;
        RECT 14.810 80.635 15.100 80.680 ;
        RECT 6.985 80.480 7.275 80.525 ;
        RECT 7.430 80.480 7.750 80.540 ;
        RECT 6.985 80.340 7.750 80.480 ;
        RECT 6.985 80.295 7.275 80.340 ;
        RECT 7.430 80.280 7.750 80.340 ;
        RECT 7.890 80.280 8.210 80.540 ;
        RECT 9.290 80.480 9.580 80.525 ;
        RECT 11.130 80.480 11.420 80.525 ;
        RECT 9.290 80.340 11.420 80.480 ;
        RECT 9.290 80.295 9.580 80.340 ;
        RECT 11.130 80.295 11.420 80.340 ;
        RECT 13.475 80.480 13.765 80.525 ;
        RECT 15.315 80.480 15.605 80.525 ;
        RECT 13.475 80.340 15.605 80.480 ;
        RECT 13.475 80.295 13.765 80.340 ;
        RECT 15.315 80.295 15.605 80.340 ;
        RECT 31.810 80.280 32.130 80.540 ;
        RECT 12.030 80.185 12.350 80.200 ;
        RECT 11.585 80.140 11.875 80.185 ;
        RECT 7.520 80.000 11.875 80.140 ;
        RECT 7.520 79.860 7.660 80.000 ;
        RECT 11.585 79.955 11.875 80.000 ;
        RECT 12.030 79.955 12.460 80.185 ;
        RECT 12.950 80.140 13.270 80.200 ;
        RECT 31.900 80.140 32.040 80.280 ;
        RECT 12.950 80.000 32.040 80.140 ;
        RECT 12.030 79.940 12.350 79.955 ;
        RECT 12.950 79.940 13.270 80.000 ;
        RECT 7.430 79.600 7.750 79.860 ;
        RECT 10.205 79.615 10.495 79.845 ;
        RECT 11.165 79.800 11.455 79.845 ;
        RECT 14.395 79.800 14.685 79.845 ;
        RECT 11.165 79.660 14.685 79.800 ;
        RECT 11.165 79.615 11.455 79.660 ;
        RECT 14.395 79.615 14.685 79.660 ;
        RECT 10.280 79.460 10.420 79.615 ;
        RECT 12.490 79.460 12.810 79.520 ;
        RECT 10.280 79.320 12.810 79.460 ;
        RECT 12.490 79.260 12.810 79.320 ;
        RECT 13.870 79.460 14.190 79.520 ;
        RECT 16.185 79.460 16.475 79.505 ;
        RECT 13.870 79.320 16.475 79.460 ;
        RECT 13.870 79.260 14.190 79.320 ;
        RECT 16.185 79.275 16.475 79.320 ;
        RECT 7.905 78.440 8.195 78.485 ;
        RECT 12.030 78.440 12.350 78.500 ;
        RECT 7.905 78.300 12.350 78.440 ;
        RECT 7.905 78.255 8.195 78.300 ;
        RECT 12.030 78.240 12.350 78.300 ;
        RECT 8.370 75.380 8.660 75.425 ;
        RECT 13.890 75.380 14.180 75.425 ;
        RECT 14.810 75.380 15.100 75.425 ;
        RECT 8.370 75.240 15.100 75.380 ;
        RECT 8.370 75.195 8.660 75.240 ;
        RECT 13.890 75.195 14.180 75.240 ;
        RECT 14.810 75.195 15.100 75.240 ;
        RECT 6.970 74.840 7.290 75.100 ;
        RECT 7.890 74.840 8.210 75.100 ;
        RECT 9.290 75.040 9.580 75.085 ;
        RECT 11.130 75.040 11.420 75.085 ;
        RECT 9.290 74.900 11.420 75.040 ;
        RECT 9.290 74.855 9.580 74.900 ;
        RECT 11.130 74.855 11.420 74.900 ;
        RECT 12.950 74.840 13.270 75.100 ;
        RECT 13.475 75.040 13.765 75.085 ;
        RECT 15.315 75.040 15.605 75.085 ;
        RECT 13.475 74.900 15.605 75.040 ;
        RECT 13.475 74.855 13.765 74.900 ;
        RECT 15.315 74.855 15.605 74.900 ;
        RECT 8.810 74.700 9.130 74.760 ;
        RECT 12.030 74.745 12.350 74.760 ;
        RECT 11.585 74.700 11.875 74.745 ;
        RECT 8.810 74.560 11.875 74.700 ;
        RECT 8.810 74.500 9.130 74.560 ;
        RECT 11.585 74.515 11.875 74.560 ;
        RECT 12.030 74.515 12.460 74.745 ;
        RECT 12.030 74.500 12.350 74.515 ;
        RECT 10.205 74.175 10.495 74.405 ;
        RECT 11.165 74.360 11.455 74.405 ;
        RECT 14.395 74.360 14.685 74.405 ;
        RECT 11.165 74.220 14.685 74.360 ;
        RECT 11.165 74.175 11.455 74.220 ;
        RECT 14.395 74.175 14.685 74.220 ;
        RECT 8.350 74.020 8.670 74.080 ;
        RECT 10.280 74.020 10.420 74.175 ;
        RECT 12.490 74.020 12.810 74.080 ;
        RECT 8.350 73.880 12.810 74.020 ;
        RECT 8.350 73.820 8.670 73.880 ;
        RECT 12.490 73.820 12.810 73.880 ;
        RECT 16.170 73.820 16.490 74.080 ;
        RECT 7.905 73.000 8.195 73.045 ;
        RECT 12.030 73.000 12.350 73.060 ;
        RECT 16.170 73.000 16.490 73.060 ;
        RECT 7.905 72.860 12.350 73.000 ;
        RECT 7.905 72.815 8.195 72.860 ;
        RECT 12.030 72.800 12.350 72.860 ;
        RECT 13.960 72.860 16.490 73.000 ;
        RECT 7.890 72.320 8.210 72.380 ;
        RECT 11.570 72.320 11.890 72.380 ;
        RECT 13.960 72.365 14.100 72.860 ;
        RECT 16.170 72.800 16.490 72.860 ;
        RECT 7.890 72.180 13.640 72.320 ;
        RECT 7.890 72.120 8.210 72.180 ;
        RECT 11.570 72.120 11.890 72.180 ;
        RECT 13.500 71.980 13.640 72.180 ;
        RECT 13.885 72.135 14.175 72.365 ;
        RECT 14.345 72.135 14.635 72.365 ;
        RECT 14.420 71.980 14.560 72.135 ;
        RECT 13.500 71.840 14.560 71.980 ;
        RECT 13.425 71.640 13.715 71.685 ;
        RECT 13.870 71.640 14.190 71.700 ;
        RECT 13.425 71.500 14.190 71.640 ;
        RECT 13.425 71.455 13.715 71.500 ;
        RECT 13.870 71.440 14.190 71.500 ;
        RECT 11.570 71.100 11.890 71.360 ;
        RECT 7.430 67.560 7.750 67.620 ;
        RECT 7.905 67.560 8.195 67.605 ;
        RECT 7.430 67.420 8.195 67.560 ;
        RECT 7.430 67.360 7.750 67.420 ;
        RECT 7.905 67.375 8.195 67.420 ;
        RECT 11.570 60.900 11.890 61.160 ;
        RECT 12.505 61.100 12.795 61.145 ;
        RECT 13.870 61.100 14.190 61.160 ;
        RECT 41.470 61.100 41.790 61.160 ;
        RECT 12.505 60.960 41.790 61.100 ;
        RECT 12.505 60.915 12.795 60.960 ;
        RECT 13.870 60.900 14.190 60.960 ;
        RECT 41.470 60.900 41.790 60.960 ;
        RECT 12.030 60.220 12.350 60.480 ;
        RECT 7.905 59.400 8.195 59.445 ;
        RECT 8.810 59.400 9.130 59.460 ;
        RECT 7.905 59.260 9.130 59.400 ;
        RECT 7.905 59.215 8.195 59.260 ;
        RECT 8.810 59.200 9.130 59.260 ;
        RECT 12.030 59.200 12.350 59.460 ;
        RECT 13.870 59.200 14.190 59.460 ;
        RECT 12.120 58.765 12.260 59.200 ;
        RECT 13.960 58.765 14.100 59.200 ;
        RECT 12.045 58.535 12.335 58.765 ;
        RECT 13.885 58.535 14.175 58.765 ;
        RECT 14.790 58.180 15.110 58.440 ;
        RECT 12.490 57.840 12.810 58.100 ;
        RECT 12.490 56.680 12.810 56.740 ;
        RECT 12.490 56.540 34.570 56.680 ;
        RECT 12.490 56.480 12.810 56.540 ;
        RECT 34.430 55.660 34.570 56.540 ;
        RECT 35.505 55.660 35.795 55.705 ;
        RECT 34.430 55.520 35.795 55.660 ;
        RECT 35.505 55.475 35.795 55.520 ;
        RECT 7.430 52.260 7.750 52.320 ;
        RECT 7.905 52.260 8.195 52.305 ;
        RECT 7.430 52.120 8.195 52.260 ;
        RECT 7.430 52.060 7.750 52.120 ;
        RECT 7.905 52.075 8.195 52.120 ;
        RECT 7.890 47.640 8.210 47.900 ;
        RECT 8.350 47.640 8.670 47.900 ;
        RECT 7.430 47.300 7.750 47.560 ;
        RECT 7.980 47.500 8.120 47.640 ;
        RECT 12.030 47.500 12.350 47.560 ;
        RECT 7.980 47.360 12.350 47.500 ;
        RECT 12.030 47.300 12.350 47.360 ;
        RECT 9.285 46.820 9.575 46.865 ;
        RECT 12.950 46.820 13.270 46.880 ;
        RECT 9.285 46.680 13.270 46.820 ;
        RECT 9.285 46.635 9.575 46.680 ;
        RECT 12.950 46.620 13.270 46.680 ;
        RECT 7.890 43.900 8.210 44.160 ;
        RECT 7.890 43.080 8.210 43.140 ;
        RECT 8.825 43.080 9.115 43.125 ;
        RECT 7.890 42.940 9.115 43.080 ;
        RECT 7.890 42.880 8.210 42.940 ;
        RECT 8.825 42.895 9.115 42.940 ;
        RECT 10.665 43.080 10.955 43.125 ;
        RECT 11.585 43.080 11.875 43.125 ;
        RECT 10.665 42.940 11.875 43.080 ;
        RECT 10.665 42.895 10.955 42.940 ;
        RECT 11.585 42.895 11.875 42.940 ;
        RECT 12.030 42.880 12.350 43.140 ;
        RECT 12.950 42.880 13.270 43.140 ;
        RECT 13.410 42.880 13.730 43.140 ;
        RECT 8.350 42.740 8.670 42.800 ;
        RECT 7.980 42.600 8.670 42.740 ;
        RECT 7.980 42.105 8.120 42.600 ;
        RECT 8.350 42.540 8.670 42.600 ;
        RECT 12.120 42.445 12.260 42.880 ;
        RECT 12.045 42.215 12.335 42.445 ;
        RECT 12.490 42.200 12.810 42.460 ;
        RECT 13.040 42.445 13.180 42.880 ;
        RECT 12.965 42.215 13.255 42.445 ;
        RECT 7.905 41.875 8.195 42.105 ;
        RECT 8.350 41.860 8.670 42.120 ;
        RECT 12.580 42.060 12.720 42.200 ;
        RECT 13.425 42.060 13.715 42.105 ;
        RECT 12.580 41.920 13.715 42.060 ;
        RECT 13.425 41.875 13.715 41.920 ;
        RECT 12.490 41.180 12.810 41.440 ;
        RECT 8.810 40.160 9.130 40.420 ;
        RECT 9.745 40.360 10.035 40.405 ;
        RECT 12.490 40.360 12.810 40.420 ;
        RECT 9.745 40.220 12.810 40.360 ;
        RECT 9.745 40.175 10.035 40.220 ;
        RECT 12.490 40.160 12.810 40.220 ;
        RECT 6.985 40.020 7.275 40.065 ;
        RECT 7.430 40.020 7.750 40.080 ;
        RECT 6.985 39.880 7.750 40.020 ;
        RECT 8.900 40.020 9.040 40.160 ;
        RECT 12.030 40.020 12.350 40.080 ;
        RECT 8.900 39.880 12.350 40.020 ;
        RECT 6.985 39.835 7.275 39.880 ;
        RECT 7.430 39.820 7.750 39.880 ;
        RECT 12.030 39.820 12.350 39.880 ;
        RECT 8.810 38.460 9.130 38.720 ;
        RECT 7.905 37.640 8.195 37.685 ;
        RECT 8.810 37.640 9.130 37.700 ;
        RECT 7.905 37.500 9.130 37.640 ;
        RECT 7.905 37.455 8.195 37.500 ;
        RECT 8.810 37.440 9.130 37.500 ;
        RECT 10.205 34.240 10.495 34.285 ;
        RECT 11.570 34.240 11.890 34.300 ;
        RECT 10.205 34.100 11.890 34.240 ;
        RECT 10.205 34.055 10.495 34.100 ;
        RECT 11.570 34.040 11.890 34.100 ;
        RECT 8.365 33.900 8.655 33.945 ;
        RECT 9.730 33.900 10.050 33.960 ;
        RECT 8.365 33.760 10.050 33.900 ;
        RECT 8.365 33.715 8.655 33.760 ;
        RECT 9.730 33.700 10.050 33.760 ;
        RECT 10.665 33.900 10.955 33.945 ;
        RECT 13.410 33.900 13.730 33.960 ;
        RECT 10.665 33.760 13.730 33.900 ;
        RECT 10.665 33.715 10.955 33.760 ;
        RECT 13.410 33.700 13.730 33.760 ;
        RECT 6.970 33.560 7.290 33.620 ;
        RECT 12.030 33.560 12.350 33.620 ;
        RECT 6.970 33.420 12.350 33.560 ;
        RECT 6.970 33.360 7.290 33.420 ;
        RECT 12.030 33.360 12.350 33.420 ;
        RECT 8.810 33.020 9.130 33.280 ;
        RECT 9.270 33.020 9.590 33.280 ;
        RECT 11.585 33.220 11.875 33.265 ;
        RECT 13.870 33.220 14.190 33.280 ;
        RECT 11.585 33.080 14.190 33.220 ;
        RECT 11.585 33.035 11.875 33.080 ;
        RECT 13.870 33.020 14.190 33.080 ;
        RECT 8.810 32.200 9.130 32.260 ;
        RECT 11.125 32.200 11.415 32.245 ;
        RECT 8.810 32.060 11.415 32.200 ;
        RECT 8.810 32.000 9.130 32.060 ;
        RECT 11.125 32.015 11.415 32.060 ;
        RECT 9.730 31.860 10.050 31.920 ;
        RECT 7.520 31.720 9.500 31.860 ;
        RECT 7.520 31.580 7.660 31.720 ;
        RECT 7.430 31.320 7.750 31.580 ;
        RECT 7.890 31.320 8.210 31.580 ;
        RECT 9.360 31.225 9.500 31.720 ;
        RECT 9.730 31.720 10.880 31.860 ;
        RECT 9.730 31.660 10.050 31.720 ;
        RECT 9.285 30.995 9.575 31.225 ;
        RECT 6.970 30.500 7.290 30.560 ;
        RECT 8.365 30.500 8.655 30.545 ;
        RECT 6.970 30.360 8.655 30.500 ;
        RECT 9.360 30.500 9.500 30.995 ;
        RECT 10.740 30.885 10.880 31.720 ;
        RECT 12.030 31.320 12.350 31.580 ;
        RECT 12.490 31.320 12.810 31.580 ;
        RECT 12.965 31.335 13.255 31.565 ;
        RECT 13.040 31.180 13.180 31.335 ;
        RECT 12.580 31.040 13.180 31.180 ;
        RECT 10.665 30.655 10.955 30.885 ;
        RECT 12.580 30.500 12.720 31.040 ;
        RECT 9.360 30.360 12.720 30.500 ;
        RECT 6.970 30.300 7.290 30.360 ;
        RECT 8.365 30.315 8.655 30.360 ;
        RECT 7.905 29.480 8.195 29.525 ;
        RECT 8.350 29.480 8.670 29.540 ;
        RECT 7.905 29.340 8.670 29.480 ;
        RECT 7.905 29.295 8.195 29.340 ;
        RECT 8.350 29.280 8.670 29.340 ;
        RECT 8.810 29.480 9.130 29.540 ;
        RECT 9.285 29.480 9.575 29.525 ;
        RECT 8.810 29.340 9.575 29.480 ;
        RECT 8.810 29.280 9.130 29.340 ;
        RECT 9.285 29.295 9.575 29.340 ;
        RECT 7.430 28.460 7.750 28.520 ;
        RECT 8.825 28.460 9.115 28.505 ;
        RECT 7.430 28.320 9.115 28.460 ;
        RECT 7.430 28.260 7.750 28.320 ;
        RECT 8.825 28.275 9.115 28.320 ;
        RECT 9.730 28.260 10.050 28.520 ;
        RECT 9.730 26.760 10.050 26.820 ;
        RECT 10.665 26.760 10.955 26.805 ;
        RECT 9.730 26.620 10.955 26.760 ;
        RECT 9.730 26.560 10.050 26.620 ;
        RECT 10.665 26.575 10.955 26.620 ;
        RECT 8.810 25.880 9.130 26.140 ;
        RECT 6.970 25.740 7.290 25.800 ;
        RECT 7.445 25.740 7.735 25.785 ;
        RECT 6.970 25.600 7.735 25.740 ;
        RECT 6.970 25.540 7.290 25.600 ;
        RECT 7.445 25.555 7.735 25.600 ;
        RECT 8.350 25.540 8.670 25.800 ;
        RECT 7.890 23.840 8.210 24.100 ;
        RECT 7.905 18.600 8.195 18.645 ;
        RECT 8.810 18.600 9.130 18.660 ;
        RECT 7.905 18.460 9.130 18.600 ;
        RECT 7.905 18.415 8.195 18.460 ;
        RECT 8.810 18.400 9.130 18.460 ;
        RECT 8.350 13.160 8.670 13.220 ;
        RECT 9.285 13.160 9.575 13.205 ;
        RECT 8.350 13.020 9.575 13.160 ;
        RECT 8.350 12.960 8.670 13.020 ;
        RECT 9.285 12.975 9.575 13.020 ;
        RECT 12.490 12.960 12.810 13.220 ;
        RECT 7.905 12.820 8.195 12.865 ;
        RECT 12.580 12.820 12.720 12.960 ;
        RECT 7.905 12.680 12.720 12.820 ;
        RECT 7.905 12.635 8.195 12.680 ;
      LAYER met2 ;
        RECT 8.840 97.250 9.100 97.570 ;
        RECT 12.520 97.250 12.780 97.570 ;
        RECT 8.380 95.550 8.640 95.870 ;
        RECT 8.440 93.570 8.580 95.550 ;
        RECT 7.520 93.430 8.580 93.570 ;
        RECT 7.000 84.670 7.260 84.990 ;
        RECT 7.520 84.730 7.660 93.430 ;
        RECT 7.920 92.830 8.180 93.150 ;
        RECT 7.980 85.410 8.120 92.830 ;
        RECT 7.980 85.270 8.580 85.410 ;
        RECT 7.060 75.130 7.200 84.670 ;
        RECT 7.520 84.590 8.120 84.730 ;
        RECT 7.460 82.970 7.720 83.290 ;
        RECT 7.520 80.570 7.660 82.970 ;
        RECT 7.980 80.570 8.120 84.590 ;
        RECT 8.440 83.290 8.580 85.270 ;
        RECT 8.380 82.970 8.640 83.290 ;
        RECT 7.460 80.250 7.720 80.570 ;
        RECT 7.920 80.250 8.180 80.570 ;
        RECT 7.460 79.570 7.720 79.890 ;
        RECT 7.000 74.810 7.260 75.130 ;
        RECT 7.520 67.650 7.660 79.570 ;
        RECT 8.900 78.610 9.040 97.250 ;
        RECT 11.600 96.230 11.860 96.550 ;
        RECT 7.980 78.470 9.040 78.610 ;
        RECT 7.980 75.130 8.120 78.470 ;
        RECT 7.920 74.810 8.180 75.130 ;
        RECT 8.840 74.470 9.100 74.790 ;
        RECT 8.380 73.790 8.640 74.110 ;
        RECT 7.920 72.090 8.180 72.410 ;
        RECT 7.460 67.330 7.720 67.650 ;
        RECT 7.460 52.030 7.720 52.350 ;
        RECT 7.520 47.590 7.660 52.030 ;
        RECT 7.980 47.930 8.120 72.090 ;
        RECT 8.440 47.930 8.580 73.790 ;
        RECT 8.900 59.490 9.040 74.470 ;
        RECT 11.660 72.410 11.800 96.230 ;
        RECT 12.060 79.910 12.320 80.230 ;
        RECT 12.120 78.530 12.260 79.910 ;
        RECT 12.580 79.550 12.720 97.250 ;
        RECT 31.840 95.890 32.100 96.210 ;
        RECT 31.900 80.570 32.040 95.890 ;
        RECT 41.500 95.550 41.760 95.870 ;
        RECT 31.840 80.250 32.100 80.570 ;
        RECT 12.980 79.910 13.240 80.230 ;
        RECT 12.520 79.230 12.780 79.550 ;
        RECT 12.060 78.210 12.320 78.530 ;
        RECT 12.060 74.470 12.320 74.790 ;
        RECT 12.120 73.090 12.260 74.470 ;
        RECT 12.580 74.110 12.720 79.230 ;
        RECT 13.040 75.130 13.180 79.910 ;
        RECT 13.900 79.230 14.160 79.550 ;
        RECT 12.980 74.810 13.240 75.130 ;
        RECT 12.520 73.790 12.780 74.110 ;
        RECT 12.060 72.770 12.320 73.090 ;
        RECT 11.600 72.090 11.860 72.410 ;
        RECT 11.600 71.070 11.860 71.390 ;
        RECT 11.660 61.190 11.800 71.070 ;
        RECT 11.600 60.870 11.860 61.190 ;
        RECT 12.060 60.190 12.320 60.510 ;
        RECT 12.120 59.490 12.260 60.190 ;
        RECT 8.840 59.170 9.100 59.490 ;
        RECT 12.060 59.170 12.320 59.490 ;
        RECT 12.520 57.810 12.780 58.130 ;
        RECT 12.580 56.770 12.720 57.810 ;
        RECT 12.520 56.450 12.780 56.770 ;
        RECT 7.920 47.610 8.180 47.930 ;
        RECT 8.380 47.610 8.640 47.930 ;
        RECT 7.460 47.270 7.720 47.590 ;
        RECT 7.980 44.610 8.120 47.610 ;
        RECT 7.520 44.470 8.120 44.610 ;
        RECT 7.520 40.110 7.660 44.470 ;
        RECT 7.920 43.870 8.180 44.190 ;
        RECT 7.980 43.170 8.120 43.870 ;
        RECT 7.920 42.850 8.180 43.170 ;
        RECT 8.440 42.830 8.580 47.610 ;
        RECT 12.060 47.270 12.320 47.590 ;
        RECT 13.040 47.330 13.180 74.810 ;
        RECT 13.960 71.730 14.100 79.230 ;
        RECT 16.200 73.790 16.460 74.110 ;
        RECT 16.260 73.090 16.400 73.790 ;
        RECT 16.200 72.770 16.460 73.090 ;
        RECT 13.900 71.410 14.160 71.730 ;
        RECT 41.560 61.190 41.700 95.550 ;
        RECT 13.900 60.870 14.160 61.190 ;
        RECT 41.500 60.870 41.760 61.190 ;
        RECT 13.960 59.490 14.100 60.870 ;
        RECT 13.900 59.170 14.160 59.490 ;
        RECT 14.820 58.150 15.080 58.470 ;
        RECT 14.880 55.490 15.020 58.150 ;
        RECT 12.120 43.170 12.260 47.270 ;
        RECT 12.580 47.190 13.180 47.330 ;
        RECT 13.960 55.350 15.020 55.490 ;
        RECT 12.060 42.850 12.320 43.170 ;
        RECT 8.380 42.570 8.640 42.830 ;
        RECT 8.380 42.510 9.040 42.570 ;
        RECT 8.440 42.430 9.040 42.510 ;
        RECT 12.580 42.490 12.720 47.190 ;
        RECT 12.980 46.590 13.240 46.910 ;
        RECT 13.040 43.170 13.180 46.590 ;
        RECT 12.980 42.850 13.240 43.170 ;
        RECT 13.440 42.850 13.700 43.170 ;
        RECT 8.380 41.830 8.640 42.150 ;
        RECT 7.460 39.790 7.720 40.110 ;
        RECT 7.000 33.330 7.260 33.650 ;
        RECT 7.060 30.590 7.200 33.330 ;
        RECT 7.520 31.610 7.660 39.790 ;
        RECT 7.460 31.290 7.720 31.610 ;
        RECT 7.920 31.290 8.180 31.610 ;
        RECT 7.000 30.270 7.260 30.590 ;
        RECT 7.060 25.830 7.200 30.270 ;
        RECT 7.520 28.550 7.660 31.290 ;
        RECT 7.460 28.230 7.720 28.550 ;
        RECT 7.000 25.510 7.260 25.830 ;
        RECT 7.980 24.130 8.120 31.290 ;
        RECT 8.440 29.570 8.580 41.830 ;
        RECT 8.900 40.450 9.040 42.430 ;
        RECT 12.520 42.170 12.780 42.490 ;
        RECT 12.580 41.890 12.720 42.170 ;
        RECT 11.660 41.750 12.720 41.890 ;
        RECT 8.840 40.130 9.100 40.450 ;
        RECT 8.840 38.430 9.100 38.750 ;
        RECT 8.900 37.730 9.040 38.430 ;
        RECT 8.840 37.410 9.100 37.730 ;
        RECT 11.660 34.330 11.800 41.750 ;
        RECT 12.520 41.150 12.780 41.470 ;
        RECT 12.580 40.450 12.720 41.150 ;
        RECT 12.520 40.130 12.780 40.450 ;
        RECT 12.060 39.790 12.320 40.110 ;
        RECT 11.600 34.010 11.860 34.330 ;
        RECT 9.760 33.670 10.020 33.990 ;
        RECT 8.840 32.990 9.100 33.310 ;
        RECT 9.300 32.990 9.560 33.310 ;
        RECT 8.900 32.290 9.040 32.990 ;
        RECT 8.840 31.970 9.100 32.290 ;
        RECT 9.360 31.010 9.500 32.990 ;
        RECT 9.820 31.950 9.960 33.670 ;
        RECT 12.120 33.650 12.260 39.790 ;
        RECT 13.500 33.990 13.640 42.850 ;
        RECT 13.440 33.670 13.700 33.990 ;
        RECT 12.060 33.330 12.320 33.650 ;
        RECT 9.760 31.630 10.020 31.950 ;
        RECT 12.120 31.610 12.260 33.330 ;
        RECT 13.960 33.310 14.100 55.350 ;
        RECT 13.900 32.990 14.160 33.310 ;
        RECT 12.060 31.290 12.320 31.610 ;
        RECT 12.520 31.290 12.780 31.610 ;
        RECT 8.900 30.870 9.500 31.010 ;
        RECT 8.900 29.570 9.040 30.870 ;
        RECT 8.380 29.250 8.640 29.570 ;
        RECT 8.840 29.250 9.100 29.570 ;
        RECT 9.760 28.230 10.020 28.550 ;
        RECT 9.820 26.850 9.960 28.230 ;
        RECT 9.760 26.530 10.020 26.850 ;
        RECT 8.840 25.850 9.100 26.170 ;
        RECT 8.380 25.510 8.640 25.830 ;
        RECT 7.920 23.810 8.180 24.130 ;
        RECT 8.440 13.250 8.580 25.510 ;
        RECT 8.900 18.690 9.040 25.850 ;
        RECT 8.840 18.370 9.100 18.690 ;
        RECT 12.580 13.250 12.720 31.290 ;
        RECT 8.380 12.930 8.640 13.250 ;
        RECT 12.520 12.930 12.780 13.250 ;
  END
END mux16x1_project
MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r2
  CLASS BLOCK ;
  FOREIGN sky130_osu_ring_oscillator_mpr2xa_8_b0r2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 104.095 BY 12.465 ;
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 32.740 8.240 32.910 9.510 ;
        RECT 38.355 8.240 38.525 9.510 ;
        RECT 38.355 2.955 38.525 4.225 ;
      LAYER met1 ;
        RECT 32.650 8.410 33.000 8.470 ;
        RECT 38.280 8.410 38.620 8.500 ;
        RECT 32.650 8.380 33.140 8.410 ;
        RECT 38.280 8.405 38.755 8.410 ;
        RECT 38.260 8.380 38.755 8.405 ;
        RECT 32.650 8.240 38.755 8.380 ;
        RECT 32.650 8.205 38.620 8.240 ;
        RECT 32.650 8.180 33.000 8.205 ;
        RECT 38.280 8.150 38.620 8.205 ;
        RECT 38.280 4.225 38.620 4.350 ;
        RECT 38.280 4.055 38.755 4.225 ;
        RECT 38.280 4.000 38.620 4.055 ;
      LAYER met2 ;
        RECT 32.680 8.135 32.970 8.515 ;
        RECT 38.280 8.150 38.620 8.500 ;
        RECT 38.360 4.350 38.530 8.150 ;
        RECT 38.280 4.000 38.620 4.350 ;
      LAYER met3 ;
        RECT 32.650 8.135 33.000 12.465 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 48.000 8.240 48.170 9.510 ;
        RECT 53.615 8.240 53.785 9.510 ;
        RECT 53.615 2.955 53.785 4.225 ;
      LAYER met1 ;
        RECT 47.910 8.410 48.260 8.470 ;
        RECT 53.540 8.410 53.880 8.500 ;
        RECT 47.910 8.380 48.400 8.410 ;
        RECT 53.540 8.405 54.015 8.410 ;
        RECT 53.520 8.380 54.015 8.405 ;
        RECT 47.910 8.240 54.015 8.380 ;
        RECT 47.910 8.205 53.880 8.240 ;
        RECT 47.910 8.180 48.260 8.205 ;
        RECT 53.540 8.150 53.880 8.205 ;
        RECT 53.540 4.225 53.880 4.350 ;
        RECT 53.540 4.055 54.015 4.225 ;
        RECT 53.540 4.000 53.880 4.055 ;
      LAYER met2 ;
        RECT 47.940 8.135 48.230 8.515 ;
        RECT 53.540 8.150 53.880 8.500 ;
        RECT 53.620 4.350 53.790 8.150 ;
        RECT 53.540 4.000 53.880 4.350 ;
      LAYER met3 ;
        RECT 47.910 8.135 48.260 12.465 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 63.260 8.240 63.430 9.510 ;
        RECT 68.875 8.240 69.045 9.510 ;
        RECT 68.875 2.955 69.045 4.225 ;
      LAYER met1 ;
        RECT 63.170 8.410 63.520 8.470 ;
        RECT 68.800 8.410 69.140 8.500 ;
        RECT 63.170 8.380 63.660 8.410 ;
        RECT 68.800 8.405 69.275 8.410 ;
        RECT 68.780 8.380 69.275 8.405 ;
        RECT 63.170 8.240 69.275 8.380 ;
        RECT 63.170 8.205 69.140 8.240 ;
        RECT 63.170 8.180 63.520 8.205 ;
        RECT 68.800 8.150 69.140 8.205 ;
        RECT 68.800 4.225 69.140 4.350 ;
        RECT 68.800 4.055 69.275 4.225 ;
        RECT 68.800 4.000 69.140 4.055 ;
      LAYER met2 ;
        RECT 63.200 8.135 63.490 8.515 ;
        RECT 68.800 8.150 69.140 8.500 ;
        RECT 68.880 4.350 69.050 8.150 ;
        RECT 68.800 4.000 69.140 4.350 ;
      LAYER met3 ;
        RECT 63.170 8.135 63.520 12.465 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 78.520 8.240 78.690 9.510 ;
        RECT 84.135 8.240 84.305 9.510 ;
        RECT 84.135 2.955 84.305 4.225 ;
      LAYER met1 ;
        RECT 78.430 8.410 78.780 8.470 ;
        RECT 84.060 8.410 84.400 8.500 ;
        RECT 78.430 8.380 78.920 8.410 ;
        RECT 84.060 8.405 84.535 8.410 ;
        RECT 84.040 8.380 84.535 8.405 ;
        RECT 78.430 8.240 84.535 8.380 ;
        RECT 78.430 8.205 84.400 8.240 ;
        RECT 78.430 8.180 78.780 8.205 ;
        RECT 84.060 8.150 84.400 8.205 ;
        RECT 84.060 4.225 84.400 4.350 ;
        RECT 84.060 4.055 84.535 4.225 ;
        RECT 84.060 4.000 84.400 4.055 ;
      LAYER met2 ;
        RECT 78.460 8.135 78.750 8.515 ;
        RECT 84.060 8.150 84.400 8.500 ;
        RECT 84.140 4.350 84.310 8.150 ;
        RECT 84.060 4.000 84.400 4.350 ;
      LAYER met3 ;
        RECT 78.430 8.135 78.780 12.465 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 93.780 8.240 93.950 9.510 ;
        RECT 99.395 8.240 99.565 9.510 ;
        RECT 99.395 2.955 99.565 4.225 ;
      LAYER met1 ;
        RECT 93.690 8.410 94.040 8.470 ;
        RECT 99.320 8.410 99.660 8.500 ;
        RECT 93.690 8.380 94.180 8.410 ;
        RECT 99.320 8.405 99.795 8.410 ;
        RECT 99.300 8.380 99.795 8.405 ;
        RECT 93.690 8.240 99.795 8.380 ;
        RECT 93.690 8.205 99.660 8.240 ;
        RECT 93.690 8.180 94.040 8.205 ;
        RECT 99.320 8.150 99.660 8.205 ;
        RECT 99.320 4.225 99.660 4.350 ;
        RECT 99.320 4.055 99.795 4.225 ;
        RECT 99.320 4.000 99.660 4.055 ;
      LAYER met2 ;
        RECT 93.720 8.135 94.010 8.515 ;
        RECT 99.320 8.150 99.660 8.500 ;
        RECT 99.400 4.350 99.570 8.150 ;
        RECT 99.320 4.000 99.660 4.350 ;
      LAYER met3 ;
        RECT 93.690 8.135 94.040 12.465 ;
    END
  END s5
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 42.505 4.010 42.680 5.155 ;
        RECT 42.505 3.575 42.675 4.010 ;
        RECT 42.510 1.865 42.680 2.375 ;
      LAYER met1 ;
        RECT 42.445 3.540 42.735 3.775 ;
        RECT 42.445 3.535 42.675 3.540 ;
        RECT 42.505 2.435 42.675 3.535 ;
        RECT 42.445 2.175 42.740 2.435 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 57.765 4.010 57.940 5.155 ;
        RECT 57.765 3.575 57.935 4.010 ;
        RECT 57.770 1.865 57.940 2.375 ;
      LAYER met1 ;
        RECT 57.705 3.540 57.995 3.775 ;
        RECT 57.705 3.535 57.935 3.540 ;
        RECT 57.765 2.435 57.935 3.535 ;
        RECT 57.705 2.175 58.000 2.435 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 73.025 4.010 73.200 5.155 ;
        RECT 73.025 3.575 73.195 4.010 ;
        RECT 73.030 1.865 73.200 2.375 ;
      LAYER met1 ;
        RECT 72.965 3.540 73.255 3.775 ;
        RECT 72.965 3.535 73.195 3.540 ;
        RECT 73.025 2.435 73.195 3.535 ;
        RECT 72.965 2.175 73.260 2.435 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 88.285 4.010 88.460 5.155 ;
        RECT 88.285 3.575 88.455 4.010 ;
        RECT 88.290 1.865 88.460 2.375 ;
      LAYER met1 ;
        RECT 88.225 3.540 88.515 3.775 ;
        RECT 88.225 3.535 88.455 3.540 ;
        RECT 88.285 2.435 88.455 3.535 ;
        RECT 88.225 2.175 88.520 2.435 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 103.545 4.010 103.720 5.155 ;
        RECT 103.545 3.575 103.715 4.010 ;
        RECT 103.550 1.865 103.720 2.375 ;
      LAYER met1 ;
        RECT 103.485 3.540 103.775 3.775 ;
        RECT 103.485 3.535 103.715 3.540 ;
        RECT 103.545 2.435 103.715 3.535 ;
        RECT 103.485 2.175 103.780 2.435 ;
    END
  END X5_Y1
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 25.225 8.240 25.395 9.510 ;
      LAYER met1 ;
        RECT 25.165 8.435 25.455 8.440 ;
        RECT 25.165 8.410 25.460 8.435 ;
        RECT 25.165 8.240 25.625 8.410 ;
        RECT 25.165 8.210 25.460 8.240 ;
        RECT 25.170 8.205 25.460 8.210 ;
    END
  END start
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 10.865 104.095 12.465 ;
        RECT 25.215 10.240 25.385 10.865 ;
        RECT 32.730 10.240 32.900 10.865 ;
        RECT 33.685 10.320 33.855 10.600 ;
        RECT 33.685 10.150 33.915 10.320 ;
        RECT 38.345 10.240 38.515 10.865 ;
        RECT 41.090 10.240 41.260 10.865 ;
        RECT 42.080 10.240 42.250 10.865 ;
        RECT 47.990 10.240 48.160 10.865 ;
        RECT 48.945 10.320 49.115 10.600 ;
        RECT 48.945 10.150 49.175 10.320 ;
        RECT 53.605 10.240 53.775 10.865 ;
        RECT 56.350 10.240 56.520 10.865 ;
        RECT 57.340 10.240 57.510 10.865 ;
        RECT 63.250 10.240 63.420 10.865 ;
        RECT 64.205 10.320 64.375 10.600 ;
        RECT 64.205 10.150 64.435 10.320 ;
        RECT 68.865 10.240 69.035 10.865 ;
        RECT 71.610 10.240 71.780 10.865 ;
        RECT 72.600 10.240 72.770 10.865 ;
        RECT 78.510 10.240 78.680 10.865 ;
        RECT 79.465 10.320 79.635 10.600 ;
        RECT 79.465 10.150 79.695 10.320 ;
        RECT 84.125 10.240 84.295 10.865 ;
        RECT 86.870 10.240 87.040 10.865 ;
        RECT 87.860 10.240 88.030 10.865 ;
        RECT 93.770 10.240 93.940 10.865 ;
        RECT 94.725 10.320 94.895 10.600 ;
        RECT 94.725 10.150 94.955 10.320 ;
        RECT 99.385 10.240 99.555 10.865 ;
        RECT 102.130 10.240 102.300 10.865 ;
        RECT 103.120 10.240 103.290 10.865 ;
        RECT 33.745 8.540 33.915 10.150 ;
        RECT 49.005 8.540 49.175 10.150 ;
        RECT 64.265 8.540 64.435 10.150 ;
        RECT 79.525 8.540 79.695 10.150 ;
        RECT 94.785 8.540 94.955 10.150 ;
        RECT 33.685 8.370 33.915 8.540 ;
        RECT 48.945 8.370 49.175 8.540 ;
        RECT 64.205 8.370 64.435 8.540 ;
        RECT 79.465 8.370 79.695 8.540 ;
        RECT 94.725 8.370 94.955 8.540 ;
        RECT 33.685 7.310 33.855 8.370 ;
        RECT 48.945 7.310 49.115 8.370 ;
        RECT 64.205 7.310 64.375 8.370 ;
        RECT 79.465 7.310 79.635 8.370 ;
        RECT 94.725 7.310 94.895 8.370 ;
      LAYER met1 ;
        RECT 0.000 10.865 104.095 12.465 ;
        RECT 33.515 8.820 33.685 10.865 ;
        RECT 48.775 8.820 48.945 10.865 ;
        RECT 64.035 8.820 64.205 10.865 ;
        RECT 79.295 8.820 79.465 10.865 ;
        RECT 94.555 8.820 94.725 10.865 ;
        RECT 33.515 8.790 33.975 8.820 ;
        RECT 48.775 8.790 49.235 8.820 ;
        RECT 64.035 8.790 64.495 8.820 ;
        RECT 79.295 8.790 79.755 8.820 ;
        RECT 94.555 8.790 95.015 8.820 ;
        RECT 33.510 8.620 33.975 8.790 ;
        RECT 48.770 8.620 49.235 8.790 ;
        RECT 64.030 8.620 64.495 8.790 ;
        RECT 79.290 8.620 79.755 8.790 ;
        RECT 94.550 8.620 95.015 8.790 ;
        RECT 33.515 8.605 33.975 8.620 ;
        RECT 48.775 8.605 49.235 8.620 ;
        RECT 64.035 8.605 64.495 8.620 ;
        RECT 79.295 8.605 79.755 8.620 ;
        RECT 94.555 8.605 95.015 8.620 ;
        RECT 33.685 8.590 33.975 8.605 ;
        RECT 48.945 8.590 49.235 8.605 ;
        RECT 64.205 8.590 64.495 8.605 ;
        RECT 79.465 8.590 79.755 8.605 ;
        RECT 94.725 8.590 95.015 8.605 ;
    END
    PORT
      LAYER li1 ;
        RECT 29.095 3.785 29.265 4.235 ;
        RECT 30.415 3.865 30.785 4.035 ;
        RECT 30.415 3.395 30.585 3.865 ;
        RECT 44.355 3.785 44.525 4.235 ;
        RECT 45.675 3.865 46.045 4.035 ;
        RECT 45.675 3.395 45.845 3.865 ;
        RECT 59.615 3.785 59.785 4.235 ;
        RECT 60.935 3.865 61.305 4.035 ;
        RECT 60.935 3.395 61.105 3.865 ;
        RECT 74.875 3.785 75.045 4.235 ;
        RECT 76.195 3.865 76.565 4.035 ;
        RECT 76.195 3.395 76.365 3.865 ;
        RECT 90.135 3.785 90.305 4.235 ;
        RECT 91.455 3.865 91.825 4.035 ;
        RECT 91.455 3.395 91.625 3.865 ;
        RECT 29.815 2.890 29.985 3.375 ;
        RECT 30.295 3.225 30.585 3.395 ;
        RECT 29.815 2.875 30.090 2.890 ;
        RECT 31.735 2.875 31.905 3.375 ;
        RECT 32.695 2.875 32.865 3.375 ;
        RECT 33.570 2.875 33.765 2.890 ;
        RECT 34.615 2.875 34.785 3.375 ;
        RECT 35.575 2.880 35.745 3.375 ;
        RECT 35.420 2.875 35.745 2.880 ;
        RECT 36.515 2.875 36.685 3.375 ;
        RECT 45.075 2.890 45.245 3.375 ;
        RECT 45.555 3.225 45.845 3.395 ;
        RECT 37.090 2.875 37.285 2.880 ;
        RECT 45.075 2.875 45.350 2.890 ;
        RECT 46.995 2.875 47.165 3.375 ;
        RECT 47.955 2.875 48.125 3.375 ;
        RECT 48.830 2.875 49.025 2.890 ;
        RECT 49.875 2.875 50.045 3.375 ;
        RECT 50.835 2.880 51.005 3.375 ;
        RECT 50.680 2.875 51.005 2.880 ;
        RECT 51.775 2.875 51.945 3.375 ;
        RECT 60.335 2.890 60.505 3.375 ;
        RECT 60.815 3.225 61.105 3.395 ;
        RECT 52.350 2.875 52.545 2.880 ;
        RECT 60.335 2.875 60.610 2.890 ;
        RECT 62.255 2.875 62.425 3.375 ;
        RECT 63.215 2.875 63.385 3.375 ;
        RECT 64.090 2.875 64.285 2.890 ;
        RECT 65.135 2.875 65.305 3.375 ;
        RECT 66.095 2.880 66.265 3.375 ;
        RECT 65.940 2.875 66.265 2.880 ;
        RECT 67.035 2.875 67.205 3.375 ;
        RECT 75.595 2.890 75.765 3.375 ;
        RECT 76.075 3.225 76.365 3.395 ;
        RECT 67.610 2.875 67.805 2.880 ;
        RECT 75.595 2.875 75.870 2.890 ;
        RECT 77.515 2.875 77.685 3.375 ;
        RECT 78.475 2.875 78.645 3.375 ;
        RECT 79.350 2.875 79.545 2.890 ;
        RECT 80.395 2.875 80.565 3.375 ;
        RECT 81.355 2.880 81.525 3.375 ;
        RECT 81.200 2.875 81.525 2.880 ;
        RECT 82.295 2.875 82.465 3.375 ;
        RECT 90.855 2.890 91.025 3.375 ;
        RECT 91.335 3.225 91.625 3.395 ;
        RECT 82.870 2.875 83.065 2.880 ;
        RECT 90.855 2.875 91.130 2.890 ;
        RECT 92.775 2.875 92.945 3.375 ;
        RECT 93.735 2.875 93.905 3.375 ;
        RECT 94.610 2.875 94.805 2.890 ;
        RECT 95.655 2.875 95.825 3.375 ;
        RECT 96.615 2.880 96.785 3.375 ;
        RECT 96.460 2.875 96.785 2.880 ;
        RECT 97.555 2.875 97.725 3.375 ;
        RECT 98.130 2.875 98.325 2.880 ;
        RECT 28.545 1.600 37.285 2.875 ;
        RECT 38.345 1.600 38.515 2.225 ;
        RECT 41.090 1.600 41.260 2.225 ;
        RECT 42.075 1.600 42.245 2.225 ;
        RECT 43.805 1.600 52.545 2.875 ;
        RECT 53.605 1.600 53.775 2.225 ;
        RECT 56.350 1.600 56.520 2.225 ;
        RECT 57.335 1.600 57.505 2.225 ;
        RECT 59.065 1.600 67.805 2.875 ;
        RECT 68.865 1.600 69.035 2.225 ;
        RECT 71.610 1.600 71.780 2.225 ;
        RECT 72.595 1.600 72.765 2.225 ;
        RECT 74.325 1.600 83.065 2.875 ;
        RECT 84.125 1.600 84.295 2.225 ;
        RECT 86.870 1.600 87.040 2.225 ;
        RECT 87.855 1.600 88.025 2.225 ;
        RECT 89.585 1.600 98.325 2.875 ;
        RECT 99.385 1.600 99.555 2.225 ;
        RECT 102.130 1.600 102.300 2.225 ;
        RECT 103.115 1.600 103.285 2.225 ;
        RECT 0.000 0.000 104.095 1.600 ;
      LAYER met1 ;
        RECT 29.035 4.035 29.325 4.265 ;
        RECT 44.295 4.035 44.585 4.265 ;
        RECT 59.555 4.035 59.845 4.265 ;
        RECT 74.815 4.035 75.105 4.265 ;
        RECT 90.075 4.035 90.365 4.265 ;
        RECT 29.105 3.805 29.245 4.035 ;
        RECT 44.365 3.805 44.505 4.035 ;
        RECT 59.625 3.805 59.765 4.035 ;
        RECT 74.885 3.805 75.025 4.035 ;
        RECT 90.145 3.805 90.285 4.035 ;
        RECT 29.105 3.665 29.725 3.805 ;
        RECT 44.365 3.665 44.985 3.805 ;
        RECT 59.625 3.665 60.245 3.805 ;
        RECT 74.885 3.665 75.505 3.805 ;
        RECT 90.145 3.665 90.765 3.805 ;
        RECT 29.585 3.505 29.725 3.665 ;
        RECT 44.845 3.505 44.985 3.665 ;
        RECT 60.105 3.505 60.245 3.665 ;
        RECT 75.365 3.505 75.505 3.665 ;
        RECT 90.625 3.505 90.765 3.665 ;
        RECT 29.345 3.445 29.725 3.505 ;
        RECT 44.605 3.445 44.985 3.505 ;
        RECT 59.865 3.445 60.245 3.505 ;
        RECT 75.125 3.445 75.505 3.505 ;
        RECT 90.385 3.445 90.765 3.505 ;
        RECT 29.345 3.385 29.935 3.445 ;
        RECT 30.235 3.385 30.525 3.425 ;
        RECT 29.345 3.245 30.525 3.385 ;
        RECT 44.605 3.385 45.195 3.445 ;
        RECT 45.495 3.385 45.785 3.425 ;
        RECT 44.605 3.245 45.785 3.385 ;
        RECT 59.865 3.385 60.455 3.445 ;
        RECT 60.755 3.385 61.045 3.425 ;
        RECT 59.865 3.245 61.045 3.385 ;
        RECT 75.125 3.385 75.715 3.445 ;
        RECT 76.015 3.385 76.305 3.425 ;
        RECT 75.125 3.245 76.305 3.385 ;
        RECT 90.385 3.385 90.975 3.445 ;
        RECT 91.275 3.385 91.565 3.425 ;
        RECT 90.385 3.245 91.565 3.385 ;
        RECT 29.530 3.185 29.935 3.245 ;
        RECT 30.235 3.195 30.525 3.245 ;
        RECT 44.790 3.185 45.195 3.245 ;
        RECT 45.495 3.195 45.785 3.245 ;
        RECT 60.050 3.185 60.455 3.245 ;
        RECT 60.755 3.195 61.045 3.245 ;
        RECT 75.310 3.185 75.715 3.245 ;
        RECT 76.015 3.195 76.305 3.245 ;
        RECT 90.570 3.185 90.975 3.245 ;
        RECT 91.275 3.195 91.565 3.245 ;
        RECT 29.530 2.915 29.820 3.185 ;
        RECT 44.790 2.915 45.080 3.185 ;
        RECT 60.050 2.915 60.340 3.185 ;
        RECT 75.310 2.915 75.600 3.185 ;
        RECT 90.570 2.915 90.860 3.185 ;
        RECT 28.545 1.600 37.285 2.915 ;
        RECT 43.805 1.600 52.545 2.915 ;
        RECT 59.065 1.600 67.805 2.915 ;
        RECT 74.325 1.600 83.065 2.915 ;
        RECT 89.585 1.600 98.325 2.915 ;
        RECT 0.000 0.000 104.095 1.600 ;
      LAYER met2 ;
        RECT 29.515 3.475 29.795 3.500 ;
        RECT 44.775 3.475 45.055 3.500 ;
        RECT 60.035 3.475 60.315 3.500 ;
        RECT 75.295 3.475 75.575 3.500 ;
        RECT 90.555 3.475 90.835 3.500 ;
        RECT 29.515 3.155 29.905 3.475 ;
        RECT 44.775 3.155 45.165 3.475 ;
        RECT 60.035 3.155 60.425 3.475 ;
        RECT 75.295 3.155 75.685 3.475 ;
        RECT 90.555 3.155 90.945 3.475 ;
        RECT 29.515 3.125 29.795 3.155 ;
        RECT 44.775 3.125 45.055 3.155 ;
        RECT 60.035 3.125 60.315 3.155 ;
        RECT 75.295 3.125 75.575 3.155 ;
        RECT 90.555 3.125 90.835 3.155 ;
      LAYER met3 ;
        RECT 29.475 3.475 29.830 3.480 ;
        RECT 44.735 3.475 45.090 3.480 ;
        RECT 59.995 3.475 60.350 3.480 ;
        RECT 75.255 3.475 75.610 3.480 ;
        RECT 90.515 3.475 90.870 3.480 ;
        RECT 29.375 3.145 30.105 3.475 ;
        RECT 44.635 3.145 45.365 3.475 ;
        RECT 59.895 3.145 60.625 3.475 ;
        RECT 75.155 3.145 75.885 3.475 ;
        RECT 90.415 3.145 91.145 3.475 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 24.995 8.745 27.805 8.750 ;
        RECT 32.510 8.745 35.320 8.750 ;
        RECT 38.125 8.745 42.905 8.750 ;
        RECT 47.770 8.745 50.580 8.750 ;
        RECT 53.385 8.745 58.165 8.750 ;
        RECT 63.030 8.745 65.840 8.750 ;
        RECT 68.645 8.745 73.425 8.750 ;
        RECT 78.290 8.745 81.100 8.750 ;
        RECT 83.905 8.745 88.685 8.750 ;
        RECT 93.550 8.745 96.360 8.750 ;
        RECT 99.165 8.745 103.945 8.750 ;
        RECT 24.995 6.660 104.095 8.745 ;
        RECT 25.000 5.095 104.095 6.660 ;
        RECT 25.010 4.100 104.095 5.095 ;
        RECT 27.795 4.095 104.095 4.100 ;
        RECT 37.105 3.720 43.055 4.095 ;
        RECT 52.365 3.720 58.315 4.095 ;
        RECT 67.625 3.720 73.575 4.095 ;
        RECT 82.885 3.720 88.835 4.095 ;
        RECT 98.145 3.720 104.095 4.095 ;
        RECT 38.125 3.715 42.900 3.720 ;
        RECT 53.385 3.715 58.160 3.720 ;
        RECT 68.645 3.715 73.420 3.720 ;
        RECT 83.905 3.715 88.680 3.720 ;
        RECT 99.165 3.715 103.940 3.720 ;
      LAYER li1 ;
        RECT 27.030 10.050 27.205 10.600 ;
        RECT 27.030 8.450 27.200 10.050 ;
        RECT 25.215 7.040 25.385 7.770 ;
        RECT 27.030 7.310 27.205 8.450 ;
        RECT 27.030 7.040 27.200 7.310 ;
        RECT 32.730 7.040 32.900 7.770 ;
        RECT 38.345 7.040 38.515 7.770 ;
        RECT 41.090 7.040 41.260 7.770 ;
        RECT 42.080 7.040 42.250 7.770 ;
        RECT 47.990 7.040 48.160 7.770 ;
        RECT 53.605 7.040 53.775 7.770 ;
        RECT 56.350 7.040 56.520 7.770 ;
        RECT 57.340 7.040 57.510 7.770 ;
        RECT 63.250 7.040 63.420 7.770 ;
        RECT 68.865 7.040 69.035 7.770 ;
        RECT 71.610 7.040 71.780 7.770 ;
        RECT 72.600 7.040 72.770 7.770 ;
        RECT 78.510 7.040 78.680 7.770 ;
        RECT 84.125 7.040 84.295 7.770 ;
        RECT 86.870 7.040 87.040 7.770 ;
        RECT 87.860 7.040 88.030 7.770 ;
        RECT 93.770 7.040 93.940 7.770 ;
        RECT 99.385 7.040 99.555 7.770 ;
        RECT 102.130 7.040 102.300 7.770 ;
        RECT 103.120 7.040 103.290 7.770 ;
        RECT 25.045 7.035 27.795 7.040 ;
        RECT 32.560 7.035 35.310 7.040 ;
        RECT 38.175 7.035 42.900 7.040 ;
        RECT 47.820 7.035 50.570 7.040 ;
        RECT 53.435 7.035 58.160 7.040 ;
        RECT 63.080 7.035 65.830 7.040 ;
        RECT 68.695 7.035 73.420 7.040 ;
        RECT 78.340 7.035 81.090 7.040 ;
        RECT 83.955 7.035 88.680 7.040 ;
        RECT 93.600 7.035 96.350 7.040 ;
        RECT 99.215 7.035 103.940 7.040 ;
        RECT 0.000 5.435 104.095 7.035 ;
        RECT 28.545 5.430 43.055 5.435 ;
        RECT 43.805 5.430 58.315 5.435 ;
        RECT 59.065 5.430 73.575 5.435 ;
        RECT 74.325 5.430 88.835 5.435 ;
        RECT 89.585 5.430 104.095 5.435 ;
        RECT 28.545 5.425 37.285 5.430 ;
        RECT 38.175 5.425 42.895 5.430 ;
        RECT 43.805 5.425 52.545 5.430 ;
        RECT 53.435 5.425 58.155 5.430 ;
        RECT 59.065 5.425 67.805 5.430 ;
        RECT 68.695 5.425 73.415 5.430 ;
        RECT 74.325 5.425 83.065 5.430 ;
        RECT 83.955 5.425 88.675 5.430 ;
        RECT 89.585 5.425 98.325 5.430 ;
        RECT 99.215 5.425 103.935 5.430 ;
        RECT 29.335 4.925 29.505 5.425 ;
        RECT 31.255 4.925 31.425 5.425 ;
        RECT 32.715 4.925 32.885 5.425 ;
        RECT 33.655 4.925 33.825 5.425 ;
        RECT 35.575 4.925 35.745 5.425 ;
        RECT 38.345 4.695 38.515 5.425 ;
        RECT 41.090 4.695 41.260 5.425 ;
        RECT 42.075 4.695 42.245 5.425 ;
        RECT 44.595 4.925 44.765 5.425 ;
        RECT 46.515 4.925 46.685 5.425 ;
        RECT 47.975 4.925 48.145 5.425 ;
        RECT 48.915 4.925 49.085 5.425 ;
        RECT 50.835 4.925 51.005 5.425 ;
        RECT 53.605 4.695 53.775 5.425 ;
        RECT 56.350 4.695 56.520 5.425 ;
        RECT 57.335 4.695 57.505 5.425 ;
        RECT 59.855 4.925 60.025 5.425 ;
        RECT 61.775 4.925 61.945 5.425 ;
        RECT 63.235 4.925 63.405 5.425 ;
        RECT 64.175 4.925 64.345 5.425 ;
        RECT 66.095 4.925 66.265 5.425 ;
        RECT 68.865 4.695 69.035 5.425 ;
        RECT 71.610 4.695 71.780 5.425 ;
        RECT 72.595 4.695 72.765 5.425 ;
        RECT 75.115 4.925 75.285 5.425 ;
        RECT 77.035 4.925 77.205 5.425 ;
        RECT 78.495 4.925 78.665 5.425 ;
        RECT 79.435 4.925 79.605 5.425 ;
        RECT 81.355 4.925 81.525 5.425 ;
        RECT 84.125 4.695 84.295 5.425 ;
        RECT 86.870 4.695 87.040 5.425 ;
        RECT 87.855 4.695 88.025 5.425 ;
        RECT 90.375 4.925 90.545 5.425 ;
        RECT 92.295 4.925 92.465 5.425 ;
        RECT 93.755 4.925 93.925 5.425 ;
        RECT 94.695 4.925 94.865 5.425 ;
        RECT 96.615 4.925 96.785 5.425 ;
        RECT 99.385 4.695 99.555 5.425 ;
        RECT 102.130 4.695 102.300 5.425 ;
        RECT 103.115 4.695 103.285 5.425 ;
      LAYER met1 ;
        RECT 26.970 9.150 27.260 9.180 ;
        RECT 26.800 8.980 27.260 9.150 ;
        RECT 26.970 8.950 27.260 8.980 ;
        RECT 25.045 7.035 27.795 7.040 ;
        RECT 32.560 7.035 35.310 7.040 ;
        RECT 38.175 7.035 42.900 7.040 ;
        RECT 47.820 7.035 50.570 7.040 ;
        RECT 53.435 7.035 58.160 7.040 ;
        RECT 63.080 7.035 65.830 7.040 ;
        RECT 68.695 7.035 73.420 7.040 ;
        RECT 78.340 7.035 81.090 7.040 ;
        RECT 83.955 7.035 88.680 7.040 ;
        RECT 93.600 7.035 96.350 7.040 ;
        RECT 99.215 7.035 103.940 7.040 ;
        RECT 0.000 5.435 104.095 7.035 ;
        RECT 28.545 5.430 43.055 5.435 ;
        RECT 43.805 5.430 58.315 5.435 ;
        RECT 59.065 5.430 73.575 5.435 ;
        RECT 74.325 5.430 88.835 5.435 ;
        RECT 89.585 5.430 104.095 5.435 ;
        RECT 28.545 5.395 37.285 5.430 ;
        RECT 38.175 5.425 42.895 5.430 ;
        RECT 43.805 5.395 52.545 5.430 ;
        RECT 53.435 5.425 58.155 5.430 ;
        RECT 59.065 5.395 67.805 5.430 ;
        RECT 68.695 5.425 73.415 5.430 ;
        RECT 74.325 5.395 83.065 5.430 ;
        RECT 83.955 5.425 88.675 5.430 ;
        RECT 89.585 5.395 98.325 5.430 ;
        RECT 99.215 5.425 103.935 5.430 ;
    END
  END vccd1
  OBS
      LAYER pwell ;
        RECT 28.925 2.715 29.095 2.875 ;
        RECT 44.185 2.715 44.355 2.875 ;
        RECT 59.445 2.715 59.615 2.875 ;
        RECT 74.705 2.715 74.875 2.875 ;
        RECT 89.965 2.715 90.135 2.875 ;
      LAYER li1 ;
        RECT 25.645 10.110 25.820 10.600 ;
        RECT 26.170 10.320 26.340 10.600 ;
        RECT 26.170 10.150 26.400 10.320 ;
        RECT 25.645 9.940 25.815 10.110 ;
        RECT 25.645 9.610 26.055 9.940 ;
        RECT 25.645 9.100 25.815 9.610 ;
        RECT 25.645 8.770 26.055 9.100 ;
        RECT 25.645 8.570 25.815 8.770 ;
        RECT 25.645 7.310 25.820 8.570 ;
        RECT 26.230 8.540 26.400 10.150 ;
        RECT 26.600 10.090 26.775 10.600 ;
        RECT 33.160 10.110 33.335 10.600 ;
        RECT 33.160 9.940 33.330 10.110 ;
        RECT 34.115 10.090 34.290 10.600 ;
        RECT 34.545 10.050 34.720 10.600 ;
        RECT 38.775 10.110 38.950 10.600 ;
        RECT 39.300 10.320 39.470 10.600 ;
        RECT 39.300 10.150 39.530 10.320 ;
        RECT 33.160 9.610 33.570 9.940 ;
        RECT 26.170 8.370 26.400 8.540 ;
        RECT 26.600 8.570 26.770 9.520 ;
        RECT 33.160 9.100 33.330 9.610 ;
        RECT 33.160 8.770 33.570 9.100 ;
        RECT 33.160 8.570 33.330 8.770 ;
        RECT 34.115 8.570 34.285 9.520 ;
        RECT 26.170 7.310 26.340 8.370 ;
        RECT 26.600 7.310 26.775 8.570 ;
        RECT 33.160 7.310 33.335 8.570 ;
        RECT 34.115 7.310 34.290 8.570 ;
        RECT 34.545 8.450 34.715 10.050 ;
        RECT 38.775 9.940 38.945 10.110 ;
        RECT 38.775 9.610 39.185 9.940 ;
        RECT 38.775 9.100 38.945 9.610 ;
        RECT 38.775 8.770 39.185 9.100 ;
        RECT 38.775 8.570 38.945 8.770 ;
        RECT 34.545 7.310 34.720 8.450 ;
        RECT 38.775 7.310 38.950 8.570 ;
        RECT 39.360 8.540 39.530 10.150 ;
        RECT 39.730 10.090 39.905 10.600 ;
        RECT 40.160 10.050 40.335 10.600 ;
        RECT 41.525 10.090 41.695 10.600 ;
        RECT 42.515 10.090 42.685 10.600 ;
        RECT 48.420 10.110 48.595 10.600 ;
        RECT 39.300 8.370 39.530 8.540 ;
        RECT 39.730 8.570 39.900 9.520 ;
        RECT 39.300 7.310 39.470 8.370 ;
        RECT 39.730 7.310 39.905 8.570 ;
        RECT 40.160 8.450 40.330 10.050 ;
        RECT 48.420 9.940 48.590 10.110 ;
        RECT 49.375 10.090 49.550 10.600 ;
        RECT 49.805 10.050 49.980 10.600 ;
        RECT 54.035 10.110 54.210 10.600 ;
        RECT 54.560 10.320 54.730 10.600 ;
        RECT 54.560 10.150 54.790 10.320 ;
        RECT 48.420 9.610 48.830 9.940 ;
        RECT 41.090 9.430 41.320 9.585 ;
        RECT 41.090 9.355 41.620 9.430 ;
        RECT 41.150 9.260 41.620 9.355 ;
        RECT 42.140 9.260 42.610 9.430 ;
        RECT 41.150 8.570 41.320 9.260 ;
        RECT 41.520 8.810 41.690 8.890 ;
        RECT 42.140 8.810 42.310 9.260 ;
        RECT 48.420 9.100 48.590 9.610 ;
        RECT 41.520 8.610 42.310 8.810 ;
        RECT 40.160 7.310 40.335 8.450 ;
        RECT 41.520 7.310 41.695 8.610 ;
        RECT 42.140 8.570 42.310 8.610 ;
        RECT 42.510 8.455 42.680 8.890 ;
        RECT 48.420 8.770 48.830 9.100 ;
        RECT 48.420 8.570 48.590 8.770 ;
        RECT 49.375 8.570 49.545 9.520 ;
        RECT 42.510 7.310 42.685 8.455 ;
        RECT 48.420 7.310 48.595 8.570 ;
        RECT 49.375 7.310 49.550 8.570 ;
        RECT 49.805 8.450 49.975 10.050 ;
        RECT 54.035 9.940 54.205 10.110 ;
        RECT 54.035 9.610 54.445 9.940 ;
        RECT 54.035 9.100 54.205 9.610 ;
        RECT 54.035 8.770 54.445 9.100 ;
        RECT 54.035 8.570 54.205 8.770 ;
        RECT 49.805 7.310 49.980 8.450 ;
        RECT 54.035 7.310 54.210 8.570 ;
        RECT 54.620 8.540 54.790 10.150 ;
        RECT 54.990 10.090 55.165 10.600 ;
        RECT 55.420 10.050 55.595 10.600 ;
        RECT 56.785 10.090 56.955 10.600 ;
        RECT 57.775 10.090 57.945 10.600 ;
        RECT 63.680 10.110 63.855 10.600 ;
        RECT 54.560 8.370 54.790 8.540 ;
        RECT 54.990 8.570 55.160 9.520 ;
        RECT 54.560 7.310 54.730 8.370 ;
        RECT 54.990 7.310 55.165 8.570 ;
        RECT 55.420 8.450 55.590 10.050 ;
        RECT 63.680 9.940 63.850 10.110 ;
        RECT 64.635 10.090 64.810 10.600 ;
        RECT 65.065 10.050 65.240 10.600 ;
        RECT 69.295 10.110 69.470 10.600 ;
        RECT 69.820 10.320 69.990 10.600 ;
        RECT 69.820 10.150 70.050 10.320 ;
        RECT 63.680 9.610 64.090 9.940 ;
        RECT 56.350 9.430 56.580 9.585 ;
        RECT 56.350 9.355 56.880 9.430 ;
        RECT 56.410 9.260 56.880 9.355 ;
        RECT 57.400 9.260 57.870 9.430 ;
        RECT 56.410 8.570 56.580 9.260 ;
        RECT 56.780 8.810 56.950 8.890 ;
        RECT 57.400 8.810 57.570 9.260 ;
        RECT 63.680 9.100 63.850 9.610 ;
        RECT 56.780 8.610 57.570 8.810 ;
        RECT 55.420 7.310 55.595 8.450 ;
        RECT 56.780 7.310 56.955 8.610 ;
        RECT 57.400 8.570 57.570 8.610 ;
        RECT 57.770 8.455 57.940 8.890 ;
        RECT 63.680 8.770 64.090 9.100 ;
        RECT 63.680 8.570 63.850 8.770 ;
        RECT 64.635 8.570 64.805 9.520 ;
        RECT 57.770 7.310 57.945 8.455 ;
        RECT 63.680 7.310 63.855 8.570 ;
        RECT 64.635 7.310 64.810 8.570 ;
        RECT 65.065 8.450 65.235 10.050 ;
        RECT 69.295 9.940 69.465 10.110 ;
        RECT 69.295 9.610 69.705 9.940 ;
        RECT 69.295 9.100 69.465 9.610 ;
        RECT 69.295 8.770 69.705 9.100 ;
        RECT 69.295 8.570 69.465 8.770 ;
        RECT 65.065 7.310 65.240 8.450 ;
        RECT 69.295 7.310 69.470 8.570 ;
        RECT 69.880 8.540 70.050 10.150 ;
        RECT 70.250 10.090 70.425 10.600 ;
        RECT 70.680 10.050 70.855 10.600 ;
        RECT 72.045 10.090 72.215 10.600 ;
        RECT 73.035 10.090 73.205 10.600 ;
        RECT 78.940 10.110 79.115 10.600 ;
        RECT 69.820 8.370 70.050 8.540 ;
        RECT 70.250 8.570 70.420 9.520 ;
        RECT 69.820 7.310 69.990 8.370 ;
        RECT 70.250 7.310 70.425 8.570 ;
        RECT 70.680 8.450 70.850 10.050 ;
        RECT 78.940 9.940 79.110 10.110 ;
        RECT 79.895 10.090 80.070 10.600 ;
        RECT 80.325 10.050 80.500 10.600 ;
        RECT 84.555 10.110 84.730 10.600 ;
        RECT 85.080 10.320 85.250 10.600 ;
        RECT 85.080 10.150 85.310 10.320 ;
        RECT 78.940 9.610 79.350 9.940 ;
        RECT 71.610 9.430 71.840 9.585 ;
        RECT 71.610 9.355 72.140 9.430 ;
        RECT 71.670 9.260 72.140 9.355 ;
        RECT 72.660 9.260 73.130 9.430 ;
        RECT 71.670 8.570 71.840 9.260 ;
        RECT 72.040 8.810 72.210 8.890 ;
        RECT 72.660 8.810 72.830 9.260 ;
        RECT 78.940 9.100 79.110 9.610 ;
        RECT 72.040 8.610 72.830 8.810 ;
        RECT 70.680 7.310 70.855 8.450 ;
        RECT 72.040 7.310 72.215 8.610 ;
        RECT 72.660 8.570 72.830 8.610 ;
        RECT 73.030 8.455 73.200 8.890 ;
        RECT 78.940 8.770 79.350 9.100 ;
        RECT 78.940 8.570 79.110 8.770 ;
        RECT 79.895 8.570 80.065 9.520 ;
        RECT 73.030 7.310 73.205 8.455 ;
        RECT 78.940 7.310 79.115 8.570 ;
        RECT 79.895 7.310 80.070 8.570 ;
        RECT 80.325 8.450 80.495 10.050 ;
        RECT 84.555 9.940 84.725 10.110 ;
        RECT 84.555 9.610 84.965 9.940 ;
        RECT 84.555 9.100 84.725 9.610 ;
        RECT 84.555 8.770 84.965 9.100 ;
        RECT 84.555 8.570 84.725 8.770 ;
        RECT 80.325 7.310 80.500 8.450 ;
        RECT 84.555 7.310 84.730 8.570 ;
        RECT 85.140 8.540 85.310 10.150 ;
        RECT 85.510 10.090 85.685 10.600 ;
        RECT 85.940 10.050 86.115 10.600 ;
        RECT 87.305 10.090 87.475 10.600 ;
        RECT 88.295 10.090 88.465 10.600 ;
        RECT 94.200 10.110 94.375 10.600 ;
        RECT 85.080 8.370 85.310 8.540 ;
        RECT 85.510 8.570 85.680 9.520 ;
        RECT 85.080 7.310 85.250 8.370 ;
        RECT 85.510 7.310 85.685 8.570 ;
        RECT 85.940 8.450 86.110 10.050 ;
        RECT 94.200 9.940 94.370 10.110 ;
        RECT 95.155 10.090 95.330 10.600 ;
        RECT 95.585 10.050 95.760 10.600 ;
        RECT 99.815 10.110 99.990 10.600 ;
        RECT 100.340 10.320 100.510 10.600 ;
        RECT 100.340 10.150 100.570 10.320 ;
        RECT 94.200 9.610 94.610 9.940 ;
        RECT 86.870 9.430 87.100 9.585 ;
        RECT 86.870 9.355 87.400 9.430 ;
        RECT 86.930 9.260 87.400 9.355 ;
        RECT 87.920 9.260 88.390 9.430 ;
        RECT 86.930 8.570 87.100 9.260 ;
        RECT 87.300 8.810 87.470 8.890 ;
        RECT 87.920 8.810 88.090 9.260 ;
        RECT 94.200 9.100 94.370 9.610 ;
        RECT 87.300 8.610 88.090 8.810 ;
        RECT 85.940 7.310 86.115 8.450 ;
        RECT 87.300 7.310 87.475 8.610 ;
        RECT 87.920 8.570 88.090 8.610 ;
        RECT 88.290 8.455 88.460 8.890 ;
        RECT 94.200 8.770 94.610 9.100 ;
        RECT 94.200 8.570 94.370 8.770 ;
        RECT 95.155 8.570 95.325 9.520 ;
        RECT 88.290 7.310 88.465 8.455 ;
        RECT 94.200 7.310 94.375 8.570 ;
        RECT 95.155 7.310 95.330 8.570 ;
        RECT 95.585 8.450 95.755 10.050 ;
        RECT 99.815 9.940 99.985 10.110 ;
        RECT 99.815 9.610 100.225 9.940 ;
        RECT 99.815 9.100 99.985 9.610 ;
        RECT 99.815 8.770 100.225 9.100 ;
        RECT 99.815 8.570 99.985 8.770 ;
        RECT 95.585 7.310 95.760 8.450 ;
        RECT 99.815 7.310 99.990 8.570 ;
        RECT 100.400 8.540 100.570 10.150 ;
        RECT 100.770 10.090 100.945 10.600 ;
        RECT 101.200 10.050 101.375 10.600 ;
        RECT 102.565 10.090 102.735 10.600 ;
        RECT 103.555 10.090 103.725 10.600 ;
        RECT 100.340 8.370 100.570 8.540 ;
        RECT 100.770 8.570 100.940 9.520 ;
        RECT 100.340 7.310 100.510 8.370 ;
        RECT 100.770 7.310 100.945 8.570 ;
        RECT 101.200 8.450 101.370 10.050 ;
        RECT 102.130 9.430 102.360 9.585 ;
        RECT 102.130 9.355 102.660 9.430 ;
        RECT 102.190 9.260 102.660 9.355 ;
        RECT 103.180 9.260 103.650 9.430 ;
        RECT 102.190 8.570 102.360 9.260 ;
        RECT 102.560 8.810 102.730 8.890 ;
        RECT 103.180 8.810 103.350 9.260 ;
        RECT 102.560 8.610 103.350 8.810 ;
        RECT 101.200 7.310 101.375 8.450 ;
        RECT 102.560 7.310 102.735 8.610 ;
        RECT 103.180 8.570 103.350 8.610 ;
        RECT 103.550 8.455 103.720 8.890 ;
        RECT 103.550 7.310 103.725 8.455 ;
        RECT 28.875 4.435 29.045 4.795 ;
        RECT 29.815 4.435 29.985 4.795 ;
        RECT 30.295 4.345 30.465 4.765 ;
        RECT 30.655 4.515 30.945 5.075 ;
        RECT 31.735 4.775 31.905 5.105 ;
        RECT 32.215 4.685 32.385 5.075 ;
        RECT 34.110 4.775 34.285 5.105 ;
        RECT 36.055 4.905 36.565 5.075 ;
        RECT 34.635 4.685 34.815 4.795 ;
        RECT 36.395 4.765 36.565 4.905 ;
        RECT 32.105 4.515 32.440 4.685 ;
        RECT 32.935 4.515 33.425 4.685 ;
        RECT 34.635 4.515 35.985 4.685 ;
        RECT 36.395 4.515 36.680 4.765 ;
        RECT 30.775 4.435 30.945 4.515 ;
        RECT 29.575 3.785 29.745 4.235 ;
        RECT 30.055 3.785 30.225 4.115 ;
        RECT 31.015 3.785 31.185 4.115 ;
        RECT 31.495 3.785 31.665 4.515 ;
        RECT 32.935 4.345 33.105 4.515 ;
        RECT 34.635 4.435 34.815 4.515 ;
        RECT 35.815 4.345 35.985 4.515 ;
        RECT 36.505 4.435 36.680 4.515 ;
        RECT 31.975 3.785 32.145 4.235 ;
        RECT 32.455 3.785 32.625 4.115 ;
        RECT 32.935 3.785 33.105 4.115 ;
        RECT 33.415 3.785 33.585 4.235 ;
        RECT 34.375 4.135 34.545 4.235 ;
        RECT 33.895 4.035 34.545 4.135 ;
        RECT 33.815 3.865 34.625 4.035 ;
        RECT 34.855 3.785 35.025 4.115 ;
        RECT 35.335 3.785 35.505 4.235 ;
        RECT 35.815 3.785 35.985 4.115 ;
        RECT 36.295 4.035 36.565 4.235 ;
        RECT 36.175 3.825 36.565 4.035 ;
        RECT 38.775 3.895 38.950 5.155 ;
        RECT 39.300 4.095 39.470 5.155 ;
        RECT 39.300 3.925 39.530 4.095 ;
        RECT 38.775 3.695 38.945 3.895 ;
        RECT 33.895 3.615 34.065 3.655 ;
        RECT 33.535 3.445 34.065 3.615 ;
        RECT 28.875 3.045 29.045 3.395 ;
        RECT 30.775 3.045 30.945 3.395 ;
        RECT 32.175 3.375 32.345 3.395 ;
        RECT 32.175 3.345 32.385 3.375 ;
        RECT 32.075 3.125 32.385 3.345 ;
        RECT 32.215 3.045 32.385 3.125 ;
        RECT 33.175 3.275 33.345 3.395 ;
        RECT 33.175 3.105 34.415 3.275 ;
        RECT 35.095 3.045 35.265 3.395 ;
        RECT 36.055 3.045 36.225 3.395 ;
        RECT 38.775 3.365 39.185 3.695 ;
        RECT 38.775 2.855 38.945 3.365 ;
        RECT 38.775 2.525 39.185 2.855 ;
        RECT 38.775 2.355 38.945 2.525 ;
        RECT 38.775 1.865 38.950 2.355 ;
        RECT 39.360 2.315 39.530 3.925 ;
        RECT 39.730 3.895 39.905 5.155 ;
        RECT 40.160 4.015 40.335 5.155 ;
        RECT 39.730 2.945 39.900 3.895 ;
        RECT 40.160 2.415 40.330 4.015 ;
        RECT 41.520 4.010 41.695 5.155 ;
        RECT 44.135 4.435 44.305 4.795 ;
        RECT 45.075 4.435 45.245 4.795 ;
        RECT 45.555 4.345 45.725 4.765 ;
        RECT 45.915 4.515 46.205 5.075 ;
        RECT 46.995 4.775 47.165 5.105 ;
        RECT 47.475 4.685 47.645 5.075 ;
        RECT 49.370 4.775 49.545 5.105 ;
        RECT 51.315 4.905 51.825 5.075 ;
        RECT 49.895 4.685 50.075 4.795 ;
        RECT 51.655 4.765 51.825 4.905 ;
        RECT 47.365 4.515 47.700 4.685 ;
        RECT 48.195 4.515 48.685 4.685 ;
        RECT 49.895 4.515 51.245 4.685 ;
        RECT 51.655 4.515 51.940 4.765 ;
        RECT 46.035 4.435 46.205 4.515 ;
        RECT 41.150 3.205 41.320 3.895 ;
        RECT 41.520 3.820 41.690 4.010 ;
        RECT 42.135 3.820 42.305 3.895 ;
        RECT 41.520 3.625 42.305 3.820 ;
        RECT 44.835 3.785 45.005 4.235 ;
        RECT 45.315 3.785 45.485 4.115 ;
        RECT 46.275 3.785 46.445 4.115 ;
        RECT 46.755 3.785 46.925 4.515 ;
        RECT 48.195 4.345 48.365 4.515 ;
        RECT 49.895 4.435 50.075 4.515 ;
        RECT 51.075 4.345 51.245 4.515 ;
        RECT 51.765 4.435 51.940 4.515 ;
        RECT 47.235 3.785 47.405 4.235 ;
        RECT 47.715 3.785 47.885 4.115 ;
        RECT 48.195 3.785 48.365 4.115 ;
        RECT 48.675 3.785 48.845 4.235 ;
        RECT 49.635 4.135 49.805 4.235 ;
        RECT 49.155 4.035 49.805 4.135 ;
        RECT 49.075 3.865 49.885 4.035 ;
        RECT 50.115 3.785 50.285 4.115 ;
        RECT 50.595 3.785 50.765 4.235 ;
        RECT 51.075 3.785 51.245 4.115 ;
        RECT 51.555 4.035 51.825 4.235 ;
        RECT 51.435 3.825 51.825 4.035 ;
        RECT 54.035 3.895 54.210 5.155 ;
        RECT 54.560 4.095 54.730 5.155 ;
        RECT 54.560 3.925 54.790 4.095 ;
        RECT 54.035 3.695 54.205 3.895 ;
        RECT 41.520 3.575 41.690 3.625 ;
        RECT 42.135 3.205 42.305 3.625 ;
        RECT 49.155 3.615 49.325 3.655 ;
        RECT 48.795 3.445 49.325 3.615 ;
        RECT 41.150 3.170 41.620 3.205 ;
        RECT 41.090 3.035 41.620 3.170 ;
        RECT 42.135 3.035 42.605 3.205 ;
        RECT 44.135 3.045 44.305 3.395 ;
        RECT 46.035 3.045 46.205 3.395 ;
        RECT 47.435 3.375 47.605 3.395 ;
        RECT 47.435 3.345 47.645 3.375 ;
        RECT 47.335 3.125 47.645 3.345 ;
        RECT 47.475 3.045 47.645 3.125 ;
        RECT 48.435 3.275 48.605 3.395 ;
        RECT 48.435 3.105 49.675 3.275 ;
        RECT 50.355 3.045 50.525 3.395 ;
        RECT 51.315 3.045 51.485 3.395 ;
        RECT 54.035 3.365 54.445 3.695 ;
        RECT 41.090 2.940 41.320 3.035 ;
        RECT 54.035 2.855 54.205 3.365 ;
        RECT 54.035 2.525 54.445 2.855 ;
        RECT 39.300 2.145 39.530 2.315 ;
        RECT 39.300 1.865 39.470 2.145 ;
        RECT 39.730 1.865 39.905 2.375 ;
        RECT 40.160 1.865 40.335 2.415 ;
        RECT 41.525 1.865 41.695 2.375 ;
        RECT 54.035 2.355 54.205 2.525 ;
        RECT 54.035 1.865 54.210 2.355 ;
        RECT 54.620 2.315 54.790 3.925 ;
        RECT 54.990 3.895 55.165 5.155 ;
        RECT 55.420 4.015 55.595 5.155 ;
        RECT 54.990 2.945 55.160 3.895 ;
        RECT 55.420 2.415 55.590 4.015 ;
        RECT 56.780 4.010 56.955 5.155 ;
        RECT 59.395 4.435 59.565 4.795 ;
        RECT 60.335 4.435 60.505 4.795 ;
        RECT 60.815 4.345 60.985 4.765 ;
        RECT 61.175 4.515 61.465 5.075 ;
        RECT 62.255 4.775 62.425 5.105 ;
        RECT 62.735 4.685 62.905 5.075 ;
        RECT 64.630 4.775 64.805 5.105 ;
        RECT 66.575 4.905 67.085 5.075 ;
        RECT 65.155 4.685 65.335 4.795 ;
        RECT 66.915 4.765 67.085 4.905 ;
        RECT 62.625 4.515 62.960 4.685 ;
        RECT 63.455 4.515 63.945 4.685 ;
        RECT 65.155 4.515 66.505 4.685 ;
        RECT 66.915 4.515 67.200 4.765 ;
        RECT 61.295 4.435 61.465 4.515 ;
        RECT 56.410 3.205 56.580 3.895 ;
        RECT 56.780 3.820 56.950 4.010 ;
        RECT 57.395 3.820 57.565 3.895 ;
        RECT 56.780 3.625 57.565 3.820 ;
        RECT 60.095 3.785 60.265 4.235 ;
        RECT 60.575 3.785 60.745 4.115 ;
        RECT 61.535 3.785 61.705 4.115 ;
        RECT 62.015 3.785 62.185 4.515 ;
        RECT 63.455 4.345 63.625 4.515 ;
        RECT 65.155 4.435 65.335 4.515 ;
        RECT 66.335 4.345 66.505 4.515 ;
        RECT 67.025 4.435 67.200 4.515 ;
        RECT 62.495 3.785 62.665 4.235 ;
        RECT 62.975 3.785 63.145 4.115 ;
        RECT 63.455 3.785 63.625 4.115 ;
        RECT 63.935 3.785 64.105 4.235 ;
        RECT 64.895 4.135 65.065 4.235 ;
        RECT 64.415 4.035 65.065 4.135 ;
        RECT 64.335 3.865 65.145 4.035 ;
        RECT 65.375 3.785 65.545 4.115 ;
        RECT 65.855 3.785 66.025 4.235 ;
        RECT 66.335 3.785 66.505 4.115 ;
        RECT 66.815 4.035 67.085 4.235 ;
        RECT 66.695 3.825 67.085 4.035 ;
        RECT 69.295 3.895 69.470 5.155 ;
        RECT 69.820 4.095 69.990 5.155 ;
        RECT 69.820 3.925 70.050 4.095 ;
        RECT 69.295 3.695 69.465 3.895 ;
        RECT 56.780 3.575 56.950 3.625 ;
        RECT 57.395 3.205 57.565 3.625 ;
        RECT 64.415 3.615 64.585 3.655 ;
        RECT 64.055 3.445 64.585 3.615 ;
        RECT 56.410 3.170 56.880 3.205 ;
        RECT 56.350 3.035 56.880 3.170 ;
        RECT 57.395 3.035 57.865 3.205 ;
        RECT 59.395 3.045 59.565 3.395 ;
        RECT 61.295 3.045 61.465 3.395 ;
        RECT 62.695 3.375 62.865 3.395 ;
        RECT 62.695 3.345 62.905 3.375 ;
        RECT 62.595 3.125 62.905 3.345 ;
        RECT 62.735 3.045 62.905 3.125 ;
        RECT 63.695 3.275 63.865 3.395 ;
        RECT 63.695 3.105 64.935 3.275 ;
        RECT 65.615 3.045 65.785 3.395 ;
        RECT 66.575 3.045 66.745 3.395 ;
        RECT 69.295 3.365 69.705 3.695 ;
        RECT 56.350 2.940 56.580 3.035 ;
        RECT 69.295 2.855 69.465 3.365 ;
        RECT 69.295 2.525 69.705 2.855 ;
        RECT 54.560 2.145 54.790 2.315 ;
        RECT 54.560 1.865 54.730 2.145 ;
        RECT 54.990 1.865 55.165 2.375 ;
        RECT 55.420 1.865 55.595 2.415 ;
        RECT 56.785 1.865 56.955 2.375 ;
        RECT 69.295 2.355 69.465 2.525 ;
        RECT 69.295 1.865 69.470 2.355 ;
        RECT 69.880 2.315 70.050 3.925 ;
        RECT 70.250 3.895 70.425 5.155 ;
        RECT 70.680 4.015 70.855 5.155 ;
        RECT 70.250 2.945 70.420 3.895 ;
        RECT 70.680 2.415 70.850 4.015 ;
        RECT 72.040 4.010 72.215 5.155 ;
        RECT 74.655 4.435 74.825 4.795 ;
        RECT 75.595 4.435 75.765 4.795 ;
        RECT 76.075 4.345 76.245 4.765 ;
        RECT 76.435 4.515 76.725 5.075 ;
        RECT 77.515 4.775 77.685 5.105 ;
        RECT 77.995 4.685 78.165 5.075 ;
        RECT 79.890 4.775 80.065 5.105 ;
        RECT 81.835 4.905 82.345 5.075 ;
        RECT 80.415 4.685 80.595 4.795 ;
        RECT 82.175 4.765 82.345 4.905 ;
        RECT 77.885 4.515 78.220 4.685 ;
        RECT 78.715 4.515 79.205 4.685 ;
        RECT 80.415 4.515 81.765 4.685 ;
        RECT 82.175 4.515 82.460 4.765 ;
        RECT 76.555 4.435 76.725 4.515 ;
        RECT 71.670 3.205 71.840 3.895 ;
        RECT 72.040 3.820 72.210 4.010 ;
        RECT 72.655 3.820 72.825 3.895 ;
        RECT 72.040 3.625 72.825 3.820 ;
        RECT 75.355 3.785 75.525 4.235 ;
        RECT 75.835 3.785 76.005 4.115 ;
        RECT 76.795 3.785 76.965 4.115 ;
        RECT 77.275 3.785 77.445 4.515 ;
        RECT 78.715 4.345 78.885 4.515 ;
        RECT 80.415 4.435 80.595 4.515 ;
        RECT 81.595 4.345 81.765 4.515 ;
        RECT 82.285 4.435 82.460 4.515 ;
        RECT 77.755 3.785 77.925 4.235 ;
        RECT 78.235 3.785 78.405 4.115 ;
        RECT 78.715 3.785 78.885 4.115 ;
        RECT 79.195 3.785 79.365 4.235 ;
        RECT 80.155 4.135 80.325 4.235 ;
        RECT 79.675 4.035 80.325 4.135 ;
        RECT 79.595 3.865 80.405 4.035 ;
        RECT 80.635 3.785 80.805 4.115 ;
        RECT 81.115 3.785 81.285 4.235 ;
        RECT 81.595 3.785 81.765 4.115 ;
        RECT 82.075 4.035 82.345 4.235 ;
        RECT 81.955 3.825 82.345 4.035 ;
        RECT 84.555 3.895 84.730 5.155 ;
        RECT 85.080 4.095 85.250 5.155 ;
        RECT 85.080 3.925 85.310 4.095 ;
        RECT 84.555 3.695 84.725 3.895 ;
        RECT 72.040 3.575 72.210 3.625 ;
        RECT 72.655 3.205 72.825 3.625 ;
        RECT 79.675 3.615 79.845 3.655 ;
        RECT 79.315 3.445 79.845 3.615 ;
        RECT 71.670 3.170 72.140 3.205 ;
        RECT 71.610 3.035 72.140 3.170 ;
        RECT 72.655 3.035 73.125 3.205 ;
        RECT 74.655 3.045 74.825 3.395 ;
        RECT 76.555 3.045 76.725 3.395 ;
        RECT 77.955 3.375 78.125 3.395 ;
        RECT 77.955 3.345 78.165 3.375 ;
        RECT 77.855 3.125 78.165 3.345 ;
        RECT 77.995 3.045 78.165 3.125 ;
        RECT 78.955 3.275 79.125 3.395 ;
        RECT 78.955 3.105 80.195 3.275 ;
        RECT 80.875 3.045 81.045 3.395 ;
        RECT 81.835 3.045 82.005 3.395 ;
        RECT 84.555 3.365 84.965 3.695 ;
        RECT 71.610 2.940 71.840 3.035 ;
        RECT 84.555 2.855 84.725 3.365 ;
        RECT 84.555 2.525 84.965 2.855 ;
        RECT 69.820 2.145 70.050 2.315 ;
        RECT 69.820 1.865 69.990 2.145 ;
        RECT 70.250 1.865 70.425 2.375 ;
        RECT 70.680 1.865 70.855 2.415 ;
        RECT 72.045 1.865 72.215 2.375 ;
        RECT 84.555 2.355 84.725 2.525 ;
        RECT 84.555 1.865 84.730 2.355 ;
        RECT 85.140 2.315 85.310 3.925 ;
        RECT 85.510 3.895 85.685 5.155 ;
        RECT 85.940 4.015 86.115 5.155 ;
        RECT 85.510 2.945 85.680 3.895 ;
        RECT 85.940 2.415 86.110 4.015 ;
        RECT 87.300 4.010 87.475 5.155 ;
        RECT 89.915 4.435 90.085 4.795 ;
        RECT 90.855 4.435 91.025 4.795 ;
        RECT 91.335 4.345 91.505 4.765 ;
        RECT 91.695 4.515 91.985 5.075 ;
        RECT 92.775 4.775 92.945 5.105 ;
        RECT 93.255 4.685 93.425 5.075 ;
        RECT 95.150 4.775 95.325 5.105 ;
        RECT 97.095 4.905 97.605 5.075 ;
        RECT 95.675 4.685 95.855 4.795 ;
        RECT 97.435 4.765 97.605 4.905 ;
        RECT 93.145 4.515 93.480 4.685 ;
        RECT 93.975 4.515 94.465 4.685 ;
        RECT 95.675 4.515 97.025 4.685 ;
        RECT 97.435 4.515 97.720 4.765 ;
        RECT 91.815 4.435 91.985 4.515 ;
        RECT 86.930 3.205 87.100 3.895 ;
        RECT 87.300 3.820 87.470 4.010 ;
        RECT 87.915 3.820 88.085 3.895 ;
        RECT 87.300 3.625 88.085 3.820 ;
        RECT 90.615 3.785 90.785 4.235 ;
        RECT 91.095 3.785 91.265 4.115 ;
        RECT 92.055 3.785 92.225 4.115 ;
        RECT 92.535 3.785 92.705 4.515 ;
        RECT 93.975 4.345 94.145 4.515 ;
        RECT 95.675 4.435 95.855 4.515 ;
        RECT 96.855 4.345 97.025 4.515 ;
        RECT 97.545 4.435 97.720 4.515 ;
        RECT 93.015 3.785 93.185 4.235 ;
        RECT 93.495 3.785 93.665 4.115 ;
        RECT 93.975 3.785 94.145 4.115 ;
        RECT 94.455 3.785 94.625 4.235 ;
        RECT 95.415 4.135 95.585 4.235 ;
        RECT 94.935 4.035 95.585 4.135 ;
        RECT 94.855 3.865 95.665 4.035 ;
        RECT 95.895 3.785 96.065 4.115 ;
        RECT 96.375 3.785 96.545 4.235 ;
        RECT 96.855 3.785 97.025 4.115 ;
        RECT 97.335 4.035 97.605 4.235 ;
        RECT 97.215 3.825 97.605 4.035 ;
        RECT 99.815 3.895 99.990 5.155 ;
        RECT 100.340 4.095 100.510 5.155 ;
        RECT 100.340 3.925 100.570 4.095 ;
        RECT 99.815 3.695 99.985 3.895 ;
        RECT 87.300 3.575 87.470 3.625 ;
        RECT 87.915 3.205 88.085 3.625 ;
        RECT 94.935 3.615 95.105 3.655 ;
        RECT 94.575 3.445 95.105 3.615 ;
        RECT 86.930 3.170 87.400 3.205 ;
        RECT 86.870 3.035 87.400 3.170 ;
        RECT 87.915 3.035 88.385 3.205 ;
        RECT 89.915 3.045 90.085 3.395 ;
        RECT 91.815 3.045 91.985 3.395 ;
        RECT 93.215 3.375 93.385 3.395 ;
        RECT 93.215 3.345 93.425 3.375 ;
        RECT 93.115 3.125 93.425 3.345 ;
        RECT 93.255 3.045 93.425 3.125 ;
        RECT 94.215 3.275 94.385 3.395 ;
        RECT 94.215 3.105 95.455 3.275 ;
        RECT 96.135 3.045 96.305 3.395 ;
        RECT 97.095 3.045 97.265 3.395 ;
        RECT 99.815 3.365 100.225 3.695 ;
        RECT 86.870 2.940 87.100 3.035 ;
        RECT 99.815 2.855 99.985 3.365 ;
        RECT 99.815 2.525 100.225 2.855 ;
        RECT 85.080 2.145 85.310 2.315 ;
        RECT 85.080 1.865 85.250 2.145 ;
        RECT 85.510 1.865 85.685 2.375 ;
        RECT 85.940 1.865 86.115 2.415 ;
        RECT 87.305 1.865 87.475 2.375 ;
        RECT 99.815 2.355 99.985 2.525 ;
        RECT 99.815 1.865 99.990 2.355 ;
        RECT 100.400 2.315 100.570 3.925 ;
        RECT 100.770 3.895 100.945 5.155 ;
        RECT 101.200 4.015 101.375 5.155 ;
        RECT 100.770 2.945 100.940 3.895 ;
        RECT 101.200 2.415 101.370 4.015 ;
        RECT 102.560 4.010 102.735 5.155 ;
        RECT 102.190 3.205 102.360 3.895 ;
        RECT 102.560 3.820 102.730 4.010 ;
        RECT 103.175 3.820 103.345 3.895 ;
        RECT 102.560 3.625 103.345 3.820 ;
        RECT 102.560 3.575 102.730 3.625 ;
        RECT 103.175 3.205 103.345 3.625 ;
        RECT 102.190 3.170 102.660 3.205 ;
        RECT 102.130 3.035 102.660 3.170 ;
        RECT 103.175 3.035 103.645 3.205 ;
        RECT 102.130 2.940 102.360 3.035 ;
        RECT 100.340 2.145 100.570 2.315 ;
        RECT 100.340 1.865 100.510 2.145 ;
        RECT 100.770 1.865 100.945 2.375 ;
        RECT 101.200 1.865 101.375 2.415 ;
        RECT 102.565 1.865 102.735 2.375 ;
      LAYER met1 ;
        RECT 26.540 10.060 26.830 10.290 ;
        RECT 34.055 10.060 34.345 10.290 ;
        RECT 39.670 10.060 39.960 10.290 ;
        RECT 26.600 9.610 26.770 10.060 ;
        RECT 34.115 9.715 34.285 10.060 ;
        RECT 26.510 9.320 26.860 9.610 ;
        RECT 34.015 9.345 34.385 9.715 ;
        RECT 39.730 9.580 39.900 10.060 ;
        RECT 41.460 10.030 41.755 10.290 ;
        RECT 42.450 10.030 42.745 10.290 ;
        RECT 49.315 10.060 49.605 10.290 ;
        RECT 54.930 10.060 55.220 10.290 ;
        RECT 41.090 9.630 41.320 9.645 ;
        RECT 41.045 9.580 41.355 9.630 ;
        RECT 39.730 9.550 41.355 9.580 ;
        RECT 39.670 9.410 41.355 9.550 ;
        RECT 34.055 9.320 34.345 9.345 ;
        RECT 39.670 9.320 39.960 9.410 ;
        RECT 41.045 9.320 41.355 9.410 ;
        RECT 41.090 9.290 41.320 9.320 ;
        RECT 34.685 9.180 35.035 9.245 ;
        RECT 40.125 9.180 40.450 9.270 ;
        RECT 34.485 9.150 35.035 9.180 ;
        RECT 40.100 9.150 40.450 9.180 ;
        RECT 34.315 9.145 35.035 9.150 ;
        RECT 39.930 9.145 40.450 9.150 ;
        RECT 34.315 8.980 40.450 9.145 ;
        RECT 34.375 8.975 40.450 8.980 ;
        RECT 34.485 8.950 35.035 8.975 ;
        RECT 40.100 8.950 40.450 8.975 ;
        RECT 34.685 8.895 35.035 8.950 ;
        RECT 40.125 8.945 40.450 8.950 ;
        RECT 41.520 8.930 41.690 10.030 ;
        RECT 42.510 9.300 42.680 10.030 ;
        RECT 49.375 9.715 49.545 10.060 ;
        RECT 49.275 9.345 49.645 9.715 ;
        RECT 54.990 9.580 55.160 10.060 ;
        RECT 56.720 10.030 57.015 10.290 ;
        RECT 57.710 10.030 58.005 10.290 ;
        RECT 64.575 10.060 64.865 10.290 ;
        RECT 70.190 10.060 70.480 10.290 ;
        RECT 56.350 9.630 56.580 9.645 ;
        RECT 56.305 9.580 56.615 9.630 ;
        RECT 54.990 9.550 56.615 9.580 ;
        RECT 54.930 9.410 56.615 9.550 ;
        RECT 49.315 9.320 49.605 9.345 ;
        RECT 54.930 9.320 55.220 9.410 ;
        RECT 56.305 9.320 56.615 9.410 ;
        RECT 42.505 8.950 42.855 9.300 ;
        RECT 56.350 9.290 56.580 9.320 ;
        RECT 49.945 9.180 50.295 9.255 ;
        RECT 55.385 9.180 55.710 9.270 ;
        RECT 49.745 9.150 50.295 9.180 ;
        RECT 55.360 9.150 55.710 9.180 ;
        RECT 49.575 9.145 50.295 9.150 ;
        RECT 55.190 9.145 55.710 9.150 ;
        RECT 49.575 8.980 55.710 9.145 ;
        RECT 49.635 8.975 55.710 8.980 ;
        RECT 49.745 8.950 50.295 8.975 ;
        RECT 55.360 8.950 55.710 8.975 ;
        RECT 42.505 8.930 42.800 8.950 ;
        RECT 41.460 8.925 41.690 8.930 ;
        RECT 26.135 8.790 26.485 8.865 ;
        RECT 39.325 8.820 39.645 8.835 ;
        RECT 39.300 8.790 39.645 8.820 ;
        RECT 25.995 8.620 26.485 8.790 ;
        RECT 39.125 8.620 39.645 8.790 ;
        RECT 41.460 8.690 41.750 8.925 ;
        RECT 42.450 8.860 42.800 8.930 ;
        RECT 49.945 8.905 50.295 8.950 ;
        RECT 55.385 8.945 55.710 8.950 ;
        RECT 56.780 8.930 56.950 10.030 ;
        RECT 57.770 9.305 57.940 10.030 ;
        RECT 64.635 9.715 64.805 10.060 ;
        RECT 64.535 9.345 64.905 9.715 ;
        RECT 70.250 9.580 70.420 10.060 ;
        RECT 71.980 10.030 72.275 10.290 ;
        RECT 72.970 10.030 73.265 10.290 ;
        RECT 79.835 10.060 80.125 10.290 ;
        RECT 85.450 10.060 85.740 10.290 ;
        RECT 71.610 9.630 71.840 9.645 ;
        RECT 71.565 9.580 71.875 9.630 ;
        RECT 70.250 9.550 71.875 9.580 ;
        RECT 70.190 9.410 71.875 9.550 ;
        RECT 64.575 9.320 64.865 9.345 ;
        RECT 70.190 9.320 70.480 9.410 ;
        RECT 71.565 9.320 71.875 9.410 ;
        RECT 57.760 8.950 58.115 9.305 ;
        RECT 71.610 9.290 71.840 9.320 ;
        RECT 65.205 9.180 65.555 9.255 ;
        RECT 70.645 9.180 70.970 9.270 ;
        RECT 65.005 9.150 65.555 9.180 ;
        RECT 70.620 9.150 70.970 9.180 ;
        RECT 64.835 9.145 65.555 9.150 ;
        RECT 70.450 9.145 70.970 9.150 ;
        RECT 64.835 8.980 70.970 9.145 ;
        RECT 64.895 8.975 70.970 8.980 ;
        RECT 65.005 8.950 65.555 8.975 ;
        RECT 70.620 8.950 70.970 8.975 ;
        RECT 57.760 8.930 58.060 8.950 ;
        RECT 56.720 8.925 56.950 8.930 ;
        RECT 42.450 8.690 42.740 8.860 ;
        RECT 54.585 8.820 54.905 8.835 ;
        RECT 54.560 8.790 54.905 8.820 ;
        RECT 54.385 8.620 54.905 8.790 ;
        RECT 56.720 8.690 57.010 8.925 ;
        RECT 57.710 8.865 58.060 8.930 ;
        RECT 65.205 8.905 65.555 8.950 ;
        RECT 70.645 8.945 70.970 8.950 ;
        RECT 72.040 8.930 72.210 10.030 ;
        RECT 73.030 9.300 73.200 10.030 ;
        RECT 79.895 9.715 80.065 10.060 ;
        RECT 79.795 9.345 80.165 9.715 ;
        RECT 85.510 9.580 85.680 10.060 ;
        RECT 87.240 10.030 87.535 10.290 ;
        RECT 88.230 10.030 88.525 10.290 ;
        RECT 95.095 10.060 95.385 10.290 ;
        RECT 100.710 10.060 101.000 10.290 ;
        RECT 86.870 9.630 87.100 9.645 ;
        RECT 86.825 9.580 87.135 9.630 ;
        RECT 85.510 9.550 87.135 9.580 ;
        RECT 85.450 9.410 87.135 9.550 ;
        RECT 79.835 9.320 80.125 9.345 ;
        RECT 85.450 9.320 85.740 9.410 ;
        RECT 86.825 9.320 87.135 9.410 ;
        RECT 72.980 8.950 73.330 9.300 ;
        RECT 86.870 9.290 87.100 9.320 ;
        RECT 80.470 9.180 80.820 9.255 ;
        RECT 85.905 9.180 86.230 9.270 ;
        RECT 80.265 9.150 80.820 9.180 ;
        RECT 85.880 9.150 86.230 9.180 ;
        RECT 80.095 9.145 80.820 9.150 ;
        RECT 85.710 9.145 86.230 9.150 ;
        RECT 80.095 8.980 86.230 9.145 ;
        RECT 80.155 8.975 86.230 8.980 ;
        RECT 80.265 8.950 80.820 8.975 ;
        RECT 85.880 8.950 86.230 8.975 ;
        RECT 72.980 8.930 73.320 8.950 ;
        RECT 71.980 8.925 72.210 8.930 ;
        RECT 57.710 8.690 58.000 8.865 ;
        RECT 69.845 8.820 70.165 8.835 ;
        RECT 69.820 8.790 70.165 8.820 ;
        RECT 69.645 8.620 70.165 8.790 ;
        RECT 71.980 8.690 72.270 8.925 ;
        RECT 72.970 8.860 73.320 8.930 ;
        RECT 80.470 8.905 80.820 8.950 ;
        RECT 85.905 8.945 86.230 8.950 ;
        RECT 87.300 8.930 87.470 10.030 ;
        RECT 88.290 9.300 88.460 10.030 ;
        RECT 95.155 9.715 95.325 10.060 ;
        RECT 95.055 9.345 95.425 9.715 ;
        RECT 100.770 9.580 100.940 10.060 ;
        RECT 102.500 10.030 102.795 10.290 ;
        RECT 103.490 10.030 103.785 10.290 ;
        RECT 102.130 9.630 102.360 9.645 ;
        RECT 102.085 9.580 102.395 9.630 ;
        RECT 100.770 9.550 102.395 9.580 ;
        RECT 100.710 9.410 102.395 9.550 ;
        RECT 95.095 9.320 95.385 9.345 ;
        RECT 100.710 9.320 101.000 9.410 ;
        RECT 102.085 9.320 102.395 9.410 ;
        RECT 88.240 8.950 88.590 9.300 ;
        RECT 102.130 9.290 102.360 9.320 ;
        RECT 95.725 9.180 96.075 9.255 ;
        RECT 101.165 9.180 101.490 9.270 ;
        RECT 95.525 9.150 96.075 9.180 ;
        RECT 101.140 9.150 101.490 9.180 ;
        RECT 95.355 9.145 96.075 9.150 ;
        RECT 100.970 9.145 101.490 9.150 ;
        RECT 95.355 8.980 101.490 9.145 ;
        RECT 95.415 8.975 101.490 8.980 ;
        RECT 95.525 8.950 96.075 8.975 ;
        RECT 101.140 8.950 101.490 8.975 ;
        RECT 88.240 8.930 88.580 8.950 ;
        RECT 87.240 8.925 87.470 8.930 ;
        RECT 72.970 8.690 73.260 8.860 ;
        RECT 85.105 8.820 85.425 8.835 ;
        RECT 85.080 8.790 85.425 8.820 ;
        RECT 84.905 8.620 85.425 8.790 ;
        RECT 87.240 8.690 87.530 8.925 ;
        RECT 88.230 8.860 88.580 8.930 ;
        RECT 95.725 8.905 96.075 8.950 ;
        RECT 101.165 8.945 101.490 8.950 ;
        RECT 102.560 8.930 102.730 10.030 ;
        RECT 103.525 9.995 103.785 10.030 ;
        RECT 103.525 9.915 103.845 9.995 ;
        RECT 103.525 9.565 103.875 9.915 ;
        RECT 103.550 8.930 103.720 9.565 ;
        RECT 102.500 8.925 102.730 8.930 ;
        RECT 103.490 8.925 103.720 8.930 ;
        RECT 88.230 8.690 88.520 8.860 ;
        RECT 100.365 8.820 100.685 8.835 ;
        RECT 100.340 8.790 100.685 8.820 ;
        RECT 100.165 8.620 100.685 8.790 ;
        RECT 102.500 8.690 102.790 8.925 ;
        RECT 103.490 8.690 103.780 8.925 ;
        RECT 26.135 8.575 26.485 8.620 ;
        RECT 39.300 8.590 39.645 8.620 ;
        RECT 54.560 8.590 54.905 8.620 ;
        RECT 69.820 8.590 70.165 8.620 ;
        RECT 85.080 8.590 85.425 8.620 ;
        RECT 100.340 8.590 100.685 8.620 ;
        RECT 39.325 8.545 39.645 8.590 ;
        RECT 54.585 8.545 54.905 8.590 ;
        RECT 69.845 8.545 70.165 8.590 ;
        RECT 85.105 8.545 85.425 8.590 ;
        RECT 100.365 8.545 100.685 8.590 ;
        RECT 30.715 4.895 31.005 5.105 ;
        RECT 29.825 4.875 31.005 4.895 ;
        RECT 28.805 4.585 29.125 4.845 ;
        RECT 29.825 4.825 30.925 4.875 ;
        RECT 31.655 4.865 31.975 5.125 ;
        RECT 32.255 5.105 32.575 5.125 ;
        RECT 32.155 4.875 32.575 5.105 ;
        RECT 32.255 4.865 32.575 4.875 ;
        RECT 33.815 5.105 34.150 5.125 ;
        RECT 33.815 4.875 34.340 5.105 ;
        RECT 35.995 5.065 36.285 5.105 ;
        RECT 36.425 5.065 36.745 5.125 ;
        RECT 35.995 4.925 36.745 5.065 ;
        RECT 35.995 4.875 36.285 4.925 ;
        RECT 33.815 4.865 34.150 4.875 ;
        RECT 36.425 4.865 36.745 4.925 ;
        RECT 45.975 4.895 46.265 5.105 ;
        RECT 45.085 4.875 46.265 4.895 ;
        RECT 29.755 4.755 30.925 4.825 ;
        RECT 29.755 4.595 30.045 4.755 ;
        RECT 32.185 4.585 32.355 4.685 ;
        RECT 34.565 4.585 34.885 4.845 ;
        RECT 44.065 4.585 44.385 4.845 ;
        RECT 45.085 4.825 46.185 4.875 ;
        RECT 46.915 4.865 47.235 5.125 ;
        RECT 47.515 5.105 47.835 5.125 ;
        RECT 47.415 4.875 47.835 5.105 ;
        RECT 47.515 4.865 47.835 4.875 ;
        RECT 49.075 5.105 49.410 5.125 ;
        RECT 49.075 4.875 49.600 5.105 ;
        RECT 51.255 5.065 51.545 5.105 ;
        RECT 51.685 5.065 52.005 5.125 ;
        RECT 51.255 4.925 52.005 5.065 ;
        RECT 51.255 4.875 51.545 4.925 ;
        RECT 49.075 4.865 49.410 4.875 ;
        RECT 51.685 4.865 52.005 4.925 ;
        RECT 61.235 4.895 61.525 5.105 ;
        RECT 60.345 4.875 61.525 4.895 ;
        RECT 45.015 4.755 46.185 4.825 ;
        RECT 45.015 4.595 45.305 4.755 ;
        RECT 47.445 4.585 47.615 4.685 ;
        RECT 49.825 4.585 50.145 4.845 ;
        RECT 59.325 4.585 59.645 4.845 ;
        RECT 60.345 4.825 61.445 4.875 ;
        RECT 62.175 4.865 62.495 5.125 ;
        RECT 62.775 5.105 63.095 5.125 ;
        RECT 62.675 4.875 63.095 5.105 ;
        RECT 62.775 4.865 63.095 4.875 ;
        RECT 64.335 5.105 64.670 5.125 ;
        RECT 64.335 4.875 64.860 5.105 ;
        RECT 66.515 5.065 66.805 5.105 ;
        RECT 66.945 5.065 67.265 5.125 ;
        RECT 66.515 4.925 67.265 5.065 ;
        RECT 66.515 4.875 66.805 4.925 ;
        RECT 64.335 4.865 64.670 4.875 ;
        RECT 66.945 4.865 67.265 4.925 ;
        RECT 76.495 4.895 76.785 5.105 ;
        RECT 75.605 4.875 76.785 4.895 ;
        RECT 60.275 4.755 61.445 4.825 ;
        RECT 60.275 4.595 60.565 4.755 ;
        RECT 62.705 4.585 62.875 4.685 ;
        RECT 65.085 4.585 65.405 4.845 ;
        RECT 74.585 4.585 74.905 4.845 ;
        RECT 75.605 4.825 76.705 4.875 ;
        RECT 77.435 4.865 77.755 5.125 ;
        RECT 78.035 5.105 78.355 5.125 ;
        RECT 77.935 4.875 78.355 5.105 ;
        RECT 78.035 4.865 78.355 4.875 ;
        RECT 79.595 5.105 79.930 5.125 ;
        RECT 79.595 4.875 80.120 5.105 ;
        RECT 81.775 5.065 82.065 5.105 ;
        RECT 82.205 5.065 82.525 5.125 ;
        RECT 81.775 4.925 82.525 5.065 ;
        RECT 81.775 4.875 82.065 4.925 ;
        RECT 79.595 4.865 79.930 4.875 ;
        RECT 82.205 4.865 82.525 4.925 ;
        RECT 91.755 4.895 92.045 5.105 ;
        RECT 90.865 4.875 92.045 4.895 ;
        RECT 75.535 4.755 76.705 4.825 ;
        RECT 75.535 4.595 75.825 4.755 ;
        RECT 77.965 4.585 78.135 4.685 ;
        RECT 80.345 4.585 80.665 4.845 ;
        RECT 89.845 4.585 90.165 4.845 ;
        RECT 90.865 4.825 91.965 4.875 ;
        RECT 92.695 4.865 93.015 5.125 ;
        RECT 93.295 5.105 93.615 5.125 ;
        RECT 93.195 4.875 93.615 5.105 ;
        RECT 93.295 4.865 93.615 4.875 ;
        RECT 94.855 5.105 95.190 5.125 ;
        RECT 94.855 4.875 95.380 5.105 ;
        RECT 97.035 5.065 97.325 5.105 ;
        RECT 97.465 5.065 97.785 5.125 ;
        RECT 97.035 4.925 97.785 5.065 ;
        RECT 97.035 4.875 97.325 4.925 ;
        RECT 94.855 4.865 95.190 4.875 ;
        RECT 97.465 4.865 97.785 4.925 ;
        RECT 90.795 4.755 91.965 4.825 ;
        RECT 90.795 4.595 91.085 4.755 ;
        RECT 93.225 4.585 93.395 4.685 ;
        RECT 95.605 4.585 95.925 4.845 ;
        RECT 31.175 4.545 31.495 4.565 ;
        RECT 30.235 4.505 30.525 4.545 ;
        RECT 30.235 4.315 30.685 4.505 ;
        RECT 29.495 4.025 29.815 4.285 ;
        RECT 29.975 3.745 30.295 4.005 ;
        RECT 30.545 3.985 30.685 4.315 ;
        RECT 31.175 4.315 31.725 4.545 ;
        RECT 31.865 4.445 34.045 4.585 ;
        RECT 46.435 4.545 46.755 4.565 ;
        RECT 31.865 4.365 33.165 4.445 ;
        RECT 31.175 4.305 31.495 4.315 ;
        RECT 31.865 4.085 32.205 4.365 ;
        RECT 32.875 4.315 33.165 4.365 ;
        RECT 31.915 4.035 32.205 4.085 ;
        RECT 33.335 4.025 33.655 4.285 ;
        RECT 30.545 3.845 30.805 3.985 ;
        RECT 28.805 3.185 29.125 3.445 ;
        RECT 30.665 3.425 30.805 3.845 ;
        RECT 30.955 3.945 31.245 3.985 ;
        RECT 31.415 3.945 31.735 4.005 ;
        RECT 30.955 3.805 31.735 3.945 ;
        RECT 30.955 3.755 31.245 3.805 ;
        RECT 31.415 3.745 31.735 3.805 ;
        RECT 32.395 3.755 32.685 3.985 ;
        RECT 32.545 3.505 32.685 3.755 ;
        RECT 32.855 3.745 33.175 4.005 ;
        RECT 33.905 3.805 34.045 4.445 ;
        RECT 35.755 4.505 36.045 4.545 ;
        RECT 45.495 4.505 45.785 4.545 ;
        RECT 35.755 4.365 36.325 4.505 ;
        RECT 34.385 4.285 35.485 4.365 ;
        RECT 35.755 4.315 36.045 4.365 ;
        RECT 34.195 4.265 35.485 4.285 ;
        RECT 36.185 4.265 36.445 4.365 ;
        RECT 34.195 4.225 35.565 4.265 ;
        RECT 36.185 4.225 36.525 4.265 ;
        RECT 34.195 4.035 34.605 4.225 ;
        RECT 35.275 4.035 35.565 4.225 ;
        RECT 36.235 4.035 36.525 4.225 ;
        RECT 34.195 4.025 34.515 4.035 ;
        RECT 34.795 3.805 35.085 3.985 ;
        RECT 33.905 3.755 35.085 3.805 ;
        RECT 33.905 3.705 35.005 3.755 ;
        RECT 35.735 3.745 36.055 4.005 ;
        RECT 37.720 3.995 38.060 4.345 ;
        RECT 45.495 4.315 45.945 4.505 ;
        RECT 44.755 4.025 45.075 4.285 ;
        RECT 33.835 3.665 35.005 3.705 ;
        RECT 32.545 3.445 32.845 3.505 ;
        RECT 33.835 3.455 34.125 3.665 ;
        RECT 37.810 3.490 37.980 3.995 ;
        RECT 39.325 3.875 39.645 3.980 ;
        RECT 39.300 3.860 39.645 3.875 ;
        RECT 39.290 3.845 39.645 3.860 ;
        RECT 39.125 3.675 39.645 3.845 ;
        RECT 39.300 3.660 39.645 3.675 ;
        RECT 39.300 3.645 39.590 3.660 ;
        RECT 40.100 3.490 40.450 3.610 ;
        RECT 41.460 3.540 41.750 3.775 ;
        RECT 45.235 3.745 45.555 4.005 ;
        RECT 45.805 3.985 45.945 4.315 ;
        RECT 46.435 4.315 46.985 4.545 ;
        RECT 47.125 4.445 49.305 4.585 ;
        RECT 61.695 4.545 62.015 4.565 ;
        RECT 47.125 4.365 48.425 4.445 ;
        RECT 46.435 4.305 46.755 4.315 ;
        RECT 47.125 4.085 47.465 4.365 ;
        RECT 48.135 4.315 48.425 4.365 ;
        RECT 47.175 4.035 47.465 4.085 ;
        RECT 48.595 4.025 48.915 4.285 ;
        RECT 45.805 3.845 46.065 3.985 ;
        RECT 41.460 3.535 41.690 3.540 ;
        RECT 30.665 3.385 31.005 3.425 ;
        RECT 31.535 3.385 31.855 3.445 ;
        RECT 30.665 3.245 31.855 3.385 ;
        RECT 30.715 3.195 31.005 3.245 ;
        RECT 31.535 3.185 31.855 3.245 ;
        RECT 32.005 3.185 32.405 3.445 ;
        RECT 32.545 3.385 32.935 3.445 ;
        RECT 33.335 3.425 33.655 3.445 ;
        RECT 33.115 3.385 33.655 3.425 ;
        RECT 32.545 3.365 33.655 3.385 ;
        RECT 32.615 3.245 33.655 3.365 ;
        RECT 32.615 3.185 32.935 3.245 ;
        RECT 33.115 3.195 33.655 3.245 ;
        RECT 33.335 3.185 33.655 3.195 ;
        RECT 34.565 3.385 34.885 3.445 ;
        RECT 35.035 3.385 35.325 3.425 ;
        RECT 34.565 3.245 35.325 3.385 ;
        RECT 34.565 3.185 34.885 3.245 ;
        RECT 35.035 3.195 35.325 3.245 ;
        RECT 35.995 3.385 36.285 3.425 ;
        RECT 36.425 3.385 36.745 3.445 ;
        RECT 35.995 3.245 36.745 3.385 ;
        RECT 37.810 3.320 40.450 3.490 ;
        RECT 39.930 3.315 40.450 3.320 ;
        RECT 40.100 3.260 40.450 3.315 ;
        RECT 35.995 3.195 36.285 3.245 ;
        RECT 36.425 3.185 36.745 3.245 ;
        RECT 41.090 3.205 41.320 3.230 ;
        RECT 39.670 3.120 39.960 3.145 ;
        RECT 41.060 3.120 41.350 3.205 ;
        RECT 39.670 2.950 41.350 3.120 ;
        RECT 39.670 2.915 39.960 2.950 ;
        RECT 39.730 2.405 39.900 2.915 ;
        RECT 41.060 2.900 41.350 2.950 ;
        RECT 41.090 2.880 41.320 2.900 ;
        RECT 41.520 2.435 41.690 3.535 ;
        RECT 44.065 3.185 44.385 3.445 ;
        RECT 45.925 3.425 46.065 3.845 ;
        RECT 46.215 3.945 46.505 3.985 ;
        RECT 46.675 3.945 46.995 4.005 ;
        RECT 46.215 3.805 46.995 3.945 ;
        RECT 46.215 3.755 46.505 3.805 ;
        RECT 46.675 3.745 46.995 3.805 ;
        RECT 47.655 3.755 47.945 3.985 ;
        RECT 47.805 3.505 47.945 3.755 ;
        RECT 48.115 3.745 48.435 4.005 ;
        RECT 49.165 3.805 49.305 4.445 ;
        RECT 51.015 4.505 51.305 4.545 ;
        RECT 60.755 4.505 61.045 4.545 ;
        RECT 51.015 4.365 51.585 4.505 ;
        RECT 49.645 4.285 50.745 4.365 ;
        RECT 51.015 4.315 51.305 4.365 ;
        RECT 49.455 4.265 50.745 4.285 ;
        RECT 51.445 4.265 51.705 4.365 ;
        RECT 49.455 4.225 50.825 4.265 ;
        RECT 51.445 4.225 51.785 4.265 ;
        RECT 49.455 4.035 49.865 4.225 ;
        RECT 50.535 4.035 50.825 4.225 ;
        RECT 51.495 4.035 51.785 4.225 ;
        RECT 49.455 4.025 49.775 4.035 ;
        RECT 50.055 3.805 50.345 3.985 ;
        RECT 49.165 3.755 50.345 3.805 ;
        RECT 49.165 3.705 50.265 3.755 ;
        RECT 50.995 3.745 51.315 4.005 ;
        RECT 52.980 3.995 53.320 4.345 ;
        RECT 60.755 4.315 61.205 4.505 ;
        RECT 60.015 4.025 60.335 4.285 ;
        RECT 49.095 3.665 50.265 3.705 ;
        RECT 47.805 3.445 48.105 3.505 ;
        RECT 49.095 3.455 49.385 3.665 ;
        RECT 53.070 3.490 53.240 3.995 ;
        RECT 54.585 3.875 54.905 3.980 ;
        RECT 54.560 3.860 54.905 3.875 ;
        RECT 54.550 3.845 54.905 3.860 ;
        RECT 54.385 3.675 54.905 3.845 ;
        RECT 54.560 3.660 54.905 3.675 ;
        RECT 54.560 3.645 54.850 3.660 ;
        RECT 55.360 3.490 55.710 3.610 ;
        RECT 56.720 3.540 57.010 3.775 ;
        RECT 60.495 3.745 60.815 4.005 ;
        RECT 61.065 3.985 61.205 4.315 ;
        RECT 61.695 4.315 62.245 4.545 ;
        RECT 62.385 4.445 64.565 4.585 ;
        RECT 76.955 4.545 77.275 4.565 ;
        RECT 62.385 4.365 63.685 4.445 ;
        RECT 61.695 4.305 62.015 4.315 ;
        RECT 62.385 4.085 62.725 4.365 ;
        RECT 63.395 4.315 63.685 4.365 ;
        RECT 62.435 4.035 62.725 4.085 ;
        RECT 63.855 4.025 64.175 4.285 ;
        RECT 61.065 3.845 61.325 3.985 ;
        RECT 56.720 3.535 56.950 3.540 ;
        RECT 45.925 3.385 46.265 3.425 ;
        RECT 46.795 3.385 47.115 3.445 ;
        RECT 45.925 3.245 47.115 3.385 ;
        RECT 45.975 3.195 46.265 3.245 ;
        RECT 46.795 3.185 47.115 3.245 ;
        RECT 47.265 3.185 47.665 3.445 ;
        RECT 47.805 3.385 48.195 3.445 ;
        RECT 48.595 3.425 48.915 3.445 ;
        RECT 48.375 3.385 48.915 3.425 ;
        RECT 47.805 3.365 48.915 3.385 ;
        RECT 47.875 3.245 48.915 3.365 ;
        RECT 47.875 3.185 48.195 3.245 ;
        RECT 48.375 3.195 48.915 3.245 ;
        RECT 48.595 3.185 48.915 3.195 ;
        RECT 49.825 3.385 50.145 3.445 ;
        RECT 50.295 3.385 50.585 3.425 ;
        RECT 49.825 3.245 50.585 3.385 ;
        RECT 49.825 3.185 50.145 3.245 ;
        RECT 50.295 3.195 50.585 3.245 ;
        RECT 51.255 3.385 51.545 3.425 ;
        RECT 51.685 3.385 52.005 3.445 ;
        RECT 51.255 3.245 52.005 3.385 ;
        RECT 53.070 3.320 55.710 3.490 ;
        RECT 55.190 3.315 55.710 3.320 ;
        RECT 55.360 3.260 55.710 3.315 ;
        RECT 51.255 3.195 51.545 3.245 ;
        RECT 51.685 3.185 52.005 3.245 ;
        RECT 56.350 3.205 56.580 3.230 ;
        RECT 54.930 3.120 55.220 3.145 ;
        RECT 56.320 3.120 56.610 3.205 ;
        RECT 54.930 2.950 56.610 3.120 ;
        RECT 54.930 2.915 55.220 2.950 ;
        RECT 39.670 2.175 39.960 2.405 ;
        RECT 41.460 2.175 41.755 2.435 ;
        RECT 54.990 2.405 55.160 2.915 ;
        RECT 56.320 2.900 56.610 2.950 ;
        RECT 56.350 2.880 56.580 2.900 ;
        RECT 56.780 2.435 56.950 3.535 ;
        RECT 59.325 3.185 59.645 3.445 ;
        RECT 61.185 3.425 61.325 3.845 ;
        RECT 61.475 3.945 61.765 3.985 ;
        RECT 61.935 3.945 62.255 4.005 ;
        RECT 61.475 3.805 62.255 3.945 ;
        RECT 61.475 3.755 61.765 3.805 ;
        RECT 61.935 3.745 62.255 3.805 ;
        RECT 62.915 3.755 63.205 3.985 ;
        RECT 63.065 3.505 63.205 3.755 ;
        RECT 63.375 3.745 63.695 4.005 ;
        RECT 64.425 3.805 64.565 4.445 ;
        RECT 66.275 4.505 66.565 4.545 ;
        RECT 76.015 4.505 76.305 4.545 ;
        RECT 66.275 4.365 66.845 4.505 ;
        RECT 64.905 4.285 66.005 4.365 ;
        RECT 66.275 4.315 66.565 4.365 ;
        RECT 64.715 4.265 66.005 4.285 ;
        RECT 66.705 4.265 66.965 4.365 ;
        RECT 64.715 4.225 66.085 4.265 ;
        RECT 66.705 4.225 67.045 4.265 ;
        RECT 64.715 4.035 65.125 4.225 ;
        RECT 65.795 4.035 66.085 4.225 ;
        RECT 66.755 4.035 67.045 4.225 ;
        RECT 64.715 4.025 65.035 4.035 ;
        RECT 65.315 3.805 65.605 3.985 ;
        RECT 64.425 3.755 65.605 3.805 ;
        RECT 64.425 3.705 65.525 3.755 ;
        RECT 66.255 3.745 66.575 4.005 ;
        RECT 68.240 3.995 68.580 4.345 ;
        RECT 76.015 4.315 76.465 4.505 ;
        RECT 75.275 4.025 75.595 4.285 ;
        RECT 64.355 3.665 65.525 3.705 ;
        RECT 63.065 3.445 63.365 3.505 ;
        RECT 64.355 3.455 64.645 3.665 ;
        RECT 68.330 3.490 68.500 3.995 ;
        RECT 69.845 3.875 70.165 3.980 ;
        RECT 69.820 3.860 70.165 3.875 ;
        RECT 69.810 3.845 70.165 3.860 ;
        RECT 69.645 3.675 70.165 3.845 ;
        RECT 69.820 3.660 70.165 3.675 ;
        RECT 69.820 3.645 70.110 3.660 ;
        RECT 70.620 3.490 70.970 3.610 ;
        RECT 71.980 3.540 72.270 3.775 ;
        RECT 75.755 3.745 76.075 4.005 ;
        RECT 76.325 3.985 76.465 4.315 ;
        RECT 76.955 4.315 77.505 4.545 ;
        RECT 77.645 4.445 79.825 4.585 ;
        RECT 92.215 4.545 92.535 4.565 ;
        RECT 77.645 4.365 78.945 4.445 ;
        RECT 76.955 4.305 77.275 4.315 ;
        RECT 77.645 4.085 77.985 4.365 ;
        RECT 78.655 4.315 78.945 4.365 ;
        RECT 77.695 4.035 77.985 4.085 ;
        RECT 79.115 4.025 79.435 4.285 ;
        RECT 76.325 3.845 76.585 3.985 ;
        RECT 71.980 3.535 72.210 3.540 ;
        RECT 61.185 3.385 61.525 3.425 ;
        RECT 62.055 3.385 62.375 3.445 ;
        RECT 61.185 3.245 62.375 3.385 ;
        RECT 61.235 3.195 61.525 3.245 ;
        RECT 62.055 3.185 62.375 3.245 ;
        RECT 62.525 3.185 62.925 3.445 ;
        RECT 63.065 3.385 63.455 3.445 ;
        RECT 63.855 3.425 64.175 3.445 ;
        RECT 63.635 3.385 64.175 3.425 ;
        RECT 63.065 3.365 64.175 3.385 ;
        RECT 63.135 3.245 64.175 3.365 ;
        RECT 63.135 3.185 63.455 3.245 ;
        RECT 63.635 3.195 64.175 3.245 ;
        RECT 63.855 3.185 64.175 3.195 ;
        RECT 65.085 3.385 65.405 3.445 ;
        RECT 65.555 3.385 65.845 3.425 ;
        RECT 65.085 3.245 65.845 3.385 ;
        RECT 65.085 3.185 65.405 3.245 ;
        RECT 65.555 3.195 65.845 3.245 ;
        RECT 66.515 3.385 66.805 3.425 ;
        RECT 66.945 3.385 67.265 3.445 ;
        RECT 66.515 3.245 67.265 3.385 ;
        RECT 68.330 3.320 70.970 3.490 ;
        RECT 70.450 3.315 70.970 3.320 ;
        RECT 70.620 3.260 70.970 3.315 ;
        RECT 66.515 3.195 66.805 3.245 ;
        RECT 66.945 3.185 67.265 3.245 ;
        RECT 71.610 3.205 71.840 3.230 ;
        RECT 70.190 3.120 70.480 3.145 ;
        RECT 71.580 3.120 71.870 3.205 ;
        RECT 70.190 2.950 71.870 3.120 ;
        RECT 70.190 2.915 70.480 2.950 ;
        RECT 54.930 2.175 55.220 2.405 ;
        RECT 56.720 2.175 57.015 2.435 ;
        RECT 70.250 2.405 70.420 2.915 ;
        RECT 71.580 2.900 71.870 2.950 ;
        RECT 71.610 2.880 71.840 2.900 ;
        RECT 72.040 2.435 72.210 3.535 ;
        RECT 74.585 3.185 74.905 3.445 ;
        RECT 76.445 3.425 76.585 3.845 ;
        RECT 76.735 3.945 77.025 3.985 ;
        RECT 77.195 3.945 77.515 4.005 ;
        RECT 76.735 3.805 77.515 3.945 ;
        RECT 76.735 3.755 77.025 3.805 ;
        RECT 77.195 3.745 77.515 3.805 ;
        RECT 78.175 3.755 78.465 3.985 ;
        RECT 78.325 3.505 78.465 3.755 ;
        RECT 78.635 3.745 78.955 4.005 ;
        RECT 79.685 3.805 79.825 4.445 ;
        RECT 81.535 4.505 81.825 4.545 ;
        RECT 91.275 4.505 91.565 4.545 ;
        RECT 81.535 4.365 82.105 4.505 ;
        RECT 80.165 4.285 81.265 4.365 ;
        RECT 81.535 4.315 81.825 4.365 ;
        RECT 79.975 4.265 81.265 4.285 ;
        RECT 81.965 4.265 82.225 4.365 ;
        RECT 79.975 4.225 81.345 4.265 ;
        RECT 81.965 4.225 82.305 4.265 ;
        RECT 79.975 4.035 80.385 4.225 ;
        RECT 81.055 4.035 81.345 4.225 ;
        RECT 82.015 4.035 82.305 4.225 ;
        RECT 79.975 4.025 80.295 4.035 ;
        RECT 80.575 3.805 80.865 3.985 ;
        RECT 79.685 3.755 80.865 3.805 ;
        RECT 79.685 3.705 80.785 3.755 ;
        RECT 81.515 3.745 81.835 4.005 ;
        RECT 83.500 3.995 83.840 4.345 ;
        RECT 91.275 4.315 91.725 4.505 ;
        RECT 90.535 4.025 90.855 4.285 ;
        RECT 79.615 3.665 80.785 3.705 ;
        RECT 78.325 3.445 78.625 3.505 ;
        RECT 79.615 3.455 79.905 3.665 ;
        RECT 83.590 3.490 83.760 3.995 ;
        RECT 85.105 3.875 85.425 3.980 ;
        RECT 85.080 3.860 85.425 3.875 ;
        RECT 85.070 3.845 85.425 3.860 ;
        RECT 84.905 3.675 85.425 3.845 ;
        RECT 85.080 3.660 85.425 3.675 ;
        RECT 85.080 3.645 85.370 3.660 ;
        RECT 85.880 3.490 86.230 3.610 ;
        RECT 87.240 3.540 87.530 3.775 ;
        RECT 91.015 3.745 91.335 4.005 ;
        RECT 91.585 3.985 91.725 4.315 ;
        RECT 92.215 4.315 92.765 4.545 ;
        RECT 92.905 4.445 95.085 4.585 ;
        RECT 92.905 4.365 94.205 4.445 ;
        RECT 92.215 4.305 92.535 4.315 ;
        RECT 92.905 4.085 93.245 4.365 ;
        RECT 93.915 4.315 94.205 4.365 ;
        RECT 92.955 4.035 93.245 4.085 ;
        RECT 94.375 4.025 94.695 4.285 ;
        RECT 91.585 3.845 91.845 3.985 ;
        RECT 87.240 3.535 87.470 3.540 ;
        RECT 76.445 3.385 76.785 3.425 ;
        RECT 77.315 3.385 77.635 3.445 ;
        RECT 76.445 3.245 77.635 3.385 ;
        RECT 76.495 3.195 76.785 3.245 ;
        RECT 77.315 3.185 77.635 3.245 ;
        RECT 77.785 3.185 78.185 3.445 ;
        RECT 78.325 3.385 78.715 3.445 ;
        RECT 79.115 3.425 79.435 3.445 ;
        RECT 78.895 3.385 79.435 3.425 ;
        RECT 78.325 3.365 79.435 3.385 ;
        RECT 78.395 3.245 79.435 3.365 ;
        RECT 78.395 3.185 78.715 3.245 ;
        RECT 78.895 3.195 79.435 3.245 ;
        RECT 79.115 3.185 79.435 3.195 ;
        RECT 80.345 3.385 80.665 3.445 ;
        RECT 80.815 3.385 81.105 3.425 ;
        RECT 80.345 3.245 81.105 3.385 ;
        RECT 80.345 3.185 80.665 3.245 ;
        RECT 80.815 3.195 81.105 3.245 ;
        RECT 81.775 3.385 82.065 3.425 ;
        RECT 82.205 3.385 82.525 3.445 ;
        RECT 81.775 3.245 82.525 3.385 ;
        RECT 83.590 3.320 86.230 3.490 ;
        RECT 85.710 3.315 86.230 3.320 ;
        RECT 85.880 3.260 86.230 3.315 ;
        RECT 81.775 3.195 82.065 3.245 ;
        RECT 82.205 3.185 82.525 3.245 ;
        RECT 86.870 3.205 87.100 3.230 ;
        RECT 85.450 3.120 85.740 3.145 ;
        RECT 86.840 3.120 87.130 3.205 ;
        RECT 85.450 2.950 87.130 3.120 ;
        RECT 85.450 2.915 85.740 2.950 ;
        RECT 70.190 2.175 70.480 2.405 ;
        RECT 71.980 2.175 72.275 2.435 ;
        RECT 85.510 2.405 85.680 2.915 ;
        RECT 86.840 2.900 87.130 2.950 ;
        RECT 86.870 2.880 87.100 2.900 ;
        RECT 87.300 2.435 87.470 3.535 ;
        RECT 89.845 3.185 90.165 3.445 ;
        RECT 91.705 3.425 91.845 3.845 ;
        RECT 91.995 3.945 92.285 3.985 ;
        RECT 92.455 3.945 92.775 4.005 ;
        RECT 91.995 3.805 92.775 3.945 ;
        RECT 91.995 3.755 92.285 3.805 ;
        RECT 92.455 3.745 92.775 3.805 ;
        RECT 93.435 3.755 93.725 3.985 ;
        RECT 93.585 3.505 93.725 3.755 ;
        RECT 93.895 3.745 94.215 4.005 ;
        RECT 94.945 3.805 95.085 4.445 ;
        RECT 96.795 4.505 97.085 4.545 ;
        RECT 96.795 4.365 97.365 4.505 ;
        RECT 95.425 4.285 96.525 4.365 ;
        RECT 96.795 4.315 97.085 4.365 ;
        RECT 95.235 4.265 96.525 4.285 ;
        RECT 97.225 4.265 97.485 4.365 ;
        RECT 95.235 4.225 96.605 4.265 ;
        RECT 97.225 4.225 97.565 4.265 ;
        RECT 95.235 4.035 95.645 4.225 ;
        RECT 96.315 4.035 96.605 4.225 ;
        RECT 97.275 4.035 97.565 4.225 ;
        RECT 95.235 4.025 95.555 4.035 ;
        RECT 95.835 3.805 96.125 3.985 ;
        RECT 94.945 3.755 96.125 3.805 ;
        RECT 94.945 3.705 96.045 3.755 ;
        RECT 96.775 3.745 97.095 4.005 ;
        RECT 98.760 3.995 99.100 4.345 ;
        RECT 94.875 3.665 96.045 3.705 ;
        RECT 93.585 3.445 93.885 3.505 ;
        RECT 94.875 3.455 95.165 3.665 ;
        RECT 98.850 3.490 99.020 3.995 ;
        RECT 100.365 3.875 100.685 3.980 ;
        RECT 100.340 3.860 100.685 3.875 ;
        RECT 100.330 3.845 100.685 3.860 ;
        RECT 100.165 3.675 100.685 3.845 ;
        RECT 100.340 3.660 100.685 3.675 ;
        RECT 100.340 3.645 100.630 3.660 ;
        RECT 101.140 3.490 101.490 3.610 ;
        RECT 102.500 3.540 102.790 3.775 ;
        RECT 102.500 3.535 102.730 3.540 ;
        RECT 91.705 3.385 92.045 3.425 ;
        RECT 92.575 3.385 92.895 3.445 ;
        RECT 91.705 3.245 92.895 3.385 ;
        RECT 91.755 3.195 92.045 3.245 ;
        RECT 92.575 3.185 92.895 3.245 ;
        RECT 93.045 3.185 93.445 3.445 ;
        RECT 93.585 3.385 93.975 3.445 ;
        RECT 94.375 3.425 94.695 3.445 ;
        RECT 94.155 3.385 94.695 3.425 ;
        RECT 93.585 3.365 94.695 3.385 ;
        RECT 93.655 3.245 94.695 3.365 ;
        RECT 93.655 3.185 93.975 3.245 ;
        RECT 94.155 3.195 94.695 3.245 ;
        RECT 94.375 3.185 94.695 3.195 ;
        RECT 95.605 3.385 95.925 3.445 ;
        RECT 96.075 3.385 96.365 3.425 ;
        RECT 95.605 3.245 96.365 3.385 ;
        RECT 95.605 3.185 95.925 3.245 ;
        RECT 96.075 3.195 96.365 3.245 ;
        RECT 97.035 3.385 97.325 3.425 ;
        RECT 97.465 3.385 97.785 3.445 ;
        RECT 97.035 3.245 97.785 3.385 ;
        RECT 98.850 3.320 101.490 3.490 ;
        RECT 100.970 3.315 101.490 3.320 ;
        RECT 101.140 3.260 101.490 3.315 ;
        RECT 97.035 3.195 97.325 3.245 ;
        RECT 97.465 3.185 97.785 3.245 ;
        RECT 102.130 3.205 102.360 3.230 ;
        RECT 100.710 3.120 101.000 3.145 ;
        RECT 102.100 3.120 102.390 3.205 ;
        RECT 100.710 2.950 102.390 3.120 ;
        RECT 100.710 2.915 101.000 2.950 ;
        RECT 85.450 2.175 85.740 2.405 ;
        RECT 87.240 2.175 87.535 2.435 ;
        RECT 100.770 2.405 100.940 2.915 ;
        RECT 102.100 2.900 102.390 2.950 ;
        RECT 102.130 2.880 102.360 2.900 ;
        RECT 102.560 2.435 102.730 3.535 ;
        RECT 100.710 2.175 101.000 2.405 ;
        RECT 102.500 2.175 102.795 2.435 ;
      LAYER met2 ;
        RECT 26.230 10.690 103.725 10.860 ;
        RECT 26.230 8.895 26.400 10.690 ;
        RECT 103.555 9.915 103.725 10.690 ;
        RECT 26.540 9.515 26.830 9.640 ;
        RECT 26.540 9.510 26.860 9.515 ;
        RECT 26.540 9.340 27.795 9.510 ;
        RECT 34.015 9.345 34.385 9.715 ;
        RECT 49.275 9.345 49.645 9.715 ;
        RECT 64.535 9.345 64.905 9.715 ;
        RECT 79.795 9.345 80.165 9.715 ;
        RECT 95.055 9.345 95.425 9.715 ;
        RECT 103.525 9.565 103.875 9.915 ;
        RECT 26.540 9.290 26.830 9.340 ;
        RECT 27.625 9.145 27.795 9.340 ;
        RECT 34.685 9.145 35.035 9.245 ;
        RECT 40.125 9.205 40.450 9.270 ;
        RECT 27.625 8.975 35.035 9.145 ;
        RECT 34.685 8.895 35.035 8.975 ;
        RECT 39.010 9.035 40.450 9.205 ;
        RECT 26.165 8.545 26.455 8.895 ;
        RECT 31.985 5.305 34.425 5.445 ;
        RECT 31.985 5.155 32.125 5.305 ;
        RECT 31.685 5.065 32.125 5.155 ;
        RECT 29.345 4.925 32.125 5.065 ;
        RECT 28.835 4.785 29.095 4.875 ;
        RECT 29.345 4.785 29.485 4.925 ;
        RECT 31.685 4.835 31.945 4.925 ;
        RECT 32.285 4.835 32.545 5.155 ;
        RECT 32.285 4.785 32.485 4.835 ;
        RECT 28.835 4.645 29.485 4.785 ;
        RECT 32.095 4.645 32.485 4.785 ;
        RECT 33.355 4.775 33.635 5.155 ;
        RECT 33.845 4.835 34.120 5.155 ;
        RECT 28.835 4.555 29.095 4.645 ;
        RECT 28.895 3.475 29.035 4.555 ;
        RECT 29.755 4.505 30.035 4.620 ;
        RECT 31.205 4.505 31.465 4.595 ;
        RECT 29.585 4.365 31.465 4.505 ;
        RECT 29.585 4.315 30.035 4.365 ;
        RECT 29.525 4.245 30.035 4.315 ;
        RECT 31.205 4.275 31.465 4.365 ;
        RECT 29.525 4.055 29.785 4.245 ;
        RECT 30.700 4.055 31.005 4.060 ;
        RECT 29.515 3.685 29.795 4.055 ;
        RECT 30.005 3.945 30.265 4.035 ;
        RECT 30.595 3.945 31.005 4.055 ;
        RECT 30.005 3.805 31.005 3.945 ;
        RECT 30.005 3.715 30.265 3.805 ;
        RECT 30.595 3.685 31.005 3.805 ;
        RECT 31.435 3.685 31.715 4.060 ;
        RECT 32.095 3.525 32.235 4.645 ;
        RECT 33.425 4.315 33.565 4.775 ;
        RECT 32.875 3.685 33.155 4.155 ;
        RECT 33.365 4.055 33.625 4.315 ;
        RECT 33.355 3.685 33.635 4.055 ;
        RECT 32.095 3.475 32.405 3.525 ;
        RECT 33.905 3.515 34.045 4.835 ;
        RECT 34.285 4.315 34.425 5.305 ;
        RECT 34.595 4.555 34.855 4.875 ;
        RECT 36.455 4.835 36.715 5.155 ;
        RECT 34.225 3.995 34.485 4.315 ;
        RECT 34.655 3.515 34.795 4.555 ;
        RECT 36.515 4.055 36.655 4.835 ;
        RECT 37.750 4.345 38.040 4.360 ;
        RECT 35.765 3.945 36.025 4.035 ;
        RECT 35.105 3.805 36.025 3.945 ;
        RECT 33.565 3.495 34.045 3.515 ;
        RECT 28.835 3.155 29.095 3.475 ;
        RECT 31.565 3.385 31.825 3.475 ;
        RECT 32.035 3.445 32.405 3.475 ;
        RECT 31.565 3.155 31.885 3.385 ;
        RECT 31.745 3.005 31.885 3.155 ;
        RECT 32.035 3.150 32.445 3.445 ;
        RECT 32.635 3.155 32.915 3.495 ;
        RECT 33.365 3.245 34.045 3.495 ;
        RECT 34.585 3.445 34.865 3.515 ;
        RECT 33.365 3.145 33.845 3.245 ;
        RECT 34.535 3.185 34.910 3.445 ;
        RECT 34.585 3.145 34.865 3.185 ;
        RECT 35.105 3.005 35.245 3.805 ;
        RECT 35.765 3.715 36.025 3.805 ;
        RECT 36.345 3.685 36.655 4.055 ;
        RECT 37.720 3.995 38.060 4.345 ;
        RECT 37.750 3.980 38.040 3.995 ;
        RECT 39.010 3.860 39.170 9.035 ;
        RECT 40.125 8.945 40.450 9.035 ;
        RECT 42.505 9.180 42.855 9.300 ;
        RECT 49.945 9.180 50.295 9.255 ;
        RECT 55.385 9.205 55.710 9.270 ;
        RECT 42.505 8.980 50.295 9.180 ;
        RECT 42.505 8.950 42.855 8.980 ;
        RECT 49.945 8.905 50.295 8.980 ;
        RECT 54.270 9.035 55.710 9.205 ;
        RECT 39.325 8.510 39.645 8.835 ;
        RECT 39.355 8.335 39.525 8.510 ;
        RECT 39.355 8.160 39.530 8.335 ;
        RECT 39.355 7.985 40.330 8.160 ;
        RECT 39.325 3.860 39.645 3.980 ;
        RECT 39.010 3.690 39.645 3.860 ;
        RECT 36.415 3.500 36.655 3.685 ;
        RECT 39.325 3.660 39.645 3.690 ;
        RECT 40.155 3.610 40.330 7.985 ;
        RECT 47.245 5.305 49.685 5.445 ;
        RECT 47.245 5.155 47.385 5.305 ;
        RECT 46.945 5.065 47.385 5.155 ;
        RECT 44.605 4.925 47.385 5.065 ;
        RECT 44.095 4.785 44.355 4.875 ;
        RECT 44.605 4.785 44.745 4.925 ;
        RECT 46.945 4.835 47.205 4.925 ;
        RECT 47.545 4.835 47.805 5.155 ;
        RECT 47.545 4.785 47.745 4.835 ;
        RECT 44.095 4.645 44.745 4.785 ;
        RECT 47.355 4.645 47.745 4.785 ;
        RECT 48.615 4.775 48.895 5.155 ;
        RECT 49.105 4.835 49.380 5.155 ;
        RECT 44.095 4.555 44.355 4.645 ;
        RECT 36.415 3.435 36.725 3.500 ;
        RECT 36.415 3.245 36.730 3.435 ;
        RECT 40.100 3.260 40.450 3.610 ;
        RECT 44.155 3.475 44.295 4.555 ;
        RECT 45.015 4.505 45.295 4.620 ;
        RECT 46.465 4.505 46.725 4.595 ;
        RECT 44.845 4.365 46.725 4.505 ;
        RECT 44.845 4.315 45.295 4.365 ;
        RECT 44.785 4.245 45.295 4.315 ;
        RECT 46.465 4.275 46.725 4.365 ;
        RECT 44.785 4.055 45.045 4.245 ;
        RECT 45.960 4.055 46.265 4.060 ;
        RECT 44.775 3.685 45.055 4.055 ;
        RECT 45.265 3.945 45.525 4.035 ;
        RECT 45.855 3.945 46.265 4.055 ;
        RECT 45.265 3.805 46.265 3.945 ;
        RECT 45.265 3.715 45.525 3.805 ;
        RECT 45.855 3.685 46.265 3.805 ;
        RECT 46.695 3.685 46.975 4.060 ;
        RECT 47.355 3.525 47.495 4.645 ;
        RECT 48.685 4.315 48.825 4.775 ;
        RECT 48.135 3.685 48.415 4.155 ;
        RECT 48.625 4.055 48.885 4.315 ;
        RECT 48.615 3.685 48.895 4.055 ;
        RECT 47.355 3.475 47.665 3.525 ;
        RECT 49.165 3.515 49.305 4.835 ;
        RECT 49.545 4.315 49.685 5.305 ;
        RECT 49.855 4.555 50.115 4.875 ;
        RECT 51.715 4.835 51.975 5.155 ;
        RECT 49.485 3.995 49.745 4.315 ;
        RECT 49.915 3.515 50.055 4.555 ;
        RECT 51.775 4.055 51.915 4.835 ;
        RECT 53.010 4.345 53.300 4.360 ;
        RECT 51.025 3.945 51.285 4.035 ;
        RECT 50.365 3.805 51.285 3.945 ;
        RECT 48.825 3.495 49.305 3.515 ;
        RECT 36.445 3.235 36.730 3.245 ;
        RECT 36.445 3.125 36.725 3.235 ;
        RECT 44.095 3.155 44.355 3.475 ;
        RECT 46.825 3.385 47.085 3.475 ;
        RECT 47.295 3.445 47.665 3.475 ;
        RECT 46.825 3.155 47.145 3.385 ;
        RECT 31.745 2.865 35.245 3.005 ;
        RECT 47.005 3.005 47.145 3.155 ;
        RECT 47.295 3.150 47.705 3.445 ;
        RECT 47.895 3.155 48.175 3.495 ;
        RECT 48.625 3.245 49.305 3.495 ;
        RECT 49.845 3.445 50.125 3.515 ;
        RECT 48.625 3.145 49.105 3.245 ;
        RECT 49.795 3.185 50.170 3.445 ;
        RECT 49.845 3.145 50.125 3.185 ;
        RECT 50.365 3.005 50.505 3.805 ;
        RECT 51.025 3.715 51.285 3.805 ;
        RECT 51.605 3.685 51.915 4.055 ;
        RECT 52.980 3.995 53.320 4.345 ;
        RECT 53.010 3.980 53.300 3.995 ;
        RECT 54.270 3.860 54.430 9.035 ;
        RECT 55.385 8.945 55.710 9.035 ;
        RECT 57.765 9.180 58.115 9.300 ;
        RECT 65.205 9.180 65.555 9.255 ;
        RECT 70.645 9.205 70.970 9.270 ;
        RECT 57.765 8.980 65.555 9.180 ;
        RECT 57.765 8.950 58.115 8.980 ;
        RECT 65.205 8.905 65.555 8.980 ;
        RECT 69.530 9.035 70.970 9.205 ;
        RECT 54.585 8.510 54.905 8.835 ;
        RECT 54.615 8.335 54.785 8.510 ;
        RECT 54.615 8.160 54.790 8.335 ;
        RECT 54.615 7.985 55.590 8.160 ;
        RECT 54.585 3.860 54.905 3.980 ;
        RECT 54.270 3.690 54.905 3.860 ;
        RECT 51.675 3.500 51.915 3.685 ;
        RECT 54.585 3.660 54.905 3.690 ;
        RECT 55.415 3.610 55.590 7.985 ;
        RECT 62.505 5.305 64.945 5.445 ;
        RECT 62.505 5.155 62.645 5.305 ;
        RECT 62.205 5.065 62.645 5.155 ;
        RECT 59.865 4.925 62.645 5.065 ;
        RECT 59.355 4.785 59.615 4.875 ;
        RECT 59.865 4.785 60.005 4.925 ;
        RECT 62.205 4.835 62.465 4.925 ;
        RECT 62.805 4.835 63.065 5.155 ;
        RECT 62.805 4.785 63.005 4.835 ;
        RECT 59.355 4.645 60.005 4.785 ;
        RECT 62.615 4.645 63.005 4.785 ;
        RECT 63.875 4.775 64.155 5.155 ;
        RECT 64.365 4.835 64.640 5.155 ;
        RECT 59.355 4.555 59.615 4.645 ;
        RECT 51.675 3.435 51.985 3.500 ;
        RECT 51.675 3.245 51.990 3.435 ;
        RECT 55.360 3.260 55.710 3.610 ;
        RECT 59.415 3.475 59.555 4.555 ;
        RECT 60.275 4.505 60.555 4.620 ;
        RECT 61.725 4.505 61.985 4.595 ;
        RECT 60.105 4.365 61.985 4.505 ;
        RECT 60.105 4.315 60.555 4.365 ;
        RECT 60.045 4.245 60.555 4.315 ;
        RECT 61.725 4.275 61.985 4.365 ;
        RECT 60.045 4.055 60.305 4.245 ;
        RECT 61.220 4.055 61.525 4.060 ;
        RECT 60.035 3.685 60.315 4.055 ;
        RECT 60.525 3.945 60.785 4.035 ;
        RECT 61.115 3.945 61.525 4.055 ;
        RECT 60.525 3.805 61.525 3.945 ;
        RECT 60.525 3.715 60.785 3.805 ;
        RECT 61.115 3.685 61.525 3.805 ;
        RECT 61.955 3.685 62.235 4.060 ;
        RECT 62.615 3.525 62.755 4.645 ;
        RECT 63.945 4.315 64.085 4.775 ;
        RECT 63.395 3.685 63.675 4.155 ;
        RECT 63.885 4.055 64.145 4.315 ;
        RECT 63.875 3.685 64.155 4.055 ;
        RECT 62.615 3.475 62.925 3.525 ;
        RECT 64.425 3.515 64.565 4.835 ;
        RECT 64.805 4.315 64.945 5.305 ;
        RECT 65.115 4.555 65.375 4.875 ;
        RECT 66.975 4.835 67.235 5.155 ;
        RECT 64.745 3.995 65.005 4.315 ;
        RECT 65.175 3.515 65.315 4.555 ;
        RECT 67.035 4.055 67.175 4.835 ;
        RECT 68.270 4.345 68.560 4.360 ;
        RECT 66.285 3.945 66.545 4.035 ;
        RECT 65.625 3.805 66.545 3.945 ;
        RECT 64.085 3.495 64.565 3.515 ;
        RECT 51.705 3.235 51.990 3.245 ;
        RECT 51.705 3.125 51.985 3.235 ;
        RECT 59.355 3.155 59.615 3.475 ;
        RECT 62.085 3.385 62.345 3.475 ;
        RECT 62.555 3.445 62.925 3.475 ;
        RECT 62.085 3.155 62.405 3.385 ;
        RECT 47.005 2.865 50.505 3.005 ;
        RECT 62.265 3.005 62.405 3.155 ;
        RECT 62.555 3.150 62.965 3.445 ;
        RECT 63.155 3.155 63.435 3.495 ;
        RECT 63.885 3.245 64.565 3.495 ;
        RECT 65.105 3.445 65.385 3.515 ;
        RECT 63.885 3.145 64.365 3.245 ;
        RECT 65.055 3.185 65.430 3.445 ;
        RECT 65.105 3.145 65.385 3.185 ;
        RECT 65.625 3.005 65.765 3.805 ;
        RECT 66.285 3.715 66.545 3.805 ;
        RECT 66.865 3.685 67.175 4.055 ;
        RECT 68.240 3.995 68.580 4.345 ;
        RECT 68.270 3.980 68.560 3.995 ;
        RECT 69.530 3.860 69.690 9.035 ;
        RECT 70.645 8.945 70.970 9.035 ;
        RECT 72.980 9.180 73.330 9.300 ;
        RECT 80.470 9.180 80.820 9.255 ;
        RECT 85.905 9.205 86.230 9.270 ;
        RECT 72.980 8.980 80.820 9.180 ;
        RECT 72.980 8.950 73.330 8.980 ;
        RECT 80.470 8.905 80.820 8.980 ;
        RECT 84.790 9.035 86.230 9.205 ;
        RECT 69.845 8.510 70.165 8.835 ;
        RECT 69.875 8.335 70.045 8.510 ;
        RECT 69.875 8.160 70.050 8.335 ;
        RECT 69.875 7.985 70.850 8.160 ;
        RECT 69.845 3.860 70.165 3.980 ;
        RECT 69.530 3.690 70.165 3.860 ;
        RECT 66.935 3.500 67.175 3.685 ;
        RECT 69.845 3.660 70.165 3.690 ;
        RECT 70.675 3.610 70.850 7.985 ;
        RECT 77.765 5.305 80.205 5.445 ;
        RECT 77.765 5.155 77.905 5.305 ;
        RECT 77.465 5.065 77.905 5.155 ;
        RECT 75.125 4.925 77.905 5.065 ;
        RECT 74.615 4.785 74.875 4.875 ;
        RECT 75.125 4.785 75.265 4.925 ;
        RECT 77.465 4.835 77.725 4.925 ;
        RECT 78.065 4.835 78.325 5.155 ;
        RECT 78.065 4.785 78.265 4.835 ;
        RECT 74.615 4.645 75.265 4.785 ;
        RECT 77.875 4.645 78.265 4.785 ;
        RECT 79.135 4.775 79.415 5.155 ;
        RECT 79.625 4.835 79.900 5.155 ;
        RECT 74.615 4.555 74.875 4.645 ;
        RECT 66.935 3.435 67.245 3.500 ;
        RECT 66.935 3.245 67.250 3.435 ;
        RECT 70.620 3.260 70.970 3.610 ;
        RECT 74.675 3.475 74.815 4.555 ;
        RECT 75.535 4.505 75.815 4.620 ;
        RECT 76.985 4.505 77.245 4.595 ;
        RECT 75.365 4.365 77.245 4.505 ;
        RECT 75.365 4.315 75.815 4.365 ;
        RECT 75.305 4.245 75.815 4.315 ;
        RECT 76.985 4.275 77.245 4.365 ;
        RECT 75.305 4.055 75.565 4.245 ;
        RECT 76.480 4.055 76.785 4.060 ;
        RECT 75.295 3.685 75.575 4.055 ;
        RECT 75.785 3.945 76.045 4.035 ;
        RECT 76.375 3.945 76.785 4.055 ;
        RECT 75.785 3.805 76.785 3.945 ;
        RECT 75.785 3.715 76.045 3.805 ;
        RECT 76.375 3.685 76.785 3.805 ;
        RECT 77.215 3.685 77.495 4.060 ;
        RECT 77.875 3.525 78.015 4.645 ;
        RECT 79.205 4.315 79.345 4.775 ;
        RECT 78.655 3.685 78.935 4.155 ;
        RECT 79.145 4.055 79.405 4.315 ;
        RECT 79.135 3.685 79.415 4.055 ;
        RECT 77.875 3.475 78.185 3.525 ;
        RECT 79.685 3.515 79.825 4.835 ;
        RECT 80.065 4.315 80.205 5.305 ;
        RECT 80.375 4.555 80.635 4.875 ;
        RECT 82.235 4.835 82.495 5.155 ;
        RECT 80.005 3.995 80.265 4.315 ;
        RECT 80.435 3.515 80.575 4.555 ;
        RECT 82.295 4.055 82.435 4.835 ;
        RECT 83.530 4.345 83.820 4.360 ;
        RECT 81.545 3.945 81.805 4.035 ;
        RECT 80.885 3.805 81.805 3.945 ;
        RECT 79.345 3.495 79.825 3.515 ;
        RECT 66.965 3.235 67.250 3.245 ;
        RECT 66.965 3.125 67.245 3.235 ;
        RECT 74.615 3.155 74.875 3.475 ;
        RECT 77.345 3.385 77.605 3.475 ;
        RECT 77.815 3.445 78.185 3.475 ;
        RECT 77.345 3.155 77.665 3.385 ;
        RECT 62.265 2.865 65.765 3.005 ;
        RECT 77.525 3.005 77.665 3.155 ;
        RECT 77.815 3.150 78.225 3.445 ;
        RECT 78.415 3.155 78.695 3.495 ;
        RECT 79.145 3.245 79.825 3.495 ;
        RECT 80.365 3.445 80.645 3.515 ;
        RECT 79.145 3.145 79.625 3.245 ;
        RECT 80.315 3.185 80.690 3.445 ;
        RECT 80.365 3.145 80.645 3.185 ;
        RECT 80.885 3.005 81.025 3.805 ;
        RECT 81.545 3.715 81.805 3.805 ;
        RECT 82.125 3.685 82.435 4.055 ;
        RECT 83.500 3.995 83.840 4.345 ;
        RECT 83.530 3.980 83.820 3.995 ;
        RECT 84.790 3.860 84.950 9.035 ;
        RECT 85.905 8.945 86.230 9.035 ;
        RECT 88.240 9.180 88.590 9.300 ;
        RECT 95.725 9.180 96.075 9.255 ;
        RECT 101.165 9.205 101.490 9.270 ;
        RECT 88.240 8.980 96.075 9.180 ;
        RECT 88.240 8.950 88.590 8.980 ;
        RECT 95.725 8.905 96.075 8.980 ;
        RECT 100.050 9.035 101.490 9.205 ;
        RECT 85.105 8.510 85.425 8.835 ;
        RECT 85.135 8.335 85.305 8.510 ;
        RECT 85.135 8.160 85.310 8.335 ;
        RECT 85.135 7.985 86.110 8.160 ;
        RECT 85.105 3.860 85.425 3.980 ;
        RECT 84.790 3.690 85.425 3.860 ;
        RECT 82.195 3.500 82.435 3.685 ;
        RECT 85.105 3.660 85.425 3.690 ;
        RECT 85.935 3.610 86.110 7.985 ;
        RECT 93.025 5.305 95.465 5.445 ;
        RECT 93.025 5.155 93.165 5.305 ;
        RECT 92.725 5.065 93.165 5.155 ;
        RECT 90.385 4.925 93.165 5.065 ;
        RECT 89.875 4.785 90.135 4.875 ;
        RECT 90.385 4.785 90.525 4.925 ;
        RECT 92.725 4.835 92.985 4.925 ;
        RECT 93.325 4.835 93.585 5.155 ;
        RECT 93.325 4.785 93.525 4.835 ;
        RECT 89.875 4.645 90.525 4.785 ;
        RECT 93.135 4.645 93.525 4.785 ;
        RECT 94.395 4.775 94.675 5.155 ;
        RECT 94.885 4.835 95.160 5.155 ;
        RECT 89.875 4.555 90.135 4.645 ;
        RECT 82.195 3.435 82.505 3.500 ;
        RECT 82.195 3.245 82.510 3.435 ;
        RECT 85.880 3.260 86.230 3.610 ;
        RECT 89.935 3.475 90.075 4.555 ;
        RECT 90.795 4.505 91.075 4.620 ;
        RECT 92.245 4.505 92.505 4.595 ;
        RECT 90.625 4.365 92.505 4.505 ;
        RECT 90.625 4.315 91.075 4.365 ;
        RECT 90.565 4.245 91.075 4.315 ;
        RECT 92.245 4.275 92.505 4.365 ;
        RECT 90.565 4.055 90.825 4.245 ;
        RECT 91.740 4.055 92.045 4.060 ;
        RECT 90.555 3.685 90.835 4.055 ;
        RECT 91.045 3.945 91.305 4.035 ;
        RECT 91.635 3.945 92.045 4.055 ;
        RECT 91.045 3.805 92.045 3.945 ;
        RECT 91.045 3.715 91.305 3.805 ;
        RECT 91.635 3.685 92.045 3.805 ;
        RECT 92.475 3.685 92.755 4.060 ;
        RECT 93.135 3.525 93.275 4.645 ;
        RECT 94.465 4.315 94.605 4.775 ;
        RECT 93.915 3.685 94.195 4.155 ;
        RECT 94.405 4.055 94.665 4.315 ;
        RECT 94.395 3.685 94.675 4.055 ;
        RECT 93.135 3.475 93.445 3.525 ;
        RECT 94.945 3.515 95.085 4.835 ;
        RECT 95.325 4.315 95.465 5.305 ;
        RECT 95.635 4.555 95.895 4.875 ;
        RECT 97.495 4.835 97.755 5.155 ;
        RECT 95.265 3.995 95.525 4.315 ;
        RECT 95.695 3.515 95.835 4.555 ;
        RECT 97.555 4.055 97.695 4.835 ;
        RECT 98.790 4.345 99.080 4.360 ;
        RECT 96.805 3.945 97.065 4.035 ;
        RECT 96.145 3.805 97.065 3.945 ;
        RECT 94.605 3.495 95.085 3.515 ;
        RECT 82.225 3.235 82.510 3.245 ;
        RECT 82.225 3.125 82.505 3.235 ;
        RECT 89.875 3.155 90.135 3.475 ;
        RECT 92.605 3.385 92.865 3.475 ;
        RECT 93.075 3.445 93.445 3.475 ;
        RECT 92.605 3.155 92.925 3.385 ;
        RECT 77.525 2.865 81.025 3.005 ;
        RECT 92.785 3.005 92.925 3.155 ;
        RECT 93.075 3.150 93.485 3.445 ;
        RECT 93.675 3.155 93.955 3.495 ;
        RECT 94.405 3.245 95.085 3.495 ;
        RECT 95.625 3.445 95.905 3.515 ;
        RECT 94.405 3.145 94.885 3.245 ;
        RECT 95.575 3.185 95.950 3.445 ;
        RECT 95.625 3.145 95.905 3.185 ;
        RECT 96.145 3.005 96.285 3.805 ;
        RECT 96.805 3.715 97.065 3.805 ;
        RECT 97.385 3.685 97.695 4.055 ;
        RECT 98.760 3.995 99.100 4.345 ;
        RECT 98.790 3.980 99.080 3.995 ;
        RECT 100.050 3.860 100.210 9.035 ;
        RECT 101.165 8.945 101.490 9.035 ;
        RECT 100.365 8.510 100.685 8.835 ;
        RECT 100.395 8.335 100.565 8.510 ;
        RECT 100.395 8.160 100.570 8.335 ;
        RECT 100.395 7.985 101.370 8.160 ;
        RECT 100.365 3.860 100.685 3.980 ;
        RECT 100.050 3.690 100.685 3.860 ;
        RECT 97.455 3.500 97.695 3.685 ;
        RECT 100.365 3.660 100.685 3.690 ;
        RECT 101.195 3.610 101.370 7.985 ;
        RECT 97.455 3.435 97.765 3.500 ;
        RECT 97.455 3.245 97.770 3.435 ;
        RECT 101.140 3.260 101.490 3.610 ;
        RECT 97.485 3.235 97.770 3.245 ;
        RECT 97.485 3.125 97.765 3.235 ;
        RECT 92.785 2.865 96.285 3.005 ;
      LAYER met3 ;
        RECT 34.015 9.345 34.385 9.715 ;
        RECT 49.275 9.345 49.645 9.715 ;
        RECT 64.535 9.345 64.905 9.715 ;
        RECT 79.795 9.345 80.165 9.715 ;
        RECT 95.055 9.345 95.425 9.715 ;
        RECT 34.050 6.070 34.350 9.345 ;
        RECT 49.310 6.070 49.610 9.345 ;
        RECT 64.570 6.070 64.870 9.345 ;
        RECT 79.830 6.070 80.130 9.345 ;
        RECT 95.090 6.070 95.390 9.345 ;
        RECT 29.815 5.770 34.350 6.070 ;
        RECT 45.075 5.770 49.610 6.070 ;
        RECT 60.335 5.770 64.870 6.070 ;
        RECT 75.595 5.770 80.130 6.070 ;
        RECT 90.855 5.770 95.390 6.070 ;
        RECT 29.815 5.550 32.910 5.770 ;
        RECT 29.815 4.600 30.115 5.550 ;
        RECT 32.610 5.145 32.910 5.550 ;
        RECT 45.075 5.550 48.170 5.770 ;
        RECT 33.335 5.145 33.665 5.155 ;
        RECT 31.425 4.845 33.665 5.145 ;
        RECT 29.735 4.595 30.115 4.600 ;
        RECT 29.505 4.265 30.235 4.595 ;
        RECT 30.695 4.245 31.015 4.625 ;
        RECT 30.695 4.055 31.025 4.245 ;
        RECT 31.425 4.055 31.725 4.845 ;
        RECT 32.610 4.155 32.910 4.845 ;
        RECT 33.325 4.795 33.665 4.845 ;
        RECT 45.075 4.600 45.375 5.550 ;
        RECT 47.870 5.145 48.170 5.550 ;
        RECT 60.335 5.550 63.430 5.770 ;
        RECT 48.595 5.145 48.925 5.155 ;
        RECT 46.685 4.845 48.925 5.145 ;
        RECT 44.995 4.595 45.375 4.600 ;
        RECT 30.695 3.705 31.030 4.055 ;
        RECT 31.405 4.040 31.725 4.055 ;
        RECT 31.405 3.705 31.745 4.040 ;
        RECT 32.405 3.815 33.185 4.155 ;
        RECT 32.610 3.810 33.185 3.815 ;
        RECT 32.845 3.805 33.185 3.810 ;
        RECT 32.855 3.775 33.185 3.805 ;
        RECT 37.720 3.940 38.080 4.365 ;
        RECT 44.765 4.265 45.495 4.595 ;
        RECT 45.955 4.245 46.275 4.625 ;
        RECT 45.955 4.055 46.285 4.245 ;
        RECT 46.685 4.055 46.985 4.845 ;
        RECT 47.870 4.155 48.170 4.845 ;
        RECT 48.585 4.795 48.925 4.845 ;
        RECT 60.335 4.600 60.635 5.550 ;
        RECT 63.130 5.145 63.430 5.550 ;
        RECT 75.595 5.550 78.690 5.770 ;
        RECT 63.855 5.145 64.185 5.155 ;
        RECT 61.945 4.845 64.185 5.145 ;
        RECT 60.255 4.595 60.635 4.600 ;
        RECT 31.975 3.175 32.705 3.505 ;
        RECT 33.520 3.495 33.870 3.500 ;
        RECT 31.975 3.165 32.455 3.175 ;
        RECT 32.130 2.700 32.430 3.165 ;
        RECT 33.520 3.145 34.255 3.495 ;
        RECT 34.555 3.165 35.295 3.495 ;
        RECT 36.415 3.475 36.775 3.480 ;
        RECT 34.555 3.155 34.885 3.165 ;
        RECT 36.255 3.145 36.985 3.475 ;
        RECT 33.520 3.140 33.870 3.145 ;
        RECT 36.415 3.140 36.775 3.145 ;
        RECT 37.720 2.700 38.060 3.940 ;
        RECT 45.955 3.705 46.290 4.055 ;
        RECT 46.665 4.040 46.985 4.055 ;
        RECT 46.665 3.705 47.005 4.040 ;
        RECT 47.665 3.815 48.445 4.155 ;
        RECT 47.870 3.810 48.445 3.815 ;
        RECT 48.105 3.805 48.445 3.810 ;
        RECT 48.115 3.775 48.445 3.805 ;
        RECT 52.980 3.940 53.340 4.365 ;
        RECT 60.025 4.265 60.755 4.595 ;
        RECT 61.215 4.245 61.535 4.625 ;
        RECT 61.215 4.055 61.545 4.245 ;
        RECT 61.945 4.055 62.245 4.845 ;
        RECT 63.130 4.155 63.430 4.845 ;
        RECT 63.845 4.795 64.185 4.845 ;
        RECT 75.595 4.600 75.895 5.550 ;
        RECT 78.390 5.145 78.690 5.550 ;
        RECT 90.855 5.550 93.950 5.770 ;
        RECT 79.115 5.145 79.445 5.155 ;
        RECT 77.205 4.845 79.445 5.145 ;
        RECT 75.515 4.595 75.895 4.600 ;
        RECT 47.235 3.175 47.965 3.505 ;
        RECT 48.780 3.495 49.130 3.500 ;
        RECT 47.235 3.165 47.715 3.175 ;
        RECT 32.130 2.400 38.060 2.700 ;
        RECT 47.390 2.700 47.690 3.165 ;
        RECT 48.780 3.145 49.515 3.495 ;
        RECT 49.815 3.165 50.555 3.495 ;
        RECT 51.675 3.475 52.035 3.480 ;
        RECT 49.815 3.155 50.145 3.165 ;
        RECT 51.515 3.145 52.245 3.475 ;
        RECT 48.780 3.140 49.130 3.145 ;
        RECT 51.675 3.140 52.035 3.145 ;
        RECT 52.980 2.700 53.320 3.940 ;
        RECT 61.215 3.705 61.550 4.055 ;
        RECT 61.925 4.040 62.245 4.055 ;
        RECT 61.925 3.705 62.265 4.040 ;
        RECT 62.925 3.815 63.705 4.155 ;
        RECT 63.130 3.810 63.705 3.815 ;
        RECT 63.365 3.805 63.705 3.810 ;
        RECT 63.375 3.775 63.705 3.805 ;
        RECT 68.240 3.940 68.600 4.365 ;
        RECT 75.285 4.265 76.015 4.595 ;
        RECT 76.475 4.245 76.795 4.625 ;
        RECT 76.475 4.055 76.805 4.245 ;
        RECT 77.205 4.055 77.505 4.845 ;
        RECT 78.390 4.155 78.690 4.845 ;
        RECT 79.105 4.795 79.445 4.845 ;
        RECT 90.855 4.600 91.155 5.550 ;
        RECT 93.650 5.145 93.950 5.550 ;
        RECT 94.375 5.145 94.705 5.155 ;
        RECT 92.465 4.845 94.705 5.145 ;
        RECT 90.775 4.595 91.155 4.600 ;
        RECT 62.495 3.175 63.225 3.505 ;
        RECT 64.040 3.495 64.390 3.500 ;
        RECT 62.495 3.165 62.975 3.175 ;
        RECT 47.390 2.400 53.320 2.700 ;
        RECT 62.650 2.700 62.950 3.165 ;
        RECT 64.040 3.145 64.775 3.495 ;
        RECT 65.075 3.165 65.815 3.495 ;
        RECT 66.935 3.475 67.295 3.480 ;
        RECT 65.075 3.155 65.405 3.165 ;
        RECT 66.775 3.145 67.505 3.475 ;
        RECT 64.040 3.140 64.390 3.145 ;
        RECT 66.935 3.140 67.295 3.145 ;
        RECT 68.240 2.700 68.580 3.940 ;
        RECT 76.475 3.705 76.810 4.055 ;
        RECT 77.185 4.040 77.505 4.055 ;
        RECT 77.185 3.705 77.525 4.040 ;
        RECT 78.185 3.815 78.965 4.155 ;
        RECT 78.390 3.810 78.965 3.815 ;
        RECT 78.625 3.805 78.965 3.810 ;
        RECT 78.635 3.775 78.965 3.805 ;
        RECT 83.500 3.940 83.860 4.365 ;
        RECT 90.545 4.265 91.275 4.595 ;
        RECT 91.735 4.245 92.055 4.625 ;
        RECT 91.735 4.055 92.065 4.245 ;
        RECT 92.465 4.055 92.765 4.845 ;
        RECT 93.650 4.155 93.950 4.845 ;
        RECT 94.365 4.795 94.705 4.845 ;
        RECT 77.755 3.175 78.485 3.505 ;
        RECT 79.300 3.495 79.650 3.500 ;
        RECT 77.755 3.165 78.235 3.175 ;
        RECT 62.650 2.400 68.580 2.700 ;
        RECT 77.910 2.700 78.210 3.165 ;
        RECT 79.300 3.145 80.035 3.495 ;
        RECT 80.335 3.165 81.075 3.495 ;
        RECT 82.195 3.475 82.555 3.480 ;
        RECT 80.335 3.155 80.665 3.165 ;
        RECT 82.035 3.145 82.765 3.475 ;
        RECT 79.300 3.140 79.650 3.145 ;
        RECT 82.195 3.140 82.555 3.145 ;
        RECT 83.500 2.700 83.840 3.940 ;
        RECT 91.735 3.705 92.070 4.055 ;
        RECT 92.445 4.040 92.765 4.055 ;
        RECT 92.445 3.705 92.785 4.040 ;
        RECT 93.445 3.815 94.225 4.155 ;
        RECT 93.650 3.810 94.225 3.815 ;
        RECT 93.885 3.805 94.225 3.810 ;
        RECT 93.895 3.775 94.225 3.805 ;
        RECT 98.760 3.940 99.120 4.365 ;
        RECT 93.015 3.175 93.745 3.505 ;
        RECT 94.560 3.495 94.910 3.500 ;
        RECT 93.015 3.165 93.495 3.175 ;
        RECT 77.910 2.400 83.840 2.700 ;
        RECT 93.170 2.700 93.470 3.165 ;
        RECT 94.560 3.145 95.295 3.495 ;
        RECT 95.595 3.165 96.335 3.495 ;
        RECT 97.455 3.475 97.815 3.480 ;
        RECT 95.595 3.155 95.925 3.165 ;
        RECT 97.295 3.145 98.025 3.475 ;
        RECT 94.560 3.140 94.910 3.145 ;
        RECT 97.455 3.140 97.815 3.145 ;
        RECT 98.760 2.700 99.100 3.940 ;
        RECT 93.170 2.400 99.100 2.700 ;
      LAYER met4 ;
        RECT 30.685 4.265 31.025 4.600 ;
        RECT 45.945 4.265 46.285 4.600 ;
        RECT 61.205 4.265 61.545 4.600 ;
        RECT 76.465 4.265 76.805 4.600 ;
        RECT 91.725 4.265 92.065 4.600 ;
        RECT 30.705 4.095 31.025 4.265 ;
        RECT 32.845 4.095 33.185 4.135 ;
        RECT 30.705 3.795 33.185 4.095 ;
        RECT 45.965 4.095 46.285 4.265 ;
        RECT 48.105 4.095 48.445 4.135 ;
        RECT 45.965 3.795 48.445 4.095 ;
        RECT 61.225 4.095 61.545 4.265 ;
        RECT 63.365 4.095 63.705 4.135 ;
        RECT 61.225 3.795 63.705 4.095 ;
        RECT 76.485 4.095 76.805 4.265 ;
        RECT 78.625 4.095 78.965 4.135 ;
        RECT 76.485 3.795 78.965 4.095 ;
        RECT 91.745 4.095 92.065 4.265 ;
        RECT 93.885 4.095 94.225 4.135 ;
        RECT 91.745 3.795 94.225 4.095 ;
        RECT 32.855 3.775 33.185 3.795 ;
        RECT 48.115 3.775 48.445 3.795 ;
        RECT 63.375 3.775 63.705 3.795 ;
        RECT 78.635 3.775 78.965 3.795 ;
        RECT 93.895 3.775 94.225 3.795 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r2
MACRO sky130_fd_sc_hd__conb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__conb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.775 0.085 1.115 0.745 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.275 1.910 0.605 2.635 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.605 1.740 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775 0.915 1.295 2.465 ;
    END
  END LO
END sky130_fd_sc_hd__conb_1
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.430000 ;
    PORT
      LAYER li1 ;
        RECT 2358.235 2253.225 2358.405 2254.495 ;
        RECT 2358.250 2161.235 2358.420 2162.505 ;
        RECT 2358.230 2056.235 2358.400 2057.505 ;
        RECT 2358.230 1951.240 2358.400 1952.510 ;
        RECT 2368.175 1788.240 2368.345 1789.510 ;
        RECT 2358.595 1708.225 2358.765 1709.495 ;
        RECT 2358.225 1608.235 2358.395 1609.505 ;
        RECT 2358.225 1531.235 2358.395 1532.505 ;
        RECT 2358.225 1433.240 2358.395 1434.510 ;
        RECT 2368.225 1333.240 2368.395 1334.510 ;
      LAYER met1 ;
        RECT 2358.490 2266.680 2358.810 2266.740 ;
        RECT 2900.830 2266.680 2901.150 2266.740 ;
        RECT 2358.490 2266.540 2901.150 2266.680 ;
        RECT 2358.490 2266.480 2358.810 2266.540 ;
        RECT 2900.830 2266.480 2901.150 2266.540 ;
        RECT 2358.175 2253.395 2358.470 2253.425 ;
        RECT 2358.175 2253.310 2358.635 2253.395 ;
        RECT 2358.120 2253.225 2358.635 2253.310 ;
        RECT 2358.120 2253.195 2358.470 2253.225 ;
        RECT 2358.120 2252.400 2358.260 2253.195 ;
        RECT 2358.490 2252.400 2358.810 2252.460 ;
        RECT 2358.120 2252.260 2358.810 2252.400 ;
        RECT 2358.490 2252.200 2358.810 2252.260 ;
        RECT 2358.060 2161.435 2358.320 2161.480 ;
        RECT 2358.060 2161.430 2358.480 2161.435 ;
        RECT 2358.060 2161.405 2358.485 2161.430 ;
        RECT 2358.060 2161.235 2358.650 2161.405 ;
        RECT 2358.060 2161.200 2358.485 2161.235 ;
        RECT 2358.060 2161.160 2358.320 2161.200 ;
        RECT 2358.170 2056.430 2358.460 2056.435 ;
        RECT 2358.170 2056.405 2358.465 2056.430 ;
        RECT 2358.170 2056.315 2358.630 2056.405 ;
        RECT 2356.190 2056.220 2356.510 2056.280 ;
        RECT 2358.120 2056.235 2358.630 2056.315 ;
        RECT 2358.120 2056.220 2358.465 2056.235 ;
        RECT 2356.190 2056.200 2358.465 2056.220 ;
        RECT 2356.190 2056.080 2358.260 2056.200 ;
        RECT 2356.190 2056.020 2356.510 2056.080 ;
        RECT 2356.190 1951.500 2356.510 1951.560 ;
        RECT 2356.190 1951.440 2358.260 1951.500 ;
        RECT 2356.190 1951.435 2358.460 1951.440 ;
        RECT 2356.190 1951.410 2358.465 1951.435 ;
        RECT 2356.190 1951.360 2358.630 1951.410 ;
        RECT 2356.190 1951.300 2356.510 1951.360 ;
        RECT 2358.120 1951.240 2358.630 1951.360 ;
        RECT 2358.120 1951.205 2358.465 1951.240 ;
        RECT 2358.120 1950.480 2358.260 1951.205 ;
        RECT 2358.490 1950.480 2358.810 1950.540 ;
        RECT 2358.120 1950.340 2358.810 1950.480 ;
        RECT 2358.490 1950.280 2358.810 1950.340 ;
        RECT 2368.115 1788.435 2368.405 1788.440 ;
        RECT 2368.115 1788.410 2368.410 1788.435 ;
        RECT 2368.115 1788.240 2368.575 1788.410 ;
        RECT 2368.115 1788.210 2368.410 1788.240 ;
        RECT 2368.120 1788.205 2368.410 1788.210 ;
        RECT 2358.490 1787.960 2358.810 1788.020 ;
        RECT 2368.240 1787.960 2368.380 1788.205 ;
        RECT 2358.490 1787.820 2368.380 1787.960 ;
        RECT 2358.490 1787.760 2358.810 1787.820 ;
        RECT 2358.490 1708.880 2358.810 1709.140 ;
        RECT 2356.190 1708.740 2356.510 1708.800 ;
        RECT 2358.580 1708.740 2358.720 1708.880 ;
        RECT 2356.190 1708.600 2358.720 1708.740 ;
        RECT 2356.190 1708.540 2356.510 1708.600 ;
        RECT 2358.580 1708.430 2358.720 1708.600 ;
        RECT 2358.540 1708.425 2358.830 1708.430 ;
        RECT 2358.535 1708.395 2358.830 1708.425 ;
        RECT 2358.535 1708.225 2358.995 1708.395 ;
        RECT 2358.535 1708.200 2358.830 1708.225 ;
        RECT 2358.535 1708.195 2358.825 1708.200 ;
        RECT 2358.165 1608.430 2358.455 1608.435 ;
        RECT 2358.165 1608.405 2358.460 1608.430 ;
        RECT 2358.165 1608.315 2358.625 1608.405 ;
        RECT 2358.120 1608.235 2358.625 1608.315 ;
        RECT 2358.120 1608.200 2358.460 1608.235 ;
        RECT 2356.190 1608.100 2356.510 1608.160 ;
        RECT 2358.120 1608.100 2358.260 1608.200 ;
        RECT 2356.190 1607.960 2358.260 1608.100 ;
        RECT 2356.190 1607.900 2356.510 1607.960 ;
        RECT 2356.190 1531.600 2356.510 1531.660 ;
        RECT 2356.190 1531.460 2358.260 1531.600 ;
        RECT 2356.190 1531.400 2356.510 1531.460 ;
        RECT 2358.120 1531.435 2358.260 1531.460 ;
        RECT 2358.120 1531.430 2358.455 1531.435 ;
        RECT 2358.120 1531.405 2358.460 1531.430 ;
        RECT 2358.120 1531.320 2358.625 1531.405 ;
        RECT 2358.165 1531.235 2358.625 1531.320 ;
        RECT 2358.165 1531.205 2358.460 1531.235 ;
        RECT 2358.170 1531.200 2358.460 1531.205 ;
        RECT 2358.140 1433.410 2358.480 1433.455 ;
        RECT 2356.190 1433.340 2356.510 1433.400 ;
        RECT 2358.140 1433.340 2358.625 1433.410 ;
        RECT 2356.190 1433.240 2358.625 1433.340 ;
        RECT 2356.190 1433.200 2358.480 1433.240 ;
        RECT 2356.190 1433.140 2356.510 1433.200 ;
        RECT 2358.120 1433.195 2358.480 1433.200 ;
        RECT 2358.120 1432.660 2358.260 1433.195 ;
        RECT 2358.490 1432.660 2358.810 1432.720 ;
        RECT 2358.120 1432.520 2358.810 1432.660 ;
        RECT 2358.490 1432.460 2358.810 1432.520 ;
        RECT 2358.490 1345.620 2358.810 1345.680 ;
        RECT 2368.150 1345.620 2368.470 1345.680 ;
        RECT 2358.490 1345.480 2368.470 1345.620 ;
        RECT 2358.490 1345.420 2358.810 1345.480 ;
        RECT 2368.150 1345.420 2368.470 1345.480 ;
        RECT 2368.150 1333.410 2368.470 1333.455 ;
        RECT 2368.150 1333.240 2368.625 1333.410 ;
        RECT 2368.150 1333.195 2368.470 1333.240 ;
      LAYER met2 ;
        RECT 2900.850 2290.395 2901.130 2290.765 ;
        RECT 2900.920 2266.770 2901.060 2290.395 ;
        RECT 2358.520 2266.450 2358.780 2266.770 ;
        RECT 2900.860 2266.450 2901.120 2266.770 ;
        RECT 2358.580 2252.490 2358.720 2266.450 ;
        RECT 2358.520 2252.170 2358.780 2252.490 ;
        RECT 2358.580 2208.070 2358.720 2252.170 ;
        RECT 2358.120 2207.930 2358.720 2208.070 ;
        RECT 2358.120 2161.480 2358.260 2207.930 ;
        RECT 2358.060 2161.160 2358.320 2161.480 ;
        RECT 2358.120 2159.770 2358.260 2161.160 ;
        RECT 2356.280 2159.630 2358.260 2159.770 ;
        RECT 2356.280 2056.310 2356.420 2159.630 ;
        RECT 2356.220 2055.990 2356.480 2056.310 ;
        RECT 2356.280 1951.590 2356.420 2055.990 ;
        RECT 2356.220 1951.270 2356.480 1951.590 ;
        RECT 2358.520 1950.250 2358.780 1950.570 ;
        RECT 2358.580 1788.050 2358.720 1950.250 ;
        RECT 2358.520 1787.730 2358.780 1788.050 ;
        RECT 2358.580 1773.370 2358.720 1787.730 ;
        RECT 2358.580 1773.230 2359.640 1773.370 ;
        RECT 2359.500 1725.070 2359.640 1773.230 ;
        RECT 2358.580 1724.930 2359.640 1725.070 ;
        RECT 2358.580 1709.170 2358.720 1724.930 ;
        RECT 2358.520 1708.850 2358.780 1709.170 ;
        RECT 2356.220 1708.510 2356.480 1708.830 ;
        RECT 2356.280 1608.190 2356.420 1708.510 ;
        RECT 2356.220 1607.870 2356.480 1608.190 ;
        RECT 2356.280 1531.690 2356.420 1607.870 ;
        RECT 2356.220 1531.370 2356.480 1531.690 ;
        RECT 2356.280 1433.430 2356.420 1531.370 ;
        RECT 2356.220 1433.110 2356.480 1433.430 ;
        RECT 2358.520 1432.430 2358.780 1432.750 ;
        RECT 2358.580 1345.710 2358.720 1432.430 ;
        RECT 2358.520 1345.390 2358.780 1345.710 ;
        RECT 2368.180 1345.390 2368.440 1345.710 ;
        RECT 2368.240 1333.485 2368.380 1345.390 ;
        RECT 2368.180 1333.165 2368.440 1333.485 ;
      LAYER met3 ;
        RECT 2900.825 2290.730 2901.155 2290.745 ;
        RECT 2917.600 2290.730 2924.800 2291.180 ;
        RECT 2900.825 2290.430 2924.800 2290.730 ;
        RECT 2900.825 2290.415 2901.155 2290.430 ;
        RECT 2917.600 2289.980 2924.800 2290.430 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.065000 ;
    PORT
      LAYER li1 ;
        RECT 2697.325 2215.595 2697.685 2216.175 ;
        RECT 2697.325 2035.595 2697.685 2036.175 ;
        RECT 2697.325 1855.595 2697.685 1856.175 ;
        RECT 2697.325 1675.595 2697.685 1676.175 ;
        RECT 2697.325 1495.595 2697.685 1496.175 ;
      LAYER met1 ;
        RECT 2696.970 2216.140 2697.290 2216.200 ;
        RECT 2697.445 2216.140 2697.735 2216.185 ;
        RECT 2696.970 2216.000 2697.735 2216.140 ;
        RECT 2696.970 2215.940 2697.290 2216.000 ;
        RECT 2697.445 2215.955 2697.735 2216.000 ;
        RECT 2696.970 2036.140 2697.290 2036.200 ;
        RECT 2697.445 2036.140 2697.735 2036.185 ;
        RECT 2696.970 2036.000 2697.735 2036.140 ;
        RECT 2696.970 2035.940 2697.290 2036.000 ;
        RECT 2697.445 2035.955 2697.735 2036.000 ;
        RECT 2696.970 1856.140 2697.290 1856.200 ;
        RECT 2697.445 1856.140 2697.735 1856.185 ;
        RECT 2696.970 1856.000 2697.735 1856.140 ;
        RECT 2696.970 1855.940 2697.290 1856.000 ;
        RECT 2697.445 1855.955 2697.735 1856.000 ;
        RECT 2696.970 1676.140 2697.290 1676.200 ;
        RECT 2697.445 1676.140 2697.735 1676.185 ;
        RECT 2696.970 1676.000 2697.735 1676.140 ;
        RECT 2696.970 1675.940 2697.290 1676.000 ;
        RECT 2697.445 1675.955 2697.735 1676.000 ;
        RECT 2696.970 1496.140 2697.290 1496.200 ;
        RECT 2697.445 1496.140 2697.735 1496.185 ;
        RECT 2696.970 1496.000 2697.735 1496.140 ;
        RECT 2696.970 1495.940 2697.290 1496.000 ;
        RECT 2697.445 1495.955 2697.735 1496.000 ;
      LAYER met2 ;
        RECT 2904.070 2556.275 2904.350 2556.645 ;
        RECT 2904.140 2239.085 2904.280 2556.275 ;
        RECT 2696.150 2238.715 2696.430 2239.085 ;
        RECT 2904.070 2238.715 2904.350 2239.085 ;
        RECT 2696.220 2229.000 2696.360 2238.715 ;
        RECT 2696.070 2228.770 2696.360 2229.000 ;
        RECT 2693.460 2228.700 2696.360 2228.770 ;
        RECT 2693.460 2228.630 2696.350 2228.700 ;
        RECT 2693.460 2111.470 2693.600 2228.630 ;
        RECT 2696.070 2225.490 2696.350 2228.630 ;
        RECT 2696.070 2225.350 2697.200 2225.490 ;
        RECT 2696.070 2225.000 2696.350 2225.350 ;
        RECT 2697.060 2216.230 2697.200 2225.350 ;
        RECT 2697.000 2215.910 2697.260 2216.230 ;
        RECT 2693.460 2111.330 2694.520 2111.470 ;
        RECT 2694.380 2045.850 2694.520 2111.330 ;
        RECT 2696.070 2045.850 2696.350 2049.000 ;
        RECT 2693.920 2045.710 2696.350 2045.850 ;
        RECT 2693.920 1966.570 2694.060 2045.710 ;
        RECT 2696.070 2045.490 2696.350 2045.710 ;
        RECT 2696.070 2045.350 2697.200 2045.490 ;
        RECT 2696.070 2045.000 2696.350 2045.350 ;
        RECT 2697.060 2036.230 2697.200 2045.350 ;
        RECT 2697.000 2035.910 2697.260 2036.230 ;
        RECT 2693.460 1966.430 2694.060 1966.570 ;
        RECT 2693.460 1918.270 2693.600 1966.430 ;
        RECT 2693.460 1918.130 2694.060 1918.270 ;
        RECT 2693.920 1866.330 2694.060 1918.130 ;
        RECT 2696.070 1866.330 2696.350 1869.000 ;
        RECT 2693.920 1866.190 2696.350 1866.330 ;
        RECT 2693.920 1773.370 2694.060 1866.190 ;
        RECT 2696.070 1865.490 2696.350 1866.190 ;
        RECT 2696.070 1865.350 2697.200 1865.490 ;
        RECT 2696.070 1865.000 2696.350 1865.350 ;
        RECT 2697.060 1856.230 2697.200 1865.350 ;
        RECT 2697.000 1855.910 2697.260 1856.230 ;
        RECT 2693.460 1773.230 2694.060 1773.370 ;
        RECT 2693.460 1725.070 2693.600 1773.230 ;
        RECT 2693.460 1724.930 2694.520 1725.070 ;
        RECT 2694.380 1688.850 2694.520 1724.930 ;
        RECT 2696.070 1688.850 2696.350 1689.000 ;
        RECT 2693.920 1688.710 2696.350 1688.850 ;
        RECT 2693.920 1580.170 2694.060 1688.710 ;
        RECT 2696.070 1685.490 2696.350 1688.710 ;
        RECT 2696.070 1685.350 2697.200 1685.490 ;
        RECT 2696.070 1685.000 2696.350 1685.350 ;
        RECT 2697.060 1676.230 2697.200 1685.350 ;
        RECT 2697.000 1675.910 2697.260 1676.230 ;
        RECT 2693.920 1580.030 2694.520 1580.170 ;
        RECT 2694.380 1508.650 2694.520 1580.030 ;
        RECT 2696.070 1508.650 2696.350 1509.000 ;
        RECT 2694.380 1508.510 2696.350 1508.650 ;
        RECT 2696.070 1505.490 2696.350 1508.510 ;
        RECT 2696.070 1505.350 2697.200 1505.490 ;
        RECT 2696.070 1505.000 2696.350 1505.350 ;
        RECT 2697.060 1496.230 2697.200 1505.350 ;
        RECT 2697.000 1495.910 2697.260 1496.230 ;
      LAYER met3 ;
        RECT 2904.045 2556.610 2904.375 2556.625 ;
        RECT 2917.600 2556.610 2924.800 2557.060 ;
        RECT 2904.045 2556.310 2924.800 2556.610 ;
        RECT 2904.045 2556.295 2904.375 2556.310 ;
        RECT 2917.600 2555.860 2924.800 2556.310 ;
        RECT 2696.125 2239.050 2696.455 2239.065 ;
        RECT 2904.045 2239.050 2904.375 2239.065 ;
        RECT 2696.125 2238.750 2904.375 2239.050 ;
        RECT 2696.125 2238.735 2696.455 2238.750 ;
        RECT 2904.045 2238.735 2904.375 2238.750 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 2708.945 2215.565 2709.300 2215.935 ;
        RECT 2708.945 2035.565 2709.300 2035.935 ;
        RECT 2708.945 1855.565 2709.300 1855.935 ;
        RECT 2708.945 1675.565 2709.300 1675.935 ;
        RECT 2708.945 1495.565 2709.300 1495.935 ;
      LAYER met1 ;
        RECT 2708.470 2215.800 2708.790 2215.860 ;
        RECT 2708.945 2215.800 2709.235 2215.845 ;
        RECT 2708.470 2215.660 2709.235 2215.800 ;
        RECT 2708.470 2215.600 2708.790 2215.660 ;
        RECT 2708.945 2215.615 2709.235 2215.660 ;
        RECT 2708.470 2035.800 2708.790 2035.860 ;
        RECT 2708.945 2035.800 2709.235 2035.845 ;
        RECT 2708.470 2035.660 2709.235 2035.800 ;
        RECT 2708.470 2035.600 2708.790 2035.660 ;
        RECT 2708.945 2035.615 2709.235 2035.660 ;
        RECT 2708.470 1855.800 2708.790 1855.860 ;
        RECT 2708.945 1855.800 2709.235 1855.845 ;
        RECT 2708.470 1855.660 2709.235 1855.800 ;
        RECT 2708.470 1855.600 2708.790 1855.660 ;
        RECT 2708.945 1855.615 2709.235 1855.660 ;
        RECT 2708.470 1675.800 2708.790 1675.860 ;
        RECT 2708.945 1675.800 2709.235 1675.845 ;
        RECT 2708.470 1675.660 2709.235 1675.800 ;
        RECT 2708.470 1675.600 2708.790 1675.660 ;
        RECT 2708.945 1675.615 2709.235 1675.660 ;
        RECT 2708.470 1495.800 2708.790 1495.860 ;
        RECT 2708.945 1495.800 2709.235 1495.845 ;
        RECT 2708.470 1495.660 2709.235 1495.800 ;
        RECT 2708.470 1495.600 2708.790 1495.660 ;
        RECT 2708.945 1495.615 2709.235 1495.660 ;
      LAYER met2 ;
        RECT 2903.150 2821.475 2903.430 2821.845 ;
        RECT 2903.220 2236.365 2903.360 2821.475 ;
        RECT 2708.570 2235.995 2708.850 2236.365 ;
        RECT 2903.150 2235.995 2903.430 2236.365 ;
        RECT 2708.640 2229.000 2708.780 2235.995 ;
        RECT 2708.490 2226.845 2708.780 2229.000 ;
        RECT 2708.490 2226.475 2708.850 2226.845 ;
        RECT 2708.490 2225.000 2708.770 2226.475 ;
        RECT 2708.560 2215.890 2708.700 2225.000 ;
        RECT 2708.500 2215.570 2708.760 2215.890 ;
        RECT 2708.490 2046.645 2708.770 2049.000 ;
        RECT 2708.490 2046.275 2708.850 2046.645 ;
        RECT 2708.490 2045.000 2708.770 2046.275 ;
        RECT 2708.560 2035.890 2708.700 2045.000 ;
        RECT 2708.500 2035.570 2708.760 2035.890 ;
        RECT 2708.490 1865.765 2708.770 1869.000 ;
        RECT 2708.490 1865.395 2708.850 1865.765 ;
        RECT 2708.490 1865.000 2708.770 1865.395 ;
        RECT 2708.560 1855.890 2708.700 1865.000 ;
        RECT 2708.500 1855.570 2708.760 1855.890 ;
        RECT 2708.570 1697.435 2708.850 1697.805 ;
        RECT 2708.640 1689.000 2708.780 1697.435 ;
        RECT 2708.490 1688.780 2708.780 1689.000 ;
        RECT 2708.490 1685.000 2708.770 1688.780 ;
        RECT 2708.560 1675.890 2708.700 1685.000 ;
        RECT 2708.500 1675.570 2708.760 1675.890 ;
        RECT 2708.570 1518.595 2708.850 1518.965 ;
        RECT 2708.640 1509.000 2708.780 1518.595 ;
        RECT 2708.490 1508.580 2708.780 1509.000 ;
        RECT 2708.490 1505.000 2708.770 1508.580 ;
        RECT 2708.560 1495.890 2708.700 1505.000 ;
        RECT 2708.500 1495.570 2708.760 1495.890 ;
      LAYER met3 ;
        RECT 2903.125 2821.810 2903.455 2821.825 ;
        RECT 2917.600 2821.810 2924.800 2822.260 ;
        RECT 2903.125 2821.510 2924.800 2821.810 ;
        RECT 2903.125 2821.495 2903.455 2821.510 ;
        RECT 2917.600 2821.060 2924.800 2821.510 ;
        RECT 2708.545 2236.330 2708.875 2236.345 ;
        RECT 2903.125 2236.330 2903.455 2236.345 ;
        RECT 2708.545 2236.030 2903.455 2236.330 ;
        RECT 2708.545 2236.015 2708.875 2236.030 ;
        RECT 2903.125 2236.015 2903.455 2236.030 ;
        RECT 2707.830 2226.810 2708.210 2226.820 ;
        RECT 2708.545 2226.810 2708.875 2226.825 ;
        RECT 2707.830 2226.510 2708.875 2226.810 ;
        RECT 2707.830 2226.500 2708.210 2226.510 ;
        RECT 2708.545 2226.495 2708.875 2226.510 ;
        RECT 2707.830 2046.610 2708.210 2046.620 ;
        RECT 2708.545 2046.610 2708.875 2046.625 ;
        RECT 2707.830 2046.310 2708.875 2046.610 ;
        RECT 2707.830 2046.300 2708.210 2046.310 ;
        RECT 2708.545 2046.295 2708.875 2046.310 ;
        RECT 2707.830 1865.730 2708.210 1865.740 ;
        RECT 2708.545 1865.730 2708.875 1865.745 ;
        RECT 2707.830 1865.430 2708.875 1865.730 ;
        RECT 2707.830 1865.420 2708.210 1865.430 ;
        RECT 2708.545 1865.415 2708.875 1865.430 ;
        RECT 2707.830 1697.770 2708.210 1697.780 ;
        RECT 2708.545 1697.770 2708.875 1697.785 ;
        RECT 2707.830 1697.470 2708.875 1697.770 ;
        RECT 2707.830 1697.460 2708.210 1697.470 ;
        RECT 2708.545 1697.455 2708.875 1697.470 ;
        RECT 2707.830 1518.930 2708.210 1518.940 ;
        RECT 2708.545 1518.930 2708.875 1518.945 ;
        RECT 2707.830 1518.630 2708.875 1518.930 ;
        RECT 2707.830 1518.620 2708.210 1518.630 ;
        RECT 2708.545 1518.615 2708.875 1518.630 ;
      LAYER met4 ;
        RECT 2707.855 2226.495 2708.185 2226.825 ;
        RECT 2707.870 2046.625 2708.170 2226.495 ;
        RECT 2707.855 2046.295 2708.185 2046.625 ;
        RECT 2707.870 1865.745 2708.170 2046.295 ;
        RECT 2707.855 1865.415 2708.185 1865.745 ;
        RECT 2707.870 1697.785 2708.170 1865.415 ;
        RECT 2707.855 1697.455 2708.185 1697.785 ;
        RECT 2707.870 1518.945 2708.170 1697.455 ;
        RECT 2707.855 1518.615 2708.185 1518.945 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.065000 ;
    PORT
      LAYER li1 ;
        RECT 2722.795 2215.595 2723.155 2216.175 ;
        RECT 2722.795 2035.595 2723.155 2036.175 ;
        RECT 2722.795 1855.595 2723.155 1856.175 ;
        RECT 2722.795 1675.595 2723.155 1676.175 ;
        RECT 2722.795 1495.595 2723.155 1496.175 ;
      LAYER met1 ;
        RECT 2720.890 2216.140 2721.210 2216.200 ;
        RECT 2722.745 2216.140 2723.035 2216.185 ;
        RECT 2720.890 2216.000 2723.035 2216.140 ;
        RECT 2720.890 2215.940 2721.210 2216.000 ;
        RECT 2722.745 2215.955 2723.035 2216.000 ;
        RECT 2720.890 2036.140 2721.210 2036.200 ;
        RECT 2722.745 2036.140 2723.035 2036.185 ;
        RECT 2720.890 2036.000 2723.035 2036.140 ;
        RECT 2720.890 2035.940 2721.210 2036.000 ;
        RECT 2722.745 2035.955 2723.035 2036.000 ;
        RECT 2720.890 1856.140 2721.210 1856.200 ;
        RECT 2722.745 1856.140 2723.035 1856.185 ;
        RECT 2720.890 1856.000 2723.035 1856.140 ;
        RECT 2720.890 1855.940 2721.210 1856.000 ;
        RECT 2722.745 1855.955 2723.035 1856.000 ;
        RECT 2720.890 1676.140 2721.210 1676.200 ;
        RECT 2722.745 1676.140 2723.035 1676.185 ;
        RECT 2720.890 1676.000 2723.035 1676.140 ;
        RECT 2720.890 1675.940 2721.210 1676.000 ;
        RECT 2722.745 1675.955 2723.035 1676.000 ;
        RECT 2720.890 1496.140 2721.210 1496.200 ;
        RECT 2722.745 1496.140 2723.035 1496.185 ;
        RECT 2720.890 1496.000 2723.035 1496.140 ;
        RECT 2720.890 1495.940 2721.210 1496.000 ;
        RECT 2722.745 1495.955 2723.035 1496.000 ;
      LAYER met2 ;
        RECT 2902.230 3087.355 2902.510 3087.725 ;
        RECT 2902.300 2239.765 2902.440 3087.355 ;
        RECT 2720.990 2239.395 2721.270 2239.765 ;
        RECT 2902.230 2239.395 2902.510 2239.765 ;
        RECT 2721.060 2229.000 2721.200 2239.395 ;
        RECT 2720.910 2228.885 2721.200 2229.000 ;
        RECT 2720.910 2228.515 2721.270 2228.885 ;
        RECT 2720.910 2225.000 2721.190 2228.515 ;
        RECT 2720.980 2216.230 2721.120 2225.000 ;
        RECT 2720.920 2215.910 2721.180 2216.230 ;
        RECT 2720.910 2046.530 2721.190 2049.000 ;
        RECT 2721.450 2046.530 2721.730 2046.645 ;
        RECT 2720.910 2046.390 2721.730 2046.530 ;
        RECT 2720.910 2045.000 2721.190 2046.390 ;
        RECT 2721.450 2046.275 2721.730 2046.390 ;
        RECT 2720.980 2036.230 2721.120 2045.000 ;
        RECT 2720.920 2035.910 2721.180 2036.230 ;
        RECT 2720.910 1865.765 2721.190 1869.000 ;
        RECT 2720.910 1865.395 2721.270 1865.765 ;
        RECT 2720.910 1865.000 2721.190 1865.395 ;
        RECT 2720.980 1856.230 2721.120 1865.000 ;
        RECT 2720.920 1855.910 2721.180 1856.230 ;
        RECT 2720.990 1697.435 2721.270 1697.805 ;
        RECT 2721.060 1689.000 2721.200 1697.435 ;
        RECT 2720.910 1688.780 2721.200 1689.000 ;
        RECT 2720.910 1685.000 2721.190 1688.780 ;
        RECT 2720.980 1676.230 2721.120 1685.000 ;
        RECT 2720.920 1675.910 2721.180 1676.230 ;
        RECT 2720.990 1518.595 2721.270 1518.965 ;
        RECT 2721.060 1509.000 2721.200 1518.595 ;
        RECT 2720.910 1508.580 2721.200 1509.000 ;
        RECT 2720.910 1505.000 2721.190 1508.580 ;
        RECT 2720.980 1496.230 2721.120 1505.000 ;
        RECT 2720.920 1495.910 2721.180 1496.230 ;
      LAYER met3 ;
        RECT 2902.205 3087.690 2902.535 3087.705 ;
        RECT 2917.600 3087.690 2924.800 3088.140 ;
        RECT 2902.205 3087.390 2924.800 3087.690 ;
        RECT 2902.205 3087.375 2902.535 3087.390 ;
        RECT 2917.600 3086.940 2924.800 3087.390 ;
        RECT 2720.965 2239.730 2721.295 2239.745 ;
        RECT 2902.205 2239.730 2902.535 2239.745 ;
        RECT 2720.965 2239.430 2902.535 2239.730 ;
        RECT 2720.965 2239.415 2721.295 2239.430 ;
        RECT 2902.205 2239.415 2902.535 2239.430 ;
        RECT 2720.965 2228.850 2721.295 2228.865 ;
        RECT 2721.630 2228.850 2722.010 2228.860 ;
        RECT 2720.965 2228.550 2722.010 2228.850 ;
        RECT 2720.965 2228.535 2721.295 2228.550 ;
        RECT 2721.630 2228.540 2722.010 2228.550 ;
        RECT 2721.425 2046.620 2721.755 2046.625 ;
        RECT 2721.425 2046.610 2722.010 2046.620 ;
        RECT 2721.200 2046.310 2722.010 2046.610 ;
        RECT 2721.425 2046.300 2722.010 2046.310 ;
        RECT 2721.425 2046.295 2721.755 2046.300 ;
        RECT 2720.965 1865.730 2721.295 1865.745 ;
        RECT 2721.630 1865.730 2722.010 1865.740 ;
        RECT 2720.965 1865.430 2722.010 1865.730 ;
        RECT 2720.965 1865.415 2721.295 1865.430 ;
        RECT 2721.630 1865.420 2722.010 1865.430 ;
        RECT 2720.965 1697.770 2721.295 1697.785 ;
        RECT 2721.630 1697.770 2722.010 1697.780 ;
        RECT 2720.965 1697.470 2722.010 1697.770 ;
        RECT 2720.965 1697.455 2721.295 1697.470 ;
        RECT 2721.630 1697.460 2722.010 1697.470 ;
        RECT 2720.965 1518.930 2721.295 1518.945 ;
        RECT 2721.630 1518.930 2722.010 1518.940 ;
        RECT 2720.965 1518.630 2722.010 1518.930 ;
        RECT 2720.965 1518.615 2721.295 1518.630 ;
        RECT 2721.630 1518.620 2722.010 1518.630 ;
      LAYER met4 ;
        RECT 2721.655 2228.535 2721.985 2228.865 ;
        RECT 2721.670 2046.625 2721.970 2228.535 ;
        RECT 2721.655 2046.295 2721.985 2046.625 ;
        RECT 2721.670 1865.745 2721.970 2046.295 ;
        RECT 2721.655 1865.415 2721.985 1865.745 ;
        RECT 2721.670 1697.785 2721.970 1865.415 ;
        RECT 2721.655 1697.455 2721.985 1697.785 ;
        RECT 2721.670 1518.945 2721.970 1697.455 ;
        RECT 2721.655 1518.615 2721.985 1518.945 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.982500 ;
    PORT
      LAYER li1 ;
        RECT 2732.335 2215.565 2732.675 2215.935 ;
        RECT 2732.335 2035.565 2732.675 2035.935 ;
        RECT 2732.335 1855.565 2732.675 1855.935 ;
        RECT 2732.335 1675.565 2732.675 1675.935 ;
        RECT 2732.335 1495.565 2732.675 1495.935 ;
      LAYER met1 ;
        RECT 2734.770 2225.880 2735.090 2225.940 ;
        RECT 2737.530 2225.880 2737.850 2225.940 ;
        RECT 2734.770 2225.740 2737.850 2225.880 ;
        RECT 2734.770 2225.680 2735.090 2225.740 ;
        RECT 2737.530 2225.680 2737.850 2225.740 ;
        RECT 2732.850 2216.280 2733.170 2216.540 ;
        RECT 2732.405 2215.800 2732.695 2215.845 ;
        RECT 2732.940 2215.800 2733.080 2216.280 ;
        RECT 2732.405 2215.660 2733.080 2215.800 ;
        RECT 2732.405 2215.615 2732.695 2215.660 ;
        RECT 2736.150 2040.920 2736.470 2040.980 ;
        RECT 2737.530 2040.920 2737.850 2040.980 ;
        RECT 2736.150 2040.780 2737.850 2040.920 ;
        RECT 2736.150 2040.720 2736.470 2040.780 ;
        RECT 2737.530 2040.720 2737.850 2040.780 ;
        RECT 2732.850 2036.280 2733.170 2036.540 ;
        RECT 2732.405 2035.800 2732.695 2035.845 ;
        RECT 2732.940 2035.800 2733.080 2036.280 ;
        RECT 2732.405 2035.660 2733.080 2035.800 ;
        RECT 2732.405 2035.615 2732.695 2035.660 ;
        RECT 2735.230 1866.500 2735.550 1866.560 ;
        RECT 2737.530 1866.500 2737.850 1866.560 ;
        RECT 2735.230 1866.360 2737.850 1866.500 ;
        RECT 2735.230 1866.300 2735.550 1866.360 ;
        RECT 2737.530 1866.300 2737.850 1866.360 ;
        RECT 2732.850 1856.280 2733.170 1856.540 ;
        RECT 2732.405 1855.800 2732.695 1855.845 ;
        RECT 2732.940 1855.800 2733.080 1856.280 ;
        RECT 2732.405 1855.660 2733.080 1855.800 ;
        RECT 2732.405 1855.615 2732.695 1855.660 ;
        RECT 2735.690 1725.060 2736.010 1725.120 ;
        RECT 2737.530 1725.060 2737.850 1725.120 ;
        RECT 2735.690 1724.920 2737.850 1725.060 ;
        RECT 2735.690 1724.860 2736.010 1724.920 ;
        RECT 2737.530 1724.860 2737.850 1724.920 ;
        RECT 2734.770 1688.680 2735.090 1688.740 ;
        RECT 2737.530 1688.680 2737.850 1688.740 ;
        RECT 2734.770 1688.540 2737.850 1688.680 ;
        RECT 2734.770 1688.480 2735.090 1688.540 ;
        RECT 2737.530 1688.480 2737.850 1688.540 ;
        RECT 2732.850 1676.280 2733.170 1676.540 ;
        RECT 2732.405 1675.800 2732.695 1675.845 ;
        RECT 2732.940 1675.800 2733.080 1676.280 ;
        RECT 2732.405 1675.660 2733.080 1675.800 ;
        RECT 2732.405 1675.615 2732.695 1675.660 ;
        RECT 2735.230 1518.680 2735.550 1518.740 ;
        RECT 2737.530 1518.680 2737.850 1518.740 ;
        RECT 2735.230 1518.540 2737.850 1518.680 ;
        RECT 2735.230 1518.480 2735.550 1518.540 ;
        RECT 2737.530 1518.480 2737.850 1518.540 ;
        RECT 2732.850 1496.280 2733.170 1496.540 ;
        RECT 2732.405 1495.800 2732.695 1495.845 ;
        RECT 2732.940 1495.800 2733.080 1496.280 ;
        RECT 2732.405 1495.660 2733.080 1495.800 ;
        RECT 2732.405 1495.615 2732.695 1495.660 ;
      LAYER met2 ;
        RECT 2901.310 3353.235 2901.590 3353.605 ;
        RECT 2901.380 2240.445 2901.520 3353.235 ;
        RECT 2733.410 2240.075 2733.690 2240.445 ;
        RECT 2901.310 2240.075 2901.590 2240.445 ;
        RECT 2733.480 2229.000 2733.620 2240.075 ;
        RECT 2733.330 2228.770 2733.620 2229.000 ;
        RECT 2733.330 2228.630 2735.000 2228.770 ;
        RECT 2733.330 2225.490 2733.610 2228.630 ;
        RECT 2734.860 2225.970 2735.000 2228.630 ;
        RECT 2734.800 2225.650 2735.060 2225.970 ;
        RECT 2737.560 2225.650 2737.820 2225.970 ;
        RECT 2732.940 2225.350 2733.610 2225.490 ;
        RECT 2732.940 2216.570 2733.080 2225.350 ;
        RECT 2733.330 2225.000 2733.610 2225.350 ;
        RECT 2732.880 2216.250 2733.140 2216.570 ;
        RECT 2733.330 2045.850 2733.610 2049.000 ;
        RECT 2733.330 2045.710 2736.380 2045.850 ;
        RECT 2733.330 2045.490 2733.610 2045.710 ;
        RECT 2732.940 2045.350 2733.610 2045.490 ;
        RECT 2732.940 2036.570 2733.080 2045.350 ;
        RECT 2733.330 2045.000 2733.610 2045.350 ;
        RECT 2736.240 2041.010 2736.380 2045.710 ;
        RECT 2737.620 2041.010 2737.760 2225.650 ;
        RECT 2736.180 2040.690 2736.440 2041.010 ;
        RECT 2737.560 2040.690 2737.820 2041.010 ;
        RECT 2732.880 2036.250 2733.140 2036.570 ;
        RECT 2733.330 1867.010 2733.610 1869.000 ;
        RECT 2733.330 1866.870 2735.460 1867.010 ;
        RECT 2733.330 1865.490 2733.610 1866.870 ;
        RECT 2735.320 1866.590 2735.460 1866.870 ;
        RECT 2737.620 1866.590 2737.760 2040.690 ;
        RECT 2735.260 1866.270 2735.520 1866.590 ;
        RECT 2737.560 1866.270 2737.820 1866.590 ;
        RECT 2732.940 1865.350 2733.610 1865.490 ;
        RECT 2732.940 1856.570 2733.080 1865.350 ;
        RECT 2733.330 1865.000 2733.610 1865.350 ;
        RECT 2732.880 1856.250 2733.140 1856.570 ;
        RECT 2737.620 1725.150 2737.760 1866.270 ;
        RECT 2735.720 1725.070 2735.980 1725.150 ;
        RECT 2734.860 1724.930 2735.980 1725.070 ;
        RECT 2733.330 1688.850 2733.610 1689.000 ;
        RECT 2734.860 1688.850 2735.000 1724.930 ;
        RECT 2735.720 1724.830 2735.980 1724.930 ;
        RECT 2737.560 1724.830 2737.820 1725.150 ;
        RECT 2733.330 1688.770 2735.000 1688.850 ;
        RECT 2733.330 1688.710 2735.060 1688.770 ;
        RECT 2733.330 1685.490 2733.610 1688.710 ;
        RECT 2734.800 1688.450 2735.060 1688.710 ;
        RECT 2737.560 1688.450 2737.820 1688.770 ;
        RECT 2732.940 1685.350 2733.610 1685.490 ;
        RECT 2732.940 1676.570 2733.080 1685.350 ;
        RECT 2733.330 1685.000 2733.610 1685.350 ;
        RECT 2732.880 1676.250 2733.140 1676.570 ;
        RECT 2737.620 1518.770 2737.760 1688.450 ;
        RECT 2735.260 1518.450 2735.520 1518.770 ;
        RECT 2737.560 1518.450 2737.820 1518.770 ;
        RECT 2733.330 1508.650 2733.610 1509.000 ;
        RECT 2735.320 1508.650 2735.460 1518.450 ;
        RECT 2733.330 1508.510 2735.460 1508.650 ;
        RECT 2733.330 1505.490 2733.610 1508.510 ;
        RECT 2732.940 1505.350 2733.610 1505.490 ;
        RECT 2732.940 1496.570 2733.080 1505.350 ;
        RECT 2733.330 1505.000 2733.610 1505.350 ;
        RECT 2732.880 1496.250 2733.140 1496.570 ;
      LAYER met3 ;
        RECT 2901.285 3353.570 2901.615 3353.585 ;
        RECT 2917.600 3353.570 2924.800 3354.020 ;
        RECT 2901.285 3353.270 2924.800 3353.570 ;
        RECT 2901.285 3353.255 2901.615 3353.270 ;
        RECT 2917.600 3352.820 2924.800 3353.270 ;
        RECT 2733.385 2240.410 2733.715 2240.425 ;
        RECT 2901.285 2240.410 2901.615 2240.425 ;
        RECT 2733.385 2240.110 2901.615 2240.410 ;
        RECT 2733.385 2240.095 2733.715 2240.110 ;
        RECT 2901.285 2240.095 2901.615 2240.110 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.289999 ;
    PORT
      LAYER li1 ;
        RECT 2361.465 2253.225 2361.635 2254.495 ;
        RECT 2372.690 2253.230 2372.860 2254.500 ;
        RECT 2372.690 2247.960 2372.860 2249.230 ;
        RECT 2361.660 2161.225 2361.830 2162.495 ;
        RECT 2373.345 2161.465 2373.515 2162.505 ;
        RECT 2373.340 2161.225 2373.520 2161.465 ;
        RECT 2373.345 2155.955 2373.515 2157.225 ;
        RECT 2366.810 2056.235 2366.980 2057.505 ;
        RECT 2372.425 2056.235 2372.595 2057.505 ;
        RECT 2372.425 2050.955 2372.595 2052.225 ;
        RECT 2369.045 1951.240 2369.215 1952.510 ;
        RECT 2374.660 1951.240 2374.830 1952.510 ;
        RECT 2374.660 1945.955 2374.830 1947.225 ;
        RECT 2375.690 1788.240 2375.860 1789.510 ;
        RECT 2381.305 1788.240 2381.475 1789.510 ;
        RECT 2381.305 1782.955 2381.475 1784.225 ;
        RECT 2361.825 1708.225 2361.995 1709.495 ;
        RECT 2373.050 1708.230 2373.220 1709.500 ;
        RECT 2373.050 1702.960 2373.220 1704.230 ;
        RECT 2361.635 1608.235 2361.805 1609.505 ;
        RECT 2373.320 1608.465 2373.490 1609.505 ;
        RECT 2373.315 1608.225 2373.495 1608.465 ;
        RECT 2373.320 1602.955 2373.490 1604.225 ;
        RECT 2366.805 1531.235 2366.975 1532.505 ;
        RECT 2372.420 1531.235 2372.590 1532.505 ;
        RECT 2372.420 1525.955 2372.590 1527.225 ;
        RECT 2369.040 1433.240 2369.210 1434.510 ;
        RECT 2374.655 1433.240 2374.825 1434.510 ;
        RECT 2374.655 1427.955 2374.825 1429.225 ;
        RECT 2375.740 1333.240 2375.910 1334.510 ;
        RECT 2381.355 1333.240 2381.525 1334.510 ;
        RECT 2381.355 1327.955 2381.525 1329.225 ;
      LAYER met1 ;
        RECT 2361.380 2253.400 2361.720 2253.450 ;
        RECT 2361.380 2253.395 2361.725 2253.400 ;
        RECT 2361.380 2253.365 2361.865 2253.395 ;
        RECT 2363.690 2253.365 2364.030 2253.455 ;
        RECT 2361.380 2253.190 2364.030 2253.365 ;
        RECT 2361.380 2253.170 2361.720 2253.190 ;
        RECT 2363.690 2253.175 2364.030 2253.190 ;
        RECT 2372.620 2253.400 2372.945 2253.475 ;
        RECT 2372.620 2253.230 2373.090 2253.400 ;
        RECT 2372.620 2253.150 2372.945 2253.230 ;
        RECT 2372.615 2249.930 2372.940 2250.255 ;
        RECT 2372.690 2249.260 2372.870 2249.930 ;
        RECT 2372.630 2249.230 2372.920 2249.260 ;
        RECT 2372.630 2249.060 2373.090 2249.230 ;
        RECT 2372.630 2249.030 2372.920 2249.060 ;
        RECT 2361.565 2161.400 2361.905 2161.495 ;
        RECT 2361.565 2161.395 2361.920 2161.400 ;
        RECT 2361.565 2161.365 2362.060 2161.395 ;
        RECT 2363.885 2161.365 2364.225 2161.455 ;
        RECT 2361.565 2161.200 2364.225 2161.365 ;
        RECT 2361.565 2161.155 2361.905 2161.200 ;
        RECT 2363.885 2161.175 2364.225 2161.200 ;
        RECT 2373.270 2161.405 2373.595 2161.465 ;
        RECT 2373.270 2161.235 2373.745 2161.405 ;
        RECT 2373.270 2161.140 2373.595 2161.235 ;
        RECT 2373.270 2157.790 2373.595 2158.115 ;
        RECT 2373.350 2157.255 2373.520 2157.790 ;
        RECT 2373.285 2157.225 2373.575 2157.255 ;
        RECT 2373.285 2157.055 2373.745 2157.225 ;
        RECT 2373.285 2157.025 2373.575 2157.055 ;
        RECT 2366.735 2056.405 2367.055 2056.465 ;
        RECT 2366.735 2056.375 2367.210 2056.405 ;
        RECT 2368.610 2056.375 2368.930 2056.420 ;
        RECT 2372.345 2056.405 2372.685 2056.475 ;
        RECT 2372.345 2056.400 2372.825 2056.405 ;
        RECT 2372.330 2056.375 2372.825 2056.400 ;
        RECT 2366.735 2056.235 2372.825 2056.375 ;
        RECT 2366.735 2056.205 2372.685 2056.235 ;
        RECT 2366.735 2056.175 2367.055 2056.205 ;
        RECT 2368.610 2056.160 2368.930 2056.205 ;
        RECT 2372.345 2056.125 2372.685 2056.205 ;
        RECT 2372.355 2052.225 2372.695 2052.370 ;
        RECT 2372.355 2052.055 2372.825 2052.225 ;
        RECT 2372.355 2052.015 2372.695 2052.055 ;
        RECT 2368.960 1951.410 2369.310 1951.500 ;
        RECT 2374.580 1951.410 2374.920 1951.485 ;
        RECT 2368.960 1951.380 2369.445 1951.410 ;
        RECT 2374.580 1951.405 2375.060 1951.410 ;
        RECT 2374.565 1951.380 2375.065 1951.405 ;
        RECT 2368.960 1951.235 2375.065 1951.380 ;
        RECT 2368.960 1951.200 2374.920 1951.235 ;
        RECT 2368.960 1951.150 2369.310 1951.200 ;
        RECT 2374.580 1951.135 2374.920 1951.200 ;
        RECT 2374.590 1947.225 2374.930 1947.350 ;
        RECT 2374.590 1947.055 2375.060 1947.225 ;
        RECT 2374.590 1947.000 2374.930 1947.055 ;
        RECT 2375.600 1788.410 2375.950 1788.470 ;
        RECT 2381.230 1788.410 2381.570 1788.500 ;
        RECT 2375.600 1788.370 2376.090 1788.410 ;
        RECT 2381.230 1788.405 2381.705 1788.410 ;
        RECT 2381.210 1788.370 2381.705 1788.405 ;
        RECT 2375.600 1788.360 2381.705 1788.370 ;
        RECT 2375.510 1788.240 2381.705 1788.360 ;
        RECT 2375.510 1788.205 2381.570 1788.240 ;
        RECT 2375.510 1788.180 2375.950 1788.205 ;
        RECT 2375.510 1788.100 2375.830 1788.180 ;
        RECT 2381.230 1788.150 2381.570 1788.205 ;
        RECT 2381.230 1784.225 2381.570 1784.350 ;
        RECT 2381.230 1784.055 2381.705 1784.225 ;
        RECT 2381.230 1784.000 2381.570 1784.055 ;
        RECT 2361.740 1708.395 2362.080 1708.455 ;
        RECT 2361.740 1708.365 2362.225 1708.395 ;
        RECT 2364.050 1708.365 2364.390 1708.455 ;
        RECT 2361.740 1708.195 2364.390 1708.365 ;
        RECT 2361.740 1708.175 2362.080 1708.195 ;
        RECT 2364.050 1708.175 2364.390 1708.195 ;
        RECT 2372.980 1708.400 2373.305 1708.475 ;
        RECT 2372.980 1708.230 2373.450 1708.400 ;
        RECT 2372.980 1708.150 2373.305 1708.230 ;
        RECT 2372.975 1704.930 2373.300 1705.255 ;
        RECT 2373.050 1704.275 2373.230 1704.930 ;
        RECT 2373.050 1704.260 2373.530 1704.275 ;
        RECT 2372.990 1704.030 2373.530 1704.260 ;
        RECT 2373.210 1704.015 2373.530 1704.030 ;
        RECT 2361.545 1608.405 2361.885 1608.490 ;
        RECT 2361.545 1608.375 2362.035 1608.405 ;
        RECT 2363.860 1608.375 2364.200 1608.455 ;
        RECT 2361.545 1608.200 2364.200 1608.375 ;
        RECT 2361.545 1608.150 2361.885 1608.200 ;
        RECT 2363.860 1608.175 2364.200 1608.200 ;
        RECT 2373.245 1608.405 2373.570 1608.465 ;
        RECT 2373.245 1608.235 2373.720 1608.405 ;
        RECT 2373.245 1608.140 2373.570 1608.235 ;
        RECT 2373.245 1604.790 2373.570 1605.115 ;
        RECT 2373.325 1604.255 2373.495 1604.790 ;
        RECT 2373.260 1604.225 2373.550 1604.255 ;
        RECT 2373.260 1604.055 2373.720 1604.225 ;
        RECT 2373.260 1604.025 2373.550 1604.055 ;
        RECT 2366.720 1531.405 2367.070 1531.465 ;
        RECT 2366.720 1531.375 2367.205 1531.405 ;
        RECT 2368.610 1531.375 2368.930 1531.420 ;
        RECT 2372.340 1531.405 2372.680 1531.475 ;
        RECT 2372.340 1531.400 2372.820 1531.405 ;
        RECT 2372.325 1531.375 2372.820 1531.400 ;
        RECT 2366.720 1531.235 2372.820 1531.375 ;
        RECT 2366.720 1531.205 2372.680 1531.235 ;
        RECT 2366.720 1531.175 2367.070 1531.205 ;
        RECT 2368.610 1531.160 2368.930 1531.205 ;
        RECT 2372.340 1531.125 2372.680 1531.205 ;
        RECT 2372.350 1527.225 2372.690 1527.350 ;
        RECT 2372.350 1527.055 2372.820 1527.225 ;
        RECT 2372.350 1527.000 2372.690 1527.055 ;
        RECT 2368.950 1433.410 2369.300 1433.495 ;
        RECT 2374.575 1433.410 2374.915 1433.485 ;
        RECT 2368.950 1433.380 2369.440 1433.410 ;
        RECT 2374.575 1433.405 2375.055 1433.410 ;
        RECT 2374.560 1433.380 2375.060 1433.405 ;
        RECT 2368.950 1433.235 2375.060 1433.380 ;
        RECT 2368.950 1433.210 2374.915 1433.235 ;
        RECT 2368.950 1433.145 2369.300 1433.210 ;
        RECT 2374.575 1433.135 2374.915 1433.210 ;
        RECT 2374.585 1429.225 2374.925 1429.350 ;
        RECT 2374.585 1429.055 2375.055 1429.225 ;
        RECT 2374.585 1429.000 2374.925 1429.055 ;
        RECT 2375.650 1333.410 2376.000 1333.470 ;
        RECT 2381.280 1333.410 2381.620 1333.500 ;
        RECT 2375.650 1333.380 2376.140 1333.410 ;
        RECT 2381.280 1333.405 2381.755 1333.410 ;
        RECT 2381.260 1333.380 2381.755 1333.405 ;
        RECT 2375.650 1333.240 2381.755 1333.380 ;
        RECT 2375.650 1333.205 2381.620 1333.240 ;
        RECT 2375.650 1333.180 2376.000 1333.205 ;
        RECT 2381.280 1333.150 2381.620 1333.205 ;
        RECT 2381.280 1329.225 2381.620 1329.350 ;
        RECT 2381.280 1329.055 2381.755 1329.225 ;
        RECT 2381.280 1329.000 2381.620 1329.055 ;
      LAYER met2 ;
        RECT 2363.775 2254.315 2372.860 2254.485 ;
        RECT 2361.410 2253.125 2361.690 2253.495 ;
        RECT 2363.775 2253.485 2363.945 2254.315 ;
        RECT 2363.720 2253.145 2364.000 2253.485 ;
        RECT 2372.685 2253.475 2372.860 2254.315 ;
        RECT 2372.620 2253.150 2372.945 2253.475 ;
        RECT 2372.685 2251.890 2372.860 2253.150 ;
        RECT 2370.540 2251.750 2372.860 2251.890 ;
        RECT 2370.540 2248.605 2370.680 2251.750 ;
        RECT 2372.685 2250.255 2372.860 2251.750 ;
        RECT 2372.615 2249.930 2372.940 2250.255 ;
        RECT 2370.470 2248.235 2370.750 2248.605 ;
        RECT 2363.970 2162.320 2373.520 2162.490 ;
        RECT 2361.545 2161.140 2361.920 2161.510 ;
        RECT 2363.970 2161.485 2364.140 2162.320 ;
        RECT 2363.915 2161.145 2364.195 2161.485 ;
        RECT 2373.350 2161.465 2373.520 2162.320 ;
        RECT 2373.270 2161.140 2373.595 2161.465 ;
        RECT 2373.340 2160.090 2373.510 2161.140 ;
        RECT 2371.460 2159.950 2373.510 2160.090 ;
        RECT 2371.460 2159.525 2371.600 2159.950 ;
        RECT 2371.390 2159.155 2371.670 2159.525 ;
        RECT 2373.340 2158.115 2373.510 2159.950 ;
        RECT 2373.270 2157.790 2373.595 2158.115 ;
        RECT 2368.640 2056.130 2368.900 2056.450 ;
        RECT 2368.700 2054.805 2368.840 2056.130 ;
        RECT 2372.345 2056.125 2372.685 2056.475 ;
        RECT 2368.630 2054.435 2368.910 2054.805 ;
        RECT 2372.430 2052.370 2372.600 2056.125 ;
        RECT 2372.355 2052.020 2372.695 2052.370 ;
        RECT 2368.945 1951.135 2369.325 1951.515 ;
        RECT 2374.580 1951.135 2374.920 1951.485 ;
        RECT 2374.665 1947.350 2374.835 1951.135 ;
        RECT 2374.590 1947.000 2374.930 1947.350 ;
        RECT 2374.680 1946.685 2374.820 1947.000 ;
        RECT 2374.610 1946.315 2374.890 1946.685 ;
        RECT 2375.540 1788.070 2375.800 1788.390 ;
        RECT 2381.230 1788.150 2381.570 1788.500 ;
        RECT 2375.070 1787.450 2375.350 1787.565 ;
        RECT 2375.600 1787.450 2375.740 1788.070 ;
        RECT 2375.070 1787.310 2375.740 1787.450 ;
        RECT 2375.070 1787.195 2375.350 1787.310 ;
        RECT 2381.310 1784.350 2381.480 1788.150 ;
        RECT 2381.230 1784.000 2381.570 1784.350 ;
        RECT 2364.135 1709.300 2373.220 1709.470 ;
        RECT 2361.770 1708.130 2362.050 1708.500 ;
        RECT 2364.135 1708.485 2364.305 1709.300 ;
        RECT 2364.080 1708.145 2364.360 1708.485 ;
        RECT 2373.045 1708.475 2373.220 1709.300 ;
        RECT 2372.980 1708.150 2373.305 1708.475 ;
        RECT 2373.045 1705.255 2373.220 1708.150 ;
        RECT 2372.975 1704.930 2373.300 1705.255 ;
        RECT 2373.240 1703.985 2373.500 1704.305 ;
        RECT 2372.770 1702.450 2373.050 1702.565 ;
        RECT 2373.300 1702.450 2373.440 1703.985 ;
        RECT 2372.770 1702.310 2373.440 1702.450 ;
        RECT 2372.770 1702.195 2373.050 1702.310 ;
        RECT 2363.945 1609.240 2373.495 1609.410 ;
        RECT 2361.525 1608.135 2361.900 1608.505 ;
        RECT 2363.945 1608.485 2364.115 1609.240 ;
        RECT 2363.890 1608.145 2364.170 1608.485 ;
        RECT 2373.325 1608.465 2373.495 1609.240 ;
        RECT 2373.245 1608.140 2373.570 1608.465 ;
        RECT 2371.390 1606.570 2371.670 1606.685 ;
        RECT 2373.315 1606.570 2373.485 1608.140 ;
        RECT 2371.390 1606.430 2373.485 1606.570 ;
        RECT 2371.390 1606.315 2371.670 1606.430 ;
        RECT 2373.315 1605.115 2373.485 1606.430 ;
        RECT 2373.245 1604.790 2373.570 1605.115 ;
        RECT 2366.750 1531.130 2367.040 1531.510 ;
        RECT 2368.640 1531.130 2368.900 1531.450 ;
        RECT 2368.700 1529.845 2368.840 1531.130 ;
        RECT 2372.340 1531.125 2372.680 1531.475 ;
        RECT 2368.630 1529.475 2368.910 1529.845 ;
        RECT 2372.425 1527.350 2372.595 1531.125 ;
        RECT 2372.350 1527.000 2372.690 1527.350 ;
        RECT 2374.575 1433.240 2374.915 1433.485 ;
        RECT 2374.560 1432.960 2374.930 1433.240 ;
        RECT 2374.660 1429.350 2374.830 1432.960 ;
        RECT 2374.585 1429.000 2374.925 1429.350 ;
        RECT 2375.680 1333.135 2375.970 1333.515 ;
        RECT 2381.280 1333.150 2381.620 1333.500 ;
        RECT 2381.360 1329.350 2381.530 1333.150 ;
        RECT 2381.280 1329.000 2381.620 1329.350 ;
        RECT 2381.375 1328.450 2381.515 1329.000 ;
        RECT 2381.375 1328.310 2381.720 1328.450 ;
        RECT 2381.580 1325.050 2381.720 1328.310 ;
        RECT 2382.430 1325.050 2382.710 1325.165 ;
        RECT 2381.580 1324.910 2382.710 1325.050 ;
        RECT 2382.430 1324.795 2382.710 1324.910 ;
      LAYER met3 ;
        RECT 2361.380 2253.125 2361.720 2257.455 ;
        RECT 2368.350 2248.570 2368.730 2248.580 ;
        RECT 2370.445 2248.570 2370.775 2248.585 ;
        RECT 2368.350 2248.270 2370.775 2248.570 ;
        RECT 2368.350 2248.260 2368.730 2248.270 ;
        RECT 2370.445 2248.255 2370.775 2248.270 ;
        RECT 2361.570 2161.510 2361.900 2165.445 ;
        RECT 2361.545 2161.140 2361.920 2161.510 ;
        RECT 2368.350 2159.490 2368.730 2159.500 ;
        RECT 2371.365 2159.490 2371.695 2159.505 ;
        RECT 2368.350 2159.190 2371.695 2159.490 ;
        RECT 2368.350 2159.180 2368.730 2159.190 ;
        RECT 2371.365 2159.175 2371.695 2159.190 ;
        RECT 2368.605 2054.780 2368.935 2054.785 ;
        RECT 2368.350 2054.770 2368.935 2054.780 ;
        RECT 2368.350 2054.470 2369.160 2054.770 ;
        RECT 2368.350 2054.460 2368.935 2054.470 ;
        RECT 2368.605 2054.455 2368.935 2054.460 ;
        RECT 2368.350 1960.250 2368.730 1960.260 ;
        RECT 2374.790 1960.250 2375.170 1960.260 ;
        RECT 2368.350 1959.950 2375.170 1960.250 ;
        RECT 2368.350 1959.940 2368.730 1959.950 ;
        RECT 2374.790 1959.940 2375.170 1959.950 ;
        RECT 2368.970 1951.515 2369.295 1955.360 ;
        RECT 2368.945 1951.135 2369.325 1951.515 ;
        RECT 2374.585 1946.660 2374.915 1946.665 ;
        RECT 2374.585 1946.650 2375.170 1946.660 ;
        RECT 2374.360 1946.350 2375.170 1946.650 ;
        RECT 2374.585 1946.340 2375.170 1946.350 ;
        RECT 2374.585 1946.335 2374.915 1946.340 ;
        RECT 2375.045 1787.540 2375.375 1787.545 ;
        RECT 2374.790 1787.530 2375.375 1787.540 ;
        RECT 2374.790 1787.230 2375.600 1787.530 ;
        RECT 2374.790 1787.220 2375.375 1787.230 ;
        RECT 2375.045 1787.215 2375.375 1787.220 ;
        RECT 2368.350 1718.850 2368.730 1718.860 ;
        RECT 2374.790 1718.850 2375.170 1718.860 ;
        RECT 2368.350 1718.550 2375.170 1718.850 ;
        RECT 2368.350 1718.540 2368.730 1718.550 ;
        RECT 2374.790 1718.540 2375.170 1718.550 ;
        RECT 2361.740 1708.130 2362.080 1712.460 ;
        RECT 2368.350 1702.530 2368.730 1702.540 ;
        RECT 2372.745 1702.530 2373.075 1702.545 ;
        RECT 2368.350 1702.230 2373.075 1702.530 ;
        RECT 2368.350 1702.220 2368.730 1702.230 ;
        RECT 2372.745 1702.215 2373.075 1702.230 ;
        RECT 2361.545 1608.505 2361.880 1612.385 ;
        RECT 2361.525 1608.135 2361.900 1608.505 ;
        RECT 2368.350 1606.650 2368.730 1606.660 ;
        RECT 2371.365 1606.650 2371.695 1606.665 ;
        RECT 2368.350 1606.350 2371.695 1606.650 ;
        RECT 2368.350 1606.340 2368.730 1606.350 ;
        RECT 2371.365 1606.335 2371.695 1606.350 ;
        RECT 2366.715 1531.465 2367.065 1535.460 ;
        RECT 2366.720 1531.130 2367.070 1531.465 ;
        RECT 2368.605 1529.820 2368.935 1529.825 ;
        RECT 2368.350 1529.810 2368.935 1529.820 ;
        RECT 2368.350 1529.510 2369.160 1529.810 ;
        RECT 2368.350 1529.500 2368.935 1529.510 ;
        RECT 2368.605 1529.495 2368.935 1529.500 ;
        RECT 2368.350 1448.890 2368.730 1448.900 ;
        RECT 2380.310 1448.890 2380.690 1448.900 ;
        RECT 2368.350 1448.590 2380.690 1448.890 ;
        RECT 2368.350 1448.580 2368.730 1448.590 ;
        RECT 2380.310 1448.580 2380.690 1448.590 ;
        RECT 2374.580 1433.250 2374.910 1433.265 ;
        RECT 2380.310 1433.250 2380.690 1433.260 ;
        RECT 2374.580 1432.950 2380.690 1433.250 ;
        RECT 2374.580 1432.935 2374.910 1432.950 ;
        RECT 2380.310 1432.940 2380.690 1432.950 ;
        RECT 2375.650 1333.135 2376.000 1337.465 ;
        RECT 2382.405 1325.140 2382.735 1325.145 ;
        RECT 2382.150 1325.130 2382.735 1325.140 ;
        RECT 2386.750 1325.130 2387.130 1325.140 ;
        RECT 2381.770 1324.830 2387.130 1325.130 ;
        RECT 2382.150 1324.820 2382.735 1324.830 ;
        RECT 2386.750 1324.820 2387.130 1324.830 ;
        RECT 2382.405 1324.815 2382.735 1324.820 ;
        RECT 2386.750 1028.650 2387.130 1028.660 ;
        RECT 2917.600 1028.650 2924.800 1029.100 ;
        RECT 2386.750 1028.350 2924.800 1028.650 ;
        RECT 2386.750 1028.340 2387.130 1028.350 ;
        RECT 2917.600 1027.900 2924.800 1028.350 ;
      LAYER met4 ;
        RECT 2368.375 2248.255 2368.705 2248.585 ;
        RECT 2368.390 2159.505 2368.690 2248.255 ;
        RECT 2368.375 2159.175 2368.705 2159.505 ;
        RECT 2368.390 2054.785 2368.690 2159.175 ;
        RECT 2368.375 2054.455 2368.705 2054.785 ;
        RECT 2368.390 1960.265 2368.690 2054.455 ;
        RECT 2368.375 1959.935 2368.705 1960.265 ;
        RECT 2374.815 1959.935 2375.145 1960.265 ;
        RECT 2374.830 1946.665 2375.130 1959.935 ;
        RECT 2374.815 1946.335 2375.145 1946.665 ;
        RECT 2374.830 1787.545 2375.130 1946.335 ;
        RECT 2374.815 1787.215 2375.145 1787.545 ;
        RECT 2374.830 1786.850 2375.130 1787.215 ;
        RECT 2374.830 1786.550 2376.970 1786.850 ;
        RECT 2376.670 1783.450 2376.970 1786.550 ;
        RECT 2374.830 1783.150 2376.970 1783.450 ;
        RECT 2374.830 1718.865 2375.130 1783.150 ;
        RECT 2368.375 1718.535 2368.705 1718.865 ;
        RECT 2374.815 1718.535 2375.145 1718.865 ;
        RECT 2368.390 1702.545 2368.690 1718.535 ;
        RECT 2368.375 1702.215 2368.705 1702.545 ;
        RECT 2368.390 1606.665 2368.690 1702.215 ;
        RECT 2368.375 1606.335 2368.705 1606.665 ;
        RECT 2368.390 1529.825 2368.690 1606.335 ;
        RECT 2368.375 1529.495 2368.705 1529.825 ;
        RECT 2368.390 1448.905 2368.690 1529.495 ;
        RECT 2368.375 1448.575 2368.705 1448.905 ;
        RECT 2380.335 1448.575 2380.665 1448.905 ;
        RECT 2380.350 1433.265 2380.650 1448.575 ;
        RECT 2380.335 1432.935 2380.665 1433.265 ;
        RECT 2380.350 1338.750 2380.650 1432.935 ;
        RECT 2380.350 1338.450 2382.490 1338.750 ;
        RECT 2382.190 1325.145 2382.490 1338.450 ;
        RECT 2382.175 1324.815 2382.505 1325.145 ;
        RECT 2386.775 1324.815 2387.105 1325.145 ;
        RECT 2386.790 1028.665 2387.090 1324.815 ;
        RECT 2386.775 1028.335 2387.105 1028.665 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.289999 ;
    PORT
      LAYER li1 ;
        RECT 2378.050 2253.225 2378.220 2254.495 ;
        RECT 2389.275 2253.230 2389.445 2254.500 ;
        RECT 2389.275 2247.960 2389.445 2249.230 ;
        RECT 2378.880 2161.225 2379.050 2162.495 ;
        RECT 2390.565 2161.465 2390.735 2162.505 ;
        RECT 2390.560 2161.225 2390.740 2161.465 ;
        RECT 2390.565 2155.955 2390.735 2157.225 ;
        RECT 2383.135 2056.235 2383.305 2057.505 ;
        RECT 2388.750 2056.235 2388.920 2057.505 ;
        RECT 2388.750 2050.955 2388.920 2052.225 ;
        RECT 2387.605 1951.240 2387.775 1952.510 ;
        RECT 2393.220 1951.240 2393.390 1952.510 ;
        RECT 2393.220 1945.955 2393.390 1947.225 ;
        RECT 2390.950 1788.240 2391.120 1789.510 ;
        RECT 2396.565 1788.240 2396.735 1789.510 ;
        RECT 2396.565 1782.955 2396.735 1784.225 ;
        RECT 2378.410 1708.225 2378.580 1709.495 ;
        RECT 2389.635 1708.230 2389.805 1709.500 ;
        RECT 2389.635 1702.960 2389.805 1704.230 ;
        RECT 2378.855 1608.235 2379.025 1609.505 ;
        RECT 2390.540 1608.465 2390.710 1609.505 ;
        RECT 2390.535 1608.225 2390.715 1608.465 ;
        RECT 2390.540 1602.955 2390.710 1604.225 ;
        RECT 2383.130 1531.235 2383.300 1532.505 ;
        RECT 2388.745 1531.235 2388.915 1532.505 ;
        RECT 2388.745 1525.955 2388.915 1527.225 ;
        RECT 2387.600 1433.240 2387.770 1434.510 ;
        RECT 2393.215 1433.240 2393.385 1434.510 ;
        RECT 2393.215 1427.955 2393.385 1429.225 ;
        RECT 2391.000 1333.240 2391.170 1334.510 ;
        RECT 2396.615 1333.240 2396.785 1334.510 ;
        RECT 2396.615 1327.955 2396.785 1329.225 ;
      LAYER met1 ;
        RECT 2377.965 2253.400 2378.305 2253.450 ;
        RECT 2377.965 2253.395 2378.310 2253.400 ;
        RECT 2377.965 2253.365 2378.450 2253.395 ;
        RECT 2380.275 2253.365 2380.615 2253.455 ;
        RECT 2377.965 2253.190 2380.615 2253.365 ;
        RECT 2377.965 2253.170 2378.305 2253.190 ;
        RECT 2380.275 2253.175 2380.615 2253.190 ;
        RECT 2389.205 2253.400 2389.530 2253.475 ;
        RECT 2389.205 2253.230 2389.675 2253.400 ;
        RECT 2389.205 2253.150 2389.530 2253.230 ;
        RECT 2389.200 2249.930 2389.525 2250.255 ;
        RECT 2389.275 2249.260 2389.455 2249.930 ;
        RECT 2389.215 2249.230 2389.505 2249.260 ;
        RECT 2389.215 2249.060 2389.675 2249.230 ;
        RECT 2389.215 2249.030 2389.505 2249.060 ;
        RECT 2378.785 2161.400 2379.125 2161.495 ;
        RECT 2378.785 2161.395 2379.140 2161.400 ;
        RECT 2378.785 2161.365 2379.280 2161.395 ;
        RECT 2381.105 2161.365 2381.445 2161.455 ;
        RECT 2378.785 2161.200 2381.445 2161.365 ;
        RECT 2378.785 2161.155 2379.125 2161.200 ;
        RECT 2381.105 2161.175 2381.445 2161.200 ;
        RECT 2390.490 2161.405 2390.815 2161.465 ;
        RECT 2390.490 2161.235 2390.965 2161.405 ;
        RECT 2390.490 2161.140 2390.815 2161.235 ;
        RECT 2390.490 2157.790 2390.815 2158.115 ;
        RECT 2390.570 2157.255 2390.740 2157.790 ;
        RECT 2390.505 2157.225 2390.795 2157.255 ;
        RECT 2390.505 2157.055 2390.965 2157.225 ;
        RECT 2390.505 2157.025 2390.795 2157.055 ;
        RECT 2383.035 2056.405 2383.405 2056.505 ;
        RECT 2388.670 2056.405 2389.010 2056.475 ;
        RECT 2383.035 2056.375 2383.535 2056.405 ;
        RECT 2388.670 2056.400 2389.150 2056.405 ;
        RECT 2388.655 2056.375 2389.150 2056.400 ;
        RECT 2383.035 2056.235 2389.150 2056.375 ;
        RECT 2383.035 2056.205 2389.010 2056.235 ;
        RECT 2383.035 2056.135 2383.405 2056.205 ;
        RECT 2388.670 2056.125 2389.010 2056.205 ;
        RECT 2388.680 2052.225 2389.020 2052.370 ;
        RECT 2388.680 2052.200 2392.360 2052.225 ;
        RECT 2388.680 2052.085 2392.390 2052.200 ;
        RECT 2388.680 2052.055 2389.150 2052.085 ;
        RECT 2388.680 2052.015 2389.020 2052.055 ;
        RECT 2392.070 2051.940 2392.390 2052.085 ;
        RECT 2387.520 1951.410 2387.870 1951.500 ;
        RECT 2393.140 1951.410 2393.480 1951.485 ;
        RECT 2387.520 1951.380 2388.005 1951.410 ;
        RECT 2393.140 1951.405 2393.620 1951.410 ;
        RECT 2393.125 1951.380 2393.625 1951.405 ;
        RECT 2387.520 1951.235 2393.625 1951.380 ;
        RECT 2387.520 1951.200 2393.480 1951.235 ;
        RECT 2387.520 1951.150 2387.870 1951.200 ;
        RECT 2393.140 1951.135 2393.480 1951.200 ;
        RECT 2393.150 1947.225 2393.490 1947.350 ;
        RECT 2393.150 1947.055 2393.620 1947.225 ;
        RECT 2393.150 1947.000 2393.490 1947.055 ;
        RECT 2390.860 1788.410 2391.210 1788.470 ;
        RECT 2390.860 1788.370 2391.350 1788.410 ;
        RECT 2394.370 1788.370 2394.690 1788.415 ;
        RECT 2396.490 1788.410 2396.830 1788.500 ;
        RECT 2396.490 1788.405 2396.965 1788.410 ;
        RECT 2396.470 1788.370 2396.965 1788.405 ;
        RECT 2390.860 1788.240 2396.965 1788.370 ;
        RECT 2390.860 1788.205 2396.830 1788.240 ;
        RECT 2390.860 1788.180 2391.210 1788.205 ;
        RECT 2394.370 1788.155 2394.690 1788.205 ;
        RECT 2396.490 1788.150 2396.830 1788.205 ;
        RECT 2396.490 1784.225 2396.830 1784.350 ;
        RECT 2396.490 1784.055 2396.965 1784.225 ;
        RECT 2396.490 1784.000 2396.830 1784.055 ;
        RECT 2378.325 1708.395 2378.665 1708.455 ;
        RECT 2378.325 1708.365 2378.810 1708.395 ;
        RECT 2380.635 1708.365 2380.975 1708.455 ;
        RECT 2378.325 1708.195 2380.975 1708.365 ;
        RECT 2378.325 1708.175 2378.665 1708.195 ;
        RECT 2380.635 1708.175 2380.975 1708.195 ;
        RECT 2389.565 1708.400 2389.890 1708.475 ;
        RECT 2389.565 1708.230 2390.035 1708.400 ;
        RECT 2389.565 1708.150 2389.890 1708.230 ;
        RECT 2389.560 1704.930 2389.885 1705.255 ;
        RECT 2389.635 1704.260 2389.815 1704.930 ;
        RECT 2389.575 1704.230 2389.865 1704.260 ;
        RECT 2389.575 1704.060 2390.035 1704.230 ;
        RECT 2389.575 1704.030 2389.865 1704.060 ;
        RECT 2378.765 1608.405 2379.105 1608.490 ;
        RECT 2378.765 1608.375 2379.255 1608.405 ;
        RECT 2381.080 1608.375 2381.420 1608.455 ;
        RECT 2378.765 1608.200 2381.420 1608.375 ;
        RECT 2378.765 1608.150 2379.105 1608.200 ;
        RECT 2381.080 1608.175 2381.420 1608.200 ;
        RECT 2390.465 1608.405 2390.790 1608.465 ;
        RECT 2390.465 1608.235 2390.940 1608.405 ;
        RECT 2390.465 1608.140 2390.790 1608.235 ;
        RECT 2390.465 1604.790 2390.790 1605.115 ;
        RECT 2390.545 1604.255 2390.715 1604.790 ;
        RECT 2390.480 1604.225 2390.770 1604.255 ;
        RECT 2390.480 1604.055 2390.940 1604.225 ;
        RECT 2390.480 1604.025 2390.770 1604.055 ;
        RECT 2383.045 1531.405 2383.395 1531.465 ;
        RECT 2388.665 1531.405 2389.005 1531.475 ;
        RECT 2383.045 1531.375 2383.530 1531.405 ;
        RECT 2388.665 1531.400 2389.145 1531.405 ;
        RECT 2388.650 1531.375 2389.145 1531.400 ;
        RECT 2383.045 1531.235 2389.145 1531.375 ;
        RECT 2383.045 1531.205 2389.005 1531.235 ;
        RECT 2383.045 1531.175 2383.395 1531.205 ;
        RECT 2388.665 1531.125 2389.005 1531.205 ;
        RECT 2388.675 1527.225 2389.015 1527.350 ;
        RECT 2388.675 1527.055 2389.145 1527.225 ;
        RECT 2388.675 1527.000 2389.015 1527.055 ;
        RECT 2387.510 1433.410 2387.860 1433.495 ;
        RECT 2393.135 1433.410 2393.475 1433.485 ;
        RECT 2387.510 1433.380 2388.000 1433.410 ;
        RECT 2393.135 1433.405 2393.615 1433.410 ;
        RECT 2393.120 1433.380 2393.620 1433.405 ;
        RECT 2387.510 1433.235 2393.620 1433.380 ;
        RECT 2387.510 1433.210 2393.475 1433.235 ;
        RECT 2387.510 1433.145 2387.860 1433.210 ;
        RECT 2393.135 1433.135 2393.475 1433.210 ;
        RECT 2393.145 1429.225 2393.485 1429.350 ;
        RECT 2393.145 1429.055 2393.615 1429.225 ;
        RECT 2393.145 1429.000 2393.485 1429.055 ;
        RECT 2390.910 1333.410 2391.260 1333.470 ;
        RECT 2396.540 1333.410 2396.880 1333.500 ;
        RECT 2390.910 1333.380 2391.400 1333.410 ;
        RECT 2396.540 1333.405 2397.015 1333.410 ;
        RECT 2396.520 1333.380 2397.015 1333.405 ;
        RECT 2390.910 1333.240 2397.015 1333.380 ;
        RECT 2390.910 1333.205 2396.880 1333.240 ;
        RECT 2390.910 1333.180 2391.260 1333.205 ;
        RECT 2396.540 1333.150 2396.880 1333.205 ;
        RECT 2396.540 1329.225 2396.880 1329.350 ;
        RECT 2396.540 1329.055 2397.015 1329.225 ;
        RECT 2396.540 1329.000 2396.880 1329.055 ;
      LAYER met2 ;
        RECT 2380.360 2254.315 2389.445 2254.485 ;
        RECT 2377.995 2253.125 2378.275 2253.495 ;
        RECT 2380.360 2253.485 2380.530 2254.315 ;
        RECT 2380.305 2253.145 2380.585 2253.485 ;
        RECT 2389.270 2253.475 2389.445 2254.315 ;
        RECT 2389.205 2253.150 2389.530 2253.475 ;
        RECT 2389.270 2251.325 2389.445 2253.150 ;
        RECT 2389.215 2250.955 2389.495 2251.325 ;
        RECT 2389.270 2250.255 2389.445 2250.955 ;
        RECT 2389.200 2249.930 2389.525 2250.255 ;
        RECT 2381.190 2162.320 2390.740 2162.490 ;
        RECT 2378.765 2161.140 2379.140 2161.510 ;
        RECT 2381.190 2161.485 2381.360 2162.320 ;
        RECT 2381.135 2161.145 2381.415 2161.485 ;
        RECT 2390.570 2161.465 2390.740 2162.320 ;
        RECT 2390.490 2161.140 2390.815 2161.465 ;
        RECT 2390.560 2158.165 2390.730 2161.140 ;
        RECT 2390.510 2158.115 2390.790 2158.165 ;
        RECT 2390.490 2157.790 2390.815 2158.115 ;
        RECT 2383.035 2056.135 2383.405 2056.505 ;
        RECT 2388.670 2056.125 2389.010 2056.475 ;
        RECT 2388.755 2052.370 2388.925 2056.125 ;
        RECT 2388.680 2052.020 2389.020 2052.370 ;
        RECT 2392.100 2051.910 2392.360 2052.230 ;
        RECT 2392.160 2050.725 2392.300 2051.910 ;
        RECT 2392.090 2050.355 2392.370 2050.725 ;
        RECT 2387.505 1951.135 2387.885 1951.515 ;
        RECT 2393.140 1951.135 2393.480 1951.485 ;
        RECT 2393.225 1947.350 2393.395 1951.135 ;
        RECT 2393.150 1947.000 2393.490 1947.350 ;
        RECT 2393.240 1946.685 2393.380 1947.000 ;
        RECT 2393.170 1946.315 2393.450 1946.685 ;
        RECT 2394.390 1789.915 2394.670 1790.285 ;
        RECT 2394.460 1788.445 2394.600 1789.915 ;
        RECT 2394.400 1788.125 2394.660 1788.445 ;
        RECT 2396.490 1788.150 2396.830 1788.500 ;
        RECT 2396.570 1784.350 2396.740 1788.150 ;
        RECT 2396.490 1784.000 2396.830 1784.350 ;
        RECT 2380.720 1709.300 2389.805 1709.470 ;
        RECT 2378.355 1708.130 2378.635 1708.500 ;
        RECT 2380.720 1708.485 2380.890 1709.300 ;
        RECT 2380.665 1708.145 2380.945 1708.485 ;
        RECT 2389.630 1708.475 2389.805 1709.300 ;
        RECT 2389.565 1708.150 2389.890 1708.475 ;
        RECT 2389.630 1705.255 2389.805 1708.150 ;
        RECT 2389.560 1705.240 2389.885 1705.255 ;
        RECT 2389.530 1704.960 2389.900 1705.240 ;
        RECT 2389.560 1704.930 2389.885 1704.960 ;
        RECT 2381.165 1609.240 2390.715 1609.410 ;
        RECT 2378.745 1608.135 2379.120 1608.505 ;
        RECT 2381.165 1608.485 2381.335 1609.240 ;
        RECT 2381.110 1608.145 2381.390 1608.485 ;
        RECT 2390.545 1608.465 2390.715 1609.240 ;
        RECT 2390.465 1608.140 2390.790 1608.465 ;
        RECT 2390.535 1605.210 2390.705 1608.140 ;
        RECT 2390.535 1605.115 2390.920 1605.210 ;
        RECT 2390.465 1604.790 2390.920 1605.115 ;
        RECT 2390.780 1604.645 2390.920 1604.790 ;
        RECT 2390.710 1604.275 2390.990 1604.645 ;
        RECT 2383.075 1531.130 2383.365 1531.510 ;
        RECT 2388.665 1531.125 2389.005 1531.475 ;
        RECT 2388.750 1528.485 2388.920 1531.125 ;
        RECT 2388.695 1528.115 2388.975 1528.485 ;
        RECT 2388.750 1527.350 2388.920 1528.115 ;
        RECT 2388.675 1527.000 2389.015 1527.350 ;
        RECT 2393.165 1434.275 2393.445 1434.645 ;
        RECT 2393.235 1433.485 2393.375 1434.275 ;
        RECT 2393.135 1433.135 2393.475 1433.485 ;
        RECT 2393.220 1429.350 2393.390 1433.135 ;
        RECT 2393.145 1429.000 2393.485 1429.350 ;
        RECT 2390.940 1333.135 2391.230 1333.515 ;
        RECT 2396.540 1333.150 2396.880 1333.500 ;
        RECT 2395.310 1329.810 2395.590 1329.925 ;
        RECT 2396.620 1329.810 2396.790 1333.150 ;
        RECT 2395.310 1329.670 2396.790 1329.810 ;
        RECT 2395.310 1329.555 2395.590 1329.670 ;
        RECT 2396.620 1329.350 2396.790 1329.670 ;
        RECT 2396.540 1329.000 2396.880 1329.350 ;
        RECT 2396.635 1328.450 2396.775 1329.000 ;
        RECT 2396.635 1328.310 2396.900 1328.450 ;
        RECT 2396.760 1325.050 2396.900 1328.310 ;
        RECT 2397.610 1325.050 2397.890 1325.165 ;
        RECT 2396.760 1324.910 2397.890 1325.050 ;
        RECT 2397.610 1324.795 2397.890 1324.910 ;
      LAYER met3 ;
        RECT 2377.965 2253.125 2378.305 2257.455 ;
        RECT 2389.190 2251.290 2389.520 2251.305 ;
        RECT 2392.270 2251.290 2392.650 2251.300 ;
        RECT 2389.190 2250.990 2392.650 2251.290 ;
        RECT 2389.190 2250.975 2389.520 2250.990 ;
        RECT 2392.270 2250.980 2392.650 2250.990 ;
        RECT 2378.790 2161.510 2379.120 2165.445 ;
        RECT 2378.765 2161.140 2379.140 2161.510 ;
        RECT 2390.485 2158.130 2390.815 2158.145 ;
        RECT 2392.270 2158.130 2392.650 2158.140 ;
        RECT 2390.485 2157.830 2392.650 2158.130 ;
        RECT 2390.485 2157.815 2390.815 2157.830 ;
        RECT 2392.270 2157.820 2392.650 2157.830 ;
        RECT 2392.065 2050.700 2392.395 2050.705 ;
        RECT 2392.065 2050.690 2392.650 2050.700 ;
        RECT 2391.840 2050.390 2392.650 2050.690 ;
        RECT 2392.065 2050.380 2392.650 2050.390 ;
        RECT 2392.065 2050.375 2392.395 2050.380 ;
        RECT 2387.530 1951.515 2387.855 1955.360 ;
        RECT 2387.505 1951.135 2387.885 1951.515 ;
        RECT 2393.145 1946.660 2393.475 1946.665 ;
        RECT 2393.145 1946.650 2393.570 1946.660 ;
        RECT 2392.760 1946.350 2393.570 1946.650 ;
        RECT 2393.145 1946.340 2393.570 1946.350 ;
        RECT 2393.145 1946.335 2393.475 1946.340 ;
        RECT 2393.190 1790.250 2393.570 1790.260 ;
        RECT 2394.365 1790.250 2394.695 1790.265 ;
        RECT 2393.190 1789.950 2394.695 1790.250 ;
        RECT 2393.190 1789.940 2393.570 1789.950 ;
        RECT 2394.365 1789.935 2394.695 1789.950 ;
        RECT 2378.325 1708.130 2378.665 1712.460 ;
        RECT 2389.550 1705.250 2389.880 1705.265 ;
        RECT 2392.270 1705.250 2392.650 1705.260 ;
        RECT 2389.550 1704.950 2392.650 1705.250 ;
        RECT 2389.550 1704.935 2389.880 1704.950 ;
        RECT 2392.270 1704.940 2392.650 1704.950 ;
        RECT 2378.765 1608.505 2379.100 1612.385 ;
        RECT 2378.745 1608.135 2379.120 1608.505 ;
        RECT 2390.685 1604.610 2391.015 1604.625 ;
        RECT 2393.190 1604.610 2393.570 1604.620 ;
        RECT 2390.685 1604.310 2393.570 1604.610 ;
        RECT 2390.685 1604.295 2391.015 1604.310 ;
        RECT 2393.190 1604.300 2393.570 1604.310 ;
        RECT 2383.040 1531.465 2383.390 1535.460 ;
        RECT 2383.045 1531.130 2383.395 1531.465 ;
        RECT 2388.670 1528.450 2389.000 1528.465 ;
        RECT 2394.110 1528.450 2394.490 1528.460 ;
        RECT 2388.670 1528.150 2394.490 1528.450 ;
        RECT 2388.670 1528.135 2389.000 1528.150 ;
        RECT 2394.110 1528.140 2394.490 1528.150 ;
        RECT 2393.140 1434.610 2393.470 1434.625 ;
        RECT 2394.110 1434.610 2394.490 1434.620 ;
        RECT 2393.140 1434.310 2394.490 1434.610 ;
        RECT 2393.140 1434.295 2393.470 1434.310 ;
        RECT 2394.110 1434.300 2394.490 1434.310 ;
        RECT 2390.910 1333.135 2391.260 1337.465 ;
        RECT 2395.285 1329.900 2395.615 1329.905 ;
        RECT 2395.030 1329.890 2395.615 1329.900 ;
        RECT 2394.830 1329.590 2395.615 1329.890 ;
        RECT 2395.030 1329.580 2395.615 1329.590 ;
        RECT 2395.285 1329.575 2395.615 1329.580 ;
        RECT 2397.585 1325.130 2397.915 1325.145 ;
        RECT 2400.550 1325.130 2400.930 1325.140 ;
        RECT 2397.585 1324.830 2400.930 1325.130 ;
        RECT 2397.585 1324.815 2397.915 1324.830 ;
        RECT 2400.550 1324.820 2400.930 1324.830 ;
        RECT 2400.550 1227.890 2400.930 1227.900 ;
        RECT 2917.600 1227.890 2924.800 1228.340 ;
        RECT 2400.550 1227.590 2924.800 1227.890 ;
        RECT 2400.550 1227.580 2400.930 1227.590 ;
        RECT 2917.600 1227.140 2924.800 1227.590 ;
      LAYER met4 ;
        RECT 2392.295 2250.975 2392.625 2251.305 ;
        RECT 2392.310 2158.145 2392.610 2250.975 ;
        RECT 2392.295 2157.815 2392.625 2158.145 ;
        RECT 2392.310 2050.705 2392.610 2157.815 ;
        RECT 2392.295 2050.375 2392.625 2050.705 ;
        RECT 2392.310 2014.950 2392.610 2050.375 ;
        RECT 2392.310 2014.650 2393.530 2014.950 ;
        RECT 2393.230 1946.665 2393.530 2014.650 ;
        RECT 2393.215 1946.335 2393.545 1946.665 ;
        RECT 2393.230 1790.265 2393.530 1946.335 ;
        RECT 2393.215 1789.935 2393.545 1790.265 ;
        RECT 2393.230 1725.150 2393.530 1789.935 ;
        RECT 2392.310 1724.850 2393.530 1725.150 ;
        RECT 2392.310 1705.265 2392.610 1724.850 ;
        RECT 2392.295 1704.935 2392.625 1705.265 ;
        RECT 2392.310 1628.550 2392.610 1704.935 ;
        RECT 2392.310 1628.250 2393.530 1628.550 ;
        RECT 2393.230 1604.625 2393.530 1628.250 ;
        RECT 2393.215 1604.295 2393.545 1604.625 ;
        RECT 2393.230 1531.950 2393.530 1604.295 ;
        RECT 2393.230 1531.650 2394.450 1531.950 ;
        RECT 2394.150 1528.465 2394.450 1531.650 ;
        RECT 2394.135 1528.135 2394.465 1528.465 ;
        RECT 2394.150 1435.350 2394.450 1528.135 ;
        RECT 2394.150 1435.050 2395.370 1435.350 ;
        RECT 2394.150 1434.625 2394.450 1435.050 ;
        RECT 2394.135 1434.295 2394.465 1434.625 ;
        RECT 2395.070 1329.905 2395.370 1435.050 ;
        RECT 2395.055 1329.575 2395.385 1329.905 ;
        RECT 2400.575 1324.815 2400.905 1325.145 ;
        RECT 2400.590 1227.905 2400.890 1324.815 ;
        RECT 2400.575 1227.575 2400.905 1227.905 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.289999 ;
    PORT
      LAYER li1 ;
        RECT 2394.635 2253.225 2394.805 2254.495 ;
        RECT 2405.860 2253.230 2406.030 2254.500 ;
        RECT 2405.860 2247.960 2406.030 2249.230 ;
        RECT 2396.100 2161.225 2396.270 2162.495 ;
        RECT 2407.785 2161.465 2407.955 2162.505 ;
        RECT 2407.780 2161.225 2407.960 2161.465 ;
        RECT 2407.785 2155.955 2407.955 2157.225 ;
        RECT 2399.460 2056.235 2399.630 2057.505 ;
        RECT 2405.075 2056.235 2405.245 2057.505 ;
        RECT 2405.075 2050.955 2405.245 2052.225 ;
        RECT 2406.165 1951.240 2406.335 1952.510 ;
        RECT 2411.780 1951.240 2411.950 1952.510 ;
        RECT 2411.780 1945.955 2411.950 1947.225 ;
        RECT 2406.210 1788.240 2406.380 1789.510 ;
        RECT 2411.825 1788.240 2411.995 1789.510 ;
        RECT 2411.825 1782.955 2411.995 1784.225 ;
        RECT 2394.995 1708.230 2395.165 1709.500 ;
        RECT 2406.220 1708.235 2406.390 1709.505 ;
        RECT 2406.220 1702.965 2406.390 1704.235 ;
        RECT 2396.075 1608.240 2396.245 1609.510 ;
        RECT 2407.760 1608.470 2407.930 1609.510 ;
        RECT 2407.755 1608.230 2407.935 1608.470 ;
        RECT 2407.760 1602.960 2407.930 1604.230 ;
        RECT 2399.455 1531.235 2399.625 1532.505 ;
        RECT 2405.070 1531.235 2405.240 1532.505 ;
        RECT 2405.070 1525.955 2405.240 1527.225 ;
        RECT 2406.160 1433.240 2406.330 1434.510 ;
        RECT 2411.775 1433.240 2411.945 1434.510 ;
        RECT 2411.775 1427.955 2411.945 1429.225 ;
        RECT 2406.260 1333.240 2406.430 1334.510 ;
        RECT 2411.875 1333.240 2412.045 1334.510 ;
        RECT 2411.875 1327.955 2412.045 1329.225 ;
      LAYER met1 ;
        RECT 2394.550 2253.400 2394.890 2253.450 ;
        RECT 2394.550 2253.395 2394.895 2253.400 ;
        RECT 2394.550 2253.365 2395.035 2253.395 ;
        RECT 2396.860 2253.365 2397.200 2253.455 ;
        RECT 2394.550 2253.190 2397.200 2253.365 ;
        RECT 2394.550 2253.170 2394.890 2253.190 ;
        RECT 2396.860 2253.175 2397.200 2253.190 ;
        RECT 2405.790 2253.400 2406.115 2253.475 ;
        RECT 2405.790 2253.230 2406.260 2253.400 ;
        RECT 2405.790 2253.150 2406.115 2253.230 ;
        RECT 2405.785 2249.930 2406.110 2250.255 ;
        RECT 2405.860 2249.260 2406.040 2249.930 ;
        RECT 2405.800 2249.230 2406.090 2249.260 ;
        RECT 2405.800 2249.060 2406.260 2249.230 ;
        RECT 2405.800 2249.030 2406.090 2249.060 ;
        RECT 2396.005 2161.400 2396.345 2161.495 ;
        RECT 2396.005 2161.395 2396.360 2161.400 ;
        RECT 2396.005 2161.365 2396.500 2161.395 ;
        RECT 2398.325 2161.365 2398.665 2161.455 ;
        RECT 2396.005 2161.200 2398.665 2161.365 ;
        RECT 2396.005 2161.155 2396.345 2161.200 ;
        RECT 2398.325 2161.175 2398.665 2161.200 ;
        RECT 2407.710 2161.405 2408.035 2161.465 ;
        RECT 2407.710 2161.235 2408.185 2161.405 ;
        RECT 2407.710 2161.140 2408.035 2161.235 ;
        RECT 2407.710 2157.790 2408.035 2158.115 ;
        RECT 2407.790 2157.255 2407.960 2157.790 ;
        RECT 2407.725 2157.225 2408.015 2157.255 ;
        RECT 2407.725 2157.055 2408.185 2157.225 ;
        RECT 2407.725 2157.025 2408.015 2157.055 ;
        RECT 2399.385 2056.405 2399.705 2056.465 ;
        RECT 2404.995 2056.405 2405.335 2056.475 ;
        RECT 2399.385 2056.375 2399.860 2056.405 ;
        RECT 2404.995 2056.400 2405.475 2056.405 ;
        RECT 2404.980 2056.375 2405.475 2056.400 ;
        RECT 2399.385 2056.235 2405.475 2056.375 ;
        RECT 2399.385 2056.205 2405.335 2056.235 ;
        RECT 2399.385 2056.175 2399.705 2056.205 ;
        RECT 2404.995 2056.125 2405.335 2056.205 ;
        RECT 2405.005 2052.225 2405.345 2052.370 ;
        RECT 2405.005 2052.055 2405.475 2052.225 ;
        RECT 2405.005 2052.015 2405.345 2052.055 ;
        RECT 2406.080 1951.410 2406.430 1951.500 ;
        RECT 2411.700 1951.410 2412.040 1951.485 ;
        RECT 2406.080 1951.380 2406.565 1951.410 ;
        RECT 2411.700 1951.405 2412.180 1951.410 ;
        RECT 2411.685 1951.380 2412.185 1951.405 ;
        RECT 2406.080 1951.235 2412.185 1951.380 ;
        RECT 2406.080 1951.200 2412.040 1951.235 ;
        RECT 2406.080 1951.150 2406.430 1951.200 ;
        RECT 2411.700 1951.135 2412.040 1951.200 ;
        RECT 2411.710 1947.225 2412.050 1947.350 ;
        RECT 2411.710 1947.055 2412.180 1947.225 ;
        RECT 2411.710 1947.000 2412.050 1947.055 ;
        RECT 2406.120 1788.410 2406.470 1788.470 ;
        RECT 2406.120 1788.370 2406.610 1788.410 ;
        RECT 2409.090 1788.370 2409.410 1788.415 ;
        RECT 2411.750 1788.410 2412.090 1788.500 ;
        RECT 2411.750 1788.405 2412.225 1788.410 ;
        RECT 2411.730 1788.370 2412.225 1788.405 ;
        RECT 2406.120 1788.240 2412.225 1788.370 ;
        RECT 2406.120 1788.205 2412.090 1788.240 ;
        RECT 2406.120 1788.180 2406.470 1788.205 ;
        RECT 2409.090 1788.155 2409.410 1788.205 ;
        RECT 2411.750 1788.150 2412.090 1788.205 ;
        RECT 2411.750 1784.225 2412.090 1784.350 ;
        RECT 2411.750 1784.055 2412.225 1784.225 ;
        RECT 2411.750 1784.000 2412.090 1784.055 ;
        RECT 2394.910 1708.400 2395.250 1708.460 ;
        RECT 2394.910 1708.370 2395.395 1708.400 ;
        RECT 2397.220 1708.370 2397.560 1708.460 ;
        RECT 2394.910 1708.200 2397.560 1708.370 ;
        RECT 2394.910 1708.180 2395.250 1708.200 ;
        RECT 2397.220 1708.180 2397.560 1708.200 ;
        RECT 2406.150 1708.405 2406.475 1708.480 ;
        RECT 2406.150 1708.235 2406.620 1708.405 ;
        RECT 2406.150 1708.155 2406.475 1708.235 ;
        RECT 2406.145 1704.935 2406.470 1705.260 ;
        RECT 2406.220 1704.265 2406.400 1704.935 ;
        RECT 2406.160 1704.235 2406.450 1704.265 ;
        RECT 2406.160 1704.065 2406.620 1704.235 ;
        RECT 2406.160 1704.035 2406.450 1704.065 ;
        RECT 2395.985 1608.410 2396.325 1608.495 ;
        RECT 2395.985 1608.380 2396.475 1608.410 ;
        RECT 2398.300 1608.380 2398.640 1608.460 ;
        RECT 2395.985 1608.205 2398.640 1608.380 ;
        RECT 2395.985 1608.155 2396.325 1608.205 ;
        RECT 2398.300 1608.180 2398.640 1608.205 ;
        RECT 2407.685 1608.410 2408.010 1608.470 ;
        RECT 2407.685 1608.240 2408.160 1608.410 ;
        RECT 2407.685 1608.145 2408.010 1608.240 ;
        RECT 2407.685 1604.795 2408.010 1605.120 ;
        RECT 2407.765 1604.260 2407.935 1604.795 ;
        RECT 2407.700 1604.230 2407.990 1604.260 ;
        RECT 2407.700 1604.060 2408.160 1604.230 ;
        RECT 2407.700 1604.030 2407.990 1604.060 ;
        RECT 2399.370 1531.405 2399.720 1531.465 ;
        RECT 2404.990 1531.405 2405.330 1531.475 ;
        RECT 2399.370 1531.375 2399.855 1531.405 ;
        RECT 2404.990 1531.400 2405.470 1531.405 ;
        RECT 2404.975 1531.375 2405.470 1531.400 ;
        RECT 2399.370 1531.235 2405.470 1531.375 ;
        RECT 2399.370 1531.205 2405.330 1531.235 ;
        RECT 2399.370 1531.175 2399.720 1531.205 ;
        RECT 2404.990 1531.125 2405.330 1531.205 ;
        RECT 2405.000 1527.225 2405.340 1527.350 ;
        RECT 2405.000 1527.055 2405.470 1527.225 ;
        RECT 2405.000 1527.000 2405.340 1527.055 ;
        RECT 2406.070 1433.410 2406.420 1433.495 ;
        RECT 2411.695 1433.410 2412.035 1433.485 ;
        RECT 2406.070 1433.380 2406.560 1433.410 ;
        RECT 2411.695 1433.405 2412.175 1433.410 ;
        RECT 2411.680 1433.380 2412.180 1433.405 ;
        RECT 2406.070 1433.235 2412.180 1433.380 ;
        RECT 2406.070 1433.210 2412.035 1433.235 ;
        RECT 2406.070 1433.145 2406.420 1433.210 ;
        RECT 2411.695 1433.135 2412.035 1433.210 ;
        RECT 2411.705 1429.225 2412.045 1429.350 ;
        RECT 2411.705 1429.055 2412.175 1429.225 ;
        RECT 2411.705 1429.000 2412.045 1429.055 ;
        RECT 2406.170 1333.410 2406.520 1333.470 ;
        RECT 2411.800 1333.410 2412.140 1333.500 ;
        RECT 2406.170 1333.380 2406.660 1333.410 ;
        RECT 2411.800 1333.405 2412.275 1333.410 ;
        RECT 2411.780 1333.380 2412.275 1333.405 ;
        RECT 2406.170 1333.240 2412.275 1333.380 ;
        RECT 2406.170 1333.205 2412.140 1333.240 ;
        RECT 2406.170 1333.180 2406.520 1333.205 ;
        RECT 2411.800 1333.150 2412.140 1333.205 ;
        RECT 2411.800 1329.225 2412.140 1329.350 ;
        RECT 2411.800 1329.055 2412.275 1329.225 ;
        RECT 2411.800 1329.000 2412.140 1329.055 ;
      LAYER met2 ;
        RECT 2396.945 2254.315 2406.030 2254.485 ;
        RECT 2394.580 2253.125 2394.860 2253.495 ;
        RECT 2396.945 2253.485 2397.115 2254.315 ;
        RECT 2396.890 2253.145 2397.170 2253.485 ;
        RECT 2405.855 2253.475 2406.030 2254.315 ;
        RECT 2405.790 2253.150 2406.115 2253.475 ;
        RECT 2405.855 2251.325 2406.030 2253.150 ;
        RECT 2405.800 2250.955 2406.080 2251.325 ;
        RECT 2405.855 2250.255 2406.030 2250.955 ;
        RECT 2405.785 2249.930 2406.110 2250.255 ;
        RECT 2398.410 2162.320 2407.960 2162.490 ;
        RECT 2395.985 2161.140 2396.360 2161.510 ;
        RECT 2398.410 2161.485 2398.580 2162.320 ;
        RECT 2398.355 2161.145 2398.635 2161.485 ;
        RECT 2407.790 2161.465 2407.960 2162.320 ;
        RECT 2407.710 2161.140 2408.035 2161.465 ;
        RECT 2406.350 2160.770 2406.630 2160.885 ;
        RECT 2407.780 2160.770 2407.950 2161.140 ;
        RECT 2406.350 2160.630 2407.950 2160.770 ;
        RECT 2406.350 2160.515 2406.630 2160.630 ;
        RECT 2407.780 2158.115 2407.950 2160.630 ;
        RECT 2407.710 2157.790 2408.035 2158.115 ;
        RECT 2404.995 2056.125 2405.335 2056.475 ;
        RECT 2405.080 2052.370 2405.250 2056.125 ;
        RECT 2405.005 2052.020 2405.345 2052.370 ;
        RECT 2405.095 2051.290 2405.235 2052.020 ;
        RECT 2405.095 2051.150 2405.640 2051.290 ;
        RECT 2405.500 2050.610 2405.640 2051.150 ;
        RECT 2406.810 2050.610 2407.090 2050.725 ;
        RECT 2405.500 2050.470 2407.090 2050.610 ;
        RECT 2406.810 2050.355 2407.090 2050.470 ;
        RECT 2406.065 1951.135 2406.445 1951.515 ;
        RECT 2411.700 1951.135 2412.040 1951.485 ;
        RECT 2410.490 1947.250 2410.770 1947.365 ;
        RECT 2411.785 1947.350 2411.955 1951.135 ;
        RECT 2411.710 1947.250 2412.050 1947.350 ;
        RECT 2410.490 1947.110 2412.050 1947.250 ;
        RECT 2410.490 1946.995 2410.770 1947.110 ;
        RECT 2411.710 1947.000 2412.050 1947.110 ;
        RECT 2409.110 1789.915 2409.390 1790.285 ;
        RECT 2409.180 1788.445 2409.320 1789.915 ;
        RECT 2409.120 1788.125 2409.380 1788.445 ;
        RECT 2411.750 1788.150 2412.090 1788.500 ;
        RECT 2411.830 1784.350 2412.000 1788.150 ;
        RECT 2411.750 1784.000 2412.090 1784.350 ;
        RECT 2397.305 1709.305 2406.390 1709.475 ;
        RECT 2394.940 1708.135 2395.220 1708.505 ;
        RECT 2397.305 1708.490 2397.475 1709.305 ;
        RECT 2397.250 1708.150 2397.530 1708.490 ;
        RECT 2406.215 1708.480 2406.390 1709.305 ;
        RECT 2406.150 1708.155 2406.475 1708.480 ;
        RECT 2406.215 1705.260 2406.390 1708.155 ;
        RECT 2406.145 1705.240 2406.470 1705.260 ;
        RECT 2406.115 1704.960 2406.485 1705.240 ;
        RECT 2406.145 1704.935 2406.470 1704.960 ;
        RECT 2398.385 1609.245 2407.935 1609.415 ;
        RECT 2395.965 1608.140 2396.340 1608.510 ;
        RECT 2398.385 1608.490 2398.555 1609.245 ;
        RECT 2398.330 1608.150 2398.610 1608.490 ;
        RECT 2407.765 1608.470 2407.935 1609.245 ;
        RECT 2407.685 1608.145 2408.010 1608.470 ;
        RECT 2405.890 1605.210 2406.170 1605.325 ;
        RECT 2407.755 1605.210 2407.925 1608.145 ;
        RECT 2405.890 1605.120 2407.925 1605.210 ;
        RECT 2405.890 1605.070 2408.010 1605.120 ;
        RECT 2405.890 1604.955 2406.170 1605.070 ;
        RECT 2407.685 1604.795 2408.010 1605.070 ;
        RECT 2404.510 1532.195 2404.790 1532.565 ;
        RECT 2399.400 1531.130 2399.690 1531.510 ;
        RECT 2404.580 1530.410 2404.720 1532.195 ;
        RECT 2404.990 1531.125 2405.330 1531.475 ;
        RECT 2405.075 1530.410 2405.245 1531.125 ;
        RECT 2404.580 1530.270 2405.245 1530.410 ;
        RECT 2405.075 1527.350 2405.245 1530.270 ;
        RECT 2405.000 1527.000 2405.340 1527.350 ;
        RECT 2411.410 1511.115 2411.690 1511.485 ;
        RECT 2900.850 1511.115 2901.130 1511.485 ;
        RECT 2411.480 1442.125 2411.620 1511.115 ;
        RECT 2900.920 1493.805 2901.060 1511.115 ;
        RECT 2900.850 1493.435 2901.130 1493.805 ;
        RECT 2411.410 1441.755 2411.690 1442.125 ;
        RECT 2411.695 1433.135 2412.035 1433.485 ;
        RECT 2411.780 1429.350 2411.950 1433.135 ;
        RECT 2411.705 1429.090 2412.045 1429.350 ;
        RECT 2411.020 1429.000 2412.045 1429.090 ;
        RECT 2411.020 1428.950 2411.865 1429.000 ;
        RECT 2411.020 1428.525 2411.160 1428.950 ;
        RECT 2410.950 1428.155 2411.230 1428.525 ;
        RECT 2411.870 1366.275 2412.150 1366.645 ;
        RECT 2411.940 1336.725 2412.080 1366.275 ;
        RECT 2411.870 1336.355 2412.150 1336.725 ;
        RECT 2411.870 1334.995 2412.150 1335.365 ;
        RECT 2411.940 1333.890 2412.080 1334.995 ;
        RECT 2411.895 1333.750 2412.080 1333.890 ;
        RECT 2406.200 1333.135 2406.490 1333.515 ;
        RECT 2411.895 1333.500 2412.035 1333.750 ;
        RECT 2411.800 1333.150 2412.140 1333.500 ;
        RECT 2411.880 1329.350 2412.050 1333.150 ;
        RECT 2411.800 1329.000 2412.140 1329.350 ;
      LAYER met3 ;
        RECT 2394.550 2253.125 2394.890 2257.455 ;
        RECT 2405.775 2251.300 2406.105 2251.305 ;
        RECT 2405.775 2251.290 2406.450 2251.300 ;
        RECT 2405.775 2250.990 2406.560 2251.290 ;
        RECT 2405.775 2250.980 2406.450 2250.990 ;
        RECT 2405.775 2250.975 2406.105 2250.980 ;
        RECT 2396.010 2161.510 2396.340 2165.445 ;
        RECT 2395.985 2161.140 2396.360 2161.510 ;
        RECT 2406.325 2160.860 2406.655 2160.865 ;
        RECT 2406.070 2160.850 2406.655 2160.860 ;
        RECT 2406.070 2160.550 2406.880 2160.850 ;
        RECT 2406.070 2160.540 2406.655 2160.550 ;
        RECT 2406.325 2160.535 2406.655 2160.540 ;
        RECT 2406.785 2050.700 2407.115 2050.705 ;
        RECT 2406.785 2050.690 2407.370 2050.700 ;
        RECT 2406.560 2050.390 2407.370 2050.690 ;
        RECT 2406.785 2050.380 2407.370 2050.390 ;
        RECT 2406.785 2050.375 2407.115 2050.380 ;
        RECT 2406.090 1951.515 2406.415 1955.360 ;
        RECT 2406.065 1951.135 2406.445 1951.515 ;
        RECT 2408.830 1947.330 2409.210 1947.340 ;
        RECT 2410.465 1947.330 2410.795 1947.345 ;
        RECT 2408.830 1947.030 2410.795 1947.330 ;
        RECT 2408.830 1947.020 2409.210 1947.030 ;
        RECT 2410.465 1947.015 2410.795 1947.030 ;
        RECT 2409.085 1790.260 2409.415 1790.265 ;
        RECT 2408.830 1790.250 2409.415 1790.260 ;
        RECT 2408.830 1789.950 2409.640 1790.250 ;
        RECT 2408.830 1789.940 2409.415 1789.950 ;
        RECT 2409.085 1789.935 2409.415 1789.940 ;
        RECT 2394.910 1708.135 2395.250 1712.465 ;
        RECT 2406.135 1705.250 2406.465 1705.265 ;
        RECT 2406.990 1705.250 2407.370 1705.260 ;
        RECT 2406.135 1704.950 2407.370 1705.250 ;
        RECT 2406.135 1704.935 2406.465 1704.950 ;
        RECT 2406.990 1704.940 2407.370 1704.950 ;
        RECT 2395.985 1608.510 2396.320 1612.390 ;
        RECT 2395.965 1608.140 2396.340 1608.510 ;
        RECT 2405.150 1605.290 2405.530 1605.300 ;
        RECT 2405.865 1605.290 2406.195 1605.305 ;
        RECT 2405.150 1604.990 2406.195 1605.290 ;
        RECT 2405.150 1604.980 2405.530 1604.990 ;
        RECT 2405.865 1604.975 2406.195 1604.990 ;
        RECT 2399.365 1531.465 2399.715 1535.460 ;
        RECT 2404.485 1532.540 2404.815 1532.545 ;
        RECT 2404.230 1532.530 2404.815 1532.540 ;
        RECT 2404.230 1532.230 2405.040 1532.530 ;
        RECT 2404.230 1532.220 2404.815 1532.230 ;
        RECT 2404.485 1532.215 2404.815 1532.220 ;
        RECT 2399.370 1531.130 2399.720 1531.465 ;
        RECT 2404.230 1511.450 2404.610 1511.460 ;
        RECT 2411.385 1511.450 2411.715 1511.465 ;
        RECT 2900.825 1511.450 2901.155 1511.465 ;
        RECT 2404.230 1511.150 2901.155 1511.450 ;
        RECT 2404.230 1511.140 2404.610 1511.150 ;
        RECT 2411.385 1511.135 2411.715 1511.150 ;
        RECT 2900.825 1511.135 2901.155 1511.150 ;
        RECT 2900.825 1493.770 2901.155 1493.785 ;
        RECT 2917.600 1493.770 2924.800 1494.220 ;
        RECT 2900.825 1493.470 2924.800 1493.770 ;
        RECT 2900.825 1493.455 2901.155 1493.470 ;
        RECT 2917.600 1493.020 2924.800 1493.470 ;
        RECT 2410.670 1442.090 2411.050 1442.100 ;
        RECT 2411.385 1442.090 2411.715 1442.105 ;
        RECT 2410.670 1441.790 2411.715 1442.090 ;
        RECT 2410.670 1441.780 2411.050 1441.790 ;
        RECT 2411.385 1441.775 2411.715 1441.790 ;
        RECT 2410.925 1428.500 2411.255 1428.505 ;
        RECT 2410.670 1428.490 2411.255 1428.500 ;
        RECT 2410.670 1428.190 2411.480 1428.490 ;
        RECT 2410.670 1428.180 2411.255 1428.190 ;
        RECT 2410.925 1428.175 2411.255 1428.180 ;
        RECT 2410.670 1366.610 2411.050 1366.620 ;
        RECT 2411.845 1366.610 2412.175 1366.625 ;
        RECT 2410.670 1366.310 2412.175 1366.610 ;
        RECT 2410.670 1366.300 2411.050 1366.310 ;
        RECT 2411.845 1366.295 2412.175 1366.310 ;
        RECT 2406.170 1333.135 2406.520 1337.465 ;
        RECT 2411.845 1336.690 2412.175 1336.705 ;
        RECT 2411.630 1336.375 2412.175 1336.690 ;
        RECT 2411.630 1335.345 2411.930 1336.375 ;
        RECT 2411.630 1335.030 2412.175 1335.345 ;
        RECT 2411.845 1335.015 2412.175 1335.030 ;
      LAYER met4 ;
        RECT 2406.095 2250.975 2406.425 2251.305 ;
        RECT 2406.110 2160.865 2406.410 2250.975 ;
        RECT 2406.095 2160.535 2406.425 2160.865 ;
        RECT 2406.110 2159.850 2406.410 2160.535 ;
        RECT 2405.190 2159.550 2406.410 2159.850 ;
        RECT 2405.190 2111.550 2405.490 2159.550 ;
        RECT 2405.190 2111.250 2407.330 2111.550 ;
        RECT 2407.030 2050.705 2407.330 2111.250 ;
        RECT 2407.015 2050.375 2407.345 2050.705 ;
        RECT 2407.030 1966.650 2407.330 2050.375 ;
        RECT 2407.030 1966.350 2409.170 1966.650 ;
        RECT 2408.870 1947.345 2409.170 1966.350 ;
        RECT 2408.855 1947.015 2409.185 1947.345 ;
        RECT 2408.870 1790.265 2409.170 1947.015 ;
        RECT 2408.855 1789.935 2409.185 1790.265 ;
        RECT 2408.870 1773.450 2409.170 1789.935 ;
        RECT 2407.950 1773.150 2409.170 1773.450 ;
        RECT 2407.950 1725.150 2408.250 1773.150 ;
        RECT 2407.030 1724.850 2408.250 1725.150 ;
        RECT 2407.030 1705.265 2407.330 1724.850 ;
        RECT 2407.015 1704.935 2407.345 1705.265 ;
        RECT 2407.030 1628.550 2407.330 1704.935 ;
        RECT 2405.190 1628.250 2407.330 1628.550 ;
        RECT 2405.190 1605.305 2405.490 1628.250 ;
        RECT 2405.175 1604.975 2405.505 1605.305 ;
        RECT 2405.190 1580.250 2405.490 1604.975 ;
        RECT 2404.270 1579.950 2405.490 1580.250 ;
        RECT 2404.270 1532.545 2404.570 1579.950 ;
        RECT 2404.255 1532.215 2404.585 1532.545 ;
        RECT 2404.270 1511.465 2404.570 1532.215 ;
        RECT 2404.255 1511.135 2404.585 1511.465 ;
        RECT 2410.695 1441.775 2411.025 1442.105 ;
        RECT 2410.710 1428.505 2411.010 1441.775 ;
        RECT 2410.695 1428.175 2411.025 1428.505 ;
        RECT 2410.710 1366.625 2411.010 1428.175 ;
        RECT 2410.695 1366.295 2411.025 1366.625 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.289999 ;
    PORT
      LAYER li1 ;
        RECT 2411.220 2253.225 2411.390 2254.495 ;
        RECT 2422.445 2253.230 2422.615 2254.500 ;
        RECT 2422.445 2247.960 2422.615 2249.230 ;
        RECT 2413.320 2161.225 2413.490 2162.495 ;
        RECT 2425.005 2161.465 2425.175 2162.505 ;
        RECT 2425.000 2161.225 2425.180 2161.465 ;
        RECT 2425.005 2155.955 2425.175 2157.225 ;
        RECT 2415.785 2056.235 2415.955 2057.505 ;
        RECT 2421.400 2056.235 2421.570 2057.505 ;
        RECT 2421.400 2050.955 2421.570 2052.225 ;
        RECT 2424.725 1951.240 2424.895 1952.510 ;
        RECT 2430.340 1951.240 2430.510 1952.510 ;
        RECT 2430.340 1945.955 2430.510 1947.225 ;
        RECT 2421.470 1788.240 2421.640 1789.510 ;
        RECT 2427.085 1788.240 2427.255 1789.510 ;
        RECT 2427.085 1782.955 2427.255 1784.225 ;
        RECT 2411.580 1708.235 2411.750 1709.505 ;
        RECT 2422.805 1708.240 2422.975 1709.510 ;
        RECT 2422.805 1702.970 2422.975 1704.240 ;
        RECT 2413.295 1608.235 2413.465 1609.505 ;
        RECT 2424.980 1608.465 2425.150 1609.505 ;
        RECT 2424.975 1608.225 2425.155 1608.465 ;
        RECT 2424.980 1602.955 2425.150 1604.225 ;
        RECT 2415.780 1531.235 2415.950 1532.505 ;
        RECT 2421.395 1531.235 2421.565 1532.505 ;
        RECT 2421.395 1525.955 2421.565 1527.225 ;
        RECT 2424.720 1433.240 2424.890 1434.510 ;
        RECT 2430.335 1433.240 2430.505 1434.510 ;
        RECT 2430.335 1427.955 2430.505 1429.225 ;
        RECT 2421.520 1333.240 2421.690 1334.510 ;
        RECT 2427.135 1333.240 2427.305 1334.510 ;
        RECT 2427.135 1327.955 2427.305 1329.225 ;
      LAYER met1 ;
        RECT 2411.135 2253.400 2411.475 2253.450 ;
        RECT 2411.135 2253.395 2411.480 2253.400 ;
        RECT 2411.135 2253.365 2411.620 2253.395 ;
        RECT 2413.445 2253.365 2413.785 2253.455 ;
        RECT 2411.135 2253.190 2413.785 2253.365 ;
        RECT 2411.135 2253.170 2411.475 2253.190 ;
        RECT 2413.445 2253.175 2413.785 2253.190 ;
        RECT 2422.375 2253.400 2422.700 2253.475 ;
        RECT 2422.375 2253.230 2422.845 2253.400 ;
        RECT 2422.375 2253.150 2422.700 2253.230 ;
        RECT 2422.370 2249.930 2422.695 2250.255 ;
        RECT 2422.445 2249.260 2422.625 2249.930 ;
        RECT 2422.385 2249.230 2422.675 2249.260 ;
        RECT 2422.385 2249.060 2422.845 2249.230 ;
        RECT 2422.385 2249.030 2422.675 2249.060 ;
        RECT 2413.225 2161.400 2413.565 2161.495 ;
        RECT 2413.225 2161.395 2413.580 2161.400 ;
        RECT 2413.225 2161.365 2413.720 2161.395 ;
        RECT 2415.545 2161.365 2415.885 2161.455 ;
        RECT 2413.225 2161.200 2415.885 2161.365 ;
        RECT 2413.225 2161.155 2413.565 2161.200 ;
        RECT 2415.545 2161.175 2415.885 2161.200 ;
        RECT 2424.930 2161.405 2425.255 2161.465 ;
        RECT 2424.930 2161.235 2425.405 2161.405 ;
        RECT 2424.930 2161.140 2425.255 2161.235 ;
        RECT 2424.930 2157.790 2425.255 2158.115 ;
        RECT 2425.010 2157.255 2425.180 2157.790 ;
        RECT 2424.945 2157.225 2425.235 2157.255 ;
        RECT 2424.945 2157.055 2425.405 2157.225 ;
        RECT 2424.945 2157.025 2425.235 2157.055 ;
        RECT 2415.710 2056.405 2416.030 2056.465 ;
        RECT 2421.320 2056.405 2421.660 2056.475 ;
        RECT 2415.710 2056.375 2416.185 2056.405 ;
        RECT 2421.320 2056.400 2421.800 2056.405 ;
        RECT 2421.305 2056.375 2421.800 2056.400 ;
        RECT 2415.710 2056.235 2421.800 2056.375 ;
        RECT 2415.710 2056.205 2421.660 2056.235 ;
        RECT 2415.710 2056.175 2416.030 2056.205 ;
        RECT 2421.320 2056.125 2421.660 2056.205 ;
        RECT 2421.330 2052.225 2421.670 2052.370 ;
        RECT 2421.330 2052.055 2421.800 2052.225 ;
        RECT 2421.330 2052.015 2421.670 2052.055 ;
        RECT 2424.640 1951.410 2424.990 1951.500 ;
        RECT 2430.260 1951.410 2430.600 1951.485 ;
        RECT 2424.640 1951.380 2425.125 1951.410 ;
        RECT 2430.260 1951.405 2430.740 1951.410 ;
        RECT 2430.245 1951.380 2430.745 1951.405 ;
        RECT 2424.640 1951.235 2430.745 1951.380 ;
        RECT 2424.640 1951.200 2430.600 1951.235 ;
        RECT 2424.640 1951.150 2424.990 1951.200 ;
        RECT 2430.260 1951.135 2430.600 1951.200 ;
        RECT 2430.270 1947.225 2430.610 1947.350 ;
        RECT 2430.270 1947.055 2430.740 1947.225 ;
        RECT 2430.270 1947.000 2430.610 1947.055 ;
        RECT 2421.380 1788.410 2421.730 1788.470 ;
        RECT 2421.380 1788.370 2421.870 1788.410 ;
        RECT 2424.730 1788.370 2425.050 1788.415 ;
        RECT 2427.010 1788.410 2427.350 1788.500 ;
        RECT 2427.010 1788.405 2427.485 1788.410 ;
        RECT 2426.990 1788.370 2427.485 1788.405 ;
        RECT 2421.380 1788.240 2427.485 1788.370 ;
        RECT 2421.380 1788.205 2427.350 1788.240 ;
        RECT 2421.380 1788.180 2421.730 1788.205 ;
        RECT 2424.730 1788.155 2425.050 1788.205 ;
        RECT 2427.010 1788.150 2427.350 1788.205 ;
        RECT 2427.010 1784.225 2427.350 1784.350 ;
        RECT 2427.010 1784.055 2427.485 1784.225 ;
        RECT 2427.010 1784.000 2427.350 1784.055 ;
        RECT 2411.495 1708.405 2411.835 1708.465 ;
        RECT 2411.495 1708.375 2411.980 1708.405 ;
        RECT 2413.805 1708.375 2414.145 1708.465 ;
        RECT 2411.495 1708.205 2414.145 1708.375 ;
        RECT 2411.495 1708.185 2411.835 1708.205 ;
        RECT 2413.805 1708.185 2414.145 1708.205 ;
        RECT 2422.735 1708.410 2423.060 1708.485 ;
        RECT 2422.735 1708.240 2423.205 1708.410 ;
        RECT 2422.735 1708.160 2423.060 1708.240 ;
        RECT 2421.970 1704.980 2422.290 1705.240 ;
        RECT 2422.730 1704.940 2423.055 1705.265 ;
        RECT 2422.805 1704.270 2422.985 1704.940 ;
        RECT 2422.745 1704.240 2423.035 1704.270 ;
        RECT 2422.745 1704.070 2423.205 1704.240 ;
        RECT 2422.745 1704.040 2423.035 1704.070 ;
        RECT 2413.205 1608.405 2413.545 1608.490 ;
        RECT 2413.205 1608.375 2413.695 1608.405 ;
        RECT 2415.520 1608.375 2415.860 1608.455 ;
        RECT 2413.205 1608.200 2415.860 1608.375 ;
        RECT 2413.205 1608.150 2413.545 1608.200 ;
        RECT 2415.520 1608.175 2415.860 1608.200 ;
        RECT 2424.905 1608.405 2425.230 1608.465 ;
        RECT 2424.905 1608.235 2425.380 1608.405 ;
        RECT 2424.905 1608.140 2425.230 1608.235 ;
        RECT 2424.905 1604.790 2425.230 1605.115 ;
        RECT 2424.985 1604.255 2425.155 1604.790 ;
        RECT 2424.920 1604.225 2425.210 1604.255 ;
        RECT 2424.920 1604.055 2425.380 1604.225 ;
        RECT 2424.920 1604.025 2425.210 1604.055 ;
        RECT 2415.695 1531.405 2416.045 1531.465 ;
        RECT 2421.315 1531.405 2421.655 1531.475 ;
        RECT 2415.695 1531.375 2416.180 1531.405 ;
        RECT 2421.315 1531.400 2421.795 1531.405 ;
        RECT 2421.300 1531.375 2421.795 1531.400 ;
        RECT 2415.695 1531.235 2421.795 1531.375 ;
        RECT 2415.695 1531.205 2421.655 1531.235 ;
        RECT 2415.695 1531.175 2416.045 1531.205 ;
        RECT 2421.315 1531.125 2421.655 1531.205 ;
        RECT 2421.325 1527.225 2421.665 1527.350 ;
        RECT 2421.325 1527.055 2421.795 1527.225 ;
        RECT 2421.325 1527.000 2421.665 1527.055 ;
        RECT 2424.630 1433.410 2424.980 1433.495 ;
        RECT 2430.255 1433.410 2430.595 1433.485 ;
        RECT 2424.630 1433.380 2425.120 1433.410 ;
        RECT 2430.255 1433.405 2430.735 1433.410 ;
        RECT 2430.240 1433.380 2430.740 1433.405 ;
        RECT 2424.630 1433.235 2430.740 1433.380 ;
        RECT 2424.630 1433.210 2430.595 1433.235 ;
        RECT 2424.630 1433.145 2425.050 1433.210 ;
        RECT 2424.730 1433.140 2425.050 1433.145 ;
        RECT 2430.255 1433.135 2430.595 1433.210 ;
        RECT 2430.265 1429.225 2430.605 1429.350 ;
        RECT 2430.265 1429.055 2430.735 1429.225 ;
        RECT 2430.265 1429.000 2430.605 1429.055 ;
        RECT 2421.430 1333.410 2421.780 1333.470 ;
        RECT 2427.060 1333.410 2427.400 1333.500 ;
        RECT 2421.430 1333.380 2421.920 1333.410 ;
        RECT 2427.060 1333.405 2427.535 1333.410 ;
        RECT 2427.040 1333.380 2427.535 1333.405 ;
        RECT 2421.430 1333.240 2427.535 1333.380 ;
        RECT 2421.430 1333.205 2427.400 1333.240 ;
        RECT 2421.430 1333.180 2421.780 1333.205 ;
        RECT 2427.060 1333.150 2427.400 1333.205 ;
        RECT 2427.060 1329.225 2427.400 1329.350 ;
        RECT 2427.060 1329.055 2427.535 1329.225 ;
        RECT 2427.060 1329.000 2427.400 1329.055 ;
      LAYER met2 ;
        RECT 2413.530 2254.315 2422.615 2254.485 ;
        RECT 2411.165 2253.125 2411.445 2253.495 ;
        RECT 2413.530 2253.485 2413.700 2254.315 ;
        RECT 2413.475 2253.145 2413.755 2253.485 ;
        RECT 2422.440 2253.475 2422.615 2254.315 ;
        RECT 2422.375 2253.150 2422.700 2253.475 ;
        RECT 2422.440 2250.255 2422.615 2253.150 ;
        RECT 2422.370 2249.930 2422.695 2250.255 ;
        RECT 2422.555 2247.650 2422.695 2249.930 ;
        RECT 2418.380 2247.510 2422.695 2247.650 ;
        RECT 2418.380 2164.285 2418.520 2247.510 ;
        RECT 2418.310 2163.915 2418.590 2164.285 ;
        RECT 2415.630 2162.320 2425.180 2162.490 ;
        RECT 2413.205 2161.140 2413.580 2161.510 ;
        RECT 2415.630 2161.485 2415.800 2162.320 ;
        RECT 2415.575 2161.450 2415.855 2161.485 ;
        RECT 2417.850 2161.450 2418.130 2161.565 ;
        RECT 2425.010 2161.465 2425.180 2162.320 ;
        RECT 2415.575 2161.310 2418.130 2161.450 ;
        RECT 2415.575 2161.145 2415.855 2161.310 ;
        RECT 2417.850 2161.195 2418.130 2161.310 ;
        RECT 2424.930 2161.140 2425.255 2161.465 ;
        RECT 2425.000 2158.115 2425.170 2161.140 ;
        RECT 2424.930 2157.790 2425.255 2158.115 ;
        RECT 2421.320 2056.125 2421.660 2056.475 ;
        RECT 2421.405 2052.650 2421.575 2056.125 ;
        RECT 2420.680 2052.510 2421.575 2052.650 ;
        RECT 2420.680 2052.085 2420.820 2052.510 ;
        RECT 2421.405 2052.370 2421.575 2052.510 ;
        RECT 2420.610 2051.715 2420.890 2052.085 ;
        RECT 2421.330 2052.020 2421.670 2052.370 ;
        RECT 2424.625 1951.135 2425.005 1951.515 ;
        RECT 2430.260 1951.135 2430.600 1951.485 ;
        RECT 2430.345 1947.350 2430.515 1951.135 ;
        RECT 2430.270 1947.000 2430.610 1947.350 ;
        RECT 2424.750 1789.915 2425.030 1790.285 ;
        RECT 2424.820 1788.445 2424.960 1789.915 ;
        RECT 2424.760 1788.125 2425.020 1788.445 ;
        RECT 2427.010 1788.150 2427.350 1788.500 ;
        RECT 2427.090 1784.350 2427.260 1788.150 ;
        RECT 2427.010 1784.000 2427.350 1784.350 ;
        RECT 2422.910 1759.315 2423.190 1759.685 ;
        RECT 2422.980 1711.405 2423.120 1759.315 ;
        RECT 2422.910 1711.035 2423.190 1711.405 ;
        RECT 2413.890 1709.310 2422.975 1709.480 ;
        RECT 2411.525 1708.140 2411.805 1708.510 ;
        RECT 2413.890 1708.495 2414.060 1709.310 ;
        RECT 2413.835 1708.155 2414.115 1708.495 ;
        RECT 2421.990 1708.315 2422.270 1708.685 ;
        RECT 2422.800 1708.485 2422.975 1709.310 ;
        RECT 2422.060 1705.270 2422.200 1708.315 ;
        RECT 2422.735 1708.160 2423.060 1708.485 ;
        RECT 2422.000 1705.175 2422.260 1705.270 ;
        RECT 2422.800 1705.265 2422.975 1708.160 ;
        RECT 2422.730 1705.175 2423.055 1705.265 ;
        RECT 2422.000 1705.035 2423.055 1705.175 ;
        RECT 2422.000 1704.950 2422.260 1705.035 ;
        RECT 2422.730 1704.940 2423.055 1705.035 ;
        RECT 2422.835 1702.490 2422.975 1704.940 ;
        RECT 2422.060 1702.350 2422.975 1702.490 ;
        RECT 2422.060 1697.010 2422.200 1702.350 ;
        RECT 2421.600 1696.870 2422.200 1697.010 ;
        RECT 2421.600 1610.765 2421.740 1696.870 ;
        RECT 2421.530 1610.395 2421.810 1610.765 ;
        RECT 2415.605 1609.240 2425.155 1609.410 ;
        RECT 2415.605 1608.610 2415.775 1609.240 ;
        RECT 2413.185 1608.135 2413.560 1608.505 ;
        RECT 2415.605 1608.485 2417.600 1608.610 ;
        RECT 2415.550 1608.470 2417.600 1608.485 ;
        RECT 2415.550 1608.145 2415.830 1608.470 ;
        RECT 2417.460 1608.045 2417.600 1608.470 ;
        RECT 2424.985 1608.465 2425.155 1609.240 ;
        RECT 2424.905 1608.140 2425.230 1608.465 ;
        RECT 2417.390 1607.675 2417.670 1608.045 ;
        RECT 2424.975 1605.115 2425.145 1608.140 ;
        RECT 2424.905 1604.790 2425.230 1605.115 ;
        RECT 2415.725 1531.130 2416.015 1531.510 ;
        RECT 2421.315 1531.125 2421.655 1531.475 ;
        RECT 2420.610 1527.690 2420.890 1527.805 ;
        RECT 2421.400 1527.690 2421.570 1531.125 ;
        RECT 2420.610 1527.550 2421.570 1527.690 ;
        RECT 2420.610 1527.435 2420.890 1527.550 ;
        RECT 2421.400 1527.350 2421.570 1527.550 ;
        RECT 2421.325 1527.000 2421.665 1527.350 ;
        RECT 2423.830 1433.170 2424.110 1433.285 ;
        RECT 2424.760 1433.170 2425.020 1433.430 ;
        RECT 2423.830 1433.110 2425.020 1433.170 ;
        RECT 2430.255 1433.135 2430.595 1433.485 ;
        RECT 2423.830 1433.030 2424.960 1433.110 ;
        RECT 2423.830 1432.915 2424.110 1433.030 ;
        RECT 2430.340 1429.350 2430.510 1433.135 ;
        RECT 2430.265 1429.000 2430.605 1429.350 ;
        RECT 2427.510 1362.875 2427.790 1363.245 ;
        RECT 2427.580 1336.725 2427.720 1362.875 ;
        RECT 2427.510 1336.355 2427.790 1336.725 ;
        RECT 2427.050 1334.995 2427.330 1335.365 ;
        RECT 2421.460 1333.135 2421.750 1333.515 ;
        RECT 2427.120 1333.500 2427.260 1334.995 ;
        RECT 2427.060 1333.150 2427.400 1333.500 ;
        RECT 2427.120 1333.070 2427.310 1333.150 ;
        RECT 2427.140 1329.350 2427.310 1333.070 ;
        RECT 2427.060 1329.000 2427.400 1329.350 ;
      LAYER met3 ;
        RECT 2411.135 2253.125 2411.475 2257.455 ;
        RECT 2413.230 2161.510 2413.560 2165.445 ;
        RECT 2418.285 2164.260 2418.615 2164.265 ;
        RECT 2418.030 2164.250 2418.615 2164.260 ;
        RECT 2417.830 2163.950 2418.615 2164.250 ;
        RECT 2418.030 2163.940 2418.615 2163.950 ;
        RECT 2418.285 2163.935 2418.615 2163.940 ;
        RECT 2417.825 2161.540 2418.155 2161.545 ;
        RECT 2417.825 2161.530 2418.410 2161.540 ;
        RECT 2413.205 2161.140 2413.580 2161.510 ;
        RECT 2417.600 2161.230 2418.410 2161.530 ;
        RECT 2417.825 2161.220 2418.410 2161.230 ;
        RECT 2417.825 2161.215 2418.155 2161.220 ;
        RECT 2420.585 2052.060 2420.915 2052.065 ;
        RECT 2420.585 2052.050 2421.170 2052.060 ;
        RECT 2420.360 2051.750 2421.170 2052.050 ;
        RECT 2420.585 2051.740 2421.170 2051.750 ;
        RECT 2420.585 2051.735 2420.915 2051.740 ;
        RECT 2424.650 1951.515 2424.975 1955.360 ;
        RECT 2424.500 1951.135 2425.005 1951.515 ;
        RECT 2424.725 1790.260 2425.055 1790.265 ;
        RECT 2424.470 1790.250 2425.055 1790.260 ;
        RECT 2424.470 1789.950 2425.280 1790.250 ;
        RECT 2424.470 1789.940 2425.055 1789.950 ;
        RECT 2424.725 1789.935 2425.055 1789.940 ;
        RECT 2422.885 1759.650 2423.215 1759.665 ;
        RECT 2427.230 1759.650 2427.610 1759.660 ;
        RECT 2917.600 1759.650 2924.800 1760.100 ;
        RECT 2422.885 1759.350 2924.800 1759.650 ;
        RECT 2422.885 1759.335 2423.215 1759.350 ;
        RECT 2427.230 1759.340 2427.610 1759.350 ;
        RECT 2917.600 1758.900 2924.800 1759.350 ;
        RECT 2411.495 1708.140 2411.835 1712.470 ;
        RECT 2422.885 1711.370 2423.215 1711.385 ;
        RECT 2422.670 1711.055 2423.215 1711.370 ;
        RECT 2421.965 1708.650 2422.295 1708.665 ;
        RECT 2422.670 1708.650 2422.970 1711.055 ;
        RECT 2421.965 1708.350 2422.970 1708.650 ;
        RECT 2421.965 1708.335 2422.295 1708.350 ;
        RECT 2413.205 1608.505 2413.540 1612.385 ;
        RECT 2418.030 1610.730 2418.410 1610.740 ;
        RECT 2421.505 1610.730 2421.835 1610.745 ;
        RECT 2418.030 1610.430 2421.835 1610.730 ;
        RECT 2418.030 1610.420 2418.410 1610.430 ;
        RECT 2421.505 1610.415 2421.835 1610.430 ;
        RECT 2413.185 1608.135 2413.560 1608.505 ;
        RECT 2417.365 1608.010 2417.695 1608.025 ;
        RECT 2418.030 1608.010 2418.410 1608.020 ;
        RECT 2417.365 1607.710 2418.410 1608.010 ;
        RECT 2417.365 1607.695 2417.695 1607.710 ;
        RECT 2418.030 1607.700 2418.410 1607.710 ;
        RECT 2415.690 1531.465 2416.040 1535.460 ;
        RECT 2415.695 1531.130 2416.045 1531.465 ;
        RECT 2420.585 1527.780 2420.915 1527.785 ;
        RECT 2420.585 1527.770 2421.170 1527.780 ;
        RECT 2420.360 1527.470 2421.170 1527.770 ;
        RECT 2420.585 1527.460 2421.170 1527.470 ;
        RECT 2420.585 1527.455 2420.915 1527.460 ;
        RECT 2420.790 1433.250 2421.170 1433.260 ;
        RECT 2423.805 1433.250 2424.135 1433.265 ;
        RECT 2420.790 1432.950 2424.135 1433.250 ;
        RECT 2420.790 1432.940 2421.170 1432.950 ;
        RECT 2423.805 1432.935 2424.135 1432.950 ;
        RECT 2420.790 1363.210 2421.170 1363.220 ;
        RECT 2427.485 1363.210 2427.815 1363.225 ;
        RECT 2420.790 1362.910 2427.815 1363.210 ;
        RECT 2420.790 1362.900 2421.170 1362.910 ;
        RECT 2427.485 1362.895 2427.815 1362.910 ;
        RECT 2421.430 1333.135 2421.780 1337.465 ;
        RECT 2427.485 1336.690 2427.815 1336.705 ;
        RECT 2427.270 1336.375 2427.815 1336.690 ;
        RECT 2427.270 1335.345 2427.570 1336.375 ;
        RECT 2427.025 1335.030 2427.570 1335.345 ;
        RECT 2427.025 1335.015 2427.355 1335.030 ;
      LAYER met4 ;
        RECT 2418.055 2163.935 2418.385 2164.265 ;
        RECT 2418.070 2161.545 2418.370 2163.935 ;
        RECT 2418.055 2161.215 2418.385 2161.545 ;
        RECT 2418.070 2159.850 2418.370 2161.215 ;
        RECT 2418.070 2159.550 2421.130 2159.850 ;
        RECT 2420.830 2052.065 2421.130 2159.550 ;
        RECT 2420.815 2051.735 2421.145 2052.065 ;
        RECT 2420.830 1966.650 2421.130 2051.735 ;
        RECT 2420.830 1966.350 2424.810 1966.650 ;
        RECT 2424.510 1951.490 2424.810 1966.350 ;
        RECT 2424.495 1951.160 2424.825 1951.490 ;
        RECT 2424.510 1790.265 2424.810 1951.160 ;
        RECT 2424.495 1789.935 2424.825 1790.265 ;
        RECT 2424.510 1773.450 2424.810 1789.935 ;
        RECT 2424.510 1773.150 2427.570 1773.450 ;
        RECT 2427.270 1759.665 2427.570 1773.150 ;
        RECT 2427.255 1759.335 2427.585 1759.665 ;
        RECT 2418.055 1610.415 2418.385 1610.745 ;
        RECT 2418.070 1608.025 2418.370 1610.415 ;
        RECT 2418.055 1607.695 2418.385 1608.025 ;
        RECT 2418.070 1580.250 2418.370 1607.695 ;
        RECT 2418.070 1579.950 2421.130 1580.250 ;
        RECT 2420.830 1527.785 2421.130 1579.950 ;
        RECT 2420.815 1527.455 2421.145 1527.785 ;
        RECT 2420.830 1433.265 2421.130 1527.455 ;
        RECT 2420.815 1432.935 2421.145 1433.265 ;
        RECT 2420.830 1363.225 2421.130 1432.935 ;
        RECT 2420.815 1362.895 2421.145 1363.225 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.289999 ;
    PORT
      LAYER li1 ;
        RECT 2427.800 2253.225 2427.970 2254.495 ;
        RECT 2439.025 2253.230 2439.195 2254.500 ;
        RECT 2439.025 2247.960 2439.195 2249.230 ;
        RECT 2430.540 2161.225 2430.710 2162.495 ;
        RECT 2442.225 2161.465 2442.395 2162.505 ;
        RECT 2442.220 2161.225 2442.400 2161.465 ;
        RECT 2442.225 2155.955 2442.395 2157.225 ;
        RECT 2432.110 2056.235 2432.280 2057.505 ;
        RECT 2437.725 2056.235 2437.895 2057.505 ;
        RECT 2437.725 2050.955 2437.895 2052.225 ;
        RECT 2443.285 1951.240 2443.455 1952.510 ;
        RECT 2448.900 1951.240 2449.070 1952.510 ;
        RECT 2448.900 1945.955 2449.070 1947.225 ;
        RECT 2436.730 1788.240 2436.900 1789.510 ;
        RECT 2442.345 1788.240 2442.515 1789.510 ;
        RECT 2442.345 1782.955 2442.515 1784.225 ;
        RECT 2428.160 1708.235 2428.330 1709.505 ;
        RECT 2439.385 1708.240 2439.555 1709.510 ;
        RECT 2439.385 1702.970 2439.555 1704.240 ;
        RECT 2430.515 1608.235 2430.685 1609.505 ;
        RECT 2442.200 1608.465 2442.370 1609.505 ;
        RECT 2442.195 1608.225 2442.375 1608.465 ;
        RECT 2442.200 1602.955 2442.370 1604.225 ;
        RECT 2432.105 1531.235 2432.275 1532.505 ;
        RECT 2437.720 1531.235 2437.890 1532.505 ;
        RECT 2437.720 1525.955 2437.890 1527.225 ;
        RECT 2443.280 1433.240 2443.450 1434.510 ;
        RECT 2448.895 1433.240 2449.065 1434.510 ;
        RECT 2448.895 1427.955 2449.065 1429.225 ;
        RECT 2436.780 1333.240 2436.950 1334.510 ;
        RECT 2442.395 1333.240 2442.565 1334.510 ;
        RECT 2442.395 1327.955 2442.565 1329.225 ;
      LAYER met1 ;
        RECT 2427.715 2253.400 2428.055 2253.450 ;
        RECT 2427.715 2253.395 2428.060 2253.400 ;
        RECT 2427.715 2253.365 2428.200 2253.395 ;
        RECT 2430.025 2253.365 2430.365 2253.455 ;
        RECT 2427.715 2253.190 2430.365 2253.365 ;
        RECT 2427.715 2253.170 2428.055 2253.190 ;
        RECT 2430.025 2253.175 2430.365 2253.190 ;
        RECT 2438.955 2253.400 2439.280 2253.475 ;
        RECT 2438.955 2253.230 2439.425 2253.400 ;
        RECT 2438.955 2253.150 2439.280 2253.230 ;
        RECT 2438.950 2249.930 2439.275 2250.255 ;
        RECT 2439.025 2249.260 2439.205 2249.930 ;
        RECT 2438.965 2249.230 2439.255 2249.260 ;
        RECT 2438.965 2249.060 2439.425 2249.230 ;
        RECT 2438.965 2249.030 2439.255 2249.060 ;
        RECT 2430.445 2161.400 2430.785 2161.495 ;
        RECT 2430.445 2161.395 2430.800 2161.400 ;
        RECT 2430.445 2161.365 2430.940 2161.395 ;
        RECT 2432.765 2161.365 2433.105 2161.455 ;
        RECT 2430.445 2161.200 2433.105 2161.365 ;
        RECT 2430.445 2161.155 2430.785 2161.200 ;
        RECT 2432.765 2161.175 2433.105 2161.200 ;
        RECT 2442.150 2161.405 2442.475 2161.465 ;
        RECT 2442.150 2161.235 2442.625 2161.405 ;
        RECT 2442.150 2161.140 2442.475 2161.235 ;
        RECT 2442.150 2157.790 2442.475 2158.115 ;
        RECT 2442.230 2157.255 2442.400 2157.790 ;
        RECT 2442.165 2157.225 2442.455 2157.255 ;
        RECT 2442.165 2157.055 2442.625 2157.225 ;
        RECT 2442.165 2157.025 2442.455 2157.055 ;
        RECT 2432.035 2056.405 2432.355 2056.465 ;
        RECT 2437.645 2056.405 2437.985 2056.475 ;
        RECT 2432.035 2056.375 2432.510 2056.405 ;
        RECT 2437.645 2056.400 2438.125 2056.405 ;
        RECT 2437.630 2056.375 2438.125 2056.400 ;
        RECT 2432.035 2056.235 2438.125 2056.375 ;
        RECT 2432.035 2056.205 2437.985 2056.235 ;
        RECT 2432.035 2056.175 2432.355 2056.205 ;
        RECT 2437.645 2056.125 2437.985 2056.205 ;
        RECT 2437.655 2052.225 2437.995 2052.370 ;
        RECT 2437.655 2052.055 2438.125 2052.225 ;
        RECT 2437.655 2052.015 2437.995 2052.055 ;
        RECT 2443.200 1951.410 2443.550 1951.500 ;
        RECT 2448.820 1951.410 2449.160 1951.485 ;
        RECT 2443.200 1951.380 2443.685 1951.410 ;
        RECT 2448.820 1951.405 2449.300 1951.410 ;
        RECT 2448.805 1951.380 2449.305 1951.405 ;
        RECT 2443.200 1951.235 2449.305 1951.380 ;
        RECT 2443.200 1951.200 2449.160 1951.235 ;
        RECT 2443.200 1951.150 2443.550 1951.200 ;
        RECT 2448.820 1951.135 2449.160 1951.200 ;
        RECT 2448.830 1947.225 2449.170 1947.350 ;
        RECT 2448.830 1947.055 2449.300 1947.225 ;
        RECT 2448.830 1947.000 2449.170 1947.055 ;
        RECT 2436.640 1788.410 2436.990 1788.470 ;
        RECT 2442.270 1788.410 2442.610 1788.500 ;
        RECT 2436.640 1788.370 2437.130 1788.410 ;
        RECT 2442.270 1788.405 2442.745 1788.410 ;
        RECT 2442.250 1788.370 2442.745 1788.405 ;
        RECT 2436.640 1788.240 2442.745 1788.370 ;
        RECT 2436.640 1788.205 2442.610 1788.240 ;
        RECT 2436.640 1788.180 2436.990 1788.205 ;
        RECT 2442.270 1788.150 2442.610 1788.205 ;
        RECT 2442.270 1784.225 2442.610 1784.350 ;
        RECT 2442.270 1784.055 2442.745 1784.225 ;
        RECT 2442.270 1784.000 2442.610 1784.055 ;
        RECT 2428.075 1708.405 2428.415 1708.465 ;
        RECT 2428.075 1708.375 2428.560 1708.405 ;
        RECT 2430.385 1708.375 2430.725 1708.465 ;
        RECT 2428.075 1708.205 2430.725 1708.375 ;
        RECT 2428.075 1708.185 2428.415 1708.205 ;
        RECT 2430.385 1708.185 2430.725 1708.205 ;
        RECT 2439.315 1708.410 2439.640 1708.485 ;
        RECT 2439.315 1708.240 2439.785 1708.410 ;
        RECT 2439.315 1708.160 2439.640 1708.240 ;
        RECT 2439.310 1704.940 2439.635 1705.265 ;
        RECT 2439.385 1704.270 2439.565 1704.940 ;
        RECT 2439.325 1704.240 2439.615 1704.270 ;
        RECT 2439.325 1704.070 2439.785 1704.240 ;
        RECT 2439.325 1704.040 2439.615 1704.070 ;
        RECT 2430.425 1608.405 2430.765 1608.490 ;
        RECT 2430.425 1608.375 2430.915 1608.405 ;
        RECT 2432.740 1608.375 2433.080 1608.455 ;
        RECT 2430.425 1608.200 2433.080 1608.375 ;
        RECT 2430.425 1608.150 2430.765 1608.200 ;
        RECT 2432.740 1608.175 2433.080 1608.200 ;
        RECT 2442.125 1608.405 2442.450 1608.465 ;
        RECT 2442.125 1608.235 2442.600 1608.405 ;
        RECT 2442.125 1608.140 2442.450 1608.235 ;
        RECT 2442.125 1604.790 2442.450 1605.115 ;
        RECT 2442.205 1604.255 2442.375 1604.790 ;
        RECT 2442.140 1604.225 2442.430 1604.255 ;
        RECT 2442.140 1604.055 2442.600 1604.225 ;
        RECT 2442.140 1604.025 2442.430 1604.055 ;
        RECT 2432.020 1531.405 2432.370 1531.465 ;
        RECT 2437.640 1531.405 2437.980 1531.475 ;
        RECT 2432.020 1531.375 2432.505 1531.405 ;
        RECT 2437.640 1531.400 2438.120 1531.405 ;
        RECT 2437.625 1531.375 2438.120 1531.400 ;
        RECT 2432.020 1531.235 2438.120 1531.375 ;
        RECT 2432.020 1531.205 2437.980 1531.235 ;
        RECT 2432.020 1531.175 2432.370 1531.205 ;
        RECT 2437.640 1531.125 2437.980 1531.205 ;
        RECT 2437.650 1527.225 2437.990 1527.350 ;
        RECT 2437.650 1527.055 2438.120 1527.225 ;
        RECT 2437.650 1527.000 2437.990 1527.055 ;
        RECT 2443.190 1433.430 2443.540 1433.495 ;
        RECT 2443.160 1433.410 2443.540 1433.430 ;
        RECT 2448.815 1433.410 2449.155 1433.485 ;
        RECT 2443.160 1433.380 2443.680 1433.410 ;
        RECT 2448.815 1433.405 2449.295 1433.410 ;
        RECT 2448.800 1433.380 2449.300 1433.405 ;
        RECT 2443.160 1433.235 2449.300 1433.380 ;
        RECT 2443.160 1433.210 2449.155 1433.235 ;
        RECT 2443.160 1433.145 2443.540 1433.210 ;
        RECT 2443.160 1433.110 2443.420 1433.145 ;
        RECT 2448.815 1433.135 2449.155 1433.210 ;
        RECT 2448.825 1429.225 2449.165 1429.350 ;
        RECT 2448.825 1429.055 2449.295 1429.225 ;
        RECT 2448.825 1429.000 2449.165 1429.055 ;
        RECT 2436.690 1333.410 2437.040 1333.470 ;
        RECT 2442.320 1333.410 2442.660 1333.500 ;
        RECT 2436.690 1333.380 2437.180 1333.410 ;
        RECT 2442.320 1333.405 2442.795 1333.410 ;
        RECT 2442.300 1333.380 2442.795 1333.405 ;
        RECT 2436.690 1333.240 2442.795 1333.380 ;
        RECT 2436.690 1333.205 2442.660 1333.240 ;
        RECT 2436.690 1333.180 2437.040 1333.205 ;
        RECT 2442.320 1333.150 2442.660 1333.205 ;
        RECT 2442.320 1329.225 2442.660 1329.350 ;
        RECT 2442.320 1329.055 2442.795 1329.225 ;
        RECT 2442.320 1329.000 2442.660 1329.055 ;
      LAYER met2 ;
        RECT 2430.110 2254.315 2439.195 2254.485 ;
        RECT 2427.745 2253.125 2428.025 2253.495 ;
        RECT 2430.110 2253.485 2430.280 2254.315 ;
        RECT 2430.055 2253.145 2430.335 2253.485 ;
        RECT 2439.020 2253.475 2439.195 2254.315 ;
        RECT 2438.955 2253.150 2439.280 2253.475 ;
        RECT 2439.020 2251.325 2439.195 2253.150 ;
        RECT 2438.965 2250.955 2439.245 2251.325 ;
        RECT 2439.020 2250.255 2439.195 2250.955 ;
        RECT 2438.950 2249.930 2439.275 2250.255 ;
        RECT 2432.850 2162.320 2442.400 2162.490 ;
        RECT 2430.425 2161.140 2430.800 2161.510 ;
        RECT 2432.850 2161.485 2433.020 2162.320 ;
        RECT 2432.795 2161.145 2433.075 2161.485 ;
        RECT 2442.230 2161.465 2442.400 2162.320 ;
        RECT 2442.150 2161.140 2442.475 2161.465 ;
        RECT 2442.220 2158.165 2442.390 2161.140 ;
        RECT 2442.165 2158.115 2442.445 2158.165 ;
        RECT 2442.150 2157.790 2442.475 2158.115 ;
        RECT 2442.690 2069.395 2442.970 2069.765 ;
        RECT 2437.645 2056.125 2437.985 2056.475 ;
        RECT 2437.730 2052.370 2437.900 2056.125 ;
        RECT 2437.655 2052.020 2437.995 2052.370 ;
        RECT 2437.745 2051.290 2437.885 2052.020 ;
        RECT 2437.745 2051.150 2438.300 2051.290 ;
        RECT 2438.160 2050.045 2438.300 2051.150 ;
        RECT 2442.760 2050.045 2442.900 2069.395 ;
        RECT 2438.090 2049.675 2438.370 2050.045 ;
        RECT 2442.690 2049.675 2442.970 2050.045 ;
        RECT 2449.130 2049.675 2449.410 2050.045 ;
        RECT 2900.850 2049.675 2901.130 2050.045 ;
        RECT 2449.200 1960.285 2449.340 2049.675 ;
        RECT 2900.920 2024.885 2901.060 2049.675 ;
        RECT 2900.850 2024.515 2901.130 2024.885 ;
        RECT 2449.130 1959.915 2449.410 1960.285 ;
        RECT 2443.185 1951.135 2443.565 1951.515 ;
        RECT 2448.820 1951.135 2449.160 1951.485 ;
        RECT 2446.830 1947.250 2447.110 1947.365 ;
        RECT 2448.905 1947.350 2449.075 1951.135 ;
        RECT 2448.830 1947.250 2449.170 1947.350 ;
        RECT 2446.830 1947.110 2449.170 1947.250 ;
        RECT 2446.830 1946.995 2447.110 1947.110 ;
        RECT 2448.830 1947.000 2449.170 1947.110 ;
        RECT 2442.230 1789.915 2442.510 1790.285 ;
        RECT 2442.300 1788.810 2442.440 1789.915 ;
        RECT 2442.300 1788.670 2442.505 1788.810 ;
        RECT 2442.365 1788.500 2442.505 1788.670 ;
        RECT 2442.270 1788.150 2442.610 1788.500 ;
        RECT 2442.350 1784.350 2442.520 1788.150 ;
        RECT 2442.270 1784.000 2442.610 1784.350 ;
        RECT 2430.470 1709.310 2439.555 1709.480 ;
        RECT 2428.105 1708.140 2428.385 1708.510 ;
        RECT 2430.470 1708.495 2430.640 1709.310 ;
        RECT 2430.415 1708.155 2430.695 1708.495 ;
        RECT 2439.380 1708.485 2439.555 1709.310 ;
        RECT 2439.315 1708.160 2439.640 1708.485 ;
        RECT 2439.380 1705.265 2439.555 1708.160 ;
        RECT 2439.310 1705.240 2439.635 1705.265 ;
        RECT 2439.310 1704.960 2439.795 1705.240 ;
        RECT 2439.310 1704.940 2439.635 1704.960 ;
        RECT 2432.825 1609.240 2442.375 1609.410 ;
        RECT 2430.405 1608.135 2430.780 1608.505 ;
        RECT 2432.825 1608.485 2432.995 1609.240 ;
        RECT 2432.770 1608.145 2433.050 1608.485 ;
        RECT 2442.205 1608.465 2442.375 1609.240 ;
        RECT 2442.125 1608.140 2442.450 1608.465 ;
        RECT 2440.850 1605.210 2441.130 1605.325 ;
        RECT 2442.195 1605.210 2442.365 1608.140 ;
        RECT 2440.850 1605.115 2442.365 1605.210 ;
        RECT 2440.850 1605.070 2442.450 1605.115 ;
        RECT 2440.850 1604.955 2441.130 1605.070 ;
        RECT 2442.125 1604.790 2442.450 1605.070 ;
        RECT 2432.050 1531.130 2432.340 1531.510 ;
        RECT 2437.640 1531.160 2437.980 1531.475 ;
        RECT 2437.625 1530.880 2437.995 1531.160 ;
        RECT 2437.725 1527.350 2437.895 1530.880 ;
        RECT 2437.650 1527.000 2437.990 1527.350 ;
        RECT 2442.690 1433.170 2442.970 1433.285 ;
        RECT 2443.160 1433.170 2443.420 1433.430 ;
        RECT 2442.690 1433.110 2443.420 1433.170 ;
        RECT 2448.815 1433.135 2449.155 1433.485 ;
        RECT 2442.690 1433.030 2443.360 1433.110 ;
        RECT 2442.690 1432.915 2442.970 1433.030 ;
        RECT 2448.900 1429.350 2449.070 1433.135 ;
        RECT 2448.825 1429.000 2449.165 1429.350 ;
        RECT 2442.230 1334.995 2442.510 1335.365 ;
        RECT 2436.720 1333.135 2437.010 1333.515 ;
        RECT 2442.300 1333.500 2442.440 1334.995 ;
        RECT 2442.300 1333.150 2442.660 1333.500 ;
        RECT 2442.300 1333.070 2442.570 1333.150 ;
        RECT 2442.400 1329.350 2442.570 1333.070 ;
        RECT 2442.320 1329.000 2442.660 1329.350 ;
      LAYER met3 ;
        RECT 2427.715 2253.125 2428.055 2257.455 ;
        RECT 2438.940 2251.300 2439.270 2251.305 ;
        RECT 2438.940 2251.290 2439.570 2251.300 ;
        RECT 2438.940 2250.990 2439.725 2251.290 ;
        RECT 2438.940 2250.980 2439.570 2250.990 ;
        RECT 2438.940 2250.975 2439.270 2250.980 ;
        RECT 2430.450 2161.510 2430.780 2165.445 ;
        RECT 2430.425 2161.140 2430.800 2161.510 ;
        RECT 2442.140 2158.140 2442.470 2158.145 ;
        RECT 2441.950 2158.130 2442.470 2158.140 ;
        RECT 2441.950 2157.830 2442.760 2158.130 ;
        RECT 2441.950 2157.820 2442.470 2157.830 ;
        RECT 2442.140 2157.815 2442.470 2157.820 ;
        RECT 2441.950 2069.730 2442.330 2069.740 ;
        RECT 2442.665 2069.730 2442.995 2069.745 ;
        RECT 2441.950 2069.430 2442.995 2069.730 ;
        RECT 2441.950 2069.420 2442.330 2069.430 ;
        RECT 2442.665 2069.415 2442.995 2069.430 ;
        RECT 2438.065 2050.010 2438.395 2050.025 ;
        RECT 2442.665 2050.010 2442.995 2050.025 ;
        RECT 2449.105 2050.010 2449.435 2050.025 ;
        RECT 2900.825 2050.010 2901.155 2050.025 ;
        RECT 2438.065 2049.710 2901.155 2050.010 ;
        RECT 2438.065 2049.695 2438.395 2049.710 ;
        RECT 2442.665 2049.695 2442.995 2049.710 ;
        RECT 2449.105 2049.695 2449.435 2049.710 ;
        RECT 2900.825 2049.695 2901.155 2049.710 ;
        RECT 2900.825 2024.850 2901.155 2024.865 ;
        RECT 2917.600 2024.850 2924.800 2025.300 ;
        RECT 2900.825 2024.550 2924.800 2024.850 ;
        RECT 2900.825 2024.535 2901.155 2024.550 ;
        RECT 2917.600 2024.100 2924.800 2024.550 ;
        RECT 2446.550 1960.250 2446.930 1960.260 ;
        RECT 2449.105 1960.250 2449.435 1960.265 ;
        RECT 2446.550 1959.950 2449.435 1960.250 ;
        RECT 2446.550 1959.940 2446.930 1959.950 ;
        RECT 2449.105 1959.935 2449.435 1959.950 ;
        RECT 2443.210 1951.515 2443.535 1955.360 ;
        RECT 2443.185 1951.135 2443.565 1951.515 ;
        RECT 2446.805 1947.340 2447.135 1947.345 ;
        RECT 2446.550 1947.330 2447.135 1947.340 ;
        RECT 2446.550 1947.030 2447.360 1947.330 ;
        RECT 2446.550 1947.020 2447.135 1947.030 ;
        RECT 2446.805 1947.015 2447.135 1947.020 ;
        RECT 2442.205 1790.260 2442.535 1790.265 ;
        RECT 2441.950 1790.250 2442.535 1790.260 ;
        RECT 2446.550 1790.250 2446.930 1790.260 ;
        RECT 2441.570 1789.950 2446.930 1790.250 ;
        RECT 2441.950 1789.940 2442.535 1789.950 ;
        RECT 2446.550 1789.940 2446.930 1789.950 ;
        RECT 2442.205 1789.935 2442.535 1789.940 ;
        RECT 2428.075 1708.140 2428.415 1712.470 ;
        RECT 2439.445 1705.250 2439.775 1705.265 ;
        RECT 2440.110 1705.250 2440.490 1705.260 ;
        RECT 2439.445 1704.950 2440.490 1705.250 ;
        RECT 2439.445 1704.935 2439.775 1704.950 ;
        RECT 2440.110 1704.940 2440.490 1704.950 ;
        RECT 2430.425 1608.505 2430.760 1612.385 ;
        RECT 2430.405 1608.135 2430.780 1608.505 ;
        RECT 2440.110 1605.290 2440.490 1605.300 ;
        RECT 2440.825 1605.290 2441.155 1605.305 ;
        RECT 2440.110 1604.990 2441.155 1605.290 ;
        RECT 2440.110 1604.980 2440.490 1604.990 ;
        RECT 2440.825 1604.975 2441.155 1604.990 ;
        RECT 2432.015 1531.465 2432.365 1535.460 ;
        RECT 2438.270 1531.540 2438.650 1531.860 ;
        RECT 2432.020 1531.130 2432.370 1531.465 ;
        RECT 2437.645 1531.170 2437.975 1531.185 ;
        RECT 2438.310 1531.170 2438.610 1531.540 ;
        RECT 2437.645 1530.870 2438.610 1531.170 ;
        RECT 2437.645 1530.855 2437.975 1530.870 ;
        RECT 2441.950 1433.620 2442.330 1433.940 ;
        RECT 2441.990 1433.250 2442.290 1433.620 ;
        RECT 2442.665 1433.250 2442.995 1433.265 ;
        RECT 2441.990 1432.950 2442.995 1433.250 ;
        RECT 2442.665 1432.935 2442.995 1432.950 ;
        RECT 2436.690 1333.135 2437.040 1337.465 ;
        RECT 2442.205 1335.340 2442.535 1335.345 ;
        RECT 2441.950 1335.330 2442.535 1335.340 ;
        RECT 2441.750 1335.030 2442.535 1335.330 ;
        RECT 2441.950 1335.020 2442.535 1335.030 ;
        RECT 2442.205 1335.015 2442.535 1335.020 ;
      LAYER met4 ;
        RECT 2439.215 2250.975 2439.545 2251.305 ;
        RECT 2439.230 2208.150 2439.530 2250.975 ;
        RECT 2439.230 2207.850 2442.290 2208.150 ;
        RECT 2441.990 2158.145 2442.290 2207.850 ;
        RECT 2441.975 2157.815 2442.305 2158.145 ;
        RECT 2441.990 2069.745 2442.290 2157.815 ;
        RECT 2441.975 2069.415 2442.305 2069.745 ;
        RECT 2446.575 1959.935 2446.905 1960.265 ;
        RECT 2446.590 1947.345 2446.890 1959.935 ;
        RECT 2446.575 1947.015 2446.905 1947.345 ;
        RECT 2446.590 1790.265 2446.890 1947.015 ;
        RECT 2441.975 1789.935 2442.305 1790.265 ;
        RECT 2446.575 1789.935 2446.905 1790.265 ;
        RECT 2441.990 1725.150 2442.290 1789.935 ;
        RECT 2440.150 1724.850 2442.290 1725.150 ;
        RECT 2440.150 1705.265 2440.450 1724.850 ;
        RECT 2440.135 1704.935 2440.465 1705.265 ;
        RECT 2440.150 1605.305 2440.450 1704.935 ;
        RECT 2440.135 1604.975 2440.465 1605.305 ;
        RECT 2440.150 1580.250 2440.450 1604.975 ;
        RECT 2438.310 1579.950 2440.450 1580.250 ;
        RECT 2438.310 1531.950 2438.610 1579.950 ;
        RECT 2438.310 1531.865 2442.290 1531.950 ;
        RECT 2438.295 1531.650 2442.290 1531.865 ;
        RECT 2438.295 1531.535 2438.625 1531.650 ;
        RECT 2441.990 1433.945 2442.290 1531.650 ;
        RECT 2441.975 1433.615 2442.305 1433.945 ;
        RECT 2441.990 1335.345 2442.290 1433.615 ;
        RECT 2441.975 1335.015 2442.305 1335.345 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2882.775 2422.920 2883.295 2424.405 ;
      LAYER met1 ;
        RECT 2882.985 2423.045 2883.305 2423.305 ;
      LAYER met2 ;
        RECT 2883.025 2423.335 2883.305 2423.375 ;
        RECT 2883.015 2423.015 2883.305 2423.335 ;
        RECT 2883.025 2423.005 2883.305 2423.015 ;
      LAYER met3 ;
        RECT 2883.000 2423.345 2883.330 2423.355 ;
        RECT 2883.000 2423.330 2908.700 2423.345 ;
        RECT 2917.600 2423.330 2924.800 2423.780 ;
        RECT 2883.000 2423.035 2924.800 2423.330 ;
        RECT 2883.000 2423.025 2883.330 2423.035 ;
        RECT 2904.935 2423.030 2924.800 2423.035 ;
        RECT 2917.600 2422.580 2924.800 2423.030 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2882.775 2688.800 2883.295 2690.285 ;
      LAYER met1 ;
        RECT 2882.985 2688.925 2883.305 2689.185 ;
      LAYER met2 ;
        RECT 2883.025 2689.215 2883.305 2689.255 ;
        RECT 2883.015 2688.895 2883.305 2689.215 ;
        RECT 2883.025 2688.885 2883.305 2688.895 ;
      LAYER met3 ;
        RECT 2883.000 2689.225 2883.330 2689.235 ;
        RECT 2883.000 2689.210 2907.740 2689.225 ;
        RECT 2917.600 2689.210 2924.800 2689.660 ;
        RECT 2883.000 2688.915 2924.800 2689.210 ;
        RECT 2883.000 2688.905 2883.330 2688.915 ;
        RECT 2904.950 2688.910 2924.800 2688.915 ;
        RECT 2917.600 2688.460 2924.800 2688.910 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2882.775 2954.680 2883.295 2956.165 ;
      LAYER met1 ;
        RECT 2882.985 2954.805 2883.305 2955.065 ;
      LAYER met2 ;
        RECT 2883.025 2955.095 2883.305 2955.135 ;
        RECT 2883.015 2954.775 2883.305 2955.095 ;
        RECT 2883.025 2954.765 2883.305 2954.775 ;
      LAYER met3 ;
        RECT 2883.000 2955.105 2883.330 2955.115 ;
        RECT 2883.000 2955.090 2908.325 2955.105 ;
        RECT 2917.600 2955.090 2924.800 2955.540 ;
        RECT 2883.000 2954.795 2924.800 2955.090 ;
        RECT 2883.000 2954.785 2883.330 2954.795 ;
        RECT 2904.950 2954.790 2924.800 2954.795 ;
        RECT 2917.600 2954.340 2924.800 2954.790 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2882.775 3219.880 2883.295 3221.365 ;
      LAYER met1 ;
        RECT 2882.985 3220.005 2883.305 3220.265 ;
      LAYER met2 ;
        RECT 2883.025 3220.295 2883.305 3220.335 ;
        RECT 2883.015 3219.975 2883.305 3220.295 ;
        RECT 2883.025 3219.965 2883.305 3219.975 ;
      LAYER met3 ;
        RECT 2883.000 3220.305 2883.330 3220.315 ;
        RECT 2883.000 3220.290 2906.310 3220.305 ;
        RECT 2917.600 3220.290 2924.800 3220.740 ;
        RECT 2883.000 3219.995 2924.800 3220.290 ;
        RECT 2883.000 3219.985 2883.330 3219.995 ;
        RECT 2905.140 3219.990 2924.800 3219.995 ;
        RECT 2917.600 3219.540 2924.800 3219.990 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2882.775 3485.760 2883.295 3487.245 ;
      LAYER met1 ;
        RECT 2882.985 3485.885 2883.305 3486.145 ;
      LAYER met2 ;
        RECT 2883.025 3486.175 2883.305 3486.215 ;
        RECT 2883.015 3485.855 2883.305 3486.175 ;
        RECT 2883.025 3485.845 2883.305 3485.855 ;
        RECT 2904.530 3485.835 2904.810 3486.205 ;
      LAYER met3 ;
        RECT 2883.000 3486.185 2883.330 3486.195 ;
        RECT 2883.000 3486.170 2906.190 3486.185 ;
        RECT 2917.600 3486.170 2924.800 3486.620 ;
        RECT 2883.000 3485.875 2924.800 3486.170 ;
        RECT 2883.000 3485.865 2883.330 3485.875 ;
        RECT 2904.505 3485.870 2924.800 3485.875 ;
        RECT 2904.505 3485.855 2904.835 3485.870 ;
        RECT 2917.600 3485.420 2924.800 3485.870 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2523.580 3508.780 2524.100 3510.330 ;
      LAYER met1 ;
        RECT 2523.630 3508.905 2523.950 3509.165 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2523.660 3509.165 2523.915 3509.195 ;
        RECT 2523.630 3509.110 2523.950 3509.165 ;
        RECT 2635.960 3509.110 2636.100 3517.600 ;
        RECT 2523.630 3508.945 2636.100 3509.110 ;
        RECT 2523.630 3508.905 2523.950 3508.945 ;
        RECT 2635.960 3508.930 2636.100 3508.945 ;
        RECT 2523.660 3508.875 2523.915 3508.905 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2163.580 3508.095 2164.100 3509.645 ;
      LAYER met1 ;
        RECT 2163.630 3508.220 2163.950 3508.480 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2163.660 3508.480 2163.915 3508.510 ;
        RECT 2163.630 3508.425 2163.950 3508.480 ;
        RECT 2311.660 3508.425 2311.800 3517.600 ;
        RECT 2163.630 3508.260 2311.800 3508.425 ;
        RECT 2163.630 3508.220 2163.950 3508.260 ;
        RECT 2311.660 3508.255 2311.800 3508.260 ;
        RECT 2163.660 3508.190 2163.915 3508.220 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1803.580 3508.455 1804.100 3510.005 ;
      LAYER met1 ;
        RECT 1803.630 3508.580 1803.950 3508.840 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1803.660 3508.840 1803.915 3508.870 ;
        RECT 1803.630 3508.785 1803.950 3508.840 ;
        RECT 1987.360 3508.785 1987.500 3517.600 ;
        RECT 1803.630 3508.625 1987.500 3508.785 ;
        RECT 1803.630 3508.620 1987.085 3508.625 ;
        RECT 1803.630 3508.580 1803.950 3508.620 ;
        RECT 1803.660 3508.550 1803.915 3508.580 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1623.580 3510.375 1624.100 3511.925 ;
      LAYER met1 ;
        RECT 1623.630 3510.500 1623.950 3510.760 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1623.660 3510.760 1623.915 3510.790 ;
        RECT 1623.630 3510.705 1623.950 3510.760 ;
        RECT 1662.600 3510.705 1662.740 3517.600 ;
        RECT 1623.630 3510.550 1662.740 3510.705 ;
        RECT 1623.630 3510.540 1662.405 3510.550 ;
        RECT 1623.630 3510.500 1623.950 3510.540 ;
        RECT 1623.660 3510.470 1623.915 3510.500 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1263.580 3509.925 1264.100 3511.475 ;
      LAYER met1 ;
        RECT 1263.630 3510.050 1263.950 3510.310 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1263.660 3510.310 1263.915 3510.340 ;
        RECT 1263.630 3510.255 1263.950 3510.310 ;
        RECT 1338.300 3510.255 1338.440 3517.600 ;
        RECT 1263.630 3510.090 1338.440 3510.255 ;
        RECT 1263.630 3510.050 1263.950 3510.090 ;
        RECT 1338.300 3510.085 1338.440 3510.090 ;
        RECT 1263.660 3510.020 1263.915 3510.050 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2882.775 1161.520 2883.295 1163.005 ;
      LAYER met1 ;
        RECT 2882.985 1161.645 2883.305 1161.905 ;
      LAYER met2 ;
        RECT 2883.025 1161.935 2883.305 1161.975 ;
        RECT 2883.015 1161.615 2883.305 1161.935 ;
        RECT 2883.025 1161.605 2883.305 1161.615 ;
      LAYER met3 ;
        RECT 2883.000 1161.945 2883.330 1161.955 ;
        RECT 2883.000 1161.930 2907.110 1161.945 ;
        RECT 2917.600 1161.930 2924.800 1162.380 ;
        RECT 2883.000 1161.635 2924.800 1161.930 ;
        RECT 2883.000 1161.625 2883.330 1161.635 ;
        RECT 2905.145 1161.630 2924.800 1161.635 ;
        RECT 2917.600 1161.180 2924.800 1161.630 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2882.775 1360.760 2883.295 1362.245 ;
      LAYER met1 ;
        RECT 2882.985 1360.885 2883.305 1361.145 ;
      LAYER met2 ;
        RECT 2883.025 1361.175 2883.305 1361.215 ;
        RECT 2883.015 1360.855 2883.305 1361.175 ;
        RECT 2883.025 1360.845 2883.305 1360.855 ;
      LAYER met3 ;
        RECT 2883.000 1361.185 2883.330 1361.195 ;
        RECT 2883.000 1361.170 2908.560 1361.185 ;
        RECT 2917.600 1361.170 2924.800 1361.620 ;
        RECT 2883.000 1360.875 2924.800 1361.170 ;
        RECT 2883.000 1360.865 2883.330 1360.875 ;
        RECT 2904.990 1360.870 2924.800 1360.875 ;
        RECT 2917.600 1360.420 2924.800 1360.870 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2882.775 1625.960 2883.295 1627.445 ;
      LAYER met1 ;
        RECT 2882.985 1626.085 2883.305 1626.345 ;
      LAYER met2 ;
        RECT 2883.025 1626.375 2883.305 1626.415 ;
        RECT 2883.015 1626.055 2883.305 1626.375 ;
        RECT 2883.025 1626.045 2883.305 1626.055 ;
      LAYER met3 ;
        RECT 2883.000 1626.385 2883.330 1626.395 ;
        RECT 2883.000 1626.370 2906.955 1626.385 ;
        RECT 2917.600 1626.370 2924.800 1626.820 ;
        RECT 2883.000 1626.075 2924.800 1626.370 ;
        RECT 2883.000 1626.065 2883.330 1626.075 ;
        RECT 2905.005 1626.070 2924.800 1626.075 ;
        RECT 2917.600 1625.620 2924.800 1626.070 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2882.775 1891.840 2883.295 1893.325 ;
      LAYER met1 ;
        RECT 2882.985 1891.965 2883.305 1892.225 ;
      LAYER met2 ;
        RECT 2883.025 1892.255 2883.305 1892.295 ;
        RECT 2883.015 1891.935 2883.305 1892.255 ;
        RECT 2883.025 1891.925 2883.305 1891.935 ;
      LAYER met3 ;
        RECT 2883.000 1892.265 2883.330 1892.275 ;
        RECT 2883.000 1892.250 2906.915 1892.265 ;
        RECT 2917.600 1892.250 2924.800 1892.700 ;
        RECT 2883.000 1891.955 2924.800 1892.250 ;
        RECT 2883.000 1891.945 2883.330 1891.955 ;
        RECT 2905.015 1891.950 2924.800 1891.955 ;
        RECT 2917.600 1891.500 2924.800 1891.950 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2882.775 2157.720 2883.295 2159.205 ;
      LAYER met1 ;
        RECT 2882.985 2157.845 2883.305 2158.105 ;
      LAYER met2 ;
        RECT 2883.025 2158.135 2883.305 2158.175 ;
        RECT 2883.015 2157.815 2883.305 2158.135 ;
        RECT 2883.025 2157.805 2883.305 2157.815 ;
      LAYER met3 ;
        RECT 2883.000 2158.145 2883.330 2158.155 ;
        RECT 2883.000 2158.130 2907.090 2158.145 ;
        RECT 2917.600 2158.130 2924.800 2158.580 ;
        RECT 2883.000 2157.835 2924.800 2158.130 ;
        RECT 2883.000 2157.825 2883.330 2157.835 ;
        RECT 2905.020 2157.830 2924.800 2157.835 ;
        RECT 2917.600 2157.380 2924.800 2157.830 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER li1 ;
        RECT 2727.695 2175.015 2727.865 2175.865 ;
        RECT 2728.535 2175.015 2728.705 2175.865 ;
        RECT 2729.375 2175.015 2729.545 2175.865 ;
        RECT 2730.215 2175.015 2730.385 2175.865 ;
        RECT 2731.055 2175.015 2731.225 2175.865 ;
        RECT 2731.895 2175.015 2732.065 2175.865 ;
        RECT 2727.695 2174.845 2732.065 2175.015 ;
        RECT 2730.130 2174.305 2732.065 2174.845 ;
        RECT 2727.695 2174.135 2732.065 2174.305 ;
        RECT 2727.695 2173.655 2727.865 2174.135 ;
        RECT 2728.535 2173.655 2728.705 2174.135 ;
        RECT 2729.375 2173.655 2729.545 2174.135 ;
        RECT 2730.215 2173.655 2730.385 2174.135 ;
        RECT 2731.055 2173.655 2731.225 2174.135 ;
        RECT 2731.895 2173.655 2732.065 2174.135 ;
      LAYER met1 ;
        RECT 2731.010 2174.120 2731.330 2174.380 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3499.125 2717.520 3517.600 ;
        RECT 2717.310 3498.755 2717.590 3499.125 ;
        RECT 2740.310 3498.755 2740.590 3499.125 ;
        RECT 2740.380 2177.205 2740.520 3498.755 ;
        RECT 2740.310 2176.835 2740.590 2177.205 ;
        RECT 2731.040 2174.090 2731.300 2174.410 ;
        RECT 2731.100 2172.565 2731.240 2174.090 ;
        RECT 2731.030 2172.195 2731.310 2172.565 ;
      LAYER met3 ;
        RECT 2717.285 3499.090 2717.615 3499.105 ;
        RECT 2740.285 3499.090 2740.615 3499.105 ;
        RECT 2717.285 3498.790 2740.615 3499.090 ;
        RECT 2717.285 3498.775 2717.615 3498.790 ;
        RECT 2740.285 3498.775 2740.615 3498.790 ;
        RECT 2740.285 2177.170 2740.615 2177.185 ;
        RECT 2739.150 2176.870 2740.615 2177.170 ;
        RECT 2739.150 2174.040 2739.450 2176.870 ;
        RECT 2740.285 2176.855 2740.615 2176.870 ;
        RECT 2736.000 2173.890 2740.000 2174.040 ;
        RECT 2735.390 2173.590 2740.000 2173.890 ;
        RECT 2731.005 2172.530 2731.335 2172.545 ;
        RECT 2735.390 2172.530 2735.690 2173.590 ;
        RECT 2736.000 2173.440 2740.000 2173.590 ;
        RECT 2731.005 2172.230 2735.690 2172.530 ;
        RECT 2731.005 2172.215 2731.335 2172.230 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER li1 ;
        RECT 2727.695 1995.015 2727.865 1995.865 ;
        RECT 2728.535 1995.015 2728.705 1995.865 ;
        RECT 2729.375 1995.015 2729.545 1995.865 ;
        RECT 2730.215 1995.015 2730.385 1995.865 ;
        RECT 2731.055 1995.015 2731.225 1995.865 ;
        RECT 2731.895 1995.015 2732.065 1995.865 ;
        RECT 2727.695 1994.845 2732.065 1995.015 ;
        RECT 2730.130 1994.305 2732.065 1994.845 ;
        RECT 2727.695 1994.135 2732.065 1994.305 ;
        RECT 2727.695 1993.655 2727.865 1994.135 ;
        RECT 2728.535 1993.655 2728.705 1994.135 ;
        RECT 2729.375 1993.655 2729.545 1994.135 ;
        RECT 2730.215 1993.655 2730.385 1994.135 ;
        RECT 2731.055 1993.655 2731.225 1994.135 ;
        RECT 2731.895 1993.655 2732.065 1994.135 ;
      LAYER met1 ;
        RECT 2731.010 1994.120 2731.330 1994.380 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3503.885 2392.760 3517.600 ;
        RECT 2392.550 3503.515 2392.830 3503.885 ;
        RECT 2739.850 3503.515 2740.130 3503.885 ;
        RECT 2731.040 1994.090 2731.300 1994.410 ;
        RECT 2731.100 1992.565 2731.240 1994.090 ;
        RECT 2739.920 1992.925 2740.060 3503.515 ;
        RECT 2731.030 1992.195 2731.310 1992.565 ;
        RECT 2739.850 1992.555 2740.130 1992.925 ;
      LAYER met3 ;
        RECT 2392.525 3503.850 2392.855 3503.865 ;
        RECT 2739.825 3503.850 2740.155 3503.865 ;
        RECT 2392.525 3503.550 2740.155 3503.850 ;
        RECT 2392.525 3503.535 2392.855 3503.550 ;
        RECT 2739.825 3503.535 2740.155 3503.550 ;
        RECT 2736.000 1993.890 2740.000 1994.040 ;
        RECT 2735.390 1993.590 2740.000 1993.890 ;
        RECT 2731.005 1992.530 2731.335 1992.545 ;
        RECT 2735.390 1992.530 2735.690 1993.590 ;
        RECT 2736.000 1993.440 2740.000 1993.590 ;
        RECT 2739.150 1992.890 2739.450 1993.440 ;
        RECT 2739.825 1992.890 2740.155 1992.905 ;
        RECT 2739.150 1992.590 2740.155 1992.890 ;
        RECT 2739.825 1992.575 2740.155 1992.590 ;
        RECT 2731.005 1992.230 2735.690 1992.530 ;
        RECT 2731.005 1992.215 2731.335 1992.230 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER li1 ;
        RECT 2727.695 1815.015 2727.865 1815.865 ;
        RECT 2728.535 1815.015 2728.705 1815.865 ;
        RECT 2729.375 1815.015 2729.545 1815.865 ;
        RECT 2730.215 1815.015 2730.385 1815.865 ;
        RECT 2731.055 1815.015 2731.225 1815.865 ;
        RECT 2731.895 1815.015 2732.065 1815.865 ;
        RECT 2727.695 1814.845 2732.065 1815.015 ;
        RECT 2730.130 1814.305 2732.065 1814.845 ;
        RECT 2727.695 1814.135 2732.065 1814.305 ;
        RECT 2727.695 1813.655 2727.865 1814.135 ;
        RECT 2728.535 1813.655 2728.705 1814.135 ;
        RECT 2729.375 1813.655 2729.545 1814.135 ;
        RECT 2730.215 1813.655 2730.385 1814.135 ;
        RECT 2731.055 1813.655 2731.225 1814.135 ;
        RECT 2731.895 1813.655 2732.065 1814.135 ;
      LAYER met1 ;
        RECT 2731.010 1814.120 2731.330 1814.380 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3503.205 2068.460 3517.600 ;
        RECT 2068.250 3502.835 2068.530 3503.205 ;
        RECT 2739.390 3502.835 2739.670 3503.205 ;
        RECT 2739.460 1814.765 2739.600 3502.835 ;
        RECT 2731.040 1814.090 2731.300 1814.410 ;
        RECT 2739.390 1814.395 2739.670 1814.765 ;
        RECT 2731.100 1812.565 2731.240 1814.090 ;
        RECT 2731.030 1812.195 2731.310 1812.565 ;
      LAYER met3 ;
        RECT 2068.225 3503.170 2068.555 3503.185 ;
        RECT 2739.365 3503.170 2739.695 3503.185 ;
        RECT 2068.225 3502.870 2739.695 3503.170 ;
        RECT 2068.225 3502.855 2068.555 3502.870 ;
        RECT 2739.365 3502.855 2739.695 3502.870 ;
        RECT 2739.365 1814.730 2739.695 1814.745 ;
        RECT 2739.150 1814.415 2739.695 1814.730 ;
        RECT 2739.150 1814.040 2739.450 1814.415 ;
        RECT 2736.000 1813.890 2740.000 1814.040 ;
        RECT 2735.390 1813.590 2740.000 1813.890 ;
        RECT 2731.005 1812.530 2731.335 1812.545 ;
        RECT 2735.390 1812.530 2735.690 1813.590 ;
        RECT 2736.000 1813.440 2740.000 1813.590 ;
        RECT 2731.005 1812.230 2735.690 1812.530 ;
        RECT 2731.005 1812.215 2731.335 1812.230 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER li1 ;
        RECT 2727.695 1635.015 2727.865 1635.865 ;
        RECT 2728.535 1635.015 2728.705 1635.865 ;
        RECT 2729.375 1635.015 2729.545 1635.865 ;
        RECT 2730.215 1635.015 2730.385 1635.865 ;
        RECT 2731.055 1635.015 2731.225 1635.865 ;
        RECT 2731.895 1635.015 2732.065 1635.865 ;
        RECT 2727.695 1634.845 2732.065 1635.015 ;
        RECT 2730.130 1634.305 2732.065 1634.845 ;
        RECT 2727.695 1634.135 2732.065 1634.305 ;
        RECT 2727.695 1633.655 2727.865 1634.135 ;
        RECT 2728.535 1633.655 2728.705 1634.135 ;
        RECT 2729.375 1633.655 2729.545 1634.135 ;
        RECT 2730.215 1633.655 2730.385 1634.135 ;
        RECT 2731.055 1633.655 2731.225 1634.135 ;
        RECT 2731.895 1633.655 2732.065 1634.135 ;
      LAYER met1 ;
        RECT 2731.010 1634.120 2731.330 1634.380 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3502.525 1744.160 3517.600 ;
        RECT 1743.950 3502.155 1744.230 3502.525 ;
        RECT 2737.090 3502.155 2737.370 3502.525 ;
        RECT 2737.160 1635.245 2737.300 3502.155 ;
        RECT 2737.090 1634.875 2737.370 1635.245 ;
        RECT 2731.040 1634.090 2731.300 1634.410 ;
        RECT 2731.100 1632.565 2731.240 1634.090 ;
        RECT 2731.030 1632.195 2731.310 1632.565 ;
      LAYER met3 ;
        RECT 1743.925 3502.490 1744.255 3502.505 ;
        RECT 2737.065 3502.490 2737.395 3502.505 ;
        RECT 1743.925 3502.190 2737.395 3502.490 ;
        RECT 1743.925 3502.175 1744.255 3502.190 ;
        RECT 2737.065 3502.175 2737.395 3502.190 ;
        RECT 2737.065 1635.210 2737.395 1635.225 ;
        RECT 2737.065 1634.895 2737.610 1635.210 ;
        RECT 2737.310 1634.040 2737.610 1634.895 ;
        RECT 2736.000 1633.890 2740.000 1634.040 ;
        RECT 2735.390 1633.590 2740.000 1633.890 ;
        RECT 2731.005 1632.530 2731.335 1632.545 ;
        RECT 2735.390 1632.530 2735.690 1633.590 ;
        RECT 2736.000 1633.440 2740.000 1633.590 ;
        RECT 2731.005 1632.230 2735.690 1632.530 ;
        RECT 2731.005 1632.215 2731.335 1632.230 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER li1 ;
        RECT 2727.695 1455.015 2727.865 1455.865 ;
        RECT 2728.535 1455.015 2728.705 1455.865 ;
        RECT 2729.375 1455.015 2729.545 1455.865 ;
        RECT 2730.215 1455.015 2730.385 1455.865 ;
        RECT 2731.055 1455.015 2731.225 1455.865 ;
        RECT 2731.895 1455.015 2732.065 1455.865 ;
        RECT 2727.695 1454.845 2732.065 1455.015 ;
        RECT 2730.130 1454.305 2732.065 1454.845 ;
        RECT 2727.695 1454.135 2732.065 1454.305 ;
        RECT 2727.695 1453.655 2727.865 1454.135 ;
        RECT 2728.535 1453.655 2728.705 1454.135 ;
        RECT 2729.375 1453.655 2729.545 1454.135 ;
        RECT 2730.215 1453.655 2730.385 1454.135 ;
        RECT 2731.055 1453.655 2731.225 1454.135 ;
        RECT 2731.895 1453.655 2732.065 1454.135 ;
      LAYER met1 ;
        RECT 2731.010 1454.120 2731.330 1454.380 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3501.845 1419.400 3517.600 ;
        RECT 1419.190 3501.475 1419.470 3501.845 ;
        RECT 2736.630 3501.475 2736.910 3501.845 ;
        RECT 2736.700 1455.725 2736.840 3501.475 ;
        RECT 2736.630 1455.355 2736.910 1455.725 ;
        RECT 2731.040 1454.090 2731.300 1454.410 ;
        RECT 2731.100 1452.565 2731.240 1454.090 ;
        RECT 2731.030 1452.195 2731.310 1452.565 ;
      LAYER met3 ;
        RECT 1419.165 3501.810 1419.495 3501.825 ;
        RECT 2736.605 3501.810 2736.935 3501.825 ;
        RECT 1419.165 3501.510 2736.935 3501.810 ;
        RECT 1419.165 3501.495 1419.495 3501.510 ;
        RECT 2736.605 3501.495 2736.935 3501.510 ;
        RECT 2736.605 1455.690 2736.935 1455.705 ;
        RECT 2736.390 1455.375 2736.935 1455.690 ;
        RECT 2736.390 1454.040 2736.690 1455.375 ;
        RECT 2736.000 1453.890 2740.000 1454.040 ;
        RECT 2735.390 1453.590 2740.000 1453.890 ;
        RECT 2731.005 1452.530 2731.335 1452.545 ;
        RECT 2735.390 1452.530 2735.690 1453.590 ;
        RECT 2736.000 1453.440 2740.000 1453.590 ;
        RECT 2731.005 1452.230 2735.690 1452.530 ;
        RECT 2731.005 1452.215 2731.335 1452.230 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1262.215 3508.915 1264.410 3511.090 ;
        RECT 1622.215 3509.365 1624.410 3511.540 ;
        RECT 1802.215 3507.445 1804.410 3509.620 ;
        RECT 2162.215 3507.085 2164.410 3509.260 ;
        RECT 2522.215 3507.770 2524.410 3509.945 ;
        RECT 2881.390 3486.805 2883.585 3488.980 ;
        RECT 2881.390 3220.925 2883.585 3223.100 ;
        RECT 2881.390 2955.725 2883.585 2957.900 ;
        RECT 2881.390 2689.845 2883.585 2692.020 ;
        RECT 2881.390 2423.965 2883.585 2426.140 ;
        RECT 2360.765 2253.735 2364.310 2253.740 ;
        RECT 2357.985 2253.130 2364.310 2253.735 ;
        RECT 2371.535 2253.130 2380.895 2253.740 ;
        RECT 2388.120 2253.130 2397.480 2253.740 ;
        RECT 2404.705 2253.130 2414.065 2253.740 ;
        RECT 2421.290 2253.130 2430.645 2253.740 ;
        RECT 2357.985 2252.620 2364.330 2253.130 ;
        RECT 2357.995 2252.135 2364.330 2252.620 ;
        RECT 2371.535 2252.135 2380.915 2253.130 ;
        RECT 2388.120 2252.135 2397.500 2253.130 ;
        RECT 2404.705 2252.135 2414.085 2253.130 ;
        RECT 2421.290 2252.135 2430.665 2253.130 ;
        RECT 2437.870 2252.135 2443.725 2253.740 ;
        RECT 2357.995 2250.425 2443.725 2252.135 ;
        RECT 2357.985 2249.305 2443.725 2250.425 ;
        RECT 2357.985 2248.715 2364.005 2249.305 ;
        RECT 2371.695 2248.720 2380.590 2249.305 ;
        RECT 2388.280 2248.720 2397.175 2249.305 ;
        RECT 2404.865 2248.720 2413.760 2249.305 ;
        RECT 2421.450 2248.720 2430.340 2249.305 ;
        RECT 2438.030 2248.720 2443.725 2249.305 ;
        RECT 2377.240 2248.715 2380.590 2248.720 ;
        RECT 2393.810 2248.715 2397.175 2248.720 ;
        RECT 2410.405 2248.715 2413.760 2248.720 ;
        RECT 2426.960 2248.715 2430.340 2248.720 ;
        RECT 2360.800 2248.710 2363.775 2248.715 ;
        RECT 2377.385 2248.710 2380.360 2248.715 ;
        RECT 2393.810 2248.710 2396.945 2248.715 ;
        RECT 2410.405 2248.710 2413.530 2248.715 ;
        RECT 2426.960 2248.710 2430.110 2248.715 ;
        RECT 2695.330 2212.785 2734.350 2215.615 ;
        RECT 2695.330 2207.345 2734.350 2210.175 ;
        RECT 2695.330 2201.905 2734.350 2204.735 ;
        RECT 2695.330 2196.465 2734.350 2199.295 ;
        RECT 2695.330 2191.025 2734.350 2193.855 ;
        RECT 2695.330 2185.585 2734.350 2188.415 ;
        RECT 2695.330 2180.145 2734.350 2182.975 ;
        RECT 2695.330 2174.705 2734.350 2177.535 ;
        RECT 2695.330 2169.265 2734.350 2172.095 ;
        RECT 2695.330 2163.825 2734.350 2166.655 ;
        RECT 2358.015 2161.745 2359.010 2162.015 ;
        RECT 2358.015 2161.740 2361.495 2161.745 ;
        RECT 2373.115 2161.740 2378.680 2161.745 ;
        RECT 2390.335 2161.740 2396.030 2161.745 ;
        RECT 2407.555 2161.740 2413.105 2161.745 ;
        RECT 2424.775 2161.740 2430.320 2161.745 ;
        RECT 2441.995 2161.740 2446.775 2161.745 ;
        RECT 2358.015 2160.145 2364.410 2161.740 ;
        RECT 2372.350 2161.130 2381.465 2161.740 ;
        RECT 2389.570 2161.130 2398.685 2161.740 ;
        RECT 2406.790 2161.130 2415.905 2161.740 ;
        RECT 2424.010 2161.130 2433.125 2161.740 ;
        RECT 2441.230 2161.130 2446.925 2161.740 ;
        RECT 2372.155 2160.145 2381.465 2161.130 ;
        RECT 2389.375 2160.145 2398.685 2161.130 ;
        RECT 2406.595 2160.145 2415.905 2161.130 ;
        RECT 2423.815 2160.145 2433.125 2161.130 ;
        RECT 2358.015 2160.140 2364.455 2160.145 ;
        RECT 2372.155 2160.140 2381.675 2160.145 ;
        RECT 2389.375 2160.140 2398.895 2160.145 ;
        RECT 2406.595 2160.140 2416.115 2160.145 ;
        RECT 2423.815 2160.140 2433.335 2160.145 ;
        RECT 2441.035 2160.140 2446.925 2161.130 ;
        RECT 2358.015 2157.310 2446.925 2160.140 ;
        RECT 2695.330 2158.385 2734.350 2161.215 ;
        RECT 2881.390 2158.765 2883.585 2160.940 ;
        RECT 2358.015 2156.710 2364.410 2157.310 ;
        RECT 2372.350 2156.720 2381.630 2157.310 ;
        RECT 2389.570 2156.720 2398.850 2157.310 ;
        RECT 2406.790 2156.720 2416.070 2157.310 ;
        RECT 2424.010 2156.720 2433.290 2157.310 ;
        RECT 2441.230 2156.720 2446.925 2157.310 ;
        RECT 2373.115 2156.715 2381.630 2156.720 ;
        RECT 2390.335 2156.715 2398.850 2156.720 ;
        RECT 2407.555 2156.715 2416.070 2156.720 ;
        RECT 2424.775 2156.715 2433.290 2156.720 ;
        RECT 2441.995 2156.715 2446.770 2156.720 ;
        RECT 2378.035 2156.710 2381.630 2156.715 ;
        RECT 2395.255 2156.710 2398.850 2156.715 ;
        RECT 2412.475 2156.710 2416.070 2156.715 ;
        RECT 2429.695 2156.710 2433.290 2156.715 ;
        RECT 2695.330 2152.945 2734.350 2155.775 ;
        RECT 2695.330 2147.505 2734.350 2150.335 ;
        RECT 2695.330 2142.065 2734.350 2144.895 ;
        RECT 2521.945 2135.255 2524.140 2137.430 ;
        RECT 2695.330 2136.625 2734.350 2139.455 ;
        RECT 2695.330 2131.185 2734.350 2134.015 ;
        RECT 2521.945 2127.725 2524.140 2129.900 ;
        RECT 2521.945 2121.745 2524.140 2123.920 ;
        RECT 2521.945 2115.800 2524.140 2117.975 ;
        RECT 2521.945 2110.155 2524.140 2112.330 ;
        RECT 2521.945 2104.150 2524.140 2106.325 ;
        RECT 2358.000 2056.740 2360.810 2056.745 ;
        RECT 2366.580 2056.740 2369.390 2056.745 ;
        RECT 2372.195 2056.740 2375.985 2056.745 ;
        RECT 2382.905 2056.740 2385.715 2056.745 ;
        RECT 2388.520 2056.740 2392.310 2056.745 ;
        RECT 2399.230 2056.740 2402.040 2056.745 ;
        RECT 2404.845 2056.740 2408.635 2056.745 ;
        RECT 2415.555 2056.740 2418.365 2056.745 ;
        RECT 2421.170 2056.740 2424.960 2056.745 ;
        RECT 2431.880 2056.740 2434.690 2056.745 ;
        RECT 2437.495 2056.740 2441.285 2056.745 ;
        RECT 2358.000 2052.100 2442.425 2056.740 ;
        RECT 2360.790 2052.095 2442.425 2052.100 ;
        RECT 2371.175 2052.020 2377.125 2052.095 ;
        RECT 2387.500 2052.020 2393.450 2052.095 ;
        RECT 2403.825 2052.020 2409.775 2052.095 ;
        RECT 2420.150 2052.020 2426.100 2052.095 ;
        RECT 2436.475 2052.020 2442.425 2052.095 ;
        RECT 2371.180 2051.720 2377.125 2052.020 ;
        RECT 2387.505 2051.720 2393.450 2052.020 ;
        RECT 2403.830 2051.720 2409.775 2052.020 ;
        RECT 2420.155 2051.720 2426.100 2052.020 ;
        RECT 2436.480 2051.720 2442.425 2052.020 ;
        RECT 2372.195 2051.715 2375.985 2051.720 ;
        RECT 2388.520 2051.715 2392.310 2051.720 ;
        RECT 2404.845 2051.715 2408.635 2051.720 ;
        RECT 2421.170 2051.715 2424.960 2051.720 ;
        RECT 2437.495 2051.715 2441.285 2051.720 ;
        RECT 2695.330 2032.785 2734.350 2035.615 ;
        RECT 2695.330 2027.345 2734.350 2030.175 ;
        RECT 2695.330 2021.905 2734.350 2024.735 ;
        RECT 2695.330 2016.465 2734.350 2019.295 ;
        RECT 2695.330 2011.025 2734.350 2013.855 ;
        RECT 2695.330 2005.585 2734.350 2008.415 ;
        RECT 2695.330 2000.145 2734.350 2002.975 ;
        RECT 2695.330 1994.705 2734.350 1997.535 ;
        RECT 2695.330 1989.265 2734.350 1992.095 ;
        RECT 2521.945 1983.000 2524.140 1985.175 ;
        RECT 2695.330 1983.825 2734.350 1986.655 ;
        RECT 2695.330 1978.385 2734.350 1981.215 ;
        RECT 2521.945 1975.470 2524.140 1977.645 ;
        RECT 2695.330 1972.945 2734.350 1975.775 ;
        RECT 2521.945 1969.490 2524.140 1971.665 ;
        RECT 2695.330 1967.505 2734.350 1970.335 ;
        RECT 2521.945 1963.545 2524.140 1965.720 ;
        RECT 2695.330 1962.065 2734.350 1964.895 ;
        RECT 2521.945 1957.900 2524.140 1960.075 ;
        RECT 2695.330 1956.625 2734.350 1959.455 ;
        RECT 2521.945 1951.895 2524.140 1954.070 ;
        RECT 2358.000 1951.745 2363.165 1951.750 ;
        RECT 2368.815 1951.745 2371.625 1951.750 ;
        RECT 2374.430 1951.745 2377.240 1951.750 ;
        RECT 2379.360 1951.745 2381.725 1951.750 ;
        RECT 2387.375 1951.745 2390.185 1951.750 ;
        RECT 2392.990 1951.745 2395.800 1951.750 ;
        RECT 2397.920 1951.745 2400.285 1951.750 ;
        RECT 2405.935 1951.745 2408.745 1951.750 ;
        RECT 2411.550 1951.745 2414.360 1951.750 ;
        RECT 2416.480 1951.745 2418.845 1951.750 ;
        RECT 2424.495 1951.745 2427.305 1951.750 ;
        RECT 2430.110 1951.745 2432.920 1951.750 ;
        RECT 2435.040 1951.745 2437.405 1951.750 ;
        RECT 2443.055 1951.745 2445.865 1951.750 ;
        RECT 2448.670 1951.745 2451.480 1951.750 ;
        RECT 2358.000 1948.450 2453.600 1951.745 ;
        RECT 2695.330 1951.185 2734.350 1954.015 ;
        RECT 2358.005 1948.095 2453.600 1948.450 ;
        RECT 2360.800 1947.100 2453.600 1948.095 ;
        RECT 2361.305 1947.095 2453.600 1947.100 ;
        RECT 2373.410 1946.720 2379.360 1947.095 ;
        RECT 2391.970 1946.720 2397.920 1947.095 ;
        RECT 2410.530 1947.090 2417.800 1947.095 ;
        RECT 2410.530 1946.720 2416.480 1947.090 ;
        RECT 2429.090 1946.720 2435.040 1947.095 ;
        RECT 2447.650 1946.720 2453.600 1947.095 ;
        RECT 2374.430 1946.715 2377.240 1946.720 ;
        RECT 2392.990 1946.715 2395.800 1946.720 ;
        RECT 2411.550 1946.715 2414.360 1946.720 ;
        RECT 2430.110 1946.715 2432.920 1946.720 ;
        RECT 2448.670 1946.715 2451.480 1946.720 ;
        RECT 2881.390 1892.885 2883.585 1895.060 ;
        RECT 2695.330 1852.785 2734.350 1855.615 ;
        RECT 2695.330 1847.345 2734.350 1850.175 ;
        RECT 2695.330 1841.905 2734.350 1844.735 ;
        RECT 2695.330 1836.465 2734.350 1839.295 ;
        RECT 2695.330 1831.025 2734.350 1833.855 ;
        RECT 2695.330 1825.585 2734.350 1828.415 ;
        RECT 2695.330 1820.145 2734.350 1822.975 ;
        RECT 2695.330 1814.705 2734.350 1817.535 ;
        RECT 2695.330 1809.265 2734.350 1812.095 ;
        RECT 2521.945 1806.030 2524.140 1808.205 ;
        RECT 2695.330 1803.825 2734.350 1806.655 ;
        RECT 2521.945 1798.500 2524.140 1800.675 ;
        RECT 2695.330 1798.385 2734.350 1801.215 ;
        RECT 2521.945 1792.520 2524.140 1794.695 ;
        RECT 2695.330 1792.945 2734.350 1795.775 ;
        RECT 2367.945 1788.745 2370.755 1788.750 ;
        RECT 2375.460 1788.745 2378.270 1788.750 ;
        RECT 2381.075 1788.745 2385.855 1788.750 ;
        RECT 2390.720 1788.745 2393.530 1788.750 ;
        RECT 2396.335 1788.745 2401.115 1788.750 ;
        RECT 2405.980 1788.745 2408.790 1788.750 ;
        RECT 2411.595 1788.745 2416.375 1788.750 ;
        RECT 2421.240 1788.745 2424.050 1788.750 ;
        RECT 2426.855 1788.745 2431.635 1788.750 ;
        RECT 2436.500 1788.745 2439.310 1788.750 ;
        RECT 2442.115 1788.745 2446.895 1788.750 ;
        RECT 2367.945 1786.660 2447.045 1788.745 ;
        RECT 2367.980 1784.100 2447.045 1786.660 ;
        RECT 2521.945 1786.575 2524.140 1788.750 ;
        RECT 2695.330 1787.505 2734.350 1790.335 ;
        RECT 2370.745 1784.095 2447.045 1784.100 ;
        RECT 2380.055 1783.720 2386.005 1784.095 ;
        RECT 2395.315 1783.720 2401.265 1784.095 ;
        RECT 2410.575 1783.720 2416.525 1784.095 ;
        RECT 2425.835 1783.720 2431.785 1784.095 ;
        RECT 2441.095 1783.720 2447.045 1784.095 ;
        RECT 2381.075 1783.715 2385.850 1783.720 ;
        RECT 2396.335 1783.715 2401.110 1783.720 ;
        RECT 2411.595 1783.715 2416.370 1783.720 ;
        RECT 2426.855 1783.715 2431.630 1783.720 ;
        RECT 2442.115 1783.715 2446.890 1783.720 ;
        RECT 2521.945 1780.930 2524.140 1783.105 ;
        RECT 2695.330 1782.065 2734.350 1784.895 ;
        RECT 2695.330 1776.625 2734.350 1779.455 ;
        RECT 2521.945 1769.460 2524.140 1771.635 ;
        RECT 2695.330 1771.185 2734.350 1774.015 ;
        RECT 2410.750 1708.745 2414.425 1708.750 ;
        RECT 2394.180 1708.740 2397.840 1708.745 ;
        RECT 2358.205 1708.130 2364.670 1708.740 ;
        RECT 2371.895 1708.130 2381.255 1708.740 ;
        RECT 2388.480 1708.135 2397.840 1708.740 ;
        RECT 2405.065 1708.140 2414.425 1708.745 ;
        RECT 2421.650 1708.140 2431.005 1708.750 ;
        RECT 2358.205 1707.135 2364.690 1708.130 ;
        RECT 2371.895 1707.135 2381.275 1708.130 ;
        RECT 2388.480 1707.140 2397.860 1708.135 ;
        RECT 2405.065 1707.145 2414.445 1708.140 ;
        RECT 2421.650 1707.145 2431.025 1708.140 ;
        RECT 2438.230 1707.145 2444.085 1708.750 ;
        RECT 2405.065 1707.140 2444.085 1707.145 ;
        RECT 2388.480 1707.135 2444.085 1707.140 ;
        RECT 2358.205 1704.705 2444.085 1707.135 ;
        RECT 2358.210 1704.315 2444.085 1704.705 ;
        RECT 2358.210 1704.310 2414.115 1704.315 ;
        RECT 2358.210 1704.305 2397.530 1704.310 ;
        RECT 2358.210 1704.225 2364.670 1704.305 ;
        RECT 2358.210 1703.715 2364.360 1704.225 ;
        RECT 2372.055 1703.720 2380.945 1704.305 ;
        RECT 2388.640 1703.720 2397.530 1704.305 ;
        RECT 2405.225 1703.725 2414.115 1704.310 ;
        RECT 2421.810 1703.730 2430.695 1704.315 ;
        RECT 2438.390 1703.730 2444.085 1704.315 ;
        RECT 2410.915 1703.720 2414.115 1703.725 ;
        RECT 2427.495 1703.720 2430.695 1703.730 ;
        RECT 2361.160 1703.710 2364.360 1703.715 ;
        RECT 2377.745 1703.710 2380.945 1703.720 ;
        RECT 2394.330 1703.715 2397.530 1703.720 ;
        RECT 2695.330 1672.785 2734.350 1675.615 ;
        RECT 2695.330 1667.345 2734.350 1670.175 ;
        RECT 2695.330 1661.905 2734.350 1664.735 ;
        RECT 2695.330 1656.465 2734.350 1659.295 ;
        RECT 2695.330 1651.025 2734.350 1653.855 ;
        RECT 2695.330 1645.585 2734.350 1648.415 ;
        RECT 2695.330 1640.145 2734.350 1642.975 ;
        RECT 2695.330 1634.705 2734.350 1637.535 ;
        RECT 2695.330 1629.265 2734.350 1632.095 ;
        RECT 2521.945 1624.895 2524.140 1627.070 ;
        RECT 2881.390 1627.005 2883.585 1629.180 ;
        RECT 2695.330 1623.825 2734.350 1626.655 ;
        RECT 2521.945 1618.480 2524.140 1620.655 ;
        RECT 2695.330 1618.385 2734.350 1621.215 ;
        RECT 2695.330 1612.945 2734.350 1615.775 ;
        RECT 2395.845 1608.745 2398.655 1608.750 ;
        RECT 2407.530 1608.745 2412.310 1608.750 ;
        RECT 2357.995 1608.740 2364.215 1608.745 ;
        RECT 2373.090 1608.740 2381.435 1608.745 ;
        RECT 2390.310 1608.740 2398.800 1608.745 ;
        RECT 2357.995 1607.140 2364.385 1608.740 ;
        RECT 2372.325 1608.130 2381.580 1608.740 ;
        RECT 2389.545 1608.130 2398.800 1608.740 ;
        RECT 2406.765 1608.740 2415.875 1608.745 ;
        RECT 2424.750 1608.740 2433.095 1608.745 ;
        RECT 2441.970 1608.740 2446.750 1608.745 ;
        RECT 2406.765 1608.135 2416.020 1608.740 ;
        RECT 2372.130 1607.140 2381.580 1608.130 ;
        RECT 2389.350 1607.145 2398.800 1608.130 ;
        RECT 2406.570 1607.145 2416.020 1608.135 ;
        RECT 2423.985 1608.130 2433.240 1608.740 ;
        RECT 2441.205 1608.130 2446.900 1608.740 ;
        RECT 2389.350 1607.140 2416.020 1607.145 ;
        RECT 2423.790 1607.140 2433.240 1608.130 ;
        RECT 2441.010 1607.140 2446.900 1608.130 ;
        RECT 2695.330 1607.505 2734.350 1610.335 ;
        RECT 2357.995 1606.655 2446.900 1607.140 ;
        RECT 2358.000 1604.775 2446.900 1606.655 ;
        RECT 2357.995 1604.315 2446.900 1604.775 ;
        RECT 2357.995 1604.310 2398.825 1604.315 ;
        RECT 2357.995 1603.710 2364.385 1604.310 ;
        RECT 2372.325 1603.720 2381.605 1604.310 ;
        RECT 2389.545 1603.720 2398.825 1604.310 ;
        RECT 2406.765 1604.310 2446.900 1604.315 ;
        RECT 2406.765 1603.725 2416.045 1604.310 ;
        RECT 2407.530 1603.720 2416.045 1603.725 ;
        RECT 2423.985 1603.720 2433.265 1604.310 ;
        RECT 2441.205 1603.720 2446.900 1604.310 ;
        RECT 2373.090 1603.715 2381.605 1603.720 ;
        RECT 2390.310 1603.715 2398.825 1603.720 ;
        RECT 2378.010 1603.710 2381.605 1603.715 ;
        RECT 2412.300 1603.710 2416.045 1603.720 ;
        RECT 2424.750 1603.715 2433.265 1603.720 ;
        RECT 2441.970 1603.715 2446.745 1603.720 ;
        RECT 2429.525 1603.710 2433.265 1603.715 ;
        RECT 2695.330 1602.065 2734.350 1604.895 ;
        RECT 2695.330 1596.625 2734.350 1599.455 ;
        RECT 2521.945 1589.235 2524.140 1591.410 ;
        RECT 2695.330 1591.185 2734.350 1594.015 ;
        RECT 2521.945 1581.705 2524.140 1583.880 ;
        RECT 2521.945 1575.725 2524.140 1577.900 ;
        RECT 2521.945 1567.310 2524.140 1569.485 ;
        RECT 2357.995 1531.740 2360.805 1531.745 ;
        RECT 2366.575 1531.740 2369.385 1531.745 ;
        RECT 2372.190 1531.740 2375.980 1531.745 ;
        RECT 2382.900 1531.740 2385.710 1531.745 ;
        RECT 2388.515 1531.740 2392.305 1531.745 ;
        RECT 2399.225 1531.740 2402.035 1531.745 ;
        RECT 2404.840 1531.740 2408.630 1531.745 ;
        RECT 2415.550 1531.740 2418.360 1531.745 ;
        RECT 2421.165 1531.740 2424.955 1531.745 ;
        RECT 2431.875 1531.740 2434.685 1531.745 ;
        RECT 2437.490 1531.740 2441.280 1531.745 ;
        RECT 2357.995 1529.655 2442.420 1531.740 ;
        RECT 2358.000 1527.000 2442.420 1529.655 ;
        RECT 2360.785 1526.985 2442.420 1527.000 ;
        RECT 2371.175 1526.720 2377.120 1526.985 ;
        RECT 2387.500 1526.720 2393.445 1526.985 ;
        RECT 2403.825 1526.720 2409.770 1526.985 ;
        RECT 2420.150 1526.720 2426.095 1526.985 ;
        RECT 2436.475 1526.720 2442.420 1526.985 ;
        RECT 2372.190 1526.715 2375.980 1526.720 ;
        RECT 2388.515 1526.715 2392.305 1526.720 ;
        RECT 2404.840 1526.715 2408.630 1526.720 ;
        RECT 2421.165 1526.715 2424.955 1526.720 ;
        RECT 2437.490 1526.715 2441.280 1526.720 ;
        RECT 2695.330 1492.785 2734.350 1495.615 ;
        RECT 2695.330 1487.345 2734.350 1490.175 ;
        RECT 2695.330 1481.905 2734.350 1484.735 ;
        RECT 2695.330 1476.465 2734.350 1479.295 ;
        RECT 2695.330 1471.025 2734.350 1473.855 ;
        RECT 2695.330 1465.585 2734.350 1468.415 ;
        RECT 2695.330 1460.145 2734.350 1462.975 ;
        RECT 2695.330 1454.705 2734.350 1457.535 ;
        RECT 2695.330 1449.265 2734.350 1452.095 ;
        RECT 2695.330 1443.825 2734.350 1446.655 ;
        RECT 2521.945 1437.610 2524.140 1439.785 ;
        RECT 2695.330 1438.385 2734.350 1441.215 ;
        RECT 2377.545 1433.750 2379.580 1433.755 ;
        RECT 2357.995 1433.745 2363.160 1433.750 ;
        RECT 2368.810 1433.745 2371.620 1433.750 ;
        RECT 2374.425 1433.745 2381.720 1433.750 ;
        RECT 2387.370 1433.745 2390.180 1433.750 ;
        RECT 2392.985 1433.745 2400.280 1433.750 ;
        RECT 2405.930 1433.745 2408.740 1433.750 ;
        RECT 2411.545 1433.745 2418.840 1433.750 ;
        RECT 2424.490 1433.745 2427.300 1433.750 ;
        RECT 2430.105 1433.745 2437.400 1433.750 ;
        RECT 2443.050 1433.745 2445.860 1433.750 ;
        RECT 2448.665 1433.745 2452.455 1433.750 ;
        RECT 2357.995 1431.660 2453.595 1433.745 ;
        RECT 2358.000 1429.100 2453.595 1431.660 ;
        RECT 2521.945 1431.195 2524.140 1433.370 ;
        RECT 2695.330 1432.945 2734.350 1435.775 ;
        RECT 2361.300 1429.095 2453.595 1429.100 ;
        RECT 2373.405 1428.720 2379.355 1429.095 ;
        RECT 2391.965 1428.720 2397.915 1429.095 ;
        RECT 2410.525 1428.720 2416.475 1429.095 ;
        RECT 2429.085 1428.720 2435.035 1429.095 ;
        RECT 2447.645 1428.720 2453.595 1429.095 ;
        RECT 2374.425 1428.715 2378.215 1428.720 ;
        RECT 2392.985 1428.715 2396.775 1428.720 ;
        RECT 2411.545 1428.715 2415.335 1428.720 ;
        RECT 2430.105 1428.715 2433.895 1428.720 ;
        RECT 2448.665 1428.715 2452.455 1428.720 ;
        RECT 2695.330 1427.505 2734.350 1430.335 ;
        RECT 2695.330 1422.065 2734.350 1424.895 ;
        RECT 2521.945 1417.005 2524.140 1419.180 ;
        RECT 2695.330 1416.625 2734.350 1419.455 ;
        RECT 2521.945 1409.475 2524.140 1411.650 ;
        RECT 2695.330 1411.185 2734.350 1414.015 ;
        RECT 2521.945 1403.495 2524.140 1405.670 ;
        RECT 2521.945 1395.080 2524.140 1397.255 ;
        RECT 2881.390 1361.805 2883.585 1363.980 ;
        RECT 2367.995 1333.745 2370.805 1333.750 ;
        RECT 2375.510 1333.745 2378.320 1333.750 ;
        RECT 2381.125 1333.745 2385.905 1333.750 ;
        RECT 2390.770 1333.745 2393.580 1333.750 ;
        RECT 2396.385 1333.745 2401.165 1333.750 ;
        RECT 2406.030 1333.745 2408.840 1333.750 ;
        RECT 2411.645 1333.745 2416.425 1333.750 ;
        RECT 2421.290 1333.745 2424.100 1333.750 ;
        RECT 2426.905 1333.745 2431.685 1333.750 ;
        RECT 2436.550 1333.745 2439.360 1333.750 ;
        RECT 2442.165 1333.745 2446.945 1333.750 ;
        RECT 2367.995 1331.660 2447.095 1333.745 ;
        RECT 2368.000 1330.095 2447.095 1331.660 ;
        RECT 2368.010 1329.100 2447.095 1330.095 ;
        RECT 2370.795 1329.095 2447.095 1329.100 ;
        RECT 2380.105 1328.720 2386.055 1329.095 ;
        RECT 2395.365 1328.720 2401.315 1329.095 ;
        RECT 2410.625 1328.720 2416.575 1329.095 ;
        RECT 2425.885 1328.720 2431.835 1329.095 ;
        RECT 2441.145 1328.720 2447.095 1329.095 ;
        RECT 2381.125 1328.715 2385.900 1328.720 ;
        RECT 2396.385 1328.715 2401.160 1328.720 ;
        RECT 2411.645 1328.715 2416.420 1328.720 ;
        RECT 2426.905 1328.715 2431.680 1328.720 ;
        RECT 2442.165 1328.715 2446.940 1328.720 ;
        RECT 2881.390 1162.565 2883.585 1164.740 ;
      LAYER li1 ;
        RECT 1263.080 3509.755 1263.410 3510.480 ;
        RECT 1623.080 3510.205 1623.410 3510.930 ;
        RECT 1622.405 3510.035 1624.185 3510.205 ;
        RECT 1262.405 3509.585 1264.185 3509.755 ;
        RECT 1803.080 3508.285 1803.410 3509.010 ;
        RECT 1802.405 3508.115 1804.185 3508.285 ;
        RECT 2163.080 3507.925 2163.410 3508.650 ;
        RECT 2523.080 3508.610 2523.410 3509.335 ;
        RECT 2522.405 3508.440 2524.185 3508.610 ;
        RECT 2162.405 3507.755 2164.185 3507.925 ;
        RECT 2881.580 3488.140 2883.380 3488.310 ;
        RECT 2882.775 3487.415 2883.105 3488.140 ;
        RECT 2881.580 3222.260 2883.380 3222.430 ;
        RECT 2882.775 3221.535 2883.105 3222.260 ;
        RECT 2881.580 2957.060 2883.380 2957.230 ;
        RECT 2882.775 2956.335 2883.105 2957.060 ;
        RECT 2881.580 2691.180 2883.380 2691.350 ;
        RECT 2882.775 2690.455 2883.105 2691.180 ;
        RECT 2881.580 2425.300 2883.380 2425.470 ;
        RECT 2882.775 2424.575 2883.105 2425.300 ;
        RECT 2360.040 2255.035 2360.215 2255.585 ;
        RECT 2360.040 2253.435 2360.210 2255.035 ;
        RECT 2358.225 2252.025 2358.395 2252.755 ;
        RECT 2360.040 2252.295 2360.215 2253.435 ;
        RECT 2360.040 2252.025 2360.210 2252.295 ;
        RECT 2361.455 2252.025 2361.625 2252.755 ;
        RECT 2372.680 2252.030 2372.850 2252.760 ;
        RECT 2375.425 2252.030 2375.595 2252.760 ;
        RECT 2376.415 2252.030 2376.585 2252.760 ;
        RECT 2378.040 2252.030 2378.210 2252.755 ;
        RECT 2389.265 2252.030 2389.435 2252.760 ;
        RECT 2392.010 2252.030 2392.180 2252.760 ;
        RECT 2393.000 2252.030 2393.170 2252.760 ;
        RECT 2394.625 2252.030 2394.795 2252.755 ;
        RECT 2405.850 2252.030 2406.020 2252.760 ;
        RECT 2408.595 2252.030 2408.765 2252.760 ;
        RECT 2409.585 2252.030 2409.755 2252.760 ;
        RECT 2411.210 2252.030 2411.380 2252.755 ;
        RECT 2422.435 2252.030 2422.605 2252.760 ;
        RECT 2425.180 2252.030 2425.350 2252.760 ;
        RECT 2426.170 2252.030 2426.340 2252.760 ;
        RECT 2427.790 2252.030 2427.960 2252.755 ;
        RECT 2439.015 2252.030 2439.185 2252.760 ;
        RECT 2441.760 2252.030 2441.930 2252.760 ;
        RECT 2442.750 2252.030 2442.920 2252.760 ;
        RECT 2343.000 2250.805 2364.620 2252.025 ;
        RECT 2365.710 2250.805 2366.040 2251.525 ;
        RECT 2366.725 2250.805 2367.005 2251.265 ;
        RECT 2367.870 2250.805 2368.140 2251.585 ;
        RECT 2368.690 2250.805 2369.060 2251.185 ;
        RECT 2371.450 2250.965 2381.205 2252.030 ;
        RECT 2371.320 2250.805 2381.205 2250.965 ;
        RECT 2382.295 2250.805 2382.625 2251.525 ;
        RECT 2383.310 2250.805 2383.590 2251.265 ;
        RECT 2384.455 2250.805 2384.725 2251.585 ;
        RECT 2385.275 2250.805 2385.645 2251.185 ;
        RECT 2388.035 2250.965 2397.790 2252.030 ;
        RECT 2387.905 2250.805 2397.790 2250.965 ;
        RECT 2398.880 2250.805 2399.210 2251.525 ;
        RECT 2399.895 2250.805 2400.175 2251.265 ;
        RECT 2401.040 2250.805 2401.310 2251.585 ;
        RECT 2401.860 2250.805 2402.230 2251.185 ;
        RECT 2404.620 2250.965 2414.375 2252.030 ;
        RECT 2404.490 2250.805 2414.375 2250.965 ;
        RECT 2415.465 2250.805 2415.795 2251.525 ;
        RECT 2416.480 2250.805 2416.760 2251.265 ;
        RECT 2417.625 2250.805 2417.895 2251.585 ;
        RECT 2418.445 2250.805 2418.815 2251.185 ;
        RECT 2421.205 2250.965 2430.960 2252.030 ;
        RECT 2421.075 2250.805 2430.960 2250.965 ;
        RECT 2432.045 2250.805 2432.375 2251.525 ;
        RECT 2433.060 2250.805 2433.340 2251.265 ;
        RECT 2434.205 2250.805 2434.475 2251.585 ;
        RECT 2435.025 2250.805 2435.395 2251.185 ;
        RECT 2437.785 2250.965 2443.725 2252.030 ;
        RECT 2437.655 2250.805 2443.725 2250.965 ;
        RECT 2343.000 2250.635 2443.725 2250.805 ;
        RECT 2343.000 2250.425 2364.620 2250.635 ;
        RECT 2364.295 2250.125 2364.555 2250.425 ;
        RECT 2365.520 2250.135 2366.140 2250.635 ;
        RECT 2365.940 2249.955 2366.140 2250.135 ;
        RECT 2366.950 2250.095 2367.170 2250.635 ;
        RECT 2367.820 2249.985 2368.430 2250.635 ;
        RECT 2369.250 2250.095 2369.510 2250.635 ;
        RECT 2370.990 2250.430 2381.205 2250.635 ;
        RECT 2368.250 2249.955 2368.440 2249.985 ;
        RECT 2365.940 2249.765 2366.270 2249.955 ;
        RECT 2368.250 2249.715 2368.580 2249.955 ;
        RECT 2370.990 2249.495 2371.320 2250.430 ;
        RECT 2372.680 2249.700 2372.850 2250.430 ;
        RECT 2375.425 2249.700 2375.595 2250.430 ;
        RECT 2376.415 2249.700 2376.585 2250.430 ;
        RECT 2377.225 2250.425 2381.205 2250.430 ;
        RECT 2380.880 2250.125 2381.140 2250.425 ;
        RECT 2382.105 2250.135 2382.725 2250.635 ;
        RECT 2382.525 2249.955 2382.725 2250.135 ;
        RECT 2383.535 2250.095 2383.755 2250.635 ;
        RECT 2384.405 2249.985 2385.015 2250.635 ;
        RECT 2385.835 2250.095 2386.095 2250.635 ;
        RECT 2387.575 2250.430 2397.790 2250.635 ;
        RECT 2384.835 2249.955 2385.025 2249.985 ;
        RECT 2382.525 2249.765 2382.855 2249.955 ;
        RECT 2384.835 2249.715 2385.165 2249.955 ;
        RECT 2387.575 2249.495 2387.905 2250.430 ;
        RECT 2389.265 2249.700 2389.435 2250.430 ;
        RECT 2392.010 2249.700 2392.180 2250.430 ;
        RECT 2393.000 2249.700 2393.170 2250.430 ;
        RECT 2393.805 2250.425 2397.790 2250.430 ;
        RECT 2397.465 2250.125 2397.725 2250.425 ;
        RECT 2398.690 2250.135 2399.310 2250.635 ;
        RECT 2399.110 2249.955 2399.310 2250.135 ;
        RECT 2400.120 2250.095 2400.340 2250.635 ;
        RECT 2400.990 2249.985 2401.600 2250.635 ;
        RECT 2402.420 2250.095 2402.680 2250.635 ;
        RECT 2404.160 2250.430 2414.375 2250.635 ;
        RECT 2401.420 2249.955 2401.610 2249.985 ;
        RECT 2399.110 2249.765 2399.440 2249.955 ;
        RECT 2401.420 2249.715 2401.750 2249.955 ;
        RECT 2404.160 2249.495 2404.490 2250.430 ;
        RECT 2405.850 2249.700 2406.020 2250.430 ;
        RECT 2408.595 2249.700 2408.765 2250.430 ;
        RECT 2409.585 2249.700 2409.755 2250.430 ;
        RECT 2410.385 2250.425 2414.375 2250.430 ;
        RECT 2414.050 2250.125 2414.310 2250.425 ;
        RECT 2415.275 2250.135 2415.895 2250.635 ;
        RECT 2415.695 2249.955 2415.895 2250.135 ;
        RECT 2416.705 2250.095 2416.925 2250.635 ;
        RECT 2417.575 2249.985 2418.185 2250.635 ;
        RECT 2419.005 2250.095 2419.265 2250.635 ;
        RECT 2420.745 2250.430 2430.960 2250.635 ;
        RECT 2418.005 2249.955 2418.195 2249.985 ;
        RECT 2415.695 2249.765 2416.025 2249.955 ;
        RECT 2418.005 2249.715 2418.335 2249.955 ;
        RECT 2420.745 2249.495 2421.075 2250.430 ;
        RECT 2422.435 2249.700 2422.605 2250.430 ;
        RECT 2425.180 2249.700 2425.350 2250.430 ;
        RECT 2426.170 2249.700 2426.340 2250.430 ;
        RECT 2426.965 2250.425 2430.955 2250.430 ;
        RECT 2430.630 2250.125 2430.890 2250.425 ;
        RECT 2431.855 2250.135 2432.475 2250.635 ;
        RECT 2432.275 2249.955 2432.475 2250.135 ;
        RECT 2433.285 2250.095 2433.505 2250.635 ;
        RECT 2434.155 2249.985 2434.765 2250.635 ;
        RECT 2435.585 2250.095 2435.845 2250.635 ;
        RECT 2437.325 2250.430 2443.725 2250.635 ;
        RECT 2434.585 2249.955 2434.775 2249.985 ;
        RECT 2432.275 2249.765 2432.605 2249.955 ;
        RECT 2434.585 2249.715 2434.915 2249.955 ;
        RECT 2437.325 2249.495 2437.655 2250.430 ;
        RECT 2439.015 2249.700 2439.185 2250.430 ;
        RECT 2441.760 2249.700 2441.930 2250.430 ;
        RECT 2442.750 2249.700 2442.920 2250.430 ;
        RECT 2696.295 2215.375 2696.815 2215.915 ;
        RECT 2695.605 2214.285 2696.815 2215.375 ;
        RECT 2697.425 2214.285 2697.755 2215.065 ;
        RECT 2698.315 2214.285 2698.650 2214.710 ;
        RECT 2699.265 2214.285 2699.595 2215.045 ;
        RECT 2700.645 2214.285 2700.975 2215.045 ;
        RECT 2704.990 2214.720 2705.340 2215.970 ;
        RECT 2707.795 2215.375 2708.315 2215.915 ;
        RECT 2701.585 2214.285 2706.930 2214.720 ;
        RECT 2707.105 2214.285 2708.315 2215.375 ;
        RECT 2708.485 2214.285 2708.775 2215.450 ;
        RECT 2709.420 2214.285 2709.750 2215.045 ;
        RECT 2710.350 2214.285 2710.610 2215.435 ;
        RECT 2714.190 2214.720 2714.540 2215.970 ;
        RECT 2718.125 2215.375 2719.815 2215.895 ;
        RECT 2720.675 2215.375 2721.195 2215.915 ;
        RECT 2710.785 2214.285 2716.130 2214.720 ;
        RECT 2716.305 2214.285 2719.815 2215.375 ;
        RECT 2719.985 2214.285 2721.195 2215.375 ;
        RECT 2721.365 2214.285 2721.655 2215.450 ;
        RECT 2721.830 2214.285 2722.165 2214.710 ;
        RECT 2722.725 2214.285 2723.055 2215.065 ;
        RECT 2727.070 2214.720 2727.420 2215.970 ;
        RECT 2730.105 2215.375 2730.855 2215.895 ;
        RECT 2723.665 2214.285 2729.010 2214.720 ;
        RECT 2729.185 2214.285 2730.855 2215.375 ;
        RECT 2732.865 2215.375 2733.385 2215.915 ;
        RECT 2731.925 2214.285 2732.255 2215.045 ;
        RECT 2732.865 2214.285 2734.075 2215.375 ;
        RECT 2695.520 2214.115 2734.160 2214.285 ;
        RECT 2695.605 2213.025 2696.815 2214.115 ;
        RECT 2697.425 2213.355 2697.755 2214.115 ;
        RECT 2698.365 2213.680 2703.710 2214.115 ;
        RECT 2696.295 2212.485 2696.815 2213.025 ;
        RECT 2701.770 2212.430 2702.120 2213.680 ;
        RECT 2703.885 2213.025 2707.395 2214.115 ;
        RECT 2705.705 2212.505 2707.395 2213.025 ;
        RECT 2708.485 2212.950 2708.775 2214.115 ;
        RECT 2708.945 2213.680 2714.290 2214.115 ;
        RECT 2714.465 2213.680 2719.810 2214.115 ;
        RECT 2719.985 2213.680 2725.330 2214.115 ;
        RECT 2725.505 2213.680 2730.850 2214.115 ;
        RECT 2712.350 2212.430 2712.700 2213.680 ;
        RECT 2717.870 2212.430 2718.220 2213.680 ;
        RECT 2723.390 2212.430 2723.740 2213.680 ;
        RECT 2728.910 2212.430 2729.260 2213.680 ;
        RECT 2731.025 2213.025 2732.695 2214.115 ;
        RECT 2731.945 2212.505 2732.695 2213.025 ;
        RECT 2732.865 2213.025 2734.075 2214.115 ;
        RECT 2732.865 2212.485 2733.385 2213.025 ;
        RECT 2696.295 2209.935 2696.815 2210.475 ;
        RECT 2695.605 2208.845 2696.815 2209.935 ;
        RECT 2700.390 2209.280 2700.740 2210.530 ;
        RECT 2705.910 2209.280 2706.260 2210.530 ;
        RECT 2711.430 2209.280 2711.780 2210.530 ;
        RECT 2716.950 2209.280 2717.300 2210.530 ;
        RECT 2719.985 2209.935 2720.735 2210.455 ;
        RECT 2696.985 2208.845 2702.330 2209.280 ;
        RECT 2702.505 2208.845 2707.850 2209.280 ;
        RECT 2708.025 2208.845 2713.370 2209.280 ;
        RECT 2713.545 2208.845 2718.890 2209.280 ;
        RECT 2719.065 2208.845 2720.735 2209.935 ;
        RECT 2721.365 2208.845 2721.655 2210.010 ;
        RECT 2725.230 2209.280 2725.580 2210.530 ;
        RECT 2730.750 2209.280 2731.100 2210.530 ;
        RECT 2732.865 2209.935 2733.385 2210.475 ;
        RECT 2721.825 2208.845 2727.170 2209.280 ;
        RECT 2727.345 2208.845 2732.690 2209.280 ;
        RECT 2732.865 2208.845 2734.075 2209.935 ;
        RECT 2695.520 2208.675 2734.160 2208.845 ;
        RECT 2695.605 2207.585 2696.815 2208.675 ;
        RECT 2696.985 2208.240 2702.330 2208.675 ;
        RECT 2702.505 2208.240 2707.850 2208.675 ;
        RECT 2696.295 2207.045 2696.815 2207.585 ;
        RECT 2700.390 2206.990 2700.740 2208.240 ;
        RECT 2705.910 2206.990 2706.260 2208.240 ;
        RECT 2708.485 2207.510 2708.775 2208.675 ;
        RECT 2708.945 2208.240 2714.290 2208.675 ;
        RECT 2714.465 2208.240 2719.810 2208.675 ;
        RECT 2719.985 2208.240 2725.330 2208.675 ;
        RECT 2725.505 2208.240 2730.850 2208.675 ;
        RECT 2712.350 2206.990 2712.700 2208.240 ;
        RECT 2717.870 2206.990 2718.220 2208.240 ;
        RECT 2723.390 2206.990 2723.740 2208.240 ;
        RECT 2728.910 2206.990 2729.260 2208.240 ;
        RECT 2731.025 2207.585 2732.695 2208.675 ;
        RECT 2731.945 2207.065 2732.695 2207.585 ;
        RECT 2732.865 2207.585 2734.075 2208.675 ;
        RECT 2732.865 2207.045 2733.385 2207.585 ;
        RECT 2696.295 2204.495 2696.815 2205.035 ;
        RECT 2695.605 2203.405 2696.815 2204.495 ;
        RECT 2697.425 2203.405 2697.755 2204.165 ;
        RECT 2701.770 2203.840 2702.120 2205.090 ;
        RECT 2707.290 2203.840 2707.640 2205.090 ;
        RECT 2712.810 2203.840 2713.160 2205.090 ;
        RECT 2718.330 2203.840 2718.680 2205.090 ;
        RECT 2698.365 2203.405 2703.710 2203.840 ;
        RECT 2703.885 2203.405 2709.230 2203.840 ;
        RECT 2709.405 2203.405 2714.750 2203.840 ;
        RECT 2714.925 2203.405 2720.270 2203.840 ;
        RECT 2721.365 2203.405 2721.655 2204.570 ;
        RECT 2725.230 2203.840 2725.580 2205.090 ;
        RECT 2730.750 2203.840 2731.100 2205.090 ;
        RECT 2732.865 2204.495 2733.385 2205.035 ;
        RECT 2721.825 2203.405 2727.170 2203.840 ;
        RECT 2727.345 2203.405 2732.690 2203.840 ;
        RECT 2732.865 2203.405 2734.075 2204.495 ;
        RECT 2695.520 2203.235 2734.160 2203.405 ;
        RECT 2695.605 2202.145 2696.815 2203.235 ;
        RECT 2696.985 2202.800 2702.330 2203.235 ;
        RECT 2702.505 2202.800 2707.850 2203.235 ;
        RECT 2696.295 2201.605 2696.815 2202.145 ;
        RECT 2700.390 2201.550 2700.740 2202.800 ;
        RECT 2705.910 2201.550 2706.260 2202.800 ;
        RECT 2708.485 2202.070 2708.775 2203.235 ;
        RECT 2708.945 2202.800 2714.290 2203.235 ;
        RECT 2714.465 2202.800 2719.810 2203.235 ;
        RECT 2719.985 2202.800 2725.330 2203.235 ;
        RECT 2725.505 2202.800 2730.850 2203.235 ;
        RECT 2712.350 2201.550 2712.700 2202.800 ;
        RECT 2717.870 2201.550 2718.220 2202.800 ;
        RECT 2723.390 2201.550 2723.740 2202.800 ;
        RECT 2728.910 2201.550 2729.260 2202.800 ;
        RECT 2731.025 2202.145 2732.695 2203.235 ;
        RECT 2731.945 2201.625 2732.695 2202.145 ;
        RECT 2732.865 2202.145 2734.075 2203.235 ;
        RECT 2732.865 2201.605 2733.385 2202.145 ;
        RECT 2696.295 2199.055 2696.815 2199.595 ;
        RECT 2695.605 2197.965 2696.815 2199.055 ;
        RECT 2710.050 2198.400 2710.400 2199.650 ;
        RECT 2715.570 2198.400 2715.920 2199.650 ;
        RECT 2719.505 2199.055 2721.195 2199.575 ;
        RECT 2697.415 2197.965 2697.745 2198.345 ;
        RECT 2700.135 2197.965 2700.465 2198.345 ;
        RECT 2701.960 2197.965 2702.290 2198.345 ;
        RECT 2702.880 2197.965 2703.230 2198.345 ;
        RECT 2705.715 2197.965 2706.045 2198.345 ;
        RECT 2706.645 2197.965 2711.990 2198.400 ;
        RECT 2712.165 2197.965 2717.510 2198.400 ;
        RECT 2717.685 2197.965 2721.195 2199.055 ;
        RECT 2721.365 2197.965 2721.655 2199.130 ;
        RECT 2725.230 2198.400 2725.580 2199.650 ;
        RECT 2730.750 2198.400 2731.100 2199.650 ;
        RECT 2732.865 2199.055 2733.385 2199.595 ;
        RECT 2721.825 2197.965 2727.170 2198.400 ;
        RECT 2727.345 2197.965 2732.690 2198.400 ;
        RECT 2732.865 2197.965 2734.075 2199.055 ;
        RECT 2695.520 2197.795 2734.160 2197.965 ;
        RECT 2695.605 2196.705 2696.815 2197.795 ;
        RECT 2697.425 2197.035 2697.755 2197.795 ;
        RECT 2698.365 2197.360 2703.710 2197.795 ;
        RECT 2696.295 2196.165 2696.815 2196.705 ;
        RECT 2701.770 2196.110 2702.120 2197.360 ;
        RECT 2703.885 2196.705 2707.395 2197.795 ;
        RECT 2705.705 2196.185 2707.395 2196.705 ;
        RECT 2708.485 2196.630 2708.775 2197.795 ;
        RECT 2708.945 2197.360 2714.290 2197.795 ;
        RECT 2714.465 2197.360 2719.810 2197.795 ;
        RECT 2719.985 2197.360 2725.330 2197.795 ;
        RECT 2725.505 2197.360 2730.850 2197.795 ;
        RECT 2712.350 2196.110 2712.700 2197.360 ;
        RECT 2717.870 2196.110 2718.220 2197.360 ;
        RECT 2723.390 2196.110 2723.740 2197.360 ;
        RECT 2728.910 2196.110 2729.260 2197.360 ;
        RECT 2731.025 2196.705 2732.695 2197.795 ;
        RECT 2731.945 2196.185 2732.695 2196.705 ;
        RECT 2732.865 2196.705 2734.075 2197.795 ;
        RECT 2732.865 2196.165 2733.385 2196.705 ;
        RECT 2696.295 2193.615 2696.815 2194.155 ;
        RECT 2695.605 2192.525 2696.815 2193.615 ;
        RECT 2710.050 2192.960 2710.400 2194.210 ;
        RECT 2715.570 2192.960 2715.920 2194.210 ;
        RECT 2719.505 2193.615 2721.195 2194.135 ;
        RECT 2697.415 2192.525 2697.745 2192.905 ;
        RECT 2700.135 2192.525 2700.465 2192.905 ;
        RECT 2701.960 2192.525 2702.290 2192.905 ;
        RECT 2702.880 2192.525 2703.230 2192.905 ;
        RECT 2705.715 2192.525 2706.045 2192.905 ;
        RECT 2706.645 2192.525 2711.990 2192.960 ;
        RECT 2712.165 2192.525 2717.510 2192.960 ;
        RECT 2717.685 2192.525 2721.195 2193.615 ;
        RECT 2721.365 2192.525 2721.655 2193.690 ;
        RECT 2725.230 2192.960 2725.580 2194.210 ;
        RECT 2730.750 2192.960 2731.100 2194.210 ;
        RECT 2732.865 2193.615 2733.385 2194.155 ;
        RECT 2721.825 2192.525 2727.170 2192.960 ;
        RECT 2727.345 2192.525 2732.690 2192.960 ;
        RECT 2732.865 2192.525 2734.075 2193.615 ;
        RECT 2695.520 2192.355 2734.160 2192.525 ;
        RECT 2695.605 2191.265 2696.815 2192.355 ;
        RECT 2697.425 2191.595 2697.755 2192.355 ;
        RECT 2698.365 2191.265 2700.955 2192.355 ;
        RECT 2696.295 2190.725 2696.815 2191.265 ;
        RECT 2699.745 2190.745 2700.955 2191.265 ;
        RECT 2702.095 2191.215 2702.265 2192.355 ;
        RECT 2704.635 2191.595 2704.805 2192.355 ;
        RECT 2705.725 2191.265 2708.315 2192.355 ;
        RECT 2707.105 2190.745 2708.315 2191.265 ;
        RECT 2708.485 2191.190 2708.775 2192.355 ;
        RECT 2708.945 2191.920 2714.290 2192.355 ;
        RECT 2714.465 2191.920 2719.810 2192.355 ;
        RECT 2719.985 2191.920 2725.330 2192.355 ;
        RECT 2725.505 2191.920 2730.850 2192.355 ;
        RECT 2712.350 2190.670 2712.700 2191.920 ;
        RECT 2717.870 2190.670 2718.220 2191.920 ;
        RECT 2723.390 2190.670 2723.740 2191.920 ;
        RECT 2728.910 2190.670 2729.260 2191.920 ;
        RECT 2731.025 2191.265 2732.695 2192.355 ;
        RECT 2731.945 2190.745 2732.695 2191.265 ;
        RECT 2732.865 2191.265 2734.075 2192.355 ;
        RECT 2732.865 2190.725 2733.385 2191.265 ;
        RECT 2696.295 2188.175 2696.815 2188.715 ;
        RECT 2695.605 2187.085 2696.815 2188.175 ;
        RECT 2700.390 2187.520 2700.740 2188.770 ;
        RECT 2705.910 2187.520 2706.260 2188.770 ;
        RECT 2711.430 2187.520 2711.780 2188.770 ;
        RECT 2716.950 2187.520 2717.300 2188.770 ;
        RECT 2719.985 2188.175 2720.735 2188.695 ;
        RECT 2696.985 2187.085 2702.330 2187.520 ;
        RECT 2702.505 2187.085 2707.850 2187.520 ;
        RECT 2708.025 2187.085 2713.370 2187.520 ;
        RECT 2713.545 2187.085 2718.890 2187.520 ;
        RECT 2719.065 2187.085 2720.735 2188.175 ;
        RECT 2721.365 2187.085 2721.655 2188.250 ;
        RECT 2725.230 2187.520 2725.580 2188.770 ;
        RECT 2730.750 2187.520 2731.100 2188.770 ;
        RECT 2732.865 2188.175 2733.385 2188.715 ;
        RECT 2721.825 2187.085 2727.170 2187.520 ;
        RECT 2727.345 2187.085 2732.690 2187.520 ;
        RECT 2732.865 2187.085 2734.075 2188.175 ;
        RECT 2695.520 2186.915 2734.160 2187.085 ;
        RECT 2695.605 2185.825 2696.815 2186.915 ;
        RECT 2697.425 2186.155 2697.755 2186.915 ;
        RECT 2698.365 2186.480 2703.710 2186.915 ;
        RECT 2696.295 2185.285 2696.815 2185.825 ;
        RECT 2701.770 2185.230 2702.120 2186.480 ;
        RECT 2703.885 2185.825 2707.395 2186.915 ;
        RECT 2705.705 2185.305 2707.395 2185.825 ;
        RECT 2708.485 2185.750 2708.775 2186.915 ;
        RECT 2708.945 2186.480 2714.290 2186.915 ;
        RECT 2714.465 2186.480 2719.810 2186.915 ;
        RECT 2719.985 2186.480 2725.330 2186.915 ;
        RECT 2725.505 2186.480 2730.850 2186.915 ;
        RECT 2712.350 2185.230 2712.700 2186.480 ;
        RECT 2717.870 2185.230 2718.220 2186.480 ;
        RECT 2723.390 2185.230 2723.740 2186.480 ;
        RECT 2728.910 2185.230 2729.260 2186.480 ;
        RECT 2731.025 2185.825 2732.695 2186.915 ;
        RECT 2731.945 2185.305 2732.695 2185.825 ;
        RECT 2732.865 2185.825 2734.075 2186.915 ;
        RECT 2732.865 2185.285 2733.385 2185.825 ;
        RECT 2696.295 2182.735 2696.815 2183.275 ;
        RECT 2695.605 2181.645 2696.815 2182.735 ;
        RECT 2700.390 2182.080 2700.740 2183.330 ;
        RECT 2705.910 2182.080 2706.260 2183.330 ;
        RECT 2711.430 2182.080 2711.780 2183.330 ;
        RECT 2716.950 2182.080 2717.300 2183.330 ;
        RECT 2719.985 2182.735 2720.735 2183.255 ;
        RECT 2696.985 2181.645 2702.330 2182.080 ;
        RECT 2702.505 2181.645 2707.850 2182.080 ;
        RECT 2708.025 2181.645 2713.370 2182.080 ;
        RECT 2713.545 2181.645 2718.890 2182.080 ;
        RECT 2719.065 2181.645 2720.735 2182.735 ;
        RECT 2721.365 2181.645 2721.655 2182.810 ;
        RECT 2725.230 2182.080 2725.580 2183.330 ;
        RECT 2730.750 2182.080 2731.100 2183.330 ;
        RECT 2732.865 2182.735 2733.385 2183.275 ;
        RECT 2721.825 2181.645 2727.170 2182.080 ;
        RECT 2727.345 2181.645 2732.690 2182.080 ;
        RECT 2732.865 2181.645 2734.075 2182.735 ;
        RECT 2695.520 2181.475 2734.160 2181.645 ;
        RECT 2695.605 2180.385 2696.815 2181.475 ;
        RECT 2696.985 2180.385 2700.495 2181.475 ;
        RECT 2696.295 2179.845 2696.815 2180.385 ;
        RECT 2698.805 2179.865 2700.495 2180.385 ;
        RECT 2702.455 2180.335 2702.785 2181.475 ;
        RECT 2702.965 2181.040 2708.310 2181.475 ;
        RECT 2706.370 2179.790 2706.720 2181.040 ;
        RECT 2708.485 2180.310 2708.775 2181.475 ;
        RECT 2708.945 2181.040 2714.290 2181.475 ;
        RECT 2714.465 2181.040 2719.810 2181.475 ;
        RECT 2719.985 2181.040 2725.330 2181.475 ;
        RECT 2725.505 2181.040 2730.850 2181.475 ;
        RECT 2712.350 2179.790 2712.700 2181.040 ;
        RECT 2717.870 2179.790 2718.220 2181.040 ;
        RECT 2723.390 2179.790 2723.740 2181.040 ;
        RECT 2728.910 2179.790 2729.260 2181.040 ;
        RECT 2731.025 2180.385 2732.695 2181.475 ;
        RECT 2731.945 2179.865 2732.695 2180.385 ;
        RECT 2732.865 2180.385 2734.075 2181.475 ;
        RECT 2732.865 2179.845 2733.385 2180.385 ;
        RECT 2696.295 2177.295 2696.815 2177.835 ;
        RECT 2700.185 2177.295 2701.875 2177.815 ;
        RECT 2695.605 2176.205 2696.815 2177.295 ;
        RECT 2697.425 2176.205 2697.755 2176.965 ;
        RECT 2698.365 2176.205 2701.875 2177.295 ;
        RECT 2703.535 2176.205 2703.705 2176.645 ;
        RECT 2708.670 2176.640 2709.020 2177.890 ;
        RECT 2714.190 2176.640 2714.540 2177.890 ;
        RECT 2718.125 2177.295 2719.815 2177.815 ;
        RECT 2720.675 2177.295 2721.195 2177.835 ;
        RECT 2704.310 2176.205 2704.640 2176.565 ;
        RECT 2705.265 2176.205 2710.610 2176.640 ;
        RECT 2710.785 2176.205 2716.130 2176.640 ;
        RECT 2716.305 2176.205 2719.815 2177.295 ;
        RECT 2719.985 2176.205 2721.195 2177.295 ;
        RECT 2721.365 2176.205 2721.655 2177.370 ;
        RECT 2725.230 2176.640 2725.580 2177.890 ;
        RECT 2730.750 2176.640 2731.100 2177.890 ;
        RECT 2732.865 2177.295 2733.385 2177.835 ;
        RECT 2721.825 2176.205 2727.170 2176.640 ;
        RECT 2727.345 2176.205 2732.690 2176.640 ;
        RECT 2732.865 2176.205 2734.075 2177.295 ;
        RECT 2695.520 2176.035 2734.160 2176.205 ;
        RECT 2695.605 2174.945 2696.815 2176.035 ;
        RECT 2696.985 2175.600 2702.330 2176.035 ;
        RECT 2702.505 2175.600 2707.850 2176.035 ;
        RECT 2696.295 2174.405 2696.815 2174.945 ;
        RECT 2700.390 2174.350 2700.740 2175.600 ;
        RECT 2705.910 2174.350 2706.260 2175.600 ;
        RECT 2708.485 2174.870 2708.775 2176.035 ;
        RECT 2708.945 2175.600 2714.290 2176.035 ;
        RECT 2714.465 2175.600 2719.810 2176.035 ;
        RECT 2719.985 2175.600 2725.330 2176.035 ;
        RECT 2712.350 2174.350 2712.700 2175.600 ;
        RECT 2717.870 2174.350 2718.220 2175.600 ;
        RECT 2723.390 2174.350 2723.740 2175.600 ;
        RECT 2725.595 2175.235 2725.765 2176.035 ;
        RECT 2726.435 2175.235 2726.605 2176.035 ;
        RECT 2727.275 2175.235 2727.445 2176.035 ;
        RECT 2728.035 2175.235 2728.365 2176.035 ;
        RECT 2728.875 2175.235 2729.205 2176.035 ;
        RECT 2729.715 2175.235 2730.045 2176.035 ;
        RECT 2730.555 2175.235 2730.885 2176.035 ;
        RECT 2731.395 2175.235 2731.725 2176.035 ;
        RECT 2732.235 2174.885 2732.565 2176.035 ;
        RECT 2732.865 2174.945 2734.075 2176.035 ;
        RECT 2732.865 2174.405 2733.385 2174.945 ;
        RECT 2696.295 2171.855 2696.815 2172.395 ;
        RECT 2695.605 2170.765 2696.815 2171.855 ;
        RECT 2697.425 2170.765 2697.755 2171.525 ;
        RECT 2701.770 2171.200 2702.120 2172.450 ;
        RECT 2707.290 2171.200 2707.640 2172.450 ;
        RECT 2712.810 2171.200 2713.160 2172.450 ;
        RECT 2718.330 2171.200 2718.680 2172.450 ;
        RECT 2698.365 2170.765 2703.710 2171.200 ;
        RECT 2703.885 2170.765 2709.230 2171.200 ;
        RECT 2709.405 2170.765 2714.750 2171.200 ;
        RECT 2714.925 2170.765 2720.270 2171.200 ;
        RECT 2721.365 2170.765 2721.655 2171.930 ;
        RECT 2725.230 2171.200 2725.580 2172.450 ;
        RECT 2730.750 2171.200 2731.100 2172.450 ;
        RECT 2732.865 2171.855 2733.385 2172.395 ;
        RECT 2721.825 2170.765 2727.170 2171.200 ;
        RECT 2727.345 2170.765 2732.690 2171.200 ;
        RECT 2732.865 2170.765 2734.075 2171.855 ;
        RECT 2695.520 2170.595 2734.160 2170.765 ;
        RECT 2695.605 2169.505 2696.815 2170.595 ;
        RECT 2696.985 2170.160 2702.330 2170.595 ;
        RECT 2702.505 2170.160 2707.850 2170.595 ;
        RECT 2696.295 2168.965 2696.815 2169.505 ;
        RECT 2700.390 2168.910 2700.740 2170.160 ;
        RECT 2705.910 2168.910 2706.260 2170.160 ;
        RECT 2708.485 2169.430 2708.775 2170.595 ;
        RECT 2708.945 2170.160 2714.290 2170.595 ;
        RECT 2714.465 2170.160 2719.810 2170.595 ;
        RECT 2719.985 2170.160 2725.330 2170.595 ;
        RECT 2725.505 2170.160 2730.850 2170.595 ;
        RECT 2712.350 2168.910 2712.700 2170.160 ;
        RECT 2717.870 2168.910 2718.220 2170.160 ;
        RECT 2723.390 2168.910 2723.740 2170.160 ;
        RECT 2728.910 2168.910 2729.260 2170.160 ;
        RECT 2731.025 2169.505 2732.695 2170.595 ;
        RECT 2731.945 2168.985 2732.695 2169.505 ;
        RECT 2732.865 2169.505 2734.075 2170.595 ;
        RECT 2732.865 2168.965 2733.385 2169.505 ;
        RECT 2696.295 2166.415 2696.815 2166.955 ;
        RECT 2695.605 2165.325 2696.815 2166.415 ;
        RECT 2697.715 2165.325 2698.045 2165.835 ;
        RECT 2703.150 2165.760 2703.500 2167.010 ;
        RECT 2708.670 2165.760 2709.020 2167.010 ;
        RECT 2714.190 2165.760 2714.540 2167.010 ;
        RECT 2718.125 2166.415 2719.815 2166.935 ;
        RECT 2720.675 2166.415 2721.195 2166.955 ;
        RECT 2699.745 2165.325 2705.090 2165.760 ;
        RECT 2705.265 2165.325 2710.610 2165.760 ;
        RECT 2710.785 2165.325 2716.130 2165.760 ;
        RECT 2716.305 2165.325 2719.815 2166.415 ;
        RECT 2719.985 2165.325 2721.195 2166.415 ;
        RECT 2721.365 2165.325 2721.655 2166.490 ;
        RECT 2725.230 2165.760 2725.580 2167.010 ;
        RECT 2730.750 2165.760 2731.100 2167.010 ;
        RECT 2732.865 2166.415 2733.385 2166.955 ;
        RECT 2721.825 2165.325 2727.170 2165.760 ;
        RECT 2727.345 2165.325 2732.690 2165.760 ;
        RECT 2732.865 2165.325 2734.075 2166.415 ;
        RECT 2695.520 2165.155 2734.160 2165.325 ;
        RECT 2695.605 2164.065 2696.815 2165.155 ;
        RECT 2697.425 2164.395 2697.755 2165.155 ;
        RECT 2698.365 2164.720 2703.710 2165.155 ;
        RECT 2360.055 2163.045 2360.230 2163.595 ;
        RECT 2696.295 2163.525 2696.815 2164.065 ;
        RECT 2701.770 2163.470 2702.120 2164.720 ;
        RECT 2703.885 2164.065 2707.395 2165.155 ;
        RECT 2705.705 2163.545 2707.395 2164.065 ;
        RECT 2708.485 2163.990 2708.775 2165.155 ;
        RECT 2708.945 2164.720 2714.290 2165.155 ;
        RECT 2714.465 2164.720 2719.810 2165.155 ;
        RECT 2719.985 2164.720 2725.330 2165.155 ;
        RECT 2725.505 2164.720 2730.850 2165.155 ;
        RECT 2712.350 2163.470 2712.700 2164.720 ;
        RECT 2717.870 2163.470 2718.220 2164.720 ;
        RECT 2723.390 2163.470 2723.740 2164.720 ;
        RECT 2728.910 2163.470 2729.260 2164.720 ;
        RECT 2731.025 2164.065 2732.695 2165.155 ;
        RECT 2731.945 2163.545 2732.695 2164.065 ;
        RECT 2732.865 2164.065 2734.075 2165.155 ;
        RECT 2732.865 2163.525 2733.385 2164.065 ;
        RECT 2360.055 2161.445 2360.225 2163.045 ;
        RECT 2358.240 2160.035 2358.410 2160.765 ;
        RECT 2360.055 2160.305 2360.230 2161.445 ;
        RECT 2696.295 2160.975 2696.815 2161.515 ;
        RECT 2360.055 2160.035 2360.225 2160.305 ;
        RECT 2358.070 2160.030 2360.820 2160.035 ;
        RECT 2361.650 2160.030 2361.820 2160.755 ;
        RECT 2373.335 2160.035 2373.505 2160.765 ;
        RECT 2376.080 2160.035 2376.250 2160.765 ;
        RECT 2377.070 2160.035 2377.240 2160.765 ;
        RECT 2373.165 2160.030 2377.890 2160.035 ;
        RECT 2378.870 2160.030 2379.040 2160.755 ;
        RECT 2390.555 2160.035 2390.725 2160.765 ;
        RECT 2393.300 2160.035 2393.470 2160.765 ;
        RECT 2394.290 2160.035 2394.460 2160.765 ;
        RECT 2390.385 2160.030 2395.110 2160.035 ;
        RECT 2396.090 2160.030 2396.260 2160.755 ;
        RECT 2407.775 2160.035 2407.945 2160.765 ;
        RECT 2410.520 2160.035 2410.690 2160.765 ;
        RECT 2411.510 2160.035 2411.680 2160.765 ;
        RECT 2407.605 2160.030 2412.330 2160.035 ;
        RECT 2413.310 2160.030 2413.480 2160.755 ;
        RECT 2424.995 2160.035 2425.165 2160.765 ;
        RECT 2427.740 2160.035 2427.910 2160.765 ;
        RECT 2428.730 2160.035 2428.900 2160.765 ;
        RECT 2424.825 2160.030 2429.550 2160.035 ;
        RECT 2430.530 2160.030 2430.700 2160.755 ;
        RECT 2442.215 2160.035 2442.385 2160.765 ;
        RECT 2444.960 2160.035 2445.130 2160.765 ;
        RECT 2445.950 2160.035 2446.120 2160.765 ;
        RECT 2442.045 2160.030 2446.770 2160.035 ;
        RECT 2358.070 2160.025 2364.495 2160.030 ;
        RECT 2343.015 2160.000 2364.500 2160.025 ;
        RECT 2371.960 2160.000 2381.715 2160.030 ;
        RECT 2389.180 2160.000 2398.935 2160.030 ;
        RECT 2406.400 2160.000 2416.155 2160.030 ;
        RECT 2423.620 2160.000 2433.375 2160.030 ;
        RECT 2343.015 2158.810 2364.625 2160.000 ;
        RECT 2365.155 2158.810 2365.435 2159.950 ;
        RECT 2366.105 2158.810 2366.365 2159.950 ;
        RECT 2367.455 2158.810 2367.735 2159.950 ;
        RECT 2368.405 2158.810 2368.665 2159.950 ;
        RECT 2368.835 2158.810 2369.095 2159.950 ;
        RECT 2369.765 2158.810 2370.045 2159.950 ;
        RECT 2370.215 2158.810 2370.475 2159.950 ;
        RECT 2371.145 2158.810 2371.425 2159.950 ;
        RECT 2371.960 2158.810 2381.845 2160.000 ;
        RECT 2382.375 2158.810 2382.655 2159.950 ;
        RECT 2383.325 2158.810 2383.585 2159.950 ;
        RECT 2384.675 2158.810 2384.955 2159.950 ;
        RECT 2385.625 2158.810 2385.885 2159.950 ;
        RECT 2386.055 2158.810 2386.315 2159.950 ;
        RECT 2386.985 2158.810 2387.265 2159.950 ;
        RECT 2387.435 2158.810 2387.695 2159.950 ;
        RECT 2388.365 2158.810 2388.645 2159.950 ;
        RECT 2389.180 2158.810 2399.065 2160.000 ;
        RECT 2399.595 2158.810 2399.875 2159.950 ;
        RECT 2400.545 2158.810 2400.805 2159.950 ;
        RECT 2401.895 2158.810 2402.175 2159.950 ;
        RECT 2402.845 2158.810 2403.105 2159.950 ;
        RECT 2403.275 2158.810 2403.535 2159.950 ;
        RECT 2404.205 2158.810 2404.485 2159.950 ;
        RECT 2404.655 2158.810 2404.915 2159.950 ;
        RECT 2405.585 2158.810 2405.865 2159.950 ;
        RECT 2406.400 2158.810 2416.285 2160.000 ;
        RECT 2416.815 2158.810 2417.095 2159.950 ;
        RECT 2417.765 2158.810 2418.025 2159.950 ;
        RECT 2419.115 2158.810 2419.395 2159.950 ;
        RECT 2420.065 2158.810 2420.325 2159.950 ;
        RECT 2420.495 2158.810 2420.755 2159.950 ;
        RECT 2421.425 2158.810 2421.705 2159.950 ;
        RECT 2421.875 2158.810 2422.135 2159.950 ;
        RECT 2422.805 2158.810 2423.085 2159.950 ;
        RECT 2423.620 2158.810 2433.505 2160.000 ;
        RECT 2434.035 2158.810 2434.315 2159.950 ;
        RECT 2434.985 2158.810 2435.245 2159.950 ;
        RECT 2436.335 2158.810 2436.615 2159.950 ;
        RECT 2437.285 2158.810 2437.545 2159.950 ;
        RECT 2437.715 2158.810 2437.975 2159.950 ;
        RECT 2438.645 2158.810 2438.925 2159.950 ;
        RECT 2439.095 2158.810 2439.355 2159.950 ;
        RECT 2440.025 2158.810 2440.305 2159.950 ;
        RECT 2440.840 2158.810 2446.925 2160.030 ;
        RECT 2695.605 2159.885 2696.815 2160.975 ;
        RECT 2697.735 2159.885 2697.905 2160.645 ;
        RECT 2700.275 2159.885 2700.445 2161.025 ;
        RECT 2701.590 2159.885 2701.920 2160.600 ;
        RECT 2708.210 2160.320 2708.560 2161.570 ;
        RECT 2713.730 2160.320 2714.080 2161.570 ;
        RECT 2719.250 2160.320 2719.600 2161.570 ;
        RECT 2704.805 2159.885 2710.150 2160.320 ;
        RECT 2710.325 2159.885 2715.670 2160.320 ;
        RECT 2715.845 2159.885 2721.190 2160.320 ;
        RECT 2721.365 2159.885 2721.655 2161.050 ;
        RECT 2725.230 2160.320 2725.580 2161.570 ;
        RECT 2730.750 2160.320 2731.100 2161.570 ;
        RECT 2732.865 2160.975 2733.385 2161.515 ;
        RECT 2721.825 2159.885 2727.170 2160.320 ;
        RECT 2727.345 2159.885 2732.690 2160.320 ;
        RECT 2732.865 2159.885 2734.075 2160.975 ;
        RECT 2881.580 2160.100 2883.380 2160.270 ;
        RECT 2695.520 2159.715 2734.160 2159.885 ;
        RECT 2343.015 2158.640 2446.925 2158.810 ;
        RECT 2343.015 2158.425 2364.965 2158.640 ;
        RECT 2364.755 2157.500 2364.965 2158.425 ;
        RECT 2365.635 2157.500 2365.865 2158.640 ;
        RECT 2366.085 2157.500 2366.415 2158.640 ;
        RECT 2368.325 2157.500 2368.655 2158.640 ;
        RECT 2369.905 2158.130 2370.075 2158.640 ;
        RECT 2370.745 2157.790 2370.915 2158.640 ;
        RECT 2372.055 2158.430 2382.185 2158.640 ;
        RECT 2373.165 2158.425 2382.185 2158.430 ;
        RECT 2373.335 2157.695 2373.505 2158.425 ;
        RECT 2376.080 2157.695 2376.250 2158.425 ;
        RECT 2377.065 2157.695 2377.235 2158.425 ;
        RECT 2381.975 2157.500 2382.185 2158.425 ;
        RECT 2382.855 2157.500 2383.085 2158.640 ;
        RECT 2383.305 2157.500 2383.635 2158.640 ;
        RECT 2385.545 2157.500 2385.875 2158.640 ;
        RECT 2387.125 2158.130 2387.295 2158.640 ;
        RECT 2387.965 2157.790 2388.135 2158.640 ;
        RECT 2389.275 2158.430 2399.405 2158.640 ;
        RECT 2390.385 2158.425 2399.405 2158.430 ;
        RECT 2390.555 2157.695 2390.725 2158.425 ;
        RECT 2393.300 2157.695 2393.470 2158.425 ;
        RECT 2394.285 2157.695 2394.455 2158.425 ;
        RECT 2399.195 2157.500 2399.405 2158.425 ;
        RECT 2400.075 2157.500 2400.305 2158.640 ;
        RECT 2400.525 2157.500 2400.855 2158.640 ;
        RECT 2402.765 2157.500 2403.095 2158.640 ;
        RECT 2404.345 2158.130 2404.515 2158.640 ;
        RECT 2405.185 2157.790 2405.355 2158.640 ;
        RECT 2406.495 2158.430 2416.625 2158.640 ;
        RECT 2407.605 2158.425 2416.625 2158.430 ;
        RECT 2407.775 2157.695 2407.945 2158.425 ;
        RECT 2410.520 2157.695 2410.690 2158.425 ;
        RECT 2411.505 2157.695 2411.675 2158.425 ;
        RECT 2416.415 2157.500 2416.625 2158.425 ;
        RECT 2417.295 2157.500 2417.525 2158.640 ;
        RECT 2417.745 2157.500 2418.075 2158.640 ;
        RECT 2419.985 2157.500 2420.315 2158.640 ;
        RECT 2421.565 2158.130 2421.735 2158.640 ;
        RECT 2422.405 2157.790 2422.575 2158.640 ;
        RECT 2423.715 2158.430 2433.845 2158.640 ;
        RECT 2424.825 2158.425 2433.845 2158.430 ;
        RECT 2424.995 2157.695 2425.165 2158.425 ;
        RECT 2427.740 2157.695 2427.910 2158.425 ;
        RECT 2428.725 2157.695 2428.895 2158.425 ;
        RECT 2433.635 2157.500 2433.845 2158.425 ;
        RECT 2434.515 2157.500 2434.745 2158.640 ;
        RECT 2434.965 2157.500 2435.295 2158.640 ;
        RECT 2437.205 2157.500 2437.535 2158.640 ;
        RECT 2438.785 2158.130 2438.955 2158.640 ;
        RECT 2439.625 2157.790 2439.795 2158.640 ;
        RECT 2440.935 2158.430 2446.925 2158.640 ;
        RECT 2695.605 2158.625 2696.815 2159.715 ;
        RECT 2696.985 2159.205 2697.245 2159.715 ;
        RECT 2697.905 2159.210 2698.520 2159.715 ;
        RECT 2698.325 2159.035 2698.520 2159.210 ;
        RECT 2699.335 2159.170 2699.550 2159.715 ;
        RECT 2700.205 2159.280 2705.550 2159.715 ;
        RECT 2698.325 2158.845 2698.655 2159.035 ;
        RECT 2442.045 2158.425 2446.765 2158.430 ;
        RECT 2442.215 2157.695 2442.385 2158.425 ;
        RECT 2444.960 2157.695 2445.130 2158.425 ;
        RECT 2445.945 2157.695 2446.115 2158.425 ;
        RECT 2696.295 2158.085 2696.815 2158.625 ;
        RECT 2703.610 2158.030 2703.960 2159.280 ;
        RECT 2705.725 2158.625 2708.315 2159.715 ;
        RECT 2707.105 2158.105 2708.315 2158.625 ;
        RECT 2708.485 2158.550 2708.775 2159.715 ;
        RECT 2708.945 2159.280 2714.290 2159.715 ;
        RECT 2714.465 2159.280 2719.810 2159.715 ;
        RECT 2719.985 2159.280 2725.330 2159.715 ;
        RECT 2725.505 2159.280 2730.850 2159.715 ;
        RECT 2712.350 2158.030 2712.700 2159.280 ;
        RECT 2717.870 2158.030 2718.220 2159.280 ;
        RECT 2723.390 2158.030 2723.740 2159.280 ;
        RECT 2728.910 2158.030 2729.260 2159.280 ;
        RECT 2731.025 2158.625 2732.695 2159.715 ;
        RECT 2731.945 2158.105 2732.695 2158.625 ;
        RECT 2732.865 2158.625 2734.075 2159.715 ;
        RECT 2882.775 2159.375 2883.105 2160.100 ;
        RECT 2732.865 2158.085 2733.385 2158.625 ;
        RECT 2696.295 2155.535 2696.815 2156.075 ;
        RECT 2695.605 2154.445 2696.815 2155.535 ;
        RECT 2697.425 2154.445 2697.755 2155.205 ;
        RECT 2701.770 2154.880 2702.120 2156.130 ;
        RECT 2707.290 2154.880 2707.640 2156.130 ;
        RECT 2712.810 2154.880 2713.160 2156.130 ;
        RECT 2718.330 2154.880 2718.680 2156.130 ;
        RECT 2698.365 2154.445 2703.710 2154.880 ;
        RECT 2703.885 2154.445 2709.230 2154.880 ;
        RECT 2709.405 2154.445 2714.750 2154.880 ;
        RECT 2714.925 2154.445 2720.270 2154.880 ;
        RECT 2721.365 2154.445 2721.655 2155.610 ;
        RECT 2725.230 2154.880 2725.580 2156.130 ;
        RECT 2730.750 2154.880 2731.100 2156.130 ;
        RECT 2732.865 2155.535 2733.385 2156.075 ;
        RECT 2721.825 2154.445 2727.170 2154.880 ;
        RECT 2727.345 2154.445 2732.690 2154.880 ;
        RECT 2732.865 2154.445 2734.075 2155.535 ;
        RECT 2695.520 2154.275 2734.160 2154.445 ;
        RECT 2695.605 2153.185 2696.815 2154.275 ;
        RECT 2696.985 2153.185 2698.195 2154.275 ;
        RECT 2698.865 2153.815 2699.115 2154.275 ;
        RECT 2699.795 2153.815 2700.045 2154.275 ;
        RECT 2701.115 2153.815 2701.365 2154.275 ;
        RECT 2702.045 2153.840 2707.390 2154.275 ;
        RECT 2696.295 2152.645 2696.815 2153.185 ;
        RECT 2697.675 2152.645 2698.195 2153.185 ;
        RECT 2705.450 2152.590 2705.800 2153.840 ;
        RECT 2708.485 2153.110 2708.775 2154.275 ;
        RECT 2708.945 2153.840 2714.290 2154.275 ;
        RECT 2714.465 2153.840 2719.810 2154.275 ;
        RECT 2719.985 2153.840 2725.330 2154.275 ;
        RECT 2725.505 2153.840 2730.850 2154.275 ;
        RECT 2712.350 2152.590 2712.700 2153.840 ;
        RECT 2717.870 2152.590 2718.220 2153.840 ;
        RECT 2723.390 2152.590 2723.740 2153.840 ;
        RECT 2728.910 2152.590 2729.260 2153.840 ;
        RECT 2731.025 2153.185 2732.695 2154.275 ;
        RECT 2731.945 2152.665 2732.695 2153.185 ;
        RECT 2732.865 2153.185 2734.075 2154.275 ;
        RECT 2732.865 2152.645 2733.385 2153.185 ;
        RECT 2696.295 2150.095 2696.815 2150.635 ;
        RECT 2695.605 2149.005 2696.815 2150.095 ;
        RECT 2697.905 2149.005 2698.165 2150.145 ;
        RECT 2700.190 2149.005 2700.470 2149.805 ;
        RECT 2701.885 2149.005 2702.170 2149.805 ;
        RECT 2702.840 2149.005 2703.090 2150.145 ;
        RECT 2707.290 2149.440 2707.640 2150.690 ;
        RECT 2712.810 2149.440 2713.160 2150.690 ;
        RECT 2718.330 2149.440 2718.680 2150.690 ;
        RECT 2703.885 2149.005 2709.230 2149.440 ;
        RECT 2709.405 2149.005 2714.750 2149.440 ;
        RECT 2714.925 2149.005 2720.270 2149.440 ;
        RECT 2721.365 2149.005 2721.655 2150.170 ;
        RECT 2725.230 2149.440 2725.580 2150.690 ;
        RECT 2730.750 2149.440 2731.100 2150.690 ;
        RECT 2732.865 2150.095 2733.385 2150.635 ;
        RECT 2721.825 2149.005 2727.170 2149.440 ;
        RECT 2727.345 2149.005 2732.690 2149.440 ;
        RECT 2732.865 2149.005 2734.075 2150.095 ;
        RECT 2695.520 2148.835 2734.160 2149.005 ;
        RECT 2695.605 2147.745 2696.815 2148.835 ;
        RECT 2697.425 2148.075 2697.755 2148.835 ;
        RECT 2696.295 2147.205 2696.815 2147.745 ;
        RECT 2698.825 2147.695 2699.085 2148.835 ;
        RECT 2699.755 2147.695 2700.035 2148.835 ;
        RECT 2700.205 2148.400 2705.550 2148.835 ;
        RECT 2703.610 2147.150 2703.960 2148.400 ;
        RECT 2705.725 2147.745 2708.315 2148.835 ;
        RECT 2707.105 2147.225 2708.315 2147.745 ;
        RECT 2708.485 2147.670 2708.775 2148.835 ;
        RECT 2708.945 2148.400 2714.290 2148.835 ;
        RECT 2714.465 2148.400 2719.810 2148.835 ;
        RECT 2719.985 2148.400 2725.330 2148.835 ;
        RECT 2725.505 2148.400 2730.850 2148.835 ;
        RECT 2712.350 2147.150 2712.700 2148.400 ;
        RECT 2717.870 2147.150 2718.220 2148.400 ;
        RECT 2723.390 2147.150 2723.740 2148.400 ;
        RECT 2728.910 2147.150 2729.260 2148.400 ;
        RECT 2731.025 2147.745 2732.695 2148.835 ;
        RECT 2731.945 2147.225 2732.695 2147.745 ;
        RECT 2732.865 2147.745 2734.075 2148.835 ;
        RECT 2732.865 2147.205 2733.385 2147.745 ;
        RECT 2696.295 2144.655 2696.815 2145.195 ;
        RECT 2695.605 2143.565 2696.815 2144.655 ;
        RECT 2697.735 2143.565 2697.905 2144.325 ;
        RECT 2700.275 2143.565 2700.445 2144.705 ;
        RECT 2704.530 2144.000 2704.880 2145.250 ;
        RECT 2710.050 2144.000 2710.400 2145.250 ;
        RECT 2715.570 2144.000 2715.920 2145.250 ;
        RECT 2719.505 2144.655 2721.195 2145.175 ;
        RECT 2701.125 2143.565 2706.470 2144.000 ;
        RECT 2706.645 2143.565 2711.990 2144.000 ;
        RECT 2712.165 2143.565 2717.510 2144.000 ;
        RECT 2717.685 2143.565 2721.195 2144.655 ;
        RECT 2721.365 2143.565 2721.655 2144.730 ;
        RECT 2725.230 2144.000 2725.580 2145.250 ;
        RECT 2730.750 2144.000 2731.100 2145.250 ;
        RECT 2732.865 2144.655 2733.385 2145.195 ;
        RECT 2721.825 2143.565 2727.170 2144.000 ;
        RECT 2727.345 2143.565 2732.690 2144.000 ;
        RECT 2732.865 2143.565 2734.075 2144.655 ;
        RECT 2695.520 2143.395 2734.160 2143.565 ;
        RECT 2695.605 2142.305 2696.815 2143.395 ;
        RECT 2697.425 2142.635 2697.755 2143.395 ;
        RECT 2698.365 2142.960 2703.710 2143.395 ;
        RECT 2696.295 2141.765 2696.815 2142.305 ;
        RECT 2701.770 2141.710 2702.120 2142.960 ;
        RECT 2703.885 2142.305 2707.395 2143.395 ;
        RECT 2705.705 2141.785 2707.395 2142.305 ;
        RECT 2708.485 2142.230 2708.775 2143.395 ;
        RECT 2708.945 2142.960 2714.290 2143.395 ;
        RECT 2714.465 2142.960 2719.810 2143.395 ;
        RECT 2719.985 2142.960 2725.330 2143.395 ;
        RECT 2725.505 2142.960 2730.850 2143.395 ;
        RECT 2712.350 2141.710 2712.700 2142.960 ;
        RECT 2717.870 2141.710 2718.220 2142.960 ;
        RECT 2723.390 2141.710 2723.740 2142.960 ;
        RECT 2728.910 2141.710 2729.260 2142.960 ;
        RECT 2731.025 2142.305 2732.695 2143.395 ;
        RECT 2731.945 2141.785 2732.695 2142.305 ;
        RECT 2732.865 2142.305 2734.075 2143.395 ;
        RECT 2732.865 2141.765 2733.385 2142.305 ;
        RECT 2696.295 2139.215 2696.815 2139.755 ;
        RECT 2695.605 2138.125 2696.815 2139.215 ;
        RECT 2700.390 2138.560 2700.740 2139.810 ;
        RECT 2705.910 2138.560 2706.260 2139.810 ;
        RECT 2711.430 2138.560 2711.780 2139.810 ;
        RECT 2716.950 2138.560 2717.300 2139.810 ;
        RECT 2719.985 2139.215 2720.735 2139.735 ;
        RECT 2696.985 2138.125 2702.330 2138.560 ;
        RECT 2702.505 2138.125 2707.850 2138.560 ;
        RECT 2708.025 2138.125 2713.370 2138.560 ;
        RECT 2713.545 2138.125 2718.890 2138.560 ;
        RECT 2719.065 2138.125 2720.735 2139.215 ;
        RECT 2721.365 2138.125 2721.655 2139.290 ;
        RECT 2725.230 2138.560 2725.580 2139.810 ;
        RECT 2730.750 2138.560 2731.100 2139.810 ;
        RECT 2732.865 2139.215 2733.385 2139.755 ;
        RECT 2721.825 2138.125 2727.170 2138.560 ;
        RECT 2727.345 2138.125 2732.690 2138.560 ;
        RECT 2732.865 2138.125 2734.075 2139.215 ;
        RECT 2695.520 2137.955 2734.160 2138.125 ;
        RECT 2695.605 2136.865 2696.815 2137.955 ;
        RECT 2697.425 2137.195 2697.755 2137.955 ;
        RECT 2698.365 2137.520 2703.710 2137.955 ;
        RECT 2522.135 2136.590 2523.935 2136.760 ;
        RECT 2522.830 2135.865 2523.160 2136.590 ;
        RECT 2696.295 2136.325 2696.815 2136.865 ;
        RECT 2701.770 2136.270 2702.120 2137.520 ;
        RECT 2703.885 2136.865 2707.395 2137.955 ;
        RECT 2705.705 2136.345 2707.395 2136.865 ;
        RECT 2708.485 2136.790 2708.775 2137.955 ;
        RECT 2708.945 2137.520 2714.290 2137.955 ;
        RECT 2714.465 2137.520 2719.810 2137.955 ;
        RECT 2719.985 2137.520 2725.330 2137.955 ;
        RECT 2725.505 2137.520 2730.850 2137.955 ;
        RECT 2712.350 2136.270 2712.700 2137.520 ;
        RECT 2717.870 2136.270 2718.220 2137.520 ;
        RECT 2723.390 2136.270 2723.740 2137.520 ;
        RECT 2728.910 2136.270 2729.260 2137.520 ;
        RECT 2731.025 2136.865 2732.695 2137.955 ;
        RECT 2731.945 2136.345 2732.695 2136.865 ;
        RECT 2732.865 2136.865 2734.075 2137.955 ;
        RECT 2732.865 2136.325 2733.385 2136.865 ;
        RECT 2696.295 2133.775 2696.815 2134.315 ;
        RECT 2695.605 2132.685 2696.815 2133.775 ;
        RECT 2700.390 2133.120 2700.740 2134.370 ;
        RECT 2705.910 2133.120 2706.260 2134.370 ;
        RECT 2711.430 2133.120 2711.780 2134.370 ;
        RECT 2716.950 2133.120 2717.300 2134.370 ;
        RECT 2719.985 2133.775 2720.735 2134.295 ;
        RECT 2696.985 2132.685 2702.330 2133.120 ;
        RECT 2702.505 2132.685 2707.850 2133.120 ;
        RECT 2708.025 2132.685 2713.370 2133.120 ;
        RECT 2713.545 2132.685 2718.890 2133.120 ;
        RECT 2719.065 2132.685 2720.735 2133.775 ;
        RECT 2721.365 2132.685 2721.655 2133.850 ;
        RECT 2725.230 2133.120 2725.580 2134.370 ;
        RECT 2730.750 2133.120 2731.100 2134.370 ;
        RECT 2732.865 2133.775 2733.385 2134.315 ;
        RECT 2721.825 2132.685 2727.170 2133.120 ;
        RECT 2727.345 2132.685 2732.690 2133.120 ;
        RECT 2732.865 2132.685 2734.075 2133.775 ;
        RECT 2695.520 2132.515 2734.160 2132.685 ;
        RECT 2695.605 2131.425 2696.815 2132.515 ;
        RECT 2697.425 2131.755 2697.755 2132.515 ;
        RECT 2698.805 2131.755 2699.135 2132.515 ;
        RECT 2699.745 2132.080 2705.090 2132.515 ;
        RECT 2696.295 2130.885 2696.815 2131.425 ;
        RECT 2703.150 2130.830 2703.500 2132.080 ;
        RECT 2705.265 2131.425 2707.855 2132.515 ;
        RECT 2706.645 2130.905 2707.855 2131.425 ;
        RECT 2708.485 2131.350 2708.775 2132.515 ;
        RECT 2708.945 2132.080 2714.290 2132.515 ;
        RECT 2714.465 2132.080 2719.810 2132.515 ;
        RECT 2712.350 2130.830 2712.700 2132.080 ;
        RECT 2717.870 2130.830 2718.220 2132.080 ;
        RECT 2719.985 2131.425 2721.195 2132.515 ;
        RECT 2720.675 2130.885 2721.195 2131.425 ;
        RECT 2721.365 2131.350 2721.655 2132.515 ;
        RECT 2721.825 2132.080 2727.170 2132.515 ;
        RECT 2727.345 2132.080 2732.690 2132.515 ;
        RECT 2725.230 2130.830 2725.580 2132.080 ;
        RECT 2730.750 2130.830 2731.100 2132.080 ;
        RECT 2732.865 2131.425 2734.075 2132.515 ;
        RECT 2732.865 2130.885 2733.385 2131.425 ;
        RECT 2522.135 2129.060 2523.935 2129.230 ;
        RECT 2522.830 2128.335 2523.160 2129.060 ;
        RECT 2522.135 2123.080 2523.935 2123.250 ;
        RECT 2522.830 2122.355 2523.160 2123.080 ;
        RECT 2522.135 2117.135 2523.935 2117.305 ;
        RECT 2522.830 2116.410 2523.160 2117.135 ;
        RECT 2522.135 2111.490 2523.935 2111.660 ;
        RECT 2522.830 2110.765 2523.160 2111.490 ;
        RECT 2522.135 2105.485 2523.935 2105.655 ;
        RECT 2522.830 2104.760 2523.160 2105.485 ;
        RECT 2360.035 2058.045 2360.210 2058.595 ;
        RECT 2360.035 2056.445 2360.205 2058.045 ;
        RECT 2358.220 2055.035 2358.390 2055.765 ;
        RECT 2360.035 2055.305 2360.210 2056.445 ;
        RECT 2360.035 2055.035 2360.205 2055.305 ;
        RECT 2366.800 2055.035 2366.970 2055.765 ;
        RECT 2372.415 2055.035 2372.585 2055.765 ;
        RECT 2375.160 2055.035 2375.330 2055.765 ;
        RECT 2358.050 2055.030 2360.800 2055.035 ;
        RECT 2366.630 2055.030 2369.380 2055.035 ;
        RECT 2372.245 2055.030 2375.980 2055.035 ;
        RECT 2376.155 2055.030 2376.325 2055.760 ;
        RECT 2383.125 2055.035 2383.295 2055.765 ;
        RECT 2388.740 2055.035 2388.910 2055.765 ;
        RECT 2391.485 2055.035 2391.655 2055.765 ;
        RECT 2382.955 2055.030 2385.705 2055.035 ;
        RECT 2388.570 2055.030 2392.305 2055.035 ;
        RECT 2392.480 2055.030 2392.650 2055.760 ;
        RECT 2399.450 2055.035 2399.620 2055.765 ;
        RECT 2405.065 2055.035 2405.235 2055.765 ;
        RECT 2407.810 2055.035 2407.980 2055.765 ;
        RECT 2399.280 2055.030 2402.030 2055.035 ;
        RECT 2404.895 2055.030 2408.630 2055.035 ;
        RECT 2408.805 2055.030 2408.975 2055.760 ;
        RECT 2415.775 2055.035 2415.945 2055.765 ;
        RECT 2421.390 2055.035 2421.560 2055.765 ;
        RECT 2424.135 2055.035 2424.305 2055.765 ;
        RECT 2415.605 2055.030 2418.355 2055.035 ;
        RECT 2421.220 2055.030 2424.955 2055.035 ;
        RECT 2425.130 2055.030 2425.300 2055.760 ;
        RECT 2432.100 2055.035 2432.270 2055.765 ;
        RECT 2437.715 2055.035 2437.885 2055.765 ;
        RECT 2440.460 2055.035 2440.630 2055.765 ;
        RECT 2431.930 2055.030 2434.680 2055.035 ;
        RECT 2437.545 2055.030 2441.280 2055.035 ;
        RECT 2441.455 2055.030 2441.625 2055.760 ;
        RECT 2343.005 2053.430 2442.425 2055.030 ;
        RECT 2361.540 2053.425 2371.200 2053.430 ;
        RECT 2372.245 2053.425 2375.980 2053.430 ;
        RECT 2362.830 2052.925 2363.000 2053.425 ;
        RECT 2365.270 2052.925 2365.440 2053.425 ;
        RECT 2366.230 2052.925 2366.400 2053.425 ;
        RECT 2367.230 2052.925 2367.400 2053.425 ;
        RECT 2369.670 2052.925 2369.840 2053.425 ;
        RECT 2370.630 2052.925 2370.800 2053.425 ;
        RECT 2372.415 2052.695 2372.585 2053.425 ;
        RECT 2375.160 2052.695 2375.330 2053.425 ;
        RECT 2376.150 2052.700 2376.320 2053.430 ;
        RECT 2377.865 2053.425 2387.525 2053.430 ;
        RECT 2388.570 2053.425 2392.305 2053.430 ;
        RECT 2379.155 2052.925 2379.325 2053.425 ;
        RECT 2381.595 2052.925 2381.765 2053.425 ;
        RECT 2382.555 2052.925 2382.725 2053.425 ;
        RECT 2383.555 2052.925 2383.725 2053.425 ;
        RECT 2385.995 2052.925 2386.165 2053.425 ;
        RECT 2386.955 2052.925 2387.125 2053.425 ;
        RECT 2388.740 2052.695 2388.910 2053.425 ;
        RECT 2391.485 2052.695 2391.655 2053.425 ;
        RECT 2392.475 2052.700 2392.645 2053.430 ;
        RECT 2394.190 2053.425 2403.850 2053.430 ;
        RECT 2404.895 2053.425 2408.630 2053.430 ;
        RECT 2395.480 2052.925 2395.650 2053.425 ;
        RECT 2397.920 2052.925 2398.090 2053.425 ;
        RECT 2398.880 2052.925 2399.050 2053.425 ;
        RECT 2399.880 2052.925 2400.050 2053.425 ;
        RECT 2402.320 2052.925 2402.490 2053.425 ;
        RECT 2403.280 2052.925 2403.450 2053.425 ;
        RECT 2405.065 2052.695 2405.235 2053.425 ;
        RECT 2407.810 2052.695 2407.980 2053.425 ;
        RECT 2408.800 2052.700 2408.970 2053.430 ;
        RECT 2410.515 2053.425 2420.175 2053.430 ;
        RECT 2421.220 2053.425 2424.955 2053.430 ;
        RECT 2411.805 2052.925 2411.975 2053.425 ;
        RECT 2414.245 2052.925 2414.415 2053.425 ;
        RECT 2415.205 2052.925 2415.375 2053.425 ;
        RECT 2416.205 2052.925 2416.375 2053.425 ;
        RECT 2418.645 2052.925 2418.815 2053.425 ;
        RECT 2419.605 2052.925 2419.775 2053.425 ;
        RECT 2421.390 2052.695 2421.560 2053.425 ;
        RECT 2424.135 2052.695 2424.305 2053.425 ;
        RECT 2425.125 2052.700 2425.295 2053.430 ;
        RECT 2426.840 2053.425 2436.500 2053.430 ;
        RECT 2437.545 2053.425 2441.280 2053.430 ;
        RECT 2428.130 2052.925 2428.300 2053.425 ;
        RECT 2430.570 2052.925 2430.740 2053.425 ;
        RECT 2431.530 2052.925 2431.700 2053.425 ;
        RECT 2432.530 2052.925 2432.700 2053.425 ;
        RECT 2434.970 2052.925 2435.140 2053.425 ;
        RECT 2435.930 2052.925 2436.100 2053.425 ;
        RECT 2437.715 2052.695 2437.885 2053.425 ;
        RECT 2440.460 2052.695 2440.630 2053.425 ;
        RECT 2441.450 2052.700 2441.620 2053.430 ;
        RECT 2696.295 2035.375 2696.815 2035.915 ;
        RECT 2695.605 2034.285 2696.815 2035.375 ;
        RECT 2697.425 2034.285 2697.755 2035.065 ;
        RECT 2698.315 2034.285 2698.650 2034.710 ;
        RECT 2699.265 2034.285 2699.595 2035.045 ;
        RECT 2700.645 2034.285 2700.975 2035.045 ;
        RECT 2704.990 2034.720 2705.340 2035.970 ;
        RECT 2707.795 2035.375 2708.315 2035.915 ;
        RECT 2701.585 2034.285 2706.930 2034.720 ;
        RECT 2707.105 2034.285 2708.315 2035.375 ;
        RECT 2708.485 2034.285 2708.775 2035.450 ;
        RECT 2709.420 2034.285 2709.750 2035.045 ;
        RECT 2710.350 2034.285 2710.610 2035.435 ;
        RECT 2714.190 2034.720 2714.540 2035.970 ;
        RECT 2718.125 2035.375 2719.815 2035.895 ;
        RECT 2720.675 2035.375 2721.195 2035.915 ;
        RECT 2710.785 2034.285 2716.130 2034.720 ;
        RECT 2716.305 2034.285 2719.815 2035.375 ;
        RECT 2719.985 2034.285 2721.195 2035.375 ;
        RECT 2721.365 2034.285 2721.655 2035.450 ;
        RECT 2721.830 2034.285 2722.165 2034.710 ;
        RECT 2722.725 2034.285 2723.055 2035.065 ;
        RECT 2727.070 2034.720 2727.420 2035.970 ;
        RECT 2730.105 2035.375 2730.855 2035.895 ;
        RECT 2723.665 2034.285 2729.010 2034.720 ;
        RECT 2729.185 2034.285 2730.855 2035.375 ;
        RECT 2732.865 2035.375 2733.385 2035.915 ;
        RECT 2731.925 2034.285 2732.255 2035.045 ;
        RECT 2732.865 2034.285 2734.075 2035.375 ;
        RECT 2695.520 2034.115 2734.160 2034.285 ;
        RECT 2695.605 2033.025 2696.815 2034.115 ;
        RECT 2697.425 2033.355 2697.755 2034.115 ;
        RECT 2698.365 2033.680 2703.710 2034.115 ;
        RECT 2696.295 2032.485 2696.815 2033.025 ;
        RECT 2701.770 2032.430 2702.120 2033.680 ;
        RECT 2703.885 2033.025 2707.395 2034.115 ;
        RECT 2705.705 2032.505 2707.395 2033.025 ;
        RECT 2708.485 2032.950 2708.775 2034.115 ;
        RECT 2708.945 2033.680 2714.290 2034.115 ;
        RECT 2714.465 2033.680 2719.810 2034.115 ;
        RECT 2719.985 2033.680 2725.330 2034.115 ;
        RECT 2725.505 2033.680 2730.850 2034.115 ;
        RECT 2712.350 2032.430 2712.700 2033.680 ;
        RECT 2717.870 2032.430 2718.220 2033.680 ;
        RECT 2723.390 2032.430 2723.740 2033.680 ;
        RECT 2728.910 2032.430 2729.260 2033.680 ;
        RECT 2731.025 2033.025 2732.695 2034.115 ;
        RECT 2731.945 2032.505 2732.695 2033.025 ;
        RECT 2732.865 2033.025 2734.075 2034.115 ;
        RECT 2732.865 2032.485 2733.385 2033.025 ;
        RECT 2696.295 2029.935 2696.815 2030.475 ;
        RECT 2695.605 2028.845 2696.815 2029.935 ;
        RECT 2700.390 2029.280 2700.740 2030.530 ;
        RECT 2705.910 2029.280 2706.260 2030.530 ;
        RECT 2711.430 2029.280 2711.780 2030.530 ;
        RECT 2716.950 2029.280 2717.300 2030.530 ;
        RECT 2719.985 2029.935 2720.735 2030.455 ;
        RECT 2696.985 2028.845 2702.330 2029.280 ;
        RECT 2702.505 2028.845 2707.850 2029.280 ;
        RECT 2708.025 2028.845 2713.370 2029.280 ;
        RECT 2713.545 2028.845 2718.890 2029.280 ;
        RECT 2719.065 2028.845 2720.735 2029.935 ;
        RECT 2721.365 2028.845 2721.655 2030.010 ;
        RECT 2725.230 2029.280 2725.580 2030.530 ;
        RECT 2730.750 2029.280 2731.100 2030.530 ;
        RECT 2732.865 2029.935 2733.385 2030.475 ;
        RECT 2721.825 2028.845 2727.170 2029.280 ;
        RECT 2727.345 2028.845 2732.690 2029.280 ;
        RECT 2732.865 2028.845 2734.075 2029.935 ;
        RECT 2695.520 2028.675 2734.160 2028.845 ;
        RECT 2695.605 2027.585 2696.815 2028.675 ;
        RECT 2696.985 2028.240 2702.330 2028.675 ;
        RECT 2702.505 2028.240 2707.850 2028.675 ;
        RECT 2696.295 2027.045 2696.815 2027.585 ;
        RECT 2700.390 2026.990 2700.740 2028.240 ;
        RECT 2705.910 2026.990 2706.260 2028.240 ;
        RECT 2708.485 2027.510 2708.775 2028.675 ;
        RECT 2708.945 2028.240 2714.290 2028.675 ;
        RECT 2714.465 2028.240 2719.810 2028.675 ;
        RECT 2719.985 2028.240 2725.330 2028.675 ;
        RECT 2725.505 2028.240 2730.850 2028.675 ;
        RECT 2712.350 2026.990 2712.700 2028.240 ;
        RECT 2717.870 2026.990 2718.220 2028.240 ;
        RECT 2723.390 2026.990 2723.740 2028.240 ;
        RECT 2728.910 2026.990 2729.260 2028.240 ;
        RECT 2731.025 2027.585 2732.695 2028.675 ;
        RECT 2731.945 2027.065 2732.695 2027.585 ;
        RECT 2732.865 2027.585 2734.075 2028.675 ;
        RECT 2732.865 2027.045 2733.385 2027.585 ;
        RECT 2696.295 2024.495 2696.815 2025.035 ;
        RECT 2695.605 2023.405 2696.815 2024.495 ;
        RECT 2697.425 2023.405 2697.755 2024.165 ;
        RECT 2701.770 2023.840 2702.120 2025.090 ;
        RECT 2707.290 2023.840 2707.640 2025.090 ;
        RECT 2712.810 2023.840 2713.160 2025.090 ;
        RECT 2718.330 2023.840 2718.680 2025.090 ;
        RECT 2698.365 2023.405 2703.710 2023.840 ;
        RECT 2703.885 2023.405 2709.230 2023.840 ;
        RECT 2709.405 2023.405 2714.750 2023.840 ;
        RECT 2714.925 2023.405 2720.270 2023.840 ;
        RECT 2721.365 2023.405 2721.655 2024.570 ;
        RECT 2725.230 2023.840 2725.580 2025.090 ;
        RECT 2730.750 2023.840 2731.100 2025.090 ;
        RECT 2732.865 2024.495 2733.385 2025.035 ;
        RECT 2721.825 2023.405 2727.170 2023.840 ;
        RECT 2727.345 2023.405 2732.690 2023.840 ;
        RECT 2732.865 2023.405 2734.075 2024.495 ;
        RECT 2695.520 2023.235 2734.160 2023.405 ;
        RECT 2695.605 2022.145 2696.815 2023.235 ;
        RECT 2696.985 2022.800 2702.330 2023.235 ;
        RECT 2702.505 2022.800 2707.850 2023.235 ;
        RECT 2696.295 2021.605 2696.815 2022.145 ;
        RECT 2700.390 2021.550 2700.740 2022.800 ;
        RECT 2705.910 2021.550 2706.260 2022.800 ;
        RECT 2708.485 2022.070 2708.775 2023.235 ;
        RECT 2708.945 2022.800 2714.290 2023.235 ;
        RECT 2714.465 2022.800 2719.810 2023.235 ;
        RECT 2719.985 2022.800 2725.330 2023.235 ;
        RECT 2725.505 2022.800 2730.850 2023.235 ;
        RECT 2712.350 2021.550 2712.700 2022.800 ;
        RECT 2717.870 2021.550 2718.220 2022.800 ;
        RECT 2723.390 2021.550 2723.740 2022.800 ;
        RECT 2728.910 2021.550 2729.260 2022.800 ;
        RECT 2731.025 2022.145 2732.695 2023.235 ;
        RECT 2731.945 2021.625 2732.695 2022.145 ;
        RECT 2732.865 2022.145 2734.075 2023.235 ;
        RECT 2732.865 2021.605 2733.385 2022.145 ;
        RECT 2696.295 2019.055 2696.815 2019.595 ;
        RECT 2695.605 2017.965 2696.815 2019.055 ;
        RECT 2710.050 2018.400 2710.400 2019.650 ;
        RECT 2715.570 2018.400 2715.920 2019.650 ;
        RECT 2719.505 2019.055 2721.195 2019.575 ;
        RECT 2697.415 2017.965 2697.745 2018.345 ;
        RECT 2700.135 2017.965 2700.465 2018.345 ;
        RECT 2701.960 2017.965 2702.290 2018.345 ;
        RECT 2702.880 2017.965 2703.230 2018.345 ;
        RECT 2705.715 2017.965 2706.045 2018.345 ;
        RECT 2706.645 2017.965 2711.990 2018.400 ;
        RECT 2712.165 2017.965 2717.510 2018.400 ;
        RECT 2717.685 2017.965 2721.195 2019.055 ;
        RECT 2721.365 2017.965 2721.655 2019.130 ;
        RECT 2725.230 2018.400 2725.580 2019.650 ;
        RECT 2730.750 2018.400 2731.100 2019.650 ;
        RECT 2732.865 2019.055 2733.385 2019.595 ;
        RECT 2721.825 2017.965 2727.170 2018.400 ;
        RECT 2727.345 2017.965 2732.690 2018.400 ;
        RECT 2732.865 2017.965 2734.075 2019.055 ;
        RECT 2695.520 2017.795 2734.160 2017.965 ;
        RECT 2695.605 2016.705 2696.815 2017.795 ;
        RECT 2697.425 2017.035 2697.755 2017.795 ;
        RECT 2698.365 2017.360 2703.710 2017.795 ;
        RECT 2696.295 2016.165 2696.815 2016.705 ;
        RECT 2701.770 2016.110 2702.120 2017.360 ;
        RECT 2703.885 2016.705 2707.395 2017.795 ;
        RECT 2705.705 2016.185 2707.395 2016.705 ;
        RECT 2708.485 2016.630 2708.775 2017.795 ;
        RECT 2708.945 2017.360 2714.290 2017.795 ;
        RECT 2714.465 2017.360 2719.810 2017.795 ;
        RECT 2719.985 2017.360 2725.330 2017.795 ;
        RECT 2725.505 2017.360 2730.850 2017.795 ;
        RECT 2712.350 2016.110 2712.700 2017.360 ;
        RECT 2717.870 2016.110 2718.220 2017.360 ;
        RECT 2723.390 2016.110 2723.740 2017.360 ;
        RECT 2728.910 2016.110 2729.260 2017.360 ;
        RECT 2731.025 2016.705 2732.695 2017.795 ;
        RECT 2731.945 2016.185 2732.695 2016.705 ;
        RECT 2732.865 2016.705 2734.075 2017.795 ;
        RECT 2732.865 2016.165 2733.385 2016.705 ;
        RECT 2696.295 2013.615 2696.815 2014.155 ;
        RECT 2695.605 2012.525 2696.815 2013.615 ;
        RECT 2710.050 2012.960 2710.400 2014.210 ;
        RECT 2715.570 2012.960 2715.920 2014.210 ;
        RECT 2719.505 2013.615 2721.195 2014.135 ;
        RECT 2697.415 2012.525 2697.745 2012.905 ;
        RECT 2700.135 2012.525 2700.465 2012.905 ;
        RECT 2701.960 2012.525 2702.290 2012.905 ;
        RECT 2702.880 2012.525 2703.230 2012.905 ;
        RECT 2705.715 2012.525 2706.045 2012.905 ;
        RECT 2706.645 2012.525 2711.990 2012.960 ;
        RECT 2712.165 2012.525 2717.510 2012.960 ;
        RECT 2717.685 2012.525 2721.195 2013.615 ;
        RECT 2721.365 2012.525 2721.655 2013.690 ;
        RECT 2725.230 2012.960 2725.580 2014.210 ;
        RECT 2730.750 2012.960 2731.100 2014.210 ;
        RECT 2732.865 2013.615 2733.385 2014.155 ;
        RECT 2721.825 2012.525 2727.170 2012.960 ;
        RECT 2727.345 2012.525 2732.690 2012.960 ;
        RECT 2732.865 2012.525 2734.075 2013.615 ;
        RECT 2695.520 2012.355 2734.160 2012.525 ;
        RECT 2695.605 2011.265 2696.815 2012.355 ;
        RECT 2697.425 2011.595 2697.755 2012.355 ;
        RECT 2698.365 2011.265 2700.955 2012.355 ;
        RECT 2696.295 2010.725 2696.815 2011.265 ;
        RECT 2699.745 2010.745 2700.955 2011.265 ;
        RECT 2702.095 2011.215 2702.265 2012.355 ;
        RECT 2704.635 2011.595 2704.805 2012.355 ;
        RECT 2705.725 2011.265 2708.315 2012.355 ;
        RECT 2707.105 2010.745 2708.315 2011.265 ;
        RECT 2708.485 2011.190 2708.775 2012.355 ;
        RECT 2708.945 2011.920 2714.290 2012.355 ;
        RECT 2714.465 2011.920 2719.810 2012.355 ;
        RECT 2719.985 2011.920 2725.330 2012.355 ;
        RECT 2725.505 2011.920 2730.850 2012.355 ;
        RECT 2712.350 2010.670 2712.700 2011.920 ;
        RECT 2717.870 2010.670 2718.220 2011.920 ;
        RECT 2723.390 2010.670 2723.740 2011.920 ;
        RECT 2728.910 2010.670 2729.260 2011.920 ;
        RECT 2731.025 2011.265 2732.695 2012.355 ;
        RECT 2731.945 2010.745 2732.695 2011.265 ;
        RECT 2732.865 2011.265 2734.075 2012.355 ;
        RECT 2732.865 2010.725 2733.385 2011.265 ;
        RECT 2696.295 2008.175 2696.815 2008.715 ;
        RECT 2695.605 2007.085 2696.815 2008.175 ;
        RECT 2700.390 2007.520 2700.740 2008.770 ;
        RECT 2705.910 2007.520 2706.260 2008.770 ;
        RECT 2711.430 2007.520 2711.780 2008.770 ;
        RECT 2716.950 2007.520 2717.300 2008.770 ;
        RECT 2719.985 2008.175 2720.735 2008.695 ;
        RECT 2696.985 2007.085 2702.330 2007.520 ;
        RECT 2702.505 2007.085 2707.850 2007.520 ;
        RECT 2708.025 2007.085 2713.370 2007.520 ;
        RECT 2713.545 2007.085 2718.890 2007.520 ;
        RECT 2719.065 2007.085 2720.735 2008.175 ;
        RECT 2721.365 2007.085 2721.655 2008.250 ;
        RECT 2725.230 2007.520 2725.580 2008.770 ;
        RECT 2730.750 2007.520 2731.100 2008.770 ;
        RECT 2732.865 2008.175 2733.385 2008.715 ;
        RECT 2721.825 2007.085 2727.170 2007.520 ;
        RECT 2727.345 2007.085 2732.690 2007.520 ;
        RECT 2732.865 2007.085 2734.075 2008.175 ;
        RECT 2695.520 2006.915 2734.160 2007.085 ;
        RECT 2695.605 2005.825 2696.815 2006.915 ;
        RECT 2697.425 2006.155 2697.755 2006.915 ;
        RECT 2698.365 2006.480 2703.710 2006.915 ;
        RECT 2696.295 2005.285 2696.815 2005.825 ;
        RECT 2701.770 2005.230 2702.120 2006.480 ;
        RECT 2703.885 2005.825 2707.395 2006.915 ;
        RECT 2705.705 2005.305 2707.395 2005.825 ;
        RECT 2708.485 2005.750 2708.775 2006.915 ;
        RECT 2708.945 2006.480 2714.290 2006.915 ;
        RECT 2714.465 2006.480 2719.810 2006.915 ;
        RECT 2719.985 2006.480 2725.330 2006.915 ;
        RECT 2725.505 2006.480 2730.850 2006.915 ;
        RECT 2712.350 2005.230 2712.700 2006.480 ;
        RECT 2717.870 2005.230 2718.220 2006.480 ;
        RECT 2723.390 2005.230 2723.740 2006.480 ;
        RECT 2728.910 2005.230 2729.260 2006.480 ;
        RECT 2731.025 2005.825 2732.695 2006.915 ;
        RECT 2731.945 2005.305 2732.695 2005.825 ;
        RECT 2732.865 2005.825 2734.075 2006.915 ;
        RECT 2732.865 2005.285 2733.385 2005.825 ;
        RECT 2696.295 2002.735 2696.815 2003.275 ;
        RECT 2695.605 2001.645 2696.815 2002.735 ;
        RECT 2700.390 2002.080 2700.740 2003.330 ;
        RECT 2705.910 2002.080 2706.260 2003.330 ;
        RECT 2711.430 2002.080 2711.780 2003.330 ;
        RECT 2716.950 2002.080 2717.300 2003.330 ;
        RECT 2719.985 2002.735 2720.735 2003.255 ;
        RECT 2696.985 2001.645 2702.330 2002.080 ;
        RECT 2702.505 2001.645 2707.850 2002.080 ;
        RECT 2708.025 2001.645 2713.370 2002.080 ;
        RECT 2713.545 2001.645 2718.890 2002.080 ;
        RECT 2719.065 2001.645 2720.735 2002.735 ;
        RECT 2721.365 2001.645 2721.655 2002.810 ;
        RECT 2725.230 2002.080 2725.580 2003.330 ;
        RECT 2730.750 2002.080 2731.100 2003.330 ;
        RECT 2732.865 2002.735 2733.385 2003.275 ;
        RECT 2721.825 2001.645 2727.170 2002.080 ;
        RECT 2727.345 2001.645 2732.690 2002.080 ;
        RECT 2732.865 2001.645 2734.075 2002.735 ;
        RECT 2695.520 2001.475 2734.160 2001.645 ;
        RECT 2695.605 2000.385 2696.815 2001.475 ;
        RECT 2696.985 2000.385 2700.495 2001.475 ;
        RECT 2696.295 1999.845 2696.815 2000.385 ;
        RECT 2698.805 1999.865 2700.495 2000.385 ;
        RECT 2702.455 2000.335 2702.785 2001.475 ;
        RECT 2702.965 2001.040 2708.310 2001.475 ;
        RECT 2706.370 1999.790 2706.720 2001.040 ;
        RECT 2708.485 2000.310 2708.775 2001.475 ;
        RECT 2708.945 2001.040 2714.290 2001.475 ;
        RECT 2714.465 2001.040 2719.810 2001.475 ;
        RECT 2719.985 2001.040 2725.330 2001.475 ;
        RECT 2725.505 2001.040 2730.850 2001.475 ;
        RECT 2712.350 1999.790 2712.700 2001.040 ;
        RECT 2717.870 1999.790 2718.220 2001.040 ;
        RECT 2723.390 1999.790 2723.740 2001.040 ;
        RECT 2728.910 1999.790 2729.260 2001.040 ;
        RECT 2731.025 2000.385 2732.695 2001.475 ;
        RECT 2731.945 1999.865 2732.695 2000.385 ;
        RECT 2732.865 2000.385 2734.075 2001.475 ;
        RECT 2732.865 1999.845 2733.385 2000.385 ;
        RECT 2696.295 1997.295 2696.815 1997.835 ;
        RECT 2700.185 1997.295 2701.875 1997.815 ;
        RECT 2695.605 1996.205 2696.815 1997.295 ;
        RECT 2697.425 1996.205 2697.755 1996.965 ;
        RECT 2698.365 1996.205 2701.875 1997.295 ;
        RECT 2703.535 1996.205 2703.705 1996.645 ;
        RECT 2708.670 1996.640 2709.020 1997.890 ;
        RECT 2714.190 1996.640 2714.540 1997.890 ;
        RECT 2718.125 1997.295 2719.815 1997.815 ;
        RECT 2720.675 1997.295 2721.195 1997.835 ;
        RECT 2704.310 1996.205 2704.640 1996.565 ;
        RECT 2705.265 1996.205 2710.610 1996.640 ;
        RECT 2710.785 1996.205 2716.130 1996.640 ;
        RECT 2716.305 1996.205 2719.815 1997.295 ;
        RECT 2719.985 1996.205 2721.195 1997.295 ;
        RECT 2721.365 1996.205 2721.655 1997.370 ;
        RECT 2725.230 1996.640 2725.580 1997.890 ;
        RECT 2730.750 1996.640 2731.100 1997.890 ;
        RECT 2732.865 1997.295 2733.385 1997.835 ;
        RECT 2721.825 1996.205 2727.170 1996.640 ;
        RECT 2727.345 1996.205 2732.690 1996.640 ;
        RECT 2732.865 1996.205 2734.075 1997.295 ;
        RECT 2695.520 1996.035 2734.160 1996.205 ;
        RECT 2695.605 1994.945 2696.815 1996.035 ;
        RECT 2696.985 1995.600 2702.330 1996.035 ;
        RECT 2702.505 1995.600 2707.850 1996.035 ;
        RECT 2696.295 1994.405 2696.815 1994.945 ;
        RECT 2700.390 1994.350 2700.740 1995.600 ;
        RECT 2705.910 1994.350 2706.260 1995.600 ;
        RECT 2708.485 1994.870 2708.775 1996.035 ;
        RECT 2708.945 1995.600 2714.290 1996.035 ;
        RECT 2714.465 1995.600 2719.810 1996.035 ;
        RECT 2719.985 1995.600 2725.330 1996.035 ;
        RECT 2712.350 1994.350 2712.700 1995.600 ;
        RECT 2717.870 1994.350 2718.220 1995.600 ;
        RECT 2723.390 1994.350 2723.740 1995.600 ;
        RECT 2725.595 1995.235 2725.765 1996.035 ;
        RECT 2726.435 1995.235 2726.605 1996.035 ;
        RECT 2727.275 1995.235 2727.445 1996.035 ;
        RECT 2728.035 1995.235 2728.365 1996.035 ;
        RECT 2728.875 1995.235 2729.205 1996.035 ;
        RECT 2729.715 1995.235 2730.045 1996.035 ;
        RECT 2730.555 1995.235 2730.885 1996.035 ;
        RECT 2731.395 1995.235 2731.725 1996.035 ;
        RECT 2732.235 1994.885 2732.565 1996.035 ;
        RECT 2732.865 1994.945 2734.075 1996.035 ;
        RECT 2732.865 1994.405 2733.385 1994.945 ;
        RECT 2696.295 1991.855 2696.815 1992.395 ;
        RECT 2695.605 1990.765 2696.815 1991.855 ;
        RECT 2697.425 1990.765 2697.755 1991.525 ;
        RECT 2701.770 1991.200 2702.120 1992.450 ;
        RECT 2707.290 1991.200 2707.640 1992.450 ;
        RECT 2712.810 1991.200 2713.160 1992.450 ;
        RECT 2718.330 1991.200 2718.680 1992.450 ;
        RECT 2698.365 1990.765 2703.710 1991.200 ;
        RECT 2703.885 1990.765 2709.230 1991.200 ;
        RECT 2709.405 1990.765 2714.750 1991.200 ;
        RECT 2714.925 1990.765 2720.270 1991.200 ;
        RECT 2721.365 1990.765 2721.655 1991.930 ;
        RECT 2725.230 1991.200 2725.580 1992.450 ;
        RECT 2730.750 1991.200 2731.100 1992.450 ;
        RECT 2732.865 1991.855 2733.385 1992.395 ;
        RECT 2721.825 1990.765 2727.170 1991.200 ;
        RECT 2727.345 1990.765 2732.690 1991.200 ;
        RECT 2732.865 1990.765 2734.075 1991.855 ;
        RECT 2695.520 1990.595 2734.160 1990.765 ;
        RECT 2695.605 1989.505 2696.815 1990.595 ;
        RECT 2696.985 1990.160 2702.330 1990.595 ;
        RECT 2702.505 1990.160 2707.850 1990.595 ;
        RECT 2696.295 1988.965 2696.815 1989.505 ;
        RECT 2700.390 1988.910 2700.740 1990.160 ;
        RECT 2705.910 1988.910 2706.260 1990.160 ;
        RECT 2708.485 1989.430 2708.775 1990.595 ;
        RECT 2708.945 1990.160 2714.290 1990.595 ;
        RECT 2714.465 1990.160 2719.810 1990.595 ;
        RECT 2719.985 1990.160 2725.330 1990.595 ;
        RECT 2725.505 1990.160 2730.850 1990.595 ;
        RECT 2712.350 1988.910 2712.700 1990.160 ;
        RECT 2717.870 1988.910 2718.220 1990.160 ;
        RECT 2723.390 1988.910 2723.740 1990.160 ;
        RECT 2728.910 1988.910 2729.260 1990.160 ;
        RECT 2731.025 1989.505 2732.695 1990.595 ;
        RECT 2731.945 1988.985 2732.695 1989.505 ;
        RECT 2732.865 1989.505 2734.075 1990.595 ;
        RECT 2732.865 1988.965 2733.385 1989.505 ;
        RECT 2696.295 1986.415 2696.815 1986.955 ;
        RECT 2695.605 1985.325 2696.815 1986.415 ;
        RECT 2697.715 1985.325 2698.045 1985.835 ;
        RECT 2703.150 1985.760 2703.500 1987.010 ;
        RECT 2708.670 1985.760 2709.020 1987.010 ;
        RECT 2714.190 1985.760 2714.540 1987.010 ;
        RECT 2718.125 1986.415 2719.815 1986.935 ;
        RECT 2720.675 1986.415 2721.195 1986.955 ;
        RECT 2699.745 1985.325 2705.090 1985.760 ;
        RECT 2705.265 1985.325 2710.610 1985.760 ;
        RECT 2710.785 1985.325 2716.130 1985.760 ;
        RECT 2716.305 1985.325 2719.815 1986.415 ;
        RECT 2719.985 1985.325 2721.195 1986.415 ;
        RECT 2721.365 1985.325 2721.655 1986.490 ;
        RECT 2725.230 1985.760 2725.580 1987.010 ;
        RECT 2730.750 1985.760 2731.100 1987.010 ;
        RECT 2732.865 1986.415 2733.385 1986.955 ;
        RECT 2721.825 1985.325 2727.170 1985.760 ;
        RECT 2727.345 1985.325 2732.690 1985.760 ;
        RECT 2732.865 1985.325 2734.075 1986.415 ;
        RECT 2695.520 1985.155 2734.160 1985.325 ;
        RECT 2522.135 1984.335 2523.935 1984.505 ;
        RECT 2522.830 1983.610 2523.160 1984.335 ;
        RECT 2695.605 1984.065 2696.815 1985.155 ;
        RECT 2697.425 1984.395 2697.755 1985.155 ;
        RECT 2698.365 1984.720 2703.710 1985.155 ;
        RECT 2696.295 1983.525 2696.815 1984.065 ;
        RECT 2701.770 1983.470 2702.120 1984.720 ;
        RECT 2703.885 1984.065 2707.395 1985.155 ;
        RECT 2705.705 1983.545 2707.395 1984.065 ;
        RECT 2708.485 1983.990 2708.775 1985.155 ;
        RECT 2708.945 1984.720 2714.290 1985.155 ;
        RECT 2714.465 1984.720 2719.810 1985.155 ;
        RECT 2719.985 1984.720 2725.330 1985.155 ;
        RECT 2725.505 1984.720 2730.850 1985.155 ;
        RECT 2712.350 1983.470 2712.700 1984.720 ;
        RECT 2717.870 1983.470 2718.220 1984.720 ;
        RECT 2723.390 1983.470 2723.740 1984.720 ;
        RECT 2728.910 1983.470 2729.260 1984.720 ;
        RECT 2731.025 1984.065 2732.695 1985.155 ;
        RECT 2731.945 1983.545 2732.695 1984.065 ;
        RECT 2732.865 1984.065 2734.075 1985.155 ;
        RECT 2732.865 1983.525 2733.385 1984.065 ;
        RECT 2696.295 1980.975 2696.815 1981.515 ;
        RECT 2695.605 1979.885 2696.815 1980.975 ;
        RECT 2697.735 1979.885 2697.905 1980.645 ;
        RECT 2700.275 1979.885 2700.445 1981.025 ;
        RECT 2701.590 1979.885 2701.920 1980.600 ;
        RECT 2708.210 1980.320 2708.560 1981.570 ;
        RECT 2713.730 1980.320 2714.080 1981.570 ;
        RECT 2719.250 1980.320 2719.600 1981.570 ;
        RECT 2704.805 1979.885 2710.150 1980.320 ;
        RECT 2710.325 1979.885 2715.670 1980.320 ;
        RECT 2715.845 1979.885 2721.190 1980.320 ;
        RECT 2721.365 1979.885 2721.655 1981.050 ;
        RECT 2725.230 1980.320 2725.580 1981.570 ;
        RECT 2730.750 1980.320 2731.100 1981.570 ;
        RECT 2732.865 1980.975 2733.385 1981.515 ;
        RECT 2721.825 1979.885 2727.170 1980.320 ;
        RECT 2727.345 1979.885 2732.690 1980.320 ;
        RECT 2732.865 1979.885 2734.075 1980.975 ;
        RECT 2695.520 1979.715 2734.160 1979.885 ;
        RECT 2695.605 1978.625 2696.815 1979.715 ;
        RECT 2696.985 1979.205 2697.245 1979.715 ;
        RECT 2697.905 1979.210 2698.520 1979.715 ;
        RECT 2698.325 1979.035 2698.520 1979.210 ;
        RECT 2699.335 1979.170 2699.550 1979.715 ;
        RECT 2700.205 1979.280 2705.550 1979.715 ;
        RECT 2698.325 1978.845 2698.655 1979.035 ;
        RECT 2696.295 1978.085 2696.815 1978.625 ;
        RECT 2703.610 1978.030 2703.960 1979.280 ;
        RECT 2705.725 1978.625 2708.315 1979.715 ;
        RECT 2707.105 1978.105 2708.315 1978.625 ;
        RECT 2708.485 1978.550 2708.775 1979.715 ;
        RECT 2708.945 1979.280 2714.290 1979.715 ;
        RECT 2714.465 1979.280 2719.810 1979.715 ;
        RECT 2719.985 1979.280 2725.330 1979.715 ;
        RECT 2725.505 1979.280 2730.850 1979.715 ;
        RECT 2712.350 1978.030 2712.700 1979.280 ;
        RECT 2717.870 1978.030 2718.220 1979.280 ;
        RECT 2723.390 1978.030 2723.740 1979.280 ;
        RECT 2728.910 1978.030 2729.260 1979.280 ;
        RECT 2731.025 1978.625 2732.695 1979.715 ;
        RECT 2731.945 1978.105 2732.695 1978.625 ;
        RECT 2732.865 1978.625 2734.075 1979.715 ;
        RECT 2732.865 1978.085 2733.385 1978.625 ;
        RECT 2522.135 1976.805 2523.935 1976.975 ;
        RECT 2522.830 1976.080 2523.160 1976.805 ;
        RECT 2696.295 1975.535 2696.815 1976.075 ;
        RECT 2695.605 1974.445 2696.815 1975.535 ;
        RECT 2697.425 1974.445 2697.755 1975.205 ;
        RECT 2701.770 1974.880 2702.120 1976.130 ;
        RECT 2707.290 1974.880 2707.640 1976.130 ;
        RECT 2712.810 1974.880 2713.160 1976.130 ;
        RECT 2718.330 1974.880 2718.680 1976.130 ;
        RECT 2698.365 1974.445 2703.710 1974.880 ;
        RECT 2703.885 1974.445 2709.230 1974.880 ;
        RECT 2709.405 1974.445 2714.750 1974.880 ;
        RECT 2714.925 1974.445 2720.270 1974.880 ;
        RECT 2721.365 1974.445 2721.655 1975.610 ;
        RECT 2725.230 1974.880 2725.580 1976.130 ;
        RECT 2730.750 1974.880 2731.100 1976.130 ;
        RECT 2732.865 1975.535 2733.385 1976.075 ;
        RECT 2721.825 1974.445 2727.170 1974.880 ;
        RECT 2727.345 1974.445 2732.690 1974.880 ;
        RECT 2732.865 1974.445 2734.075 1975.535 ;
        RECT 2695.520 1974.275 2734.160 1974.445 ;
        RECT 2695.605 1973.185 2696.815 1974.275 ;
        RECT 2696.985 1973.185 2698.195 1974.275 ;
        RECT 2698.865 1973.815 2699.115 1974.275 ;
        RECT 2699.795 1973.815 2700.045 1974.275 ;
        RECT 2701.115 1973.815 2701.365 1974.275 ;
        RECT 2702.045 1973.840 2707.390 1974.275 ;
        RECT 2696.295 1972.645 2696.815 1973.185 ;
        RECT 2697.675 1972.645 2698.195 1973.185 ;
        RECT 2705.450 1972.590 2705.800 1973.840 ;
        RECT 2708.485 1973.110 2708.775 1974.275 ;
        RECT 2708.945 1973.840 2714.290 1974.275 ;
        RECT 2714.465 1973.840 2719.810 1974.275 ;
        RECT 2719.985 1973.840 2725.330 1974.275 ;
        RECT 2725.505 1973.840 2730.850 1974.275 ;
        RECT 2712.350 1972.590 2712.700 1973.840 ;
        RECT 2717.870 1972.590 2718.220 1973.840 ;
        RECT 2723.390 1972.590 2723.740 1973.840 ;
        RECT 2728.910 1972.590 2729.260 1973.840 ;
        RECT 2731.025 1973.185 2732.695 1974.275 ;
        RECT 2731.945 1972.665 2732.695 1973.185 ;
        RECT 2732.865 1973.185 2734.075 1974.275 ;
        RECT 2732.865 1972.645 2733.385 1973.185 ;
        RECT 2522.135 1970.825 2523.935 1970.995 ;
        RECT 2522.830 1970.100 2523.160 1970.825 ;
        RECT 2696.295 1970.095 2696.815 1970.635 ;
        RECT 2695.605 1969.005 2696.815 1970.095 ;
        RECT 2697.905 1969.005 2698.165 1970.145 ;
        RECT 2700.190 1969.005 2700.470 1969.805 ;
        RECT 2701.885 1969.005 2702.170 1969.805 ;
        RECT 2702.840 1969.005 2703.090 1970.145 ;
        RECT 2707.290 1969.440 2707.640 1970.690 ;
        RECT 2712.810 1969.440 2713.160 1970.690 ;
        RECT 2718.330 1969.440 2718.680 1970.690 ;
        RECT 2703.885 1969.005 2709.230 1969.440 ;
        RECT 2709.405 1969.005 2714.750 1969.440 ;
        RECT 2714.925 1969.005 2720.270 1969.440 ;
        RECT 2721.365 1969.005 2721.655 1970.170 ;
        RECT 2725.230 1969.440 2725.580 1970.690 ;
        RECT 2730.750 1969.440 2731.100 1970.690 ;
        RECT 2732.865 1970.095 2733.385 1970.635 ;
        RECT 2721.825 1969.005 2727.170 1969.440 ;
        RECT 2727.345 1969.005 2732.690 1969.440 ;
        RECT 2732.865 1969.005 2734.075 1970.095 ;
        RECT 2695.520 1968.835 2734.160 1969.005 ;
        RECT 2695.605 1967.745 2696.815 1968.835 ;
        RECT 2697.425 1968.075 2697.755 1968.835 ;
        RECT 2696.295 1967.205 2696.815 1967.745 ;
        RECT 2698.825 1967.695 2699.085 1968.835 ;
        RECT 2699.755 1967.695 2700.035 1968.835 ;
        RECT 2700.205 1968.400 2705.550 1968.835 ;
        RECT 2703.610 1967.150 2703.960 1968.400 ;
        RECT 2705.725 1967.745 2708.315 1968.835 ;
        RECT 2707.105 1967.225 2708.315 1967.745 ;
        RECT 2708.485 1967.670 2708.775 1968.835 ;
        RECT 2708.945 1968.400 2714.290 1968.835 ;
        RECT 2714.465 1968.400 2719.810 1968.835 ;
        RECT 2719.985 1968.400 2725.330 1968.835 ;
        RECT 2725.505 1968.400 2730.850 1968.835 ;
        RECT 2712.350 1967.150 2712.700 1968.400 ;
        RECT 2717.870 1967.150 2718.220 1968.400 ;
        RECT 2723.390 1967.150 2723.740 1968.400 ;
        RECT 2728.910 1967.150 2729.260 1968.400 ;
        RECT 2731.025 1967.745 2732.695 1968.835 ;
        RECT 2731.945 1967.225 2732.695 1967.745 ;
        RECT 2732.865 1967.745 2734.075 1968.835 ;
        RECT 2732.865 1967.205 2733.385 1967.745 ;
        RECT 2522.135 1964.880 2523.935 1965.050 ;
        RECT 2522.830 1964.155 2523.160 1964.880 ;
        RECT 2696.295 1964.655 2696.815 1965.195 ;
        RECT 2695.605 1963.565 2696.815 1964.655 ;
        RECT 2697.735 1963.565 2697.905 1964.325 ;
        RECT 2700.275 1963.565 2700.445 1964.705 ;
        RECT 2704.530 1964.000 2704.880 1965.250 ;
        RECT 2710.050 1964.000 2710.400 1965.250 ;
        RECT 2715.570 1964.000 2715.920 1965.250 ;
        RECT 2719.505 1964.655 2721.195 1965.175 ;
        RECT 2701.125 1963.565 2706.470 1964.000 ;
        RECT 2706.645 1963.565 2711.990 1964.000 ;
        RECT 2712.165 1963.565 2717.510 1964.000 ;
        RECT 2717.685 1963.565 2721.195 1964.655 ;
        RECT 2721.365 1963.565 2721.655 1964.730 ;
        RECT 2725.230 1964.000 2725.580 1965.250 ;
        RECT 2730.750 1964.000 2731.100 1965.250 ;
        RECT 2732.865 1964.655 2733.385 1965.195 ;
        RECT 2721.825 1963.565 2727.170 1964.000 ;
        RECT 2727.345 1963.565 2732.690 1964.000 ;
        RECT 2732.865 1963.565 2734.075 1964.655 ;
        RECT 2695.520 1963.395 2734.160 1963.565 ;
        RECT 2695.605 1962.305 2696.815 1963.395 ;
        RECT 2697.425 1962.635 2697.755 1963.395 ;
        RECT 2698.365 1962.960 2703.710 1963.395 ;
        RECT 2696.295 1961.765 2696.815 1962.305 ;
        RECT 2701.770 1961.710 2702.120 1962.960 ;
        RECT 2703.885 1962.305 2707.395 1963.395 ;
        RECT 2705.705 1961.785 2707.395 1962.305 ;
        RECT 2708.485 1962.230 2708.775 1963.395 ;
        RECT 2708.945 1962.960 2714.290 1963.395 ;
        RECT 2714.465 1962.960 2719.810 1963.395 ;
        RECT 2719.985 1962.960 2725.330 1963.395 ;
        RECT 2725.505 1962.960 2730.850 1963.395 ;
        RECT 2712.350 1961.710 2712.700 1962.960 ;
        RECT 2717.870 1961.710 2718.220 1962.960 ;
        RECT 2723.390 1961.710 2723.740 1962.960 ;
        RECT 2728.910 1961.710 2729.260 1962.960 ;
        RECT 2731.025 1962.305 2732.695 1963.395 ;
        RECT 2731.945 1961.785 2732.695 1962.305 ;
        RECT 2732.865 1962.305 2734.075 1963.395 ;
        RECT 2732.865 1961.765 2733.385 1962.305 ;
        RECT 2522.135 1959.235 2523.935 1959.405 ;
        RECT 2522.830 1958.510 2523.160 1959.235 ;
        RECT 2696.295 1959.215 2696.815 1959.755 ;
        RECT 2695.605 1958.125 2696.815 1959.215 ;
        RECT 2700.390 1958.560 2700.740 1959.810 ;
        RECT 2705.910 1958.560 2706.260 1959.810 ;
        RECT 2711.430 1958.560 2711.780 1959.810 ;
        RECT 2716.950 1958.560 2717.300 1959.810 ;
        RECT 2719.985 1959.215 2720.735 1959.735 ;
        RECT 2696.985 1958.125 2702.330 1958.560 ;
        RECT 2702.505 1958.125 2707.850 1958.560 ;
        RECT 2708.025 1958.125 2713.370 1958.560 ;
        RECT 2713.545 1958.125 2718.890 1958.560 ;
        RECT 2719.065 1958.125 2720.735 1959.215 ;
        RECT 2721.365 1958.125 2721.655 1959.290 ;
        RECT 2725.230 1958.560 2725.580 1959.810 ;
        RECT 2730.750 1958.560 2731.100 1959.810 ;
        RECT 2732.865 1959.215 2733.385 1959.755 ;
        RECT 2721.825 1958.125 2727.170 1958.560 ;
        RECT 2727.345 1958.125 2732.690 1958.560 ;
        RECT 2732.865 1958.125 2734.075 1959.215 ;
        RECT 2695.520 1957.955 2734.160 1958.125 ;
        RECT 2695.605 1956.865 2696.815 1957.955 ;
        RECT 2697.425 1957.195 2697.755 1957.955 ;
        RECT 2698.365 1957.520 2703.710 1957.955 ;
        RECT 2696.295 1956.325 2696.815 1956.865 ;
        RECT 2701.770 1956.270 2702.120 1957.520 ;
        RECT 2703.885 1956.865 2707.395 1957.955 ;
        RECT 2705.705 1956.345 2707.395 1956.865 ;
        RECT 2708.485 1956.790 2708.775 1957.955 ;
        RECT 2708.945 1957.520 2714.290 1957.955 ;
        RECT 2714.465 1957.520 2719.810 1957.955 ;
        RECT 2719.985 1957.520 2725.330 1957.955 ;
        RECT 2725.505 1957.520 2730.850 1957.955 ;
        RECT 2712.350 1956.270 2712.700 1957.520 ;
        RECT 2717.870 1956.270 2718.220 1957.520 ;
        RECT 2723.390 1956.270 2723.740 1957.520 ;
        RECT 2728.910 1956.270 2729.260 1957.520 ;
        RECT 2731.025 1956.865 2732.695 1957.955 ;
        RECT 2731.945 1956.345 2732.695 1956.865 ;
        RECT 2732.865 1956.865 2734.075 1957.955 ;
        RECT 2732.865 1956.325 2733.385 1956.865 ;
        RECT 2696.295 1953.775 2696.815 1954.315 ;
        RECT 2360.035 1953.050 2360.210 1953.600 ;
        RECT 2522.135 1953.230 2523.935 1953.400 ;
        RECT 2360.035 1951.450 2360.205 1953.050 ;
        RECT 2522.830 1952.505 2523.160 1953.230 ;
        RECT 2695.605 1952.685 2696.815 1953.775 ;
        RECT 2700.390 1953.120 2700.740 1954.370 ;
        RECT 2705.910 1953.120 2706.260 1954.370 ;
        RECT 2711.430 1953.120 2711.780 1954.370 ;
        RECT 2716.950 1953.120 2717.300 1954.370 ;
        RECT 2719.985 1953.775 2720.735 1954.295 ;
        RECT 2696.985 1952.685 2702.330 1953.120 ;
        RECT 2702.505 1952.685 2707.850 1953.120 ;
        RECT 2708.025 1952.685 2713.370 1953.120 ;
        RECT 2713.545 1952.685 2718.890 1953.120 ;
        RECT 2719.065 1952.685 2720.735 1953.775 ;
        RECT 2721.365 1952.685 2721.655 1953.850 ;
        RECT 2725.230 1953.120 2725.580 1954.370 ;
        RECT 2730.750 1953.120 2731.100 1954.370 ;
        RECT 2732.865 1953.775 2733.385 1954.315 ;
        RECT 2721.825 1952.685 2727.170 1953.120 ;
        RECT 2727.345 1952.685 2732.690 1953.120 ;
        RECT 2732.865 1952.685 2734.075 1953.775 ;
        RECT 2695.520 1952.515 2734.160 1952.685 ;
        RECT 2358.220 1950.050 2358.390 1950.770 ;
        RECT 2360.035 1950.310 2360.210 1951.450 ;
        RECT 2695.605 1951.425 2696.815 1952.515 ;
        RECT 2697.425 1951.755 2697.755 1952.515 ;
        RECT 2698.805 1951.755 2699.135 1952.515 ;
        RECT 2699.745 1952.080 2705.090 1952.515 ;
        RECT 2696.295 1950.885 2696.815 1951.425 ;
        RECT 2703.150 1950.830 2703.500 1952.080 ;
        RECT 2705.265 1951.425 2707.855 1952.515 ;
        RECT 2706.645 1950.905 2707.855 1951.425 ;
        RECT 2708.485 1951.350 2708.775 1952.515 ;
        RECT 2708.945 1952.080 2714.290 1952.515 ;
        RECT 2714.465 1952.080 2719.810 1952.515 ;
        RECT 2712.350 1950.830 2712.700 1952.080 ;
        RECT 2717.870 1950.830 2718.220 1952.080 ;
        RECT 2719.985 1951.425 2721.195 1952.515 ;
        RECT 2720.675 1950.885 2721.195 1951.425 ;
        RECT 2721.365 1951.350 2721.655 1952.515 ;
        RECT 2721.825 1952.080 2727.170 1952.515 ;
        RECT 2727.345 1952.080 2732.690 1952.515 ;
        RECT 2725.230 1950.830 2725.580 1952.080 ;
        RECT 2730.750 1950.830 2731.100 1952.080 ;
        RECT 2732.865 1951.425 2734.075 1952.515 ;
        RECT 2732.865 1950.885 2733.385 1951.425 ;
        RECT 2360.035 1950.050 2360.205 1950.310 ;
        RECT 2369.035 1950.050 2369.205 1950.770 ;
        RECT 2374.650 1950.050 2374.820 1950.770 ;
        RECT 2377.395 1950.050 2377.565 1950.765 ;
        RECT 2378.385 1950.050 2378.555 1950.765 ;
        RECT 2387.595 1950.050 2387.765 1950.770 ;
        RECT 2393.210 1950.050 2393.380 1950.770 ;
        RECT 2395.955 1950.050 2396.125 1950.765 ;
        RECT 2396.945 1950.050 2397.115 1950.765 ;
        RECT 2406.155 1950.050 2406.325 1950.770 ;
        RECT 2411.770 1950.050 2411.940 1950.770 ;
        RECT 2414.515 1950.050 2414.685 1950.765 ;
        RECT 2415.505 1950.050 2415.675 1950.765 ;
        RECT 2424.715 1950.050 2424.885 1950.770 ;
        RECT 2430.330 1950.050 2430.500 1950.770 ;
        RECT 2433.075 1950.050 2433.245 1950.765 ;
        RECT 2434.065 1950.050 2434.235 1950.765 ;
        RECT 2443.275 1950.050 2443.445 1950.770 ;
        RECT 2448.890 1950.050 2449.060 1950.770 ;
        RECT 2451.635 1950.050 2451.805 1950.765 ;
        RECT 2452.625 1950.050 2452.795 1950.765 ;
        RECT 2343.000 1948.450 2453.600 1950.050 ;
        RECT 2360.800 1948.435 2453.600 1948.450 ;
        RECT 2361.545 1948.430 2379.360 1948.435 ;
        RECT 2380.105 1948.430 2397.920 1948.435 ;
        RECT 2398.665 1948.430 2416.480 1948.435 ;
        RECT 2417.225 1948.430 2435.040 1948.435 ;
        RECT 2435.785 1948.430 2453.600 1948.435 ;
        RECT 2361.545 1948.425 2373.505 1948.430 ;
        RECT 2374.480 1948.425 2377.565 1948.430 ;
        RECT 2362.355 1947.925 2362.525 1948.425 ;
        RECT 2363.315 1947.925 2363.485 1948.425 ;
        RECT 2364.315 1947.925 2364.485 1948.425 ;
        RECT 2366.275 1947.925 2366.445 1948.425 ;
        RECT 2367.235 1947.925 2367.405 1948.425 ;
        RECT 2369.195 1947.925 2369.365 1948.425 ;
        RECT 2371.635 1947.925 2371.805 1948.425 ;
        RECT 2374.650 1947.695 2374.820 1948.425 ;
        RECT 2377.395 1947.700 2377.565 1948.425 ;
        RECT 2378.380 1947.700 2378.550 1948.430 ;
        RECT 2380.105 1948.425 2392.065 1948.430 ;
        RECT 2393.040 1948.425 2396.125 1948.430 ;
        RECT 2380.915 1947.925 2381.085 1948.425 ;
        RECT 2381.875 1947.925 2382.045 1948.425 ;
        RECT 2382.875 1947.925 2383.045 1948.425 ;
        RECT 2384.835 1947.925 2385.005 1948.425 ;
        RECT 2385.795 1947.925 2385.965 1948.425 ;
        RECT 2387.755 1947.925 2387.925 1948.425 ;
        RECT 2390.195 1947.925 2390.365 1948.425 ;
        RECT 2393.210 1947.695 2393.380 1948.425 ;
        RECT 2395.955 1947.700 2396.125 1948.425 ;
        RECT 2396.940 1947.700 2397.110 1948.430 ;
        RECT 2398.665 1948.425 2410.625 1948.430 ;
        RECT 2411.600 1948.425 2414.685 1948.430 ;
        RECT 2399.475 1947.925 2399.645 1948.425 ;
        RECT 2400.435 1947.925 2400.605 1948.425 ;
        RECT 2401.435 1947.925 2401.605 1948.425 ;
        RECT 2403.395 1947.925 2403.565 1948.425 ;
        RECT 2404.355 1947.925 2404.525 1948.425 ;
        RECT 2406.315 1947.925 2406.485 1948.425 ;
        RECT 2408.755 1947.925 2408.925 1948.425 ;
        RECT 2411.770 1947.695 2411.940 1948.425 ;
        RECT 2414.515 1947.700 2414.685 1948.425 ;
        RECT 2415.500 1947.700 2415.670 1948.430 ;
        RECT 2417.225 1948.425 2429.185 1948.430 ;
        RECT 2430.160 1948.425 2433.245 1948.430 ;
        RECT 2418.035 1947.925 2418.205 1948.425 ;
        RECT 2418.995 1947.925 2419.165 1948.425 ;
        RECT 2419.995 1947.925 2420.165 1948.425 ;
        RECT 2421.955 1947.925 2422.125 1948.425 ;
        RECT 2422.915 1947.925 2423.085 1948.425 ;
        RECT 2424.875 1947.925 2425.045 1948.425 ;
        RECT 2427.315 1947.925 2427.485 1948.425 ;
        RECT 2430.330 1947.695 2430.500 1948.425 ;
        RECT 2433.075 1947.700 2433.245 1948.425 ;
        RECT 2434.060 1947.700 2434.230 1948.430 ;
        RECT 2435.785 1948.425 2447.745 1948.430 ;
        RECT 2448.720 1948.425 2451.805 1948.430 ;
        RECT 2436.595 1947.925 2436.765 1948.425 ;
        RECT 2437.555 1947.925 2437.725 1948.425 ;
        RECT 2438.555 1947.925 2438.725 1948.425 ;
        RECT 2440.515 1947.925 2440.685 1948.425 ;
        RECT 2441.475 1947.925 2441.645 1948.425 ;
        RECT 2443.435 1947.925 2443.605 1948.425 ;
        RECT 2445.875 1947.925 2446.045 1948.425 ;
        RECT 2448.890 1947.695 2449.060 1948.425 ;
        RECT 2451.635 1947.700 2451.805 1948.425 ;
        RECT 2452.620 1947.700 2452.790 1948.430 ;
        RECT 2881.580 1894.220 2883.380 1894.390 ;
        RECT 2882.775 1893.495 2883.105 1894.220 ;
        RECT 2696.295 1855.375 2696.815 1855.915 ;
        RECT 2695.605 1854.285 2696.815 1855.375 ;
        RECT 2697.425 1854.285 2697.755 1855.065 ;
        RECT 2698.315 1854.285 2698.650 1854.710 ;
        RECT 2699.265 1854.285 2699.595 1855.045 ;
        RECT 2700.645 1854.285 2700.975 1855.045 ;
        RECT 2704.990 1854.720 2705.340 1855.970 ;
        RECT 2707.795 1855.375 2708.315 1855.915 ;
        RECT 2701.585 1854.285 2706.930 1854.720 ;
        RECT 2707.105 1854.285 2708.315 1855.375 ;
        RECT 2708.485 1854.285 2708.775 1855.450 ;
        RECT 2709.420 1854.285 2709.750 1855.045 ;
        RECT 2710.350 1854.285 2710.610 1855.435 ;
        RECT 2714.190 1854.720 2714.540 1855.970 ;
        RECT 2718.125 1855.375 2719.815 1855.895 ;
        RECT 2720.675 1855.375 2721.195 1855.915 ;
        RECT 2710.785 1854.285 2716.130 1854.720 ;
        RECT 2716.305 1854.285 2719.815 1855.375 ;
        RECT 2719.985 1854.285 2721.195 1855.375 ;
        RECT 2721.365 1854.285 2721.655 1855.450 ;
        RECT 2721.830 1854.285 2722.165 1854.710 ;
        RECT 2722.725 1854.285 2723.055 1855.065 ;
        RECT 2727.070 1854.720 2727.420 1855.970 ;
        RECT 2730.105 1855.375 2730.855 1855.895 ;
        RECT 2723.665 1854.285 2729.010 1854.720 ;
        RECT 2729.185 1854.285 2730.855 1855.375 ;
        RECT 2732.865 1855.375 2733.385 1855.915 ;
        RECT 2731.925 1854.285 2732.255 1855.045 ;
        RECT 2732.865 1854.285 2734.075 1855.375 ;
        RECT 2695.520 1854.115 2734.160 1854.285 ;
        RECT 2695.605 1853.025 2696.815 1854.115 ;
        RECT 2697.425 1853.355 2697.755 1854.115 ;
        RECT 2698.365 1853.680 2703.710 1854.115 ;
        RECT 2696.295 1852.485 2696.815 1853.025 ;
        RECT 2701.770 1852.430 2702.120 1853.680 ;
        RECT 2703.885 1853.025 2707.395 1854.115 ;
        RECT 2705.705 1852.505 2707.395 1853.025 ;
        RECT 2708.485 1852.950 2708.775 1854.115 ;
        RECT 2708.945 1853.680 2714.290 1854.115 ;
        RECT 2714.465 1853.680 2719.810 1854.115 ;
        RECT 2719.985 1853.680 2725.330 1854.115 ;
        RECT 2725.505 1853.680 2730.850 1854.115 ;
        RECT 2712.350 1852.430 2712.700 1853.680 ;
        RECT 2717.870 1852.430 2718.220 1853.680 ;
        RECT 2723.390 1852.430 2723.740 1853.680 ;
        RECT 2728.910 1852.430 2729.260 1853.680 ;
        RECT 2731.025 1853.025 2732.695 1854.115 ;
        RECT 2731.945 1852.505 2732.695 1853.025 ;
        RECT 2732.865 1853.025 2734.075 1854.115 ;
        RECT 2732.865 1852.485 2733.385 1853.025 ;
        RECT 2696.295 1849.935 2696.815 1850.475 ;
        RECT 2695.605 1848.845 2696.815 1849.935 ;
        RECT 2700.390 1849.280 2700.740 1850.530 ;
        RECT 2705.910 1849.280 2706.260 1850.530 ;
        RECT 2711.430 1849.280 2711.780 1850.530 ;
        RECT 2716.950 1849.280 2717.300 1850.530 ;
        RECT 2719.985 1849.935 2720.735 1850.455 ;
        RECT 2696.985 1848.845 2702.330 1849.280 ;
        RECT 2702.505 1848.845 2707.850 1849.280 ;
        RECT 2708.025 1848.845 2713.370 1849.280 ;
        RECT 2713.545 1848.845 2718.890 1849.280 ;
        RECT 2719.065 1848.845 2720.735 1849.935 ;
        RECT 2721.365 1848.845 2721.655 1850.010 ;
        RECT 2725.230 1849.280 2725.580 1850.530 ;
        RECT 2730.750 1849.280 2731.100 1850.530 ;
        RECT 2732.865 1849.935 2733.385 1850.475 ;
        RECT 2721.825 1848.845 2727.170 1849.280 ;
        RECT 2727.345 1848.845 2732.690 1849.280 ;
        RECT 2732.865 1848.845 2734.075 1849.935 ;
        RECT 2695.520 1848.675 2734.160 1848.845 ;
        RECT 2695.605 1847.585 2696.815 1848.675 ;
        RECT 2696.985 1848.240 2702.330 1848.675 ;
        RECT 2702.505 1848.240 2707.850 1848.675 ;
        RECT 2696.295 1847.045 2696.815 1847.585 ;
        RECT 2700.390 1846.990 2700.740 1848.240 ;
        RECT 2705.910 1846.990 2706.260 1848.240 ;
        RECT 2708.485 1847.510 2708.775 1848.675 ;
        RECT 2708.945 1848.240 2714.290 1848.675 ;
        RECT 2714.465 1848.240 2719.810 1848.675 ;
        RECT 2719.985 1848.240 2725.330 1848.675 ;
        RECT 2725.505 1848.240 2730.850 1848.675 ;
        RECT 2712.350 1846.990 2712.700 1848.240 ;
        RECT 2717.870 1846.990 2718.220 1848.240 ;
        RECT 2723.390 1846.990 2723.740 1848.240 ;
        RECT 2728.910 1846.990 2729.260 1848.240 ;
        RECT 2731.025 1847.585 2732.695 1848.675 ;
        RECT 2731.945 1847.065 2732.695 1847.585 ;
        RECT 2732.865 1847.585 2734.075 1848.675 ;
        RECT 2732.865 1847.045 2733.385 1847.585 ;
        RECT 2696.295 1844.495 2696.815 1845.035 ;
        RECT 2695.605 1843.405 2696.815 1844.495 ;
        RECT 2697.425 1843.405 2697.755 1844.165 ;
        RECT 2701.770 1843.840 2702.120 1845.090 ;
        RECT 2707.290 1843.840 2707.640 1845.090 ;
        RECT 2712.810 1843.840 2713.160 1845.090 ;
        RECT 2718.330 1843.840 2718.680 1845.090 ;
        RECT 2698.365 1843.405 2703.710 1843.840 ;
        RECT 2703.885 1843.405 2709.230 1843.840 ;
        RECT 2709.405 1843.405 2714.750 1843.840 ;
        RECT 2714.925 1843.405 2720.270 1843.840 ;
        RECT 2721.365 1843.405 2721.655 1844.570 ;
        RECT 2725.230 1843.840 2725.580 1845.090 ;
        RECT 2730.750 1843.840 2731.100 1845.090 ;
        RECT 2732.865 1844.495 2733.385 1845.035 ;
        RECT 2721.825 1843.405 2727.170 1843.840 ;
        RECT 2727.345 1843.405 2732.690 1843.840 ;
        RECT 2732.865 1843.405 2734.075 1844.495 ;
        RECT 2695.520 1843.235 2734.160 1843.405 ;
        RECT 2695.605 1842.145 2696.815 1843.235 ;
        RECT 2696.985 1842.800 2702.330 1843.235 ;
        RECT 2702.505 1842.800 2707.850 1843.235 ;
        RECT 2696.295 1841.605 2696.815 1842.145 ;
        RECT 2700.390 1841.550 2700.740 1842.800 ;
        RECT 2705.910 1841.550 2706.260 1842.800 ;
        RECT 2708.485 1842.070 2708.775 1843.235 ;
        RECT 2708.945 1842.800 2714.290 1843.235 ;
        RECT 2714.465 1842.800 2719.810 1843.235 ;
        RECT 2719.985 1842.800 2725.330 1843.235 ;
        RECT 2725.505 1842.800 2730.850 1843.235 ;
        RECT 2712.350 1841.550 2712.700 1842.800 ;
        RECT 2717.870 1841.550 2718.220 1842.800 ;
        RECT 2723.390 1841.550 2723.740 1842.800 ;
        RECT 2728.910 1841.550 2729.260 1842.800 ;
        RECT 2731.025 1842.145 2732.695 1843.235 ;
        RECT 2731.945 1841.625 2732.695 1842.145 ;
        RECT 2732.865 1842.145 2734.075 1843.235 ;
        RECT 2732.865 1841.605 2733.385 1842.145 ;
        RECT 2696.295 1839.055 2696.815 1839.595 ;
        RECT 2695.605 1837.965 2696.815 1839.055 ;
        RECT 2710.050 1838.400 2710.400 1839.650 ;
        RECT 2715.570 1838.400 2715.920 1839.650 ;
        RECT 2719.505 1839.055 2721.195 1839.575 ;
        RECT 2697.415 1837.965 2697.745 1838.345 ;
        RECT 2700.135 1837.965 2700.465 1838.345 ;
        RECT 2701.960 1837.965 2702.290 1838.345 ;
        RECT 2702.880 1837.965 2703.230 1838.345 ;
        RECT 2705.715 1837.965 2706.045 1838.345 ;
        RECT 2706.645 1837.965 2711.990 1838.400 ;
        RECT 2712.165 1837.965 2717.510 1838.400 ;
        RECT 2717.685 1837.965 2721.195 1839.055 ;
        RECT 2721.365 1837.965 2721.655 1839.130 ;
        RECT 2725.230 1838.400 2725.580 1839.650 ;
        RECT 2730.750 1838.400 2731.100 1839.650 ;
        RECT 2732.865 1839.055 2733.385 1839.595 ;
        RECT 2721.825 1837.965 2727.170 1838.400 ;
        RECT 2727.345 1837.965 2732.690 1838.400 ;
        RECT 2732.865 1837.965 2734.075 1839.055 ;
        RECT 2695.520 1837.795 2734.160 1837.965 ;
        RECT 2695.605 1836.705 2696.815 1837.795 ;
        RECT 2697.425 1837.035 2697.755 1837.795 ;
        RECT 2698.365 1837.360 2703.710 1837.795 ;
        RECT 2696.295 1836.165 2696.815 1836.705 ;
        RECT 2701.770 1836.110 2702.120 1837.360 ;
        RECT 2703.885 1836.705 2707.395 1837.795 ;
        RECT 2705.705 1836.185 2707.395 1836.705 ;
        RECT 2708.485 1836.630 2708.775 1837.795 ;
        RECT 2708.945 1837.360 2714.290 1837.795 ;
        RECT 2714.465 1837.360 2719.810 1837.795 ;
        RECT 2719.985 1837.360 2725.330 1837.795 ;
        RECT 2725.505 1837.360 2730.850 1837.795 ;
        RECT 2712.350 1836.110 2712.700 1837.360 ;
        RECT 2717.870 1836.110 2718.220 1837.360 ;
        RECT 2723.390 1836.110 2723.740 1837.360 ;
        RECT 2728.910 1836.110 2729.260 1837.360 ;
        RECT 2731.025 1836.705 2732.695 1837.795 ;
        RECT 2731.945 1836.185 2732.695 1836.705 ;
        RECT 2732.865 1836.705 2734.075 1837.795 ;
        RECT 2732.865 1836.165 2733.385 1836.705 ;
        RECT 2696.295 1833.615 2696.815 1834.155 ;
        RECT 2695.605 1832.525 2696.815 1833.615 ;
        RECT 2710.050 1832.960 2710.400 1834.210 ;
        RECT 2715.570 1832.960 2715.920 1834.210 ;
        RECT 2719.505 1833.615 2721.195 1834.135 ;
        RECT 2697.415 1832.525 2697.745 1832.905 ;
        RECT 2700.135 1832.525 2700.465 1832.905 ;
        RECT 2701.960 1832.525 2702.290 1832.905 ;
        RECT 2702.880 1832.525 2703.230 1832.905 ;
        RECT 2705.715 1832.525 2706.045 1832.905 ;
        RECT 2706.645 1832.525 2711.990 1832.960 ;
        RECT 2712.165 1832.525 2717.510 1832.960 ;
        RECT 2717.685 1832.525 2721.195 1833.615 ;
        RECT 2721.365 1832.525 2721.655 1833.690 ;
        RECT 2725.230 1832.960 2725.580 1834.210 ;
        RECT 2730.750 1832.960 2731.100 1834.210 ;
        RECT 2732.865 1833.615 2733.385 1834.155 ;
        RECT 2721.825 1832.525 2727.170 1832.960 ;
        RECT 2727.345 1832.525 2732.690 1832.960 ;
        RECT 2732.865 1832.525 2734.075 1833.615 ;
        RECT 2695.520 1832.355 2734.160 1832.525 ;
        RECT 2695.605 1831.265 2696.815 1832.355 ;
        RECT 2697.425 1831.595 2697.755 1832.355 ;
        RECT 2698.365 1831.265 2700.955 1832.355 ;
        RECT 2696.295 1830.725 2696.815 1831.265 ;
        RECT 2699.745 1830.745 2700.955 1831.265 ;
        RECT 2702.095 1831.215 2702.265 1832.355 ;
        RECT 2704.635 1831.595 2704.805 1832.355 ;
        RECT 2705.725 1831.265 2708.315 1832.355 ;
        RECT 2707.105 1830.745 2708.315 1831.265 ;
        RECT 2708.485 1831.190 2708.775 1832.355 ;
        RECT 2708.945 1831.920 2714.290 1832.355 ;
        RECT 2714.465 1831.920 2719.810 1832.355 ;
        RECT 2719.985 1831.920 2725.330 1832.355 ;
        RECT 2725.505 1831.920 2730.850 1832.355 ;
        RECT 2712.350 1830.670 2712.700 1831.920 ;
        RECT 2717.870 1830.670 2718.220 1831.920 ;
        RECT 2723.390 1830.670 2723.740 1831.920 ;
        RECT 2728.910 1830.670 2729.260 1831.920 ;
        RECT 2731.025 1831.265 2732.695 1832.355 ;
        RECT 2731.945 1830.745 2732.695 1831.265 ;
        RECT 2732.865 1831.265 2734.075 1832.355 ;
        RECT 2732.865 1830.725 2733.385 1831.265 ;
        RECT 2696.295 1828.175 2696.815 1828.715 ;
        RECT 2695.605 1827.085 2696.815 1828.175 ;
        RECT 2700.390 1827.520 2700.740 1828.770 ;
        RECT 2705.910 1827.520 2706.260 1828.770 ;
        RECT 2711.430 1827.520 2711.780 1828.770 ;
        RECT 2716.950 1827.520 2717.300 1828.770 ;
        RECT 2719.985 1828.175 2720.735 1828.695 ;
        RECT 2696.985 1827.085 2702.330 1827.520 ;
        RECT 2702.505 1827.085 2707.850 1827.520 ;
        RECT 2708.025 1827.085 2713.370 1827.520 ;
        RECT 2713.545 1827.085 2718.890 1827.520 ;
        RECT 2719.065 1827.085 2720.735 1828.175 ;
        RECT 2721.365 1827.085 2721.655 1828.250 ;
        RECT 2725.230 1827.520 2725.580 1828.770 ;
        RECT 2730.750 1827.520 2731.100 1828.770 ;
        RECT 2732.865 1828.175 2733.385 1828.715 ;
        RECT 2721.825 1827.085 2727.170 1827.520 ;
        RECT 2727.345 1827.085 2732.690 1827.520 ;
        RECT 2732.865 1827.085 2734.075 1828.175 ;
        RECT 2695.520 1826.915 2734.160 1827.085 ;
        RECT 2695.605 1825.825 2696.815 1826.915 ;
        RECT 2697.425 1826.155 2697.755 1826.915 ;
        RECT 2698.365 1826.480 2703.710 1826.915 ;
        RECT 2696.295 1825.285 2696.815 1825.825 ;
        RECT 2701.770 1825.230 2702.120 1826.480 ;
        RECT 2703.885 1825.825 2707.395 1826.915 ;
        RECT 2705.705 1825.305 2707.395 1825.825 ;
        RECT 2708.485 1825.750 2708.775 1826.915 ;
        RECT 2708.945 1826.480 2714.290 1826.915 ;
        RECT 2714.465 1826.480 2719.810 1826.915 ;
        RECT 2719.985 1826.480 2725.330 1826.915 ;
        RECT 2725.505 1826.480 2730.850 1826.915 ;
        RECT 2712.350 1825.230 2712.700 1826.480 ;
        RECT 2717.870 1825.230 2718.220 1826.480 ;
        RECT 2723.390 1825.230 2723.740 1826.480 ;
        RECT 2728.910 1825.230 2729.260 1826.480 ;
        RECT 2731.025 1825.825 2732.695 1826.915 ;
        RECT 2731.945 1825.305 2732.695 1825.825 ;
        RECT 2732.865 1825.825 2734.075 1826.915 ;
        RECT 2732.865 1825.285 2733.385 1825.825 ;
        RECT 2696.295 1822.735 2696.815 1823.275 ;
        RECT 2695.605 1821.645 2696.815 1822.735 ;
        RECT 2700.390 1822.080 2700.740 1823.330 ;
        RECT 2705.910 1822.080 2706.260 1823.330 ;
        RECT 2711.430 1822.080 2711.780 1823.330 ;
        RECT 2716.950 1822.080 2717.300 1823.330 ;
        RECT 2719.985 1822.735 2720.735 1823.255 ;
        RECT 2696.985 1821.645 2702.330 1822.080 ;
        RECT 2702.505 1821.645 2707.850 1822.080 ;
        RECT 2708.025 1821.645 2713.370 1822.080 ;
        RECT 2713.545 1821.645 2718.890 1822.080 ;
        RECT 2719.065 1821.645 2720.735 1822.735 ;
        RECT 2721.365 1821.645 2721.655 1822.810 ;
        RECT 2725.230 1822.080 2725.580 1823.330 ;
        RECT 2730.750 1822.080 2731.100 1823.330 ;
        RECT 2732.865 1822.735 2733.385 1823.275 ;
        RECT 2721.825 1821.645 2727.170 1822.080 ;
        RECT 2727.345 1821.645 2732.690 1822.080 ;
        RECT 2732.865 1821.645 2734.075 1822.735 ;
        RECT 2695.520 1821.475 2734.160 1821.645 ;
        RECT 2695.605 1820.385 2696.815 1821.475 ;
        RECT 2696.985 1820.385 2700.495 1821.475 ;
        RECT 2696.295 1819.845 2696.815 1820.385 ;
        RECT 2698.805 1819.865 2700.495 1820.385 ;
        RECT 2702.455 1820.335 2702.785 1821.475 ;
        RECT 2702.965 1821.040 2708.310 1821.475 ;
        RECT 2706.370 1819.790 2706.720 1821.040 ;
        RECT 2708.485 1820.310 2708.775 1821.475 ;
        RECT 2708.945 1821.040 2714.290 1821.475 ;
        RECT 2714.465 1821.040 2719.810 1821.475 ;
        RECT 2719.985 1821.040 2725.330 1821.475 ;
        RECT 2725.505 1821.040 2730.850 1821.475 ;
        RECT 2712.350 1819.790 2712.700 1821.040 ;
        RECT 2717.870 1819.790 2718.220 1821.040 ;
        RECT 2723.390 1819.790 2723.740 1821.040 ;
        RECT 2728.910 1819.790 2729.260 1821.040 ;
        RECT 2731.025 1820.385 2732.695 1821.475 ;
        RECT 2731.945 1819.865 2732.695 1820.385 ;
        RECT 2732.865 1820.385 2734.075 1821.475 ;
        RECT 2732.865 1819.845 2733.385 1820.385 ;
        RECT 2696.295 1817.295 2696.815 1817.835 ;
        RECT 2700.185 1817.295 2701.875 1817.815 ;
        RECT 2695.605 1816.205 2696.815 1817.295 ;
        RECT 2697.425 1816.205 2697.755 1816.965 ;
        RECT 2698.365 1816.205 2701.875 1817.295 ;
        RECT 2703.535 1816.205 2703.705 1816.645 ;
        RECT 2708.670 1816.640 2709.020 1817.890 ;
        RECT 2714.190 1816.640 2714.540 1817.890 ;
        RECT 2718.125 1817.295 2719.815 1817.815 ;
        RECT 2720.675 1817.295 2721.195 1817.835 ;
        RECT 2704.310 1816.205 2704.640 1816.565 ;
        RECT 2705.265 1816.205 2710.610 1816.640 ;
        RECT 2710.785 1816.205 2716.130 1816.640 ;
        RECT 2716.305 1816.205 2719.815 1817.295 ;
        RECT 2719.985 1816.205 2721.195 1817.295 ;
        RECT 2721.365 1816.205 2721.655 1817.370 ;
        RECT 2725.230 1816.640 2725.580 1817.890 ;
        RECT 2730.750 1816.640 2731.100 1817.890 ;
        RECT 2732.865 1817.295 2733.385 1817.835 ;
        RECT 2721.825 1816.205 2727.170 1816.640 ;
        RECT 2727.345 1816.205 2732.690 1816.640 ;
        RECT 2732.865 1816.205 2734.075 1817.295 ;
        RECT 2695.520 1816.035 2734.160 1816.205 ;
        RECT 2695.605 1814.945 2696.815 1816.035 ;
        RECT 2696.985 1815.600 2702.330 1816.035 ;
        RECT 2702.505 1815.600 2707.850 1816.035 ;
        RECT 2696.295 1814.405 2696.815 1814.945 ;
        RECT 2700.390 1814.350 2700.740 1815.600 ;
        RECT 2705.910 1814.350 2706.260 1815.600 ;
        RECT 2708.485 1814.870 2708.775 1816.035 ;
        RECT 2708.945 1815.600 2714.290 1816.035 ;
        RECT 2714.465 1815.600 2719.810 1816.035 ;
        RECT 2719.985 1815.600 2725.330 1816.035 ;
        RECT 2712.350 1814.350 2712.700 1815.600 ;
        RECT 2717.870 1814.350 2718.220 1815.600 ;
        RECT 2723.390 1814.350 2723.740 1815.600 ;
        RECT 2725.595 1815.235 2725.765 1816.035 ;
        RECT 2726.435 1815.235 2726.605 1816.035 ;
        RECT 2727.275 1815.235 2727.445 1816.035 ;
        RECT 2728.035 1815.235 2728.365 1816.035 ;
        RECT 2728.875 1815.235 2729.205 1816.035 ;
        RECT 2729.715 1815.235 2730.045 1816.035 ;
        RECT 2730.555 1815.235 2730.885 1816.035 ;
        RECT 2731.395 1815.235 2731.725 1816.035 ;
        RECT 2732.235 1814.885 2732.565 1816.035 ;
        RECT 2732.865 1814.945 2734.075 1816.035 ;
        RECT 2732.865 1814.405 2733.385 1814.945 ;
        RECT 2696.295 1811.855 2696.815 1812.395 ;
        RECT 2695.605 1810.765 2696.815 1811.855 ;
        RECT 2697.425 1810.765 2697.755 1811.525 ;
        RECT 2701.770 1811.200 2702.120 1812.450 ;
        RECT 2707.290 1811.200 2707.640 1812.450 ;
        RECT 2712.810 1811.200 2713.160 1812.450 ;
        RECT 2718.330 1811.200 2718.680 1812.450 ;
        RECT 2698.365 1810.765 2703.710 1811.200 ;
        RECT 2703.885 1810.765 2709.230 1811.200 ;
        RECT 2709.405 1810.765 2714.750 1811.200 ;
        RECT 2714.925 1810.765 2720.270 1811.200 ;
        RECT 2721.365 1810.765 2721.655 1811.930 ;
        RECT 2725.230 1811.200 2725.580 1812.450 ;
        RECT 2730.750 1811.200 2731.100 1812.450 ;
        RECT 2732.865 1811.855 2733.385 1812.395 ;
        RECT 2721.825 1810.765 2727.170 1811.200 ;
        RECT 2727.345 1810.765 2732.690 1811.200 ;
        RECT 2732.865 1810.765 2734.075 1811.855 ;
        RECT 2695.520 1810.595 2734.160 1810.765 ;
        RECT 2695.605 1809.505 2696.815 1810.595 ;
        RECT 2696.985 1810.160 2702.330 1810.595 ;
        RECT 2702.505 1810.160 2707.850 1810.595 ;
        RECT 2696.295 1808.965 2696.815 1809.505 ;
        RECT 2700.390 1808.910 2700.740 1810.160 ;
        RECT 2705.910 1808.910 2706.260 1810.160 ;
        RECT 2708.485 1809.430 2708.775 1810.595 ;
        RECT 2708.945 1810.160 2714.290 1810.595 ;
        RECT 2714.465 1810.160 2719.810 1810.595 ;
        RECT 2719.985 1810.160 2725.330 1810.595 ;
        RECT 2725.505 1810.160 2730.850 1810.595 ;
        RECT 2712.350 1808.910 2712.700 1810.160 ;
        RECT 2717.870 1808.910 2718.220 1810.160 ;
        RECT 2723.390 1808.910 2723.740 1810.160 ;
        RECT 2728.910 1808.910 2729.260 1810.160 ;
        RECT 2731.025 1809.505 2732.695 1810.595 ;
        RECT 2731.945 1808.985 2732.695 1809.505 ;
        RECT 2732.865 1809.505 2734.075 1810.595 ;
        RECT 2732.865 1808.965 2733.385 1809.505 ;
        RECT 2522.135 1807.365 2523.935 1807.535 ;
        RECT 2522.830 1806.640 2523.160 1807.365 ;
        RECT 2696.295 1806.415 2696.815 1806.955 ;
        RECT 2695.605 1805.325 2696.815 1806.415 ;
        RECT 2697.715 1805.325 2698.045 1805.835 ;
        RECT 2703.150 1805.760 2703.500 1807.010 ;
        RECT 2708.670 1805.760 2709.020 1807.010 ;
        RECT 2714.190 1805.760 2714.540 1807.010 ;
        RECT 2718.125 1806.415 2719.815 1806.935 ;
        RECT 2720.675 1806.415 2721.195 1806.955 ;
        RECT 2699.745 1805.325 2705.090 1805.760 ;
        RECT 2705.265 1805.325 2710.610 1805.760 ;
        RECT 2710.785 1805.325 2716.130 1805.760 ;
        RECT 2716.305 1805.325 2719.815 1806.415 ;
        RECT 2719.985 1805.325 2721.195 1806.415 ;
        RECT 2721.365 1805.325 2721.655 1806.490 ;
        RECT 2725.230 1805.760 2725.580 1807.010 ;
        RECT 2730.750 1805.760 2731.100 1807.010 ;
        RECT 2732.865 1806.415 2733.385 1806.955 ;
        RECT 2721.825 1805.325 2727.170 1805.760 ;
        RECT 2727.345 1805.325 2732.690 1805.760 ;
        RECT 2732.865 1805.325 2734.075 1806.415 ;
        RECT 2695.520 1805.155 2734.160 1805.325 ;
        RECT 2695.605 1804.065 2696.815 1805.155 ;
        RECT 2697.425 1804.395 2697.755 1805.155 ;
        RECT 2698.365 1804.720 2703.710 1805.155 ;
        RECT 2696.295 1803.525 2696.815 1804.065 ;
        RECT 2701.770 1803.470 2702.120 1804.720 ;
        RECT 2703.885 1804.065 2707.395 1805.155 ;
        RECT 2705.705 1803.545 2707.395 1804.065 ;
        RECT 2708.485 1803.990 2708.775 1805.155 ;
        RECT 2708.945 1804.720 2714.290 1805.155 ;
        RECT 2714.465 1804.720 2719.810 1805.155 ;
        RECT 2719.985 1804.720 2725.330 1805.155 ;
        RECT 2725.505 1804.720 2730.850 1805.155 ;
        RECT 2712.350 1803.470 2712.700 1804.720 ;
        RECT 2717.870 1803.470 2718.220 1804.720 ;
        RECT 2723.390 1803.470 2723.740 1804.720 ;
        RECT 2728.910 1803.470 2729.260 1804.720 ;
        RECT 2731.025 1804.065 2732.695 1805.155 ;
        RECT 2731.945 1803.545 2732.695 1804.065 ;
        RECT 2732.865 1804.065 2734.075 1805.155 ;
        RECT 2732.865 1803.525 2733.385 1804.065 ;
        RECT 2696.295 1800.975 2696.815 1801.515 ;
        RECT 2522.135 1799.835 2523.935 1800.005 ;
        RECT 2695.605 1799.885 2696.815 1800.975 ;
        RECT 2697.735 1799.885 2697.905 1800.645 ;
        RECT 2700.275 1799.885 2700.445 1801.025 ;
        RECT 2701.590 1799.885 2701.920 1800.600 ;
        RECT 2708.210 1800.320 2708.560 1801.570 ;
        RECT 2713.730 1800.320 2714.080 1801.570 ;
        RECT 2719.250 1800.320 2719.600 1801.570 ;
        RECT 2704.805 1799.885 2710.150 1800.320 ;
        RECT 2710.325 1799.885 2715.670 1800.320 ;
        RECT 2715.845 1799.885 2721.190 1800.320 ;
        RECT 2721.365 1799.885 2721.655 1801.050 ;
        RECT 2725.230 1800.320 2725.580 1801.570 ;
        RECT 2730.750 1800.320 2731.100 1801.570 ;
        RECT 2732.865 1800.975 2733.385 1801.515 ;
        RECT 2721.825 1799.885 2727.170 1800.320 ;
        RECT 2727.345 1799.885 2732.690 1800.320 ;
        RECT 2732.865 1799.885 2734.075 1800.975 ;
        RECT 2522.830 1799.110 2523.160 1799.835 ;
        RECT 2695.520 1799.715 2734.160 1799.885 ;
        RECT 2695.605 1798.625 2696.815 1799.715 ;
        RECT 2696.985 1799.205 2697.245 1799.715 ;
        RECT 2697.905 1799.210 2698.520 1799.715 ;
        RECT 2698.325 1799.035 2698.520 1799.210 ;
        RECT 2699.335 1799.170 2699.550 1799.715 ;
        RECT 2700.205 1799.280 2705.550 1799.715 ;
        RECT 2698.325 1798.845 2698.655 1799.035 ;
        RECT 2696.295 1798.085 2696.815 1798.625 ;
        RECT 2703.610 1798.030 2703.960 1799.280 ;
        RECT 2705.725 1798.625 2708.315 1799.715 ;
        RECT 2707.105 1798.105 2708.315 1798.625 ;
        RECT 2708.485 1798.550 2708.775 1799.715 ;
        RECT 2708.945 1799.280 2714.290 1799.715 ;
        RECT 2714.465 1799.280 2719.810 1799.715 ;
        RECT 2719.985 1799.280 2725.330 1799.715 ;
        RECT 2725.505 1799.280 2730.850 1799.715 ;
        RECT 2712.350 1798.030 2712.700 1799.280 ;
        RECT 2717.870 1798.030 2718.220 1799.280 ;
        RECT 2723.390 1798.030 2723.740 1799.280 ;
        RECT 2728.910 1798.030 2729.260 1799.280 ;
        RECT 2731.025 1798.625 2732.695 1799.715 ;
        RECT 2731.945 1798.105 2732.695 1798.625 ;
        RECT 2732.865 1798.625 2734.075 1799.715 ;
        RECT 2732.865 1798.085 2733.385 1798.625 ;
        RECT 2696.295 1795.535 2696.815 1796.075 ;
        RECT 2695.605 1794.445 2696.815 1795.535 ;
        RECT 2697.425 1794.445 2697.755 1795.205 ;
        RECT 2701.770 1794.880 2702.120 1796.130 ;
        RECT 2707.290 1794.880 2707.640 1796.130 ;
        RECT 2712.810 1794.880 2713.160 1796.130 ;
        RECT 2718.330 1794.880 2718.680 1796.130 ;
        RECT 2698.365 1794.445 2703.710 1794.880 ;
        RECT 2703.885 1794.445 2709.230 1794.880 ;
        RECT 2709.405 1794.445 2714.750 1794.880 ;
        RECT 2714.925 1794.445 2720.270 1794.880 ;
        RECT 2721.365 1794.445 2721.655 1795.610 ;
        RECT 2725.230 1794.880 2725.580 1796.130 ;
        RECT 2730.750 1794.880 2731.100 1796.130 ;
        RECT 2732.865 1795.535 2733.385 1796.075 ;
        RECT 2721.825 1794.445 2727.170 1794.880 ;
        RECT 2727.345 1794.445 2732.690 1794.880 ;
        RECT 2732.865 1794.445 2734.075 1795.535 ;
        RECT 2695.520 1794.275 2734.160 1794.445 ;
        RECT 2522.135 1793.855 2523.935 1794.025 ;
        RECT 2522.830 1793.130 2523.160 1793.855 ;
        RECT 2695.605 1793.185 2696.815 1794.275 ;
        RECT 2696.985 1793.185 2698.195 1794.275 ;
        RECT 2698.865 1793.815 2699.115 1794.275 ;
        RECT 2699.795 1793.815 2700.045 1794.275 ;
        RECT 2701.115 1793.815 2701.365 1794.275 ;
        RECT 2702.045 1793.840 2707.390 1794.275 ;
        RECT 2696.295 1792.645 2696.815 1793.185 ;
        RECT 2697.675 1792.645 2698.195 1793.185 ;
        RECT 2705.450 1792.590 2705.800 1793.840 ;
        RECT 2708.485 1793.110 2708.775 1794.275 ;
        RECT 2708.945 1793.840 2714.290 1794.275 ;
        RECT 2714.465 1793.840 2719.810 1794.275 ;
        RECT 2719.985 1793.840 2725.330 1794.275 ;
        RECT 2725.505 1793.840 2730.850 1794.275 ;
        RECT 2712.350 1792.590 2712.700 1793.840 ;
        RECT 2717.870 1792.590 2718.220 1793.840 ;
        RECT 2723.390 1792.590 2723.740 1793.840 ;
        RECT 2728.910 1792.590 2729.260 1793.840 ;
        RECT 2731.025 1793.185 2732.695 1794.275 ;
        RECT 2731.945 1792.665 2732.695 1793.185 ;
        RECT 2732.865 1793.185 2734.075 1794.275 ;
        RECT 2732.865 1792.645 2733.385 1793.185 ;
        RECT 2369.980 1790.050 2370.155 1790.600 ;
        RECT 2696.295 1790.095 2696.815 1790.635 ;
        RECT 2369.980 1788.450 2370.150 1790.050 ;
        RECT 2695.605 1789.005 2696.815 1790.095 ;
        RECT 2697.905 1789.005 2698.165 1790.145 ;
        RECT 2700.190 1789.005 2700.470 1789.805 ;
        RECT 2701.885 1789.005 2702.170 1789.805 ;
        RECT 2702.840 1789.005 2703.090 1790.145 ;
        RECT 2707.290 1789.440 2707.640 1790.690 ;
        RECT 2712.810 1789.440 2713.160 1790.690 ;
        RECT 2718.330 1789.440 2718.680 1790.690 ;
        RECT 2703.885 1789.005 2709.230 1789.440 ;
        RECT 2709.405 1789.005 2714.750 1789.440 ;
        RECT 2714.925 1789.005 2720.270 1789.440 ;
        RECT 2721.365 1789.005 2721.655 1790.170 ;
        RECT 2725.230 1789.440 2725.580 1790.690 ;
        RECT 2730.750 1789.440 2731.100 1790.690 ;
        RECT 2732.865 1790.095 2733.385 1790.635 ;
        RECT 2721.825 1789.005 2727.170 1789.440 ;
        RECT 2727.345 1789.005 2732.690 1789.440 ;
        RECT 2732.865 1789.005 2734.075 1790.095 ;
        RECT 2695.520 1788.835 2734.160 1789.005 ;
        RECT 2368.165 1787.040 2368.335 1787.770 ;
        RECT 2369.980 1787.310 2370.155 1788.450 ;
        RECT 2522.135 1787.910 2523.935 1788.080 ;
        RECT 2369.980 1787.040 2370.150 1787.310 ;
        RECT 2375.680 1787.040 2375.850 1787.770 ;
        RECT 2381.295 1787.040 2381.465 1787.770 ;
        RECT 2384.040 1787.040 2384.210 1787.770 ;
        RECT 2385.030 1787.040 2385.200 1787.770 ;
        RECT 2390.940 1787.040 2391.110 1787.770 ;
        RECT 2396.555 1787.040 2396.725 1787.770 ;
        RECT 2399.300 1787.040 2399.470 1787.770 ;
        RECT 2400.290 1787.040 2400.460 1787.770 ;
        RECT 2406.200 1787.040 2406.370 1787.770 ;
        RECT 2411.815 1787.040 2411.985 1787.770 ;
        RECT 2414.560 1787.040 2414.730 1787.770 ;
        RECT 2415.550 1787.040 2415.720 1787.770 ;
        RECT 2421.460 1787.040 2421.630 1787.770 ;
        RECT 2427.075 1787.040 2427.245 1787.770 ;
        RECT 2429.820 1787.040 2429.990 1787.770 ;
        RECT 2430.810 1787.040 2430.980 1787.770 ;
        RECT 2436.720 1787.040 2436.890 1787.770 ;
        RECT 2442.335 1787.040 2442.505 1787.770 ;
        RECT 2445.080 1787.040 2445.250 1787.770 ;
        RECT 2446.070 1787.040 2446.240 1787.770 ;
        RECT 2522.830 1787.185 2523.160 1787.910 ;
        RECT 2695.605 1787.745 2696.815 1788.835 ;
        RECT 2697.425 1788.075 2697.755 1788.835 ;
        RECT 2696.295 1787.205 2696.815 1787.745 ;
        RECT 2698.825 1787.695 2699.085 1788.835 ;
        RECT 2699.755 1787.695 2700.035 1788.835 ;
        RECT 2700.205 1788.400 2705.550 1788.835 ;
        RECT 2703.610 1787.150 2703.960 1788.400 ;
        RECT 2705.725 1787.745 2708.315 1788.835 ;
        RECT 2707.105 1787.225 2708.315 1787.745 ;
        RECT 2708.485 1787.670 2708.775 1788.835 ;
        RECT 2708.945 1788.400 2714.290 1788.835 ;
        RECT 2714.465 1788.400 2719.810 1788.835 ;
        RECT 2719.985 1788.400 2725.330 1788.835 ;
        RECT 2725.505 1788.400 2730.850 1788.835 ;
        RECT 2712.350 1787.150 2712.700 1788.400 ;
        RECT 2717.870 1787.150 2718.220 1788.400 ;
        RECT 2723.390 1787.150 2723.740 1788.400 ;
        RECT 2728.910 1787.150 2729.260 1788.400 ;
        RECT 2731.025 1787.745 2732.695 1788.835 ;
        RECT 2731.945 1787.225 2732.695 1787.745 ;
        RECT 2732.865 1787.745 2734.075 1788.835 ;
        RECT 2732.865 1787.205 2733.385 1787.745 ;
        RECT 2367.995 1787.035 2370.745 1787.040 ;
        RECT 2375.510 1787.035 2378.260 1787.040 ;
        RECT 2381.125 1787.035 2385.850 1787.040 ;
        RECT 2390.770 1787.035 2393.520 1787.040 ;
        RECT 2396.385 1787.035 2401.110 1787.040 ;
        RECT 2406.030 1787.035 2408.780 1787.040 ;
        RECT 2411.645 1787.035 2416.370 1787.040 ;
        RECT 2421.290 1787.035 2424.040 1787.040 ;
        RECT 2426.905 1787.035 2431.630 1787.040 ;
        RECT 2436.550 1787.035 2439.300 1787.040 ;
        RECT 2442.165 1787.035 2446.890 1787.040 ;
        RECT 2343.000 1785.435 2447.045 1787.035 ;
        RECT 2371.495 1785.430 2386.005 1785.435 ;
        RECT 2386.755 1785.430 2401.265 1785.435 ;
        RECT 2402.015 1785.430 2416.525 1785.435 ;
        RECT 2417.275 1785.430 2431.785 1785.435 ;
        RECT 2432.535 1785.430 2447.045 1785.435 ;
        RECT 2371.495 1785.425 2380.235 1785.430 ;
        RECT 2381.125 1785.425 2385.845 1785.430 ;
        RECT 2386.755 1785.425 2395.495 1785.430 ;
        RECT 2396.385 1785.425 2401.105 1785.430 ;
        RECT 2402.015 1785.425 2410.755 1785.430 ;
        RECT 2411.645 1785.425 2416.365 1785.430 ;
        RECT 2417.275 1785.425 2426.015 1785.430 ;
        RECT 2426.905 1785.425 2431.625 1785.430 ;
        RECT 2432.535 1785.425 2441.275 1785.430 ;
        RECT 2442.165 1785.425 2446.885 1785.430 ;
        RECT 2372.285 1784.925 2372.455 1785.425 ;
        RECT 2374.205 1784.925 2374.375 1785.425 ;
        RECT 2375.665 1784.925 2375.835 1785.425 ;
        RECT 2376.605 1784.925 2376.775 1785.425 ;
        RECT 2378.525 1784.925 2378.695 1785.425 ;
        RECT 2381.295 1784.695 2381.465 1785.425 ;
        RECT 2384.040 1784.695 2384.210 1785.425 ;
        RECT 2385.025 1784.695 2385.195 1785.425 ;
        RECT 2387.545 1784.925 2387.715 1785.425 ;
        RECT 2389.465 1784.925 2389.635 1785.425 ;
        RECT 2390.925 1784.925 2391.095 1785.425 ;
        RECT 2391.865 1784.925 2392.035 1785.425 ;
        RECT 2393.785 1784.925 2393.955 1785.425 ;
        RECT 2396.555 1784.695 2396.725 1785.425 ;
        RECT 2399.300 1784.695 2399.470 1785.425 ;
        RECT 2400.285 1784.695 2400.455 1785.425 ;
        RECT 2402.805 1784.925 2402.975 1785.425 ;
        RECT 2404.725 1784.925 2404.895 1785.425 ;
        RECT 2406.185 1784.925 2406.355 1785.425 ;
        RECT 2407.125 1784.925 2407.295 1785.425 ;
        RECT 2409.045 1784.925 2409.215 1785.425 ;
        RECT 2411.815 1784.695 2411.985 1785.425 ;
        RECT 2414.560 1784.695 2414.730 1785.425 ;
        RECT 2415.545 1784.695 2415.715 1785.425 ;
        RECT 2418.065 1784.925 2418.235 1785.425 ;
        RECT 2419.985 1784.925 2420.155 1785.425 ;
        RECT 2421.445 1784.925 2421.615 1785.425 ;
        RECT 2422.385 1784.925 2422.555 1785.425 ;
        RECT 2424.305 1784.925 2424.475 1785.425 ;
        RECT 2427.075 1784.695 2427.245 1785.425 ;
        RECT 2429.820 1784.695 2429.990 1785.425 ;
        RECT 2430.805 1784.695 2430.975 1785.425 ;
        RECT 2433.325 1784.925 2433.495 1785.425 ;
        RECT 2435.245 1784.925 2435.415 1785.425 ;
        RECT 2436.705 1784.925 2436.875 1785.425 ;
        RECT 2437.645 1784.925 2437.815 1785.425 ;
        RECT 2439.565 1784.925 2439.735 1785.425 ;
        RECT 2442.335 1784.695 2442.505 1785.425 ;
        RECT 2445.080 1784.695 2445.250 1785.425 ;
        RECT 2446.065 1784.695 2446.235 1785.425 ;
        RECT 2696.295 1784.655 2696.815 1785.195 ;
        RECT 2695.605 1783.565 2696.815 1784.655 ;
        RECT 2697.735 1783.565 2697.905 1784.325 ;
        RECT 2700.275 1783.565 2700.445 1784.705 ;
        RECT 2704.530 1784.000 2704.880 1785.250 ;
        RECT 2710.050 1784.000 2710.400 1785.250 ;
        RECT 2715.570 1784.000 2715.920 1785.250 ;
        RECT 2719.505 1784.655 2721.195 1785.175 ;
        RECT 2701.125 1783.565 2706.470 1784.000 ;
        RECT 2706.645 1783.565 2711.990 1784.000 ;
        RECT 2712.165 1783.565 2717.510 1784.000 ;
        RECT 2717.685 1783.565 2721.195 1784.655 ;
        RECT 2721.365 1783.565 2721.655 1784.730 ;
        RECT 2725.230 1784.000 2725.580 1785.250 ;
        RECT 2730.750 1784.000 2731.100 1785.250 ;
        RECT 2732.865 1784.655 2733.385 1785.195 ;
        RECT 2721.825 1783.565 2727.170 1784.000 ;
        RECT 2727.345 1783.565 2732.690 1784.000 ;
        RECT 2732.865 1783.565 2734.075 1784.655 ;
        RECT 2695.520 1783.395 2734.160 1783.565 ;
        RECT 2522.135 1782.265 2523.935 1782.435 ;
        RECT 2695.605 1782.305 2696.815 1783.395 ;
        RECT 2697.425 1782.635 2697.755 1783.395 ;
        RECT 2698.365 1782.960 2703.710 1783.395 ;
        RECT 2522.830 1781.540 2523.160 1782.265 ;
        RECT 2696.295 1781.765 2696.815 1782.305 ;
        RECT 2701.770 1781.710 2702.120 1782.960 ;
        RECT 2703.885 1782.305 2707.395 1783.395 ;
        RECT 2705.705 1781.785 2707.395 1782.305 ;
        RECT 2708.485 1782.230 2708.775 1783.395 ;
        RECT 2708.945 1782.960 2714.290 1783.395 ;
        RECT 2714.465 1782.960 2719.810 1783.395 ;
        RECT 2719.985 1782.960 2725.330 1783.395 ;
        RECT 2725.505 1782.960 2730.850 1783.395 ;
        RECT 2712.350 1781.710 2712.700 1782.960 ;
        RECT 2717.870 1781.710 2718.220 1782.960 ;
        RECT 2723.390 1781.710 2723.740 1782.960 ;
        RECT 2728.910 1781.710 2729.260 1782.960 ;
        RECT 2731.025 1782.305 2732.695 1783.395 ;
        RECT 2731.945 1781.785 2732.695 1782.305 ;
        RECT 2732.865 1782.305 2734.075 1783.395 ;
        RECT 2732.865 1781.765 2733.385 1782.305 ;
        RECT 2696.295 1779.215 2696.815 1779.755 ;
        RECT 2695.605 1778.125 2696.815 1779.215 ;
        RECT 2700.390 1778.560 2700.740 1779.810 ;
        RECT 2705.910 1778.560 2706.260 1779.810 ;
        RECT 2711.430 1778.560 2711.780 1779.810 ;
        RECT 2716.950 1778.560 2717.300 1779.810 ;
        RECT 2719.985 1779.215 2720.735 1779.735 ;
        RECT 2696.985 1778.125 2702.330 1778.560 ;
        RECT 2702.505 1778.125 2707.850 1778.560 ;
        RECT 2708.025 1778.125 2713.370 1778.560 ;
        RECT 2713.545 1778.125 2718.890 1778.560 ;
        RECT 2719.065 1778.125 2720.735 1779.215 ;
        RECT 2721.365 1778.125 2721.655 1779.290 ;
        RECT 2725.230 1778.560 2725.580 1779.810 ;
        RECT 2730.750 1778.560 2731.100 1779.810 ;
        RECT 2732.865 1779.215 2733.385 1779.755 ;
        RECT 2721.825 1778.125 2727.170 1778.560 ;
        RECT 2727.345 1778.125 2732.690 1778.560 ;
        RECT 2732.865 1778.125 2734.075 1779.215 ;
        RECT 2695.520 1777.955 2734.160 1778.125 ;
        RECT 2695.605 1776.865 2696.815 1777.955 ;
        RECT 2697.425 1777.195 2697.755 1777.955 ;
        RECT 2698.365 1777.520 2703.710 1777.955 ;
        RECT 2696.295 1776.325 2696.815 1776.865 ;
        RECT 2701.770 1776.270 2702.120 1777.520 ;
        RECT 2703.885 1776.865 2707.395 1777.955 ;
        RECT 2705.705 1776.345 2707.395 1776.865 ;
        RECT 2708.485 1776.790 2708.775 1777.955 ;
        RECT 2708.945 1777.520 2714.290 1777.955 ;
        RECT 2714.465 1777.520 2719.810 1777.955 ;
        RECT 2719.985 1777.520 2725.330 1777.955 ;
        RECT 2725.505 1777.520 2730.850 1777.955 ;
        RECT 2712.350 1776.270 2712.700 1777.520 ;
        RECT 2717.870 1776.270 2718.220 1777.520 ;
        RECT 2723.390 1776.270 2723.740 1777.520 ;
        RECT 2728.910 1776.270 2729.260 1777.520 ;
        RECT 2731.025 1776.865 2732.695 1777.955 ;
        RECT 2731.945 1776.345 2732.695 1776.865 ;
        RECT 2732.865 1776.865 2734.075 1777.955 ;
        RECT 2732.865 1776.325 2733.385 1776.865 ;
        RECT 2696.295 1773.775 2696.815 1774.315 ;
        RECT 2695.605 1772.685 2696.815 1773.775 ;
        RECT 2700.390 1773.120 2700.740 1774.370 ;
        RECT 2705.910 1773.120 2706.260 1774.370 ;
        RECT 2711.430 1773.120 2711.780 1774.370 ;
        RECT 2716.950 1773.120 2717.300 1774.370 ;
        RECT 2719.985 1773.775 2720.735 1774.295 ;
        RECT 2696.985 1772.685 2702.330 1773.120 ;
        RECT 2702.505 1772.685 2707.850 1773.120 ;
        RECT 2708.025 1772.685 2713.370 1773.120 ;
        RECT 2713.545 1772.685 2718.890 1773.120 ;
        RECT 2719.065 1772.685 2720.735 1773.775 ;
        RECT 2721.365 1772.685 2721.655 1773.850 ;
        RECT 2725.230 1773.120 2725.580 1774.370 ;
        RECT 2730.750 1773.120 2731.100 1774.370 ;
        RECT 2732.865 1773.775 2733.385 1774.315 ;
        RECT 2721.825 1772.685 2727.170 1773.120 ;
        RECT 2727.345 1772.685 2732.690 1773.120 ;
        RECT 2732.865 1772.685 2734.075 1773.775 ;
        RECT 2695.520 1772.515 2734.160 1772.685 ;
        RECT 2695.605 1771.425 2696.815 1772.515 ;
        RECT 2697.425 1771.755 2697.755 1772.515 ;
        RECT 2698.805 1771.755 2699.135 1772.515 ;
        RECT 2699.745 1772.080 2705.090 1772.515 ;
        RECT 2522.135 1770.795 2523.935 1770.965 ;
        RECT 2696.295 1770.885 2696.815 1771.425 ;
        RECT 2703.150 1770.830 2703.500 1772.080 ;
        RECT 2705.265 1771.425 2707.855 1772.515 ;
        RECT 2706.645 1770.905 2707.855 1771.425 ;
        RECT 2708.485 1771.350 2708.775 1772.515 ;
        RECT 2708.945 1772.080 2714.290 1772.515 ;
        RECT 2714.465 1772.080 2719.810 1772.515 ;
        RECT 2712.350 1770.830 2712.700 1772.080 ;
        RECT 2717.870 1770.830 2718.220 1772.080 ;
        RECT 2719.985 1771.425 2721.195 1772.515 ;
        RECT 2720.675 1770.885 2721.195 1771.425 ;
        RECT 2721.365 1771.350 2721.655 1772.515 ;
        RECT 2721.825 1772.080 2727.170 1772.515 ;
        RECT 2727.345 1772.080 2732.690 1772.515 ;
        RECT 2725.230 1770.830 2725.580 1772.080 ;
        RECT 2730.750 1770.830 2731.100 1772.080 ;
        RECT 2732.865 1771.425 2734.075 1772.515 ;
        RECT 2732.865 1770.885 2733.385 1771.425 ;
        RECT 2522.830 1770.070 2523.160 1770.795 ;
        RECT 2360.400 1710.035 2360.575 1710.585 ;
        RECT 2360.400 1708.435 2360.570 1710.035 ;
        RECT 2358.585 1707.025 2358.755 1707.755 ;
        RECT 2360.400 1707.295 2360.575 1708.435 ;
        RECT 2360.400 1707.025 2360.570 1707.295 ;
        RECT 2361.815 1707.025 2361.985 1707.755 ;
        RECT 2373.040 1707.040 2373.210 1707.760 ;
        RECT 2375.785 1707.040 2375.955 1707.760 ;
        RECT 2376.775 1707.040 2376.945 1707.760 ;
        RECT 2371.810 1707.030 2377.750 1707.040 ;
        RECT 2378.400 1707.030 2378.570 1707.755 ;
        RECT 2389.625 1707.040 2389.795 1707.760 ;
        RECT 2392.370 1707.040 2392.540 1707.760 ;
        RECT 2393.360 1707.040 2393.530 1707.760 ;
        RECT 2388.395 1707.030 2394.335 1707.040 ;
        RECT 2394.985 1707.030 2395.155 1707.760 ;
        RECT 2406.210 1707.045 2406.380 1707.765 ;
        RECT 2408.955 1707.045 2409.125 1707.765 ;
        RECT 2409.945 1707.045 2410.115 1707.765 ;
        RECT 2404.980 1707.035 2410.920 1707.045 ;
        RECT 2411.570 1707.035 2411.740 1707.765 ;
        RECT 2422.795 1707.050 2422.965 1707.770 ;
        RECT 2425.540 1707.050 2425.710 1707.770 ;
        RECT 2426.530 1707.050 2426.700 1707.770 ;
        RECT 2421.565 1707.035 2427.505 1707.050 ;
        RECT 2428.150 1707.035 2428.320 1707.765 ;
        RECT 2439.375 1707.050 2439.545 1707.770 ;
        RECT 2442.120 1707.050 2442.290 1707.770 ;
        RECT 2443.110 1707.050 2443.280 1707.770 ;
        RECT 2404.980 1707.030 2414.495 1707.035 ;
        RECT 2421.565 1707.030 2431.075 1707.035 ;
        RECT 2343.000 1705.805 2364.965 1707.025 ;
        RECT 2366.070 1705.805 2366.400 1706.525 ;
        RECT 2367.085 1705.805 2367.365 1706.265 ;
        RECT 2368.230 1705.805 2368.500 1706.585 ;
        RECT 2369.050 1705.805 2369.420 1706.185 ;
        RECT 2371.810 1705.965 2381.575 1707.030 ;
        RECT 2371.680 1705.805 2381.575 1705.965 ;
        RECT 2382.655 1705.805 2382.985 1706.525 ;
        RECT 2383.670 1705.805 2383.950 1706.265 ;
        RECT 2384.815 1705.805 2385.085 1706.585 ;
        RECT 2385.635 1705.805 2386.005 1706.185 ;
        RECT 2388.395 1705.965 2398.160 1707.030 ;
        RECT 2388.265 1705.810 2398.160 1705.965 ;
        RECT 2399.240 1705.810 2399.570 1706.530 ;
        RECT 2400.255 1705.810 2400.535 1706.270 ;
        RECT 2401.400 1705.810 2401.670 1706.590 ;
        RECT 2402.220 1705.810 2402.590 1706.190 ;
        RECT 2404.980 1705.970 2414.745 1707.030 ;
        RECT 2404.850 1705.815 2414.745 1705.970 ;
        RECT 2415.825 1705.815 2416.155 1706.535 ;
        RECT 2416.840 1705.815 2417.120 1706.275 ;
        RECT 2417.985 1705.815 2418.255 1706.595 ;
        RECT 2418.805 1705.815 2419.175 1706.195 ;
        RECT 2421.565 1705.975 2431.330 1707.030 ;
        RECT 2421.435 1705.815 2431.330 1705.975 ;
        RECT 2432.405 1705.815 2432.735 1706.535 ;
        RECT 2433.420 1705.815 2433.700 1706.275 ;
        RECT 2434.565 1705.815 2434.835 1706.595 ;
        RECT 2435.385 1705.815 2435.755 1706.195 ;
        RECT 2438.145 1705.975 2444.085 1707.050 ;
        RECT 2438.015 1705.815 2444.085 1705.975 ;
        RECT 2404.850 1705.810 2444.085 1705.815 ;
        RECT 2388.265 1705.805 2444.085 1705.810 ;
        RECT 2343.000 1705.645 2444.085 1705.805 ;
        RECT 2343.000 1705.640 2414.745 1705.645 ;
        RECT 2343.000 1705.635 2398.160 1705.640 ;
        RECT 2343.000 1705.425 2364.965 1705.635 ;
        RECT 2364.655 1705.125 2364.915 1705.425 ;
        RECT 2365.880 1705.135 2366.500 1705.635 ;
        RECT 2366.300 1704.955 2366.500 1705.135 ;
        RECT 2367.310 1705.095 2367.530 1705.635 ;
        RECT 2368.180 1704.985 2368.790 1705.635 ;
        RECT 2369.610 1705.095 2369.870 1705.635 ;
        RECT 2371.350 1705.430 2381.575 1705.635 ;
        RECT 2368.610 1704.955 2368.800 1704.985 ;
        RECT 2366.300 1704.765 2366.630 1704.955 ;
        RECT 2368.610 1704.715 2368.940 1704.955 ;
        RECT 2371.350 1704.495 2371.680 1705.430 ;
        RECT 2373.040 1704.700 2373.210 1705.430 ;
        RECT 2375.785 1704.700 2375.955 1705.430 ;
        RECT 2376.775 1704.700 2376.945 1705.430 ;
        RECT 2377.750 1705.425 2381.500 1705.430 ;
        RECT 2381.240 1705.125 2381.500 1705.425 ;
        RECT 2382.465 1705.135 2383.085 1705.635 ;
        RECT 2382.885 1704.955 2383.085 1705.135 ;
        RECT 2383.895 1705.095 2384.115 1705.635 ;
        RECT 2384.765 1704.985 2385.375 1705.635 ;
        RECT 2386.195 1705.095 2386.455 1705.635 ;
        RECT 2387.935 1705.430 2398.160 1705.635 ;
        RECT 2385.195 1704.955 2385.385 1704.985 ;
        RECT 2382.885 1704.765 2383.215 1704.955 ;
        RECT 2385.195 1704.715 2385.525 1704.955 ;
        RECT 2387.935 1704.495 2388.265 1705.430 ;
        RECT 2389.625 1704.700 2389.795 1705.430 ;
        RECT 2392.370 1704.700 2392.540 1705.430 ;
        RECT 2393.360 1704.700 2393.530 1705.430 ;
        RECT 2397.825 1705.130 2398.085 1705.430 ;
        RECT 2399.050 1705.140 2399.670 1705.640 ;
        RECT 2399.470 1704.960 2399.670 1705.140 ;
        RECT 2400.480 1705.100 2400.700 1705.640 ;
        RECT 2401.350 1704.990 2401.960 1705.640 ;
        RECT 2402.780 1705.100 2403.040 1705.640 ;
        RECT 2404.520 1705.430 2414.745 1705.640 ;
        RECT 2401.780 1704.960 2401.970 1704.990 ;
        RECT 2399.470 1704.770 2399.800 1704.960 ;
        RECT 2401.780 1704.720 2402.110 1704.960 ;
        RECT 2404.520 1704.500 2404.850 1705.430 ;
        RECT 2406.210 1704.705 2406.380 1705.430 ;
        RECT 2408.955 1704.705 2409.125 1705.430 ;
        RECT 2409.945 1704.705 2410.115 1705.430 ;
        RECT 2414.410 1705.135 2414.670 1705.430 ;
        RECT 2415.635 1705.145 2416.255 1705.645 ;
        RECT 2416.055 1704.965 2416.255 1705.145 ;
        RECT 2417.065 1705.105 2417.285 1705.645 ;
        RECT 2417.935 1704.995 2418.545 1705.645 ;
        RECT 2419.365 1705.105 2419.625 1705.645 ;
        RECT 2421.105 1705.430 2431.330 1705.645 ;
        RECT 2418.365 1704.965 2418.555 1704.995 ;
        RECT 2416.055 1704.775 2416.385 1704.965 ;
        RECT 2418.365 1704.725 2418.695 1704.965 ;
        RECT 2421.105 1704.505 2421.435 1705.430 ;
        RECT 2422.795 1704.710 2422.965 1705.430 ;
        RECT 2425.540 1704.710 2425.710 1705.430 ;
        RECT 2426.530 1704.710 2426.700 1705.430 ;
        RECT 2430.990 1705.135 2431.250 1705.430 ;
        RECT 2432.215 1705.145 2432.835 1705.645 ;
        RECT 2432.635 1704.965 2432.835 1705.145 ;
        RECT 2433.645 1705.105 2433.865 1705.645 ;
        RECT 2434.515 1704.995 2435.125 1705.645 ;
        RECT 2435.945 1705.105 2436.205 1705.645 ;
        RECT 2437.685 1705.430 2444.085 1705.645 ;
        RECT 2434.945 1704.965 2435.135 1704.995 ;
        RECT 2432.635 1704.775 2432.965 1704.965 ;
        RECT 2434.945 1704.725 2435.275 1704.965 ;
        RECT 2437.685 1704.505 2438.015 1705.430 ;
        RECT 2439.375 1704.710 2439.545 1705.430 ;
        RECT 2442.120 1704.710 2442.290 1705.430 ;
        RECT 2443.110 1704.710 2443.280 1705.430 ;
        RECT 2696.295 1675.375 2696.815 1675.915 ;
        RECT 2695.605 1674.285 2696.815 1675.375 ;
        RECT 2697.425 1674.285 2697.755 1675.065 ;
        RECT 2698.315 1674.285 2698.650 1674.710 ;
        RECT 2699.265 1674.285 2699.595 1675.045 ;
        RECT 2700.645 1674.285 2700.975 1675.045 ;
        RECT 2704.990 1674.720 2705.340 1675.970 ;
        RECT 2707.795 1675.375 2708.315 1675.915 ;
        RECT 2701.585 1674.285 2706.930 1674.720 ;
        RECT 2707.105 1674.285 2708.315 1675.375 ;
        RECT 2708.485 1674.285 2708.775 1675.450 ;
        RECT 2709.420 1674.285 2709.750 1675.045 ;
        RECT 2710.350 1674.285 2710.610 1675.435 ;
        RECT 2714.190 1674.720 2714.540 1675.970 ;
        RECT 2718.125 1675.375 2719.815 1675.895 ;
        RECT 2720.675 1675.375 2721.195 1675.915 ;
        RECT 2710.785 1674.285 2716.130 1674.720 ;
        RECT 2716.305 1674.285 2719.815 1675.375 ;
        RECT 2719.985 1674.285 2721.195 1675.375 ;
        RECT 2721.365 1674.285 2721.655 1675.450 ;
        RECT 2721.830 1674.285 2722.165 1674.710 ;
        RECT 2722.725 1674.285 2723.055 1675.065 ;
        RECT 2727.070 1674.720 2727.420 1675.970 ;
        RECT 2730.105 1675.375 2730.855 1675.895 ;
        RECT 2723.665 1674.285 2729.010 1674.720 ;
        RECT 2729.185 1674.285 2730.855 1675.375 ;
        RECT 2732.865 1675.375 2733.385 1675.915 ;
        RECT 2731.925 1674.285 2732.255 1675.045 ;
        RECT 2732.865 1674.285 2734.075 1675.375 ;
        RECT 2695.520 1674.115 2734.160 1674.285 ;
        RECT 2695.605 1673.025 2696.815 1674.115 ;
        RECT 2697.425 1673.355 2697.755 1674.115 ;
        RECT 2698.365 1673.680 2703.710 1674.115 ;
        RECT 2696.295 1672.485 2696.815 1673.025 ;
        RECT 2701.770 1672.430 2702.120 1673.680 ;
        RECT 2703.885 1673.025 2707.395 1674.115 ;
        RECT 2705.705 1672.505 2707.395 1673.025 ;
        RECT 2708.485 1672.950 2708.775 1674.115 ;
        RECT 2708.945 1673.680 2714.290 1674.115 ;
        RECT 2714.465 1673.680 2719.810 1674.115 ;
        RECT 2719.985 1673.680 2725.330 1674.115 ;
        RECT 2725.505 1673.680 2730.850 1674.115 ;
        RECT 2712.350 1672.430 2712.700 1673.680 ;
        RECT 2717.870 1672.430 2718.220 1673.680 ;
        RECT 2723.390 1672.430 2723.740 1673.680 ;
        RECT 2728.910 1672.430 2729.260 1673.680 ;
        RECT 2731.025 1673.025 2732.695 1674.115 ;
        RECT 2731.945 1672.505 2732.695 1673.025 ;
        RECT 2732.865 1673.025 2734.075 1674.115 ;
        RECT 2732.865 1672.485 2733.385 1673.025 ;
        RECT 2696.295 1669.935 2696.815 1670.475 ;
        RECT 2695.605 1668.845 2696.815 1669.935 ;
        RECT 2700.390 1669.280 2700.740 1670.530 ;
        RECT 2705.910 1669.280 2706.260 1670.530 ;
        RECT 2711.430 1669.280 2711.780 1670.530 ;
        RECT 2716.950 1669.280 2717.300 1670.530 ;
        RECT 2719.985 1669.935 2720.735 1670.455 ;
        RECT 2696.985 1668.845 2702.330 1669.280 ;
        RECT 2702.505 1668.845 2707.850 1669.280 ;
        RECT 2708.025 1668.845 2713.370 1669.280 ;
        RECT 2713.545 1668.845 2718.890 1669.280 ;
        RECT 2719.065 1668.845 2720.735 1669.935 ;
        RECT 2721.365 1668.845 2721.655 1670.010 ;
        RECT 2725.230 1669.280 2725.580 1670.530 ;
        RECT 2730.750 1669.280 2731.100 1670.530 ;
        RECT 2732.865 1669.935 2733.385 1670.475 ;
        RECT 2721.825 1668.845 2727.170 1669.280 ;
        RECT 2727.345 1668.845 2732.690 1669.280 ;
        RECT 2732.865 1668.845 2734.075 1669.935 ;
        RECT 2695.520 1668.675 2734.160 1668.845 ;
        RECT 2695.605 1667.585 2696.815 1668.675 ;
        RECT 2696.985 1668.240 2702.330 1668.675 ;
        RECT 2702.505 1668.240 2707.850 1668.675 ;
        RECT 2696.295 1667.045 2696.815 1667.585 ;
        RECT 2700.390 1666.990 2700.740 1668.240 ;
        RECT 2705.910 1666.990 2706.260 1668.240 ;
        RECT 2708.485 1667.510 2708.775 1668.675 ;
        RECT 2708.945 1668.240 2714.290 1668.675 ;
        RECT 2714.465 1668.240 2719.810 1668.675 ;
        RECT 2719.985 1668.240 2725.330 1668.675 ;
        RECT 2725.505 1668.240 2730.850 1668.675 ;
        RECT 2712.350 1666.990 2712.700 1668.240 ;
        RECT 2717.870 1666.990 2718.220 1668.240 ;
        RECT 2723.390 1666.990 2723.740 1668.240 ;
        RECT 2728.910 1666.990 2729.260 1668.240 ;
        RECT 2731.025 1667.585 2732.695 1668.675 ;
        RECT 2731.945 1667.065 2732.695 1667.585 ;
        RECT 2732.865 1667.585 2734.075 1668.675 ;
        RECT 2732.865 1667.045 2733.385 1667.585 ;
        RECT 2696.295 1664.495 2696.815 1665.035 ;
        RECT 2695.605 1663.405 2696.815 1664.495 ;
        RECT 2697.425 1663.405 2697.755 1664.165 ;
        RECT 2701.770 1663.840 2702.120 1665.090 ;
        RECT 2707.290 1663.840 2707.640 1665.090 ;
        RECT 2712.810 1663.840 2713.160 1665.090 ;
        RECT 2718.330 1663.840 2718.680 1665.090 ;
        RECT 2698.365 1663.405 2703.710 1663.840 ;
        RECT 2703.885 1663.405 2709.230 1663.840 ;
        RECT 2709.405 1663.405 2714.750 1663.840 ;
        RECT 2714.925 1663.405 2720.270 1663.840 ;
        RECT 2721.365 1663.405 2721.655 1664.570 ;
        RECT 2725.230 1663.840 2725.580 1665.090 ;
        RECT 2730.750 1663.840 2731.100 1665.090 ;
        RECT 2732.865 1664.495 2733.385 1665.035 ;
        RECT 2721.825 1663.405 2727.170 1663.840 ;
        RECT 2727.345 1663.405 2732.690 1663.840 ;
        RECT 2732.865 1663.405 2734.075 1664.495 ;
        RECT 2695.520 1663.235 2734.160 1663.405 ;
        RECT 2695.605 1662.145 2696.815 1663.235 ;
        RECT 2696.985 1662.800 2702.330 1663.235 ;
        RECT 2702.505 1662.800 2707.850 1663.235 ;
        RECT 2696.295 1661.605 2696.815 1662.145 ;
        RECT 2700.390 1661.550 2700.740 1662.800 ;
        RECT 2705.910 1661.550 2706.260 1662.800 ;
        RECT 2708.485 1662.070 2708.775 1663.235 ;
        RECT 2708.945 1662.800 2714.290 1663.235 ;
        RECT 2714.465 1662.800 2719.810 1663.235 ;
        RECT 2719.985 1662.800 2725.330 1663.235 ;
        RECT 2725.505 1662.800 2730.850 1663.235 ;
        RECT 2712.350 1661.550 2712.700 1662.800 ;
        RECT 2717.870 1661.550 2718.220 1662.800 ;
        RECT 2723.390 1661.550 2723.740 1662.800 ;
        RECT 2728.910 1661.550 2729.260 1662.800 ;
        RECT 2731.025 1662.145 2732.695 1663.235 ;
        RECT 2731.945 1661.625 2732.695 1662.145 ;
        RECT 2732.865 1662.145 2734.075 1663.235 ;
        RECT 2732.865 1661.605 2733.385 1662.145 ;
        RECT 2696.295 1659.055 2696.815 1659.595 ;
        RECT 2695.605 1657.965 2696.815 1659.055 ;
        RECT 2710.050 1658.400 2710.400 1659.650 ;
        RECT 2715.570 1658.400 2715.920 1659.650 ;
        RECT 2719.505 1659.055 2721.195 1659.575 ;
        RECT 2697.415 1657.965 2697.745 1658.345 ;
        RECT 2700.135 1657.965 2700.465 1658.345 ;
        RECT 2701.960 1657.965 2702.290 1658.345 ;
        RECT 2702.880 1657.965 2703.230 1658.345 ;
        RECT 2705.715 1657.965 2706.045 1658.345 ;
        RECT 2706.645 1657.965 2711.990 1658.400 ;
        RECT 2712.165 1657.965 2717.510 1658.400 ;
        RECT 2717.685 1657.965 2721.195 1659.055 ;
        RECT 2721.365 1657.965 2721.655 1659.130 ;
        RECT 2725.230 1658.400 2725.580 1659.650 ;
        RECT 2730.750 1658.400 2731.100 1659.650 ;
        RECT 2732.865 1659.055 2733.385 1659.595 ;
        RECT 2721.825 1657.965 2727.170 1658.400 ;
        RECT 2727.345 1657.965 2732.690 1658.400 ;
        RECT 2732.865 1657.965 2734.075 1659.055 ;
        RECT 2695.520 1657.795 2734.160 1657.965 ;
        RECT 2695.605 1656.705 2696.815 1657.795 ;
        RECT 2697.425 1657.035 2697.755 1657.795 ;
        RECT 2698.365 1657.360 2703.710 1657.795 ;
        RECT 2696.295 1656.165 2696.815 1656.705 ;
        RECT 2701.770 1656.110 2702.120 1657.360 ;
        RECT 2703.885 1656.705 2707.395 1657.795 ;
        RECT 2705.705 1656.185 2707.395 1656.705 ;
        RECT 2708.485 1656.630 2708.775 1657.795 ;
        RECT 2708.945 1657.360 2714.290 1657.795 ;
        RECT 2714.465 1657.360 2719.810 1657.795 ;
        RECT 2719.985 1657.360 2725.330 1657.795 ;
        RECT 2725.505 1657.360 2730.850 1657.795 ;
        RECT 2712.350 1656.110 2712.700 1657.360 ;
        RECT 2717.870 1656.110 2718.220 1657.360 ;
        RECT 2723.390 1656.110 2723.740 1657.360 ;
        RECT 2728.910 1656.110 2729.260 1657.360 ;
        RECT 2731.025 1656.705 2732.695 1657.795 ;
        RECT 2731.945 1656.185 2732.695 1656.705 ;
        RECT 2732.865 1656.705 2734.075 1657.795 ;
        RECT 2732.865 1656.165 2733.385 1656.705 ;
        RECT 2696.295 1653.615 2696.815 1654.155 ;
        RECT 2695.605 1652.525 2696.815 1653.615 ;
        RECT 2710.050 1652.960 2710.400 1654.210 ;
        RECT 2715.570 1652.960 2715.920 1654.210 ;
        RECT 2719.505 1653.615 2721.195 1654.135 ;
        RECT 2697.415 1652.525 2697.745 1652.905 ;
        RECT 2700.135 1652.525 2700.465 1652.905 ;
        RECT 2701.960 1652.525 2702.290 1652.905 ;
        RECT 2702.880 1652.525 2703.230 1652.905 ;
        RECT 2705.715 1652.525 2706.045 1652.905 ;
        RECT 2706.645 1652.525 2711.990 1652.960 ;
        RECT 2712.165 1652.525 2717.510 1652.960 ;
        RECT 2717.685 1652.525 2721.195 1653.615 ;
        RECT 2721.365 1652.525 2721.655 1653.690 ;
        RECT 2725.230 1652.960 2725.580 1654.210 ;
        RECT 2730.750 1652.960 2731.100 1654.210 ;
        RECT 2732.865 1653.615 2733.385 1654.155 ;
        RECT 2721.825 1652.525 2727.170 1652.960 ;
        RECT 2727.345 1652.525 2732.690 1652.960 ;
        RECT 2732.865 1652.525 2734.075 1653.615 ;
        RECT 2695.520 1652.355 2734.160 1652.525 ;
        RECT 2695.605 1651.265 2696.815 1652.355 ;
        RECT 2697.425 1651.595 2697.755 1652.355 ;
        RECT 2698.365 1651.265 2700.955 1652.355 ;
        RECT 2696.295 1650.725 2696.815 1651.265 ;
        RECT 2699.745 1650.745 2700.955 1651.265 ;
        RECT 2702.095 1651.215 2702.265 1652.355 ;
        RECT 2704.635 1651.595 2704.805 1652.355 ;
        RECT 2705.725 1651.265 2708.315 1652.355 ;
        RECT 2707.105 1650.745 2708.315 1651.265 ;
        RECT 2708.485 1651.190 2708.775 1652.355 ;
        RECT 2708.945 1651.920 2714.290 1652.355 ;
        RECT 2714.465 1651.920 2719.810 1652.355 ;
        RECT 2719.985 1651.920 2725.330 1652.355 ;
        RECT 2725.505 1651.920 2730.850 1652.355 ;
        RECT 2712.350 1650.670 2712.700 1651.920 ;
        RECT 2717.870 1650.670 2718.220 1651.920 ;
        RECT 2723.390 1650.670 2723.740 1651.920 ;
        RECT 2728.910 1650.670 2729.260 1651.920 ;
        RECT 2731.025 1651.265 2732.695 1652.355 ;
        RECT 2731.945 1650.745 2732.695 1651.265 ;
        RECT 2732.865 1651.265 2734.075 1652.355 ;
        RECT 2732.865 1650.725 2733.385 1651.265 ;
        RECT 2696.295 1648.175 2696.815 1648.715 ;
        RECT 2695.605 1647.085 2696.815 1648.175 ;
        RECT 2700.390 1647.520 2700.740 1648.770 ;
        RECT 2705.910 1647.520 2706.260 1648.770 ;
        RECT 2711.430 1647.520 2711.780 1648.770 ;
        RECT 2716.950 1647.520 2717.300 1648.770 ;
        RECT 2719.985 1648.175 2720.735 1648.695 ;
        RECT 2696.985 1647.085 2702.330 1647.520 ;
        RECT 2702.505 1647.085 2707.850 1647.520 ;
        RECT 2708.025 1647.085 2713.370 1647.520 ;
        RECT 2713.545 1647.085 2718.890 1647.520 ;
        RECT 2719.065 1647.085 2720.735 1648.175 ;
        RECT 2721.365 1647.085 2721.655 1648.250 ;
        RECT 2725.230 1647.520 2725.580 1648.770 ;
        RECT 2730.750 1647.520 2731.100 1648.770 ;
        RECT 2732.865 1648.175 2733.385 1648.715 ;
        RECT 2721.825 1647.085 2727.170 1647.520 ;
        RECT 2727.345 1647.085 2732.690 1647.520 ;
        RECT 2732.865 1647.085 2734.075 1648.175 ;
        RECT 2695.520 1646.915 2734.160 1647.085 ;
        RECT 2695.605 1645.825 2696.815 1646.915 ;
        RECT 2697.425 1646.155 2697.755 1646.915 ;
        RECT 2698.365 1646.480 2703.710 1646.915 ;
        RECT 2696.295 1645.285 2696.815 1645.825 ;
        RECT 2701.770 1645.230 2702.120 1646.480 ;
        RECT 2703.885 1645.825 2707.395 1646.915 ;
        RECT 2705.705 1645.305 2707.395 1645.825 ;
        RECT 2708.485 1645.750 2708.775 1646.915 ;
        RECT 2708.945 1646.480 2714.290 1646.915 ;
        RECT 2714.465 1646.480 2719.810 1646.915 ;
        RECT 2719.985 1646.480 2725.330 1646.915 ;
        RECT 2725.505 1646.480 2730.850 1646.915 ;
        RECT 2712.350 1645.230 2712.700 1646.480 ;
        RECT 2717.870 1645.230 2718.220 1646.480 ;
        RECT 2723.390 1645.230 2723.740 1646.480 ;
        RECT 2728.910 1645.230 2729.260 1646.480 ;
        RECT 2731.025 1645.825 2732.695 1646.915 ;
        RECT 2731.945 1645.305 2732.695 1645.825 ;
        RECT 2732.865 1645.825 2734.075 1646.915 ;
        RECT 2732.865 1645.285 2733.385 1645.825 ;
        RECT 2696.295 1642.735 2696.815 1643.275 ;
        RECT 2695.605 1641.645 2696.815 1642.735 ;
        RECT 2700.390 1642.080 2700.740 1643.330 ;
        RECT 2705.910 1642.080 2706.260 1643.330 ;
        RECT 2711.430 1642.080 2711.780 1643.330 ;
        RECT 2716.950 1642.080 2717.300 1643.330 ;
        RECT 2719.985 1642.735 2720.735 1643.255 ;
        RECT 2696.985 1641.645 2702.330 1642.080 ;
        RECT 2702.505 1641.645 2707.850 1642.080 ;
        RECT 2708.025 1641.645 2713.370 1642.080 ;
        RECT 2713.545 1641.645 2718.890 1642.080 ;
        RECT 2719.065 1641.645 2720.735 1642.735 ;
        RECT 2721.365 1641.645 2721.655 1642.810 ;
        RECT 2725.230 1642.080 2725.580 1643.330 ;
        RECT 2730.750 1642.080 2731.100 1643.330 ;
        RECT 2732.865 1642.735 2733.385 1643.275 ;
        RECT 2721.825 1641.645 2727.170 1642.080 ;
        RECT 2727.345 1641.645 2732.690 1642.080 ;
        RECT 2732.865 1641.645 2734.075 1642.735 ;
        RECT 2695.520 1641.475 2734.160 1641.645 ;
        RECT 2695.605 1640.385 2696.815 1641.475 ;
        RECT 2696.985 1640.385 2700.495 1641.475 ;
        RECT 2696.295 1639.845 2696.815 1640.385 ;
        RECT 2698.805 1639.865 2700.495 1640.385 ;
        RECT 2702.455 1640.335 2702.785 1641.475 ;
        RECT 2702.965 1641.040 2708.310 1641.475 ;
        RECT 2706.370 1639.790 2706.720 1641.040 ;
        RECT 2708.485 1640.310 2708.775 1641.475 ;
        RECT 2708.945 1641.040 2714.290 1641.475 ;
        RECT 2714.465 1641.040 2719.810 1641.475 ;
        RECT 2719.985 1641.040 2725.330 1641.475 ;
        RECT 2725.505 1641.040 2730.850 1641.475 ;
        RECT 2712.350 1639.790 2712.700 1641.040 ;
        RECT 2717.870 1639.790 2718.220 1641.040 ;
        RECT 2723.390 1639.790 2723.740 1641.040 ;
        RECT 2728.910 1639.790 2729.260 1641.040 ;
        RECT 2731.025 1640.385 2732.695 1641.475 ;
        RECT 2731.945 1639.865 2732.695 1640.385 ;
        RECT 2732.865 1640.385 2734.075 1641.475 ;
        RECT 2732.865 1639.845 2733.385 1640.385 ;
        RECT 2696.295 1637.295 2696.815 1637.835 ;
        RECT 2700.185 1637.295 2701.875 1637.815 ;
        RECT 2695.605 1636.205 2696.815 1637.295 ;
        RECT 2697.425 1636.205 2697.755 1636.965 ;
        RECT 2698.365 1636.205 2701.875 1637.295 ;
        RECT 2703.535 1636.205 2703.705 1636.645 ;
        RECT 2708.670 1636.640 2709.020 1637.890 ;
        RECT 2714.190 1636.640 2714.540 1637.890 ;
        RECT 2718.125 1637.295 2719.815 1637.815 ;
        RECT 2720.675 1637.295 2721.195 1637.835 ;
        RECT 2704.310 1636.205 2704.640 1636.565 ;
        RECT 2705.265 1636.205 2710.610 1636.640 ;
        RECT 2710.785 1636.205 2716.130 1636.640 ;
        RECT 2716.305 1636.205 2719.815 1637.295 ;
        RECT 2719.985 1636.205 2721.195 1637.295 ;
        RECT 2721.365 1636.205 2721.655 1637.370 ;
        RECT 2725.230 1636.640 2725.580 1637.890 ;
        RECT 2730.750 1636.640 2731.100 1637.890 ;
        RECT 2732.865 1637.295 2733.385 1637.835 ;
        RECT 2721.825 1636.205 2727.170 1636.640 ;
        RECT 2727.345 1636.205 2732.690 1636.640 ;
        RECT 2732.865 1636.205 2734.075 1637.295 ;
        RECT 2695.520 1636.035 2734.160 1636.205 ;
        RECT 2695.605 1634.945 2696.815 1636.035 ;
        RECT 2696.985 1635.600 2702.330 1636.035 ;
        RECT 2702.505 1635.600 2707.850 1636.035 ;
        RECT 2696.295 1634.405 2696.815 1634.945 ;
        RECT 2700.390 1634.350 2700.740 1635.600 ;
        RECT 2705.910 1634.350 2706.260 1635.600 ;
        RECT 2708.485 1634.870 2708.775 1636.035 ;
        RECT 2708.945 1635.600 2714.290 1636.035 ;
        RECT 2714.465 1635.600 2719.810 1636.035 ;
        RECT 2719.985 1635.600 2725.330 1636.035 ;
        RECT 2712.350 1634.350 2712.700 1635.600 ;
        RECT 2717.870 1634.350 2718.220 1635.600 ;
        RECT 2723.390 1634.350 2723.740 1635.600 ;
        RECT 2725.595 1635.235 2725.765 1636.035 ;
        RECT 2726.435 1635.235 2726.605 1636.035 ;
        RECT 2727.275 1635.235 2727.445 1636.035 ;
        RECT 2728.035 1635.235 2728.365 1636.035 ;
        RECT 2728.875 1635.235 2729.205 1636.035 ;
        RECT 2729.715 1635.235 2730.045 1636.035 ;
        RECT 2730.555 1635.235 2730.885 1636.035 ;
        RECT 2731.395 1635.235 2731.725 1636.035 ;
        RECT 2732.235 1634.885 2732.565 1636.035 ;
        RECT 2732.865 1634.945 2734.075 1636.035 ;
        RECT 2732.865 1634.405 2733.385 1634.945 ;
        RECT 2696.295 1631.855 2696.815 1632.395 ;
        RECT 2695.605 1630.765 2696.815 1631.855 ;
        RECT 2697.425 1630.765 2697.755 1631.525 ;
        RECT 2701.770 1631.200 2702.120 1632.450 ;
        RECT 2707.290 1631.200 2707.640 1632.450 ;
        RECT 2712.810 1631.200 2713.160 1632.450 ;
        RECT 2718.330 1631.200 2718.680 1632.450 ;
        RECT 2698.365 1630.765 2703.710 1631.200 ;
        RECT 2703.885 1630.765 2709.230 1631.200 ;
        RECT 2709.405 1630.765 2714.750 1631.200 ;
        RECT 2714.925 1630.765 2720.270 1631.200 ;
        RECT 2721.365 1630.765 2721.655 1631.930 ;
        RECT 2725.230 1631.200 2725.580 1632.450 ;
        RECT 2730.750 1631.200 2731.100 1632.450 ;
        RECT 2732.865 1631.855 2733.385 1632.395 ;
        RECT 2721.825 1630.765 2727.170 1631.200 ;
        RECT 2727.345 1630.765 2732.690 1631.200 ;
        RECT 2732.865 1630.765 2734.075 1631.855 ;
        RECT 2695.520 1630.595 2734.160 1630.765 ;
        RECT 2695.605 1629.505 2696.815 1630.595 ;
        RECT 2696.985 1630.160 2702.330 1630.595 ;
        RECT 2702.505 1630.160 2707.850 1630.595 ;
        RECT 2696.295 1628.965 2696.815 1629.505 ;
        RECT 2700.390 1628.910 2700.740 1630.160 ;
        RECT 2705.910 1628.910 2706.260 1630.160 ;
        RECT 2708.485 1629.430 2708.775 1630.595 ;
        RECT 2708.945 1630.160 2714.290 1630.595 ;
        RECT 2714.465 1630.160 2719.810 1630.595 ;
        RECT 2719.985 1630.160 2725.330 1630.595 ;
        RECT 2725.505 1630.160 2730.850 1630.595 ;
        RECT 2712.350 1628.910 2712.700 1630.160 ;
        RECT 2717.870 1628.910 2718.220 1630.160 ;
        RECT 2723.390 1628.910 2723.740 1630.160 ;
        RECT 2728.910 1628.910 2729.260 1630.160 ;
        RECT 2731.025 1629.505 2732.695 1630.595 ;
        RECT 2731.945 1628.985 2732.695 1629.505 ;
        RECT 2732.865 1629.505 2734.075 1630.595 ;
        RECT 2732.865 1628.965 2733.385 1629.505 ;
        RECT 2881.580 1628.340 2883.380 1628.510 ;
        RECT 2882.775 1627.615 2883.105 1628.340 ;
        RECT 2696.295 1626.415 2696.815 1626.955 ;
        RECT 2522.135 1626.230 2523.935 1626.400 ;
        RECT 2522.830 1625.505 2523.160 1626.230 ;
        RECT 2695.605 1625.325 2696.815 1626.415 ;
        RECT 2697.715 1625.325 2698.045 1625.835 ;
        RECT 2703.150 1625.760 2703.500 1627.010 ;
        RECT 2708.670 1625.760 2709.020 1627.010 ;
        RECT 2714.190 1625.760 2714.540 1627.010 ;
        RECT 2718.125 1626.415 2719.815 1626.935 ;
        RECT 2720.675 1626.415 2721.195 1626.955 ;
        RECT 2699.745 1625.325 2705.090 1625.760 ;
        RECT 2705.265 1625.325 2710.610 1625.760 ;
        RECT 2710.785 1625.325 2716.130 1625.760 ;
        RECT 2716.305 1625.325 2719.815 1626.415 ;
        RECT 2719.985 1625.325 2721.195 1626.415 ;
        RECT 2721.365 1625.325 2721.655 1626.490 ;
        RECT 2725.230 1625.760 2725.580 1627.010 ;
        RECT 2730.750 1625.760 2731.100 1627.010 ;
        RECT 2732.865 1626.415 2733.385 1626.955 ;
        RECT 2721.825 1625.325 2727.170 1625.760 ;
        RECT 2727.345 1625.325 2732.690 1625.760 ;
        RECT 2732.865 1625.325 2734.075 1626.415 ;
        RECT 2695.520 1625.155 2734.160 1625.325 ;
        RECT 2695.605 1624.065 2696.815 1625.155 ;
        RECT 2697.425 1624.395 2697.755 1625.155 ;
        RECT 2698.365 1624.720 2703.710 1625.155 ;
        RECT 2696.295 1623.525 2696.815 1624.065 ;
        RECT 2701.770 1623.470 2702.120 1624.720 ;
        RECT 2703.885 1624.065 2707.395 1625.155 ;
        RECT 2705.705 1623.545 2707.395 1624.065 ;
        RECT 2708.485 1623.990 2708.775 1625.155 ;
        RECT 2708.945 1624.720 2714.290 1625.155 ;
        RECT 2714.465 1624.720 2719.810 1625.155 ;
        RECT 2719.985 1624.720 2725.330 1625.155 ;
        RECT 2725.505 1624.720 2730.850 1625.155 ;
        RECT 2712.350 1623.470 2712.700 1624.720 ;
        RECT 2717.870 1623.470 2718.220 1624.720 ;
        RECT 2723.390 1623.470 2723.740 1624.720 ;
        RECT 2728.910 1623.470 2729.260 1624.720 ;
        RECT 2731.025 1624.065 2732.695 1625.155 ;
        RECT 2731.945 1623.545 2732.695 1624.065 ;
        RECT 2732.865 1624.065 2734.075 1625.155 ;
        RECT 2732.865 1623.525 2733.385 1624.065 ;
        RECT 2696.295 1620.975 2696.815 1621.515 ;
        RECT 2522.135 1619.815 2523.935 1619.985 ;
        RECT 2695.605 1619.885 2696.815 1620.975 ;
        RECT 2697.735 1619.885 2697.905 1620.645 ;
        RECT 2700.275 1619.885 2700.445 1621.025 ;
        RECT 2701.590 1619.885 2701.920 1620.600 ;
        RECT 2708.210 1620.320 2708.560 1621.570 ;
        RECT 2713.730 1620.320 2714.080 1621.570 ;
        RECT 2719.250 1620.320 2719.600 1621.570 ;
        RECT 2704.805 1619.885 2710.150 1620.320 ;
        RECT 2710.325 1619.885 2715.670 1620.320 ;
        RECT 2715.845 1619.885 2721.190 1620.320 ;
        RECT 2721.365 1619.885 2721.655 1621.050 ;
        RECT 2725.230 1620.320 2725.580 1621.570 ;
        RECT 2730.750 1620.320 2731.100 1621.570 ;
        RECT 2732.865 1620.975 2733.385 1621.515 ;
        RECT 2721.825 1619.885 2727.170 1620.320 ;
        RECT 2727.345 1619.885 2732.690 1620.320 ;
        RECT 2732.865 1619.885 2734.075 1620.975 ;
        RECT 2522.830 1619.090 2523.160 1619.815 ;
        RECT 2695.520 1619.715 2734.160 1619.885 ;
        RECT 2695.605 1618.625 2696.815 1619.715 ;
        RECT 2696.985 1619.205 2697.245 1619.715 ;
        RECT 2697.905 1619.210 2698.520 1619.715 ;
        RECT 2698.325 1619.035 2698.520 1619.210 ;
        RECT 2699.335 1619.170 2699.550 1619.715 ;
        RECT 2700.205 1619.280 2705.550 1619.715 ;
        RECT 2698.325 1618.845 2698.655 1619.035 ;
        RECT 2696.295 1618.085 2696.815 1618.625 ;
        RECT 2703.610 1618.030 2703.960 1619.280 ;
        RECT 2705.725 1618.625 2708.315 1619.715 ;
        RECT 2707.105 1618.105 2708.315 1618.625 ;
        RECT 2708.485 1618.550 2708.775 1619.715 ;
        RECT 2708.945 1619.280 2714.290 1619.715 ;
        RECT 2714.465 1619.280 2719.810 1619.715 ;
        RECT 2719.985 1619.280 2725.330 1619.715 ;
        RECT 2725.505 1619.280 2730.850 1619.715 ;
        RECT 2712.350 1618.030 2712.700 1619.280 ;
        RECT 2717.870 1618.030 2718.220 1619.280 ;
        RECT 2723.390 1618.030 2723.740 1619.280 ;
        RECT 2728.910 1618.030 2729.260 1619.280 ;
        RECT 2731.025 1618.625 2732.695 1619.715 ;
        RECT 2731.945 1618.105 2732.695 1618.625 ;
        RECT 2732.865 1618.625 2734.075 1619.715 ;
        RECT 2732.865 1618.085 2733.385 1618.625 ;
        RECT 2696.295 1615.535 2696.815 1616.075 ;
        RECT 2695.605 1614.445 2696.815 1615.535 ;
        RECT 2697.425 1614.445 2697.755 1615.205 ;
        RECT 2701.770 1614.880 2702.120 1616.130 ;
        RECT 2707.290 1614.880 2707.640 1616.130 ;
        RECT 2712.810 1614.880 2713.160 1616.130 ;
        RECT 2718.330 1614.880 2718.680 1616.130 ;
        RECT 2698.365 1614.445 2703.710 1614.880 ;
        RECT 2703.885 1614.445 2709.230 1614.880 ;
        RECT 2709.405 1614.445 2714.750 1614.880 ;
        RECT 2714.925 1614.445 2720.270 1614.880 ;
        RECT 2721.365 1614.445 2721.655 1615.610 ;
        RECT 2725.230 1614.880 2725.580 1616.130 ;
        RECT 2730.750 1614.880 2731.100 1616.130 ;
        RECT 2732.865 1615.535 2733.385 1616.075 ;
        RECT 2721.825 1614.445 2727.170 1614.880 ;
        RECT 2727.345 1614.445 2732.690 1614.880 ;
        RECT 2732.865 1614.445 2734.075 1615.535 ;
        RECT 2695.520 1614.275 2734.160 1614.445 ;
        RECT 2695.605 1613.185 2696.815 1614.275 ;
        RECT 2696.985 1613.185 2698.195 1614.275 ;
        RECT 2698.865 1613.815 2699.115 1614.275 ;
        RECT 2699.795 1613.815 2700.045 1614.275 ;
        RECT 2701.115 1613.815 2701.365 1614.275 ;
        RECT 2702.045 1613.840 2707.390 1614.275 ;
        RECT 2696.295 1612.645 2696.815 1613.185 ;
        RECT 2697.675 1612.645 2698.195 1613.185 ;
        RECT 2705.450 1612.590 2705.800 1613.840 ;
        RECT 2708.485 1613.110 2708.775 1614.275 ;
        RECT 2708.945 1613.840 2714.290 1614.275 ;
        RECT 2714.465 1613.840 2719.810 1614.275 ;
        RECT 2719.985 1613.840 2725.330 1614.275 ;
        RECT 2725.505 1613.840 2730.850 1614.275 ;
        RECT 2712.350 1612.590 2712.700 1613.840 ;
        RECT 2717.870 1612.590 2718.220 1613.840 ;
        RECT 2723.390 1612.590 2723.740 1613.840 ;
        RECT 2728.910 1612.590 2729.260 1613.840 ;
        RECT 2731.025 1613.185 2732.695 1614.275 ;
        RECT 2731.945 1612.665 2732.695 1613.185 ;
        RECT 2732.865 1613.185 2734.075 1614.275 ;
        RECT 2732.865 1612.645 2733.385 1613.185 ;
        RECT 2360.030 1610.045 2360.205 1610.595 ;
        RECT 2696.295 1610.095 2696.815 1610.635 ;
        RECT 2360.030 1608.445 2360.200 1610.045 ;
        RECT 2695.605 1609.005 2696.815 1610.095 ;
        RECT 2697.905 1609.005 2698.165 1610.145 ;
        RECT 2700.190 1609.005 2700.470 1609.805 ;
        RECT 2701.885 1609.005 2702.170 1609.805 ;
        RECT 2702.840 1609.005 2703.090 1610.145 ;
        RECT 2707.290 1609.440 2707.640 1610.690 ;
        RECT 2712.810 1609.440 2713.160 1610.690 ;
        RECT 2718.330 1609.440 2718.680 1610.690 ;
        RECT 2703.885 1609.005 2709.230 1609.440 ;
        RECT 2709.405 1609.005 2714.750 1609.440 ;
        RECT 2714.925 1609.005 2720.270 1609.440 ;
        RECT 2721.365 1609.005 2721.655 1610.170 ;
        RECT 2725.230 1609.440 2725.580 1610.690 ;
        RECT 2730.750 1609.440 2731.100 1610.690 ;
        RECT 2732.865 1610.095 2733.385 1610.635 ;
        RECT 2721.825 1609.005 2727.170 1609.440 ;
        RECT 2727.345 1609.005 2732.690 1609.440 ;
        RECT 2732.865 1609.005 2734.075 1610.095 ;
        RECT 2695.520 1608.835 2734.160 1609.005 ;
        RECT 2358.215 1607.035 2358.385 1607.765 ;
        RECT 2360.030 1607.305 2360.205 1608.445 ;
        RECT 2360.030 1607.035 2360.200 1607.305 ;
        RECT 2361.625 1607.035 2361.795 1607.765 ;
        RECT 2373.310 1607.035 2373.480 1607.765 ;
        RECT 2376.055 1607.035 2376.225 1607.765 ;
        RECT 2377.045 1607.035 2377.215 1607.765 ;
        RECT 2378.845 1607.035 2379.015 1607.765 ;
        RECT 2390.530 1607.035 2390.700 1607.765 ;
        RECT 2393.275 1607.035 2393.445 1607.765 ;
        RECT 2394.265 1607.035 2394.435 1607.765 ;
        RECT 2396.065 1607.040 2396.235 1607.770 ;
        RECT 2407.750 1607.040 2407.920 1607.770 ;
        RECT 2410.495 1607.040 2410.665 1607.770 ;
        RECT 2411.485 1607.040 2411.655 1607.770 ;
        RECT 2358.045 1607.025 2360.795 1607.035 ;
        RECT 2361.455 1607.025 2364.205 1607.035 ;
        RECT 2373.140 1607.030 2377.865 1607.035 ;
        RECT 2378.675 1607.030 2381.425 1607.035 ;
        RECT 2390.360 1607.030 2395.085 1607.035 ;
        RECT 2395.895 1607.030 2398.645 1607.040 ;
        RECT 2407.580 1607.035 2412.305 1607.040 ;
        RECT 2413.285 1607.035 2413.455 1607.765 ;
        RECT 2424.970 1607.035 2425.140 1607.765 ;
        RECT 2427.715 1607.035 2427.885 1607.765 ;
        RECT 2428.705 1607.035 2428.875 1607.765 ;
        RECT 2430.505 1607.035 2430.675 1607.765 ;
        RECT 2442.190 1607.035 2442.360 1607.765 ;
        RECT 2444.935 1607.035 2445.105 1607.765 ;
        RECT 2445.925 1607.035 2446.095 1607.765 ;
        RECT 2695.605 1607.745 2696.815 1608.835 ;
        RECT 2697.425 1608.075 2697.755 1608.835 ;
        RECT 2696.295 1607.205 2696.815 1607.745 ;
        RECT 2698.825 1607.695 2699.085 1608.835 ;
        RECT 2699.755 1607.695 2700.035 1608.835 ;
        RECT 2700.205 1608.400 2705.550 1608.835 ;
        RECT 2703.610 1607.150 2703.960 1608.400 ;
        RECT 2705.725 1607.745 2708.315 1608.835 ;
        RECT 2707.105 1607.225 2708.315 1607.745 ;
        RECT 2708.485 1607.670 2708.775 1608.835 ;
        RECT 2708.945 1608.400 2714.290 1608.835 ;
        RECT 2714.465 1608.400 2719.810 1608.835 ;
        RECT 2719.985 1608.400 2725.330 1608.835 ;
        RECT 2725.505 1608.400 2730.850 1608.835 ;
        RECT 2712.350 1607.150 2712.700 1608.400 ;
        RECT 2717.870 1607.150 2718.220 1608.400 ;
        RECT 2723.390 1607.150 2723.740 1608.400 ;
        RECT 2728.910 1607.150 2729.260 1608.400 ;
        RECT 2731.025 1607.745 2732.695 1608.835 ;
        RECT 2731.945 1607.225 2732.695 1607.745 ;
        RECT 2732.865 1607.745 2734.075 1608.835 ;
        RECT 2732.865 1607.205 2733.385 1607.745 ;
        RECT 2406.475 1607.030 2412.460 1607.035 ;
        RECT 2413.115 1607.030 2415.865 1607.035 ;
        RECT 2424.800 1607.030 2429.525 1607.035 ;
        RECT 2430.335 1607.030 2433.085 1607.035 ;
        RECT 2442.020 1607.030 2446.745 1607.035 ;
        RECT 2343.000 1607.000 2364.470 1607.025 ;
        RECT 2372.035 1607.005 2381.580 1607.030 ;
        RECT 2343.000 1606.800 2364.940 1607.000 ;
        RECT 2343.000 1605.810 2364.945 1606.800 ;
        RECT 2365.130 1605.810 2365.410 1606.950 ;
        RECT 2366.080 1605.810 2366.340 1606.950 ;
        RECT 2367.430 1605.810 2367.710 1606.950 ;
        RECT 2368.380 1605.810 2368.640 1606.950 ;
        RECT 2368.810 1605.810 2369.070 1606.950 ;
        RECT 2369.740 1605.810 2370.020 1606.950 ;
        RECT 2370.190 1605.810 2370.450 1606.950 ;
        RECT 2371.120 1605.810 2371.400 1606.950 ;
        RECT 2372.035 1606.800 2381.585 1607.005 ;
        RECT 2371.935 1605.810 2382.165 1606.800 ;
        RECT 2382.350 1605.810 2382.630 1606.950 ;
        RECT 2383.300 1605.810 2383.560 1606.950 ;
        RECT 2384.650 1605.810 2384.930 1606.950 ;
        RECT 2385.600 1605.810 2385.860 1606.950 ;
        RECT 2386.030 1605.810 2386.290 1606.950 ;
        RECT 2386.960 1605.810 2387.240 1606.950 ;
        RECT 2387.410 1605.810 2387.670 1606.950 ;
        RECT 2388.340 1605.810 2388.620 1606.950 ;
        RECT 2389.255 1606.805 2398.805 1607.030 ;
        RECT 2389.255 1606.800 2399.385 1606.805 ;
        RECT 2389.155 1605.815 2399.385 1606.800 ;
        RECT 2399.570 1605.815 2399.850 1606.955 ;
        RECT 2400.520 1605.815 2400.780 1606.955 ;
        RECT 2401.870 1605.815 2402.150 1606.955 ;
        RECT 2402.820 1605.815 2403.080 1606.955 ;
        RECT 2403.250 1605.815 2403.510 1606.955 ;
        RECT 2404.180 1605.815 2404.460 1606.955 ;
        RECT 2404.630 1605.815 2404.890 1606.955 ;
        RECT 2405.560 1605.815 2405.840 1606.955 ;
        RECT 2406.475 1606.805 2416.025 1607.030 ;
        RECT 2406.375 1606.800 2416.025 1606.805 ;
        RECT 2406.375 1605.815 2416.605 1606.800 ;
        RECT 2389.155 1605.810 2416.605 1605.815 ;
        RECT 2416.790 1605.810 2417.070 1606.950 ;
        RECT 2417.740 1605.810 2418.000 1606.950 ;
        RECT 2419.090 1605.810 2419.370 1606.950 ;
        RECT 2420.040 1605.810 2420.300 1606.950 ;
        RECT 2420.470 1605.810 2420.730 1606.950 ;
        RECT 2421.400 1605.810 2421.680 1606.950 ;
        RECT 2421.850 1605.810 2422.110 1606.950 ;
        RECT 2422.780 1605.810 2423.060 1606.950 ;
        RECT 2423.695 1606.800 2433.245 1607.030 ;
        RECT 2423.595 1605.810 2433.825 1606.800 ;
        RECT 2434.010 1605.810 2434.290 1606.950 ;
        RECT 2434.960 1605.810 2435.220 1606.950 ;
        RECT 2436.310 1605.810 2436.590 1606.950 ;
        RECT 2437.260 1605.810 2437.520 1606.950 ;
        RECT 2437.690 1605.810 2437.950 1606.950 ;
        RECT 2438.620 1605.810 2438.900 1606.950 ;
        RECT 2439.070 1605.810 2439.330 1606.950 ;
        RECT 2440.000 1605.810 2440.280 1606.950 ;
        RECT 2440.915 1606.800 2446.900 1607.030 ;
        RECT 2440.815 1605.810 2446.900 1606.800 ;
        RECT 2343.000 1605.645 2446.900 1605.810 ;
        RECT 2343.000 1605.640 2399.380 1605.645 ;
        RECT 2343.000 1605.425 2364.940 1605.640 ;
        RECT 2364.730 1604.500 2364.940 1605.425 ;
        RECT 2365.610 1604.500 2365.840 1605.640 ;
        RECT 2366.060 1604.500 2366.390 1605.640 ;
        RECT 2368.300 1604.500 2368.630 1605.640 ;
        RECT 2369.880 1605.130 2370.050 1605.640 ;
        RECT 2370.720 1604.790 2370.890 1605.640 ;
        RECT 2372.030 1605.430 2382.160 1605.640 ;
        RECT 2373.140 1605.425 2382.160 1605.430 ;
        RECT 2373.310 1604.695 2373.480 1605.425 ;
        RECT 2376.055 1604.695 2376.225 1605.425 ;
        RECT 2377.040 1604.695 2377.210 1605.425 ;
        RECT 2381.950 1604.500 2382.160 1605.425 ;
        RECT 2382.830 1604.500 2383.060 1605.640 ;
        RECT 2383.280 1604.500 2383.610 1605.640 ;
        RECT 2385.520 1604.500 2385.850 1605.640 ;
        RECT 2387.100 1605.130 2387.270 1605.640 ;
        RECT 2387.940 1604.790 2388.110 1605.640 ;
        RECT 2389.250 1605.430 2399.380 1605.640 ;
        RECT 2390.360 1605.425 2395.080 1605.430 ;
        RECT 2390.530 1604.695 2390.700 1605.425 ;
        RECT 2393.275 1604.695 2393.445 1605.425 ;
        RECT 2394.260 1604.695 2394.430 1605.425 ;
        RECT 2399.170 1604.505 2399.380 1605.430 ;
        RECT 2400.050 1604.505 2400.280 1605.645 ;
        RECT 2400.500 1604.505 2400.830 1605.645 ;
        RECT 2402.740 1604.505 2403.070 1605.645 ;
        RECT 2404.320 1605.135 2404.490 1605.645 ;
        RECT 2405.160 1604.795 2405.330 1605.645 ;
        RECT 2406.470 1605.640 2446.900 1605.645 ;
        RECT 2406.470 1605.435 2416.600 1605.640 ;
        RECT 2406.475 1605.430 2416.600 1605.435 ;
        RECT 2407.750 1604.700 2407.920 1605.430 ;
        RECT 2410.495 1604.700 2410.665 1605.430 ;
        RECT 2411.480 1604.700 2411.650 1605.430 ;
        RECT 2412.455 1605.425 2416.600 1605.430 ;
        RECT 2416.390 1604.500 2416.600 1605.425 ;
        RECT 2417.270 1604.500 2417.500 1605.640 ;
        RECT 2417.720 1604.500 2418.050 1605.640 ;
        RECT 2419.960 1604.500 2420.290 1605.640 ;
        RECT 2421.540 1605.130 2421.710 1605.640 ;
        RECT 2422.380 1604.790 2422.550 1605.640 ;
        RECT 2423.690 1605.430 2433.820 1605.640 ;
        RECT 2424.800 1605.425 2433.820 1605.430 ;
        RECT 2424.970 1604.695 2425.140 1605.425 ;
        RECT 2427.715 1604.695 2427.885 1605.425 ;
        RECT 2428.700 1604.695 2428.870 1605.425 ;
        RECT 2433.610 1604.500 2433.820 1605.425 ;
        RECT 2434.490 1604.500 2434.720 1605.640 ;
        RECT 2434.940 1604.500 2435.270 1605.640 ;
        RECT 2437.180 1604.500 2437.510 1605.640 ;
        RECT 2438.760 1605.130 2438.930 1605.640 ;
        RECT 2439.600 1604.790 2439.770 1605.640 ;
        RECT 2440.910 1605.430 2446.900 1605.640 ;
        RECT 2442.020 1605.425 2446.740 1605.430 ;
        RECT 2442.190 1604.695 2442.360 1605.425 ;
        RECT 2444.935 1604.695 2445.105 1605.425 ;
        RECT 2445.920 1604.695 2446.090 1605.425 ;
        RECT 2696.295 1604.655 2696.815 1605.195 ;
        RECT 2695.605 1603.565 2696.815 1604.655 ;
        RECT 2697.735 1603.565 2697.905 1604.325 ;
        RECT 2700.275 1603.565 2700.445 1604.705 ;
        RECT 2704.530 1604.000 2704.880 1605.250 ;
        RECT 2710.050 1604.000 2710.400 1605.250 ;
        RECT 2715.570 1604.000 2715.920 1605.250 ;
        RECT 2719.505 1604.655 2721.195 1605.175 ;
        RECT 2701.125 1603.565 2706.470 1604.000 ;
        RECT 2706.645 1603.565 2711.990 1604.000 ;
        RECT 2712.165 1603.565 2717.510 1604.000 ;
        RECT 2717.685 1603.565 2721.195 1604.655 ;
        RECT 2721.365 1603.565 2721.655 1604.730 ;
        RECT 2725.230 1604.000 2725.580 1605.250 ;
        RECT 2730.750 1604.000 2731.100 1605.250 ;
        RECT 2732.865 1604.655 2733.385 1605.195 ;
        RECT 2721.825 1603.565 2727.170 1604.000 ;
        RECT 2727.345 1603.565 2732.690 1604.000 ;
        RECT 2732.865 1603.565 2734.075 1604.655 ;
        RECT 2695.520 1603.395 2734.160 1603.565 ;
        RECT 2695.605 1602.305 2696.815 1603.395 ;
        RECT 2697.425 1602.635 2697.755 1603.395 ;
        RECT 2698.365 1602.960 2703.710 1603.395 ;
        RECT 2696.295 1601.765 2696.815 1602.305 ;
        RECT 2701.770 1601.710 2702.120 1602.960 ;
        RECT 2703.885 1602.305 2707.395 1603.395 ;
        RECT 2705.705 1601.785 2707.395 1602.305 ;
        RECT 2708.485 1602.230 2708.775 1603.395 ;
        RECT 2708.945 1602.960 2714.290 1603.395 ;
        RECT 2714.465 1602.960 2719.810 1603.395 ;
        RECT 2719.985 1602.960 2725.330 1603.395 ;
        RECT 2725.505 1602.960 2730.850 1603.395 ;
        RECT 2712.350 1601.710 2712.700 1602.960 ;
        RECT 2717.870 1601.710 2718.220 1602.960 ;
        RECT 2723.390 1601.710 2723.740 1602.960 ;
        RECT 2728.910 1601.710 2729.260 1602.960 ;
        RECT 2731.025 1602.305 2732.695 1603.395 ;
        RECT 2731.945 1601.785 2732.695 1602.305 ;
        RECT 2732.865 1602.305 2734.075 1603.395 ;
        RECT 2732.865 1601.765 2733.385 1602.305 ;
        RECT 2696.295 1599.215 2696.815 1599.755 ;
        RECT 2695.605 1598.125 2696.815 1599.215 ;
        RECT 2700.390 1598.560 2700.740 1599.810 ;
        RECT 2705.910 1598.560 2706.260 1599.810 ;
        RECT 2711.430 1598.560 2711.780 1599.810 ;
        RECT 2716.950 1598.560 2717.300 1599.810 ;
        RECT 2719.985 1599.215 2720.735 1599.735 ;
        RECT 2696.985 1598.125 2702.330 1598.560 ;
        RECT 2702.505 1598.125 2707.850 1598.560 ;
        RECT 2708.025 1598.125 2713.370 1598.560 ;
        RECT 2713.545 1598.125 2718.890 1598.560 ;
        RECT 2719.065 1598.125 2720.735 1599.215 ;
        RECT 2721.365 1598.125 2721.655 1599.290 ;
        RECT 2725.230 1598.560 2725.580 1599.810 ;
        RECT 2730.750 1598.560 2731.100 1599.810 ;
        RECT 2732.865 1599.215 2733.385 1599.755 ;
        RECT 2721.825 1598.125 2727.170 1598.560 ;
        RECT 2727.345 1598.125 2732.690 1598.560 ;
        RECT 2732.865 1598.125 2734.075 1599.215 ;
        RECT 2695.520 1597.955 2734.160 1598.125 ;
        RECT 2695.605 1596.865 2696.815 1597.955 ;
        RECT 2697.425 1597.195 2697.755 1597.955 ;
        RECT 2698.365 1597.520 2703.710 1597.955 ;
        RECT 2696.295 1596.325 2696.815 1596.865 ;
        RECT 2701.770 1596.270 2702.120 1597.520 ;
        RECT 2703.885 1596.865 2707.395 1597.955 ;
        RECT 2705.705 1596.345 2707.395 1596.865 ;
        RECT 2708.485 1596.790 2708.775 1597.955 ;
        RECT 2708.945 1597.520 2714.290 1597.955 ;
        RECT 2714.465 1597.520 2719.810 1597.955 ;
        RECT 2719.985 1597.520 2725.330 1597.955 ;
        RECT 2725.505 1597.520 2730.850 1597.955 ;
        RECT 2712.350 1596.270 2712.700 1597.520 ;
        RECT 2717.870 1596.270 2718.220 1597.520 ;
        RECT 2723.390 1596.270 2723.740 1597.520 ;
        RECT 2728.910 1596.270 2729.260 1597.520 ;
        RECT 2731.025 1596.865 2732.695 1597.955 ;
        RECT 2731.945 1596.345 2732.695 1596.865 ;
        RECT 2732.865 1596.865 2734.075 1597.955 ;
        RECT 2732.865 1596.325 2733.385 1596.865 ;
        RECT 2696.295 1593.775 2696.815 1594.315 ;
        RECT 2695.605 1592.685 2696.815 1593.775 ;
        RECT 2700.390 1593.120 2700.740 1594.370 ;
        RECT 2705.910 1593.120 2706.260 1594.370 ;
        RECT 2711.430 1593.120 2711.780 1594.370 ;
        RECT 2716.950 1593.120 2717.300 1594.370 ;
        RECT 2719.985 1593.775 2720.735 1594.295 ;
        RECT 2696.985 1592.685 2702.330 1593.120 ;
        RECT 2702.505 1592.685 2707.850 1593.120 ;
        RECT 2708.025 1592.685 2713.370 1593.120 ;
        RECT 2713.545 1592.685 2718.890 1593.120 ;
        RECT 2719.065 1592.685 2720.735 1593.775 ;
        RECT 2721.365 1592.685 2721.655 1593.850 ;
        RECT 2725.230 1593.120 2725.580 1594.370 ;
        RECT 2730.750 1593.120 2731.100 1594.370 ;
        RECT 2732.865 1593.775 2733.385 1594.315 ;
        RECT 2721.825 1592.685 2727.170 1593.120 ;
        RECT 2727.345 1592.685 2732.690 1593.120 ;
        RECT 2732.865 1592.685 2734.075 1593.775 ;
        RECT 2695.520 1592.515 2734.160 1592.685 ;
        RECT 2695.605 1591.425 2696.815 1592.515 ;
        RECT 2697.425 1591.755 2697.755 1592.515 ;
        RECT 2698.805 1591.755 2699.135 1592.515 ;
        RECT 2699.745 1592.080 2705.090 1592.515 ;
        RECT 2696.295 1590.885 2696.815 1591.425 ;
        RECT 2703.150 1590.830 2703.500 1592.080 ;
        RECT 2705.265 1591.425 2707.855 1592.515 ;
        RECT 2706.645 1590.905 2707.855 1591.425 ;
        RECT 2708.485 1591.350 2708.775 1592.515 ;
        RECT 2708.945 1592.080 2714.290 1592.515 ;
        RECT 2714.465 1592.080 2719.810 1592.515 ;
        RECT 2712.350 1590.830 2712.700 1592.080 ;
        RECT 2717.870 1590.830 2718.220 1592.080 ;
        RECT 2719.985 1591.425 2721.195 1592.515 ;
        RECT 2720.675 1590.885 2721.195 1591.425 ;
        RECT 2721.365 1591.350 2721.655 1592.515 ;
        RECT 2721.825 1592.080 2727.170 1592.515 ;
        RECT 2727.345 1592.080 2732.690 1592.515 ;
        RECT 2725.230 1590.830 2725.580 1592.080 ;
        RECT 2730.750 1590.830 2731.100 1592.080 ;
        RECT 2732.865 1591.425 2734.075 1592.515 ;
        RECT 2732.865 1590.885 2733.385 1591.425 ;
        RECT 2522.135 1590.570 2523.935 1590.740 ;
        RECT 2522.830 1589.845 2523.160 1590.570 ;
        RECT 2522.135 1583.040 2523.935 1583.210 ;
        RECT 2522.830 1582.315 2523.160 1583.040 ;
        RECT 2522.135 1577.060 2523.935 1577.230 ;
        RECT 2522.830 1576.335 2523.160 1577.060 ;
        RECT 2522.135 1568.645 2523.935 1568.815 ;
        RECT 2522.830 1567.920 2523.160 1568.645 ;
        RECT 2360.030 1533.045 2360.205 1533.595 ;
        RECT 2360.030 1531.445 2360.200 1533.045 ;
        RECT 2358.215 1530.035 2358.385 1530.765 ;
        RECT 2360.030 1530.305 2360.205 1531.445 ;
        RECT 2360.030 1530.035 2360.200 1530.305 ;
        RECT 2366.795 1530.035 2366.965 1530.765 ;
        RECT 2372.410 1530.035 2372.580 1530.765 ;
        RECT 2375.155 1530.035 2375.325 1530.765 ;
        RECT 2376.150 1530.035 2376.320 1530.760 ;
        RECT 2383.120 1530.035 2383.290 1530.765 ;
        RECT 2388.735 1530.035 2388.905 1530.765 ;
        RECT 2391.480 1530.035 2391.650 1530.765 ;
        RECT 2392.475 1530.035 2392.645 1530.760 ;
        RECT 2399.445 1530.035 2399.615 1530.765 ;
        RECT 2405.060 1530.035 2405.230 1530.765 ;
        RECT 2407.805 1530.035 2407.975 1530.765 ;
        RECT 2408.800 1530.035 2408.970 1530.760 ;
        RECT 2415.770 1530.035 2415.940 1530.765 ;
        RECT 2421.385 1530.035 2421.555 1530.765 ;
        RECT 2424.130 1530.035 2424.300 1530.765 ;
        RECT 2425.125 1530.035 2425.295 1530.760 ;
        RECT 2432.095 1530.035 2432.265 1530.765 ;
        RECT 2437.710 1530.035 2437.880 1530.765 ;
        RECT 2440.455 1530.035 2440.625 1530.765 ;
        RECT 2441.450 1530.035 2441.620 1530.760 ;
        RECT 2343.000 1528.435 2442.420 1530.035 ;
        RECT 2360.790 1528.430 2442.420 1528.435 ;
        RECT 2361.535 1528.315 2371.195 1528.430 ;
        RECT 2372.240 1528.425 2375.975 1528.430 ;
        RECT 2362.825 1527.815 2362.995 1528.315 ;
        RECT 2365.265 1527.815 2365.435 1528.315 ;
        RECT 2366.225 1527.815 2366.395 1528.315 ;
        RECT 2367.225 1527.815 2367.395 1528.315 ;
        RECT 2369.665 1527.815 2369.835 1528.315 ;
        RECT 2370.625 1527.815 2370.795 1528.315 ;
        RECT 2372.410 1527.695 2372.580 1528.425 ;
        RECT 2375.155 1527.695 2375.325 1528.425 ;
        RECT 2376.145 1527.700 2376.315 1528.430 ;
        RECT 2377.860 1528.315 2387.520 1528.430 ;
        RECT 2388.565 1528.425 2392.300 1528.430 ;
        RECT 2379.150 1527.815 2379.320 1528.315 ;
        RECT 2381.590 1527.815 2381.760 1528.315 ;
        RECT 2382.550 1527.815 2382.720 1528.315 ;
        RECT 2383.550 1527.815 2383.720 1528.315 ;
        RECT 2385.990 1527.815 2386.160 1528.315 ;
        RECT 2386.950 1527.815 2387.120 1528.315 ;
        RECT 2388.735 1527.695 2388.905 1528.425 ;
        RECT 2391.480 1527.695 2391.650 1528.425 ;
        RECT 2392.470 1527.700 2392.640 1528.430 ;
        RECT 2394.185 1528.315 2403.845 1528.430 ;
        RECT 2404.890 1528.425 2408.625 1528.430 ;
        RECT 2395.475 1527.815 2395.645 1528.315 ;
        RECT 2397.915 1527.815 2398.085 1528.315 ;
        RECT 2398.875 1527.815 2399.045 1528.315 ;
        RECT 2399.875 1527.815 2400.045 1528.315 ;
        RECT 2402.315 1527.815 2402.485 1528.315 ;
        RECT 2403.275 1527.815 2403.445 1528.315 ;
        RECT 2405.060 1527.695 2405.230 1528.425 ;
        RECT 2407.805 1527.695 2407.975 1528.425 ;
        RECT 2408.795 1527.700 2408.965 1528.430 ;
        RECT 2410.510 1528.315 2420.170 1528.430 ;
        RECT 2421.215 1528.425 2424.950 1528.430 ;
        RECT 2411.800 1527.815 2411.970 1528.315 ;
        RECT 2414.240 1527.815 2414.410 1528.315 ;
        RECT 2415.200 1527.815 2415.370 1528.315 ;
        RECT 2416.200 1527.815 2416.370 1528.315 ;
        RECT 2418.640 1527.815 2418.810 1528.315 ;
        RECT 2419.600 1527.815 2419.770 1528.315 ;
        RECT 2421.385 1527.695 2421.555 1528.425 ;
        RECT 2424.130 1527.695 2424.300 1528.425 ;
        RECT 2425.120 1527.700 2425.290 1528.430 ;
        RECT 2426.835 1528.315 2436.495 1528.430 ;
        RECT 2437.540 1528.425 2441.275 1528.430 ;
        RECT 2428.125 1527.815 2428.295 1528.315 ;
        RECT 2430.565 1527.815 2430.735 1528.315 ;
        RECT 2431.525 1527.815 2431.695 1528.315 ;
        RECT 2432.525 1527.815 2432.695 1528.315 ;
        RECT 2434.965 1527.815 2435.135 1528.315 ;
        RECT 2435.925 1527.815 2436.095 1528.315 ;
        RECT 2437.710 1527.695 2437.880 1528.425 ;
        RECT 2440.455 1527.695 2440.625 1528.425 ;
        RECT 2441.445 1527.700 2441.615 1528.430 ;
        RECT 2696.295 1495.375 2696.815 1495.915 ;
        RECT 2695.605 1494.285 2696.815 1495.375 ;
        RECT 2697.425 1494.285 2697.755 1495.065 ;
        RECT 2698.315 1494.285 2698.650 1494.710 ;
        RECT 2699.265 1494.285 2699.595 1495.045 ;
        RECT 2700.645 1494.285 2700.975 1495.045 ;
        RECT 2704.990 1494.720 2705.340 1495.970 ;
        RECT 2707.795 1495.375 2708.315 1495.915 ;
        RECT 2701.585 1494.285 2706.930 1494.720 ;
        RECT 2707.105 1494.285 2708.315 1495.375 ;
        RECT 2708.485 1494.285 2708.775 1495.450 ;
        RECT 2709.420 1494.285 2709.750 1495.045 ;
        RECT 2710.350 1494.285 2710.610 1495.435 ;
        RECT 2714.190 1494.720 2714.540 1495.970 ;
        RECT 2718.125 1495.375 2719.815 1495.895 ;
        RECT 2720.675 1495.375 2721.195 1495.915 ;
        RECT 2710.785 1494.285 2716.130 1494.720 ;
        RECT 2716.305 1494.285 2719.815 1495.375 ;
        RECT 2719.985 1494.285 2721.195 1495.375 ;
        RECT 2721.365 1494.285 2721.655 1495.450 ;
        RECT 2721.830 1494.285 2722.165 1494.710 ;
        RECT 2722.725 1494.285 2723.055 1495.065 ;
        RECT 2727.070 1494.720 2727.420 1495.970 ;
        RECT 2730.105 1495.375 2730.855 1495.895 ;
        RECT 2723.665 1494.285 2729.010 1494.720 ;
        RECT 2729.185 1494.285 2730.855 1495.375 ;
        RECT 2732.865 1495.375 2733.385 1495.915 ;
        RECT 2731.925 1494.285 2732.255 1495.045 ;
        RECT 2732.865 1494.285 2734.075 1495.375 ;
        RECT 2695.520 1494.115 2734.160 1494.285 ;
        RECT 2695.605 1493.025 2696.815 1494.115 ;
        RECT 2697.425 1493.355 2697.755 1494.115 ;
        RECT 2698.365 1493.680 2703.710 1494.115 ;
        RECT 2696.295 1492.485 2696.815 1493.025 ;
        RECT 2701.770 1492.430 2702.120 1493.680 ;
        RECT 2703.885 1493.025 2707.395 1494.115 ;
        RECT 2705.705 1492.505 2707.395 1493.025 ;
        RECT 2708.485 1492.950 2708.775 1494.115 ;
        RECT 2708.945 1493.680 2714.290 1494.115 ;
        RECT 2714.465 1493.680 2719.810 1494.115 ;
        RECT 2719.985 1493.680 2725.330 1494.115 ;
        RECT 2725.505 1493.680 2730.850 1494.115 ;
        RECT 2712.350 1492.430 2712.700 1493.680 ;
        RECT 2717.870 1492.430 2718.220 1493.680 ;
        RECT 2723.390 1492.430 2723.740 1493.680 ;
        RECT 2728.910 1492.430 2729.260 1493.680 ;
        RECT 2731.025 1493.025 2732.695 1494.115 ;
        RECT 2731.945 1492.505 2732.695 1493.025 ;
        RECT 2732.865 1493.025 2734.075 1494.115 ;
        RECT 2732.865 1492.485 2733.385 1493.025 ;
        RECT 2696.295 1489.935 2696.815 1490.475 ;
        RECT 2695.605 1488.845 2696.815 1489.935 ;
        RECT 2700.390 1489.280 2700.740 1490.530 ;
        RECT 2705.910 1489.280 2706.260 1490.530 ;
        RECT 2711.430 1489.280 2711.780 1490.530 ;
        RECT 2716.950 1489.280 2717.300 1490.530 ;
        RECT 2719.985 1489.935 2720.735 1490.455 ;
        RECT 2696.985 1488.845 2702.330 1489.280 ;
        RECT 2702.505 1488.845 2707.850 1489.280 ;
        RECT 2708.025 1488.845 2713.370 1489.280 ;
        RECT 2713.545 1488.845 2718.890 1489.280 ;
        RECT 2719.065 1488.845 2720.735 1489.935 ;
        RECT 2721.365 1488.845 2721.655 1490.010 ;
        RECT 2725.230 1489.280 2725.580 1490.530 ;
        RECT 2730.750 1489.280 2731.100 1490.530 ;
        RECT 2732.865 1489.935 2733.385 1490.475 ;
        RECT 2721.825 1488.845 2727.170 1489.280 ;
        RECT 2727.345 1488.845 2732.690 1489.280 ;
        RECT 2732.865 1488.845 2734.075 1489.935 ;
        RECT 2695.520 1488.675 2734.160 1488.845 ;
        RECT 2695.605 1487.585 2696.815 1488.675 ;
        RECT 2696.985 1488.240 2702.330 1488.675 ;
        RECT 2702.505 1488.240 2707.850 1488.675 ;
        RECT 2696.295 1487.045 2696.815 1487.585 ;
        RECT 2700.390 1486.990 2700.740 1488.240 ;
        RECT 2705.910 1486.990 2706.260 1488.240 ;
        RECT 2708.485 1487.510 2708.775 1488.675 ;
        RECT 2708.945 1488.240 2714.290 1488.675 ;
        RECT 2714.465 1488.240 2719.810 1488.675 ;
        RECT 2719.985 1488.240 2725.330 1488.675 ;
        RECT 2725.505 1488.240 2730.850 1488.675 ;
        RECT 2712.350 1486.990 2712.700 1488.240 ;
        RECT 2717.870 1486.990 2718.220 1488.240 ;
        RECT 2723.390 1486.990 2723.740 1488.240 ;
        RECT 2728.910 1486.990 2729.260 1488.240 ;
        RECT 2731.025 1487.585 2732.695 1488.675 ;
        RECT 2731.945 1487.065 2732.695 1487.585 ;
        RECT 2732.865 1487.585 2734.075 1488.675 ;
        RECT 2732.865 1487.045 2733.385 1487.585 ;
        RECT 2696.295 1484.495 2696.815 1485.035 ;
        RECT 2695.605 1483.405 2696.815 1484.495 ;
        RECT 2697.425 1483.405 2697.755 1484.165 ;
        RECT 2701.770 1483.840 2702.120 1485.090 ;
        RECT 2707.290 1483.840 2707.640 1485.090 ;
        RECT 2712.810 1483.840 2713.160 1485.090 ;
        RECT 2718.330 1483.840 2718.680 1485.090 ;
        RECT 2698.365 1483.405 2703.710 1483.840 ;
        RECT 2703.885 1483.405 2709.230 1483.840 ;
        RECT 2709.405 1483.405 2714.750 1483.840 ;
        RECT 2714.925 1483.405 2720.270 1483.840 ;
        RECT 2721.365 1483.405 2721.655 1484.570 ;
        RECT 2725.230 1483.840 2725.580 1485.090 ;
        RECT 2730.750 1483.840 2731.100 1485.090 ;
        RECT 2732.865 1484.495 2733.385 1485.035 ;
        RECT 2721.825 1483.405 2727.170 1483.840 ;
        RECT 2727.345 1483.405 2732.690 1483.840 ;
        RECT 2732.865 1483.405 2734.075 1484.495 ;
        RECT 2695.520 1483.235 2734.160 1483.405 ;
        RECT 2695.605 1482.145 2696.815 1483.235 ;
        RECT 2696.985 1482.800 2702.330 1483.235 ;
        RECT 2702.505 1482.800 2707.850 1483.235 ;
        RECT 2696.295 1481.605 2696.815 1482.145 ;
        RECT 2700.390 1481.550 2700.740 1482.800 ;
        RECT 2705.910 1481.550 2706.260 1482.800 ;
        RECT 2708.485 1482.070 2708.775 1483.235 ;
        RECT 2708.945 1482.800 2714.290 1483.235 ;
        RECT 2714.465 1482.800 2719.810 1483.235 ;
        RECT 2719.985 1482.800 2725.330 1483.235 ;
        RECT 2725.505 1482.800 2730.850 1483.235 ;
        RECT 2712.350 1481.550 2712.700 1482.800 ;
        RECT 2717.870 1481.550 2718.220 1482.800 ;
        RECT 2723.390 1481.550 2723.740 1482.800 ;
        RECT 2728.910 1481.550 2729.260 1482.800 ;
        RECT 2731.025 1482.145 2732.695 1483.235 ;
        RECT 2731.945 1481.625 2732.695 1482.145 ;
        RECT 2732.865 1482.145 2734.075 1483.235 ;
        RECT 2732.865 1481.605 2733.385 1482.145 ;
        RECT 2696.295 1479.055 2696.815 1479.595 ;
        RECT 2695.605 1477.965 2696.815 1479.055 ;
        RECT 2710.050 1478.400 2710.400 1479.650 ;
        RECT 2715.570 1478.400 2715.920 1479.650 ;
        RECT 2719.505 1479.055 2721.195 1479.575 ;
        RECT 2697.415 1477.965 2697.745 1478.345 ;
        RECT 2700.135 1477.965 2700.465 1478.345 ;
        RECT 2701.960 1477.965 2702.290 1478.345 ;
        RECT 2702.880 1477.965 2703.230 1478.345 ;
        RECT 2705.715 1477.965 2706.045 1478.345 ;
        RECT 2706.645 1477.965 2711.990 1478.400 ;
        RECT 2712.165 1477.965 2717.510 1478.400 ;
        RECT 2717.685 1477.965 2721.195 1479.055 ;
        RECT 2721.365 1477.965 2721.655 1479.130 ;
        RECT 2725.230 1478.400 2725.580 1479.650 ;
        RECT 2730.750 1478.400 2731.100 1479.650 ;
        RECT 2732.865 1479.055 2733.385 1479.595 ;
        RECT 2721.825 1477.965 2727.170 1478.400 ;
        RECT 2727.345 1477.965 2732.690 1478.400 ;
        RECT 2732.865 1477.965 2734.075 1479.055 ;
        RECT 2695.520 1477.795 2734.160 1477.965 ;
        RECT 2695.605 1476.705 2696.815 1477.795 ;
        RECT 2697.425 1477.035 2697.755 1477.795 ;
        RECT 2698.365 1477.360 2703.710 1477.795 ;
        RECT 2696.295 1476.165 2696.815 1476.705 ;
        RECT 2701.770 1476.110 2702.120 1477.360 ;
        RECT 2703.885 1476.705 2707.395 1477.795 ;
        RECT 2705.705 1476.185 2707.395 1476.705 ;
        RECT 2708.485 1476.630 2708.775 1477.795 ;
        RECT 2708.945 1477.360 2714.290 1477.795 ;
        RECT 2714.465 1477.360 2719.810 1477.795 ;
        RECT 2719.985 1477.360 2725.330 1477.795 ;
        RECT 2725.505 1477.360 2730.850 1477.795 ;
        RECT 2712.350 1476.110 2712.700 1477.360 ;
        RECT 2717.870 1476.110 2718.220 1477.360 ;
        RECT 2723.390 1476.110 2723.740 1477.360 ;
        RECT 2728.910 1476.110 2729.260 1477.360 ;
        RECT 2731.025 1476.705 2732.695 1477.795 ;
        RECT 2731.945 1476.185 2732.695 1476.705 ;
        RECT 2732.865 1476.705 2734.075 1477.795 ;
        RECT 2732.865 1476.165 2733.385 1476.705 ;
        RECT 2696.295 1473.615 2696.815 1474.155 ;
        RECT 2695.605 1472.525 2696.815 1473.615 ;
        RECT 2710.050 1472.960 2710.400 1474.210 ;
        RECT 2715.570 1472.960 2715.920 1474.210 ;
        RECT 2719.505 1473.615 2721.195 1474.135 ;
        RECT 2697.415 1472.525 2697.745 1472.905 ;
        RECT 2700.135 1472.525 2700.465 1472.905 ;
        RECT 2701.960 1472.525 2702.290 1472.905 ;
        RECT 2702.880 1472.525 2703.230 1472.905 ;
        RECT 2705.715 1472.525 2706.045 1472.905 ;
        RECT 2706.645 1472.525 2711.990 1472.960 ;
        RECT 2712.165 1472.525 2717.510 1472.960 ;
        RECT 2717.685 1472.525 2721.195 1473.615 ;
        RECT 2721.365 1472.525 2721.655 1473.690 ;
        RECT 2725.230 1472.960 2725.580 1474.210 ;
        RECT 2730.750 1472.960 2731.100 1474.210 ;
        RECT 2732.865 1473.615 2733.385 1474.155 ;
        RECT 2721.825 1472.525 2727.170 1472.960 ;
        RECT 2727.345 1472.525 2732.690 1472.960 ;
        RECT 2732.865 1472.525 2734.075 1473.615 ;
        RECT 2695.520 1472.355 2734.160 1472.525 ;
        RECT 2695.605 1471.265 2696.815 1472.355 ;
        RECT 2697.425 1471.595 2697.755 1472.355 ;
        RECT 2698.365 1471.265 2700.955 1472.355 ;
        RECT 2696.295 1470.725 2696.815 1471.265 ;
        RECT 2699.745 1470.745 2700.955 1471.265 ;
        RECT 2702.095 1471.215 2702.265 1472.355 ;
        RECT 2704.635 1471.595 2704.805 1472.355 ;
        RECT 2705.725 1471.265 2708.315 1472.355 ;
        RECT 2707.105 1470.745 2708.315 1471.265 ;
        RECT 2708.485 1471.190 2708.775 1472.355 ;
        RECT 2708.945 1471.920 2714.290 1472.355 ;
        RECT 2714.465 1471.920 2719.810 1472.355 ;
        RECT 2719.985 1471.920 2725.330 1472.355 ;
        RECT 2725.505 1471.920 2730.850 1472.355 ;
        RECT 2712.350 1470.670 2712.700 1471.920 ;
        RECT 2717.870 1470.670 2718.220 1471.920 ;
        RECT 2723.390 1470.670 2723.740 1471.920 ;
        RECT 2728.910 1470.670 2729.260 1471.920 ;
        RECT 2731.025 1471.265 2732.695 1472.355 ;
        RECT 2731.945 1470.745 2732.695 1471.265 ;
        RECT 2732.865 1471.265 2734.075 1472.355 ;
        RECT 2732.865 1470.725 2733.385 1471.265 ;
        RECT 2696.295 1468.175 2696.815 1468.715 ;
        RECT 2695.605 1467.085 2696.815 1468.175 ;
        RECT 2700.390 1467.520 2700.740 1468.770 ;
        RECT 2705.910 1467.520 2706.260 1468.770 ;
        RECT 2711.430 1467.520 2711.780 1468.770 ;
        RECT 2716.950 1467.520 2717.300 1468.770 ;
        RECT 2719.985 1468.175 2720.735 1468.695 ;
        RECT 2696.985 1467.085 2702.330 1467.520 ;
        RECT 2702.505 1467.085 2707.850 1467.520 ;
        RECT 2708.025 1467.085 2713.370 1467.520 ;
        RECT 2713.545 1467.085 2718.890 1467.520 ;
        RECT 2719.065 1467.085 2720.735 1468.175 ;
        RECT 2721.365 1467.085 2721.655 1468.250 ;
        RECT 2725.230 1467.520 2725.580 1468.770 ;
        RECT 2730.750 1467.520 2731.100 1468.770 ;
        RECT 2732.865 1468.175 2733.385 1468.715 ;
        RECT 2721.825 1467.085 2727.170 1467.520 ;
        RECT 2727.345 1467.085 2732.690 1467.520 ;
        RECT 2732.865 1467.085 2734.075 1468.175 ;
        RECT 2695.520 1466.915 2734.160 1467.085 ;
        RECT 2695.605 1465.825 2696.815 1466.915 ;
        RECT 2697.425 1466.155 2697.755 1466.915 ;
        RECT 2698.365 1466.480 2703.710 1466.915 ;
        RECT 2696.295 1465.285 2696.815 1465.825 ;
        RECT 2701.770 1465.230 2702.120 1466.480 ;
        RECT 2703.885 1465.825 2707.395 1466.915 ;
        RECT 2705.705 1465.305 2707.395 1465.825 ;
        RECT 2708.485 1465.750 2708.775 1466.915 ;
        RECT 2708.945 1466.480 2714.290 1466.915 ;
        RECT 2714.465 1466.480 2719.810 1466.915 ;
        RECT 2719.985 1466.480 2725.330 1466.915 ;
        RECT 2725.505 1466.480 2730.850 1466.915 ;
        RECT 2712.350 1465.230 2712.700 1466.480 ;
        RECT 2717.870 1465.230 2718.220 1466.480 ;
        RECT 2723.390 1465.230 2723.740 1466.480 ;
        RECT 2728.910 1465.230 2729.260 1466.480 ;
        RECT 2731.025 1465.825 2732.695 1466.915 ;
        RECT 2731.945 1465.305 2732.695 1465.825 ;
        RECT 2732.865 1465.825 2734.075 1466.915 ;
        RECT 2732.865 1465.285 2733.385 1465.825 ;
        RECT 2696.295 1462.735 2696.815 1463.275 ;
        RECT 2695.605 1461.645 2696.815 1462.735 ;
        RECT 2700.390 1462.080 2700.740 1463.330 ;
        RECT 2705.910 1462.080 2706.260 1463.330 ;
        RECT 2711.430 1462.080 2711.780 1463.330 ;
        RECT 2716.950 1462.080 2717.300 1463.330 ;
        RECT 2719.985 1462.735 2720.735 1463.255 ;
        RECT 2696.985 1461.645 2702.330 1462.080 ;
        RECT 2702.505 1461.645 2707.850 1462.080 ;
        RECT 2708.025 1461.645 2713.370 1462.080 ;
        RECT 2713.545 1461.645 2718.890 1462.080 ;
        RECT 2719.065 1461.645 2720.735 1462.735 ;
        RECT 2721.365 1461.645 2721.655 1462.810 ;
        RECT 2725.230 1462.080 2725.580 1463.330 ;
        RECT 2730.750 1462.080 2731.100 1463.330 ;
        RECT 2732.865 1462.735 2733.385 1463.275 ;
        RECT 2721.825 1461.645 2727.170 1462.080 ;
        RECT 2727.345 1461.645 2732.690 1462.080 ;
        RECT 2732.865 1461.645 2734.075 1462.735 ;
        RECT 2695.520 1461.475 2734.160 1461.645 ;
        RECT 2695.605 1460.385 2696.815 1461.475 ;
        RECT 2696.985 1460.385 2700.495 1461.475 ;
        RECT 2696.295 1459.845 2696.815 1460.385 ;
        RECT 2698.805 1459.865 2700.495 1460.385 ;
        RECT 2702.455 1460.335 2702.785 1461.475 ;
        RECT 2702.965 1461.040 2708.310 1461.475 ;
        RECT 2706.370 1459.790 2706.720 1461.040 ;
        RECT 2708.485 1460.310 2708.775 1461.475 ;
        RECT 2708.945 1461.040 2714.290 1461.475 ;
        RECT 2714.465 1461.040 2719.810 1461.475 ;
        RECT 2719.985 1461.040 2725.330 1461.475 ;
        RECT 2725.505 1461.040 2730.850 1461.475 ;
        RECT 2712.350 1459.790 2712.700 1461.040 ;
        RECT 2717.870 1459.790 2718.220 1461.040 ;
        RECT 2723.390 1459.790 2723.740 1461.040 ;
        RECT 2728.910 1459.790 2729.260 1461.040 ;
        RECT 2731.025 1460.385 2732.695 1461.475 ;
        RECT 2731.945 1459.865 2732.695 1460.385 ;
        RECT 2732.865 1460.385 2734.075 1461.475 ;
        RECT 2732.865 1459.845 2733.385 1460.385 ;
        RECT 2696.295 1457.295 2696.815 1457.835 ;
        RECT 2700.185 1457.295 2701.875 1457.815 ;
        RECT 2695.605 1456.205 2696.815 1457.295 ;
        RECT 2697.425 1456.205 2697.755 1456.965 ;
        RECT 2698.365 1456.205 2701.875 1457.295 ;
        RECT 2703.535 1456.205 2703.705 1456.645 ;
        RECT 2708.670 1456.640 2709.020 1457.890 ;
        RECT 2714.190 1456.640 2714.540 1457.890 ;
        RECT 2718.125 1457.295 2719.815 1457.815 ;
        RECT 2720.675 1457.295 2721.195 1457.835 ;
        RECT 2704.310 1456.205 2704.640 1456.565 ;
        RECT 2705.265 1456.205 2710.610 1456.640 ;
        RECT 2710.785 1456.205 2716.130 1456.640 ;
        RECT 2716.305 1456.205 2719.815 1457.295 ;
        RECT 2719.985 1456.205 2721.195 1457.295 ;
        RECT 2721.365 1456.205 2721.655 1457.370 ;
        RECT 2725.230 1456.640 2725.580 1457.890 ;
        RECT 2730.750 1456.640 2731.100 1457.890 ;
        RECT 2732.865 1457.295 2733.385 1457.835 ;
        RECT 2721.825 1456.205 2727.170 1456.640 ;
        RECT 2727.345 1456.205 2732.690 1456.640 ;
        RECT 2732.865 1456.205 2734.075 1457.295 ;
        RECT 2695.520 1456.035 2734.160 1456.205 ;
        RECT 2695.605 1454.945 2696.815 1456.035 ;
        RECT 2696.985 1455.600 2702.330 1456.035 ;
        RECT 2702.505 1455.600 2707.850 1456.035 ;
        RECT 2696.295 1454.405 2696.815 1454.945 ;
        RECT 2700.390 1454.350 2700.740 1455.600 ;
        RECT 2705.910 1454.350 2706.260 1455.600 ;
        RECT 2708.485 1454.870 2708.775 1456.035 ;
        RECT 2708.945 1455.600 2714.290 1456.035 ;
        RECT 2714.465 1455.600 2719.810 1456.035 ;
        RECT 2719.985 1455.600 2725.330 1456.035 ;
        RECT 2712.350 1454.350 2712.700 1455.600 ;
        RECT 2717.870 1454.350 2718.220 1455.600 ;
        RECT 2723.390 1454.350 2723.740 1455.600 ;
        RECT 2725.595 1455.235 2725.765 1456.035 ;
        RECT 2726.435 1455.235 2726.605 1456.035 ;
        RECT 2727.275 1455.235 2727.445 1456.035 ;
        RECT 2728.035 1455.235 2728.365 1456.035 ;
        RECT 2728.875 1455.235 2729.205 1456.035 ;
        RECT 2729.715 1455.235 2730.045 1456.035 ;
        RECT 2730.555 1455.235 2730.885 1456.035 ;
        RECT 2731.395 1455.235 2731.725 1456.035 ;
        RECT 2732.235 1454.885 2732.565 1456.035 ;
        RECT 2732.865 1454.945 2734.075 1456.035 ;
        RECT 2732.865 1454.405 2733.385 1454.945 ;
        RECT 2696.295 1451.855 2696.815 1452.395 ;
        RECT 2695.605 1450.765 2696.815 1451.855 ;
        RECT 2697.425 1450.765 2697.755 1451.525 ;
        RECT 2701.770 1451.200 2702.120 1452.450 ;
        RECT 2707.290 1451.200 2707.640 1452.450 ;
        RECT 2712.810 1451.200 2713.160 1452.450 ;
        RECT 2718.330 1451.200 2718.680 1452.450 ;
        RECT 2698.365 1450.765 2703.710 1451.200 ;
        RECT 2703.885 1450.765 2709.230 1451.200 ;
        RECT 2709.405 1450.765 2714.750 1451.200 ;
        RECT 2714.925 1450.765 2720.270 1451.200 ;
        RECT 2721.365 1450.765 2721.655 1451.930 ;
        RECT 2725.230 1451.200 2725.580 1452.450 ;
        RECT 2730.750 1451.200 2731.100 1452.450 ;
        RECT 2732.865 1451.855 2733.385 1452.395 ;
        RECT 2721.825 1450.765 2727.170 1451.200 ;
        RECT 2727.345 1450.765 2732.690 1451.200 ;
        RECT 2732.865 1450.765 2734.075 1451.855 ;
        RECT 2695.520 1450.595 2734.160 1450.765 ;
        RECT 2695.605 1449.505 2696.815 1450.595 ;
        RECT 2696.985 1450.160 2702.330 1450.595 ;
        RECT 2702.505 1450.160 2707.850 1450.595 ;
        RECT 2696.295 1448.965 2696.815 1449.505 ;
        RECT 2700.390 1448.910 2700.740 1450.160 ;
        RECT 2705.910 1448.910 2706.260 1450.160 ;
        RECT 2708.485 1449.430 2708.775 1450.595 ;
        RECT 2708.945 1450.160 2714.290 1450.595 ;
        RECT 2714.465 1450.160 2719.810 1450.595 ;
        RECT 2719.985 1450.160 2725.330 1450.595 ;
        RECT 2725.505 1450.160 2730.850 1450.595 ;
        RECT 2712.350 1448.910 2712.700 1450.160 ;
        RECT 2717.870 1448.910 2718.220 1450.160 ;
        RECT 2723.390 1448.910 2723.740 1450.160 ;
        RECT 2728.910 1448.910 2729.260 1450.160 ;
        RECT 2731.025 1449.505 2732.695 1450.595 ;
        RECT 2731.945 1448.985 2732.695 1449.505 ;
        RECT 2732.865 1449.505 2734.075 1450.595 ;
        RECT 2732.865 1448.965 2733.385 1449.505 ;
        RECT 2696.295 1446.415 2696.815 1446.955 ;
        RECT 2695.605 1445.325 2696.815 1446.415 ;
        RECT 2697.715 1445.325 2698.045 1445.835 ;
        RECT 2703.150 1445.760 2703.500 1447.010 ;
        RECT 2708.670 1445.760 2709.020 1447.010 ;
        RECT 2714.190 1445.760 2714.540 1447.010 ;
        RECT 2718.125 1446.415 2719.815 1446.935 ;
        RECT 2720.675 1446.415 2721.195 1446.955 ;
        RECT 2699.745 1445.325 2705.090 1445.760 ;
        RECT 2705.265 1445.325 2710.610 1445.760 ;
        RECT 2710.785 1445.325 2716.130 1445.760 ;
        RECT 2716.305 1445.325 2719.815 1446.415 ;
        RECT 2719.985 1445.325 2721.195 1446.415 ;
        RECT 2721.365 1445.325 2721.655 1446.490 ;
        RECT 2725.230 1445.760 2725.580 1447.010 ;
        RECT 2730.750 1445.760 2731.100 1447.010 ;
        RECT 2732.865 1446.415 2733.385 1446.955 ;
        RECT 2721.825 1445.325 2727.170 1445.760 ;
        RECT 2727.345 1445.325 2732.690 1445.760 ;
        RECT 2732.865 1445.325 2734.075 1446.415 ;
        RECT 2695.520 1445.155 2734.160 1445.325 ;
        RECT 2695.605 1444.065 2696.815 1445.155 ;
        RECT 2697.425 1444.395 2697.755 1445.155 ;
        RECT 2698.365 1444.720 2703.710 1445.155 ;
        RECT 2696.295 1443.525 2696.815 1444.065 ;
        RECT 2701.770 1443.470 2702.120 1444.720 ;
        RECT 2703.885 1444.065 2707.395 1445.155 ;
        RECT 2705.705 1443.545 2707.395 1444.065 ;
        RECT 2708.485 1443.990 2708.775 1445.155 ;
        RECT 2708.945 1444.720 2714.290 1445.155 ;
        RECT 2714.465 1444.720 2719.810 1445.155 ;
        RECT 2719.985 1444.720 2725.330 1445.155 ;
        RECT 2725.505 1444.720 2730.850 1445.155 ;
        RECT 2712.350 1443.470 2712.700 1444.720 ;
        RECT 2717.870 1443.470 2718.220 1444.720 ;
        RECT 2723.390 1443.470 2723.740 1444.720 ;
        RECT 2728.910 1443.470 2729.260 1444.720 ;
        RECT 2731.025 1444.065 2732.695 1445.155 ;
        RECT 2731.945 1443.545 2732.695 1444.065 ;
        RECT 2732.865 1444.065 2734.075 1445.155 ;
        RECT 2732.865 1443.525 2733.385 1444.065 ;
        RECT 2696.295 1440.975 2696.815 1441.515 ;
        RECT 2695.605 1439.885 2696.815 1440.975 ;
        RECT 2697.735 1439.885 2697.905 1440.645 ;
        RECT 2700.275 1439.885 2700.445 1441.025 ;
        RECT 2701.590 1439.885 2701.920 1440.600 ;
        RECT 2708.210 1440.320 2708.560 1441.570 ;
        RECT 2713.730 1440.320 2714.080 1441.570 ;
        RECT 2719.250 1440.320 2719.600 1441.570 ;
        RECT 2704.805 1439.885 2710.150 1440.320 ;
        RECT 2710.325 1439.885 2715.670 1440.320 ;
        RECT 2715.845 1439.885 2721.190 1440.320 ;
        RECT 2721.365 1439.885 2721.655 1441.050 ;
        RECT 2725.230 1440.320 2725.580 1441.570 ;
        RECT 2730.750 1440.320 2731.100 1441.570 ;
        RECT 2732.865 1440.975 2733.385 1441.515 ;
        RECT 2721.825 1439.885 2727.170 1440.320 ;
        RECT 2727.345 1439.885 2732.690 1440.320 ;
        RECT 2732.865 1439.885 2734.075 1440.975 ;
        RECT 2695.520 1439.715 2734.160 1439.885 ;
        RECT 2522.135 1438.945 2523.935 1439.115 ;
        RECT 2522.830 1438.220 2523.160 1438.945 ;
        RECT 2695.605 1438.625 2696.815 1439.715 ;
        RECT 2696.985 1439.205 2697.245 1439.715 ;
        RECT 2697.905 1439.210 2698.520 1439.715 ;
        RECT 2698.325 1439.035 2698.520 1439.210 ;
        RECT 2699.335 1439.170 2699.550 1439.715 ;
        RECT 2700.205 1439.280 2705.550 1439.715 ;
        RECT 2698.325 1438.845 2698.655 1439.035 ;
        RECT 2696.295 1438.085 2696.815 1438.625 ;
        RECT 2703.610 1438.030 2703.960 1439.280 ;
        RECT 2705.725 1438.625 2708.315 1439.715 ;
        RECT 2707.105 1438.105 2708.315 1438.625 ;
        RECT 2708.485 1438.550 2708.775 1439.715 ;
        RECT 2708.945 1439.280 2714.290 1439.715 ;
        RECT 2714.465 1439.280 2719.810 1439.715 ;
        RECT 2719.985 1439.280 2725.330 1439.715 ;
        RECT 2725.505 1439.280 2730.850 1439.715 ;
        RECT 2712.350 1438.030 2712.700 1439.280 ;
        RECT 2717.870 1438.030 2718.220 1439.280 ;
        RECT 2723.390 1438.030 2723.740 1439.280 ;
        RECT 2728.910 1438.030 2729.260 1439.280 ;
        RECT 2731.025 1438.625 2732.695 1439.715 ;
        RECT 2731.945 1438.105 2732.695 1438.625 ;
        RECT 2732.865 1438.625 2734.075 1439.715 ;
        RECT 2732.865 1438.085 2733.385 1438.625 ;
        RECT 2360.030 1435.050 2360.205 1435.600 ;
        RECT 2696.295 1435.535 2696.815 1436.075 ;
        RECT 2360.030 1433.450 2360.200 1435.050 ;
        RECT 2695.605 1434.445 2696.815 1435.535 ;
        RECT 2697.425 1434.445 2697.755 1435.205 ;
        RECT 2701.770 1434.880 2702.120 1436.130 ;
        RECT 2707.290 1434.880 2707.640 1436.130 ;
        RECT 2712.810 1434.880 2713.160 1436.130 ;
        RECT 2718.330 1434.880 2718.680 1436.130 ;
        RECT 2698.365 1434.445 2703.710 1434.880 ;
        RECT 2703.885 1434.445 2709.230 1434.880 ;
        RECT 2709.405 1434.445 2714.750 1434.880 ;
        RECT 2714.925 1434.445 2720.270 1434.880 ;
        RECT 2721.365 1434.445 2721.655 1435.610 ;
        RECT 2725.230 1434.880 2725.580 1436.130 ;
        RECT 2730.750 1434.880 2731.100 1436.130 ;
        RECT 2732.865 1435.535 2733.385 1436.075 ;
        RECT 2721.825 1434.445 2727.170 1434.880 ;
        RECT 2727.345 1434.445 2732.690 1434.880 ;
        RECT 2732.865 1434.445 2734.075 1435.535 ;
        RECT 2695.520 1434.275 2734.160 1434.445 ;
        RECT 2358.215 1432.040 2358.385 1432.770 ;
        RECT 2360.030 1432.310 2360.205 1433.450 ;
        RECT 2695.605 1433.185 2696.815 1434.275 ;
        RECT 2696.985 1433.185 2698.195 1434.275 ;
        RECT 2698.865 1433.815 2699.115 1434.275 ;
        RECT 2699.795 1433.815 2700.045 1434.275 ;
        RECT 2701.115 1433.815 2701.365 1434.275 ;
        RECT 2702.045 1433.840 2707.390 1434.275 ;
        RECT 2360.030 1432.040 2360.200 1432.310 ;
        RECT 2369.030 1432.040 2369.200 1432.770 ;
        RECT 2374.645 1432.040 2374.815 1432.770 ;
        RECT 2377.390 1432.040 2377.560 1432.770 ;
        RECT 2378.385 1432.040 2378.555 1432.765 ;
        RECT 2387.590 1432.040 2387.760 1432.770 ;
        RECT 2393.205 1432.040 2393.375 1432.770 ;
        RECT 2395.950 1432.040 2396.120 1432.770 ;
        RECT 2396.945 1432.040 2397.115 1432.765 ;
        RECT 2406.150 1432.040 2406.320 1432.770 ;
        RECT 2411.765 1432.040 2411.935 1432.770 ;
        RECT 2414.510 1432.040 2414.680 1432.770 ;
        RECT 2415.505 1432.040 2415.675 1432.765 ;
        RECT 2424.710 1432.040 2424.880 1432.770 ;
        RECT 2430.325 1432.040 2430.495 1432.770 ;
        RECT 2433.070 1432.040 2433.240 1432.770 ;
        RECT 2434.065 1432.040 2434.235 1432.765 ;
        RECT 2443.270 1432.040 2443.440 1432.770 ;
        RECT 2448.885 1432.040 2449.055 1432.770 ;
        RECT 2451.630 1432.040 2451.800 1432.770 ;
        RECT 2452.625 1432.040 2452.795 1432.765 ;
        RECT 2522.135 1432.530 2523.935 1432.700 ;
        RECT 2696.295 1432.645 2696.815 1433.185 ;
        RECT 2697.675 1432.645 2698.195 1433.185 ;
        RECT 2705.450 1432.590 2705.800 1433.840 ;
        RECT 2708.485 1433.110 2708.775 1434.275 ;
        RECT 2708.945 1433.840 2714.290 1434.275 ;
        RECT 2714.465 1433.840 2719.810 1434.275 ;
        RECT 2719.985 1433.840 2725.330 1434.275 ;
        RECT 2725.505 1433.840 2730.850 1434.275 ;
        RECT 2712.350 1432.590 2712.700 1433.840 ;
        RECT 2717.870 1432.590 2718.220 1433.840 ;
        RECT 2723.390 1432.590 2723.740 1433.840 ;
        RECT 2728.910 1432.590 2729.260 1433.840 ;
        RECT 2731.025 1433.185 2732.695 1434.275 ;
        RECT 2731.945 1432.665 2732.695 1433.185 ;
        RECT 2732.865 1433.185 2734.075 1434.275 ;
        RECT 2732.865 1432.645 2733.385 1433.185 ;
        RECT 2343.000 1432.035 2453.495 1432.040 ;
        RECT 2343.000 1430.440 2453.595 1432.035 ;
        RECT 2522.830 1431.805 2523.160 1432.530 ;
        RECT 2361.540 1430.430 2379.355 1430.440 ;
        RECT 2380.100 1430.430 2397.915 1430.440 ;
        RECT 2398.660 1430.430 2416.475 1430.440 ;
        RECT 2417.220 1430.430 2435.035 1430.440 ;
        RECT 2435.780 1430.430 2453.595 1430.440 ;
        RECT 2361.540 1430.425 2373.500 1430.430 ;
        RECT 2374.475 1430.425 2378.210 1430.430 ;
        RECT 2362.350 1429.925 2362.520 1430.425 ;
        RECT 2363.310 1429.925 2363.480 1430.425 ;
        RECT 2364.310 1429.925 2364.480 1430.425 ;
        RECT 2366.270 1429.925 2366.440 1430.425 ;
        RECT 2367.230 1429.925 2367.400 1430.425 ;
        RECT 2369.190 1429.925 2369.360 1430.425 ;
        RECT 2371.630 1429.925 2371.800 1430.425 ;
        RECT 2374.645 1429.695 2374.815 1430.425 ;
        RECT 2377.390 1429.695 2377.560 1430.425 ;
        RECT 2378.380 1429.700 2378.550 1430.430 ;
        RECT 2380.100 1430.425 2392.060 1430.430 ;
        RECT 2393.035 1430.425 2396.770 1430.430 ;
        RECT 2380.910 1429.925 2381.080 1430.425 ;
        RECT 2381.870 1429.925 2382.040 1430.425 ;
        RECT 2382.870 1429.925 2383.040 1430.425 ;
        RECT 2384.830 1429.925 2385.000 1430.425 ;
        RECT 2385.790 1429.925 2385.960 1430.425 ;
        RECT 2387.750 1429.925 2387.920 1430.425 ;
        RECT 2390.190 1429.925 2390.360 1430.425 ;
        RECT 2393.205 1429.695 2393.375 1430.425 ;
        RECT 2395.950 1429.695 2396.120 1430.425 ;
        RECT 2396.940 1429.700 2397.110 1430.430 ;
        RECT 2398.660 1430.425 2410.620 1430.430 ;
        RECT 2411.595 1430.425 2415.330 1430.430 ;
        RECT 2399.470 1429.925 2399.640 1430.425 ;
        RECT 2400.430 1429.925 2400.600 1430.425 ;
        RECT 2401.430 1429.925 2401.600 1430.425 ;
        RECT 2403.390 1429.925 2403.560 1430.425 ;
        RECT 2404.350 1429.925 2404.520 1430.425 ;
        RECT 2406.310 1429.925 2406.480 1430.425 ;
        RECT 2408.750 1429.925 2408.920 1430.425 ;
        RECT 2411.765 1429.695 2411.935 1430.425 ;
        RECT 2414.510 1429.695 2414.680 1430.425 ;
        RECT 2415.500 1429.700 2415.670 1430.430 ;
        RECT 2417.220 1430.425 2429.180 1430.430 ;
        RECT 2430.155 1430.425 2433.890 1430.430 ;
        RECT 2418.030 1429.925 2418.200 1430.425 ;
        RECT 2418.990 1429.925 2419.160 1430.425 ;
        RECT 2419.990 1429.925 2420.160 1430.425 ;
        RECT 2421.950 1429.925 2422.120 1430.425 ;
        RECT 2422.910 1429.925 2423.080 1430.425 ;
        RECT 2424.870 1429.925 2425.040 1430.425 ;
        RECT 2427.310 1429.925 2427.480 1430.425 ;
        RECT 2430.325 1429.695 2430.495 1430.425 ;
        RECT 2433.070 1429.695 2433.240 1430.425 ;
        RECT 2434.060 1429.700 2434.230 1430.430 ;
        RECT 2435.780 1430.425 2447.740 1430.430 ;
        RECT 2448.715 1430.425 2452.450 1430.430 ;
        RECT 2436.590 1429.925 2436.760 1430.425 ;
        RECT 2437.550 1429.925 2437.720 1430.425 ;
        RECT 2438.550 1429.925 2438.720 1430.425 ;
        RECT 2440.510 1429.925 2440.680 1430.425 ;
        RECT 2441.470 1429.925 2441.640 1430.425 ;
        RECT 2443.430 1429.925 2443.600 1430.425 ;
        RECT 2445.870 1429.925 2446.040 1430.425 ;
        RECT 2448.885 1429.695 2449.055 1430.425 ;
        RECT 2451.630 1429.695 2451.800 1430.425 ;
        RECT 2452.620 1429.700 2452.790 1430.430 ;
        RECT 2696.295 1430.095 2696.815 1430.635 ;
        RECT 2695.605 1429.005 2696.815 1430.095 ;
        RECT 2697.905 1429.005 2698.165 1430.145 ;
        RECT 2700.190 1429.005 2700.470 1429.805 ;
        RECT 2701.885 1429.005 2702.170 1429.805 ;
        RECT 2702.840 1429.005 2703.090 1430.145 ;
        RECT 2707.290 1429.440 2707.640 1430.690 ;
        RECT 2712.810 1429.440 2713.160 1430.690 ;
        RECT 2718.330 1429.440 2718.680 1430.690 ;
        RECT 2703.885 1429.005 2709.230 1429.440 ;
        RECT 2709.405 1429.005 2714.750 1429.440 ;
        RECT 2714.925 1429.005 2720.270 1429.440 ;
        RECT 2721.365 1429.005 2721.655 1430.170 ;
        RECT 2725.230 1429.440 2725.580 1430.690 ;
        RECT 2730.750 1429.440 2731.100 1430.690 ;
        RECT 2732.865 1430.095 2733.385 1430.635 ;
        RECT 2721.825 1429.005 2727.170 1429.440 ;
        RECT 2727.345 1429.005 2732.690 1429.440 ;
        RECT 2732.865 1429.005 2734.075 1430.095 ;
        RECT 2695.520 1428.835 2734.160 1429.005 ;
        RECT 2695.605 1427.745 2696.815 1428.835 ;
        RECT 2697.425 1428.075 2697.755 1428.835 ;
        RECT 2696.295 1427.205 2696.815 1427.745 ;
        RECT 2698.825 1427.695 2699.085 1428.835 ;
        RECT 2699.755 1427.695 2700.035 1428.835 ;
        RECT 2700.205 1428.400 2705.550 1428.835 ;
        RECT 2703.610 1427.150 2703.960 1428.400 ;
        RECT 2705.725 1427.745 2708.315 1428.835 ;
        RECT 2707.105 1427.225 2708.315 1427.745 ;
        RECT 2708.485 1427.670 2708.775 1428.835 ;
        RECT 2708.945 1428.400 2714.290 1428.835 ;
        RECT 2714.465 1428.400 2719.810 1428.835 ;
        RECT 2719.985 1428.400 2725.330 1428.835 ;
        RECT 2725.505 1428.400 2730.850 1428.835 ;
        RECT 2712.350 1427.150 2712.700 1428.400 ;
        RECT 2717.870 1427.150 2718.220 1428.400 ;
        RECT 2723.390 1427.150 2723.740 1428.400 ;
        RECT 2728.910 1427.150 2729.260 1428.400 ;
        RECT 2731.025 1427.745 2732.695 1428.835 ;
        RECT 2731.945 1427.225 2732.695 1427.745 ;
        RECT 2732.865 1427.745 2734.075 1428.835 ;
        RECT 2732.865 1427.205 2733.385 1427.745 ;
        RECT 2696.295 1424.655 2696.815 1425.195 ;
        RECT 2695.605 1423.565 2696.815 1424.655 ;
        RECT 2697.735 1423.565 2697.905 1424.325 ;
        RECT 2700.275 1423.565 2700.445 1424.705 ;
        RECT 2704.530 1424.000 2704.880 1425.250 ;
        RECT 2710.050 1424.000 2710.400 1425.250 ;
        RECT 2715.570 1424.000 2715.920 1425.250 ;
        RECT 2719.505 1424.655 2721.195 1425.175 ;
        RECT 2701.125 1423.565 2706.470 1424.000 ;
        RECT 2706.645 1423.565 2711.990 1424.000 ;
        RECT 2712.165 1423.565 2717.510 1424.000 ;
        RECT 2717.685 1423.565 2721.195 1424.655 ;
        RECT 2721.365 1423.565 2721.655 1424.730 ;
        RECT 2725.230 1424.000 2725.580 1425.250 ;
        RECT 2730.750 1424.000 2731.100 1425.250 ;
        RECT 2732.865 1424.655 2733.385 1425.195 ;
        RECT 2721.825 1423.565 2727.170 1424.000 ;
        RECT 2727.345 1423.565 2732.690 1424.000 ;
        RECT 2732.865 1423.565 2734.075 1424.655 ;
        RECT 2695.520 1423.395 2734.160 1423.565 ;
        RECT 2695.605 1422.305 2696.815 1423.395 ;
        RECT 2697.425 1422.635 2697.755 1423.395 ;
        RECT 2698.365 1422.960 2703.710 1423.395 ;
        RECT 2696.295 1421.765 2696.815 1422.305 ;
        RECT 2701.770 1421.710 2702.120 1422.960 ;
        RECT 2703.885 1422.305 2707.395 1423.395 ;
        RECT 2705.705 1421.785 2707.395 1422.305 ;
        RECT 2708.485 1422.230 2708.775 1423.395 ;
        RECT 2708.945 1422.960 2714.290 1423.395 ;
        RECT 2714.465 1422.960 2719.810 1423.395 ;
        RECT 2719.985 1422.960 2725.330 1423.395 ;
        RECT 2725.505 1422.960 2730.850 1423.395 ;
        RECT 2712.350 1421.710 2712.700 1422.960 ;
        RECT 2717.870 1421.710 2718.220 1422.960 ;
        RECT 2723.390 1421.710 2723.740 1422.960 ;
        RECT 2728.910 1421.710 2729.260 1422.960 ;
        RECT 2731.025 1422.305 2732.695 1423.395 ;
        RECT 2731.945 1421.785 2732.695 1422.305 ;
        RECT 2732.865 1422.305 2734.075 1423.395 ;
        RECT 2732.865 1421.765 2733.385 1422.305 ;
        RECT 2696.295 1419.215 2696.815 1419.755 ;
        RECT 2522.135 1418.340 2523.935 1418.510 ;
        RECT 2522.830 1417.615 2523.160 1418.340 ;
        RECT 2695.605 1418.125 2696.815 1419.215 ;
        RECT 2700.390 1418.560 2700.740 1419.810 ;
        RECT 2705.910 1418.560 2706.260 1419.810 ;
        RECT 2711.430 1418.560 2711.780 1419.810 ;
        RECT 2716.950 1418.560 2717.300 1419.810 ;
        RECT 2719.985 1419.215 2720.735 1419.735 ;
        RECT 2696.985 1418.125 2702.330 1418.560 ;
        RECT 2702.505 1418.125 2707.850 1418.560 ;
        RECT 2708.025 1418.125 2713.370 1418.560 ;
        RECT 2713.545 1418.125 2718.890 1418.560 ;
        RECT 2719.065 1418.125 2720.735 1419.215 ;
        RECT 2721.365 1418.125 2721.655 1419.290 ;
        RECT 2725.230 1418.560 2725.580 1419.810 ;
        RECT 2730.750 1418.560 2731.100 1419.810 ;
        RECT 2732.865 1419.215 2733.385 1419.755 ;
        RECT 2721.825 1418.125 2727.170 1418.560 ;
        RECT 2727.345 1418.125 2732.690 1418.560 ;
        RECT 2732.865 1418.125 2734.075 1419.215 ;
        RECT 2695.520 1417.955 2734.160 1418.125 ;
        RECT 2695.605 1416.865 2696.815 1417.955 ;
        RECT 2697.425 1417.195 2697.755 1417.955 ;
        RECT 2698.365 1417.520 2703.710 1417.955 ;
        RECT 2696.295 1416.325 2696.815 1416.865 ;
        RECT 2701.770 1416.270 2702.120 1417.520 ;
        RECT 2703.885 1416.865 2707.395 1417.955 ;
        RECT 2705.705 1416.345 2707.395 1416.865 ;
        RECT 2708.485 1416.790 2708.775 1417.955 ;
        RECT 2708.945 1417.520 2714.290 1417.955 ;
        RECT 2714.465 1417.520 2719.810 1417.955 ;
        RECT 2719.985 1417.520 2725.330 1417.955 ;
        RECT 2725.505 1417.520 2730.850 1417.955 ;
        RECT 2712.350 1416.270 2712.700 1417.520 ;
        RECT 2717.870 1416.270 2718.220 1417.520 ;
        RECT 2723.390 1416.270 2723.740 1417.520 ;
        RECT 2728.910 1416.270 2729.260 1417.520 ;
        RECT 2731.025 1416.865 2732.695 1417.955 ;
        RECT 2731.945 1416.345 2732.695 1416.865 ;
        RECT 2732.865 1416.865 2734.075 1417.955 ;
        RECT 2732.865 1416.325 2733.385 1416.865 ;
        RECT 2696.295 1413.775 2696.815 1414.315 ;
        RECT 2695.605 1412.685 2696.815 1413.775 ;
        RECT 2700.390 1413.120 2700.740 1414.370 ;
        RECT 2705.910 1413.120 2706.260 1414.370 ;
        RECT 2711.430 1413.120 2711.780 1414.370 ;
        RECT 2716.950 1413.120 2717.300 1414.370 ;
        RECT 2719.985 1413.775 2720.735 1414.295 ;
        RECT 2696.985 1412.685 2702.330 1413.120 ;
        RECT 2702.505 1412.685 2707.850 1413.120 ;
        RECT 2708.025 1412.685 2713.370 1413.120 ;
        RECT 2713.545 1412.685 2718.890 1413.120 ;
        RECT 2719.065 1412.685 2720.735 1413.775 ;
        RECT 2721.365 1412.685 2721.655 1413.850 ;
        RECT 2725.230 1413.120 2725.580 1414.370 ;
        RECT 2730.750 1413.120 2731.100 1414.370 ;
        RECT 2732.865 1413.775 2733.385 1414.315 ;
        RECT 2721.825 1412.685 2727.170 1413.120 ;
        RECT 2727.345 1412.685 2732.690 1413.120 ;
        RECT 2732.865 1412.685 2734.075 1413.775 ;
        RECT 2695.520 1412.515 2734.160 1412.685 ;
        RECT 2695.605 1411.425 2696.815 1412.515 ;
        RECT 2697.425 1411.755 2697.755 1412.515 ;
        RECT 2698.805 1411.755 2699.135 1412.515 ;
        RECT 2699.745 1412.080 2705.090 1412.515 ;
        RECT 2522.135 1410.810 2523.935 1410.980 ;
        RECT 2696.295 1410.885 2696.815 1411.425 ;
        RECT 2703.150 1410.830 2703.500 1412.080 ;
        RECT 2705.265 1411.425 2707.855 1412.515 ;
        RECT 2706.645 1410.905 2707.855 1411.425 ;
        RECT 2708.485 1411.350 2708.775 1412.515 ;
        RECT 2708.945 1412.080 2714.290 1412.515 ;
        RECT 2714.465 1412.080 2719.810 1412.515 ;
        RECT 2712.350 1410.830 2712.700 1412.080 ;
        RECT 2717.870 1410.830 2718.220 1412.080 ;
        RECT 2719.985 1411.425 2721.195 1412.515 ;
        RECT 2720.675 1410.885 2721.195 1411.425 ;
        RECT 2721.365 1411.350 2721.655 1412.515 ;
        RECT 2721.825 1412.080 2727.170 1412.515 ;
        RECT 2727.345 1412.080 2732.690 1412.515 ;
        RECT 2725.230 1410.830 2725.580 1412.080 ;
        RECT 2730.750 1410.830 2731.100 1412.080 ;
        RECT 2732.865 1411.425 2734.075 1412.515 ;
        RECT 2732.865 1410.885 2733.385 1411.425 ;
        RECT 2522.830 1410.085 2523.160 1410.810 ;
        RECT 2522.135 1404.830 2523.935 1405.000 ;
        RECT 2522.830 1404.105 2523.160 1404.830 ;
        RECT 2522.135 1396.415 2523.935 1396.585 ;
        RECT 2522.830 1395.690 2523.160 1396.415 ;
        RECT 2881.580 1363.140 2883.380 1363.310 ;
        RECT 2882.775 1362.415 2883.105 1363.140 ;
        RECT 2370.030 1335.050 2370.205 1335.600 ;
        RECT 2370.030 1333.450 2370.200 1335.050 ;
        RECT 2368.215 1332.040 2368.385 1332.770 ;
        RECT 2370.030 1332.310 2370.205 1333.450 ;
        RECT 2370.030 1332.040 2370.200 1332.310 ;
        RECT 2375.730 1332.040 2375.900 1332.770 ;
        RECT 2381.345 1332.040 2381.515 1332.770 ;
        RECT 2384.090 1332.040 2384.260 1332.770 ;
        RECT 2385.080 1332.040 2385.250 1332.770 ;
        RECT 2390.990 1332.040 2391.160 1332.770 ;
        RECT 2396.605 1332.040 2396.775 1332.770 ;
        RECT 2399.350 1332.040 2399.520 1332.770 ;
        RECT 2400.340 1332.040 2400.510 1332.770 ;
        RECT 2406.250 1332.040 2406.420 1332.770 ;
        RECT 2411.865 1332.040 2412.035 1332.770 ;
        RECT 2414.610 1332.040 2414.780 1332.770 ;
        RECT 2415.600 1332.040 2415.770 1332.770 ;
        RECT 2421.510 1332.040 2421.680 1332.770 ;
        RECT 2427.125 1332.040 2427.295 1332.770 ;
        RECT 2429.870 1332.040 2430.040 1332.770 ;
        RECT 2430.860 1332.040 2431.030 1332.770 ;
        RECT 2436.770 1332.040 2436.940 1332.770 ;
        RECT 2442.385 1332.040 2442.555 1332.770 ;
        RECT 2445.130 1332.040 2445.300 1332.770 ;
        RECT 2446.120 1332.040 2446.290 1332.770 ;
        RECT 2368.045 1332.035 2370.795 1332.040 ;
        RECT 2375.560 1332.035 2378.310 1332.040 ;
        RECT 2381.175 1332.035 2385.900 1332.040 ;
        RECT 2390.820 1332.035 2393.570 1332.040 ;
        RECT 2396.435 1332.035 2401.160 1332.040 ;
        RECT 2406.080 1332.035 2408.830 1332.040 ;
        RECT 2411.695 1332.035 2416.420 1332.040 ;
        RECT 2421.340 1332.035 2424.090 1332.040 ;
        RECT 2426.955 1332.035 2431.680 1332.040 ;
        RECT 2436.600 1332.035 2439.350 1332.040 ;
        RECT 2442.215 1332.035 2446.940 1332.040 ;
        RECT 2343.000 1330.435 2447.095 1332.035 ;
        RECT 2371.545 1330.430 2386.055 1330.435 ;
        RECT 2386.805 1330.430 2401.315 1330.435 ;
        RECT 2402.065 1330.430 2416.575 1330.435 ;
        RECT 2417.325 1330.430 2431.835 1330.435 ;
        RECT 2432.585 1330.430 2447.095 1330.435 ;
        RECT 2371.545 1330.425 2380.285 1330.430 ;
        RECT 2381.175 1330.425 2385.895 1330.430 ;
        RECT 2386.805 1330.425 2395.545 1330.430 ;
        RECT 2396.435 1330.425 2401.155 1330.430 ;
        RECT 2402.065 1330.425 2410.805 1330.430 ;
        RECT 2411.695 1330.425 2416.415 1330.430 ;
        RECT 2417.325 1330.425 2426.065 1330.430 ;
        RECT 2426.955 1330.425 2431.675 1330.430 ;
        RECT 2432.585 1330.425 2441.325 1330.430 ;
        RECT 2442.215 1330.425 2446.935 1330.430 ;
        RECT 2372.335 1329.925 2372.505 1330.425 ;
        RECT 2374.255 1329.925 2374.425 1330.425 ;
        RECT 2375.715 1329.925 2375.885 1330.425 ;
        RECT 2376.655 1329.925 2376.825 1330.425 ;
        RECT 2378.575 1329.925 2378.745 1330.425 ;
        RECT 2381.345 1329.695 2381.515 1330.425 ;
        RECT 2384.090 1329.695 2384.260 1330.425 ;
        RECT 2385.075 1329.695 2385.245 1330.425 ;
        RECT 2387.595 1329.925 2387.765 1330.425 ;
        RECT 2389.515 1329.925 2389.685 1330.425 ;
        RECT 2390.975 1329.925 2391.145 1330.425 ;
        RECT 2391.915 1329.925 2392.085 1330.425 ;
        RECT 2393.835 1329.925 2394.005 1330.425 ;
        RECT 2396.605 1329.695 2396.775 1330.425 ;
        RECT 2399.350 1329.695 2399.520 1330.425 ;
        RECT 2400.335 1329.695 2400.505 1330.425 ;
        RECT 2402.855 1329.925 2403.025 1330.425 ;
        RECT 2404.775 1329.925 2404.945 1330.425 ;
        RECT 2406.235 1329.925 2406.405 1330.425 ;
        RECT 2407.175 1329.925 2407.345 1330.425 ;
        RECT 2409.095 1329.925 2409.265 1330.425 ;
        RECT 2411.865 1329.695 2412.035 1330.425 ;
        RECT 2414.610 1329.695 2414.780 1330.425 ;
        RECT 2415.595 1329.695 2415.765 1330.425 ;
        RECT 2418.115 1329.925 2418.285 1330.425 ;
        RECT 2420.035 1329.925 2420.205 1330.425 ;
        RECT 2421.495 1329.925 2421.665 1330.425 ;
        RECT 2422.435 1329.925 2422.605 1330.425 ;
        RECT 2424.355 1329.925 2424.525 1330.425 ;
        RECT 2427.125 1329.695 2427.295 1330.425 ;
        RECT 2429.870 1329.695 2430.040 1330.425 ;
        RECT 2430.855 1329.695 2431.025 1330.425 ;
        RECT 2433.375 1329.925 2433.545 1330.425 ;
        RECT 2435.295 1329.925 2435.465 1330.425 ;
        RECT 2436.755 1329.925 2436.925 1330.425 ;
        RECT 2437.695 1329.925 2437.865 1330.425 ;
        RECT 2439.615 1329.925 2439.785 1330.425 ;
        RECT 2442.385 1329.695 2442.555 1330.425 ;
        RECT 2445.130 1329.695 2445.300 1330.425 ;
        RECT 2446.115 1329.695 2446.285 1330.425 ;
        RECT 2881.580 1163.900 2883.380 1164.070 ;
        RECT 2882.775 1163.175 2883.105 1163.900 ;
      LAYER met1 ;
        RECT 1622.805 3510.325 1624.185 3510.360 ;
        RECT 1622.805 3510.205 1628.315 3510.325 ;
        RECT 1622.405 3510.035 1628.315 3510.205 ;
        RECT 1262.805 3509.875 1264.185 3509.910 ;
        RECT 1622.805 3509.880 1628.315 3510.035 ;
        RECT 1262.805 3509.755 1268.315 3509.875 ;
        RECT 1623.995 3509.845 1628.315 3509.880 ;
        RECT 1262.405 3509.585 1268.315 3509.755 ;
        RECT 1262.805 3509.430 1268.315 3509.585 ;
        RECT 1263.995 3509.395 1268.315 3509.430 ;
        RECT 1264.970 3508.275 1268.070 3509.395 ;
        RECT 1624.970 3508.725 1628.070 3509.845 ;
        RECT 2522.805 3508.730 2524.185 3508.765 ;
        RECT 2522.805 3508.610 2528.315 3508.730 ;
        RECT 2522.405 3508.440 2528.315 3508.610 ;
        RECT 1802.805 3508.405 1804.185 3508.440 ;
        RECT 1802.805 3508.285 1808.315 3508.405 ;
        RECT 2522.805 3508.285 2528.315 3508.440 ;
        RECT 1802.405 3508.115 1808.315 3508.285 ;
        RECT 2523.995 3508.250 2528.315 3508.285 ;
        RECT 1802.805 3507.960 1808.315 3508.115 ;
        RECT 1803.995 3507.925 1808.315 3507.960 ;
        RECT 2162.805 3508.045 2164.185 3508.080 ;
        RECT 2162.805 3507.925 2168.315 3508.045 ;
        RECT 1804.970 3506.805 1808.070 3507.925 ;
        RECT 2162.405 3507.755 2168.315 3507.925 ;
        RECT 2162.805 3507.600 2168.315 3507.755 ;
        RECT 2163.995 3507.565 2168.315 3507.600 ;
        RECT 2164.970 3506.445 2168.070 3507.565 ;
        RECT 2524.970 3507.130 2528.070 3508.250 ;
        RECT 2884.970 3488.465 2888.070 3489.585 ;
        RECT 2882.000 3488.310 2888.235 3488.465 ;
        RECT 2881.580 3488.140 2888.235 3488.310 ;
        RECT 2882.000 3487.985 2888.235 3488.140 ;
        RECT 2884.970 3222.585 2888.070 3223.705 ;
        RECT 2882.000 3222.430 2888.235 3222.585 ;
        RECT 2881.580 3222.260 2888.235 3222.430 ;
        RECT 2882.000 3222.105 2888.235 3222.260 ;
        RECT 2884.970 2957.385 2888.070 2958.505 ;
        RECT 2882.000 2957.230 2888.235 2957.385 ;
        RECT 2881.580 2957.060 2888.235 2957.230 ;
        RECT 2882.000 2956.905 2888.235 2957.060 ;
        RECT 2884.970 2691.505 2888.070 2692.625 ;
        RECT 2882.000 2691.350 2888.235 2691.505 ;
        RECT 2881.580 2691.180 2888.235 2691.350 ;
        RECT 2882.000 2691.025 2888.235 2691.180 ;
        RECT 2885.110 2426.680 2887.930 2426.820 ;
        RECT 2884.970 2425.625 2888.070 2426.680 ;
        RECT 2882.000 2425.470 2888.235 2425.625 ;
        RECT 2881.580 2425.300 2888.235 2425.470 ;
        RECT 2882.000 2425.145 2888.235 2425.300 ;
        RECT 2359.980 2254.135 2360.270 2254.165 ;
        RECT 2359.810 2253.965 2360.270 2254.135 ;
        RECT 2359.980 2253.935 2360.270 2253.965 ;
        RECT 2343.000 2250.965 2364.620 2252.025 ;
        RECT 2366.130 2250.965 2366.280 2250.970 ;
        RECT 2371.450 2250.965 2381.205 2252.030 ;
        RECT 2382.715 2250.965 2382.865 2250.970 ;
        RECT 2388.035 2250.965 2397.790 2252.030 ;
        RECT 2399.300 2250.965 2399.450 2250.970 ;
        RECT 2404.620 2250.965 2414.375 2252.030 ;
        RECT 2415.885 2250.965 2416.035 2250.970 ;
        RECT 2421.205 2250.965 2430.960 2252.030 ;
        RECT 2432.465 2250.965 2432.615 2250.970 ;
        RECT 2437.785 2250.965 2443.725 2252.030 ;
        RECT 2343.000 2250.485 2443.725 2250.965 ;
        RECT 2343.000 2250.425 2364.620 2250.485 ;
        RECT 2371.320 2250.430 2381.205 2250.485 ;
        RECT 2387.905 2250.430 2397.790 2250.485 ;
        RECT 2404.490 2250.430 2414.375 2250.485 ;
        RECT 2421.075 2250.430 2430.960 2250.485 ;
        RECT 2437.655 2250.430 2443.725 2250.485 ;
        RECT 2377.225 2250.425 2381.205 2250.430 ;
        RECT 2393.805 2250.425 2397.790 2250.430 ;
        RECT 2410.385 2250.425 2414.375 2250.430 ;
        RECT 2426.965 2250.425 2430.955 2250.430 ;
        RECT 2695.520 2213.960 2734.160 2214.440 ;
        RECT 2695.520 2208.520 2734.160 2209.000 ;
        RECT 2695.520 2203.080 2734.160 2203.560 ;
        RECT 2695.520 2197.640 2734.160 2198.120 ;
        RECT 2695.520 2192.200 2734.160 2192.680 ;
        RECT 2695.520 2186.760 2734.160 2187.240 ;
        RECT 2695.520 2181.320 2734.160 2181.800 ;
        RECT 2695.520 2175.880 2734.160 2176.360 ;
        RECT 2695.520 2170.440 2734.160 2170.920 ;
        RECT 2695.520 2165.000 2734.160 2165.480 ;
        RECT 2359.995 2162.145 2360.285 2162.175 ;
        RECT 2359.825 2161.975 2360.285 2162.145 ;
        RECT 2359.995 2161.945 2360.285 2161.975 ;
        RECT 2884.970 2160.425 2888.070 2161.545 ;
        RECT 2882.000 2160.270 2888.235 2160.425 ;
        RECT 2881.580 2160.100 2888.235 2160.270 ;
        RECT 2358.070 2160.030 2360.820 2160.035 ;
        RECT 2373.165 2160.030 2377.890 2160.035 ;
        RECT 2390.385 2160.030 2395.110 2160.035 ;
        RECT 2407.605 2160.030 2412.330 2160.035 ;
        RECT 2424.825 2160.030 2429.550 2160.035 ;
        RECT 2442.045 2160.030 2446.770 2160.035 ;
        RECT 2358.070 2160.025 2364.495 2160.030 ;
        RECT 2343.015 2160.000 2364.500 2160.025 ;
        RECT 2371.960 2160.000 2381.715 2160.030 ;
        RECT 2389.180 2160.000 2398.935 2160.030 ;
        RECT 2406.400 2160.000 2416.155 2160.030 ;
        RECT 2423.620 2160.000 2433.375 2160.030 ;
        RECT 2343.015 2158.965 2364.625 2160.000 ;
        RECT 2371.960 2158.965 2381.845 2160.000 ;
        RECT 2389.180 2158.965 2399.065 2160.000 ;
        RECT 2406.400 2158.965 2416.285 2160.000 ;
        RECT 2423.620 2158.965 2433.505 2160.000 ;
        RECT 2440.840 2158.965 2446.925 2160.030 ;
        RECT 2695.520 2159.560 2734.160 2160.040 ;
        RECT 2882.000 2159.945 2888.235 2160.100 ;
        RECT 2343.015 2158.485 2446.925 2158.965 ;
        RECT 2343.015 2158.425 2364.785 2158.485 ;
        RECT 2372.055 2158.430 2382.005 2158.485 ;
        RECT 2389.275 2158.430 2399.225 2158.485 ;
        RECT 2406.495 2158.430 2416.445 2158.485 ;
        RECT 2423.715 2158.430 2433.665 2158.485 ;
        RECT 2440.935 2158.430 2446.925 2158.485 ;
        RECT 2373.165 2158.425 2382.005 2158.430 ;
        RECT 2390.385 2158.425 2399.225 2158.430 ;
        RECT 2407.605 2158.425 2416.445 2158.430 ;
        RECT 2424.825 2158.425 2433.665 2158.430 ;
        RECT 2442.045 2158.425 2446.765 2158.430 ;
        RECT 2695.520 2154.120 2734.160 2154.600 ;
        RECT 2695.520 2148.680 2734.160 2149.160 ;
        RECT 2695.520 2143.240 2734.160 2143.720 ;
        RECT 2524.970 2136.915 2528.070 2138.035 ;
        RECT 2695.520 2137.800 2734.160 2138.280 ;
        RECT 2522.555 2136.760 2528.245 2136.915 ;
        RECT 2522.135 2136.590 2528.245 2136.760 ;
        RECT 2522.555 2136.435 2528.245 2136.590 ;
        RECT 2695.520 2132.360 2734.160 2132.840 ;
        RECT 2524.970 2129.385 2528.070 2130.505 ;
        RECT 2522.555 2129.230 2528.245 2129.385 ;
        RECT 2522.135 2129.060 2528.245 2129.230 ;
        RECT 2522.555 2128.905 2528.245 2129.060 ;
        RECT 2524.970 2123.405 2528.070 2124.525 ;
        RECT 2522.555 2123.250 2528.245 2123.405 ;
        RECT 2522.135 2123.080 2528.245 2123.250 ;
        RECT 2522.555 2122.925 2528.245 2123.080 ;
        RECT 2524.970 2117.460 2528.070 2118.580 ;
        RECT 2522.555 2117.305 2528.245 2117.460 ;
        RECT 2522.135 2117.135 2528.245 2117.305 ;
        RECT 2522.555 2116.980 2528.245 2117.135 ;
        RECT 2524.970 2111.815 2528.070 2112.935 ;
        RECT 2522.555 2111.660 2528.245 2111.815 ;
        RECT 2522.135 2111.490 2528.245 2111.660 ;
        RECT 2522.555 2111.335 2528.245 2111.490 ;
        RECT 2524.970 2105.810 2528.070 2106.930 ;
        RECT 2522.555 2105.655 2528.245 2105.810 ;
        RECT 2522.135 2105.485 2528.245 2105.655 ;
        RECT 2522.555 2105.330 2528.245 2105.485 ;
        RECT 2359.975 2057.145 2360.265 2057.175 ;
        RECT 2359.805 2056.975 2360.265 2057.145 ;
        RECT 2359.975 2056.945 2360.265 2056.975 ;
        RECT 2358.050 2055.030 2360.800 2055.035 ;
        RECT 2366.630 2055.030 2369.380 2055.035 ;
        RECT 2372.245 2055.030 2375.980 2055.035 ;
        RECT 2382.955 2055.030 2385.705 2055.035 ;
        RECT 2388.570 2055.030 2392.305 2055.035 ;
        RECT 2399.280 2055.030 2402.030 2055.035 ;
        RECT 2404.895 2055.030 2408.630 2055.035 ;
        RECT 2415.605 2055.030 2418.355 2055.035 ;
        RECT 2421.220 2055.030 2424.955 2055.035 ;
        RECT 2431.930 2055.030 2434.680 2055.035 ;
        RECT 2437.545 2055.030 2441.280 2055.035 ;
        RECT 2343.005 2053.430 2442.425 2055.030 ;
        RECT 2361.540 2053.395 2371.200 2053.430 ;
        RECT 2372.245 2053.425 2375.980 2053.430 ;
        RECT 2377.865 2053.395 2387.525 2053.430 ;
        RECT 2388.570 2053.425 2392.305 2053.430 ;
        RECT 2394.190 2053.395 2403.850 2053.430 ;
        RECT 2404.895 2053.425 2408.630 2053.430 ;
        RECT 2410.515 2053.395 2420.175 2053.430 ;
        RECT 2421.220 2053.425 2424.955 2053.430 ;
        RECT 2426.840 2053.395 2436.500 2053.430 ;
        RECT 2437.545 2053.425 2441.280 2053.430 ;
        RECT 2695.520 2033.960 2734.160 2034.440 ;
        RECT 2695.520 2028.520 2734.160 2029.000 ;
        RECT 2695.520 2023.080 2734.160 2023.560 ;
        RECT 2695.520 2017.640 2734.160 2018.120 ;
        RECT 2695.520 2012.200 2734.160 2012.680 ;
        RECT 2695.520 2006.760 2734.160 2007.240 ;
        RECT 2695.520 2001.320 2734.160 2001.800 ;
        RECT 2695.520 1995.880 2734.160 1996.360 ;
        RECT 2695.520 1990.440 2734.160 1990.920 ;
        RECT 2524.970 1984.660 2528.070 1985.780 ;
        RECT 2695.520 1985.000 2734.160 1985.480 ;
        RECT 2522.555 1984.505 2528.245 1984.660 ;
        RECT 2522.135 1984.335 2528.245 1984.505 ;
        RECT 2522.555 1984.180 2528.245 1984.335 ;
        RECT 2695.520 1979.560 2734.160 1980.040 ;
        RECT 2524.970 1977.130 2528.070 1978.250 ;
        RECT 2522.555 1976.975 2528.245 1977.130 ;
        RECT 2522.135 1976.805 2528.245 1976.975 ;
        RECT 2522.555 1976.650 2528.245 1976.805 ;
        RECT 2695.520 1974.120 2734.160 1974.600 ;
        RECT 2524.970 1971.150 2528.070 1972.270 ;
        RECT 2522.555 1970.995 2528.245 1971.150 ;
        RECT 2522.135 1970.825 2528.245 1970.995 ;
        RECT 2522.555 1970.670 2528.245 1970.825 ;
        RECT 2695.520 1968.680 2734.160 1969.160 ;
        RECT 2524.970 1965.205 2528.070 1966.325 ;
        RECT 2522.555 1965.050 2528.245 1965.205 ;
        RECT 2522.135 1964.880 2528.245 1965.050 ;
        RECT 2522.555 1964.725 2528.245 1964.880 ;
        RECT 2695.520 1963.240 2734.160 1963.720 ;
        RECT 2524.970 1959.560 2528.070 1960.680 ;
        RECT 2522.555 1959.405 2528.245 1959.560 ;
        RECT 2522.135 1959.235 2528.245 1959.405 ;
        RECT 2522.555 1959.080 2528.245 1959.235 ;
        RECT 2695.520 1957.800 2734.160 1958.280 ;
        RECT 2524.970 1953.555 2528.070 1954.675 ;
        RECT 2522.555 1953.400 2528.245 1953.555 ;
        RECT 2522.135 1953.230 2528.245 1953.400 ;
        RECT 2522.555 1953.075 2528.245 1953.230 ;
        RECT 2695.520 1952.360 2734.160 1952.840 ;
        RECT 2359.975 1952.150 2360.265 1952.180 ;
        RECT 2359.805 1951.980 2360.265 1952.150 ;
        RECT 2359.975 1951.950 2360.265 1951.980 ;
        RECT 2343.000 1950.025 2453.600 1950.050 ;
        RECT 2343.000 1948.450 2453.615 1950.025 ;
        RECT 2360.815 1948.425 2453.615 1948.450 ;
        RECT 2361.545 1948.395 2373.505 1948.425 ;
        RECT 2380.105 1948.395 2392.065 1948.425 ;
        RECT 2398.665 1948.395 2410.625 1948.425 ;
        RECT 2417.225 1948.395 2429.185 1948.425 ;
        RECT 2435.785 1948.395 2447.745 1948.425 ;
        RECT 2884.970 1894.545 2888.070 1895.665 ;
        RECT 2882.000 1894.390 2888.235 1894.545 ;
        RECT 2881.580 1894.220 2888.235 1894.390 ;
        RECT 2882.000 1894.065 2888.235 1894.220 ;
        RECT 2695.520 1853.960 2734.160 1854.440 ;
        RECT 2695.520 1848.520 2734.160 1849.000 ;
        RECT 2695.520 1843.080 2734.160 1843.560 ;
        RECT 2695.520 1837.640 2734.160 1838.120 ;
        RECT 2695.520 1832.200 2734.160 1832.680 ;
        RECT 2695.520 1826.760 2734.160 1827.240 ;
        RECT 2695.520 1821.320 2734.160 1821.800 ;
        RECT 2695.520 1815.880 2734.160 1816.360 ;
        RECT 2695.520 1810.440 2734.160 1810.920 ;
        RECT 2524.970 1807.690 2528.070 1808.810 ;
        RECT 2522.555 1807.535 2528.245 1807.690 ;
        RECT 2522.135 1807.365 2528.245 1807.535 ;
        RECT 2522.555 1807.210 2528.245 1807.365 ;
        RECT 2695.520 1805.000 2734.160 1805.480 ;
        RECT 2524.970 1800.160 2528.070 1801.280 ;
        RECT 2522.555 1800.005 2528.245 1800.160 ;
        RECT 2522.135 1799.835 2528.245 1800.005 ;
        RECT 2522.555 1799.680 2528.245 1799.835 ;
        RECT 2695.520 1799.560 2734.160 1800.040 ;
        RECT 2524.970 1794.180 2528.070 1795.300 ;
        RECT 2522.555 1794.025 2528.245 1794.180 ;
        RECT 2695.520 1794.120 2734.160 1794.600 ;
        RECT 2522.135 1793.855 2528.245 1794.025 ;
        RECT 2522.555 1793.700 2528.245 1793.855 ;
        RECT 2369.920 1789.150 2370.210 1789.180 ;
        RECT 2369.750 1788.980 2370.210 1789.150 ;
        RECT 2369.920 1788.950 2370.210 1788.980 ;
        RECT 2524.970 1788.235 2528.070 1789.355 ;
        RECT 2695.520 1788.680 2734.160 1789.160 ;
        RECT 2522.555 1788.080 2528.245 1788.235 ;
        RECT 2522.135 1787.910 2528.245 1788.080 ;
        RECT 2522.555 1787.755 2528.245 1787.910 ;
        RECT 2367.995 1787.035 2370.745 1787.040 ;
        RECT 2375.510 1787.035 2378.260 1787.040 ;
        RECT 2381.125 1787.035 2385.850 1787.040 ;
        RECT 2390.770 1787.035 2393.520 1787.040 ;
        RECT 2396.385 1787.035 2401.110 1787.040 ;
        RECT 2406.030 1787.035 2408.780 1787.040 ;
        RECT 2411.645 1787.035 2416.370 1787.040 ;
        RECT 2421.290 1787.035 2424.040 1787.040 ;
        RECT 2426.905 1787.035 2431.630 1787.040 ;
        RECT 2436.550 1787.035 2439.300 1787.040 ;
        RECT 2442.165 1787.035 2446.890 1787.040 ;
        RECT 2343.000 1785.435 2447.045 1787.035 ;
        RECT 2371.495 1785.430 2386.005 1785.435 ;
        RECT 2386.755 1785.430 2401.265 1785.435 ;
        RECT 2402.015 1785.430 2416.525 1785.435 ;
        RECT 2417.275 1785.430 2431.785 1785.435 ;
        RECT 2432.535 1785.430 2447.045 1785.435 ;
        RECT 2371.495 1785.395 2380.235 1785.430 ;
        RECT 2381.125 1785.425 2385.845 1785.430 ;
        RECT 2386.755 1785.395 2395.495 1785.430 ;
        RECT 2396.385 1785.425 2401.105 1785.430 ;
        RECT 2402.015 1785.395 2410.755 1785.430 ;
        RECT 2411.645 1785.425 2416.365 1785.430 ;
        RECT 2417.275 1785.395 2426.015 1785.430 ;
        RECT 2426.905 1785.425 2431.625 1785.430 ;
        RECT 2432.535 1785.395 2441.275 1785.430 ;
        RECT 2442.165 1785.425 2446.885 1785.430 ;
        RECT 2524.970 1782.590 2528.070 1783.710 ;
        RECT 2695.520 1783.240 2734.160 1783.720 ;
        RECT 2522.555 1782.435 2528.245 1782.590 ;
        RECT 2522.135 1782.265 2528.245 1782.435 ;
        RECT 2522.555 1782.110 2528.245 1782.265 ;
        RECT 2695.520 1777.800 2734.160 1778.280 ;
        RECT 2695.520 1772.360 2734.160 1772.840 ;
        RECT 2524.970 1771.120 2528.070 1772.240 ;
        RECT 2522.555 1770.965 2528.245 1771.120 ;
        RECT 2522.135 1770.795 2528.245 1770.965 ;
        RECT 2522.555 1770.640 2528.245 1770.795 ;
        RECT 2360.340 1709.135 2360.630 1709.165 ;
        RECT 2360.170 1708.965 2360.630 1709.135 ;
        RECT 2360.340 1708.935 2360.630 1708.965 ;
        RECT 2371.810 1707.030 2377.750 1707.040 ;
        RECT 2388.395 1707.030 2394.335 1707.040 ;
        RECT 2404.980 1707.035 2410.920 1707.045 ;
        RECT 2421.565 1707.035 2427.505 1707.050 ;
        RECT 2404.980 1707.030 2414.495 1707.035 ;
        RECT 2421.565 1707.030 2431.075 1707.035 ;
        RECT 2343.000 1705.965 2364.965 1707.025 ;
        RECT 2366.490 1705.965 2366.640 1705.970 ;
        RECT 2371.810 1705.965 2381.575 1707.030 ;
        RECT 2388.395 1705.970 2398.160 1707.030 ;
        RECT 2404.980 1705.975 2414.745 1707.030 ;
        RECT 2416.245 1705.975 2416.395 1705.980 ;
        RECT 2421.565 1705.975 2431.330 1707.030 ;
        RECT 2432.825 1705.975 2432.975 1705.980 ;
        RECT 2438.145 1705.975 2444.085 1707.050 ;
        RECT 2399.660 1705.970 2399.810 1705.975 ;
        RECT 2404.980 1705.970 2444.085 1705.975 ;
        RECT 2383.075 1705.965 2383.225 1705.970 ;
        RECT 2388.395 1705.965 2444.085 1705.970 ;
        RECT 2343.000 1705.495 2444.085 1705.965 ;
        RECT 2343.000 1705.490 2414.745 1705.495 ;
        RECT 2343.000 1705.485 2398.160 1705.490 ;
        RECT 2343.000 1705.425 2364.965 1705.485 ;
        RECT 2371.680 1705.445 2381.575 1705.485 ;
        RECT 2388.265 1705.445 2398.160 1705.485 ;
        RECT 2404.850 1705.450 2414.745 1705.490 ;
        RECT 2421.435 1705.455 2431.330 1705.495 ;
        RECT 2438.015 1705.455 2444.085 1705.495 ;
        RECT 2371.685 1705.430 2381.575 1705.445 ;
        RECT 2388.270 1705.430 2398.160 1705.445 ;
        RECT 2404.855 1705.435 2414.745 1705.450 ;
        RECT 2421.440 1705.440 2431.330 1705.455 ;
        RECT 2438.020 1705.440 2444.085 1705.455 ;
        RECT 2404.980 1705.430 2414.745 1705.435 ;
        RECT 2421.565 1705.430 2431.330 1705.440 ;
        RECT 2438.145 1705.430 2444.085 1705.440 ;
        RECT 2377.750 1705.425 2381.475 1705.430 ;
        RECT 2695.520 1673.960 2734.160 1674.440 ;
        RECT 2695.520 1668.520 2734.160 1669.000 ;
        RECT 2695.520 1663.080 2734.160 1663.560 ;
        RECT 2695.520 1657.640 2734.160 1658.120 ;
        RECT 2695.520 1652.200 2734.160 1652.680 ;
        RECT 2695.520 1646.760 2734.160 1647.240 ;
        RECT 2695.520 1641.320 2734.160 1641.800 ;
        RECT 2695.520 1635.880 2734.160 1636.360 ;
        RECT 2695.520 1630.440 2734.160 1630.920 ;
        RECT 2884.970 1628.665 2888.070 1629.785 ;
        RECT 2882.000 1628.510 2888.235 1628.665 ;
        RECT 2881.580 1628.340 2888.235 1628.510 ;
        RECT 2882.000 1628.185 2888.235 1628.340 ;
        RECT 2524.970 1626.555 2528.070 1627.675 ;
        RECT 2522.555 1626.400 2528.245 1626.555 ;
        RECT 2522.135 1626.230 2528.245 1626.400 ;
        RECT 2522.555 1626.075 2528.245 1626.230 ;
        RECT 2695.520 1625.000 2734.160 1625.480 ;
        RECT 2524.970 1620.140 2528.070 1621.260 ;
        RECT 2522.555 1619.985 2528.245 1620.140 ;
        RECT 2522.135 1619.815 2528.245 1619.985 ;
        RECT 2522.555 1619.660 2528.245 1619.815 ;
        RECT 2695.520 1619.560 2734.160 1620.040 ;
        RECT 2695.520 1614.120 2734.160 1614.600 ;
        RECT 2359.970 1609.145 2360.260 1609.175 ;
        RECT 2359.800 1608.975 2360.260 1609.145 ;
        RECT 2359.970 1608.945 2360.260 1608.975 ;
        RECT 2695.520 1608.680 2734.160 1609.160 ;
        RECT 2358.045 1607.025 2360.795 1607.035 ;
        RECT 2361.455 1607.025 2364.205 1607.035 ;
        RECT 2373.140 1607.030 2377.865 1607.035 ;
        RECT 2378.675 1607.030 2381.425 1607.035 ;
        RECT 2390.360 1607.030 2395.085 1607.035 ;
        RECT 2395.895 1607.030 2398.645 1607.040 ;
        RECT 2407.580 1607.035 2412.305 1607.040 ;
        RECT 2406.475 1607.030 2412.460 1607.035 ;
        RECT 2413.115 1607.030 2415.865 1607.035 ;
        RECT 2424.800 1607.030 2429.525 1607.035 ;
        RECT 2430.335 1607.030 2433.085 1607.035 ;
        RECT 2442.020 1607.030 2446.745 1607.035 ;
        RECT 2343.000 1607.000 2364.470 1607.025 ;
        RECT 2372.035 1607.005 2381.580 1607.030 ;
        RECT 2343.000 1606.800 2364.940 1607.000 ;
        RECT 2372.035 1606.955 2381.585 1607.005 ;
        RECT 2389.255 1606.955 2398.805 1607.030 ;
        RECT 2406.475 1606.960 2416.025 1607.030 ;
        RECT 2371.945 1606.800 2381.585 1606.955 ;
        RECT 2389.165 1606.805 2398.805 1606.955 ;
        RECT 2406.385 1606.805 2416.025 1606.960 ;
        RECT 2423.695 1606.955 2433.245 1607.030 ;
        RECT 2440.915 1606.955 2446.900 1607.030 ;
        RECT 2389.165 1606.800 2399.385 1606.805 ;
        RECT 2343.000 1605.965 2364.945 1606.800 ;
        RECT 2371.935 1605.965 2382.165 1606.800 ;
        RECT 2389.155 1605.970 2399.385 1606.800 ;
        RECT 2406.375 1606.800 2416.025 1606.805 ;
        RECT 2423.605 1606.800 2433.245 1606.955 ;
        RECT 2440.825 1606.800 2446.900 1606.955 ;
        RECT 2406.375 1605.970 2416.605 1606.800 ;
        RECT 2389.155 1605.965 2416.605 1605.970 ;
        RECT 2423.595 1605.965 2433.825 1606.800 ;
        RECT 2440.815 1605.965 2446.900 1606.800 ;
        RECT 2343.000 1605.490 2446.900 1605.965 ;
        RECT 2343.000 1605.485 2399.380 1605.490 ;
        RECT 2343.000 1605.425 2364.940 1605.485 ;
        RECT 2372.030 1605.430 2382.160 1605.485 ;
        RECT 2389.250 1605.430 2399.380 1605.485 ;
        RECT 2406.470 1605.485 2446.900 1605.490 ;
        RECT 2406.470 1605.435 2416.600 1605.485 ;
        RECT 2406.475 1605.430 2416.600 1605.435 ;
        RECT 2423.690 1605.430 2433.820 1605.485 ;
        RECT 2440.910 1605.430 2446.900 1605.485 ;
        RECT 2373.140 1605.425 2382.160 1605.430 ;
        RECT 2390.360 1605.425 2395.080 1605.430 ;
        RECT 2412.455 1605.425 2416.600 1605.430 ;
        RECT 2424.800 1605.425 2433.820 1605.430 ;
        RECT 2442.020 1605.425 2446.740 1605.430 ;
        RECT 2695.520 1603.240 2734.160 1603.720 ;
        RECT 2695.520 1597.800 2734.160 1598.280 ;
        RECT 2695.520 1592.360 2734.160 1592.840 ;
        RECT 2524.970 1590.895 2528.070 1592.015 ;
        RECT 2522.555 1590.740 2528.245 1590.895 ;
        RECT 2522.135 1590.570 2528.245 1590.740 ;
        RECT 2522.555 1590.415 2528.245 1590.570 ;
        RECT 2524.970 1583.365 2528.070 1584.485 ;
        RECT 2522.555 1583.210 2528.245 1583.365 ;
        RECT 2522.135 1583.040 2528.245 1583.210 ;
        RECT 2522.555 1582.885 2528.245 1583.040 ;
        RECT 2524.970 1577.385 2528.070 1578.505 ;
        RECT 2522.555 1577.230 2528.245 1577.385 ;
        RECT 2522.135 1577.060 2528.245 1577.230 ;
        RECT 2522.555 1576.905 2528.245 1577.060 ;
        RECT 2524.970 1568.970 2528.070 1570.090 ;
        RECT 2522.555 1568.815 2528.245 1568.970 ;
        RECT 2522.135 1568.645 2528.245 1568.815 ;
        RECT 2522.555 1568.490 2528.245 1568.645 ;
        RECT 2359.970 1532.145 2360.260 1532.175 ;
        RECT 2359.800 1531.975 2360.260 1532.145 ;
        RECT 2359.970 1531.945 2360.260 1531.975 ;
        RECT 2343.000 1528.435 2442.420 1530.035 ;
        RECT 2360.790 1528.430 2442.420 1528.435 ;
        RECT 2361.535 1528.285 2371.195 1528.430 ;
        RECT 2372.240 1528.425 2375.975 1528.430 ;
        RECT 2377.860 1528.285 2387.520 1528.430 ;
        RECT 2388.565 1528.425 2392.300 1528.430 ;
        RECT 2394.185 1528.285 2403.845 1528.430 ;
        RECT 2404.890 1528.425 2408.625 1528.430 ;
        RECT 2410.510 1528.285 2420.170 1528.430 ;
        RECT 2421.215 1528.425 2424.950 1528.430 ;
        RECT 2426.835 1528.285 2436.495 1528.430 ;
        RECT 2437.540 1528.425 2441.275 1528.430 ;
        RECT 2695.520 1493.960 2734.160 1494.440 ;
        RECT 2695.520 1488.520 2734.160 1489.000 ;
        RECT 2695.520 1483.080 2734.160 1483.560 ;
        RECT 2695.520 1477.640 2734.160 1478.120 ;
        RECT 2695.520 1472.200 2734.160 1472.680 ;
        RECT 2695.520 1466.760 2734.160 1467.240 ;
        RECT 2695.520 1461.320 2734.160 1461.800 ;
        RECT 2695.520 1455.880 2734.160 1456.360 ;
        RECT 2695.520 1450.440 2734.160 1450.920 ;
        RECT 2695.520 1445.000 2734.160 1445.480 ;
        RECT 2524.970 1439.270 2528.070 1440.390 ;
        RECT 2695.520 1439.560 2734.160 1440.040 ;
        RECT 2522.555 1439.115 2528.245 1439.270 ;
        RECT 2522.135 1438.945 2528.245 1439.115 ;
        RECT 2522.555 1438.790 2528.245 1438.945 ;
        RECT 2359.970 1434.150 2360.260 1434.180 ;
        RECT 2359.800 1433.980 2360.260 1434.150 ;
        RECT 2695.520 1434.120 2734.160 1434.600 ;
        RECT 2359.970 1433.950 2360.260 1433.980 ;
        RECT 2524.970 1432.855 2528.070 1433.975 ;
        RECT 2522.555 1432.700 2528.245 1432.855 ;
        RECT 2522.135 1432.530 2528.245 1432.700 ;
        RECT 2522.555 1432.375 2528.245 1432.530 ;
        RECT 2343.000 1432.035 2453.495 1432.040 ;
        RECT 2343.000 1430.440 2453.595 1432.035 ;
        RECT 2361.540 1430.430 2379.355 1430.440 ;
        RECT 2380.100 1430.430 2397.915 1430.440 ;
        RECT 2398.660 1430.430 2416.475 1430.440 ;
        RECT 2417.220 1430.430 2435.035 1430.440 ;
        RECT 2435.780 1430.430 2453.595 1430.440 ;
        RECT 2361.540 1430.395 2373.500 1430.430 ;
        RECT 2374.475 1430.425 2378.210 1430.430 ;
        RECT 2380.100 1430.395 2392.060 1430.430 ;
        RECT 2393.035 1430.425 2396.770 1430.430 ;
        RECT 2398.660 1430.395 2410.620 1430.430 ;
        RECT 2411.595 1430.425 2415.330 1430.430 ;
        RECT 2417.220 1430.395 2429.180 1430.430 ;
        RECT 2430.155 1430.425 2433.890 1430.430 ;
        RECT 2435.780 1430.395 2447.740 1430.430 ;
        RECT 2448.715 1430.425 2452.450 1430.430 ;
        RECT 2695.520 1428.680 2734.160 1429.160 ;
        RECT 2695.520 1423.240 2734.160 1423.720 ;
        RECT 2524.970 1418.665 2528.070 1419.785 ;
        RECT 2522.555 1418.510 2528.245 1418.665 ;
        RECT 2522.135 1418.340 2528.245 1418.510 ;
        RECT 2522.555 1418.185 2528.245 1418.340 ;
        RECT 2695.520 1417.800 2734.160 1418.280 ;
        RECT 2695.520 1412.360 2734.160 1412.840 ;
        RECT 2524.970 1411.135 2528.070 1412.255 ;
        RECT 2522.555 1410.980 2528.245 1411.135 ;
        RECT 2522.135 1410.810 2528.245 1410.980 ;
        RECT 2522.555 1410.655 2528.245 1410.810 ;
        RECT 2524.970 1405.155 2528.070 1406.275 ;
        RECT 2522.555 1405.000 2528.245 1405.155 ;
        RECT 2522.135 1404.830 2528.245 1405.000 ;
        RECT 2522.555 1404.675 2528.245 1404.830 ;
        RECT 2524.970 1396.740 2528.070 1397.860 ;
        RECT 2522.555 1396.585 2528.245 1396.740 ;
        RECT 2522.135 1396.415 2528.245 1396.585 ;
        RECT 2522.555 1396.260 2528.245 1396.415 ;
        RECT 2884.970 1363.465 2888.070 1364.585 ;
        RECT 2882.000 1363.310 2888.235 1363.465 ;
        RECT 2881.580 1363.140 2888.235 1363.310 ;
        RECT 2882.000 1362.985 2888.235 1363.140 ;
        RECT 2369.970 1334.150 2370.260 1334.180 ;
        RECT 2369.800 1333.980 2370.260 1334.150 ;
        RECT 2369.970 1333.950 2370.260 1333.980 ;
        RECT 2368.045 1332.035 2370.795 1332.040 ;
        RECT 2375.560 1332.035 2378.310 1332.040 ;
        RECT 2381.175 1332.035 2385.900 1332.040 ;
        RECT 2390.820 1332.035 2393.570 1332.040 ;
        RECT 2396.435 1332.035 2401.160 1332.040 ;
        RECT 2406.080 1332.035 2408.830 1332.040 ;
        RECT 2411.695 1332.035 2416.420 1332.040 ;
        RECT 2421.340 1332.035 2424.090 1332.040 ;
        RECT 2426.955 1332.035 2431.680 1332.040 ;
        RECT 2436.600 1332.035 2439.350 1332.040 ;
        RECT 2442.215 1332.035 2446.940 1332.040 ;
        RECT 2343.000 1330.435 2447.095 1332.035 ;
        RECT 2371.545 1330.430 2386.055 1330.435 ;
        RECT 2386.805 1330.430 2401.315 1330.435 ;
        RECT 2402.065 1330.430 2416.575 1330.435 ;
        RECT 2417.325 1330.430 2431.835 1330.435 ;
        RECT 2432.585 1330.430 2447.095 1330.435 ;
        RECT 2371.545 1330.395 2380.285 1330.430 ;
        RECT 2381.175 1330.425 2385.895 1330.430 ;
        RECT 2386.805 1330.395 2395.545 1330.430 ;
        RECT 2396.435 1330.425 2401.155 1330.430 ;
        RECT 2402.065 1330.395 2410.805 1330.430 ;
        RECT 2411.695 1330.425 2416.415 1330.430 ;
        RECT 2417.325 1330.395 2426.065 1330.430 ;
        RECT 2426.955 1330.425 2431.675 1330.430 ;
        RECT 2432.585 1330.395 2441.325 1330.430 ;
        RECT 2442.215 1330.425 2446.935 1330.430 ;
        RECT 2884.970 1164.225 2888.070 1165.345 ;
        RECT 2882.000 1164.070 2888.235 1164.225 ;
        RECT 2881.580 1163.900 2888.235 1164.070 ;
        RECT 2882.000 1163.745 2888.235 1163.900 ;
      LAYER met2 ;
        RECT 1265.110 3508.275 1267.930 3509.875 ;
        RECT 1625.110 3508.725 1627.930 3510.325 ;
        RECT 1805.110 3506.805 1807.930 3508.405 ;
        RECT 2165.110 3506.445 2167.930 3508.045 ;
        RECT 2525.110 3507.130 2527.930 3508.730 ;
        RECT 2885.110 3487.985 2887.930 3489.585 ;
        RECT 2885.110 3222.105 2887.930 3223.705 ;
        RECT 2885.110 2956.905 2887.930 2958.505 ;
        RECT 2885.110 2691.025 2887.930 2692.625 ;
        RECT 2885.110 2425.145 2887.930 2426.745 ;
        RECT 2345.110 2250.425 2347.930 2252.025 ;
        RECT 2699.580 2214.015 2701.120 2214.385 ;
        RECT 2709.240 2214.015 2710.780 2214.385 ;
        RECT 2718.900 2214.015 2720.440 2214.385 ;
        RECT 2728.560 2214.015 2730.100 2214.385 ;
        RECT 2699.580 2208.575 2701.120 2208.945 ;
        RECT 2709.240 2208.575 2710.780 2208.945 ;
        RECT 2718.900 2208.575 2720.440 2208.945 ;
        RECT 2728.560 2208.575 2730.100 2208.945 ;
        RECT 2699.580 2203.135 2701.120 2203.505 ;
        RECT 2709.240 2203.135 2710.780 2203.505 ;
        RECT 2718.900 2203.135 2720.440 2203.505 ;
        RECT 2728.560 2203.135 2730.100 2203.505 ;
        RECT 2699.580 2197.695 2701.120 2198.065 ;
        RECT 2709.240 2197.695 2710.780 2198.065 ;
        RECT 2718.900 2197.695 2720.440 2198.065 ;
        RECT 2728.560 2197.695 2730.100 2198.065 ;
        RECT 2699.580 2192.255 2701.120 2192.625 ;
        RECT 2709.240 2192.255 2710.780 2192.625 ;
        RECT 2718.900 2192.255 2720.440 2192.625 ;
        RECT 2728.560 2192.255 2730.100 2192.625 ;
        RECT 2699.580 2186.815 2701.120 2187.185 ;
        RECT 2709.240 2186.815 2710.780 2187.185 ;
        RECT 2718.900 2186.815 2720.440 2187.185 ;
        RECT 2728.560 2186.815 2730.100 2187.185 ;
        RECT 2699.580 2181.375 2701.120 2181.745 ;
        RECT 2709.240 2181.375 2710.780 2181.745 ;
        RECT 2718.900 2181.375 2720.440 2181.745 ;
        RECT 2728.560 2181.375 2730.100 2181.745 ;
        RECT 2699.580 2175.935 2701.120 2176.305 ;
        RECT 2709.240 2175.935 2710.780 2176.305 ;
        RECT 2718.900 2175.935 2720.440 2176.305 ;
        RECT 2728.560 2175.935 2730.100 2176.305 ;
        RECT 2699.580 2170.495 2701.120 2170.865 ;
        RECT 2709.240 2170.495 2710.780 2170.865 ;
        RECT 2718.900 2170.495 2720.440 2170.865 ;
        RECT 2728.560 2170.495 2730.100 2170.865 ;
        RECT 2699.580 2165.055 2701.120 2165.425 ;
        RECT 2709.240 2165.055 2710.780 2165.425 ;
        RECT 2718.900 2165.055 2720.440 2165.425 ;
        RECT 2728.560 2165.055 2730.100 2165.425 ;
        RECT 2345.110 2158.425 2347.930 2160.025 ;
        RECT 2699.580 2159.615 2701.120 2159.985 ;
        RECT 2709.240 2159.615 2710.780 2159.985 ;
        RECT 2718.900 2159.615 2720.440 2159.985 ;
        RECT 2728.560 2159.615 2730.100 2159.985 ;
        RECT 2885.110 2159.945 2887.930 2161.545 ;
        RECT 2699.580 2154.175 2701.120 2154.545 ;
        RECT 2709.240 2154.175 2710.780 2154.545 ;
        RECT 2718.900 2154.175 2720.440 2154.545 ;
        RECT 2728.560 2154.175 2730.100 2154.545 ;
        RECT 2699.580 2148.735 2701.120 2149.105 ;
        RECT 2709.240 2148.735 2710.780 2149.105 ;
        RECT 2718.900 2148.735 2720.440 2149.105 ;
        RECT 2728.560 2148.735 2730.100 2149.105 ;
        RECT 2699.580 2143.295 2701.120 2143.665 ;
        RECT 2709.240 2143.295 2710.780 2143.665 ;
        RECT 2718.900 2143.295 2720.440 2143.665 ;
        RECT 2728.560 2143.295 2730.100 2143.665 ;
        RECT 2525.110 2136.435 2527.930 2138.035 ;
        RECT 2699.580 2137.855 2701.120 2138.225 ;
        RECT 2709.240 2137.855 2710.780 2138.225 ;
        RECT 2718.900 2137.855 2720.440 2138.225 ;
        RECT 2728.560 2137.855 2730.100 2138.225 ;
        RECT 2699.580 2132.415 2701.120 2132.785 ;
        RECT 2709.240 2132.415 2710.780 2132.785 ;
        RECT 2718.900 2132.415 2720.440 2132.785 ;
        RECT 2728.560 2132.415 2730.100 2132.785 ;
        RECT 2525.110 2128.905 2527.930 2130.505 ;
        RECT 2525.110 2122.925 2527.930 2124.525 ;
        RECT 2525.110 2116.980 2527.930 2118.580 ;
        RECT 2525.110 2111.335 2527.930 2112.935 ;
        RECT 2525.110 2105.330 2527.930 2106.930 ;
        RECT 2345.110 2053.430 2347.930 2055.030 ;
        RECT 2699.580 2034.015 2701.120 2034.385 ;
        RECT 2709.240 2034.015 2710.780 2034.385 ;
        RECT 2718.900 2034.015 2720.440 2034.385 ;
        RECT 2728.560 2034.015 2730.100 2034.385 ;
        RECT 2699.580 2028.575 2701.120 2028.945 ;
        RECT 2709.240 2028.575 2710.780 2028.945 ;
        RECT 2718.900 2028.575 2720.440 2028.945 ;
        RECT 2728.560 2028.575 2730.100 2028.945 ;
        RECT 2699.580 2023.135 2701.120 2023.505 ;
        RECT 2709.240 2023.135 2710.780 2023.505 ;
        RECT 2718.900 2023.135 2720.440 2023.505 ;
        RECT 2728.560 2023.135 2730.100 2023.505 ;
        RECT 2699.580 2017.695 2701.120 2018.065 ;
        RECT 2709.240 2017.695 2710.780 2018.065 ;
        RECT 2718.900 2017.695 2720.440 2018.065 ;
        RECT 2728.560 2017.695 2730.100 2018.065 ;
        RECT 2699.580 2012.255 2701.120 2012.625 ;
        RECT 2709.240 2012.255 2710.780 2012.625 ;
        RECT 2718.900 2012.255 2720.440 2012.625 ;
        RECT 2728.560 2012.255 2730.100 2012.625 ;
        RECT 2699.580 2006.815 2701.120 2007.185 ;
        RECT 2709.240 2006.815 2710.780 2007.185 ;
        RECT 2718.900 2006.815 2720.440 2007.185 ;
        RECT 2728.560 2006.815 2730.100 2007.185 ;
        RECT 2699.580 2001.375 2701.120 2001.745 ;
        RECT 2709.240 2001.375 2710.780 2001.745 ;
        RECT 2718.900 2001.375 2720.440 2001.745 ;
        RECT 2728.560 2001.375 2730.100 2001.745 ;
        RECT 2699.580 1995.935 2701.120 1996.305 ;
        RECT 2709.240 1995.935 2710.780 1996.305 ;
        RECT 2718.900 1995.935 2720.440 1996.305 ;
        RECT 2728.560 1995.935 2730.100 1996.305 ;
        RECT 2699.580 1990.495 2701.120 1990.865 ;
        RECT 2709.240 1990.495 2710.780 1990.865 ;
        RECT 2718.900 1990.495 2720.440 1990.865 ;
        RECT 2728.560 1990.495 2730.100 1990.865 ;
        RECT 2525.110 1984.180 2527.930 1985.780 ;
        RECT 2699.580 1985.055 2701.120 1985.425 ;
        RECT 2709.240 1985.055 2710.780 1985.425 ;
        RECT 2718.900 1985.055 2720.440 1985.425 ;
        RECT 2728.560 1985.055 2730.100 1985.425 ;
        RECT 2699.580 1979.615 2701.120 1979.985 ;
        RECT 2709.240 1979.615 2710.780 1979.985 ;
        RECT 2718.900 1979.615 2720.440 1979.985 ;
        RECT 2728.560 1979.615 2730.100 1979.985 ;
        RECT 2525.110 1976.650 2527.930 1978.250 ;
        RECT 2699.580 1974.175 2701.120 1974.545 ;
        RECT 2709.240 1974.175 2710.780 1974.545 ;
        RECT 2718.900 1974.175 2720.440 1974.545 ;
        RECT 2728.560 1974.175 2730.100 1974.545 ;
        RECT 2525.110 1970.670 2527.930 1972.270 ;
        RECT 2699.580 1968.735 2701.120 1969.105 ;
        RECT 2709.240 1968.735 2710.780 1969.105 ;
        RECT 2718.900 1968.735 2720.440 1969.105 ;
        RECT 2728.560 1968.735 2730.100 1969.105 ;
        RECT 2525.110 1964.725 2527.930 1966.325 ;
        RECT 2699.580 1963.295 2701.120 1963.665 ;
        RECT 2709.240 1963.295 2710.780 1963.665 ;
        RECT 2718.900 1963.295 2720.440 1963.665 ;
        RECT 2728.560 1963.295 2730.100 1963.665 ;
        RECT 2525.110 1959.080 2527.930 1960.680 ;
        RECT 2699.580 1957.855 2701.120 1958.225 ;
        RECT 2709.240 1957.855 2710.780 1958.225 ;
        RECT 2718.900 1957.855 2720.440 1958.225 ;
        RECT 2728.560 1957.855 2730.100 1958.225 ;
        RECT 2525.110 1953.075 2527.930 1954.675 ;
        RECT 2699.580 1952.415 2701.120 1952.785 ;
        RECT 2709.240 1952.415 2710.780 1952.785 ;
        RECT 2718.900 1952.415 2720.440 1952.785 ;
        RECT 2728.560 1952.415 2730.100 1952.785 ;
        RECT 2345.110 1948.450 2347.930 1950.050 ;
        RECT 2885.110 1894.065 2887.930 1895.665 ;
        RECT 2699.580 1854.015 2701.120 1854.385 ;
        RECT 2709.240 1854.015 2710.780 1854.385 ;
        RECT 2718.900 1854.015 2720.440 1854.385 ;
        RECT 2728.560 1854.015 2730.100 1854.385 ;
        RECT 2699.580 1848.575 2701.120 1848.945 ;
        RECT 2709.240 1848.575 2710.780 1848.945 ;
        RECT 2718.900 1848.575 2720.440 1848.945 ;
        RECT 2728.560 1848.575 2730.100 1848.945 ;
        RECT 2699.580 1843.135 2701.120 1843.505 ;
        RECT 2709.240 1843.135 2710.780 1843.505 ;
        RECT 2718.900 1843.135 2720.440 1843.505 ;
        RECT 2728.560 1843.135 2730.100 1843.505 ;
        RECT 2699.580 1837.695 2701.120 1838.065 ;
        RECT 2709.240 1837.695 2710.780 1838.065 ;
        RECT 2718.900 1837.695 2720.440 1838.065 ;
        RECT 2728.560 1837.695 2730.100 1838.065 ;
        RECT 2699.580 1832.255 2701.120 1832.625 ;
        RECT 2709.240 1832.255 2710.780 1832.625 ;
        RECT 2718.900 1832.255 2720.440 1832.625 ;
        RECT 2728.560 1832.255 2730.100 1832.625 ;
        RECT 2699.580 1826.815 2701.120 1827.185 ;
        RECT 2709.240 1826.815 2710.780 1827.185 ;
        RECT 2718.900 1826.815 2720.440 1827.185 ;
        RECT 2728.560 1826.815 2730.100 1827.185 ;
        RECT 2699.580 1821.375 2701.120 1821.745 ;
        RECT 2709.240 1821.375 2710.780 1821.745 ;
        RECT 2718.900 1821.375 2720.440 1821.745 ;
        RECT 2728.560 1821.375 2730.100 1821.745 ;
        RECT 2699.580 1815.935 2701.120 1816.305 ;
        RECT 2709.240 1815.935 2710.780 1816.305 ;
        RECT 2718.900 1815.935 2720.440 1816.305 ;
        RECT 2728.560 1815.935 2730.100 1816.305 ;
        RECT 2699.580 1810.495 2701.120 1810.865 ;
        RECT 2709.240 1810.495 2710.780 1810.865 ;
        RECT 2718.900 1810.495 2720.440 1810.865 ;
        RECT 2728.560 1810.495 2730.100 1810.865 ;
        RECT 2525.110 1807.210 2527.930 1808.810 ;
        RECT 2699.580 1805.055 2701.120 1805.425 ;
        RECT 2709.240 1805.055 2710.780 1805.425 ;
        RECT 2718.900 1805.055 2720.440 1805.425 ;
        RECT 2728.560 1805.055 2730.100 1805.425 ;
        RECT 2525.110 1799.680 2527.930 1801.280 ;
        RECT 2699.580 1799.615 2701.120 1799.985 ;
        RECT 2709.240 1799.615 2710.780 1799.985 ;
        RECT 2718.900 1799.615 2720.440 1799.985 ;
        RECT 2728.560 1799.615 2730.100 1799.985 ;
        RECT 2525.110 1793.700 2527.930 1795.300 ;
        RECT 2699.580 1794.175 2701.120 1794.545 ;
        RECT 2709.240 1794.175 2710.780 1794.545 ;
        RECT 2718.900 1794.175 2720.440 1794.545 ;
        RECT 2728.560 1794.175 2730.100 1794.545 ;
        RECT 2525.110 1787.755 2527.930 1789.355 ;
        RECT 2699.580 1788.735 2701.120 1789.105 ;
        RECT 2709.240 1788.735 2710.780 1789.105 ;
        RECT 2718.900 1788.735 2720.440 1789.105 ;
        RECT 2728.560 1788.735 2730.100 1789.105 ;
        RECT 2345.110 1785.435 2347.930 1787.035 ;
        RECT 2525.110 1782.110 2527.930 1783.710 ;
        RECT 2699.580 1783.295 2701.120 1783.665 ;
        RECT 2709.240 1783.295 2710.780 1783.665 ;
        RECT 2718.900 1783.295 2720.440 1783.665 ;
        RECT 2728.560 1783.295 2730.100 1783.665 ;
        RECT 2699.580 1777.855 2701.120 1778.225 ;
        RECT 2709.240 1777.855 2710.780 1778.225 ;
        RECT 2718.900 1777.855 2720.440 1778.225 ;
        RECT 2728.560 1777.855 2730.100 1778.225 ;
        RECT 2699.580 1772.415 2701.120 1772.785 ;
        RECT 2709.240 1772.415 2710.780 1772.785 ;
        RECT 2718.900 1772.415 2720.440 1772.785 ;
        RECT 2728.560 1772.415 2730.100 1772.785 ;
        RECT 2525.110 1770.640 2527.930 1772.240 ;
        RECT 2345.110 1705.425 2347.930 1707.025 ;
        RECT 2699.580 1674.015 2701.120 1674.385 ;
        RECT 2709.240 1674.015 2710.780 1674.385 ;
        RECT 2718.900 1674.015 2720.440 1674.385 ;
        RECT 2728.560 1674.015 2730.100 1674.385 ;
        RECT 2699.580 1668.575 2701.120 1668.945 ;
        RECT 2709.240 1668.575 2710.780 1668.945 ;
        RECT 2718.900 1668.575 2720.440 1668.945 ;
        RECT 2728.560 1668.575 2730.100 1668.945 ;
        RECT 2699.580 1663.135 2701.120 1663.505 ;
        RECT 2709.240 1663.135 2710.780 1663.505 ;
        RECT 2718.900 1663.135 2720.440 1663.505 ;
        RECT 2728.560 1663.135 2730.100 1663.505 ;
        RECT 2699.580 1657.695 2701.120 1658.065 ;
        RECT 2709.240 1657.695 2710.780 1658.065 ;
        RECT 2718.900 1657.695 2720.440 1658.065 ;
        RECT 2728.560 1657.695 2730.100 1658.065 ;
        RECT 2699.580 1652.255 2701.120 1652.625 ;
        RECT 2709.240 1652.255 2710.780 1652.625 ;
        RECT 2718.900 1652.255 2720.440 1652.625 ;
        RECT 2728.560 1652.255 2730.100 1652.625 ;
        RECT 2699.580 1646.815 2701.120 1647.185 ;
        RECT 2709.240 1646.815 2710.780 1647.185 ;
        RECT 2718.900 1646.815 2720.440 1647.185 ;
        RECT 2728.560 1646.815 2730.100 1647.185 ;
        RECT 2699.580 1641.375 2701.120 1641.745 ;
        RECT 2709.240 1641.375 2710.780 1641.745 ;
        RECT 2718.900 1641.375 2720.440 1641.745 ;
        RECT 2728.560 1641.375 2730.100 1641.745 ;
        RECT 2699.580 1635.935 2701.120 1636.305 ;
        RECT 2709.240 1635.935 2710.780 1636.305 ;
        RECT 2718.900 1635.935 2720.440 1636.305 ;
        RECT 2728.560 1635.935 2730.100 1636.305 ;
        RECT 2699.580 1630.495 2701.120 1630.865 ;
        RECT 2709.240 1630.495 2710.780 1630.865 ;
        RECT 2718.900 1630.495 2720.440 1630.865 ;
        RECT 2728.560 1630.495 2730.100 1630.865 ;
        RECT 2885.110 1628.185 2887.930 1629.785 ;
        RECT 2525.110 1626.075 2527.930 1627.675 ;
        RECT 2699.580 1625.055 2701.120 1625.425 ;
        RECT 2709.240 1625.055 2710.780 1625.425 ;
        RECT 2718.900 1625.055 2720.440 1625.425 ;
        RECT 2728.560 1625.055 2730.100 1625.425 ;
        RECT 2525.110 1619.660 2527.930 1621.260 ;
        RECT 2699.580 1619.615 2701.120 1619.985 ;
        RECT 2709.240 1619.615 2710.780 1619.985 ;
        RECT 2718.900 1619.615 2720.440 1619.985 ;
        RECT 2728.560 1619.615 2730.100 1619.985 ;
        RECT 2699.580 1614.175 2701.120 1614.545 ;
        RECT 2709.240 1614.175 2710.780 1614.545 ;
        RECT 2718.900 1614.175 2720.440 1614.545 ;
        RECT 2728.560 1614.175 2730.100 1614.545 ;
        RECT 2699.580 1608.735 2701.120 1609.105 ;
        RECT 2709.240 1608.735 2710.780 1609.105 ;
        RECT 2718.900 1608.735 2720.440 1609.105 ;
        RECT 2728.560 1608.735 2730.100 1609.105 ;
        RECT 2345.110 1605.425 2347.930 1607.025 ;
        RECT 2699.580 1603.295 2701.120 1603.665 ;
        RECT 2709.240 1603.295 2710.780 1603.665 ;
        RECT 2718.900 1603.295 2720.440 1603.665 ;
        RECT 2728.560 1603.295 2730.100 1603.665 ;
        RECT 2699.580 1597.855 2701.120 1598.225 ;
        RECT 2709.240 1597.855 2710.780 1598.225 ;
        RECT 2718.900 1597.855 2720.440 1598.225 ;
        RECT 2728.560 1597.855 2730.100 1598.225 ;
        RECT 2699.580 1592.415 2701.120 1592.785 ;
        RECT 2709.240 1592.415 2710.780 1592.785 ;
        RECT 2718.900 1592.415 2720.440 1592.785 ;
        RECT 2728.560 1592.415 2730.100 1592.785 ;
        RECT 2525.110 1590.415 2527.930 1592.015 ;
        RECT 2525.110 1582.885 2527.930 1584.485 ;
        RECT 2525.110 1576.905 2527.930 1578.505 ;
        RECT 2525.110 1568.490 2527.930 1570.090 ;
        RECT 2345.110 1528.435 2347.930 1530.035 ;
        RECT 2699.580 1494.015 2701.120 1494.385 ;
        RECT 2709.240 1494.015 2710.780 1494.385 ;
        RECT 2718.900 1494.015 2720.440 1494.385 ;
        RECT 2728.560 1494.015 2730.100 1494.385 ;
        RECT 2699.580 1488.575 2701.120 1488.945 ;
        RECT 2709.240 1488.575 2710.780 1488.945 ;
        RECT 2718.900 1488.575 2720.440 1488.945 ;
        RECT 2728.560 1488.575 2730.100 1488.945 ;
        RECT 2699.580 1483.135 2701.120 1483.505 ;
        RECT 2709.240 1483.135 2710.780 1483.505 ;
        RECT 2718.900 1483.135 2720.440 1483.505 ;
        RECT 2728.560 1483.135 2730.100 1483.505 ;
        RECT 2699.580 1477.695 2701.120 1478.065 ;
        RECT 2709.240 1477.695 2710.780 1478.065 ;
        RECT 2718.900 1477.695 2720.440 1478.065 ;
        RECT 2728.560 1477.695 2730.100 1478.065 ;
        RECT 2699.580 1472.255 2701.120 1472.625 ;
        RECT 2709.240 1472.255 2710.780 1472.625 ;
        RECT 2718.900 1472.255 2720.440 1472.625 ;
        RECT 2728.560 1472.255 2730.100 1472.625 ;
        RECT 2699.580 1466.815 2701.120 1467.185 ;
        RECT 2709.240 1466.815 2710.780 1467.185 ;
        RECT 2718.900 1466.815 2720.440 1467.185 ;
        RECT 2728.560 1466.815 2730.100 1467.185 ;
        RECT 2699.580 1461.375 2701.120 1461.745 ;
        RECT 2709.240 1461.375 2710.780 1461.745 ;
        RECT 2718.900 1461.375 2720.440 1461.745 ;
        RECT 2728.560 1461.375 2730.100 1461.745 ;
        RECT 2699.580 1455.935 2701.120 1456.305 ;
        RECT 2709.240 1455.935 2710.780 1456.305 ;
        RECT 2718.900 1455.935 2720.440 1456.305 ;
        RECT 2728.560 1455.935 2730.100 1456.305 ;
        RECT 2699.580 1450.495 2701.120 1450.865 ;
        RECT 2709.240 1450.495 2710.780 1450.865 ;
        RECT 2718.900 1450.495 2720.440 1450.865 ;
        RECT 2728.560 1450.495 2730.100 1450.865 ;
        RECT 2699.580 1445.055 2701.120 1445.425 ;
        RECT 2709.240 1445.055 2710.780 1445.425 ;
        RECT 2718.900 1445.055 2720.440 1445.425 ;
        RECT 2728.560 1445.055 2730.100 1445.425 ;
        RECT 2525.110 1438.790 2527.930 1440.390 ;
        RECT 2699.580 1439.615 2701.120 1439.985 ;
        RECT 2709.240 1439.615 2710.780 1439.985 ;
        RECT 2718.900 1439.615 2720.440 1439.985 ;
        RECT 2728.560 1439.615 2730.100 1439.985 ;
        RECT 2699.580 1434.175 2701.120 1434.545 ;
        RECT 2709.240 1434.175 2710.780 1434.545 ;
        RECT 2718.900 1434.175 2720.440 1434.545 ;
        RECT 2728.560 1434.175 2730.100 1434.545 ;
        RECT 2525.110 1432.375 2527.930 1433.975 ;
        RECT 2345.110 1430.440 2347.930 1432.040 ;
        RECT 2699.580 1428.735 2701.120 1429.105 ;
        RECT 2709.240 1428.735 2710.780 1429.105 ;
        RECT 2718.900 1428.735 2720.440 1429.105 ;
        RECT 2728.560 1428.735 2730.100 1429.105 ;
        RECT 2699.580 1423.295 2701.120 1423.665 ;
        RECT 2709.240 1423.295 2710.780 1423.665 ;
        RECT 2718.900 1423.295 2720.440 1423.665 ;
        RECT 2728.560 1423.295 2730.100 1423.665 ;
        RECT 2525.110 1418.185 2527.930 1419.785 ;
        RECT 2699.580 1417.855 2701.120 1418.225 ;
        RECT 2709.240 1417.855 2710.780 1418.225 ;
        RECT 2718.900 1417.855 2720.440 1418.225 ;
        RECT 2728.560 1417.855 2730.100 1418.225 ;
        RECT 2699.580 1412.415 2701.120 1412.785 ;
        RECT 2709.240 1412.415 2710.780 1412.785 ;
        RECT 2718.900 1412.415 2720.440 1412.785 ;
        RECT 2728.560 1412.415 2730.100 1412.785 ;
        RECT 2525.110 1410.655 2527.930 1412.255 ;
        RECT 2525.110 1404.675 2527.930 1406.275 ;
        RECT 2525.110 1396.260 2527.930 1397.860 ;
        RECT 2885.110 1362.985 2887.930 1364.585 ;
        RECT 2345.110 1330.435 2347.930 1332.035 ;
        RECT 2885.110 1163.745 2887.930 1165.345 ;
      LAYER met3 ;
        RECT 1265.130 3508.310 1267.910 3509.840 ;
        RECT 1625.130 3508.760 1627.910 3510.290 ;
        RECT 1805.130 3506.840 1807.910 3508.370 ;
        RECT 2165.130 3506.480 2167.910 3508.010 ;
        RECT 2525.130 3507.165 2527.910 3508.695 ;
        RECT 2885.130 3488.020 2887.910 3489.550 ;
        RECT 2885.130 3222.140 2887.910 3223.670 ;
        RECT 2885.130 2956.940 2887.910 2958.470 ;
        RECT 2885.130 2691.060 2887.910 2692.590 ;
        RECT 2885.130 2425.180 2887.910 2426.710 ;
        RECT 2345.130 2250.460 2347.910 2251.990 ;
        RECT 2699.560 2214.035 2701.140 2214.365 ;
        RECT 2709.220 2214.035 2710.800 2214.365 ;
        RECT 2718.880 2214.035 2720.460 2214.365 ;
        RECT 2728.540 2214.035 2730.120 2214.365 ;
        RECT 2699.560 2208.595 2701.140 2208.925 ;
        RECT 2709.220 2208.595 2710.800 2208.925 ;
        RECT 2718.880 2208.595 2720.460 2208.925 ;
        RECT 2728.540 2208.595 2730.120 2208.925 ;
        RECT 2699.560 2203.155 2701.140 2203.485 ;
        RECT 2709.220 2203.155 2710.800 2203.485 ;
        RECT 2718.880 2203.155 2720.460 2203.485 ;
        RECT 2728.540 2203.155 2730.120 2203.485 ;
        RECT 2699.560 2197.715 2701.140 2198.045 ;
        RECT 2709.220 2197.715 2710.800 2198.045 ;
        RECT 2718.880 2197.715 2720.460 2198.045 ;
        RECT 2728.540 2197.715 2730.120 2198.045 ;
        RECT 2699.560 2192.275 2701.140 2192.605 ;
        RECT 2709.220 2192.275 2710.800 2192.605 ;
        RECT 2718.880 2192.275 2720.460 2192.605 ;
        RECT 2728.540 2192.275 2730.120 2192.605 ;
        RECT 2699.560 2186.835 2701.140 2187.165 ;
        RECT 2709.220 2186.835 2710.800 2187.165 ;
        RECT 2718.880 2186.835 2720.460 2187.165 ;
        RECT 2728.540 2186.835 2730.120 2187.165 ;
        RECT 2699.560 2181.395 2701.140 2181.725 ;
        RECT 2709.220 2181.395 2710.800 2181.725 ;
        RECT 2718.880 2181.395 2720.460 2181.725 ;
        RECT 2728.540 2181.395 2730.120 2181.725 ;
        RECT 2699.560 2175.955 2701.140 2176.285 ;
        RECT 2709.220 2175.955 2710.800 2176.285 ;
        RECT 2718.880 2175.955 2720.460 2176.285 ;
        RECT 2728.540 2175.955 2730.120 2176.285 ;
        RECT 2699.560 2170.515 2701.140 2170.845 ;
        RECT 2709.220 2170.515 2710.800 2170.845 ;
        RECT 2718.880 2170.515 2720.460 2170.845 ;
        RECT 2728.540 2170.515 2730.120 2170.845 ;
        RECT 2699.560 2165.075 2701.140 2165.405 ;
        RECT 2709.220 2165.075 2710.800 2165.405 ;
        RECT 2718.880 2165.075 2720.460 2165.405 ;
        RECT 2728.540 2165.075 2730.120 2165.405 ;
        RECT 2345.130 2158.460 2347.910 2159.990 ;
        RECT 2885.130 2159.980 2887.910 2161.510 ;
        RECT 2699.560 2159.635 2701.140 2159.965 ;
        RECT 2709.220 2159.635 2710.800 2159.965 ;
        RECT 2718.880 2159.635 2720.460 2159.965 ;
        RECT 2728.540 2159.635 2730.120 2159.965 ;
        RECT 2699.560 2154.195 2701.140 2154.525 ;
        RECT 2709.220 2154.195 2710.800 2154.525 ;
        RECT 2718.880 2154.195 2720.460 2154.525 ;
        RECT 2728.540 2154.195 2730.120 2154.525 ;
        RECT 2699.560 2148.755 2701.140 2149.085 ;
        RECT 2709.220 2148.755 2710.800 2149.085 ;
        RECT 2718.880 2148.755 2720.460 2149.085 ;
        RECT 2728.540 2148.755 2730.120 2149.085 ;
        RECT 2699.560 2143.315 2701.140 2143.645 ;
        RECT 2709.220 2143.315 2710.800 2143.645 ;
        RECT 2718.880 2143.315 2720.460 2143.645 ;
        RECT 2728.540 2143.315 2730.120 2143.645 ;
        RECT 2525.130 2136.470 2527.910 2138.000 ;
        RECT 2699.560 2137.875 2701.140 2138.205 ;
        RECT 2709.220 2137.875 2710.800 2138.205 ;
        RECT 2718.880 2137.875 2720.460 2138.205 ;
        RECT 2728.540 2137.875 2730.120 2138.205 ;
        RECT 2699.560 2132.435 2701.140 2132.765 ;
        RECT 2709.220 2132.435 2710.800 2132.765 ;
        RECT 2718.880 2132.435 2720.460 2132.765 ;
        RECT 2728.540 2132.435 2730.120 2132.765 ;
        RECT 2525.130 2128.940 2527.910 2130.470 ;
        RECT 2525.130 2122.960 2527.910 2124.490 ;
        RECT 2525.130 2117.015 2527.910 2118.545 ;
        RECT 2525.130 2111.370 2527.910 2112.900 ;
        RECT 2525.130 2105.365 2527.910 2106.895 ;
        RECT 2345.130 2053.465 2347.910 2054.995 ;
        RECT 2699.560 2034.035 2701.140 2034.365 ;
        RECT 2709.220 2034.035 2710.800 2034.365 ;
        RECT 2718.880 2034.035 2720.460 2034.365 ;
        RECT 2728.540 2034.035 2730.120 2034.365 ;
        RECT 2699.560 2028.595 2701.140 2028.925 ;
        RECT 2709.220 2028.595 2710.800 2028.925 ;
        RECT 2718.880 2028.595 2720.460 2028.925 ;
        RECT 2728.540 2028.595 2730.120 2028.925 ;
        RECT 2699.560 2023.155 2701.140 2023.485 ;
        RECT 2709.220 2023.155 2710.800 2023.485 ;
        RECT 2718.880 2023.155 2720.460 2023.485 ;
        RECT 2728.540 2023.155 2730.120 2023.485 ;
        RECT 2699.560 2017.715 2701.140 2018.045 ;
        RECT 2709.220 2017.715 2710.800 2018.045 ;
        RECT 2718.880 2017.715 2720.460 2018.045 ;
        RECT 2728.540 2017.715 2730.120 2018.045 ;
        RECT 2699.560 2012.275 2701.140 2012.605 ;
        RECT 2709.220 2012.275 2710.800 2012.605 ;
        RECT 2718.880 2012.275 2720.460 2012.605 ;
        RECT 2728.540 2012.275 2730.120 2012.605 ;
        RECT 2699.560 2006.835 2701.140 2007.165 ;
        RECT 2709.220 2006.835 2710.800 2007.165 ;
        RECT 2718.880 2006.835 2720.460 2007.165 ;
        RECT 2728.540 2006.835 2730.120 2007.165 ;
        RECT 2699.560 2001.395 2701.140 2001.725 ;
        RECT 2709.220 2001.395 2710.800 2001.725 ;
        RECT 2718.880 2001.395 2720.460 2001.725 ;
        RECT 2728.540 2001.395 2730.120 2001.725 ;
        RECT 2699.560 1995.955 2701.140 1996.285 ;
        RECT 2709.220 1995.955 2710.800 1996.285 ;
        RECT 2718.880 1995.955 2720.460 1996.285 ;
        RECT 2728.540 1995.955 2730.120 1996.285 ;
        RECT 2699.560 1990.515 2701.140 1990.845 ;
        RECT 2709.220 1990.515 2710.800 1990.845 ;
        RECT 2718.880 1990.515 2720.460 1990.845 ;
        RECT 2728.540 1990.515 2730.120 1990.845 ;
        RECT 2525.130 1984.215 2527.910 1985.745 ;
        RECT 2699.560 1985.075 2701.140 1985.405 ;
        RECT 2709.220 1985.075 2710.800 1985.405 ;
        RECT 2718.880 1985.075 2720.460 1985.405 ;
        RECT 2728.540 1985.075 2730.120 1985.405 ;
        RECT 2699.560 1979.635 2701.140 1979.965 ;
        RECT 2709.220 1979.635 2710.800 1979.965 ;
        RECT 2718.880 1979.635 2720.460 1979.965 ;
        RECT 2728.540 1979.635 2730.120 1979.965 ;
        RECT 2525.130 1976.685 2527.910 1978.215 ;
        RECT 2699.560 1974.195 2701.140 1974.525 ;
        RECT 2709.220 1974.195 2710.800 1974.525 ;
        RECT 2718.880 1974.195 2720.460 1974.525 ;
        RECT 2728.540 1974.195 2730.120 1974.525 ;
        RECT 2525.130 1970.705 2527.910 1972.235 ;
        RECT 2699.560 1968.755 2701.140 1969.085 ;
        RECT 2709.220 1968.755 2710.800 1969.085 ;
        RECT 2718.880 1968.755 2720.460 1969.085 ;
        RECT 2728.540 1968.755 2730.120 1969.085 ;
        RECT 2525.130 1964.760 2527.910 1966.290 ;
        RECT 2699.560 1963.315 2701.140 1963.645 ;
        RECT 2709.220 1963.315 2710.800 1963.645 ;
        RECT 2718.880 1963.315 2720.460 1963.645 ;
        RECT 2728.540 1963.315 2730.120 1963.645 ;
        RECT 2525.130 1959.115 2527.910 1960.645 ;
        RECT 2699.560 1957.875 2701.140 1958.205 ;
        RECT 2709.220 1957.875 2710.800 1958.205 ;
        RECT 2718.880 1957.875 2720.460 1958.205 ;
        RECT 2728.540 1957.875 2730.120 1958.205 ;
        RECT 2525.130 1953.110 2527.910 1954.640 ;
        RECT 2699.560 1952.435 2701.140 1952.765 ;
        RECT 2709.220 1952.435 2710.800 1952.765 ;
        RECT 2718.880 1952.435 2720.460 1952.765 ;
        RECT 2728.540 1952.435 2730.120 1952.765 ;
        RECT 2345.130 1948.485 2347.910 1950.015 ;
        RECT 2885.130 1894.100 2887.910 1895.630 ;
        RECT 2699.560 1854.035 2701.140 1854.365 ;
        RECT 2709.220 1854.035 2710.800 1854.365 ;
        RECT 2718.880 1854.035 2720.460 1854.365 ;
        RECT 2728.540 1854.035 2730.120 1854.365 ;
        RECT 2699.560 1848.595 2701.140 1848.925 ;
        RECT 2709.220 1848.595 2710.800 1848.925 ;
        RECT 2718.880 1848.595 2720.460 1848.925 ;
        RECT 2728.540 1848.595 2730.120 1848.925 ;
        RECT 2699.560 1843.155 2701.140 1843.485 ;
        RECT 2709.220 1843.155 2710.800 1843.485 ;
        RECT 2718.880 1843.155 2720.460 1843.485 ;
        RECT 2728.540 1843.155 2730.120 1843.485 ;
        RECT 2699.560 1837.715 2701.140 1838.045 ;
        RECT 2709.220 1837.715 2710.800 1838.045 ;
        RECT 2718.880 1837.715 2720.460 1838.045 ;
        RECT 2728.540 1837.715 2730.120 1838.045 ;
        RECT 2699.560 1832.275 2701.140 1832.605 ;
        RECT 2709.220 1832.275 2710.800 1832.605 ;
        RECT 2718.880 1832.275 2720.460 1832.605 ;
        RECT 2728.540 1832.275 2730.120 1832.605 ;
        RECT 2699.560 1826.835 2701.140 1827.165 ;
        RECT 2709.220 1826.835 2710.800 1827.165 ;
        RECT 2718.880 1826.835 2720.460 1827.165 ;
        RECT 2728.540 1826.835 2730.120 1827.165 ;
        RECT 2699.560 1821.395 2701.140 1821.725 ;
        RECT 2709.220 1821.395 2710.800 1821.725 ;
        RECT 2718.880 1821.395 2720.460 1821.725 ;
        RECT 2728.540 1821.395 2730.120 1821.725 ;
        RECT 2699.560 1815.955 2701.140 1816.285 ;
        RECT 2709.220 1815.955 2710.800 1816.285 ;
        RECT 2718.880 1815.955 2720.460 1816.285 ;
        RECT 2728.540 1815.955 2730.120 1816.285 ;
        RECT 2699.560 1810.515 2701.140 1810.845 ;
        RECT 2709.220 1810.515 2710.800 1810.845 ;
        RECT 2718.880 1810.515 2720.460 1810.845 ;
        RECT 2728.540 1810.515 2730.120 1810.845 ;
        RECT 2525.130 1807.245 2527.910 1808.775 ;
        RECT 2699.560 1805.075 2701.140 1805.405 ;
        RECT 2709.220 1805.075 2710.800 1805.405 ;
        RECT 2718.880 1805.075 2720.460 1805.405 ;
        RECT 2728.540 1805.075 2730.120 1805.405 ;
        RECT 2525.130 1799.715 2527.910 1801.245 ;
        RECT 2699.560 1799.635 2701.140 1799.965 ;
        RECT 2709.220 1799.635 2710.800 1799.965 ;
        RECT 2718.880 1799.635 2720.460 1799.965 ;
        RECT 2728.540 1799.635 2730.120 1799.965 ;
        RECT 2525.130 1793.735 2527.910 1795.265 ;
        RECT 2699.560 1794.195 2701.140 1794.525 ;
        RECT 2709.220 1794.195 2710.800 1794.525 ;
        RECT 2718.880 1794.195 2720.460 1794.525 ;
        RECT 2728.540 1794.195 2730.120 1794.525 ;
        RECT 2525.130 1787.790 2527.910 1789.320 ;
        RECT 2699.560 1788.755 2701.140 1789.085 ;
        RECT 2709.220 1788.755 2710.800 1789.085 ;
        RECT 2718.880 1788.755 2720.460 1789.085 ;
        RECT 2728.540 1788.755 2730.120 1789.085 ;
        RECT 2345.130 1785.470 2347.910 1787.000 ;
        RECT 2525.130 1782.145 2527.910 1783.675 ;
        RECT 2699.560 1783.315 2701.140 1783.645 ;
        RECT 2709.220 1783.315 2710.800 1783.645 ;
        RECT 2718.880 1783.315 2720.460 1783.645 ;
        RECT 2728.540 1783.315 2730.120 1783.645 ;
        RECT 2699.560 1777.875 2701.140 1778.205 ;
        RECT 2709.220 1777.875 2710.800 1778.205 ;
        RECT 2718.880 1777.875 2720.460 1778.205 ;
        RECT 2728.540 1777.875 2730.120 1778.205 ;
        RECT 2699.560 1772.435 2701.140 1772.765 ;
        RECT 2709.220 1772.435 2710.800 1772.765 ;
        RECT 2718.880 1772.435 2720.460 1772.765 ;
        RECT 2728.540 1772.435 2730.120 1772.765 ;
        RECT 2525.130 1770.675 2527.910 1772.205 ;
        RECT 2345.130 1705.460 2347.910 1706.990 ;
        RECT 2699.560 1674.035 2701.140 1674.365 ;
        RECT 2709.220 1674.035 2710.800 1674.365 ;
        RECT 2718.880 1674.035 2720.460 1674.365 ;
        RECT 2728.540 1674.035 2730.120 1674.365 ;
        RECT 2699.560 1668.595 2701.140 1668.925 ;
        RECT 2709.220 1668.595 2710.800 1668.925 ;
        RECT 2718.880 1668.595 2720.460 1668.925 ;
        RECT 2728.540 1668.595 2730.120 1668.925 ;
        RECT 2699.560 1663.155 2701.140 1663.485 ;
        RECT 2709.220 1663.155 2710.800 1663.485 ;
        RECT 2718.880 1663.155 2720.460 1663.485 ;
        RECT 2728.540 1663.155 2730.120 1663.485 ;
        RECT 2699.560 1657.715 2701.140 1658.045 ;
        RECT 2709.220 1657.715 2710.800 1658.045 ;
        RECT 2718.880 1657.715 2720.460 1658.045 ;
        RECT 2728.540 1657.715 2730.120 1658.045 ;
        RECT 2699.560 1652.275 2701.140 1652.605 ;
        RECT 2709.220 1652.275 2710.800 1652.605 ;
        RECT 2718.880 1652.275 2720.460 1652.605 ;
        RECT 2728.540 1652.275 2730.120 1652.605 ;
        RECT 2699.560 1646.835 2701.140 1647.165 ;
        RECT 2709.220 1646.835 2710.800 1647.165 ;
        RECT 2718.880 1646.835 2720.460 1647.165 ;
        RECT 2728.540 1646.835 2730.120 1647.165 ;
        RECT 2699.560 1641.395 2701.140 1641.725 ;
        RECT 2709.220 1641.395 2710.800 1641.725 ;
        RECT 2718.880 1641.395 2720.460 1641.725 ;
        RECT 2728.540 1641.395 2730.120 1641.725 ;
        RECT 2699.560 1635.955 2701.140 1636.285 ;
        RECT 2709.220 1635.955 2710.800 1636.285 ;
        RECT 2718.880 1635.955 2720.460 1636.285 ;
        RECT 2728.540 1635.955 2730.120 1636.285 ;
        RECT 2699.560 1630.515 2701.140 1630.845 ;
        RECT 2709.220 1630.515 2710.800 1630.845 ;
        RECT 2718.880 1630.515 2720.460 1630.845 ;
        RECT 2728.540 1630.515 2730.120 1630.845 ;
        RECT 2885.130 1628.220 2887.910 1629.750 ;
        RECT 2525.130 1626.110 2527.910 1627.640 ;
        RECT 2699.560 1625.075 2701.140 1625.405 ;
        RECT 2709.220 1625.075 2710.800 1625.405 ;
        RECT 2718.880 1625.075 2720.460 1625.405 ;
        RECT 2728.540 1625.075 2730.120 1625.405 ;
        RECT 2525.130 1619.695 2527.910 1621.225 ;
        RECT 2699.560 1619.635 2701.140 1619.965 ;
        RECT 2709.220 1619.635 2710.800 1619.965 ;
        RECT 2718.880 1619.635 2720.460 1619.965 ;
        RECT 2728.540 1619.635 2730.120 1619.965 ;
        RECT 2699.560 1614.195 2701.140 1614.525 ;
        RECT 2709.220 1614.195 2710.800 1614.525 ;
        RECT 2718.880 1614.195 2720.460 1614.525 ;
        RECT 2728.540 1614.195 2730.120 1614.525 ;
        RECT 2699.560 1608.755 2701.140 1609.085 ;
        RECT 2709.220 1608.755 2710.800 1609.085 ;
        RECT 2718.880 1608.755 2720.460 1609.085 ;
        RECT 2728.540 1608.755 2730.120 1609.085 ;
        RECT 2345.130 1605.460 2347.910 1606.990 ;
        RECT 2699.560 1603.315 2701.140 1603.645 ;
        RECT 2709.220 1603.315 2710.800 1603.645 ;
        RECT 2718.880 1603.315 2720.460 1603.645 ;
        RECT 2728.540 1603.315 2730.120 1603.645 ;
        RECT 2699.560 1597.875 2701.140 1598.205 ;
        RECT 2709.220 1597.875 2710.800 1598.205 ;
        RECT 2718.880 1597.875 2720.460 1598.205 ;
        RECT 2728.540 1597.875 2730.120 1598.205 ;
        RECT 2699.560 1592.435 2701.140 1592.765 ;
        RECT 2709.220 1592.435 2710.800 1592.765 ;
        RECT 2718.880 1592.435 2720.460 1592.765 ;
        RECT 2728.540 1592.435 2730.120 1592.765 ;
        RECT 2525.130 1590.450 2527.910 1591.980 ;
        RECT 2525.130 1582.920 2527.910 1584.450 ;
        RECT 2525.130 1576.940 2527.910 1578.470 ;
        RECT 2525.130 1568.525 2527.910 1570.055 ;
        RECT 2345.130 1528.470 2347.910 1530.000 ;
        RECT 2699.560 1494.035 2701.140 1494.365 ;
        RECT 2709.220 1494.035 2710.800 1494.365 ;
        RECT 2718.880 1494.035 2720.460 1494.365 ;
        RECT 2728.540 1494.035 2730.120 1494.365 ;
        RECT 2699.560 1488.595 2701.140 1488.925 ;
        RECT 2709.220 1488.595 2710.800 1488.925 ;
        RECT 2718.880 1488.595 2720.460 1488.925 ;
        RECT 2728.540 1488.595 2730.120 1488.925 ;
        RECT 2699.560 1483.155 2701.140 1483.485 ;
        RECT 2709.220 1483.155 2710.800 1483.485 ;
        RECT 2718.880 1483.155 2720.460 1483.485 ;
        RECT 2728.540 1483.155 2730.120 1483.485 ;
        RECT 2699.560 1477.715 2701.140 1478.045 ;
        RECT 2709.220 1477.715 2710.800 1478.045 ;
        RECT 2718.880 1477.715 2720.460 1478.045 ;
        RECT 2728.540 1477.715 2730.120 1478.045 ;
        RECT 2699.560 1472.275 2701.140 1472.605 ;
        RECT 2709.220 1472.275 2710.800 1472.605 ;
        RECT 2718.880 1472.275 2720.460 1472.605 ;
        RECT 2728.540 1472.275 2730.120 1472.605 ;
        RECT 2699.560 1466.835 2701.140 1467.165 ;
        RECT 2709.220 1466.835 2710.800 1467.165 ;
        RECT 2718.880 1466.835 2720.460 1467.165 ;
        RECT 2728.540 1466.835 2730.120 1467.165 ;
        RECT 2699.560 1461.395 2701.140 1461.725 ;
        RECT 2709.220 1461.395 2710.800 1461.725 ;
        RECT 2718.880 1461.395 2720.460 1461.725 ;
        RECT 2728.540 1461.395 2730.120 1461.725 ;
        RECT 2699.560 1455.955 2701.140 1456.285 ;
        RECT 2709.220 1455.955 2710.800 1456.285 ;
        RECT 2718.880 1455.955 2720.460 1456.285 ;
        RECT 2728.540 1455.955 2730.120 1456.285 ;
        RECT 2699.560 1450.515 2701.140 1450.845 ;
        RECT 2709.220 1450.515 2710.800 1450.845 ;
        RECT 2718.880 1450.515 2720.460 1450.845 ;
        RECT 2728.540 1450.515 2730.120 1450.845 ;
        RECT 2699.560 1445.075 2701.140 1445.405 ;
        RECT 2709.220 1445.075 2710.800 1445.405 ;
        RECT 2718.880 1445.075 2720.460 1445.405 ;
        RECT 2728.540 1445.075 2730.120 1445.405 ;
        RECT 2525.130 1438.825 2527.910 1440.355 ;
        RECT 2699.560 1439.635 2701.140 1439.965 ;
        RECT 2709.220 1439.635 2710.800 1439.965 ;
        RECT 2718.880 1439.635 2720.460 1439.965 ;
        RECT 2728.540 1439.635 2730.120 1439.965 ;
        RECT 2699.560 1434.195 2701.140 1434.525 ;
        RECT 2709.220 1434.195 2710.800 1434.525 ;
        RECT 2718.880 1434.195 2720.460 1434.525 ;
        RECT 2728.540 1434.195 2730.120 1434.525 ;
        RECT 2525.130 1432.410 2527.910 1433.940 ;
        RECT 2345.130 1430.475 2347.910 1432.005 ;
        RECT 2699.560 1428.755 2701.140 1429.085 ;
        RECT 2709.220 1428.755 2710.800 1429.085 ;
        RECT 2718.880 1428.755 2720.460 1429.085 ;
        RECT 2728.540 1428.755 2730.120 1429.085 ;
        RECT 2699.560 1423.315 2701.140 1423.645 ;
        RECT 2709.220 1423.315 2710.800 1423.645 ;
        RECT 2718.880 1423.315 2720.460 1423.645 ;
        RECT 2728.540 1423.315 2730.120 1423.645 ;
        RECT 2525.130 1418.220 2527.910 1419.750 ;
        RECT 2699.560 1417.875 2701.140 1418.205 ;
        RECT 2709.220 1417.875 2710.800 1418.205 ;
        RECT 2718.880 1417.875 2720.460 1418.205 ;
        RECT 2728.540 1417.875 2730.120 1418.205 ;
        RECT 2699.560 1412.435 2701.140 1412.765 ;
        RECT 2709.220 1412.435 2710.800 1412.765 ;
        RECT 2718.880 1412.435 2720.460 1412.765 ;
        RECT 2728.540 1412.435 2730.120 1412.765 ;
        RECT 2525.130 1410.690 2527.910 1412.220 ;
        RECT 2525.130 1404.710 2527.910 1406.240 ;
        RECT 2525.130 1396.295 2527.910 1397.825 ;
        RECT 2885.130 1363.020 2887.910 1364.550 ;
        RECT 2345.130 1330.470 2347.910 1332.000 ;
        RECT 2885.130 1163.780 2887.910 1165.310 ;
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
        RECT 4.970 -38.270 8.070 3557.950 ;
        RECT 184.970 -38.270 188.070 3557.950 ;
        RECT 364.970 -38.270 368.070 3557.950 ;
        RECT 544.970 -38.270 548.070 3557.950 ;
        RECT 724.970 -38.270 728.070 3557.950 ;
        RECT 904.970 -38.270 908.070 3557.950 ;
        RECT 1084.970 -38.270 1088.070 3557.950 ;
        RECT 1264.970 -38.270 1268.070 3557.950 ;
        RECT 1444.970 -38.270 1448.070 3557.950 ;
        RECT 1624.970 -38.270 1628.070 3557.950 ;
        RECT 1804.970 -38.270 1808.070 3557.950 ;
        RECT 1984.970 -38.270 1988.070 3557.950 ;
        RECT 2164.970 -38.270 2168.070 3557.950 ;
        RECT 2344.970 -38.270 2348.070 3557.950 ;
        RECT 2524.970 -38.270 2528.070 3557.950 ;
        RECT 2704.970 2227.860 2708.070 3557.950 ;
        RECT 2699.550 2129.640 2701.150 2217.160 ;
        RECT 2709.210 2129.640 2710.810 2217.160 ;
        RECT 2718.870 2129.640 2720.470 2217.160 ;
        RECT 2728.530 2129.640 2730.130 2217.160 ;
        RECT 2699.550 1949.640 2701.150 2037.160 ;
        RECT 2709.210 1949.640 2710.810 2037.160 ;
        RECT 2718.870 1949.640 2720.470 2037.160 ;
        RECT 2728.530 1949.640 2730.130 2037.160 ;
        RECT 2699.550 1769.640 2701.150 1857.160 ;
        RECT 2709.210 1769.640 2710.810 1857.160 ;
        RECT 2718.870 1769.640 2720.470 1857.160 ;
        RECT 2728.530 1769.640 2730.130 1857.160 ;
        RECT 2699.550 1589.640 2701.150 1677.160 ;
        RECT 2709.210 1589.640 2710.810 1677.160 ;
        RECT 2718.870 1589.640 2720.470 1677.160 ;
        RECT 2728.530 1589.640 2730.130 1677.160 ;
        RECT 2699.550 1409.640 2701.150 1497.160 ;
        RECT 2709.210 1409.640 2710.810 1497.160 ;
        RECT 2718.870 1409.640 2720.470 1497.160 ;
        RECT 2728.530 1409.640 2730.130 1497.160 ;
        RECT 2704.970 -38.270 2708.070 1398.940 ;
        RECT 2884.970 -38.270 2888.070 3557.950 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
        RECT -43.630 3430.330 2963.250 3433.430 ;
        RECT -43.630 3250.330 2963.250 3253.430 ;
        RECT -43.630 3070.330 2963.250 3073.430 ;
        RECT -43.630 2890.330 2963.250 2893.430 ;
        RECT -43.630 2710.330 2963.250 2713.430 ;
        RECT -43.630 2530.330 2963.250 2533.430 ;
        RECT -43.630 2350.330 2963.250 2353.430 ;
        RECT -43.630 2170.330 2963.250 2173.430 ;
        RECT -43.630 1990.330 2963.250 1993.430 ;
        RECT -43.630 1810.330 2963.250 1813.430 ;
        RECT -43.630 1630.330 2963.250 1633.430 ;
        RECT -43.630 1450.330 2963.250 1453.430 ;
        RECT -43.630 1270.330 2963.250 1273.430 ;
        RECT -43.630 1090.330 2963.250 1093.430 ;
        RECT -43.630 910.330 2963.250 913.430 ;
        RECT -43.630 730.330 2963.250 733.430 ;
        RECT -43.630 550.330 2963.250 553.430 ;
        RECT -43.630 370.330 2963.250 373.430 ;
        RECT -43.630 190.330 2963.250 193.430 ;
        RECT -43.630 10.330 2963.250 13.430 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
        RECT 17.370 -38.270 20.470 3557.950 ;
        RECT 197.370 -38.270 200.470 3557.950 ;
        RECT 377.370 -38.270 380.470 3557.950 ;
        RECT 557.370 -38.270 560.470 3557.950 ;
        RECT 737.370 -38.270 740.470 3557.950 ;
        RECT 917.370 -38.270 920.470 3557.950 ;
        RECT 1097.370 -38.270 1100.470 3557.950 ;
        RECT 1277.370 -38.270 1280.470 3557.950 ;
        RECT 1457.370 -38.270 1460.470 3557.950 ;
        RECT 1637.370 -38.270 1640.470 3557.950 ;
        RECT 1817.370 -38.270 1820.470 3557.950 ;
        RECT 1997.370 -38.270 2000.470 3557.950 ;
        RECT 2177.370 -38.270 2180.470 3557.950 ;
        RECT 2357.370 -38.270 2360.470 3557.950 ;
        RECT 2537.370 -38.270 2540.470 3557.950 ;
        RECT 2717.370 2227.860 2720.470 3557.950 ;
        RECT 2717.370 -38.270 2720.470 1398.940 ;
        RECT 2897.370 -38.270 2900.470 3557.950 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
        RECT -43.630 3442.730 2963.250 3445.830 ;
        RECT -43.630 3262.730 2963.250 3265.830 ;
        RECT -43.630 3082.730 2963.250 3085.830 ;
        RECT -43.630 2902.730 2963.250 2905.830 ;
        RECT -43.630 2722.730 2963.250 2725.830 ;
        RECT -43.630 2542.730 2963.250 2545.830 ;
        RECT -43.630 2362.730 2963.250 2365.830 ;
        RECT -43.630 2182.730 2963.250 2185.830 ;
        RECT -43.630 2002.730 2963.250 2005.830 ;
        RECT -43.630 1822.730 2963.250 1825.830 ;
        RECT -43.630 1642.730 2963.250 1645.830 ;
        RECT -43.630 1462.730 2963.250 1465.830 ;
        RECT -43.630 1282.730 2963.250 1285.830 ;
        RECT -43.630 1102.730 2963.250 1105.830 ;
        RECT -43.630 922.730 2963.250 925.830 ;
        RECT -43.630 742.730 2963.250 745.830 ;
        RECT -43.630 562.730 2963.250 565.830 ;
        RECT -43.630 382.730 2963.250 385.830 ;
        RECT -43.630 202.730 2963.250 205.830 ;
        RECT -43.630 22.730 2963.250 25.830 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
        RECT 29.770 -38.270 32.870 3557.950 ;
        RECT 209.770 -38.270 212.870 3557.950 ;
        RECT 389.770 -38.270 392.870 3557.950 ;
        RECT 569.770 -38.270 572.870 3557.950 ;
        RECT 749.770 -38.270 752.870 3557.950 ;
        RECT 929.770 -38.270 932.870 3557.950 ;
        RECT 1109.770 -38.270 1112.870 3557.950 ;
        RECT 1289.770 -38.270 1292.870 3557.950 ;
        RECT 1469.770 -38.270 1472.870 3557.950 ;
        RECT 1649.770 -38.270 1652.870 3557.950 ;
        RECT 1829.770 -38.270 1832.870 3557.950 ;
        RECT 2009.770 -38.270 2012.870 3557.950 ;
        RECT 2189.770 -38.270 2192.870 3557.950 ;
        RECT 2369.770 1795.300 2372.870 3557.950 ;
        RECT 2369.770 1340.300 2372.870 1773.075 ;
        RECT 2369.770 -38.270 2372.870 1318.075 ;
        RECT 2549.770 -38.270 2552.870 3557.950 ;
        RECT 2729.770 2227.860 2732.870 3557.950 ;
        RECT 2729.770 -38.270 2732.870 1398.940 ;
        RECT 2909.770 -38.270 2912.870 3557.950 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
        RECT -43.630 3455.130 2963.250 3458.230 ;
        RECT -43.630 3275.130 2963.250 3278.230 ;
        RECT -43.630 3095.130 2963.250 3098.230 ;
        RECT -43.630 2915.130 2963.250 2918.230 ;
        RECT -43.630 2735.130 2963.250 2738.230 ;
        RECT -43.630 2555.130 2963.250 2558.230 ;
        RECT -43.630 2375.130 2963.250 2378.230 ;
        RECT -43.630 2195.130 2963.250 2198.230 ;
        RECT -43.630 2015.130 2963.250 2018.230 ;
        RECT -43.630 1835.130 2963.250 1838.230 ;
        RECT -43.630 1655.130 2963.250 1658.230 ;
        RECT -43.630 1475.130 2963.250 1478.230 ;
        RECT -43.630 1295.130 2963.250 1298.230 ;
        RECT -43.630 1115.130 2963.250 1118.230 ;
        RECT -43.630 935.130 2963.250 938.230 ;
        RECT -43.630 755.130 2963.250 758.230 ;
        RECT -43.630 575.130 2963.250 578.230 ;
        RECT -43.630 395.130 2963.250 398.230 ;
        RECT -43.630 215.130 2963.250 218.230 ;
        RECT -43.630 35.130 2963.250 38.230 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
        RECT 42.170 -38.270 45.270 3557.950 ;
        RECT 222.170 -38.270 225.270 3557.950 ;
        RECT 402.170 -38.270 405.270 3557.950 ;
        RECT 582.170 -38.270 585.270 3557.950 ;
        RECT 762.170 -38.270 765.270 3557.950 ;
        RECT 942.170 -38.270 945.270 3557.950 ;
        RECT 1122.170 -38.270 1125.270 3557.950 ;
        RECT 1302.170 -38.270 1305.270 3557.950 ;
        RECT 1482.170 -38.270 1485.270 3557.950 ;
        RECT 1662.170 -38.270 1665.270 3557.950 ;
        RECT 1842.170 -38.270 1845.270 3557.950 ;
        RECT 2022.170 -38.270 2025.270 3557.950 ;
        RECT 2202.170 -38.270 2205.270 3557.950 ;
        RECT 2382.170 1795.300 2385.270 3557.950 ;
        RECT 2382.170 1340.300 2385.270 1773.075 ;
        RECT 2382.170 -38.270 2385.270 1318.075 ;
        RECT 2562.170 -38.270 2565.270 3557.950 ;
        RECT 2742.170 -38.270 2745.270 3557.950 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
        RECT -43.630 3467.530 2963.250 3470.630 ;
        RECT -43.630 3287.530 2963.250 3290.630 ;
        RECT -43.630 3107.530 2963.250 3110.630 ;
        RECT -43.630 2927.530 2963.250 2930.630 ;
        RECT -43.630 2747.530 2963.250 2750.630 ;
        RECT -43.630 2567.530 2963.250 2570.630 ;
        RECT -43.630 2387.530 2963.250 2390.630 ;
        RECT -43.630 2207.530 2963.250 2210.630 ;
        RECT -43.630 2027.530 2963.250 2030.630 ;
        RECT -43.630 1847.530 2963.250 1850.630 ;
        RECT -43.630 1667.530 2963.250 1670.630 ;
        RECT -43.630 1487.530 2963.250 1490.630 ;
        RECT -43.630 1307.530 2963.250 1310.630 ;
        RECT -43.630 1127.530 2963.250 1130.630 ;
        RECT -43.630 947.530 2963.250 950.630 ;
        RECT -43.630 767.530 2963.250 770.630 ;
        RECT -43.630 587.530 2963.250 590.630 ;
        RECT -43.630 407.530 2963.250 410.630 ;
        RECT -43.630 227.530 2963.250 230.630 ;
        RECT -43.630 47.530 2963.250 50.630 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
        RECT 35.970 -38.270 39.070 3557.950 ;
        RECT 215.970 -38.270 219.070 3557.950 ;
        RECT 395.970 -38.270 399.070 3557.950 ;
        RECT 575.970 -38.270 579.070 3557.950 ;
        RECT 755.970 -38.270 759.070 3557.950 ;
        RECT 935.970 -38.270 939.070 3557.950 ;
        RECT 1115.970 -38.270 1119.070 3557.950 ;
        RECT 1295.970 -38.270 1299.070 3557.950 ;
        RECT 1475.970 -38.270 1479.070 3557.950 ;
        RECT 1655.970 -38.270 1659.070 3557.950 ;
        RECT 1835.970 -38.270 1839.070 3557.950 ;
        RECT 2015.970 -38.270 2019.070 3557.950 ;
        RECT 2195.970 -38.270 2199.070 3557.950 ;
        RECT 2375.970 1795.300 2379.070 3557.950 ;
        RECT 2375.970 1340.300 2379.070 1773.075 ;
        RECT 2375.970 -38.270 2379.070 1318.075 ;
        RECT 2555.970 -38.270 2559.070 3557.950 ;
        RECT 2735.970 -38.270 2739.070 3557.950 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
        RECT -43.630 3461.330 2963.250 3464.430 ;
        RECT -43.630 3281.330 2963.250 3284.430 ;
        RECT -43.630 3101.330 2963.250 3104.430 ;
        RECT -43.630 2921.330 2963.250 2924.430 ;
        RECT -43.630 2741.330 2963.250 2744.430 ;
        RECT -43.630 2561.330 2963.250 2564.430 ;
        RECT -43.630 2381.330 2963.250 2384.430 ;
        RECT -43.630 2201.330 2963.250 2204.430 ;
        RECT -43.630 2021.330 2963.250 2024.430 ;
        RECT -43.630 1841.330 2963.250 1844.430 ;
        RECT -43.630 1661.330 2963.250 1664.430 ;
        RECT -43.630 1481.330 2963.250 1484.430 ;
        RECT -43.630 1301.330 2963.250 1304.430 ;
        RECT -43.630 1121.330 2963.250 1124.430 ;
        RECT -43.630 941.330 2963.250 944.430 ;
        RECT -43.630 761.330 2963.250 764.430 ;
        RECT -43.630 581.330 2963.250 584.430 ;
        RECT -43.630 401.330 2963.250 404.430 ;
        RECT -43.630 221.330 2963.250 224.430 ;
        RECT -43.630 41.330 2963.250 44.430 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
        RECT 48.370 -38.270 51.470 3557.950 ;
        RECT 228.370 -38.270 231.470 3557.950 ;
        RECT 408.370 -38.270 411.470 3557.950 ;
        RECT 588.370 -38.270 591.470 3557.950 ;
        RECT 768.370 -38.270 771.470 3557.950 ;
        RECT 948.370 -38.270 951.470 3557.950 ;
        RECT 1128.370 -38.270 1131.470 3557.950 ;
        RECT 1308.370 -38.270 1311.470 3557.950 ;
        RECT 1488.370 -38.270 1491.470 3557.950 ;
        RECT 1668.370 -38.270 1671.470 3557.950 ;
        RECT 1848.370 -38.270 1851.470 3557.950 ;
        RECT 2028.370 -38.270 2031.470 3557.950 ;
        RECT 2208.370 -38.270 2211.470 3557.950 ;
        RECT 2388.370 1795.300 2391.470 3557.950 ;
        RECT 2388.370 1340.300 2391.470 1773.075 ;
        RECT 2388.370 -38.270 2391.470 1318.075 ;
        RECT 2568.370 -38.270 2571.470 3557.950 ;
        RECT 2748.370 -38.270 2751.470 3557.950 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
        RECT -43.630 3473.730 2963.250 3476.830 ;
        RECT -43.630 3293.730 2963.250 3296.830 ;
        RECT -43.630 3113.730 2963.250 3116.830 ;
        RECT -43.630 2933.730 2963.250 2936.830 ;
        RECT -43.630 2753.730 2963.250 2756.830 ;
        RECT -43.630 2573.730 2963.250 2576.830 ;
        RECT -43.630 2393.730 2963.250 2396.830 ;
        RECT -43.630 2213.730 2963.250 2216.830 ;
        RECT -43.630 2033.730 2963.250 2036.830 ;
        RECT -43.630 1853.730 2963.250 1856.830 ;
        RECT -43.630 1673.730 2963.250 1676.830 ;
        RECT -43.630 1493.730 2963.250 1496.830 ;
        RECT -43.630 1313.730 2963.250 1316.830 ;
        RECT -43.630 1133.730 2963.250 1136.830 ;
        RECT -43.630 953.730 2963.250 956.830 ;
        RECT -43.630 773.730 2963.250 776.830 ;
        RECT -43.630 593.730 2963.250 596.830 ;
        RECT -43.630 413.730 2963.250 416.830 ;
        RECT -43.630 233.730 2963.250 236.830 ;
        RECT -43.630 53.730 2963.250 56.830 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2708.415 2215.945 2708.845 2216.730 ;
        RECT 2721.295 2215.945 2721.725 2216.730 ;
        RECT 2708.415 2211.670 2708.845 2212.455 ;
        RECT 2721.295 2210.505 2721.725 2211.290 ;
        RECT 2708.415 2206.230 2708.845 2207.015 ;
        RECT 2721.295 2205.065 2721.725 2205.850 ;
        RECT 2708.415 2200.790 2708.845 2201.575 ;
        RECT 2721.295 2199.625 2721.725 2200.410 ;
        RECT 2708.415 2195.350 2708.845 2196.135 ;
        RECT 2721.295 2194.185 2721.725 2194.970 ;
        RECT 2708.415 2189.910 2708.845 2190.695 ;
        RECT 2721.295 2188.745 2721.725 2189.530 ;
        RECT 2708.415 2184.470 2708.845 2185.255 ;
        RECT 2721.295 2183.305 2721.725 2184.090 ;
        RECT 2708.415 2179.030 2708.845 2179.815 ;
        RECT 2721.295 2177.865 2721.725 2178.650 ;
        RECT 2708.415 2173.590 2708.845 2174.375 ;
        RECT 2721.295 2172.425 2721.725 2173.210 ;
        RECT 2708.415 2168.150 2708.845 2168.935 ;
        RECT 2721.295 2166.985 2721.725 2167.770 ;
        RECT 2708.415 2162.710 2708.845 2163.495 ;
        RECT 2721.295 2161.545 2721.725 2162.330 ;
        RECT 2708.415 2157.270 2708.845 2158.055 ;
        RECT 2721.295 2156.105 2721.725 2156.890 ;
        RECT 2708.415 2151.830 2708.845 2152.615 ;
        RECT 2721.295 2150.665 2721.725 2151.450 ;
        RECT 2708.415 2146.390 2708.845 2147.175 ;
        RECT 2721.295 2145.225 2721.725 2146.010 ;
        RECT 2708.415 2140.950 2708.845 2141.735 ;
        RECT 2721.295 2139.785 2721.725 2140.570 ;
        RECT 2708.415 2135.510 2708.845 2136.295 ;
        RECT 2721.295 2134.345 2721.725 2135.130 ;
        RECT 2708.415 2130.070 2708.845 2130.855 ;
        RECT 2721.295 2130.070 2721.725 2130.855 ;
        RECT 2708.415 2035.945 2708.845 2036.730 ;
        RECT 2721.295 2035.945 2721.725 2036.730 ;
        RECT 2708.415 2031.670 2708.845 2032.455 ;
        RECT 2721.295 2030.505 2721.725 2031.290 ;
        RECT 2708.415 2026.230 2708.845 2027.015 ;
        RECT 2721.295 2025.065 2721.725 2025.850 ;
        RECT 2708.415 2020.790 2708.845 2021.575 ;
        RECT 2721.295 2019.625 2721.725 2020.410 ;
        RECT 2708.415 2015.350 2708.845 2016.135 ;
        RECT 2721.295 2014.185 2721.725 2014.970 ;
        RECT 2708.415 2009.910 2708.845 2010.695 ;
        RECT 2721.295 2008.745 2721.725 2009.530 ;
        RECT 2708.415 2004.470 2708.845 2005.255 ;
        RECT 2721.295 2003.305 2721.725 2004.090 ;
        RECT 2708.415 1999.030 2708.845 1999.815 ;
        RECT 2721.295 1997.865 2721.725 1998.650 ;
        RECT 2708.415 1993.590 2708.845 1994.375 ;
        RECT 2721.295 1992.425 2721.725 1993.210 ;
        RECT 2708.415 1988.150 2708.845 1988.935 ;
        RECT 2721.295 1986.985 2721.725 1987.770 ;
        RECT 2708.415 1982.710 2708.845 1983.495 ;
        RECT 2721.295 1981.545 2721.725 1982.330 ;
        RECT 2708.415 1977.270 2708.845 1978.055 ;
        RECT 2721.295 1976.105 2721.725 1976.890 ;
        RECT 2708.415 1971.830 2708.845 1972.615 ;
        RECT 2721.295 1970.665 2721.725 1971.450 ;
        RECT 2708.415 1966.390 2708.845 1967.175 ;
        RECT 2721.295 1965.225 2721.725 1966.010 ;
        RECT 2708.415 1960.950 2708.845 1961.735 ;
        RECT 2721.295 1959.785 2721.725 1960.570 ;
        RECT 2708.415 1955.510 2708.845 1956.295 ;
        RECT 2721.295 1954.345 2721.725 1955.130 ;
        RECT 2708.415 1950.070 2708.845 1950.855 ;
        RECT 2721.295 1950.070 2721.725 1950.855 ;
        RECT 2708.415 1855.945 2708.845 1856.730 ;
        RECT 2721.295 1855.945 2721.725 1856.730 ;
        RECT 2708.415 1851.670 2708.845 1852.455 ;
        RECT 2721.295 1850.505 2721.725 1851.290 ;
        RECT 2708.415 1846.230 2708.845 1847.015 ;
        RECT 2721.295 1845.065 2721.725 1845.850 ;
        RECT 2708.415 1840.790 2708.845 1841.575 ;
        RECT 2721.295 1839.625 2721.725 1840.410 ;
        RECT 2708.415 1835.350 2708.845 1836.135 ;
        RECT 2721.295 1834.185 2721.725 1834.970 ;
        RECT 2708.415 1829.910 2708.845 1830.695 ;
        RECT 2721.295 1828.745 2721.725 1829.530 ;
        RECT 2708.415 1824.470 2708.845 1825.255 ;
        RECT 2721.295 1823.305 2721.725 1824.090 ;
        RECT 2708.415 1819.030 2708.845 1819.815 ;
        RECT 2721.295 1817.865 2721.725 1818.650 ;
        RECT 2708.415 1813.590 2708.845 1814.375 ;
        RECT 2721.295 1812.425 2721.725 1813.210 ;
        RECT 2708.415 1808.150 2708.845 1808.935 ;
        RECT 2721.295 1806.985 2721.725 1807.770 ;
        RECT 2708.415 1802.710 2708.845 1803.495 ;
        RECT 2721.295 1801.545 2721.725 1802.330 ;
        RECT 2708.415 1797.270 2708.845 1798.055 ;
        RECT 2721.295 1796.105 2721.725 1796.890 ;
        RECT 2708.415 1791.830 2708.845 1792.615 ;
        RECT 2721.295 1790.665 2721.725 1791.450 ;
        RECT 2708.415 1786.390 2708.845 1787.175 ;
        RECT 2721.295 1785.225 2721.725 1786.010 ;
        RECT 2708.415 1780.950 2708.845 1781.735 ;
        RECT 2721.295 1779.785 2721.725 1780.570 ;
        RECT 2708.415 1775.510 2708.845 1776.295 ;
        RECT 2721.295 1774.345 2721.725 1775.130 ;
        RECT 2708.415 1770.070 2708.845 1770.855 ;
        RECT 2721.295 1770.070 2721.725 1770.855 ;
        RECT 2708.415 1675.945 2708.845 1676.730 ;
        RECT 2721.295 1675.945 2721.725 1676.730 ;
        RECT 2708.415 1671.670 2708.845 1672.455 ;
        RECT 2721.295 1670.505 2721.725 1671.290 ;
        RECT 2708.415 1666.230 2708.845 1667.015 ;
        RECT 2721.295 1665.065 2721.725 1665.850 ;
        RECT 2708.415 1660.790 2708.845 1661.575 ;
        RECT 2721.295 1659.625 2721.725 1660.410 ;
        RECT 2708.415 1655.350 2708.845 1656.135 ;
        RECT 2721.295 1654.185 2721.725 1654.970 ;
        RECT 2708.415 1649.910 2708.845 1650.695 ;
        RECT 2721.295 1648.745 2721.725 1649.530 ;
        RECT 2708.415 1644.470 2708.845 1645.255 ;
        RECT 2721.295 1643.305 2721.725 1644.090 ;
        RECT 2708.415 1639.030 2708.845 1639.815 ;
        RECT 2721.295 1637.865 2721.725 1638.650 ;
        RECT 2708.415 1633.590 2708.845 1634.375 ;
        RECT 2721.295 1632.425 2721.725 1633.210 ;
        RECT 2708.415 1628.150 2708.845 1628.935 ;
        RECT 2721.295 1626.985 2721.725 1627.770 ;
        RECT 2708.415 1622.710 2708.845 1623.495 ;
        RECT 2721.295 1621.545 2721.725 1622.330 ;
        RECT 2708.415 1617.270 2708.845 1618.055 ;
        RECT 2721.295 1616.105 2721.725 1616.890 ;
        RECT 2708.415 1611.830 2708.845 1612.615 ;
        RECT 2721.295 1610.665 2721.725 1611.450 ;
        RECT 2708.415 1606.390 2708.845 1607.175 ;
        RECT 2721.295 1605.225 2721.725 1606.010 ;
        RECT 2708.415 1600.950 2708.845 1601.735 ;
        RECT 2721.295 1599.785 2721.725 1600.570 ;
        RECT 2708.415 1595.510 2708.845 1596.295 ;
        RECT 2721.295 1594.345 2721.725 1595.130 ;
        RECT 2708.415 1590.070 2708.845 1590.855 ;
        RECT 2721.295 1590.070 2721.725 1590.855 ;
        RECT 2708.415 1495.945 2708.845 1496.730 ;
        RECT 2721.295 1495.945 2721.725 1496.730 ;
        RECT 2708.415 1491.670 2708.845 1492.455 ;
        RECT 2721.295 1490.505 2721.725 1491.290 ;
        RECT 2708.415 1486.230 2708.845 1487.015 ;
        RECT 2721.295 1485.065 2721.725 1485.850 ;
        RECT 2708.415 1480.790 2708.845 1481.575 ;
        RECT 2721.295 1479.625 2721.725 1480.410 ;
        RECT 2708.415 1475.350 2708.845 1476.135 ;
        RECT 2721.295 1474.185 2721.725 1474.970 ;
        RECT 2708.415 1469.910 2708.845 1470.695 ;
        RECT 2721.295 1468.745 2721.725 1469.530 ;
        RECT 2708.415 1464.470 2708.845 1465.255 ;
        RECT 2721.295 1463.305 2721.725 1464.090 ;
        RECT 2708.415 1459.030 2708.845 1459.815 ;
        RECT 2721.295 1457.865 2721.725 1458.650 ;
        RECT 2708.415 1453.590 2708.845 1454.375 ;
        RECT 2721.295 1452.425 2721.725 1453.210 ;
        RECT 2708.415 1448.150 2708.845 1448.935 ;
        RECT 2721.295 1446.985 2721.725 1447.770 ;
        RECT 2708.415 1442.710 2708.845 1443.495 ;
        RECT 2721.295 1441.545 2721.725 1442.330 ;
        RECT 2708.415 1437.270 2708.845 1438.055 ;
        RECT 2721.295 1436.105 2721.725 1436.890 ;
        RECT 2708.415 1431.830 2708.845 1432.615 ;
        RECT 2721.295 1430.665 2721.725 1431.450 ;
        RECT 2708.415 1426.390 2708.845 1427.175 ;
        RECT 2721.295 1425.225 2721.725 1426.010 ;
        RECT 2708.415 1420.950 2708.845 1421.735 ;
        RECT 2721.295 1419.785 2721.725 1420.570 ;
        RECT 2708.415 1415.510 2708.845 1416.295 ;
        RECT 2721.295 1414.345 2721.725 1415.130 ;
        RECT 2708.415 1410.070 2708.845 1410.855 ;
        RECT 2721.295 1410.070 2721.725 1410.855 ;
      LAYER li1 ;
        RECT 1622.380 3512.755 1624.185 3512.925 ;
        RECT 1262.805 3512.305 1264.185 3512.475 ;
        RECT 1263.580 3511.645 1263.920 3512.305 ;
        RECT 1623.580 3512.095 1623.920 3512.755 ;
        RECT 2522.380 3511.160 2524.185 3511.330 ;
        RECT 1802.380 3510.835 1804.185 3511.005 ;
        RECT 1803.580 3510.175 1803.920 3510.835 ;
        RECT 2162.380 3510.475 2164.185 3510.645 ;
        RECT 2523.580 3510.500 2523.920 3511.160 ;
        RECT 2163.580 3509.815 2163.920 3510.475 ;
        RECT 2882.265 3485.590 2882.605 3486.250 ;
        RECT 2881.575 3485.420 2883.380 3485.590 ;
        RECT 2882.265 3219.710 2882.605 3220.370 ;
        RECT 2881.575 3219.540 2883.380 3219.710 ;
        RECT 2882.265 2954.510 2882.605 2955.170 ;
        RECT 2881.575 2954.340 2883.380 2954.510 ;
        RECT 2882.265 2688.630 2882.605 2689.290 ;
        RECT 2881.575 2688.460 2883.380 2688.630 ;
        RECT 2882.265 2422.750 2882.605 2423.410 ;
        RECT 2881.575 2422.580 2883.380 2422.750 ;
        RECT 2343.055 2255.855 2443.725 2257.455 ;
        RECT 2358.225 2255.225 2358.395 2255.855 ;
        RECT 2361.455 2255.225 2361.625 2255.855 ;
        RECT 2362.410 2255.305 2362.580 2255.585 ;
        RECT 2362.410 2255.135 2362.640 2255.305 ;
        RECT 2362.470 2253.525 2362.640 2255.135 ;
        RECT 2364.515 2253.525 2364.765 2255.855 ;
        RECT 2365.040 2253.525 2365.315 2255.855 ;
        RECT 2365.590 2253.525 2365.865 2255.855 ;
        RECT 2366.140 2253.525 2366.415 2255.855 ;
        RECT 2366.690 2253.525 2366.965 2255.855 ;
        RECT 2367.240 2253.525 2367.515 2255.855 ;
        RECT 2367.790 2253.525 2368.065 2255.855 ;
        RECT 2368.340 2253.525 2368.615 2255.855 ;
        RECT 2368.890 2253.525 2369.165 2255.855 ;
        RECT 2369.440 2253.525 2369.715 2255.855 ;
        RECT 2369.990 2253.525 2370.265 2255.855 ;
        RECT 2370.540 2253.525 2370.815 2255.855 ;
        RECT 2371.090 2253.525 2371.435 2255.855 ;
        RECT 2372.680 2255.230 2372.850 2255.855 ;
        RECT 2375.425 2255.230 2375.595 2255.855 ;
        RECT 2376.415 2255.230 2376.585 2255.855 ;
        RECT 2378.040 2255.225 2378.210 2255.855 ;
        RECT 2378.995 2255.305 2379.165 2255.585 ;
        RECT 2378.995 2255.135 2379.225 2255.305 ;
        RECT 2379.055 2253.525 2379.225 2255.135 ;
        RECT 2381.100 2253.525 2381.350 2255.855 ;
        RECT 2381.625 2253.525 2381.900 2255.855 ;
        RECT 2382.175 2253.525 2382.450 2255.855 ;
        RECT 2382.725 2253.525 2383.000 2255.855 ;
        RECT 2383.275 2253.525 2383.550 2255.855 ;
        RECT 2383.825 2253.525 2384.100 2255.855 ;
        RECT 2384.375 2253.525 2384.650 2255.855 ;
        RECT 2384.925 2253.525 2385.200 2255.855 ;
        RECT 2385.475 2253.525 2385.750 2255.855 ;
        RECT 2386.025 2253.525 2386.300 2255.855 ;
        RECT 2386.575 2253.525 2386.850 2255.855 ;
        RECT 2387.125 2253.525 2387.400 2255.855 ;
        RECT 2387.675 2253.525 2388.020 2255.855 ;
        RECT 2389.265 2255.230 2389.435 2255.855 ;
        RECT 2392.010 2255.230 2392.180 2255.855 ;
        RECT 2393.000 2255.230 2393.170 2255.855 ;
        RECT 2394.625 2255.225 2394.795 2255.855 ;
        RECT 2395.580 2255.305 2395.750 2255.585 ;
        RECT 2395.580 2255.135 2395.810 2255.305 ;
        RECT 2395.640 2253.525 2395.810 2255.135 ;
        RECT 2397.685 2253.525 2397.935 2255.855 ;
        RECT 2398.210 2253.525 2398.485 2255.855 ;
        RECT 2398.760 2253.525 2399.035 2255.855 ;
        RECT 2399.310 2253.525 2399.585 2255.855 ;
        RECT 2399.860 2253.525 2400.135 2255.855 ;
        RECT 2400.410 2253.525 2400.685 2255.855 ;
        RECT 2400.960 2253.525 2401.235 2255.855 ;
        RECT 2401.510 2253.525 2401.785 2255.855 ;
        RECT 2402.060 2253.525 2402.335 2255.855 ;
        RECT 2402.610 2253.525 2402.885 2255.855 ;
        RECT 2403.160 2253.525 2403.435 2255.855 ;
        RECT 2403.710 2253.525 2403.985 2255.855 ;
        RECT 2404.260 2253.525 2404.605 2255.855 ;
        RECT 2405.850 2255.230 2406.020 2255.855 ;
        RECT 2408.595 2255.230 2408.765 2255.855 ;
        RECT 2409.585 2255.230 2409.755 2255.855 ;
        RECT 2411.210 2255.225 2411.380 2255.855 ;
        RECT 2412.165 2255.305 2412.335 2255.585 ;
        RECT 2412.165 2255.135 2412.395 2255.305 ;
        RECT 2412.225 2253.525 2412.395 2255.135 ;
        RECT 2414.270 2253.525 2414.520 2255.855 ;
        RECT 2414.795 2253.525 2415.070 2255.855 ;
        RECT 2415.345 2253.525 2415.620 2255.855 ;
        RECT 2415.895 2253.525 2416.170 2255.855 ;
        RECT 2416.445 2253.525 2416.720 2255.855 ;
        RECT 2416.995 2253.525 2417.270 2255.855 ;
        RECT 2417.545 2253.525 2417.820 2255.855 ;
        RECT 2418.095 2253.525 2418.370 2255.855 ;
        RECT 2418.645 2253.525 2418.920 2255.855 ;
        RECT 2419.195 2253.525 2419.470 2255.855 ;
        RECT 2419.745 2253.525 2420.020 2255.855 ;
        RECT 2420.295 2253.525 2420.570 2255.855 ;
        RECT 2420.845 2253.525 2421.190 2255.855 ;
        RECT 2422.435 2255.230 2422.605 2255.855 ;
        RECT 2425.180 2255.230 2425.350 2255.855 ;
        RECT 2426.170 2255.230 2426.340 2255.855 ;
        RECT 2427.790 2255.225 2427.960 2255.855 ;
        RECT 2428.745 2255.305 2428.915 2255.585 ;
        RECT 2428.745 2255.135 2428.975 2255.305 ;
        RECT 2428.805 2253.525 2428.975 2255.135 ;
        RECT 2430.850 2253.525 2431.100 2255.855 ;
        RECT 2431.375 2253.525 2431.650 2255.855 ;
        RECT 2431.925 2253.525 2432.200 2255.855 ;
        RECT 2432.475 2253.525 2432.750 2255.855 ;
        RECT 2433.025 2253.525 2433.300 2255.855 ;
        RECT 2433.575 2253.525 2433.850 2255.855 ;
        RECT 2434.125 2253.525 2434.400 2255.855 ;
        RECT 2434.675 2253.525 2434.950 2255.855 ;
        RECT 2435.225 2253.525 2435.500 2255.855 ;
        RECT 2435.775 2253.525 2436.050 2255.855 ;
        RECT 2436.325 2253.525 2436.600 2255.855 ;
        RECT 2436.875 2253.525 2437.150 2255.855 ;
        RECT 2437.425 2253.525 2437.770 2255.855 ;
        RECT 2439.015 2255.230 2439.185 2255.855 ;
        RECT 2441.760 2255.230 2441.930 2255.855 ;
        RECT 2442.750 2255.230 2442.920 2255.855 ;
        RECT 2362.410 2253.355 2362.640 2253.525 ;
        RECT 2364.380 2253.355 2371.435 2253.525 ;
        RECT 2378.995 2253.355 2379.225 2253.525 ;
        RECT 2380.965 2253.355 2388.020 2253.525 ;
        RECT 2395.580 2253.355 2395.810 2253.525 ;
        RECT 2397.550 2253.355 2404.605 2253.525 ;
        RECT 2412.165 2253.355 2412.395 2253.525 ;
        RECT 2414.135 2253.355 2421.190 2253.525 ;
        RECT 2428.745 2253.355 2428.975 2253.525 ;
        RECT 2430.715 2253.355 2437.770 2253.525 ;
        RECT 2362.410 2252.295 2362.580 2253.355 ;
        RECT 2365.790 2252.895 2366.040 2253.355 ;
        RECT 2367.860 2252.955 2368.190 2253.355 ;
        RECT 2369.950 2252.845 2370.400 2253.355 ;
        RECT 2365.940 2252.115 2366.280 2252.365 ;
        RECT 2368.160 2252.115 2368.490 2252.445 ;
        RECT 2378.995 2252.295 2379.165 2253.355 ;
        RECT 2382.375 2252.895 2382.625 2253.355 ;
        RECT 2384.445 2252.955 2384.775 2253.355 ;
        RECT 2386.535 2252.845 2386.985 2253.355 ;
        RECT 2382.525 2252.115 2382.865 2252.365 ;
        RECT 2384.745 2252.115 2385.075 2252.445 ;
        RECT 2395.580 2252.295 2395.750 2253.355 ;
        RECT 2398.960 2252.895 2399.210 2253.355 ;
        RECT 2401.030 2252.955 2401.360 2253.355 ;
        RECT 2403.120 2252.845 2403.570 2253.355 ;
        RECT 2399.110 2252.115 2399.450 2252.365 ;
        RECT 2401.330 2252.115 2401.660 2252.445 ;
        RECT 2412.165 2252.295 2412.335 2253.355 ;
        RECT 2415.545 2252.895 2415.795 2253.355 ;
        RECT 2417.615 2252.955 2417.945 2253.355 ;
        RECT 2419.705 2252.845 2420.155 2253.355 ;
        RECT 2415.695 2252.115 2416.035 2252.365 ;
        RECT 2417.915 2252.115 2418.245 2252.445 ;
        RECT 2428.745 2252.295 2428.915 2253.355 ;
        RECT 2432.125 2252.895 2432.375 2253.355 ;
        RECT 2434.195 2252.955 2434.525 2253.355 ;
        RECT 2436.285 2252.845 2436.735 2253.355 ;
        RECT 2432.275 2252.115 2432.615 2252.365 ;
        RECT 2434.495 2252.115 2434.825 2252.445 ;
        RECT 2364.300 2248.355 2364.555 2248.905 ;
        RECT 2364.300 2248.095 2364.560 2248.355 ;
        RECT 2366.890 2248.095 2367.220 2248.545 ;
        RECT 2369.270 2248.095 2369.520 2248.625 ;
        RECT 2370.140 2248.095 2370.380 2248.895 ;
        RECT 2371.050 2248.095 2371.320 2248.895 ;
        RECT 2380.885 2248.355 2381.140 2248.905 ;
        RECT 2380.885 2248.095 2381.145 2248.355 ;
        RECT 2383.475 2248.095 2383.805 2248.545 ;
        RECT 2385.855 2248.095 2386.105 2248.625 ;
        RECT 2386.725 2248.095 2386.965 2248.895 ;
        RECT 2387.635 2248.095 2387.905 2248.895 ;
        RECT 2397.470 2248.355 2397.725 2248.905 ;
        RECT 2397.470 2248.095 2397.730 2248.355 ;
        RECT 2400.060 2248.095 2400.390 2248.545 ;
        RECT 2402.440 2248.095 2402.690 2248.625 ;
        RECT 2403.310 2248.095 2403.550 2248.895 ;
        RECT 2404.220 2248.095 2404.490 2248.895 ;
        RECT 2414.055 2248.355 2414.310 2248.905 ;
        RECT 2414.055 2248.095 2414.315 2248.355 ;
        RECT 2416.645 2248.095 2416.975 2248.545 ;
        RECT 2419.025 2248.095 2419.275 2248.625 ;
        RECT 2419.895 2248.095 2420.135 2248.895 ;
        RECT 2420.805 2248.095 2421.075 2248.895 ;
        RECT 2430.635 2248.355 2430.890 2248.905 ;
        RECT 2430.635 2248.095 2430.895 2248.355 ;
        RECT 2433.225 2248.095 2433.555 2248.545 ;
        RECT 2435.605 2248.095 2435.855 2248.625 ;
        RECT 2436.475 2248.095 2436.715 2248.895 ;
        RECT 2437.385 2248.095 2437.655 2248.895 ;
        RECT 2364.220 2247.925 2371.610 2248.095 ;
        RECT 2380.805 2247.925 2388.195 2248.095 ;
        RECT 2397.390 2247.925 2404.780 2248.095 ;
        RECT 2413.975 2247.925 2421.365 2248.095 ;
        RECT 2430.555 2247.925 2437.945 2248.095 ;
        RECT 2364.265 2246.600 2364.525 2247.925 ;
        RECT 2364.815 2246.600 2365.075 2247.925 ;
        RECT 2365.355 2246.600 2365.615 2247.925 ;
        RECT 2365.895 2246.600 2366.135 2247.925 ;
        RECT 2366.435 2246.600 2366.675 2247.925 ;
        RECT 2366.955 2246.600 2367.195 2247.925 ;
        RECT 2367.475 2246.600 2367.715 2247.925 ;
        RECT 2367.995 2246.600 2368.235 2247.925 ;
        RECT 2368.515 2246.600 2368.755 2247.925 ;
        RECT 2368.995 2246.600 2369.235 2247.925 ;
        RECT 2369.475 2246.600 2369.715 2247.925 ;
        RECT 2369.955 2246.600 2370.195 2247.925 ;
        RECT 2370.435 2246.600 2370.675 2247.925 ;
        RECT 2370.915 2246.600 2371.155 2247.925 ;
        RECT 2371.395 2246.600 2371.610 2247.925 ;
        RECT 2372.680 2246.600 2372.850 2247.230 ;
        RECT 2375.425 2246.600 2375.595 2247.230 ;
        RECT 2376.415 2246.600 2376.585 2247.230 ;
        RECT 2380.850 2246.600 2381.110 2247.925 ;
        RECT 2381.400 2246.600 2381.660 2247.925 ;
        RECT 2381.940 2246.600 2382.200 2247.925 ;
        RECT 2382.480 2246.600 2382.720 2247.925 ;
        RECT 2383.020 2246.600 2383.260 2247.925 ;
        RECT 2383.540 2246.600 2383.780 2247.925 ;
        RECT 2384.060 2246.600 2384.300 2247.925 ;
        RECT 2384.580 2246.600 2384.820 2247.925 ;
        RECT 2385.100 2246.600 2385.340 2247.925 ;
        RECT 2385.580 2246.600 2385.820 2247.925 ;
        RECT 2386.060 2246.600 2386.300 2247.925 ;
        RECT 2386.540 2246.600 2386.780 2247.925 ;
        RECT 2387.020 2246.600 2387.260 2247.925 ;
        RECT 2387.500 2246.600 2387.740 2247.925 ;
        RECT 2387.980 2246.600 2388.195 2247.925 ;
        RECT 2389.265 2246.600 2389.435 2247.230 ;
        RECT 2392.010 2246.600 2392.180 2247.230 ;
        RECT 2393.000 2246.600 2393.170 2247.230 ;
        RECT 2397.435 2246.600 2397.695 2247.925 ;
        RECT 2397.985 2246.600 2398.245 2247.925 ;
        RECT 2398.525 2246.600 2398.785 2247.925 ;
        RECT 2399.065 2246.600 2399.305 2247.925 ;
        RECT 2399.605 2246.600 2399.845 2247.925 ;
        RECT 2400.125 2246.600 2400.365 2247.925 ;
        RECT 2400.645 2246.600 2400.885 2247.925 ;
        RECT 2401.165 2246.600 2401.405 2247.925 ;
        RECT 2401.685 2246.600 2401.925 2247.925 ;
        RECT 2402.165 2246.600 2402.405 2247.925 ;
        RECT 2402.645 2246.600 2402.885 2247.925 ;
        RECT 2403.125 2246.600 2403.365 2247.925 ;
        RECT 2403.605 2246.600 2403.845 2247.925 ;
        RECT 2404.085 2246.600 2404.325 2247.925 ;
        RECT 2404.565 2246.600 2404.780 2247.925 ;
        RECT 2405.850 2246.600 2406.020 2247.230 ;
        RECT 2408.595 2246.600 2408.765 2247.230 ;
        RECT 2409.585 2246.600 2409.755 2247.230 ;
        RECT 2414.020 2246.600 2414.280 2247.925 ;
        RECT 2414.570 2246.600 2414.830 2247.925 ;
        RECT 2415.110 2246.600 2415.370 2247.925 ;
        RECT 2415.650 2246.600 2415.890 2247.925 ;
        RECT 2416.190 2246.600 2416.430 2247.925 ;
        RECT 2416.710 2246.600 2416.950 2247.925 ;
        RECT 2417.230 2246.600 2417.470 2247.925 ;
        RECT 2417.750 2246.600 2417.990 2247.925 ;
        RECT 2418.270 2246.600 2418.510 2247.925 ;
        RECT 2418.750 2246.600 2418.990 2247.925 ;
        RECT 2419.230 2246.600 2419.470 2247.925 ;
        RECT 2419.710 2246.600 2419.950 2247.925 ;
        RECT 2420.190 2246.600 2420.430 2247.925 ;
        RECT 2420.670 2246.600 2420.910 2247.925 ;
        RECT 2421.150 2246.600 2421.365 2247.925 ;
        RECT 2422.435 2246.600 2422.605 2247.230 ;
        RECT 2425.180 2246.600 2425.350 2247.230 ;
        RECT 2426.170 2246.600 2426.340 2247.230 ;
        RECT 2430.600 2246.600 2430.860 2247.925 ;
        RECT 2431.150 2246.600 2431.410 2247.925 ;
        RECT 2431.690 2246.600 2431.950 2247.925 ;
        RECT 2432.230 2246.600 2432.470 2247.925 ;
        RECT 2432.770 2246.600 2433.010 2247.925 ;
        RECT 2433.290 2246.600 2433.530 2247.925 ;
        RECT 2433.810 2246.600 2434.050 2247.925 ;
        RECT 2434.330 2246.600 2434.570 2247.925 ;
        RECT 2434.850 2246.600 2435.090 2247.925 ;
        RECT 2435.330 2246.600 2435.570 2247.925 ;
        RECT 2435.810 2246.600 2436.050 2247.925 ;
        RECT 2436.290 2246.600 2436.530 2247.925 ;
        RECT 2436.770 2246.600 2437.010 2247.925 ;
        RECT 2437.250 2246.600 2437.490 2247.925 ;
        RECT 2437.730 2246.600 2437.945 2247.925 ;
        RECT 2439.015 2246.600 2439.185 2247.230 ;
        RECT 2441.760 2246.600 2441.930 2247.230 ;
        RECT 2442.750 2246.600 2442.920 2247.230 ;
        RECT 2343.000 2245.000 2443.725 2246.600 ;
        RECT 2695.520 2216.835 2734.160 2217.005 ;
        RECT 2695.605 2216.085 2696.815 2216.835 ;
        RECT 2697.455 2216.355 2697.730 2216.835 ;
        RECT 2698.315 2216.435 2698.650 2216.835 ;
        RECT 2699.265 2216.455 2699.595 2216.835 ;
        RECT 2700.645 2216.455 2700.975 2216.835 ;
        RECT 2701.585 2216.290 2706.930 2216.835 ;
        RECT 2695.605 2215.545 2696.125 2216.085 ;
        RECT 2703.170 2215.460 2703.510 2216.290 ;
        RECT 2707.105 2216.085 2708.315 2216.835 ;
        RECT 2708.485 2216.110 2708.775 2216.835 ;
        RECT 2709.420 2216.455 2709.750 2216.835 ;
        RECT 2707.105 2215.545 2707.625 2216.085 ;
        RECT 2710.350 2215.995 2710.610 2216.835 ;
        RECT 2710.785 2216.290 2716.130 2216.835 ;
        RECT 2712.370 2215.460 2712.710 2216.290 ;
        RECT 2716.305 2216.065 2719.815 2216.835 ;
        RECT 2719.985 2216.085 2721.195 2216.835 ;
        RECT 2721.365 2216.110 2721.655 2216.835 ;
        RECT 2721.830 2216.435 2722.165 2216.835 ;
        RECT 2722.750 2216.355 2723.025 2216.835 ;
        RECT 2723.665 2216.290 2729.010 2216.835 ;
        RECT 2716.305 2215.545 2717.955 2216.065 ;
        RECT 2719.985 2215.545 2720.505 2216.085 ;
        RECT 2725.250 2215.460 2725.590 2216.290 ;
        RECT 2729.185 2216.065 2730.855 2216.835 ;
        RECT 2731.925 2216.455 2732.255 2216.835 ;
        RECT 2732.865 2216.085 2734.075 2216.835 ;
        RECT 2729.185 2215.545 2729.935 2216.065 ;
        RECT 2733.555 2215.545 2734.075 2216.085 ;
        RECT 2695.605 2212.315 2696.125 2212.855 ;
        RECT 2695.605 2211.565 2696.815 2212.315 ;
        RECT 2699.950 2212.110 2700.290 2212.940 ;
        RECT 2703.885 2212.335 2705.535 2212.855 ;
        RECT 2697.425 2211.565 2697.755 2211.945 ;
        RECT 2698.365 2211.565 2703.710 2212.110 ;
        RECT 2703.885 2211.565 2707.395 2212.335 ;
        RECT 2708.485 2211.565 2708.775 2212.290 ;
        RECT 2710.530 2212.110 2710.870 2212.940 ;
        RECT 2716.050 2212.110 2716.390 2212.940 ;
        RECT 2721.570 2212.110 2721.910 2212.940 ;
        RECT 2727.090 2212.110 2727.430 2212.940 ;
        RECT 2731.025 2212.335 2731.775 2212.855 ;
        RECT 2708.945 2211.565 2714.290 2212.110 ;
        RECT 2714.465 2211.565 2719.810 2212.110 ;
        RECT 2719.985 2211.565 2725.330 2212.110 ;
        RECT 2725.505 2211.565 2730.850 2212.110 ;
        RECT 2731.025 2211.565 2732.695 2212.335 ;
        RECT 2733.555 2212.315 2734.075 2212.855 ;
        RECT 2732.865 2211.565 2734.075 2212.315 ;
        RECT 2695.520 2211.395 2734.160 2211.565 ;
        RECT 2695.605 2210.645 2696.815 2211.395 ;
        RECT 2696.985 2210.850 2702.330 2211.395 ;
        RECT 2702.505 2210.850 2707.850 2211.395 ;
        RECT 2708.025 2210.850 2713.370 2211.395 ;
        RECT 2713.545 2210.850 2718.890 2211.395 ;
        RECT 2695.605 2210.105 2696.125 2210.645 ;
        RECT 2698.570 2210.020 2698.910 2210.850 ;
        RECT 2704.090 2210.020 2704.430 2210.850 ;
        RECT 2709.610 2210.020 2709.950 2210.850 ;
        RECT 2715.130 2210.020 2715.470 2210.850 ;
        RECT 2719.065 2210.625 2720.735 2211.395 ;
        RECT 2721.365 2210.670 2721.655 2211.395 ;
        RECT 2721.825 2210.850 2727.170 2211.395 ;
        RECT 2727.345 2210.850 2732.690 2211.395 ;
        RECT 2719.065 2210.105 2719.815 2210.625 ;
        RECT 2723.410 2210.020 2723.750 2210.850 ;
        RECT 2728.930 2210.020 2729.270 2210.850 ;
        RECT 2732.865 2210.645 2734.075 2211.395 ;
        RECT 2733.555 2210.105 2734.075 2210.645 ;
        RECT 2695.605 2206.875 2696.125 2207.415 ;
        RECT 2695.605 2206.125 2696.815 2206.875 ;
        RECT 2698.570 2206.670 2698.910 2207.500 ;
        RECT 2704.090 2206.670 2704.430 2207.500 ;
        RECT 2696.985 2206.125 2702.330 2206.670 ;
        RECT 2702.505 2206.125 2707.850 2206.670 ;
        RECT 2708.485 2206.125 2708.775 2206.850 ;
        RECT 2710.530 2206.670 2710.870 2207.500 ;
        RECT 2716.050 2206.670 2716.390 2207.500 ;
        RECT 2721.570 2206.670 2721.910 2207.500 ;
        RECT 2727.090 2206.670 2727.430 2207.500 ;
        RECT 2731.025 2206.895 2731.775 2207.415 ;
        RECT 2708.945 2206.125 2714.290 2206.670 ;
        RECT 2714.465 2206.125 2719.810 2206.670 ;
        RECT 2719.985 2206.125 2725.330 2206.670 ;
        RECT 2725.505 2206.125 2730.850 2206.670 ;
        RECT 2731.025 2206.125 2732.695 2206.895 ;
        RECT 2733.555 2206.875 2734.075 2207.415 ;
        RECT 2732.865 2206.125 2734.075 2206.875 ;
        RECT 2695.520 2205.955 2734.160 2206.125 ;
        RECT 2695.605 2205.205 2696.815 2205.955 ;
        RECT 2697.425 2205.575 2697.755 2205.955 ;
        RECT 2698.365 2205.410 2703.710 2205.955 ;
        RECT 2703.885 2205.410 2709.230 2205.955 ;
        RECT 2709.405 2205.410 2714.750 2205.955 ;
        RECT 2714.925 2205.410 2720.270 2205.955 ;
        RECT 2695.605 2204.665 2696.125 2205.205 ;
        RECT 2699.950 2204.580 2700.290 2205.410 ;
        RECT 2705.470 2204.580 2705.810 2205.410 ;
        RECT 2710.990 2204.580 2711.330 2205.410 ;
        RECT 2716.510 2204.580 2716.850 2205.410 ;
        RECT 2721.365 2205.230 2721.655 2205.955 ;
        RECT 2721.825 2205.410 2727.170 2205.955 ;
        RECT 2727.345 2205.410 2732.690 2205.955 ;
        RECT 2723.410 2204.580 2723.750 2205.410 ;
        RECT 2728.930 2204.580 2729.270 2205.410 ;
        RECT 2732.865 2205.205 2734.075 2205.955 ;
        RECT 2733.555 2204.665 2734.075 2205.205 ;
        RECT 2695.605 2201.435 2696.125 2201.975 ;
        RECT 2695.605 2200.685 2696.815 2201.435 ;
        RECT 2698.570 2201.230 2698.910 2202.060 ;
        RECT 2704.090 2201.230 2704.430 2202.060 ;
        RECT 2696.985 2200.685 2702.330 2201.230 ;
        RECT 2702.505 2200.685 2707.850 2201.230 ;
        RECT 2708.485 2200.685 2708.775 2201.410 ;
        RECT 2710.530 2201.230 2710.870 2202.060 ;
        RECT 2716.050 2201.230 2716.390 2202.060 ;
        RECT 2721.570 2201.230 2721.910 2202.060 ;
        RECT 2727.090 2201.230 2727.430 2202.060 ;
        RECT 2731.025 2201.455 2731.775 2201.975 ;
        RECT 2708.945 2200.685 2714.290 2201.230 ;
        RECT 2714.465 2200.685 2719.810 2201.230 ;
        RECT 2719.985 2200.685 2725.330 2201.230 ;
        RECT 2725.505 2200.685 2730.850 2201.230 ;
        RECT 2731.025 2200.685 2732.695 2201.455 ;
        RECT 2733.555 2201.435 2734.075 2201.975 ;
        RECT 2732.865 2200.685 2734.075 2201.435 ;
        RECT 2695.520 2200.515 2734.160 2200.685 ;
        RECT 2695.605 2199.765 2696.815 2200.515 ;
        RECT 2697.415 2200.135 2697.745 2200.515 ;
        RECT 2699.700 2199.795 2699.990 2200.515 ;
        RECT 2702.050 2200.055 2702.220 2200.515 ;
        RECT 2702.910 2200.135 2703.240 2200.515 ;
        RECT 2705.795 2200.055 2705.965 2200.515 ;
        RECT 2706.645 2199.970 2711.990 2200.515 ;
        RECT 2712.165 2199.970 2717.510 2200.515 ;
        RECT 2695.605 2199.225 2696.125 2199.765 ;
        RECT 2708.230 2199.140 2708.570 2199.970 ;
        RECT 2713.750 2199.140 2714.090 2199.970 ;
        RECT 2717.685 2199.745 2721.195 2200.515 ;
        RECT 2721.365 2199.790 2721.655 2200.515 ;
        RECT 2721.825 2199.970 2727.170 2200.515 ;
        RECT 2727.345 2199.970 2732.690 2200.515 ;
        RECT 2717.685 2199.225 2719.335 2199.745 ;
        RECT 2723.410 2199.140 2723.750 2199.970 ;
        RECT 2728.930 2199.140 2729.270 2199.970 ;
        RECT 2732.865 2199.765 2734.075 2200.515 ;
        RECT 2733.555 2199.225 2734.075 2199.765 ;
        RECT 2695.605 2195.995 2696.125 2196.535 ;
        RECT 2695.605 2195.245 2696.815 2195.995 ;
        RECT 2699.950 2195.790 2700.290 2196.620 ;
        RECT 2703.885 2196.015 2705.535 2196.535 ;
        RECT 2697.425 2195.245 2697.755 2195.625 ;
        RECT 2698.365 2195.245 2703.710 2195.790 ;
        RECT 2703.885 2195.245 2707.395 2196.015 ;
        RECT 2708.485 2195.245 2708.775 2195.970 ;
        RECT 2710.530 2195.790 2710.870 2196.620 ;
        RECT 2716.050 2195.790 2716.390 2196.620 ;
        RECT 2721.570 2195.790 2721.910 2196.620 ;
        RECT 2727.090 2195.790 2727.430 2196.620 ;
        RECT 2731.025 2196.015 2731.775 2196.535 ;
        RECT 2708.945 2195.245 2714.290 2195.790 ;
        RECT 2714.465 2195.245 2719.810 2195.790 ;
        RECT 2719.985 2195.245 2725.330 2195.790 ;
        RECT 2725.505 2195.245 2730.850 2195.790 ;
        RECT 2731.025 2195.245 2732.695 2196.015 ;
        RECT 2733.555 2195.995 2734.075 2196.535 ;
        RECT 2732.865 2195.245 2734.075 2195.995 ;
        RECT 2695.520 2195.075 2734.160 2195.245 ;
        RECT 2695.605 2194.325 2696.815 2195.075 ;
        RECT 2697.415 2194.695 2697.745 2195.075 ;
        RECT 2699.700 2194.355 2699.990 2195.075 ;
        RECT 2702.050 2194.615 2702.220 2195.075 ;
        RECT 2702.910 2194.695 2703.240 2195.075 ;
        RECT 2705.795 2194.615 2705.965 2195.075 ;
        RECT 2706.645 2194.530 2711.990 2195.075 ;
        RECT 2712.165 2194.530 2717.510 2195.075 ;
        RECT 2695.605 2193.785 2696.125 2194.325 ;
        RECT 2708.230 2193.700 2708.570 2194.530 ;
        RECT 2713.750 2193.700 2714.090 2194.530 ;
        RECT 2717.685 2194.305 2721.195 2195.075 ;
        RECT 2721.365 2194.350 2721.655 2195.075 ;
        RECT 2721.825 2194.530 2727.170 2195.075 ;
        RECT 2727.345 2194.530 2732.690 2195.075 ;
        RECT 2717.685 2193.785 2719.335 2194.305 ;
        RECT 2723.410 2193.700 2723.750 2194.530 ;
        RECT 2728.930 2193.700 2729.270 2194.530 ;
        RECT 2732.865 2194.325 2734.075 2195.075 ;
        RECT 2733.555 2193.785 2734.075 2194.325 ;
        RECT 2695.605 2190.555 2696.125 2191.095 ;
        RECT 2698.365 2190.575 2699.575 2191.095 ;
        RECT 2705.725 2190.575 2706.935 2191.095 ;
        RECT 2695.605 2189.805 2696.815 2190.555 ;
        RECT 2697.425 2189.805 2697.755 2190.185 ;
        RECT 2698.365 2189.805 2700.955 2190.575 ;
        RECT 2702.015 2189.805 2702.345 2190.205 ;
        RECT 2704.305 2189.805 2704.815 2190.340 ;
        RECT 2705.725 2189.805 2708.315 2190.575 ;
        RECT 2708.485 2189.805 2708.775 2190.530 ;
        RECT 2710.530 2190.350 2710.870 2191.180 ;
        RECT 2716.050 2190.350 2716.390 2191.180 ;
        RECT 2721.570 2190.350 2721.910 2191.180 ;
        RECT 2727.090 2190.350 2727.430 2191.180 ;
        RECT 2731.025 2190.575 2731.775 2191.095 ;
        RECT 2708.945 2189.805 2714.290 2190.350 ;
        RECT 2714.465 2189.805 2719.810 2190.350 ;
        RECT 2719.985 2189.805 2725.330 2190.350 ;
        RECT 2725.505 2189.805 2730.850 2190.350 ;
        RECT 2731.025 2189.805 2732.695 2190.575 ;
        RECT 2733.555 2190.555 2734.075 2191.095 ;
        RECT 2732.865 2189.805 2734.075 2190.555 ;
        RECT 2695.520 2189.635 2734.160 2189.805 ;
        RECT 2695.605 2188.885 2696.815 2189.635 ;
        RECT 2696.985 2189.090 2702.330 2189.635 ;
        RECT 2702.505 2189.090 2707.850 2189.635 ;
        RECT 2708.025 2189.090 2713.370 2189.635 ;
        RECT 2713.545 2189.090 2718.890 2189.635 ;
        RECT 2695.605 2188.345 2696.125 2188.885 ;
        RECT 2698.570 2188.260 2698.910 2189.090 ;
        RECT 2704.090 2188.260 2704.430 2189.090 ;
        RECT 2709.610 2188.260 2709.950 2189.090 ;
        RECT 2715.130 2188.260 2715.470 2189.090 ;
        RECT 2719.065 2188.865 2720.735 2189.635 ;
        RECT 2721.365 2188.910 2721.655 2189.635 ;
        RECT 2721.825 2189.090 2727.170 2189.635 ;
        RECT 2727.345 2189.090 2732.690 2189.635 ;
        RECT 2719.065 2188.345 2719.815 2188.865 ;
        RECT 2723.410 2188.260 2723.750 2189.090 ;
        RECT 2728.930 2188.260 2729.270 2189.090 ;
        RECT 2732.865 2188.885 2734.075 2189.635 ;
        RECT 2733.555 2188.345 2734.075 2188.885 ;
        RECT 2695.605 2185.115 2696.125 2185.655 ;
        RECT 2695.605 2184.365 2696.815 2185.115 ;
        RECT 2699.950 2184.910 2700.290 2185.740 ;
        RECT 2703.885 2185.135 2705.535 2185.655 ;
        RECT 2697.425 2184.365 2697.755 2184.745 ;
        RECT 2698.365 2184.365 2703.710 2184.910 ;
        RECT 2703.885 2184.365 2707.395 2185.135 ;
        RECT 2708.485 2184.365 2708.775 2185.090 ;
        RECT 2710.530 2184.910 2710.870 2185.740 ;
        RECT 2716.050 2184.910 2716.390 2185.740 ;
        RECT 2721.570 2184.910 2721.910 2185.740 ;
        RECT 2727.090 2184.910 2727.430 2185.740 ;
        RECT 2731.025 2185.135 2731.775 2185.655 ;
        RECT 2708.945 2184.365 2714.290 2184.910 ;
        RECT 2714.465 2184.365 2719.810 2184.910 ;
        RECT 2719.985 2184.365 2725.330 2184.910 ;
        RECT 2725.505 2184.365 2730.850 2184.910 ;
        RECT 2731.025 2184.365 2732.695 2185.135 ;
        RECT 2733.555 2185.115 2734.075 2185.655 ;
        RECT 2732.865 2184.365 2734.075 2185.115 ;
        RECT 2695.520 2184.195 2734.160 2184.365 ;
        RECT 2695.605 2183.445 2696.815 2184.195 ;
        RECT 2696.985 2183.650 2702.330 2184.195 ;
        RECT 2702.505 2183.650 2707.850 2184.195 ;
        RECT 2708.025 2183.650 2713.370 2184.195 ;
        RECT 2713.545 2183.650 2718.890 2184.195 ;
        RECT 2695.605 2182.905 2696.125 2183.445 ;
        RECT 2698.570 2182.820 2698.910 2183.650 ;
        RECT 2704.090 2182.820 2704.430 2183.650 ;
        RECT 2709.610 2182.820 2709.950 2183.650 ;
        RECT 2715.130 2182.820 2715.470 2183.650 ;
        RECT 2719.065 2183.425 2720.735 2184.195 ;
        RECT 2721.365 2183.470 2721.655 2184.195 ;
        RECT 2721.825 2183.650 2727.170 2184.195 ;
        RECT 2727.345 2183.650 2732.690 2184.195 ;
        RECT 2719.065 2182.905 2719.815 2183.425 ;
        RECT 2723.410 2182.820 2723.750 2183.650 ;
        RECT 2728.930 2182.820 2729.270 2183.650 ;
        RECT 2732.865 2183.445 2734.075 2184.195 ;
        RECT 2733.555 2182.905 2734.075 2183.445 ;
        RECT 2695.605 2179.675 2696.125 2180.215 ;
        RECT 2696.985 2179.695 2698.635 2180.215 ;
        RECT 2695.605 2178.925 2696.815 2179.675 ;
        RECT 2696.985 2178.925 2700.495 2179.695 ;
        RECT 2701.605 2178.925 2701.845 2179.735 ;
        RECT 2702.515 2178.925 2702.785 2179.735 ;
        RECT 2704.550 2179.470 2704.890 2180.300 ;
        RECT 2702.965 2178.925 2708.310 2179.470 ;
        RECT 2708.485 2178.925 2708.775 2179.650 ;
        RECT 2710.530 2179.470 2710.870 2180.300 ;
        RECT 2716.050 2179.470 2716.390 2180.300 ;
        RECT 2721.570 2179.470 2721.910 2180.300 ;
        RECT 2727.090 2179.470 2727.430 2180.300 ;
        RECT 2731.025 2179.695 2731.775 2180.215 ;
        RECT 2708.945 2178.925 2714.290 2179.470 ;
        RECT 2714.465 2178.925 2719.810 2179.470 ;
        RECT 2719.985 2178.925 2725.330 2179.470 ;
        RECT 2725.505 2178.925 2730.850 2179.470 ;
        RECT 2731.025 2178.925 2732.695 2179.695 ;
        RECT 2733.555 2179.675 2734.075 2180.215 ;
        RECT 2732.865 2178.925 2734.075 2179.675 ;
        RECT 2695.520 2178.755 2734.160 2178.925 ;
        RECT 2695.605 2178.005 2696.815 2178.755 ;
        RECT 2697.425 2178.375 2697.755 2178.755 ;
        RECT 2695.605 2177.465 2696.125 2178.005 ;
        RECT 2698.365 2177.985 2701.875 2178.755 ;
        RECT 2702.055 2178.015 2702.385 2178.755 ;
        RECT 2703.090 2178.395 2703.420 2178.755 ;
        RECT 2698.365 2177.465 2700.015 2177.985 ;
        RECT 2704.785 2177.975 2705.080 2178.755 ;
        RECT 2705.265 2178.210 2710.610 2178.755 ;
        RECT 2710.785 2178.210 2716.130 2178.755 ;
        RECT 2706.850 2177.380 2707.190 2178.210 ;
        RECT 2712.370 2177.380 2712.710 2178.210 ;
        RECT 2716.305 2177.985 2719.815 2178.755 ;
        RECT 2719.985 2178.005 2721.195 2178.755 ;
        RECT 2721.365 2178.030 2721.655 2178.755 ;
        RECT 2721.825 2178.210 2727.170 2178.755 ;
        RECT 2727.345 2178.210 2732.690 2178.755 ;
        RECT 2716.305 2177.465 2717.955 2177.985 ;
        RECT 2719.985 2177.465 2720.505 2178.005 ;
        RECT 2723.410 2177.380 2723.750 2178.210 ;
        RECT 2728.930 2177.380 2729.270 2178.210 ;
        RECT 2732.865 2178.005 2734.075 2178.755 ;
        RECT 2733.555 2177.465 2734.075 2178.005 ;
        RECT 2695.605 2174.235 2696.125 2174.775 ;
        RECT 2695.605 2173.485 2696.815 2174.235 ;
        RECT 2698.570 2174.030 2698.910 2174.860 ;
        RECT 2704.090 2174.030 2704.430 2174.860 ;
        RECT 2696.985 2173.485 2702.330 2174.030 ;
        RECT 2702.505 2173.485 2707.850 2174.030 ;
        RECT 2708.485 2173.485 2708.775 2174.210 ;
        RECT 2710.530 2174.030 2710.870 2174.860 ;
        RECT 2716.050 2174.030 2716.390 2174.860 ;
        RECT 2721.570 2174.030 2721.910 2174.860 ;
        RECT 2708.945 2173.485 2714.290 2174.030 ;
        RECT 2714.465 2173.485 2719.810 2174.030 ;
        RECT 2719.985 2173.485 2725.330 2174.030 ;
        RECT 2725.515 2173.485 2725.845 2173.965 ;
        RECT 2726.355 2173.485 2726.685 2173.965 ;
        RECT 2727.195 2173.485 2727.525 2173.965 ;
        RECT 2728.035 2173.485 2728.365 2173.965 ;
        RECT 2728.875 2173.485 2729.205 2173.965 ;
        RECT 2729.715 2173.485 2730.045 2173.965 ;
        RECT 2730.555 2173.485 2730.885 2173.965 ;
        RECT 2731.395 2173.485 2731.725 2173.965 ;
        RECT 2732.235 2173.485 2732.565 2174.285 ;
        RECT 2733.555 2174.235 2734.075 2174.775 ;
        RECT 2732.865 2173.485 2734.075 2174.235 ;
        RECT 2695.520 2173.315 2734.160 2173.485 ;
        RECT 2695.605 2172.565 2696.815 2173.315 ;
        RECT 2697.425 2172.935 2697.755 2173.315 ;
        RECT 2698.365 2172.770 2703.710 2173.315 ;
        RECT 2703.885 2172.770 2709.230 2173.315 ;
        RECT 2709.405 2172.770 2714.750 2173.315 ;
        RECT 2714.925 2172.770 2720.270 2173.315 ;
        RECT 2695.605 2172.025 2696.125 2172.565 ;
        RECT 2699.950 2171.940 2700.290 2172.770 ;
        RECT 2705.470 2171.940 2705.810 2172.770 ;
        RECT 2710.990 2171.940 2711.330 2172.770 ;
        RECT 2716.510 2171.940 2716.850 2172.770 ;
        RECT 2721.365 2172.590 2721.655 2173.315 ;
        RECT 2721.825 2172.770 2727.170 2173.315 ;
        RECT 2727.345 2172.770 2732.690 2173.315 ;
        RECT 2723.410 2171.940 2723.750 2172.770 ;
        RECT 2728.930 2171.940 2729.270 2172.770 ;
        RECT 2732.865 2172.565 2734.075 2173.315 ;
        RECT 2733.555 2172.025 2734.075 2172.565 ;
        RECT 2695.605 2168.795 2696.125 2169.335 ;
        RECT 2695.605 2168.045 2696.815 2168.795 ;
        RECT 2698.570 2168.590 2698.910 2169.420 ;
        RECT 2704.090 2168.590 2704.430 2169.420 ;
        RECT 2696.985 2168.045 2702.330 2168.590 ;
        RECT 2702.505 2168.045 2707.850 2168.590 ;
        RECT 2708.485 2168.045 2708.775 2168.770 ;
        RECT 2710.530 2168.590 2710.870 2169.420 ;
        RECT 2716.050 2168.590 2716.390 2169.420 ;
        RECT 2721.570 2168.590 2721.910 2169.420 ;
        RECT 2727.090 2168.590 2727.430 2169.420 ;
        RECT 2731.025 2168.815 2731.775 2169.335 ;
        RECT 2708.945 2168.045 2714.290 2168.590 ;
        RECT 2714.465 2168.045 2719.810 2168.590 ;
        RECT 2719.985 2168.045 2725.330 2168.590 ;
        RECT 2725.505 2168.045 2730.850 2168.590 ;
        RECT 2731.025 2168.045 2732.695 2168.815 ;
        RECT 2733.555 2168.795 2734.075 2169.335 ;
        RECT 2732.865 2168.045 2734.075 2168.795 ;
        RECT 2695.520 2167.875 2734.160 2168.045 ;
        RECT 2695.605 2167.125 2696.815 2167.875 ;
        RECT 2697.715 2167.135 2698.045 2167.875 ;
        RECT 2698.555 2167.475 2698.885 2167.875 ;
        RECT 2699.745 2167.330 2705.090 2167.875 ;
        RECT 2705.265 2167.330 2710.610 2167.875 ;
        RECT 2710.785 2167.330 2716.130 2167.875 ;
        RECT 2695.605 2166.585 2696.125 2167.125 ;
        RECT 2701.330 2166.500 2701.670 2167.330 ;
        RECT 2706.850 2166.500 2707.190 2167.330 ;
        RECT 2712.370 2166.500 2712.710 2167.330 ;
        RECT 2716.305 2167.105 2719.815 2167.875 ;
        RECT 2719.985 2167.125 2721.195 2167.875 ;
        RECT 2721.365 2167.150 2721.655 2167.875 ;
        RECT 2721.825 2167.330 2727.170 2167.875 ;
        RECT 2727.345 2167.330 2732.690 2167.875 ;
        RECT 2716.305 2166.585 2717.955 2167.105 ;
        RECT 2719.985 2166.585 2720.505 2167.125 ;
        RECT 2723.410 2166.500 2723.750 2167.330 ;
        RECT 2728.930 2166.500 2729.270 2167.330 ;
        RECT 2732.865 2167.125 2734.075 2167.875 ;
        RECT 2733.555 2166.585 2734.075 2167.125 ;
        RECT 2343.000 2163.860 2446.925 2165.460 ;
        RECT 2358.240 2163.235 2358.410 2163.860 ;
        RECT 2361.480 2163.855 2364.230 2163.860 ;
        RECT 2361.650 2163.225 2361.820 2163.855 ;
        RECT 2362.605 2163.305 2362.775 2163.585 ;
        RECT 2362.605 2163.135 2362.835 2163.305 ;
        RECT 2362.665 2161.525 2362.835 2163.135 ;
        RECT 2362.605 2161.355 2362.835 2161.525 ;
        RECT 2364.610 2161.530 2364.895 2163.860 ;
        RECT 2365.180 2161.530 2365.465 2163.860 ;
        RECT 2365.750 2161.530 2366.035 2163.860 ;
        RECT 2366.320 2161.530 2366.605 2163.860 ;
        RECT 2366.890 2161.530 2367.175 2163.860 ;
        RECT 2367.460 2161.530 2367.745 2163.860 ;
        RECT 2368.030 2161.530 2368.315 2163.860 ;
        RECT 2368.600 2161.530 2368.885 2163.860 ;
        RECT 2369.170 2161.530 2369.450 2163.860 ;
        RECT 2369.735 2161.530 2370.020 2163.860 ;
        RECT 2370.305 2161.530 2370.590 2163.860 ;
        RECT 2370.875 2161.530 2371.160 2163.860 ;
        RECT 2371.730 2161.530 2371.970 2163.860 ;
        RECT 2373.335 2163.235 2373.505 2163.860 ;
        RECT 2376.080 2163.235 2376.250 2163.860 ;
        RECT 2377.070 2163.235 2377.240 2163.860 ;
        RECT 2378.700 2163.855 2381.450 2163.860 ;
        RECT 2378.870 2163.225 2379.040 2163.855 ;
        RECT 2379.825 2163.305 2379.995 2163.585 ;
        RECT 2379.825 2163.135 2380.055 2163.305 ;
        RECT 2364.610 2161.360 2371.970 2161.530 ;
        RECT 2379.885 2161.525 2380.055 2163.135 ;
        RECT 2362.605 2160.295 2362.775 2161.355 ;
        RECT 2365.155 2160.560 2365.465 2161.360 ;
        RECT 2365.165 2160.340 2365.500 2160.390 ;
        RECT 2367.085 2160.340 2367.255 2161.360 ;
        RECT 2367.455 2160.560 2367.765 2161.360 ;
        RECT 2369.735 2160.560 2370.045 2161.360 ;
        RECT 2371.115 2160.560 2371.425 2161.360 ;
        RECT 2379.825 2161.355 2380.055 2161.525 ;
        RECT 2381.830 2161.530 2382.115 2163.860 ;
        RECT 2382.400 2161.530 2382.685 2163.860 ;
        RECT 2382.970 2161.530 2383.255 2163.860 ;
        RECT 2383.540 2161.530 2383.825 2163.860 ;
        RECT 2384.110 2161.530 2384.395 2163.860 ;
        RECT 2384.680 2161.530 2384.965 2163.860 ;
        RECT 2385.250 2161.530 2385.535 2163.860 ;
        RECT 2385.820 2161.530 2386.105 2163.860 ;
        RECT 2386.390 2161.530 2386.670 2163.860 ;
        RECT 2386.955 2161.530 2387.240 2163.860 ;
        RECT 2387.525 2161.530 2387.810 2163.860 ;
        RECT 2388.095 2161.530 2388.380 2163.860 ;
        RECT 2388.950 2161.530 2389.190 2163.860 ;
        RECT 2390.555 2163.235 2390.725 2163.860 ;
        RECT 2393.300 2163.235 2393.470 2163.860 ;
        RECT 2394.290 2163.235 2394.460 2163.860 ;
        RECT 2395.920 2163.855 2398.670 2163.860 ;
        RECT 2396.090 2163.225 2396.260 2163.855 ;
        RECT 2397.045 2163.305 2397.215 2163.585 ;
        RECT 2397.045 2163.135 2397.275 2163.305 ;
        RECT 2381.830 2161.360 2389.190 2161.530 ;
        RECT 2397.105 2161.525 2397.275 2163.135 ;
        RECT 2367.465 2160.340 2367.800 2160.390 ;
        RECT 2364.695 2160.170 2365.500 2160.340 ;
        RECT 2367.075 2160.170 2367.800 2160.340 ;
        RECT 2379.825 2160.295 2379.995 2161.355 ;
        RECT 2382.375 2160.560 2382.685 2161.360 ;
        RECT 2382.385 2160.340 2382.720 2160.390 ;
        RECT 2384.305 2160.340 2384.475 2161.360 ;
        RECT 2384.675 2160.560 2384.985 2161.360 ;
        RECT 2386.955 2160.560 2387.265 2161.360 ;
        RECT 2388.335 2160.560 2388.645 2161.360 ;
        RECT 2397.045 2161.355 2397.275 2161.525 ;
        RECT 2399.050 2161.530 2399.335 2163.860 ;
        RECT 2399.620 2161.530 2399.905 2163.860 ;
        RECT 2400.190 2161.530 2400.475 2163.860 ;
        RECT 2400.760 2161.530 2401.045 2163.860 ;
        RECT 2401.330 2161.530 2401.615 2163.860 ;
        RECT 2401.900 2161.530 2402.185 2163.860 ;
        RECT 2402.470 2161.530 2402.755 2163.860 ;
        RECT 2403.040 2161.530 2403.325 2163.860 ;
        RECT 2403.610 2161.530 2403.890 2163.860 ;
        RECT 2404.175 2161.530 2404.460 2163.860 ;
        RECT 2404.745 2161.530 2405.030 2163.860 ;
        RECT 2405.315 2161.530 2405.600 2163.860 ;
        RECT 2406.170 2161.530 2406.410 2163.860 ;
        RECT 2407.775 2163.235 2407.945 2163.860 ;
        RECT 2410.520 2163.235 2410.690 2163.860 ;
        RECT 2411.510 2163.235 2411.680 2163.860 ;
        RECT 2413.140 2163.855 2415.890 2163.860 ;
        RECT 2413.310 2163.225 2413.480 2163.855 ;
        RECT 2414.265 2163.305 2414.435 2163.585 ;
        RECT 2414.265 2163.135 2414.495 2163.305 ;
        RECT 2399.050 2161.360 2406.410 2161.530 ;
        RECT 2414.325 2161.525 2414.495 2163.135 ;
        RECT 2384.685 2160.340 2385.020 2160.390 ;
        RECT 2381.915 2160.170 2382.720 2160.340 ;
        RECT 2384.295 2160.170 2385.020 2160.340 ;
        RECT 2397.045 2160.295 2397.215 2161.355 ;
        RECT 2399.595 2160.560 2399.905 2161.360 ;
        RECT 2399.605 2160.340 2399.940 2160.390 ;
        RECT 2401.525 2160.340 2401.695 2161.360 ;
        RECT 2401.895 2160.560 2402.205 2161.360 ;
        RECT 2404.175 2160.560 2404.485 2161.360 ;
        RECT 2405.555 2160.560 2405.865 2161.360 ;
        RECT 2414.265 2161.355 2414.495 2161.525 ;
        RECT 2416.270 2161.530 2416.555 2163.860 ;
        RECT 2416.840 2161.530 2417.125 2163.860 ;
        RECT 2417.410 2161.530 2417.695 2163.860 ;
        RECT 2417.980 2161.530 2418.265 2163.860 ;
        RECT 2418.550 2161.530 2418.835 2163.860 ;
        RECT 2419.120 2161.530 2419.405 2163.860 ;
        RECT 2419.690 2161.530 2419.975 2163.860 ;
        RECT 2420.260 2161.530 2420.545 2163.860 ;
        RECT 2420.830 2161.530 2421.110 2163.860 ;
        RECT 2421.395 2161.530 2421.680 2163.860 ;
        RECT 2421.965 2161.530 2422.250 2163.860 ;
        RECT 2422.535 2161.530 2422.820 2163.860 ;
        RECT 2423.390 2161.530 2423.630 2163.860 ;
        RECT 2424.995 2163.235 2425.165 2163.860 ;
        RECT 2427.740 2163.235 2427.910 2163.860 ;
        RECT 2428.730 2163.235 2428.900 2163.860 ;
        RECT 2430.360 2163.855 2433.110 2163.860 ;
        RECT 2430.530 2163.225 2430.700 2163.855 ;
        RECT 2431.485 2163.305 2431.655 2163.585 ;
        RECT 2431.485 2163.135 2431.715 2163.305 ;
        RECT 2416.270 2161.360 2423.630 2161.530 ;
        RECT 2431.545 2161.525 2431.715 2163.135 ;
        RECT 2401.905 2160.340 2402.240 2160.390 ;
        RECT 2399.135 2160.170 2399.940 2160.340 ;
        RECT 2401.515 2160.170 2402.240 2160.340 ;
        RECT 2414.265 2160.295 2414.435 2161.355 ;
        RECT 2416.815 2160.560 2417.125 2161.360 ;
        RECT 2416.825 2160.340 2417.160 2160.390 ;
        RECT 2418.745 2160.340 2418.915 2161.360 ;
        RECT 2419.115 2160.560 2419.425 2161.360 ;
        RECT 2421.395 2160.560 2421.705 2161.360 ;
        RECT 2422.775 2160.560 2423.085 2161.360 ;
        RECT 2431.485 2161.355 2431.715 2161.525 ;
        RECT 2433.490 2161.530 2433.775 2163.860 ;
        RECT 2434.060 2161.530 2434.345 2163.860 ;
        RECT 2434.630 2161.530 2434.915 2163.860 ;
        RECT 2435.200 2161.530 2435.485 2163.860 ;
        RECT 2435.770 2161.530 2436.055 2163.860 ;
        RECT 2436.340 2161.530 2436.625 2163.860 ;
        RECT 2436.910 2161.530 2437.195 2163.860 ;
        RECT 2437.480 2161.530 2437.765 2163.860 ;
        RECT 2438.050 2161.530 2438.330 2163.860 ;
        RECT 2438.615 2161.530 2438.900 2163.860 ;
        RECT 2439.185 2161.530 2439.470 2163.860 ;
        RECT 2439.755 2161.530 2440.040 2163.860 ;
        RECT 2440.610 2161.530 2440.850 2163.860 ;
        RECT 2442.215 2163.235 2442.385 2163.860 ;
        RECT 2444.960 2163.235 2445.130 2163.860 ;
        RECT 2445.950 2163.235 2446.120 2163.860 ;
        RECT 2695.605 2163.355 2696.125 2163.895 ;
        RECT 2695.605 2162.605 2696.815 2163.355 ;
        RECT 2699.950 2163.150 2700.290 2163.980 ;
        RECT 2703.885 2163.375 2705.535 2163.895 ;
        RECT 2697.425 2162.605 2697.755 2162.985 ;
        RECT 2698.365 2162.605 2703.710 2163.150 ;
        RECT 2703.885 2162.605 2707.395 2163.375 ;
        RECT 2708.485 2162.605 2708.775 2163.330 ;
        RECT 2710.530 2163.150 2710.870 2163.980 ;
        RECT 2716.050 2163.150 2716.390 2163.980 ;
        RECT 2721.570 2163.150 2721.910 2163.980 ;
        RECT 2727.090 2163.150 2727.430 2163.980 ;
        RECT 2731.025 2163.375 2731.775 2163.895 ;
        RECT 2708.945 2162.605 2714.290 2163.150 ;
        RECT 2714.465 2162.605 2719.810 2163.150 ;
        RECT 2719.985 2162.605 2725.330 2163.150 ;
        RECT 2725.505 2162.605 2730.850 2163.150 ;
        RECT 2731.025 2162.605 2732.695 2163.375 ;
        RECT 2733.555 2163.355 2734.075 2163.895 ;
        RECT 2732.865 2162.605 2734.075 2163.355 ;
        RECT 2695.520 2162.435 2734.160 2162.605 ;
        RECT 2433.490 2161.360 2440.850 2161.530 ;
        RECT 2695.605 2161.685 2696.815 2162.435 ;
        RECT 2697.725 2161.900 2698.235 2162.435 ;
        RECT 2700.195 2162.035 2700.525 2162.435 ;
        RECT 2701.210 2161.760 2701.450 2162.435 ;
        RECT 2702.840 2161.985 2703.170 2162.435 ;
        RECT 2704.090 2161.995 2704.405 2162.435 ;
        RECT 2704.805 2161.890 2710.150 2162.435 ;
        RECT 2710.325 2161.890 2715.670 2162.435 ;
        RECT 2715.845 2161.890 2721.190 2162.435 ;
        RECT 2419.125 2160.340 2419.460 2160.390 ;
        RECT 2416.355 2160.170 2417.160 2160.340 ;
        RECT 2418.735 2160.170 2419.460 2160.340 ;
        RECT 2431.485 2160.295 2431.655 2161.355 ;
        RECT 2434.035 2160.560 2434.345 2161.360 ;
        RECT 2434.045 2160.340 2434.380 2160.390 ;
        RECT 2435.965 2160.340 2436.135 2161.360 ;
        RECT 2436.335 2160.560 2436.645 2161.360 ;
        RECT 2438.615 2160.560 2438.925 2161.360 ;
        RECT 2439.995 2160.560 2440.305 2161.360 ;
        RECT 2695.605 2161.145 2696.125 2161.685 ;
        RECT 2706.390 2161.060 2706.730 2161.890 ;
        RECT 2711.910 2161.060 2712.250 2161.890 ;
        RECT 2717.430 2161.060 2717.770 2161.890 ;
        RECT 2721.365 2161.710 2721.655 2162.435 ;
        RECT 2721.825 2161.890 2727.170 2162.435 ;
        RECT 2727.345 2161.890 2732.690 2162.435 ;
        RECT 2723.410 2161.060 2723.750 2161.890 ;
        RECT 2728.930 2161.060 2729.270 2161.890 ;
        RECT 2732.865 2161.685 2734.075 2162.435 ;
        RECT 2733.555 2161.145 2734.075 2161.685 ;
        RECT 2436.345 2160.340 2436.680 2160.390 ;
        RECT 2433.575 2160.170 2434.380 2160.340 ;
        RECT 2435.955 2160.170 2436.680 2160.340 ;
        RECT 2365.165 2160.120 2365.500 2160.170 ;
        RECT 2367.465 2160.120 2367.800 2160.170 ;
        RECT 2382.385 2160.120 2382.720 2160.170 ;
        RECT 2384.685 2160.120 2385.020 2160.170 ;
        RECT 2399.605 2160.120 2399.940 2160.170 ;
        RECT 2401.905 2160.120 2402.240 2160.170 ;
        RECT 2416.825 2160.120 2417.160 2160.170 ;
        RECT 2419.125 2160.120 2419.460 2160.170 ;
        RECT 2434.045 2160.120 2434.380 2160.170 ;
        RECT 2436.345 2160.120 2436.680 2160.170 ;
        RECT 2695.605 2157.915 2696.125 2158.455 ;
        RECT 2695.605 2157.165 2696.815 2157.915 ;
        RECT 2696.985 2157.165 2697.245 2157.985 ;
        RECT 2701.790 2157.710 2702.130 2158.540 ;
        RECT 2705.725 2157.935 2706.935 2158.455 ;
        RECT 2699.275 2157.165 2699.605 2157.625 ;
        RECT 2700.205 2157.165 2705.550 2157.710 ;
        RECT 2705.725 2157.165 2708.315 2157.935 ;
        RECT 2708.485 2157.165 2708.775 2157.890 ;
        RECT 2710.530 2157.710 2710.870 2158.540 ;
        RECT 2716.050 2157.710 2716.390 2158.540 ;
        RECT 2721.570 2157.710 2721.910 2158.540 ;
        RECT 2727.090 2157.710 2727.430 2158.540 ;
        RECT 2731.025 2157.935 2731.775 2158.455 ;
        RECT 2708.945 2157.165 2714.290 2157.710 ;
        RECT 2714.465 2157.165 2719.810 2157.710 ;
        RECT 2719.985 2157.165 2725.330 2157.710 ;
        RECT 2725.505 2157.165 2730.850 2157.710 ;
        RECT 2731.025 2157.165 2732.695 2157.935 ;
        RECT 2733.555 2157.915 2734.075 2158.455 ;
        RECT 2732.865 2157.165 2734.075 2157.915 ;
        RECT 2882.265 2157.550 2882.605 2158.210 ;
        RECT 2881.575 2157.380 2883.380 2157.550 ;
        RECT 2695.520 2156.995 2734.160 2157.165 ;
        RECT 2364.755 2156.090 2364.965 2156.910 ;
        RECT 2365.635 2156.090 2365.865 2156.910 ;
        RECT 2366.085 2156.090 2366.355 2156.900 ;
        RECT 2367.025 2156.090 2367.265 2156.900 ;
        RECT 2367.475 2156.090 2367.715 2156.900 ;
        RECT 2368.385 2156.090 2368.655 2156.900 ;
        RECT 2368.835 2156.090 2369.125 2156.925 ;
        RECT 2370.665 2156.090 2370.995 2156.480 ;
        RECT 2371.505 2156.090 2371.835 2156.480 ;
        RECT 2381.975 2156.090 2382.185 2156.910 ;
        RECT 2382.855 2156.090 2383.085 2156.910 ;
        RECT 2383.305 2156.090 2383.575 2156.900 ;
        RECT 2384.245 2156.090 2384.485 2156.900 ;
        RECT 2384.695 2156.090 2384.935 2156.900 ;
        RECT 2385.605 2156.090 2385.875 2156.900 ;
        RECT 2386.055 2156.090 2386.345 2156.925 ;
        RECT 2387.885 2156.090 2388.215 2156.480 ;
        RECT 2388.725 2156.090 2389.055 2156.480 ;
        RECT 2399.195 2156.090 2399.405 2156.910 ;
        RECT 2400.075 2156.090 2400.305 2156.910 ;
        RECT 2400.525 2156.090 2400.795 2156.900 ;
        RECT 2401.465 2156.090 2401.705 2156.900 ;
        RECT 2401.915 2156.090 2402.155 2156.900 ;
        RECT 2402.825 2156.090 2403.095 2156.900 ;
        RECT 2403.275 2156.090 2403.565 2156.925 ;
        RECT 2405.105 2156.090 2405.435 2156.480 ;
        RECT 2405.945 2156.090 2406.275 2156.480 ;
        RECT 2416.415 2156.090 2416.625 2156.910 ;
        RECT 2417.295 2156.090 2417.525 2156.910 ;
        RECT 2417.745 2156.090 2418.015 2156.900 ;
        RECT 2418.685 2156.090 2418.925 2156.900 ;
        RECT 2419.135 2156.090 2419.375 2156.900 ;
        RECT 2420.045 2156.090 2420.315 2156.900 ;
        RECT 2420.495 2156.090 2420.785 2156.925 ;
        RECT 2422.325 2156.090 2422.655 2156.480 ;
        RECT 2423.165 2156.090 2423.495 2156.480 ;
        RECT 2433.635 2156.090 2433.845 2156.910 ;
        RECT 2434.515 2156.090 2434.745 2156.910 ;
        RECT 2434.965 2156.090 2435.235 2156.900 ;
        RECT 2435.905 2156.090 2436.145 2156.900 ;
        RECT 2436.355 2156.090 2436.595 2156.900 ;
        RECT 2437.265 2156.090 2437.535 2156.900 ;
        RECT 2437.715 2156.090 2438.005 2156.925 ;
        RECT 2439.545 2156.090 2439.875 2156.480 ;
        RECT 2440.385 2156.090 2440.715 2156.480 ;
        RECT 2695.605 2156.245 2696.815 2156.995 ;
        RECT 2697.425 2156.615 2697.755 2156.995 ;
        RECT 2698.365 2156.450 2703.710 2156.995 ;
        RECT 2703.885 2156.450 2709.230 2156.995 ;
        RECT 2709.405 2156.450 2714.750 2156.995 ;
        RECT 2714.925 2156.450 2720.270 2156.995 ;
        RECT 2364.605 2155.920 2372.265 2156.090 ;
        RECT 2364.605 2154.605 2364.885 2155.920 ;
        RECT 2365.170 2154.605 2365.455 2155.920 ;
        RECT 2365.740 2154.605 2366.025 2155.920 ;
        RECT 2366.310 2154.605 2366.595 2155.920 ;
        RECT 2366.880 2154.605 2367.165 2155.920 ;
        RECT 2367.450 2154.605 2367.735 2155.920 ;
        RECT 2368.020 2154.605 2368.305 2155.920 ;
        RECT 2368.590 2154.605 2368.875 2155.920 ;
        RECT 2369.160 2154.605 2369.445 2155.920 ;
        RECT 2369.730 2154.605 2370.015 2155.920 ;
        RECT 2370.300 2154.605 2370.585 2155.920 ;
        RECT 2370.870 2154.605 2371.155 2155.920 ;
        RECT 2371.440 2154.605 2371.725 2155.920 ;
        RECT 2372.010 2154.605 2372.265 2155.920 ;
        RECT 2381.825 2155.920 2389.485 2156.090 ;
        RECT 2364.605 2154.600 2372.265 2154.605 ;
        RECT 2373.335 2154.600 2373.505 2155.225 ;
        RECT 2376.080 2154.600 2376.250 2155.225 ;
        RECT 2377.065 2154.600 2377.235 2155.225 ;
        RECT 2381.825 2154.605 2382.105 2155.920 ;
        RECT 2382.390 2154.605 2382.675 2155.920 ;
        RECT 2382.960 2154.605 2383.245 2155.920 ;
        RECT 2383.530 2154.605 2383.815 2155.920 ;
        RECT 2384.100 2154.605 2384.385 2155.920 ;
        RECT 2384.670 2154.605 2384.955 2155.920 ;
        RECT 2385.240 2154.605 2385.525 2155.920 ;
        RECT 2385.810 2154.605 2386.095 2155.920 ;
        RECT 2386.380 2154.605 2386.665 2155.920 ;
        RECT 2386.950 2154.605 2387.235 2155.920 ;
        RECT 2387.520 2154.605 2387.805 2155.920 ;
        RECT 2388.090 2154.605 2388.375 2155.920 ;
        RECT 2388.660 2154.605 2388.945 2155.920 ;
        RECT 2389.230 2154.605 2389.485 2155.920 ;
        RECT 2399.045 2155.920 2406.705 2156.090 ;
        RECT 2381.825 2154.600 2389.485 2154.605 ;
        RECT 2390.555 2154.600 2390.725 2155.225 ;
        RECT 2393.300 2154.600 2393.470 2155.225 ;
        RECT 2394.285 2154.600 2394.455 2155.225 ;
        RECT 2399.045 2154.605 2399.325 2155.920 ;
        RECT 2399.610 2154.605 2399.895 2155.920 ;
        RECT 2400.180 2154.605 2400.465 2155.920 ;
        RECT 2400.750 2154.605 2401.035 2155.920 ;
        RECT 2401.320 2154.605 2401.605 2155.920 ;
        RECT 2401.890 2154.605 2402.175 2155.920 ;
        RECT 2402.460 2154.605 2402.745 2155.920 ;
        RECT 2403.030 2154.605 2403.315 2155.920 ;
        RECT 2403.600 2154.605 2403.885 2155.920 ;
        RECT 2404.170 2154.605 2404.455 2155.920 ;
        RECT 2404.740 2154.605 2405.025 2155.920 ;
        RECT 2405.310 2154.605 2405.595 2155.920 ;
        RECT 2405.880 2154.605 2406.165 2155.920 ;
        RECT 2406.450 2154.605 2406.705 2155.920 ;
        RECT 2416.265 2155.920 2423.925 2156.090 ;
        RECT 2399.045 2154.600 2406.705 2154.605 ;
        RECT 2407.775 2154.600 2407.945 2155.225 ;
        RECT 2410.520 2154.600 2410.690 2155.225 ;
        RECT 2411.505 2154.600 2411.675 2155.225 ;
        RECT 2416.265 2154.605 2416.545 2155.920 ;
        RECT 2416.830 2154.605 2417.115 2155.920 ;
        RECT 2417.400 2154.605 2417.685 2155.920 ;
        RECT 2417.970 2154.605 2418.255 2155.920 ;
        RECT 2418.540 2154.605 2418.825 2155.920 ;
        RECT 2419.110 2154.605 2419.395 2155.920 ;
        RECT 2419.680 2154.605 2419.965 2155.920 ;
        RECT 2420.250 2154.605 2420.535 2155.920 ;
        RECT 2420.820 2154.605 2421.105 2155.920 ;
        RECT 2421.390 2154.605 2421.675 2155.920 ;
        RECT 2421.960 2154.605 2422.245 2155.920 ;
        RECT 2422.530 2154.605 2422.815 2155.920 ;
        RECT 2423.100 2154.605 2423.385 2155.920 ;
        RECT 2423.670 2154.605 2423.925 2155.920 ;
        RECT 2433.485 2155.920 2441.145 2156.090 ;
        RECT 2416.265 2154.600 2423.925 2154.605 ;
        RECT 2424.995 2154.600 2425.165 2155.225 ;
        RECT 2427.740 2154.600 2427.910 2155.225 ;
        RECT 2428.725 2154.600 2428.895 2155.225 ;
        RECT 2433.485 2154.605 2433.765 2155.920 ;
        RECT 2434.050 2154.605 2434.335 2155.920 ;
        RECT 2434.620 2154.605 2434.905 2155.920 ;
        RECT 2435.190 2154.605 2435.475 2155.920 ;
        RECT 2435.760 2154.605 2436.045 2155.920 ;
        RECT 2436.330 2154.605 2436.615 2155.920 ;
        RECT 2436.900 2154.605 2437.185 2155.920 ;
        RECT 2437.470 2154.605 2437.755 2155.920 ;
        RECT 2438.040 2154.605 2438.325 2155.920 ;
        RECT 2438.610 2154.605 2438.895 2155.920 ;
        RECT 2439.180 2154.605 2439.465 2155.920 ;
        RECT 2439.750 2154.605 2440.035 2155.920 ;
        RECT 2440.320 2154.605 2440.605 2155.920 ;
        RECT 2440.890 2154.605 2441.145 2155.920 ;
        RECT 2695.605 2155.705 2696.125 2156.245 ;
        RECT 2699.950 2155.620 2700.290 2156.450 ;
        RECT 2705.470 2155.620 2705.810 2156.450 ;
        RECT 2710.990 2155.620 2711.330 2156.450 ;
        RECT 2716.510 2155.620 2716.850 2156.450 ;
        RECT 2721.365 2156.270 2721.655 2156.995 ;
        RECT 2721.825 2156.450 2727.170 2156.995 ;
        RECT 2727.345 2156.450 2732.690 2156.995 ;
        RECT 2723.410 2155.620 2723.750 2156.450 ;
        RECT 2728.930 2155.620 2729.270 2156.450 ;
        RECT 2732.865 2156.245 2734.075 2156.995 ;
        RECT 2733.555 2155.705 2734.075 2156.245 ;
        RECT 2433.485 2154.600 2441.145 2154.605 ;
        RECT 2442.215 2154.600 2442.385 2155.225 ;
        RECT 2444.960 2154.600 2445.130 2155.225 ;
        RECT 2445.945 2154.600 2446.115 2155.225 ;
        RECT 2343.015 2153.000 2446.925 2154.600 ;
        RECT 2695.605 2152.475 2696.125 2153.015 ;
        RECT 2696.985 2152.475 2697.505 2153.015 ;
        RECT 2695.605 2151.725 2696.815 2152.475 ;
        RECT 2696.985 2151.725 2698.195 2152.475 ;
        RECT 2698.365 2151.725 2698.705 2152.450 ;
        RECT 2703.630 2152.270 2703.970 2153.100 ;
        RECT 2701.035 2151.725 2701.365 2152.205 ;
        RECT 2702.045 2151.725 2707.390 2152.270 ;
        RECT 2708.485 2151.725 2708.775 2152.450 ;
        RECT 2710.530 2152.270 2710.870 2153.100 ;
        RECT 2716.050 2152.270 2716.390 2153.100 ;
        RECT 2721.570 2152.270 2721.910 2153.100 ;
        RECT 2727.090 2152.270 2727.430 2153.100 ;
        RECT 2731.025 2152.495 2731.775 2153.015 ;
        RECT 2708.945 2151.725 2714.290 2152.270 ;
        RECT 2714.465 2151.725 2719.810 2152.270 ;
        RECT 2719.985 2151.725 2725.330 2152.270 ;
        RECT 2725.505 2151.725 2730.850 2152.270 ;
        RECT 2731.025 2151.725 2732.695 2152.495 ;
        RECT 2733.555 2152.475 2734.075 2153.015 ;
        RECT 2732.865 2151.725 2734.075 2152.475 ;
        RECT 2695.520 2151.555 2734.160 2151.725 ;
        RECT 2695.605 2150.805 2696.815 2151.555 ;
        RECT 2695.605 2150.265 2696.125 2150.805 ;
        RECT 2697.905 2150.735 2698.165 2151.555 ;
        RECT 2699.275 2151.155 2699.605 2151.555 ;
        RECT 2700.115 2151.155 2700.490 2151.555 ;
        RECT 2702.760 2151.155 2703.090 2151.555 ;
        RECT 2703.885 2151.010 2709.230 2151.555 ;
        RECT 2709.405 2151.010 2714.750 2151.555 ;
        RECT 2714.925 2151.010 2720.270 2151.555 ;
        RECT 2705.470 2150.180 2705.810 2151.010 ;
        RECT 2710.990 2150.180 2711.330 2151.010 ;
        RECT 2716.510 2150.180 2716.850 2151.010 ;
        RECT 2721.365 2150.830 2721.655 2151.555 ;
        RECT 2721.825 2151.010 2727.170 2151.555 ;
        RECT 2727.345 2151.010 2732.690 2151.555 ;
        RECT 2723.410 2150.180 2723.750 2151.010 ;
        RECT 2728.930 2150.180 2729.270 2151.010 ;
        RECT 2732.865 2150.805 2734.075 2151.555 ;
        RECT 2733.555 2150.265 2734.075 2150.805 ;
        RECT 2695.605 2147.035 2696.125 2147.575 ;
        RECT 2695.605 2146.285 2696.815 2147.035 ;
        RECT 2697.425 2146.285 2697.755 2146.665 ;
        RECT 2699.725 2146.285 2700.035 2147.085 ;
        RECT 2701.790 2146.830 2702.130 2147.660 ;
        RECT 2705.725 2147.055 2706.935 2147.575 ;
        RECT 2700.205 2146.285 2705.550 2146.830 ;
        RECT 2705.725 2146.285 2708.315 2147.055 ;
        RECT 2708.485 2146.285 2708.775 2147.010 ;
        RECT 2710.530 2146.830 2710.870 2147.660 ;
        RECT 2716.050 2146.830 2716.390 2147.660 ;
        RECT 2721.570 2146.830 2721.910 2147.660 ;
        RECT 2727.090 2146.830 2727.430 2147.660 ;
        RECT 2731.025 2147.055 2731.775 2147.575 ;
        RECT 2708.945 2146.285 2714.290 2146.830 ;
        RECT 2714.465 2146.285 2719.810 2146.830 ;
        RECT 2719.985 2146.285 2725.330 2146.830 ;
        RECT 2725.505 2146.285 2730.850 2146.830 ;
        RECT 2731.025 2146.285 2732.695 2147.055 ;
        RECT 2733.555 2147.035 2734.075 2147.575 ;
        RECT 2732.865 2146.285 2734.075 2147.035 ;
        RECT 2695.520 2146.115 2734.160 2146.285 ;
        RECT 2695.605 2145.365 2696.815 2146.115 ;
        RECT 2697.725 2145.580 2698.235 2146.115 ;
        RECT 2700.195 2145.715 2700.525 2146.115 ;
        RECT 2701.125 2145.570 2706.470 2146.115 ;
        RECT 2706.645 2145.570 2711.990 2146.115 ;
        RECT 2712.165 2145.570 2717.510 2146.115 ;
        RECT 2695.605 2144.825 2696.125 2145.365 ;
        RECT 2702.710 2144.740 2703.050 2145.570 ;
        RECT 2708.230 2144.740 2708.570 2145.570 ;
        RECT 2713.750 2144.740 2714.090 2145.570 ;
        RECT 2717.685 2145.345 2721.195 2146.115 ;
        RECT 2721.365 2145.390 2721.655 2146.115 ;
        RECT 2721.825 2145.570 2727.170 2146.115 ;
        RECT 2727.345 2145.570 2732.690 2146.115 ;
        RECT 2717.685 2144.825 2719.335 2145.345 ;
        RECT 2723.410 2144.740 2723.750 2145.570 ;
        RECT 2728.930 2144.740 2729.270 2145.570 ;
        RECT 2732.865 2145.365 2734.075 2146.115 ;
        RECT 2733.555 2144.825 2734.075 2145.365 ;
        RECT 2695.605 2141.595 2696.125 2142.135 ;
        RECT 2695.605 2140.845 2696.815 2141.595 ;
        RECT 2699.950 2141.390 2700.290 2142.220 ;
        RECT 2703.885 2141.615 2705.535 2142.135 ;
        RECT 2697.425 2140.845 2697.755 2141.225 ;
        RECT 2698.365 2140.845 2703.710 2141.390 ;
        RECT 2703.885 2140.845 2707.395 2141.615 ;
        RECT 2708.485 2140.845 2708.775 2141.570 ;
        RECT 2710.530 2141.390 2710.870 2142.220 ;
        RECT 2716.050 2141.390 2716.390 2142.220 ;
        RECT 2721.570 2141.390 2721.910 2142.220 ;
        RECT 2727.090 2141.390 2727.430 2142.220 ;
        RECT 2731.025 2141.615 2731.775 2142.135 ;
        RECT 2708.945 2140.845 2714.290 2141.390 ;
        RECT 2714.465 2140.845 2719.810 2141.390 ;
        RECT 2719.985 2140.845 2725.330 2141.390 ;
        RECT 2725.505 2140.845 2730.850 2141.390 ;
        RECT 2731.025 2140.845 2732.695 2141.615 ;
        RECT 2733.555 2141.595 2734.075 2142.135 ;
        RECT 2732.865 2140.845 2734.075 2141.595 ;
        RECT 2695.520 2140.675 2734.160 2140.845 ;
        RECT 2695.605 2139.925 2696.815 2140.675 ;
        RECT 2696.985 2140.130 2702.330 2140.675 ;
        RECT 2702.505 2140.130 2707.850 2140.675 ;
        RECT 2708.025 2140.130 2713.370 2140.675 ;
        RECT 2713.545 2140.130 2718.890 2140.675 ;
        RECT 2695.605 2139.385 2696.125 2139.925 ;
        RECT 2698.570 2139.300 2698.910 2140.130 ;
        RECT 2704.090 2139.300 2704.430 2140.130 ;
        RECT 2709.610 2139.300 2709.950 2140.130 ;
        RECT 2715.130 2139.300 2715.470 2140.130 ;
        RECT 2719.065 2139.905 2720.735 2140.675 ;
        RECT 2721.365 2139.950 2721.655 2140.675 ;
        RECT 2721.825 2140.130 2727.170 2140.675 ;
        RECT 2727.345 2140.130 2732.690 2140.675 ;
        RECT 2719.065 2139.385 2719.815 2139.905 ;
        RECT 2723.410 2139.300 2723.750 2140.130 ;
        RECT 2728.930 2139.300 2729.270 2140.130 ;
        RECT 2732.865 2139.925 2734.075 2140.675 ;
        RECT 2733.555 2139.385 2734.075 2139.925 ;
        RECT 2695.605 2136.155 2696.125 2136.695 ;
        RECT 2695.605 2135.405 2696.815 2136.155 ;
        RECT 2699.950 2135.950 2700.290 2136.780 ;
        RECT 2703.885 2136.175 2705.535 2136.695 ;
        RECT 2697.425 2135.405 2697.755 2135.785 ;
        RECT 2698.365 2135.405 2703.710 2135.950 ;
        RECT 2703.885 2135.405 2707.395 2136.175 ;
        RECT 2708.485 2135.405 2708.775 2136.130 ;
        RECT 2710.530 2135.950 2710.870 2136.780 ;
        RECT 2716.050 2135.950 2716.390 2136.780 ;
        RECT 2721.570 2135.950 2721.910 2136.780 ;
        RECT 2727.090 2135.950 2727.430 2136.780 ;
        RECT 2731.025 2136.175 2731.775 2136.695 ;
        RECT 2708.945 2135.405 2714.290 2135.950 ;
        RECT 2714.465 2135.405 2719.810 2135.950 ;
        RECT 2719.985 2135.405 2725.330 2135.950 ;
        RECT 2725.505 2135.405 2730.850 2135.950 ;
        RECT 2731.025 2135.405 2732.695 2136.175 ;
        RECT 2733.555 2136.155 2734.075 2136.695 ;
        RECT 2732.865 2135.405 2734.075 2136.155 ;
        RECT 2695.520 2135.235 2734.160 2135.405 ;
        RECT 2523.330 2134.040 2523.670 2134.700 ;
        RECT 2695.605 2134.485 2696.815 2135.235 ;
        RECT 2696.985 2134.690 2702.330 2135.235 ;
        RECT 2702.505 2134.690 2707.850 2135.235 ;
        RECT 2708.025 2134.690 2713.370 2135.235 ;
        RECT 2713.545 2134.690 2718.890 2135.235 ;
        RECT 2522.130 2133.870 2523.935 2134.040 ;
        RECT 2695.605 2133.945 2696.125 2134.485 ;
        RECT 2698.570 2133.860 2698.910 2134.690 ;
        RECT 2704.090 2133.860 2704.430 2134.690 ;
        RECT 2709.610 2133.860 2709.950 2134.690 ;
        RECT 2715.130 2133.860 2715.470 2134.690 ;
        RECT 2719.065 2134.465 2720.735 2135.235 ;
        RECT 2721.365 2134.510 2721.655 2135.235 ;
        RECT 2721.825 2134.690 2727.170 2135.235 ;
        RECT 2727.345 2134.690 2732.690 2135.235 ;
        RECT 2719.065 2133.945 2719.815 2134.465 ;
        RECT 2723.410 2133.860 2723.750 2134.690 ;
        RECT 2728.930 2133.860 2729.270 2134.690 ;
        RECT 2732.865 2134.485 2734.075 2135.235 ;
        RECT 2733.555 2133.945 2734.075 2134.485 ;
        RECT 2695.605 2130.715 2696.125 2131.255 ;
        RECT 2695.605 2129.965 2696.815 2130.715 ;
        RECT 2701.330 2130.510 2701.670 2131.340 ;
        RECT 2705.265 2130.735 2706.475 2131.255 ;
        RECT 2697.425 2129.965 2697.755 2130.345 ;
        RECT 2698.805 2129.965 2699.135 2130.345 ;
        RECT 2699.745 2129.965 2705.090 2130.510 ;
        RECT 2705.265 2129.965 2707.855 2130.735 ;
        RECT 2708.485 2129.965 2708.775 2130.690 ;
        RECT 2710.530 2130.510 2710.870 2131.340 ;
        RECT 2716.050 2130.510 2716.390 2131.340 ;
        RECT 2719.985 2130.715 2720.505 2131.255 ;
        RECT 2708.945 2129.965 2714.290 2130.510 ;
        RECT 2714.465 2129.965 2719.810 2130.510 ;
        RECT 2719.985 2129.965 2721.195 2130.715 ;
        RECT 2721.365 2129.965 2721.655 2130.690 ;
        RECT 2723.410 2130.510 2723.750 2131.340 ;
        RECT 2728.930 2130.510 2729.270 2131.340 ;
        RECT 2733.555 2130.715 2734.075 2131.255 ;
        RECT 2721.825 2129.965 2727.170 2130.510 ;
        RECT 2727.345 2129.965 2732.690 2130.510 ;
        RECT 2732.865 2129.965 2734.075 2130.715 ;
        RECT 2695.520 2129.795 2734.160 2129.965 ;
        RECT 2523.330 2126.510 2523.670 2127.170 ;
        RECT 2522.130 2126.340 2523.935 2126.510 ;
        RECT 2523.330 2120.530 2523.670 2121.190 ;
        RECT 2522.130 2120.360 2523.935 2120.530 ;
        RECT 2523.330 2114.585 2523.670 2115.245 ;
        RECT 2522.130 2114.415 2523.935 2114.585 ;
        RECT 2523.330 2108.940 2523.670 2109.600 ;
        RECT 2522.130 2108.770 2523.935 2108.940 ;
        RECT 2523.330 2102.935 2523.670 2103.595 ;
        RECT 2522.130 2102.765 2523.935 2102.935 ;
        RECT 2343.050 2058.860 2442.430 2060.460 ;
        RECT 2358.220 2058.235 2358.390 2058.860 ;
        RECT 2366.800 2058.235 2366.970 2058.860 ;
        RECT 2367.755 2058.315 2367.925 2058.595 ;
        RECT 2367.755 2058.145 2367.985 2058.315 ;
        RECT 2372.415 2058.235 2372.585 2058.860 ;
        RECT 2375.160 2058.235 2375.330 2058.860 ;
        RECT 2376.155 2058.230 2376.325 2058.860 ;
        RECT 2383.125 2058.235 2383.295 2058.860 ;
        RECT 2384.080 2058.315 2384.250 2058.595 ;
        RECT 2384.080 2058.145 2384.310 2058.315 ;
        RECT 2388.740 2058.235 2388.910 2058.860 ;
        RECT 2391.485 2058.235 2391.655 2058.860 ;
        RECT 2392.480 2058.230 2392.650 2058.860 ;
        RECT 2399.450 2058.235 2399.620 2058.860 ;
        RECT 2400.405 2058.315 2400.575 2058.595 ;
        RECT 2400.405 2058.145 2400.635 2058.315 ;
        RECT 2405.065 2058.235 2405.235 2058.860 ;
        RECT 2407.810 2058.235 2407.980 2058.860 ;
        RECT 2408.805 2058.230 2408.975 2058.860 ;
        RECT 2415.775 2058.235 2415.945 2058.860 ;
        RECT 2416.730 2058.315 2416.900 2058.595 ;
        RECT 2416.730 2058.145 2416.960 2058.315 ;
        RECT 2421.390 2058.235 2421.560 2058.860 ;
        RECT 2424.135 2058.235 2424.305 2058.860 ;
        RECT 2425.130 2058.230 2425.300 2058.860 ;
        RECT 2432.100 2058.235 2432.270 2058.860 ;
        RECT 2433.055 2058.315 2433.225 2058.595 ;
        RECT 2433.055 2058.145 2433.285 2058.315 ;
        RECT 2437.715 2058.235 2437.885 2058.860 ;
        RECT 2440.460 2058.235 2440.630 2058.860 ;
        RECT 2441.455 2058.230 2441.625 2058.860 ;
        RECT 2367.815 2056.535 2367.985 2058.145 ;
        RECT 2384.140 2056.535 2384.310 2058.145 ;
        RECT 2400.465 2056.535 2400.635 2058.145 ;
        RECT 2416.790 2056.535 2416.960 2058.145 ;
        RECT 2433.115 2056.535 2433.285 2058.145 ;
        RECT 2367.755 2056.365 2367.985 2056.535 ;
        RECT 2384.080 2056.365 2384.310 2056.535 ;
        RECT 2400.405 2056.365 2400.635 2056.535 ;
        RECT 2416.730 2056.365 2416.960 2056.535 ;
        RECT 2433.055 2056.365 2433.285 2056.535 ;
        RECT 2367.755 2055.305 2367.925 2056.365 ;
        RECT 2384.080 2055.305 2384.250 2056.365 ;
        RECT 2400.405 2055.305 2400.575 2056.365 ;
        RECT 2416.730 2055.305 2416.900 2056.365 ;
        RECT 2433.055 2055.305 2433.225 2056.365 ;
        RECT 2368.670 2052.035 2368.840 2052.235 ;
        RECT 2370.630 2052.035 2370.800 2052.235 ;
        RECT 2384.995 2052.035 2385.165 2052.235 ;
        RECT 2386.955 2052.035 2387.125 2052.235 ;
        RECT 2401.320 2052.035 2401.490 2052.235 ;
        RECT 2403.280 2052.035 2403.450 2052.235 ;
        RECT 2417.645 2052.035 2417.815 2052.235 ;
        RECT 2419.605 2052.035 2419.775 2052.235 ;
        RECT 2433.970 2052.035 2434.140 2052.235 ;
        RECT 2435.930 2052.035 2436.100 2052.235 ;
        RECT 2368.350 2051.865 2368.840 2052.035 ;
        RECT 2370.310 2051.865 2370.800 2052.035 ;
        RECT 2384.675 2051.865 2385.165 2052.035 ;
        RECT 2386.635 2051.865 2387.125 2052.035 ;
        RECT 2401.000 2051.865 2401.490 2052.035 ;
        RECT 2402.960 2051.865 2403.450 2052.035 ;
        RECT 2417.325 2051.865 2417.815 2052.035 ;
        RECT 2419.285 2051.865 2419.775 2052.035 ;
        RECT 2433.650 2051.865 2434.140 2052.035 ;
        RECT 2435.610 2051.865 2436.100 2052.035 ;
        RECT 2361.870 2050.890 2362.040 2051.375 ;
        RECT 2361.665 2050.875 2362.040 2050.890 ;
        RECT 2362.830 2050.875 2363.000 2051.375 ;
        RECT 2363.790 2050.890 2363.960 2051.375 ;
        RECT 2364.310 2050.890 2364.480 2051.375 ;
        RECT 2363.790 2050.875 2364.480 2050.890 ;
        RECT 2365.270 2050.875 2365.440 2051.375 ;
        RECT 2367.710 2050.890 2367.880 2051.375 ;
        RECT 2366.090 2050.875 2366.285 2050.890 ;
        RECT 2367.640 2050.875 2367.880 2050.890 ;
        RECT 2369.670 2050.875 2369.840 2051.375 ;
        RECT 2378.195 2050.890 2378.365 2051.375 ;
        RECT 2371.165 2050.875 2371.355 2050.880 ;
        RECT 2377.990 2050.875 2378.365 2050.890 ;
        RECT 2379.155 2050.875 2379.325 2051.375 ;
        RECT 2380.115 2050.890 2380.285 2051.375 ;
        RECT 2380.635 2050.890 2380.805 2051.375 ;
        RECT 2380.115 2050.875 2380.805 2050.890 ;
        RECT 2381.595 2050.875 2381.765 2051.375 ;
        RECT 2384.035 2050.890 2384.205 2051.375 ;
        RECT 2382.415 2050.875 2382.610 2050.890 ;
        RECT 2383.965 2050.875 2384.205 2050.890 ;
        RECT 2385.995 2050.875 2386.165 2051.375 ;
        RECT 2394.520 2050.890 2394.690 2051.375 ;
        RECT 2387.490 2050.875 2387.680 2050.880 ;
        RECT 2394.315 2050.875 2394.690 2050.890 ;
        RECT 2395.480 2050.875 2395.650 2051.375 ;
        RECT 2396.440 2050.890 2396.610 2051.375 ;
        RECT 2396.960 2050.890 2397.130 2051.375 ;
        RECT 2396.440 2050.875 2397.130 2050.890 ;
        RECT 2397.920 2050.875 2398.090 2051.375 ;
        RECT 2400.360 2050.890 2400.530 2051.375 ;
        RECT 2398.740 2050.875 2398.935 2050.890 ;
        RECT 2400.290 2050.875 2400.530 2050.890 ;
        RECT 2402.320 2050.875 2402.490 2051.375 ;
        RECT 2410.845 2050.890 2411.015 2051.375 ;
        RECT 2403.815 2050.875 2404.005 2050.880 ;
        RECT 2410.640 2050.875 2411.015 2050.890 ;
        RECT 2411.805 2050.875 2411.975 2051.375 ;
        RECT 2412.765 2050.890 2412.935 2051.375 ;
        RECT 2413.285 2050.890 2413.455 2051.375 ;
        RECT 2412.765 2050.875 2413.455 2050.890 ;
        RECT 2414.245 2050.875 2414.415 2051.375 ;
        RECT 2416.685 2050.890 2416.855 2051.375 ;
        RECT 2415.065 2050.875 2415.260 2050.890 ;
        RECT 2416.615 2050.875 2416.855 2050.890 ;
        RECT 2418.645 2050.875 2418.815 2051.375 ;
        RECT 2427.170 2050.890 2427.340 2051.375 ;
        RECT 2420.140 2050.875 2420.330 2050.880 ;
        RECT 2426.965 2050.875 2427.340 2050.890 ;
        RECT 2428.130 2050.875 2428.300 2051.375 ;
        RECT 2429.090 2050.890 2429.260 2051.375 ;
        RECT 2429.610 2050.890 2429.780 2051.375 ;
        RECT 2429.090 2050.875 2429.780 2050.890 ;
        RECT 2430.570 2050.875 2430.740 2051.375 ;
        RECT 2433.010 2050.890 2433.180 2051.375 ;
        RECT 2431.390 2050.875 2431.585 2050.890 ;
        RECT 2432.940 2050.875 2433.180 2050.890 ;
        RECT 2434.970 2050.875 2435.140 2051.375 ;
        RECT 2436.465 2050.875 2436.655 2050.880 ;
        RECT 2361.540 2049.600 2371.355 2050.875 ;
        RECT 2372.415 2049.600 2372.585 2050.225 ;
        RECT 2375.160 2049.600 2375.330 2050.225 ;
        RECT 2376.150 2049.600 2376.320 2050.230 ;
        RECT 2377.865 2049.600 2387.680 2050.875 ;
        RECT 2388.740 2049.600 2388.910 2050.225 ;
        RECT 2391.485 2049.600 2391.655 2050.225 ;
        RECT 2392.475 2049.600 2392.645 2050.230 ;
        RECT 2394.190 2049.600 2404.005 2050.875 ;
        RECT 2405.065 2049.600 2405.235 2050.225 ;
        RECT 2407.810 2049.600 2407.980 2050.225 ;
        RECT 2408.800 2049.600 2408.970 2050.230 ;
        RECT 2410.515 2049.600 2420.330 2050.875 ;
        RECT 2421.390 2049.600 2421.560 2050.225 ;
        RECT 2424.135 2049.600 2424.305 2050.225 ;
        RECT 2425.125 2049.600 2425.295 2050.230 ;
        RECT 2426.840 2049.600 2436.655 2050.875 ;
        RECT 2437.715 2049.600 2437.885 2050.225 ;
        RECT 2440.460 2049.600 2440.630 2050.225 ;
        RECT 2441.450 2049.600 2441.620 2050.230 ;
        RECT 2343.000 2048.000 2442.425 2049.600 ;
        RECT 2695.520 2036.835 2734.160 2037.005 ;
        RECT 2695.605 2036.085 2696.815 2036.835 ;
        RECT 2697.455 2036.355 2697.730 2036.835 ;
        RECT 2698.315 2036.435 2698.650 2036.835 ;
        RECT 2699.265 2036.455 2699.595 2036.835 ;
        RECT 2700.645 2036.455 2700.975 2036.835 ;
        RECT 2701.585 2036.290 2706.930 2036.835 ;
        RECT 2695.605 2035.545 2696.125 2036.085 ;
        RECT 2703.170 2035.460 2703.510 2036.290 ;
        RECT 2707.105 2036.085 2708.315 2036.835 ;
        RECT 2708.485 2036.110 2708.775 2036.835 ;
        RECT 2709.420 2036.455 2709.750 2036.835 ;
        RECT 2707.105 2035.545 2707.625 2036.085 ;
        RECT 2710.350 2035.995 2710.610 2036.835 ;
        RECT 2710.785 2036.290 2716.130 2036.835 ;
        RECT 2712.370 2035.460 2712.710 2036.290 ;
        RECT 2716.305 2036.065 2719.815 2036.835 ;
        RECT 2719.985 2036.085 2721.195 2036.835 ;
        RECT 2721.365 2036.110 2721.655 2036.835 ;
        RECT 2721.830 2036.435 2722.165 2036.835 ;
        RECT 2722.750 2036.355 2723.025 2036.835 ;
        RECT 2723.665 2036.290 2729.010 2036.835 ;
        RECT 2716.305 2035.545 2717.955 2036.065 ;
        RECT 2719.985 2035.545 2720.505 2036.085 ;
        RECT 2725.250 2035.460 2725.590 2036.290 ;
        RECT 2729.185 2036.065 2730.855 2036.835 ;
        RECT 2731.925 2036.455 2732.255 2036.835 ;
        RECT 2732.865 2036.085 2734.075 2036.835 ;
        RECT 2729.185 2035.545 2729.935 2036.065 ;
        RECT 2733.555 2035.545 2734.075 2036.085 ;
        RECT 2695.605 2032.315 2696.125 2032.855 ;
        RECT 2695.605 2031.565 2696.815 2032.315 ;
        RECT 2699.950 2032.110 2700.290 2032.940 ;
        RECT 2703.885 2032.335 2705.535 2032.855 ;
        RECT 2697.425 2031.565 2697.755 2031.945 ;
        RECT 2698.365 2031.565 2703.710 2032.110 ;
        RECT 2703.885 2031.565 2707.395 2032.335 ;
        RECT 2708.485 2031.565 2708.775 2032.290 ;
        RECT 2710.530 2032.110 2710.870 2032.940 ;
        RECT 2716.050 2032.110 2716.390 2032.940 ;
        RECT 2721.570 2032.110 2721.910 2032.940 ;
        RECT 2727.090 2032.110 2727.430 2032.940 ;
        RECT 2731.025 2032.335 2731.775 2032.855 ;
        RECT 2708.945 2031.565 2714.290 2032.110 ;
        RECT 2714.465 2031.565 2719.810 2032.110 ;
        RECT 2719.985 2031.565 2725.330 2032.110 ;
        RECT 2725.505 2031.565 2730.850 2032.110 ;
        RECT 2731.025 2031.565 2732.695 2032.335 ;
        RECT 2733.555 2032.315 2734.075 2032.855 ;
        RECT 2732.865 2031.565 2734.075 2032.315 ;
        RECT 2695.520 2031.395 2734.160 2031.565 ;
        RECT 2695.605 2030.645 2696.815 2031.395 ;
        RECT 2696.985 2030.850 2702.330 2031.395 ;
        RECT 2702.505 2030.850 2707.850 2031.395 ;
        RECT 2708.025 2030.850 2713.370 2031.395 ;
        RECT 2713.545 2030.850 2718.890 2031.395 ;
        RECT 2695.605 2030.105 2696.125 2030.645 ;
        RECT 2698.570 2030.020 2698.910 2030.850 ;
        RECT 2704.090 2030.020 2704.430 2030.850 ;
        RECT 2709.610 2030.020 2709.950 2030.850 ;
        RECT 2715.130 2030.020 2715.470 2030.850 ;
        RECT 2719.065 2030.625 2720.735 2031.395 ;
        RECT 2721.365 2030.670 2721.655 2031.395 ;
        RECT 2721.825 2030.850 2727.170 2031.395 ;
        RECT 2727.345 2030.850 2732.690 2031.395 ;
        RECT 2719.065 2030.105 2719.815 2030.625 ;
        RECT 2723.410 2030.020 2723.750 2030.850 ;
        RECT 2728.930 2030.020 2729.270 2030.850 ;
        RECT 2732.865 2030.645 2734.075 2031.395 ;
        RECT 2733.555 2030.105 2734.075 2030.645 ;
        RECT 2695.605 2026.875 2696.125 2027.415 ;
        RECT 2695.605 2026.125 2696.815 2026.875 ;
        RECT 2698.570 2026.670 2698.910 2027.500 ;
        RECT 2704.090 2026.670 2704.430 2027.500 ;
        RECT 2696.985 2026.125 2702.330 2026.670 ;
        RECT 2702.505 2026.125 2707.850 2026.670 ;
        RECT 2708.485 2026.125 2708.775 2026.850 ;
        RECT 2710.530 2026.670 2710.870 2027.500 ;
        RECT 2716.050 2026.670 2716.390 2027.500 ;
        RECT 2721.570 2026.670 2721.910 2027.500 ;
        RECT 2727.090 2026.670 2727.430 2027.500 ;
        RECT 2731.025 2026.895 2731.775 2027.415 ;
        RECT 2708.945 2026.125 2714.290 2026.670 ;
        RECT 2714.465 2026.125 2719.810 2026.670 ;
        RECT 2719.985 2026.125 2725.330 2026.670 ;
        RECT 2725.505 2026.125 2730.850 2026.670 ;
        RECT 2731.025 2026.125 2732.695 2026.895 ;
        RECT 2733.555 2026.875 2734.075 2027.415 ;
        RECT 2732.865 2026.125 2734.075 2026.875 ;
        RECT 2695.520 2025.955 2734.160 2026.125 ;
        RECT 2695.605 2025.205 2696.815 2025.955 ;
        RECT 2697.425 2025.575 2697.755 2025.955 ;
        RECT 2698.365 2025.410 2703.710 2025.955 ;
        RECT 2703.885 2025.410 2709.230 2025.955 ;
        RECT 2709.405 2025.410 2714.750 2025.955 ;
        RECT 2714.925 2025.410 2720.270 2025.955 ;
        RECT 2695.605 2024.665 2696.125 2025.205 ;
        RECT 2699.950 2024.580 2700.290 2025.410 ;
        RECT 2705.470 2024.580 2705.810 2025.410 ;
        RECT 2710.990 2024.580 2711.330 2025.410 ;
        RECT 2716.510 2024.580 2716.850 2025.410 ;
        RECT 2721.365 2025.230 2721.655 2025.955 ;
        RECT 2721.825 2025.410 2727.170 2025.955 ;
        RECT 2727.345 2025.410 2732.690 2025.955 ;
        RECT 2723.410 2024.580 2723.750 2025.410 ;
        RECT 2728.930 2024.580 2729.270 2025.410 ;
        RECT 2732.865 2025.205 2734.075 2025.955 ;
        RECT 2733.555 2024.665 2734.075 2025.205 ;
        RECT 2695.605 2021.435 2696.125 2021.975 ;
        RECT 2695.605 2020.685 2696.815 2021.435 ;
        RECT 2698.570 2021.230 2698.910 2022.060 ;
        RECT 2704.090 2021.230 2704.430 2022.060 ;
        RECT 2696.985 2020.685 2702.330 2021.230 ;
        RECT 2702.505 2020.685 2707.850 2021.230 ;
        RECT 2708.485 2020.685 2708.775 2021.410 ;
        RECT 2710.530 2021.230 2710.870 2022.060 ;
        RECT 2716.050 2021.230 2716.390 2022.060 ;
        RECT 2721.570 2021.230 2721.910 2022.060 ;
        RECT 2727.090 2021.230 2727.430 2022.060 ;
        RECT 2731.025 2021.455 2731.775 2021.975 ;
        RECT 2708.945 2020.685 2714.290 2021.230 ;
        RECT 2714.465 2020.685 2719.810 2021.230 ;
        RECT 2719.985 2020.685 2725.330 2021.230 ;
        RECT 2725.505 2020.685 2730.850 2021.230 ;
        RECT 2731.025 2020.685 2732.695 2021.455 ;
        RECT 2733.555 2021.435 2734.075 2021.975 ;
        RECT 2732.865 2020.685 2734.075 2021.435 ;
        RECT 2695.520 2020.515 2734.160 2020.685 ;
        RECT 2695.605 2019.765 2696.815 2020.515 ;
        RECT 2697.415 2020.135 2697.745 2020.515 ;
        RECT 2699.700 2019.795 2699.990 2020.515 ;
        RECT 2702.050 2020.055 2702.220 2020.515 ;
        RECT 2702.910 2020.135 2703.240 2020.515 ;
        RECT 2705.795 2020.055 2705.965 2020.515 ;
        RECT 2706.645 2019.970 2711.990 2020.515 ;
        RECT 2712.165 2019.970 2717.510 2020.515 ;
        RECT 2695.605 2019.225 2696.125 2019.765 ;
        RECT 2708.230 2019.140 2708.570 2019.970 ;
        RECT 2713.750 2019.140 2714.090 2019.970 ;
        RECT 2717.685 2019.745 2721.195 2020.515 ;
        RECT 2721.365 2019.790 2721.655 2020.515 ;
        RECT 2721.825 2019.970 2727.170 2020.515 ;
        RECT 2727.345 2019.970 2732.690 2020.515 ;
        RECT 2717.685 2019.225 2719.335 2019.745 ;
        RECT 2723.410 2019.140 2723.750 2019.970 ;
        RECT 2728.930 2019.140 2729.270 2019.970 ;
        RECT 2732.865 2019.765 2734.075 2020.515 ;
        RECT 2733.555 2019.225 2734.075 2019.765 ;
        RECT 2695.605 2015.995 2696.125 2016.535 ;
        RECT 2695.605 2015.245 2696.815 2015.995 ;
        RECT 2699.950 2015.790 2700.290 2016.620 ;
        RECT 2703.885 2016.015 2705.535 2016.535 ;
        RECT 2697.425 2015.245 2697.755 2015.625 ;
        RECT 2698.365 2015.245 2703.710 2015.790 ;
        RECT 2703.885 2015.245 2707.395 2016.015 ;
        RECT 2708.485 2015.245 2708.775 2015.970 ;
        RECT 2710.530 2015.790 2710.870 2016.620 ;
        RECT 2716.050 2015.790 2716.390 2016.620 ;
        RECT 2721.570 2015.790 2721.910 2016.620 ;
        RECT 2727.090 2015.790 2727.430 2016.620 ;
        RECT 2731.025 2016.015 2731.775 2016.535 ;
        RECT 2708.945 2015.245 2714.290 2015.790 ;
        RECT 2714.465 2015.245 2719.810 2015.790 ;
        RECT 2719.985 2015.245 2725.330 2015.790 ;
        RECT 2725.505 2015.245 2730.850 2015.790 ;
        RECT 2731.025 2015.245 2732.695 2016.015 ;
        RECT 2733.555 2015.995 2734.075 2016.535 ;
        RECT 2732.865 2015.245 2734.075 2015.995 ;
        RECT 2695.520 2015.075 2734.160 2015.245 ;
        RECT 2695.605 2014.325 2696.815 2015.075 ;
        RECT 2697.415 2014.695 2697.745 2015.075 ;
        RECT 2699.700 2014.355 2699.990 2015.075 ;
        RECT 2702.050 2014.615 2702.220 2015.075 ;
        RECT 2702.910 2014.695 2703.240 2015.075 ;
        RECT 2705.795 2014.615 2705.965 2015.075 ;
        RECT 2706.645 2014.530 2711.990 2015.075 ;
        RECT 2712.165 2014.530 2717.510 2015.075 ;
        RECT 2695.605 2013.785 2696.125 2014.325 ;
        RECT 2708.230 2013.700 2708.570 2014.530 ;
        RECT 2713.750 2013.700 2714.090 2014.530 ;
        RECT 2717.685 2014.305 2721.195 2015.075 ;
        RECT 2721.365 2014.350 2721.655 2015.075 ;
        RECT 2721.825 2014.530 2727.170 2015.075 ;
        RECT 2727.345 2014.530 2732.690 2015.075 ;
        RECT 2717.685 2013.785 2719.335 2014.305 ;
        RECT 2723.410 2013.700 2723.750 2014.530 ;
        RECT 2728.930 2013.700 2729.270 2014.530 ;
        RECT 2732.865 2014.325 2734.075 2015.075 ;
        RECT 2733.555 2013.785 2734.075 2014.325 ;
        RECT 2695.605 2010.555 2696.125 2011.095 ;
        RECT 2698.365 2010.575 2699.575 2011.095 ;
        RECT 2705.725 2010.575 2706.935 2011.095 ;
        RECT 2695.605 2009.805 2696.815 2010.555 ;
        RECT 2697.425 2009.805 2697.755 2010.185 ;
        RECT 2698.365 2009.805 2700.955 2010.575 ;
        RECT 2702.015 2009.805 2702.345 2010.205 ;
        RECT 2704.305 2009.805 2704.815 2010.340 ;
        RECT 2705.725 2009.805 2708.315 2010.575 ;
        RECT 2708.485 2009.805 2708.775 2010.530 ;
        RECT 2710.530 2010.350 2710.870 2011.180 ;
        RECT 2716.050 2010.350 2716.390 2011.180 ;
        RECT 2721.570 2010.350 2721.910 2011.180 ;
        RECT 2727.090 2010.350 2727.430 2011.180 ;
        RECT 2731.025 2010.575 2731.775 2011.095 ;
        RECT 2708.945 2009.805 2714.290 2010.350 ;
        RECT 2714.465 2009.805 2719.810 2010.350 ;
        RECT 2719.985 2009.805 2725.330 2010.350 ;
        RECT 2725.505 2009.805 2730.850 2010.350 ;
        RECT 2731.025 2009.805 2732.695 2010.575 ;
        RECT 2733.555 2010.555 2734.075 2011.095 ;
        RECT 2732.865 2009.805 2734.075 2010.555 ;
        RECT 2695.520 2009.635 2734.160 2009.805 ;
        RECT 2695.605 2008.885 2696.815 2009.635 ;
        RECT 2696.985 2009.090 2702.330 2009.635 ;
        RECT 2702.505 2009.090 2707.850 2009.635 ;
        RECT 2708.025 2009.090 2713.370 2009.635 ;
        RECT 2713.545 2009.090 2718.890 2009.635 ;
        RECT 2695.605 2008.345 2696.125 2008.885 ;
        RECT 2698.570 2008.260 2698.910 2009.090 ;
        RECT 2704.090 2008.260 2704.430 2009.090 ;
        RECT 2709.610 2008.260 2709.950 2009.090 ;
        RECT 2715.130 2008.260 2715.470 2009.090 ;
        RECT 2719.065 2008.865 2720.735 2009.635 ;
        RECT 2721.365 2008.910 2721.655 2009.635 ;
        RECT 2721.825 2009.090 2727.170 2009.635 ;
        RECT 2727.345 2009.090 2732.690 2009.635 ;
        RECT 2719.065 2008.345 2719.815 2008.865 ;
        RECT 2723.410 2008.260 2723.750 2009.090 ;
        RECT 2728.930 2008.260 2729.270 2009.090 ;
        RECT 2732.865 2008.885 2734.075 2009.635 ;
        RECT 2733.555 2008.345 2734.075 2008.885 ;
        RECT 2695.605 2005.115 2696.125 2005.655 ;
        RECT 2695.605 2004.365 2696.815 2005.115 ;
        RECT 2699.950 2004.910 2700.290 2005.740 ;
        RECT 2703.885 2005.135 2705.535 2005.655 ;
        RECT 2697.425 2004.365 2697.755 2004.745 ;
        RECT 2698.365 2004.365 2703.710 2004.910 ;
        RECT 2703.885 2004.365 2707.395 2005.135 ;
        RECT 2708.485 2004.365 2708.775 2005.090 ;
        RECT 2710.530 2004.910 2710.870 2005.740 ;
        RECT 2716.050 2004.910 2716.390 2005.740 ;
        RECT 2721.570 2004.910 2721.910 2005.740 ;
        RECT 2727.090 2004.910 2727.430 2005.740 ;
        RECT 2731.025 2005.135 2731.775 2005.655 ;
        RECT 2708.945 2004.365 2714.290 2004.910 ;
        RECT 2714.465 2004.365 2719.810 2004.910 ;
        RECT 2719.985 2004.365 2725.330 2004.910 ;
        RECT 2725.505 2004.365 2730.850 2004.910 ;
        RECT 2731.025 2004.365 2732.695 2005.135 ;
        RECT 2733.555 2005.115 2734.075 2005.655 ;
        RECT 2732.865 2004.365 2734.075 2005.115 ;
        RECT 2695.520 2004.195 2734.160 2004.365 ;
        RECT 2695.605 2003.445 2696.815 2004.195 ;
        RECT 2696.985 2003.650 2702.330 2004.195 ;
        RECT 2702.505 2003.650 2707.850 2004.195 ;
        RECT 2708.025 2003.650 2713.370 2004.195 ;
        RECT 2713.545 2003.650 2718.890 2004.195 ;
        RECT 2695.605 2002.905 2696.125 2003.445 ;
        RECT 2698.570 2002.820 2698.910 2003.650 ;
        RECT 2704.090 2002.820 2704.430 2003.650 ;
        RECT 2709.610 2002.820 2709.950 2003.650 ;
        RECT 2715.130 2002.820 2715.470 2003.650 ;
        RECT 2719.065 2003.425 2720.735 2004.195 ;
        RECT 2721.365 2003.470 2721.655 2004.195 ;
        RECT 2721.825 2003.650 2727.170 2004.195 ;
        RECT 2727.345 2003.650 2732.690 2004.195 ;
        RECT 2719.065 2002.905 2719.815 2003.425 ;
        RECT 2723.410 2002.820 2723.750 2003.650 ;
        RECT 2728.930 2002.820 2729.270 2003.650 ;
        RECT 2732.865 2003.445 2734.075 2004.195 ;
        RECT 2733.555 2002.905 2734.075 2003.445 ;
        RECT 2695.605 1999.675 2696.125 2000.215 ;
        RECT 2696.985 1999.695 2698.635 2000.215 ;
        RECT 2695.605 1998.925 2696.815 1999.675 ;
        RECT 2696.985 1998.925 2700.495 1999.695 ;
        RECT 2701.605 1998.925 2701.845 1999.735 ;
        RECT 2702.515 1998.925 2702.785 1999.735 ;
        RECT 2704.550 1999.470 2704.890 2000.300 ;
        RECT 2702.965 1998.925 2708.310 1999.470 ;
        RECT 2708.485 1998.925 2708.775 1999.650 ;
        RECT 2710.530 1999.470 2710.870 2000.300 ;
        RECT 2716.050 1999.470 2716.390 2000.300 ;
        RECT 2721.570 1999.470 2721.910 2000.300 ;
        RECT 2727.090 1999.470 2727.430 2000.300 ;
        RECT 2731.025 1999.695 2731.775 2000.215 ;
        RECT 2708.945 1998.925 2714.290 1999.470 ;
        RECT 2714.465 1998.925 2719.810 1999.470 ;
        RECT 2719.985 1998.925 2725.330 1999.470 ;
        RECT 2725.505 1998.925 2730.850 1999.470 ;
        RECT 2731.025 1998.925 2732.695 1999.695 ;
        RECT 2733.555 1999.675 2734.075 2000.215 ;
        RECT 2732.865 1998.925 2734.075 1999.675 ;
        RECT 2695.520 1998.755 2734.160 1998.925 ;
        RECT 2695.605 1998.005 2696.815 1998.755 ;
        RECT 2697.425 1998.375 2697.755 1998.755 ;
        RECT 2695.605 1997.465 2696.125 1998.005 ;
        RECT 2698.365 1997.985 2701.875 1998.755 ;
        RECT 2702.055 1998.015 2702.385 1998.755 ;
        RECT 2703.090 1998.395 2703.420 1998.755 ;
        RECT 2698.365 1997.465 2700.015 1997.985 ;
        RECT 2704.785 1997.975 2705.080 1998.755 ;
        RECT 2705.265 1998.210 2710.610 1998.755 ;
        RECT 2710.785 1998.210 2716.130 1998.755 ;
        RECT 2706.850 1997.380 2707.190 1998.210 ;
        RECT 2712.370 1997.380 2712.710 1998.210 ;
        RECT 2716.305 1997.985 2719.815 1998.755 ;
        RECT 2719.985 1998.005 2721.195 1998.755 ;
        RECT 2721.365 1998.030 2721.655 1998.755 ;
        RECT 2721.825 1998.210 2727.170 1998.755 ;
        RECT 2727.345 1998.210 2732.690 1998.755 ;
        RECT 2716.305 1997.465 2717.955 1997.985 ;
        RECT 2719.985 1997.465 2720.505 1998.005 ;
        RECT 2723.410 1997.380 2723.750 1998.210 ;
        RECT 2728.930 1997.380 2729.270 1998.210 ;
        RECT 2732.865 1998.005 2734.075 1998.755 ;
        RECT 2733.555 1997.465 2734.075 1998.005 ;
        RECT 2695.605 1994.235 2696.125 1994.775 ;
        RECT 2695.605 1993.485 2696.815 1994.235 ;
        RECT 2698.570 1994.030 2698.910 1994.860 ;
        RECT 2704.090 1994.030 2704.430 1994.860 ;
        RECT 2696.985 1993.485 2702.330 1994.030 ;
        RECT 2702.505 1993.485 2707.850 1994.030 ;
        RECT 2708.485 1993.485 2708.775 1994.210 ;
        RECT 2710.530 1994.030 2710.870 1994.860 ;
        RECT 2716.050 1994.030 2716.390 1994.860 ;
        RECT 2721.570 1994.030 2721.910 1994.860 ;
        RECT 2708.945 1993.485 2714.290 1994.030 ;
        RECT 2714.465 1993.485 2719.810 1994.030 ;
        RECT 2719.985 1993.485 2725.330 1994.030 ;
        RECT 2725.515 1993.485 2725.845 1993.965 ;
        RECT 2726.355 1993.485 2726.685 1993.965 ;
        RECT 2727.195 1993.485 2727.525 1993.965 ;
        RECT 2728.035 1993.485 2728.365 1993.965 ;
        RECT 2728.875 1993.485 2729.205 1993.965 ;
        RECT 2729.715 1993.485 2730.045 1993.965 ;
        RECT 2730.555 1993.485 2730.885 1993.965 ;
        RECT 2731.395 1993.485 2731.725 1993.965 ;
        RECT 2732.235 1993.485 2732.565 1994.285 ;
        RECT 2733.555 1994.235 2734.075 1994.775 ;
        RECT 2732.865 1993.485 2734.075 1994.235 ;
        RECT 2695.520 1993.315 2734.160 1993.485 ;
        RECT 2695.605 1992.565 2696.815 1993.315 ;
        RECT 2697.425 1992.935 2697.755 1993.315 ;
        RECT 2698.365 1992.770 2703.710 1993.315 ;
        RECT 2703.885 1992.770 2709.230 1993.315 ;
        RECT 2709.405 1992.770 2714.750 1993.315 ;
        RECT 2714.925 1992.770 2720.270 1993.315 ;
        RECT 2695.605 1992.025 2696.125 1992.565 ;
        RECT 2699.950 1991.940 2700.290 1992.770 ;
        RECT 2705.470 1991.940 2705.810 1992.770 ;
        RECT 2710.990 1991.940 2711.330 1992.770 ;
        RECT 2716.510 1991.940 2716.850 1992.770 ;
        RECT 2721.365 1992.590 2721.655 1993.315 ;
        RECT 2721.825 1992.770 2727.170 1993.315 ;
        RECT 2727.345 1992.770 2732.690 1993.315 ;
        RECT 2723.410 1991.940 2723.750 1992.770 ;
        RECT 2728.930 1991.940 2729.270 1992.770 ;
        RECT 2732.865 1992.565 2734.075 1993.315 ;
        RECT 2733.555 1992.025 2734.075 1992.565 ;
        RECT 2695.605 1988.795 2696.125 1989.335 ;
        RECT 2695.605 1988.045 2696.815 1988.795 ;
        RECT 2698.570 1988.590 2698.910 1989.420 ;
        RECT 2704.090 1988.590 2704.430 1989.420 ;
        RECT 2696.985 1988.045 2702.330 1988.590 ;
        RECT 2702.505 1988.045 2707.850 1988.590 ;
        RECT 2708.485 1988.045 2708.775 1988.770 ;
        RECT 2710.530 1988.590 2710.870 1989.420 ;
        RECT 2716.050 1988.590 2716.390 1989.420 ;
        RECT 2721.570 1988.590 2721.910 1989.420 ;
        RECT 2727.090 1988.590 2727.430 1989.420 ;
        RECT 2731.025 1988.815 2731.775 1989.335 ;
        RECT 2708.945 1988.045 2714.290 1988.590 ;
        RECT 2714.465 1988.045 2719.810 1988.590 ;
        RECT 2719.985 1988.045 2725.330 1988.590 ;
        RECT 2725.505 1988.045 2730.850 1988.590 ;
        RECT 2731.025 1988.045 2732.695 1988.815 ;
        RECT 2733.555 1988.795 2734.075 1989.335 ;
        RECT 2732.865 1988.045 2734.075 1988.795 ;
        RECT 2695.520 1987.875 2734.160 1988.045 ;
        RECT 2695.605 1987.125 2696.815 1987.875 ;
        RECT 2697.715 1987.135 2698.045 1987.875 ;
        RECT 2698.555 1987.475 2698.885 1987.875 ;
        RECT 2699.745 1987.330 2705.090 1987.875 ;
        RECT 2705.265 1987.330 2710.610 1987.875 ;
        RECT 2710.785 1987.330 2716.130 1987.875 ;
        RECT 2695.605 1986.585 2696.125 1987.125 ;
        RECT 2701.330 1986.500 2701.670 1987.330 ;
        RECT 2706.850 1986.500 2707.190 1987.330 ;
        RECT 2712.370 1986.500 2712.710 1987.330 ;
        RECT 2716.305 1987.105 2719.815 1987.875 ;
        RECT 2719.985 1987.125 2721.195 1987.875 ;
        RECT 2721.365 1987.150 2721.655 1987.875 ;
        RECT 2721.825 1987.330 2727.170 1987.875 ;
        RECT 2727.345 1987.330 2732.690 1987.875 ;
        RECT 2716.305 1986.585 2717.955 1987.105 ;
        RECT 2719.985 1986.585 2720.505 1987.125 ;
        RECT 2723.410 1986.500 2723.750 1987.330 ;
        RECT 2728.930 1986.500 2729.270 1987.330 ;
        RECT 2732.865 1987.125 2734.075 1987.875 ;
        RECT 2733.555 1986.585 2734.075 1987.125 ;
        RECT 2695.605 1983.355 2696.125 1983.895 ;
        RECT 2695.605 1982.605 2696.815 1983.355 ;
        RECT 2699.950 1983.150 2700.290 1983.980 ;
        RECT 2703.885 1983.375 2705.535 1983.895 ;
        RECT 2697.425 1982.605 2697.755 1982.985 ;
        RECT 2698.365 1982.605 2703.710 1983.150 ;
        RECT 2703.885 1982.605 2707.395 1983.375 ;
        RECT 2708.485 1982.605 2708.775 1983.330 ;
        RECT 2710.530 1983.150 2710.870 1983.980 ;
        RECT 2716.050 1983.150 2716.390 1983.980 ;
        RECT 2721.570 1983.150 2721.910 1983.980 ;
        RECT 2727.090 1983.150 2727.430 1983.980 ;
        RECT 2731.025 1983.375 2731.775 1983.895 ;
        RECT 2708.945 1982.605 2714.290 1983.150 ;
        RECT 2714.465 1982.605 2719.810 1983.150 ;
        RECT 2719.985 1982.605 2725.330 1983.150 ;
        RECT 2725.505 1982.605 2730.850 1983.150 ;
        RECT 2731.025 1982.605 2732.695 1983.375 ;
        RECT 2733.555 1983.355 2734.075 1983.895 ;
        RECT 2732.865 1982.605 2734.075 1983.355 ;
        RECT 2523.330 1981.785 2523.670 1982.445 ;
        RECT 2695.520 1982.435 2734.160 1982.605 ;
        RECT 2522.130 1981.615 2523.935 1981.785 ;
        RECT 2695.605 1981.685 2696.815 1982.435 ;
        RECT 2697.725 1981.900 2698.235 1982.435 ;
        RECT 2700.195 1982.035 2700.525 1982.435 ;
        RECT 2701.210 1981.760 2701.450 1982.435 ;
        RECT 2702.840 1981.985 2703.170 1982.435 ;
        RECT 2704.090 1981.995 2704.405 1982.435 ;
        RECT 2704.805 1981.890 2710.150 1982.435 ;
        RECT 2710.325 1981.890 2715.670 1982.435 ;
        RECT 2715.845 1981.890 2721.190 1982.435 ;
        RECT 2695.605 1981.145 2696.125 1981.685 ;
        RECT 2706.390 1981.060 2706.730 1981.890 ;
        RECT 2711.910 1981.060 2712.250 1981.890 ;
        RECT 2717.430 1981.060 2717.770 1981.890 ;
        RECT 2721.365 1981.710 2721.655 1982.435 ;
        RECT 2721.825 1981.890 2727.170 1982.435 ;
        RECT 2727.345 1981.890 2732.690 1982.435 ;
        RECT 2723.410 1981.060 2723.750 1981.890 ;
        RECT 2728.930 1981.060 2729.270 1981.890 ;
        RECT 2732.865 1981.685 2734.075 1982.435 ;
        RECT 2733.555 1981.145 2734.075 1981.685 ;
        RECT 2695.605 1977.915 2696.125 1978.455 ;
        RECT 2695.605 1977.165 2696.815 1977.915 ;
        RECT 2696.985 1977.165 2697.245 1977.985 ;
        RECT 2701.790 1977.710 2702.130 1978.540 ;
        RECT 2705.725 1977.935 2706.935 1978.455 ;
        RECT 2699.275 1977.165 2699.605 1977.625 ;
        RECT 2700.205 1977.165 2705.550 1977.710 ;
        RECT 2705.725 1977.165 2708.315 1977.935 ;
        RECT 2708.485 1977.165 2708.775 1977.890 ;
        RECT 2710.530 1977.710 2710.870 1978.540 ;
        RECT 2716.050 1977.710 2716.390 1978.540 ;
        RECT 2721.570 1977.710 2721.910 1978.540 ;
        RECT 2727.090 1977.710 2727.430 1978.540 ;
        RECT 2731.025 1977.935 2731.775 1978.455 ;
        RECT 2708.945 1977.165 2714.290 1977.710 ;
        RECT 2714.465 1977.165 2719.810 1977.710 ;
        RECT 2719.985 1977.165 2725.330 1977.710 ;
        RECT 2725.505 1977.165 2730.850 1977.710 ;
        RECT 2731.025 1977.165 2732.695 1977.935 ;
        RECT 2733.555 1977.915 2734.075 1978.455 ;
        RECT 2732.865 1977.165 2734.075 1977.915 ;
        RECT 2695.520 1976.995 2734.160 1977.165 ;
        RECT 2695.605 1976.245 2696.815 1976.995 ;
        RECT 2697.425 1976.615 2697.755 1976.995 ;
        RECT 2698.365 1976.450 2703.710 1976.995 ;
        RECT 2703.885 1976.450 2709.230 1976.995 ;
        RECT 2709.405 1976.450 2714.750 1976.995 ;
        RECT 2714.925 1976.450 2720.270 1976.995 ;
        RECT 2695.605 1975.705 2696.125 1976.245 ;
        RECT 2699.950 1975.620 2700.290 1976.450 ;
        RECT 2705.470 1975.620 2705.810 1976.450 ;
        RECT 2710.990 1975.620 2711.330 1976.450 ;
        RECT 2716.510 1975.620 2716.850 1976.450 ;
        RECT 2721.365 1976.270 2721.655 1976.995 ;
        RECT 2721.825 1976.450 2727.170 1976.995 ;
        RECT 2727.345 1976.450 2732.690 1976.995 ;
        RECT 2723.410 1975.620 2723.750 1976.450 ;
        RECT 2728.930 1975.620 2729.270 1976.450 ;
        RECT 2732.865 1976.245 2734.075 1976.995 ;
        RECT 2733.555 1975.705 2734.075 1976.245 ;
        RECT 2523.330 1974.255 2523.670 1974.915 ;
        RECT 2522.130 1974.085 2523.935 1974.255 ;
        RECT 2695.605 1972.475 2696.125 1973.015 ;
        RECT 2696.985 1972.475 2697.505 1973.015 ;
        RECT 2695.605 1971.725 2696.815 1972.475 ;
        RECT 2696.985 1971.725 2698.195 1972.475 ;
        RECT 2698.365 1971.725 2698.705 1972.450 ;
        RECT 2703.630 1972.270 2703.970 1973.100 ;
        RECT 2701.035 1971.725 2701.365 1972.205 ;
        RECT 2702.045 1971.725 2707.390 1972.270 ;
        RECT 2708.485 1971.725 2708.775 1972.450 ;
        RECT 2710.530 1972.270 2710.870 1973.100 ;
        RECT 2716.050 1972.270 2716.390 1973.100 ;
        RECT 2721.570 1972.270 2721.910 1973.100 ;
        RECT 2727.090 1972.270 2727.430 1973.100 ;
        RECT 2731.025 1972.495 2731.775 1973.015 ;
        RECT 2708.945 1971.725 2714.290 1972.270 ;
        RECT 2714.465 1971.725 2719.810 1972.270 ;
        RECT 2719.985 1971.725 2725.330 1972.270 ;
        RECT 2725.505 1971.725 2730.850 1972.270 ;
        RECT 2731.025 1971.725 2732.695 1972.495 ;
        RECT 2733.555 1972.475 2734.075 1973.015 ;
        RECT 2732.865 1971.725 2734.075 1972.475 ;
        RECT 2695.520 1971.555 2734.160 1971.725 ;
        RECT 2695.605 1970.805 2696.815 1971.555 ;
        RECT 2695.605 1970.265 2696.125 1970.805 ;
        RECT 2697.905 1970.735 2698.165 1971.555 ;
        RECT 2699.275 1971.155 2699.605 1971.555 ;
        RECT 2700.115 1971.155 2700.490 1971.555 ;
        RECT 2702.760 1971.155 2703.090 1971.555 ;
        RECT 2703.885 1971.010 2709.230 1971.555 ;
        RECT 2709.405 1971.010 2714.750 1971.555 ;
        RECT 2714.925 1971.010 2720.270 1971.555 ;
        RECT 2705.470 1970.180 2705.810 1971.010 ;
        RECT 2710.990 1970.180 2711.330 1971.010 ;
        RECT 2716.510 1970.180 2716.850 1971.010 ;
        RECT 2721.365 1970.830 2721.655 1971.555 ;
        RECT 2721.825 1971.010 2727.170 1971.555 ;
        RECT 2727.345 1971.010 2732.690 1971.555 ;
        RECT 2723.410 1970.180 2723.750 1971.010 ;
        RECT 2728.930 1970.180 2729.270 1971.010 ;
        RECT 2732.865 1970.805 2734.075 1971.555 ;
        RECT 2733.555 1970.265 2734.075 1970.805 ;
        RECT 2523.330 1968.275 2523.670 1968.935 ;
        RECT 2522.130 1968.105 2523.935 1968.275 ;
        RECT 2695.605 1967.035 2696.125 1967.575 ;
        RECT 2695.605 1966.285 2696.815 1967.035 ;
        RECT 2697.425 1966.285 2697.755 1966.665 ;
        RECT 2699.725 1966.285 2700.035 1967.085 ;
        RECT 2701.790 1966.830 2702.130 1967.660 ;
        RECT 2705.725 1967.055 2706.935 1967.575 ;
        RECT 2700.205 1966.285 2705.550 1966.830 ;
        RECT 2705.725 1966.285 2708.315 1967.055 ;
        RECT 2708.485 1966.285 2708.775 1967.010 ;
        RECT 2710.530 1966.830 2710.870 1967.660 ;
        RECT 2716.050 1966.830 2716.390 1967.660 ;
        RECT 2721.570 1966.830 2721.910 1967.660 ;
        RECT 2727.090 1966.830 2727.430 1967.660 ;
        RECT 2731.025 1967.055 2731.775 1967.575 ;
        RECT 2708.945 1966.285 2714.290 1966.830 ;
        RECT 2714.465 1966.285 2719.810 1966.830 ;
        RECT 2719.985 1966.285 2725.330 1966.830 ;
        RECT 2725.505 1966.285 2730.850 1966.830 ;
        RECT 2731.025 1966.285 2732.695 1967.055 ;
        RECT 2733.555 1967.035 2734.075 1967.575 ;
        RECT 2732.865 1966.285 2734.075 1967.035 ;
        RECT 2695.520 1966.115 2734.160 1966.285 ;
        RECT 2695.605 1965.365 2696.815 1966.115 ;
        RECT 2697.725 1965.580 2698.235 1966.115 ;
        RECT 2700.195 1965.715 2700.525 1966.115 ;
        RECT 2701.125 1965.570 2706.470 1966.115 ;
        RECT 2706.645 1965.570 2711.990 1966.115 ;
        RECT 2712.165 1965.570 2717.510 1966.115 ;
        RECT 2695.605 1964.825 2696.125 1965.365 ;
        RECT 2702.710 1964.740 2703.050 1965.570 ;
        RECT 2708.230 1964.740 2708.570 1965.570 ;
        RECT 2713.750 1964.740 2714.090 1965.570 ;
        RECT 2717.685 1965.345 2721.195 1966.115 ;
        RECT 2721.365 1965.390 2721.655 1966.115 ;
        RECT 2721.825 1965.570 2727.170 1966.115 ;
        RECT 2727.345 1965.570 2732.690 1966.115 ;
        RECT 2717.685 1964.825 2719.335 1965.345 ;
        RECT 2723.410 1964.740 2723.750 1965.570 ;
        RECT 2728.930 1964.740 2729.270 1965.570 ;
        RECT 2732.865 1965.365 2734.075 1966.115 ;
        RECT 2733.555 1964.825 2734.075 1965.365 ;
        RECT 2523.330 1962.330 2523.670 1962.990 ;
        RECT 2522.130 1962.160 2523.935 1962.330 ;
        RECT 2695.605 1961.595 2696.125 1962.135 ;
        RECT 2695.605 1960.845 2696.815 1961.595 ;
        RECT 2699.950 1961.390 2700.290 1962.220 ;
        RECT 2703.885 1961.615 2705.535 1962.135 ;
        RECT 2697.425 1960.845 2697.755 1961.225 ;
        RECT 2698.365 1960.845 2703.710 1961.390 ;
        RECT 2703.885 1960.845 2707.395 1961.615 ;
        RECT 2708.485 1960.845 2708.775 1961.570 ;
        RECT 2710.530 1961.390 2710.870 1962.220 ;
        RECT 2716.050 1961.390 2716.390 1962.220 ;
        RECT 2721.570 1961.390 2721.910 1962.220 ;
        RECT 2727.090 1961.390 2727.430 1962.220 ;
        RECT 2731.025 1961.615 2731.775 1962.135 ;
        RECT 2708.945 1960.845 2714.290 1961.390 ;
        RECT 2714.465 1960.845 2719.810 1961.390 ;
        RECT 2719.985 1960.845 2725.330 1961.390 ;
        RECT 2725.505 1960.845 2730.850 1961.390 ;
        RECT 2731.025 1960.845 2732.695 1961.615 ;
        RECT 2733.555 1961.595 2734.075 1962.135 ;
        RECT 2732.865 1960.845 2734.075 1961.595 ;
        RECT 2695.520 1960.675 2734.160 1960.845 ;
        RECT 2695.605 1959.925 2696.815 1960.675 ;
        RECT 2696.985 1960.130 2702.330 1960.675 ;
        RECT 2702.505 1960.130 2707.850 1960.675 ;
        RECT 2708.025 1960.130 2713.370 1960.675 ;
        RECT 2713.545 1960.130 2718.890 1960.675 ;
        RECT 2695.605 1959.385 2696.125 1959.925 ;
        RECT 2698.570 1959.300 2698.910 1960.130 ;
        RECT 2704.090 1959.300 2704.430 1960.130 ;
        RECT 2709.610 1959.300 2709.950 1960.130 ;
        RECT 2715.130 1959.300 2715.470 1960.130 ;
        RECT 2719.065 1959.905 2720.735 1960.675 ;
        RECT 2721.365 1959.950 2721.655 1960.675 ;
        RECT 2721.825 1960.130 2727.170 1960.675 ;
        RECT 2727.345 1960.130 2732.690 1960.675 ;
        RECT 2719.065 1959.385 2719.815 1959.905 ;
        RECT 2723.410 1959.300 2723.750 1960.130 ;
        RECT 2728.930 1959.300 2729.270 1960.130 ;
        RECT 2732.865 1959.925 2734.075 1960.675 ;
        RECT 2733.555 1959.385 2734.075 1959.925 ;
        RECT 2523.330 1956.685 2523.670 1957.345 ;
        RECT 2522.130 1956.515 2523.935 1956.685 ;
        RECT 2695.605 1956.155 2696.125 1956.695 ;
        RECT 2343.005 1953.865 2453.605 1955.465 ;
        RECT 2695.605 1955.405 2696.815 1956.155 ;
        RECT 2699.950 1955.950 2700.290 1956.780 ;
        RECT 2703.885 1956.175 2705.535 1956.695 ;
        RECT 2697.425 1955.405 2697.755 1955.785 ;
        RECT 2698.365 1955.405 2703.710 1955.950 ;
        RECT 2703.885 1955.405 2707.395 1956.175 ;
        RECT 2708.485 1955.405 2708.775 1956.130 ;
        RECT 2710.530 1955.950 2710.870 1956.780 ;
        RECT 2716.050 1955.950 2716.390 1956.780 ;
        RECT 2721.570 1955.950 2721.910 1956.780 ;
        RECT 2727.090 1955.950 2727.430 1956.780 ;
        RECT 2731.025 1956.175 2731.775 1956.695 ;
        RECT 2708.945 1955.405 2714.290 1955.950 ;
        RECT 2714.465 1955.405 2719.810 1955.950 ;
        RECT 2719.985 1955.405 2725.330 1955.950 ;
        RECT 2725.505 1955.405 2730.850 1955.950 ;
        RECT 2731.025 1955.405 2732.695 1956.175 ;
        RECT 2733.555 1956.155 2734.075 1956.695 ;
        RECT 2732.865 1955.405 2734.075 1956.155 ;
        RECT 2695.520 1955.235 2734.160 1955.405 ;
        RECT 2695.605 1954.485 2696.815 1955.235 ;
        RECT 2696.985 1954.690 2702.330 1955.235 ;
        RECT 2702.505 1954.690 2707.850 1955.235 ;
        RECT 2708.025 1954.690 2713.370 1955.235 ;
        RECT 2713.545 1954.690 2718.890 1955.235 ;
        RECT 2695.605 1953.945 2696.125 1954.485 ;
        RECT 2358.220 1953.240 2358.390 1953.865 ;
        RECT 2369.035 1953.240 2369.205 1953.865 ;
        RECT 2369.990 1953.320 2370.160 1953.600 ;
        RECT 2369.990 1953.150 2370.220 1953.320 ;
        RECT 2374.650 1953.240 2374.820 1953.865 ;
        RECT 2377.395 1953.235 2377.565 1953.865 ;
        RECT 2378.385 1953.235 2378.555 1953.865 ;
        RECT 2387.595 1953.240 2387.765 1953.865 ;
        RECT 2388.550 1953.320 2388.720 1953.600 ;
        RECT 2388.550 1953.150 2388.780 1953.320 ;
        RECT 2393.210 1953.240 2393.380 1953.865 ;
        RECT 2395.955 1953.235 2396.125 1953.865 ;
        RECT 2396.945 1953.235 2397.115 1953.865 ;
        RECT 2406.155 1953.240 2406.325 1953.865 ;
        RECT 2407.110 1953.320 2407.280 1953.600 ;
        RECT 2407.110 1953.150 2407.340 1953.320 ;
        RECT 2411.770 1953.240 2411.940 1953.865 ;
        RECT 2414.515 1953.235 2414.685 1953.865 ;
        RECT 2415.505 1953.235 2415.675 1953.865 ;
        RECT 2424.715 1953.240 2424.885 1953.865 ;
        RECT 2425.670 1953.320 2425.840 1953.600 ;
        RECT 2425.670 1953.150 2425.900 1953.320 ;
        RECT 2430.330 1953.240 2430.500 1953.865 ;
        RECT 2433.075 1953.235 2433.245 1953.865 ;
        RECT 2434.065 1953.235 2434.235 1953.865 ;
        RECT 2443.275 1953.240 2443.445 1953.865 ;
        RECT 2444.230 1953.320 2444.400 1953.600 ;
        RECT 2444.230 1953.150 2444.460 1953.320 ;
        RECT 2448.890 1953.240 2449.060 1953.865 ;
        RECT 2451.635 1953.235 2451.805 1953.865 ;
        RECT 2452.625 1953.235 2452.795 1953.865 ;
        RECT 2698.570 1953.860 2698.910 1954.690 ;
        RECT 2704.090 1953.860 2704.430 1954.690 ;
        RECT 2709.610 1953.860 2709.950 1954.690 ;
        RECT 2715.130 1953.860 2715.470 1954.690 ;
        RECT 2719.065 1954.465 2720.735 1955.235 ;
        RECT 2721.365 1954.510 2721.655 1955.235 ;
        RECT 2721.825 1954.690 2727.170 1955.235 ;
        RECT 2727.345 1954.690 2732.690 1955.235 ;
        RECT 2719.065 1953.945 2719.815 1954.465 ;
        RECT 2723.410 1953.860 2723.750 1954.690 ;
        RECT 2728.930 1953.860 2729.270 1954.690 ;
        RECT 2732.865 1954.485 2734.075 1955.235 ;
        RECT 2733.555 1953.945 2734.075 1954.485 ;
        RECT 2370.050 1951.540 2370.220 1953.150 ;
        RECT 2388.610 1951.540 2388.780 1953.150 ;
        RECT 2407.170 1951.540 2407.340 1953.150 ;
        RECT 2425.730 1951.540 2425.900 1953.150 ;
        RECT 2444.290 1951.540 2444.460 1953.150 ;
        RECT 2369.990 1951.370 2370.220 1951.540 ;
        RECT 2388.550 1951.370 2388.780 1951.540 ;
        RECT 2407.110 1951.370 2407.340 1951.540 ;
        RECT 2425.670 1951.370 2425.900 1951.540 ;
        RECT 2444.230 1951.370 2444.460 1951.540 ;
        RECT 2369.990 1950.310 2370.160 1951.370 ;
        RECT 2388.550 1950.310 2388.720 1951.370 ;
        RECT 2407.110 1950.310 2407.280 1951.370 ;
        RECT 2425.670 1950.310 2425.840 1951.370 ;
        RECT 2444.230 1950.310 2444.400 1951.370 ;
        RECT 2523.330 1950.680 2523.670 1951.340 ;
        RECT 2695.605 1950.715 2696.125 1951.255 ;
        RECT 2522.130 1950.510 2523.935 1950.680 ;
        RECT 2695.605 1949.965 2696.815 1950.715 ;
        RECT 2701.330 1950.510 2701.670 1951.340 ;
        RECT 2705.265 1950.735 2706.475 1951.255 ;
        RECT 2697.425 1949.965 2697.755 1950.345 ;
        RECT 2698.805 1949.965 2699.135 1950.345 ;
        RECT 2699.745 1949.965 2705.090 1950.510 ;
        RECT 2705.265 1949.965 2707.855 1950.735 ;
        RECT 2708.485 1949.965 2708.775 1950.690 ;
        RECT 2710.530 1950.510 2710.870 1951.340 ;
        RECT 2716.050 1950.510 2716.390 1951.340 ;
        RECT 2719.985 1950.715 2720.505 1951.255 ;
        RECT 2708.945 1949.965 2714.290 1950.510 ;
        RECT 2714.465 1949.965 2719.810 1950.510 ;
        RECT 2719.985 1949.965 2721.195 1950.715 ;
        RECT 2721.365 1949.965 2721.655 1950.690 ;
        RECT 2723.410 1950.510 2723.750 1951.340 ;
        RECT 2728.930 1950.510 2729.270 1951.340 ;
        RECT 2733.555 1950.715 2734.075 1951.255 ;
        RECT 2721.825 1949.965 2727.170 1950.510 ;
        RECT 2727.345 1949.965 2732.690 1950.510 ;
        RECT 2732.865 1949.965 2734.075 1950.715 ;
        RECT 2695.520 1949.795 2734.160 1949.965 ;
        RECT 2363.195 1947.345 2363.485 1947.515 ;
        RECT 2381.755 1947.345 2382.045 1947.515 ;
        RECT 2400.315 1947.345 2400.605 1947.515 ;
        RECT 2418.875 1947.345 2419.165 1947.515 ;
        RECT 2437.435 1947.345 2437.725 1947.515 ;
        RECT 2363.195 1947.035 2363.365 1947.345 ;
        RECT 2362.995 1946.865 2363.365 1947.035 ;
        RECT 2365.035 1946.785 2365.205 1947.115 ;
        RECT 2381.755 1947.035 2381.925 1947.345 ;
        RECT 2381.555 1946.865 2381.925 1947.035 ;
        RECT 2383.595 1946.785 2383.765 1947.115 ;
        RECT 2400.315 1947.035 2400.485 1947.345 ;
        RECT 2400.115 1946.865 2400.485 1947.035 ;
        RECT 2402.155 1946.785 2402.325 1947.115 ;
        RECT 2418.875 1947.035 2419.045 1947.345 ;
        RECT 2418.675 1946.865 2419.045 1947.035 ;
        RECT 2420.715 1946.785 2420.885 1947.115 ;
        RECT 2437.435 1947.035 2437.605 1947.345 ;
        RECT 2437.235 1946.865 2437.605 1947.035 ;
        RECT 2439.275 1946.785 2439.445 1947.115 ;
        RECT 2362.355 1945.875 2362.525 1946.375 ;
        RECT 2363.835 1945.875 2364.005 1946.375 ;
        RECT 2365.755 1945.875 2365.925 1946.375 ;
        RECT 2367.235 1945.875 2367.405 1946.375 ;
        RECT 2368.195 1945.875 2368.365 1946.375 ;
        RECT 2369.195 1945.875 2369.365 1946.375 ;
        RECT 2370.155 1945.875 2370.325 1946.375 ;
        RECT 2370.675 1945.875 2370.845 1946.375 ;
        RECT 2371.635 1945.875 2371.805 1946.375 ;
        RECT 2372.595 1945.875 2372.765 1946.375 ;
        RECT 2380.915 1945.875 2381.085 1946.375 ;
        RECT 2382.395 1945.875 2382.565 1946.375 ;
        RECT 2384.315 1945.875 2384.485 1946.375 ;
        RECT 2385.795 1945.875 2385.965 1946.375 ;
        RECT 2386.755 1945.875 2386.925 1946.375 ;
        RECT 2387.755 1945.875 2387.925 1946.375 ;
        RECT 2388.715 1945.875 2388.885 1946.375 ;
        RECT 2389.235 1945.875 2389.405 1946.375 ;
        RECT 2390.195 1945.875 2390.365 1946.375 ;
        RECT 2391.155 1945.875 2391.325 1946.375 ;
        RECT 2399.475 1945.875 2399.645 1946.375 ;
        RECT 2400.955 1945.875 2401.125 1946.375 ;
        RECT 2402.875 1945.875 2403.045 1946.375 ;
        RECT 2404.355 1945.875 2404.525 1946.375 ;
        RECT 2405.315 1945.875 2405.485 1946.375 ;
        RECT 2406.315 1945.875 2406.485 1946.375 ;
        RECT 2407.275 1945.875 2407.445 1946.375 ;
        RECT 2407.795 1945.875 2407.965 1946.375 ;
        RECT 2408.755 1945.875 2408.925 1946.375 ;
        RECT 2409.715 1945.875 2409.885 1946.375 ;
        RECT 2418.035 1945.875 2418.205 1946.375 ;
        RECT 2419.515 1945.875 2419.685 1946.375 ;
        RECT 2421.435 1945.875 2421.605 1946.375 ;
        RECT 2422.915 1945.875 2423.085 1946.375 ;
        RECT 2423.875 1945.875 2424.045 1946.375 ;
        RECT 2424.875 1945.875 2425.045 1946.375 ;
        RECT 2425.835 1945.875 2426.005 1946.375 ;
        RECT 2426.355 1945.875 2426.525 1946.375 ;
        RECT 2427.315 1945.875 2427.485 1946.375 ;
        RECT 2428.275 1945.875 2428.445 1946.375 ;
        RECT 2436.595 1945.875 2436.765 1946.375 ;
        RECT 2438.075 1945.875 2438.245 1946.375 ;
        RECT 2439.995 1945.875 2440.165 1946.375 ;
        RECT 2441.475 1945.875 2441.645 1946.375 ;
        RECT 2442.435 1945.875 2442.605 1946.375 ;
        RECT 2443.435 1945.875 2443.605 1946.375 ;
        RECT 2444.395 1945.875 2444.565 1946.375 ;
        RECT 2444.915 1945.875 2445.085 1946.375 ;
        RECT 2445.875 1945.875 2446.045 1946.375 ;
        RECT 2446.835 1945.875 2447.005 1946.375 ;
        RECT 2361.545 1944.600 2373.590 1945.875 ;
        RECT 2374.650 1944.600 2374.820 1945.225 ;
        RECT 2377.395 1944.600 2377.565 1945.230 ;
        RECT 2378.380 1944.600 2378.550 1945.230 ;
        RECT 2380.105 1944.600 2392.150 1945.875 ;
        RECT 2393.210 1944.600 2393.380 1945.225 ;
        RECT 2395.955 1944.600 2396.125 1945.230 ;
        RECT 2396.940 1944.600 2397.110 1945.230 ;
        RECT 2398.665 1944.600 2410.710 1945.875 ;
        RECT 2411.770 1944.600 2411.940 1945.225 ;
        RECT 2414.515 1944.600 2414.685 1945.230 ;
        RECT 2415.500 1944.600 2415.670 1945.230 ;
        RECT 2417.225 1944.600 2429.270 1945.875 ;
        RECT 2430.330 1944.600 2430.500 1945.225 ;
        RECT 2433.075 1944.600 2433.245 1945.230 ;
        RECT 2434.060 1944.600 2434.230 1945.230 ;
        RECT 2435.785 1944.600 2447.830 1945.875 ;
        RECT 2448.890 1944.600 2449.060 1945.225 ;
        RECT 2451.635 1944.600 2451.805 1945.230 ;
        RECT 2452.620 1944.600 2452.790 1945.230 ;
        RECT 2343.005 1943.000 2453.600 1944.600 ;
        RECT 2882.265 1891.670 2882.605 1892.330 ;
        RECT 2881.575 1891.500 2883.380 1891.670 ;
        RECT 2695.520 1856.835 2734.160 1857.005 ;
        RECT 2695.605 1856.085 2696.815 1856.835 ;
        RECT 2697.455 1856.355 2697.730 1856.835 ;
        RECT 2698.315 1856.435 2698.650 1856.835 ;
        RECT 2699.265 1856.455 2699.595 1856.835 ;
        RECT 2700.645 1856.455 2700.975 1856.835 ;
        RECT 2701.585 1856.290 2706.930 1856.835 ;
        RECT 2695.605 1855.545 2696.125 1856.085 ;
        RECT 2703.170 1855.460 2703.510 1856.290 ;
        RECT 2707.105 1856.085 2708.315 1856.835 ;
        RECT 2708.485 1856.110 2708.775 1856.835 ;
        RECT 2709.420 1856.455 2709.750 1856.835 ;
        RECT 2707.105 1855.545 2707.625 1856.085 ;
        RECT 2710.350 1855.995 2710.610 1856.835 ;
        RECT 2710.785 1856.290 2716.130 1856.835 ;
        RECT 2712.370 1855.460 2712.710 1856.290 ;
        RECT 2716.305 1856.065 2719.815 1856.835 ;
        RECT 2719.985 1856.085 2721.195 1856.835 ;
        RECT 2721.365 1856.110 2721.655 1856.835 ;
        RECT 2721.830 1856.435 2722.165 1856.835 ;
        RECT 2722.750 1856.355 2723.025 1856.835 ;
        RECT 2723.665 1856.290 2729.010 1856.835 ;
        RECT 2716.305 1855.545 2717.955 1856.065 ;
        RECT 2719.985 1855.545 2720.505 1856.085 ;
        RECT 2725.250 1855.460 2725.590 1856.290 ;
        RECT 2729.185 1856.065 2730.855 1856.835 ;
        RECT 2731.925 1856.455 2732.255 1856.835 ;
        RECT 2732.865 1856.085 2734.075 1856.835 ;
        RECT 2729.185 1855.545 2729.935 1856.065 ;
        RECT 2733.555 1855.545 2734.075 1856.085 ;
        RECT 2695.605 1852.315 2696.125 1852.855 ;
        RECT 2695.605 1851.565 2696.815 1852.315 ;
        RECT 2699.950 1852.110 2700.290 1852.940 ;
        RECT 2703.885 1852.335 2705.535 1852.855 ;
        RECT 2697.425 1851.565 2697.755 1851.945 ;
        RECT 2698.365 1851.565 2703.710 1852.110 ;
        RECT 2703.885 1851.565 2707.395 1852.335 ;
        RECT 2708.485 1851.565 2708.775 1852.290 ;
        RECT 2710.530 1852.110 2710.870 1852.940 ;
        RECT 2716.050 1852.110 2716.390 1852.940 ;
        RECT 2721.570 1852.110 2721.910 1852.940 ;
        RECT 2727.090 1852.110 2727.430 1852.940 ;
        RECT 2731.025 1852.335 2731.775 1852.855 ;
        RECT 2708.945 1851.565 2714.290 1852.110 ;
        RECT 2714.465 1851.565 2719.810 1852.110 ;
        RECT 2719.985 1851.565 2725.330 1852.110 ;
        RECT 2725.505 1851.565 2730.850 1852.110 ;
        RECT 2731.025 1851.565 2732.695 1852.335 ;
        RECT 2733.555 1852.315 2734.075 1852.855 ;
        RECT 2732.865 1851.565 2734.075 1852.315 ;
        RECT 2695.520 1851.395 2734.160 1851.565 ;
        RECT 2695.605 1850.645 2696.815 1851.395 ;
        RECT 2696.985 1850.850 2702.330 1851.395 ;
        RECT 2702.505 1850.850 2707.850 1851.395 ;
        RECT 2708.025 1850.850 2713.370 1851.395 ;
        RECT 2713.545 1850.850 2718.890 1851.395 ;
        RECT 2695.605 1850.105 2696.125 1850.645 ;
        RECT 2698.570 1850.020 2698.910 1850.850 ;
        RECT 2704.090 1850.020 2704.430 1850.850 ;
        RECT 2709.610 1850.020 2709.950 1850.850 ;
        RECT 2715.130 1850.020 2715.470 1850.850 ;
        RECT 2719.065 1850.625 2720.735 1851.395 ;
        RECT 2721.365 1850.670 2721.655 1851.395 ;
        RECT 2721.825 1850.850 2727.170 1851.395 ;
        RECT 2727.345 1850.850 2732.690 1851.395 ;
        RECT 2719.065 1850.105 2719.815 1850.625 ;
        RECT 2723.410 1850.020 2723.750 1850.850 ;
        RECT 2728.930 1850.020 2729.270 1850.850 ;
        RECT 2732.865 1850.645 2734.075 1851.395 ;
        RECT 2733.555 1850.105 2734.075 1850.645 ;
        RECT 2695.605 1846.875 2696.125 1847.415 ;
        RECT 2695.605 1846.125 2696.815 1846.875 ;
        RECT 2698.570 1846.670 2698.910 1847.500 ;
        RECT 2704.090 1846.670 2704.430 1847.500 ;
        RECT 2696.985 1846.125 2702.330 1846.670 ;
        RECT 2702.505 1846.125 2707.850 1846.670 ;
        RECT 2708.485 1846.125 2708.775 1846.850 ;
        RECT 2710.530 1846.670 2710.870 1847.500 ;
        RECT 2716.050 1846.670 2716.390 1847.500 ;
        RECT 2721.570 1846.670 2721.910 1847.500 ;
        RECT 2727.090 1846.670 2727.430 1847.500 ;
        RECT 2731.025 1846.895 2731.775 1847.415 ;
        RECT 2708.945 1846.125 2714.290 1846.670 ;
        RECT 2714.465 1846.125 2719.810 1846.670 ;
        RECT 2719.985 1846.125 2725.330 1846.670 ;
        RECT 2725.505 1846.125 2730.850 1846.670 ;
        RECT 2731.025 1846.125 2732.695 1846.895 ;
        RECT 2733.555 1846.875 2734.075 1847.415 ;
        RECT 2732.865 1846.125 2734.075 1846.875 ;
        RECT 2695.520 1845.955 2734.160 1846.125 ;
        RECT 2695.605 1845.205 2696.815 1845.955 ;
        RECT 2697.425 1845.575 2697.755 1845.955 ;
        RECT 2698.365 1845.410 2703.710 1845.955 ;
        RECT 2703.885 1845.410 2709.230 1845.955 ;
        RECT 2709.405 1845.410 2714.750 1845.955 ;
        RECT 2714.925 1845.410 2720.270 1845.955 ;
        RECT 2695.605 1844.665 2696.125 1845.205 ;
        RECT 2699.950 1844.580 2700.290 1845.410 ;
        RECT 2705.470 1844.580 2705.810 1845.410 ;
        RECT 2710.990 1844.580 2711.330 1845.410 ;
        RECT 2716.510 1844.580 2716.850 1845.410 ;
        RECT 2721.365 1845.230 2721.655 1845.955 ;
        RECT 2721.825 1845.410 2727.170 1845.955 ;
        RECT 2727.345 1845.410 2732.690 1845.955 ;
        RECT 2723.410 1844.580 2723.750 1845.410 ;
        RECT 2728.930 1844.580 2729.270 1845.410 ;
        RECT 2732.865 1845.205 2734.075 1845.955 ;
        RECT 2733.555 1844.665 2734.075 1845.205 ;
        RECT 2695.605 1841.435 2696.125 1841.975 ;
        RECT 2695.605 1840.685 2696.815 1841.435 ;
        RECT 2698.570 1841.230 2698.910 1842.060 ;
        RECT 2704.090 1841.230 2704.430 1842.060 ;
        RECT 2696.985 1840.685 2702.330 1841.230 ;
        RECT 2702.505 1840.685 2707.850 1841.230 ;
        RECT 2708.485 1840.685 2708.775 1841.410 ;
        RECT 2710.530 1841.230 2710.870 1842.060 ;
        RECT 2716.050 1841.230 2716.390 1842.060 ;
        RECT 2721.570 1841.230 2721.910 1842.060 ;
        RECT 2727.090 1841.230 2727.430 1842.060 ;
        RECT 2731.025 1841.455 2731.775 1841.975 ;
        RECT 2708.945 1840.685 2714.290 1841.230 ;
        RECT 2714.465 1840.685 2719.810 1841.230 ;
        RECT 2719.985 1840.685 2725.330 1841.230 ;
        RECT 2725.505 1840.685 2730.850 1841.230 ;
        RECT 2731.025 1840.685 2732.695 1841.455 ;
        RECT 2733.555 1841.435 2734.075 1841.975 ;
        RECT 2732.865 1840.685 2734.075 1841.435 ;
        RECT 2695.520 1840.515 2734.160 1840.685 ;
        RECT 2695.605 1839.765 2696.815 1840.515 ;
        RECT 2697.415 1840.135 2697.745 1840.515 ;
        RECT 2699.700 1839.795 2699.990 1840.515 ;
        RECT 2702.050 1840.055 2702.220 1840.515 ;
        RECT 2702.910 1840.135 2703.240 1840.515 ;
        RECT 2705.795 1840.055 2705.965 1840.515 ;
        RECT 2706.645 1839.970 2711.990 1840.515 ;
        RECT 2712.165 1839.970 2717.510 1840.515 ;
        RECT 2695.605 1839.225 2696.125 1839.765 ;
        RECT 2708.230 1839.140 2708.570 1839.970 ;
        RECT 2713.750 1839.140 2714.090 1839.970 ;
        RECT 2717.685 1839.745 2721.195 1840.515 ;
        RECT 2721.365 1839.790 2721.655 1840.515 ;
        RECT 2721.825 1839.970 2727.170 1840.515 ;
        RECT 2727.345 1839.970 2732.690 1840.515 ;
        RECT 2717.685 1839.225 2719.335 1839.745 ;
        RECT 2723.410 1839.140 2723.750 1839.970 ;
        RECT 2728.930 1839.140 2729.270 1839.970 ;
        RECT 2732.865 1839.765 2734.075 1840.515 ;
        RECT 2733.555 1839.225 2734.075 1839.765 ;
        RECT 2695.605 1835.995 2696.125 1836.535 ;
        RECT 2695.605 1835.245 2696.815 1835.995 ;
        RECT 2699.950 1835.790 2700.290 1836.620 ;
        RECT 2703.885 1836.015 2705.535 1836.535 ;
        RECT 2697.425 1835.245 2697.755 1835.625 ;
        RECT 2698.365 1835.245 2703.710 1835.790 ;
        RECT 2703.885 1835.245 2707.395 1836.015 ;
        RECT 2708.485 1835.245 2708.775 1835.970 ;
        RECT 2710.530 1835.790 2710.870 1836.620 ;
        RECT 2716.050 1835.790 2716.390 1836.620 ;
        RECT 2721.570 1835.790 2721.910 1836.620 ;
        RECT 2727.090 1835.790 2727.430 1836.620 ;
        RECT 2731.025 1836.015 2731.775 1836.535 ;
        RECT 2708.945 1835.245 2714.290 1835.790 ;
        RECT 2714.465 1835.245 2719.810 1835.790 ;
        RECT 2719.985 1835.245 2725.330 1835.790 ;
        RECT 2725.505 1835.245 2730.850 1835.790 ;
        RECT 2731.025 1835.245 2732.695 1836.015 ;
        RECT 2733.555 1835.995 2734.075 1836.535 ;
        RECT 2732.865 1835.245 2734.075 1835.995 ;
        RECT 2695.520 1835.075 2734.160 1835.245 ;
        RECT 2695.605 1834.325 2696.815 1835.075 ;
        RECT 2697.415 1834.695 2697.745 1835.075 ;
        RECT 2699.700 1834.355 2699.990 1835.075 ;
        RECT 2702.050 1834.615 2702.220 1835.075 ;
        RECT 2702.910 1834.695 2703.240 1835.075 ;
        RECT 2705.795 1834.615 2705.965 1835.075 ;
        RECT 2706.645 1834.530 2711.990 1835.075 ;
        RECT 2712.165 1834.530 2717.510 1835.075 ;
        RECT 2695.605 1833.785 2696.125 1834.325 ;
        RECT 2708.230 1833.700 2708.570 1834.530 ;
        RECT 2713.750 1833.700 2714.090 1834.530 ;
        RECT 2717.685 1834.305 2721.195 1835.075 ;
        RECT 2721.365 1834.350 2721.655 1835.075 ;
        RECT 2721.825 1834.530 2727.170 1835.075 ;
        RECT 2727.345 1834.530 2732.690 1835.075 ;
        RECT 2717.685 1833.785 2719.335 1834.305 ;
        RECT 2723.410 1833.700 2723.750 1834.530 ;
        RECT 2728.930 1833.700 2729.270 1834.530 ;
        RECT 2732.865 1834.325 2734.075 1835.075 ;
        RECT 2733.555 1833.785 2734.075 1834.325 ;
        RECT 2695.605 1830.555 2696.125 1831.095 ;
        RECT 2698.365 1830.575 2699.575 1831.095 ;
        RECT 2705.725 1830.575 2706.935 1831.095 ;
        RECT 2695.605 1829.805 2696.815 1830.555 ;
        RECT 2697.425 1829.805 2697.755 1830.185 ;
        RECT 2698.365 1829.805 2700.955 1830.575 ;
        RECT 2702.015 1829.805 2702.345 1830.205 ;
        RECT 2704.305 1829.805 2704.815 1830.340 ;
        RECT 2705.725 1829.805 2708.315 1830.575 ;
        RECT 2708.485 1829.805 2708.775 1830.530 ;
        RECT 2710.530 1830.350 2710.870 1831.180 ;
        RECT 2716.050 1830.350 2716.390 1831.180 ;
        RECT 2721.570 1830.350 2721.910 1831.180 ;
        RECT 2727.090 1830.350 2727.430 1831.180 ;
        RECT 2731.025 1830.575 2731.775 1831.095 ;
        RECT 2708.945 1829.805 2714.290 1830.350 ;
        RECT 2714.465 1829.805 2719.810 1830.350 ;
        RECT 2719.985 1829.805 2725.330 1830.350 ;
        RECT 2725.505 1829.805 2730.850 1830.350 ;
        RECT 2731.025 1829.805 2732.695 1830.575 ;
        RECT 2733.555 1830.555 2734.075 1831.095 ;
        RECT 2732.865 1829.805 2734.075 1830.555 ;
        RECT 2695.520 1829.635 2734.160 1829.805 ;
        RECT 2695.605 1828.885 2696.815 1829.635 ;
        RECT 2696.985 1829.090 2702.330 1829.635 ;
        RECT 2702.505 1829.090 2707.850 1829.635 ;
        RECT 2708.025 1829.090 2713.370 1829.635 ;
        RECT 2713.545 1829.090 2718.890 1829.635 ;
        RECT 2695.605 1828.345 2696.125 1828.885 ;
        RECT 2698.570 1828.260 2698.910 1829.090 ;
        RECT 2704.090 1828.260 2704.430 1829.090 ;
        RECT 2709.610 1828.260 2709.950 1829.090 ;
        RECT 2715.130 1828.260 2715.470 1829.090 ;
        RECT 2719.065 1828.865 2720.735 1829.635 ;
        RECT 2721.365 1828.910 2721.655 1829.635 ;
        RECT 2721.825 1829.090 2727.170 1829.635 ;
        RECT 2727.345 1829.090 2732.690 1829.635 ;
        RECT 2719.065 1828.345 2719.815 1828.865 ;
        RECT 2723.410 1828.260 2723.750 1829.090 ;
        RECT 2728.930 1828.260 2729.270 1829.090 ;
        RECT 2732.865 1828.885 2734.075 1829.635 ;
        RECT 2733.555 1828.345 2734.075 1828.885 ;
        RECT 2695.605 1825.115 2696.125 1825.655 ;
        RECT 2695.605 1824.365 2696.815 1825.115 ;
        RECT 2699.950 1824.910 2700.290 1825.740 ;
        RECT 2703.885 1825.135 2705.535 1825.655 ;
        RECT 2697.425 1824.365 2697.755 1824.745 ;
        RECT 2698.365 1824.365 2703.710 1824.910 ;
        RECT 2703.885 1824.365 2707.395 1825.135 ;
        RECT 2708.485 1824.365 2708.775 1825.090 ;
        RECT 2710.530 1824.910 2710.870 1825.740 ;
        RECT 2716.050 1824.910 2716.390 1825.740 ;
        RECT 2721.570 1824.910 2721.910 1825.740 ;
        RECT 2727.090 1824.910 2727.430 1825.740 ;
        RECT 2731.025 1825.135 2731.775 1825.655 ;
        RECT 2708.945 1824.365 2714.290 1824.910 ;
        RECT 2714.465 1824.365 2719.810 1824.910 ;
        RECT 2719.985 1824.365 2725.330 1824.910 ;
        RECT 2725.505 1824.365 2730.850 1824.910 ;
        RECT 2731.025 1824.365 2732.695 1825.135 ;
        RECT 2733.555 1825.115 2734.075 1825.655 ;
        RECT 2732.865 1824.365 2734.075 1825.115 ;
        RECT 2695.520 1824.195 2734.160 1824.365 ;
        RECT 2695.605 1823.445 2696.815 1824.195 ;
        RECT 2696.985 1823.650 2702.330 1824.195 ;
        RECT 2702.505 1823.650 2707.850 1824.195 ;
        RECT 2708.025 1823.650 2713.370 1824.195 ;
        RECT 2713.545 1823.650 2718.890 1824.195 ;
        RECT 2695.605 1822.905 2696.125 1823.445 ;
        RECT 2698.570 1822.820 2698.910 1823.650 ;
        RECT 2704.090 1822.820 2704.430 1823.650 ;
        RECT 2709.610 1822.820 2709.950 1823.650 ;
        RECT 2715.130 1822.820 2715.470 1823.650 ;
        RECT 2719.065 1823.425 2720.735 1824.195 ;
        RECT 2721.365 1823.470 2721.655 1824.195 ;
        RECT 2721.825 1823.650 2727.170 1824.195 ;
        RECT 2727.345 1823.650 2732.690 1824.195 ;
        RECT 2719.065 1822.905 2719.815 1823.425 ;
        RECT 2723.410 1822.820 2723.750 1823.650 ;
        RECT 2728.930 1822.820 2729.270 1823.650 ;
        RECT 2732.865 1823.445 2734.075 1824.195 ;
        RECT 2733.555 1822.905 2734.075 1823.445 ;
        RECT 2695.605 1819.675 2696.125 1820.215 ;
        RECT 2696.985 1819.695 2698.635 1820.215 ;
        RECT 2695.605 1818.925 2696.815 1819.675 ;
        RECT 2696.985 1818.925 2700.495 1819.695 ;
        RECT 2701.605 1818.925 2701.845 1819.735 ;
        RECT 2702.515 1818.925 2702.785 1819.735 ;
        RECT 2704.550 1819.470 2704.890 1820.300 ;
        RECT 2702.965 1818.925 2708.310 1819.470 ;
        RECT 2708.485 1818.925 2708.775 1819.650 ;
        RECT 2710.530 1819.470 2710.870 1820.300 ;
        RECT 2716.050 1819.470 2716.390 1820.300 ;
        RECT 2721.570 1819.470 2721.910 1820.300 ;
        RECT 2727.090 1819.470 2727.430 1820.300 ;
        RECT 2731.025 1819.695 2731.775 1820.215 ;
        RECT 2708.945 1818.925 2714.290 1819.470 ;
        RECT 2714.465 1818.925 2719.810 1819.470 ;
        RECT 2719.985 1818.925 2725.330 1819.470 ;
        RECT 2725.505 1818.925 2730.850 1819.470 ;
        RECT 2731.025 1818.925 2732.695 1819.695 ;
        RECT 2733.555 1819.675 2734.075 1820.215 ;
        RECT 2732.865 1818.925 2734.075 1819.675 ;
        RECT 2695.520 1818.755 2734.160 1818.925 ;
        RECT 2695.605 1818.005 2696.815 1818.755 ;
        RECT 2697.425 1818.375 2697.755 1818.755 ;
        RECT 2695.605 1817.465 2696.125 1818.005 ;
        RECT 2698.365 1817.985 2701.875 1818.755 ;
        RECT 2702.055 1818.015 2702.385 1818.755 ;
        RECT 2703.090 1818.395 2703.420 1818.755 ;
        RECT 2698.365 1817.465 2700.015 1817.985 ;
        RECT 2704.785 1817.975 2705.080 1818.755 ;
        RECT 2705.265 1818.210 2710.610 1818.755 ;
        RECT 2710.785 1818.210 2716.130 1818.755 ;
        RECT 2706.850 1817.380 2707.190 1818.210 ;
        RECT 2712.370 1817.380 2712.710 1818.210 ;
        RECT 2716.305 1817.985 2719.815 1818.755 ;
        RECT 2719.985 1818.005 2721.195 1818.755 ;
        RECT 2721.365 1818.030 2721.655 1818.755 ;
        RECT 2721.825 1818.210 2727.170 1818.755 ;
        RECT 2727.345 1818.210 2732.690 1818.755 ;
        RECT 2716.305 1817.465 2717.955 1817.985 ;
        RECT 2719.985 1817.465 2720.505 1818.005 ;
        RECT 2723.410 1817.380 2723.750 1818.210 ;
        RECT 2728.930 1817.380 2729.270 1818.210 ;
        RECT 2732.865 1818.005 2734.075 1818.755 ;
        RECT 2733.555 1817.465 2734.075 1818.005 ;
        RECT 2695.605 1814.235 2696.125 1814.775 ;
        RECT 2695.605 1813.485 2696.815 1814.235 ;
        RECT 2698.570 1814.030 2698.910 1814.860 ;
        RECT 2704.090 1814.030 2704.430 1814.860 ;
        RECT 2696.985 1813.485 2702.330 1814.030 ;
        RECT 2702.505 1813.485 2707.850 1814.030 ;
        RECT 2708.485 1813.485 2708.775 1814.210 ;
        RECT 2710.530 1814.030 2710.870 1814.860 ;
        RECT 2716.050 1814.030 2716.390 1814.860 ;
        RECT 2721.570 1814.030 2721.910 1814.860 ;
        RECT 2708.945 1813.485 2714.290 1814.030 ;
        RECT 2714.465 1813.485 2719.810 1814.030 ;
        RECT 2719.985 1813.485 2725.330 1814.030 ;
        RECT 2725.515 1813.485 2725.845 1813.965 ;
        RECT 2726.355 1813.485 2726.685 1813.965 ;
        RECT 2727.195 1813.485 2727.525 1813.965 ;
        RECT 2728.035 1813.485 2728.365 1813.965 ;
        RECT 2728.875 1813.485 2729.205 1813.965 ;
        RECT 2729.715 1813.485 2730.045 1813.965 ;
        RECT 2730.555 1813.485 2730.885 1813.965 ;
        RECT 2731.395 1813.485 2731.725 1813.965 ;
        RECT 2732.235 1813.485 2732.565 1814.285 ;
        RECT 2733.555 1814.235 2734.075 1814.775 ;
        RECT 2732.865 1813.485 2734.075 1814.235 ;
        RECT 2695.520 1813.315 2734.160 1813.485 ;
        RECT 2695.605 1812.565 2696.815 1813.315 ;
        RECT 2697.425 1812.935 2697.755 1813.315 ;
        RECT 2698.365 1812.770 2703.710 1813.315 ;
        RECT 2703.885 1812.770 2709.230 1813.315 ;
        RECT 2709.405 1812.770 2714.750 1813.315 ;
        RECT 2714.925 1812.770 2720.270 1813.315 ;
        RECT 2695.605 1812.025 2696.125 1812.565 ;
        RECT 2699.950 1811.940 2700.290 1812.770 ;
        RECT 2705.470 1811.940 2705.810 1812.770 ;
        RECT 2710.990 1811.940 2711.330 1812.770 ;
        RECT 2716.510 1811.940 2716.850 1812.770 ;
        RECT 2721.365 1812.590 2721.655 1813.315 ;
        RECT 2721.825 1812.770 2727.170 1813.315 ;
        RECT 2727.345 1812.770 2732.690 1813.315 ;
        RECT 2723.410 1811.940 2723.750 1812.770 ;
        RECT 2728.930 1811.940 2729.270 1812.770 ;
        RECT 2732.865 1812.565 2734.075 1813.315 ;
        RECT 2733.555 1812.025 2734.075 1812.565 ;
        RECT 2695.605 1808.795 2696.125 1809.335 ;
        RECT 2695.605 1808.045 2696.815 1808.795 ;
        RECT 2698.570 1808.590 2698.910 1809.420 ;
        RECT 2704.090 1808.590 2704.430 1809.420 ;
        RECT 2696.985 1808.045 2702.330 1808.590 ;
        RECT 2702.505 1808.045 2707.850 1808.590 ;
        RECT 2708.485 1808.045 2708.775 1808.770 ;
        RECT 2710.530 1808.590 2710.870 1809.420 ;
        RECT 2716.050 1808.590 2716.390 1809.420 ;
        RECT 2721.570 1808.590 2721.910 1809.420 ;
        RECT 2727.090 1808.590 2727.430 1809.420 ;
        RECT 2731.025 1808.815 2731.775 1809.335 ;
        RECT 2708.945 1808.045 2714.290 1808.590 ;
        RECT 2714.465 1808.045 2719.810 1808.590 ;
        RECT 2719.985 1808.045 2725.330 1808.590 ;
        RECT 2725.505 1808.045 2730.850 1808.590 ;
        RECT 2731.025 1808.045 2732.695 1808.815 ;
        RECT 2733.555 1808.795 2734.075 1809.335 ;
        RECT 2732.865 1808.045 2734.075 1808.795 ;
        RECT 2695.520 1807.875 2734.160 1808.045 ;
        RECT 2695.605 1807.125 2696.815 1807.875 ;
        RECT 2697.715 1807.135 2698.045 1807.875 ;
        RECT 2698.555 1807.475 2698.885 1807.875 ;
        RECT 2699.745 1807.330 2705.090 1807.875 ;
        RECT 2705.265 1807.330 2710.610 1807.875 ;
        RECT 2710.785 1807.330 2716.130 1807.875 ;
        RECT 2695.605 1806.585 2696.125 1807.125 ;
        RECT 2701.330 1806.500 2701.670 1807.330 ;
        RECT 2706.850 1806.500 2707.190 1807.330 ;
        RECT 2712.370 1806.500 2712.710 1807.330 ;
        RECT 2716.305 1807.105 2719.815 1807.875 ;
        RECT 2719.985 1807.125 2721.195 1807.875 ;
        RECT 2721.365 1807.150 2721.655 1807.875 ;
        RECT 2721.825 1807.330 2727.170 1807.875 ;
        RECT 2727.345 1807.330 2732.690 1807.875 ;
        RECT 2716.305 1806.585 2717.955 1807.105 ;
        RECT 2719.985 1806.585 2720.505 1807.125 ;
        RECT 2723.410 1806.500 2723.750 1807.330 ;
        RECT 2728.930 1806.500 2729.270 1807.330 ;
        RECT 2732.865 1807.125 2734.075 1807.875 ;
        RECT 2733.555 1806.585 2734.075 1807.125 ;
        RECT 2523.330 1804.815 2523.670 1805.475 ;
        RECT 2522.130 1804.645 2523.935 1804.815 ;
        RECT 2695.605 1803.355 2696.125 1803.895 ;
        RECT 2695.605 1802.605 2696.815 1803.355 ;
        RECT 2699.950 1803.150 2700.290 1803.980 ;
        RECT 2703.885 1803.375 2705.535 1803.895 ;
        RECT 2697.425 1802.605 2697.755 1802.985 ;
        RECT 2698.365 1802.605 2703.710 1803.150 ;
        RECT 2703.885 1802.605 2707.395 1803.375 ;
        RECT 2708.485 1802.605 2708.775 1803.330 ;
        RECT 2710.530 1803.150 2710.870 1803.980 ;
        RECT 2716.050 1803.150 2716.390 1803.980 ;
        RECT 2721.570 1803.150 2721.910 1803.980 ;
        RECT 2727.090 1803.150 2727.430 1803.980 ;
        RECT 2731.025 1803.375 2731.775 1803.895 ;
        RECT 2708.945 1802.605 2714.290 1803.150 ;
        RECT 2714.465 1802.605 2719.810 1803.150 ;
        RECT 2719.985 1802.605 2725.330 1803.150 ;
        RECT 2725.505 1802.605 2730.850 1803.150 ;
        RECT 2731.025 1802.605 2732.695 1803.375 ;
        RECT 2733.555 1803.355 2734.075 1803.895 ;
        RECT 2732.865 1802.605 2734.075 1803.355 ;
        RECT 2695.520 1802.435 2734.160 1802.605 ;
        RECT 2695.605 1801.685 2696.815 1802.435 ;
        RECT 2697.725 1801.900 2698.235 1802.435 ;
        RECT 2700.195 1802.035 2700.525 1802.435 ;
        RECT 2701.210 1801.760 2701.450 1802.435 ;
        RECT 2702.840 1801.985 2703.170 1802.435 ;
        RECT 2704.090 1801.995 2704.405 1802.435 ;
        RECT 2704.805 1801.890 2710.150 1802.435 ;
        RECT 2710.325 1801.890 2715.670 1802.435 ;
        RECT 2715.845 1801.890 2721.190 1802.435 ;
        RECT 2695.605 1801.145 2696.125 1801.685 ;
        RECT 2706.390 1801.060 2706.730 1801.890 ;
        RECT 2711.910 1801.060 2712.250 1801.890 ;
        RECT 2717.430 1801.060 2717.770 1801.890 ;
        RECT 2721.365 1801.710 2721.655 1802.435 ;
        RECT 2721.825 1801.890 2727.170 1802.435 ;
        RECT 2727.345 1801.890 2732.690 1802.435 ;
        RECT 2723.410 1801.060 2723.750 1801.890 ;
        RECT 2728.930 1801.060 2729.270 1801.890 ;
        RECT 2732.865 1801.685 2734.075 1802.435 ;
        RECT 2733.555 1801.145 2734.075 1801.685 ;
        RECT 2523.330 1797.285 2523.670 1797.945 ;
        RECT 2695.605 1797.915 2696.125 1798.455 ;
        RECT 2522.130 1797.115 2523.935 1797.285 ;
        RECT 2695.605 1797.165 2696.815 1797.915 ;
        RECT 2696.985 1797.165 2697.245 1797.985 ;
        RECT 2701.790 1797.710 2702.130 1798.540 ;
        RECT 2705.725 1797.935 2706.935 1798.455 ;
        RECT 2699.275 1797.165 2699.605 1797.625 ;
        RECT 2700.205 1797.165 2705.550 1797.710 ;
        RECT 2705.725 1797.165 2708.315 1797.935 ;
        RECT 2708.485 1797.165 2708.775 1797.890 ;
        RECT 2710.530 1797.710 2710.870 1798.540 ;
        RECT 2716.050 1797.710 2716.390 1798.540 ;
        RECT 2721.570 1797.710 2721.910 1798.540 ;
        RECT 2727.090 1797.710 2727.430 1798.540 ;
        RECT 2731.025 1797.935 2731.775 1798.455 ;
        RECT 2708.945 1797.165 2714.290 1797.710 ;
        RECT 2714.465 1797.165 2719.810 1797.710 ;
        RECT 2719.985 1797.165 2725.330 1797.710 ;
        RECT 2725.505 1797.165 2730.850 1797.710 ;
        RECT 2731.025 1797.165 2732.695 1797.935 ;
        RECT 2733.555 1797.915 2734.075 1798.455 ;
        RECT 2732.865 1797.165 2734.075 1797.915 ;
        RECT 2695.520 1796.995 2734.160 1797.165 ;
        RECT 2695.605 1796.245 2696.815 1796.995 ;
        RECT 2697.425 1796.615 2697.755 1796.995 ;
        RECT 2698.365 1796.450 2703.710 1796.995 ;
        RECT 2703.885 1796.450 2709.230 1796.995 ;
        RECT 2709.405 1796.450 2714.750 1796.995 ;
        RECT 2714.925 1796.450 2720.270 1796.995 ;
        RECT 2695.605 1795.705 2696.125 1796.245 ;
        RECT 2699.950 1795.620 2700.290 1796.450 ;
        RECT 2705.470 1795.620 2705.810 1796.450 ;
        RECT 2710.990 1795.620 2711.330 1796.450 ;
        RECT 2716.510 1795.620 2716.850 1796.450 ;
        RECT 2721.365 1796.270 2721.655 1796.995 ;
        RECT 2721.825 1796.450 2727.170 1796.995 ;
        RECT 2727.345 1796.450 2732.690 1796.995 ;
        RECT 2723.410 1795.620 2723.750 1796.450 ;
        RECT 2728.930 1795.620 2729.270 1796.450 ;
        RECT 2732.865 1796.245 2734.075 1796.995 ;
        RECT 2733.555 1795.705 2734.075 1796.245 ;
        RECT 2695.605 1792.475 2696.125 1793.015 ;
        RECT 2696.985 1792.475 2697.505 1793.015 ;
        RECT 2343.000 1790.865 2447.045 1792.465 ;
        RECT 2523.330 1791.305 2523.670 1791.965 ;
        RECT 2695.605 1791.725 2696.815 1792.475 ;
        RECT 2696.985 1791.725 2698.195 1792.475 ;
        RECT 2698.365 1791.725 2698.705 1792.450 ;
        RECT 2703.630 1792.270 2703.970 1793.100 ;
        RECT 2701.035 1791.725 2701.365 1792.205 ;
        RECT 2702.045 1791.725 2707.390 1792.270 ;
        RECT 2708.485 1791.725 2708.775 1792.450 ;
        RECT 2710.530 1792.270 2710.870 1793.100 ;
        RECT 2716.050 1792.270 2716.390 1793.100 ;
        RECT 2721.570 1792.270 2721.910 1793.100 ;
        RECT 2727.090 1792.270 2727.430 1793.100 ;
        RECT 2731.025 1792.495 2731.775 1793.015 ;
        RECT 2708.945 1791.725 2714.290 1792.270 ;
        RECT 2714.465 1791.725 2719.810 1792.270 ;
        RECT 2719.985 1791.725 2725.330 1792.270 ;
        RECT 2725.505 1791.725 2730.850 1792.270 ;
        RECT 2731.025 1791.725 2732.695 1792.495 ;
        RECT 2733.555 1792.475 2734.075 1793.015 ;
        RECT 2732.865 1791.725 2734.075 1792.475 ;
        RECT 2695.520 1791.555 2734.160 1791.725 ;
        RECT 2522.130 1791.135 2523.935 1791.305 ;
        RECT 2368.165 1790.240 2368.335 1790.865 ;
        RECT 2375.680 1790.240 2375.850 1790.865 ;
        RECT 2376.635 1790.320 2376.805 1790.600 ;
        RECT 2376.635 1790.150 2376.865 1790.320 ;
        RECT 2381.295 1790.240 2381.465 1790.865 ;
        RECT 2384.040 1790.240 2384.210 1790.865 ;
        RECT 2385.030 1790.240 2385.200 1790.865 ;
        RECT 2390.940 1790.240 2391.110 1790.865 ;
        RECT 2391.895 1790.320 2392.065 1790.600 ;
        RECT 2391.895 1790.150 2392.125 1790.320 ;
        RECT 2396.555 1790.240 2396.725 1790.865 ;
        RECT 2399.300 1790.240 2399.470 1790.865 ;
        RECT 2400.290 1790.240 2400.460 1790.865 ;
        RECT 2406.200 1790.240 2406.370 1790.865 ;
        RECT 2407.155 1790.320 2407.325 1790.600 ;
        RECT 2407.155 1790.150 2407.385 1790.320 ;
        RECT 2411.815 1790.240 2411.985 1790.865 ;
        RECT 2414.560 1790.240 2414.730 1790.865 ;
        RECT 2415.550 1790.240 2415.720 1790.865 ;
        RECT 2421.460 1790.240 2421.630 1790.865 ;
        RECT 2422.415 1790.320 2422.585 1790.600 ;
        RECT 2422.415 1790.150 2422.645 1790.320 ;
        RECT 2427.075 1790.240 2427.245 1790.865 ;
        RECT 2429.820 1790.240 2429.990 1790.865 ;
        RECT 2430.810 1790.240 2430.980 1790.865 ;
        RECT 2436.720 1790.240 2436.890 1790.865 ;
        RECT 2437.675 1790.320 2437.845 1790.600 ;
        RECT 2437.675 1790.150 2437.905 1790.320 ;
        RECT 2442.335 1790.240 2442.505 1790.865 ;
        RECT 2445.080 1790.240 2445.250 1790.865 ;
        RECT 2446.070 1790.240 2446.240 1790.865 ;
        RECT 2695.605 1790.805 2696.815 1791.555 ;
        RECT 2695.605 1790.265 2696.125 1790.805 ;
        RECT 2697.905 1790.735 2698.165 1791.555 ;
        RECT 2699.275 1791.155 2699.605 1791.555 ;
        RECT 2700.115 1791.155 2700.490 1791.555 ;
        RECT 2702.760 1791.155 2703.090 1791.555 ;
        RECT 2703.885 1791.010 2709.230 1791.555 ;
        RECT 2709.405 1791.010 2714.750 1791.555 ;
        RECT 2714.925 1791.010 2720.270 1791.555 ;
        RECT 2705.470 1790.180 2705.810 1791.010 ;
        RECT 2710.990 1790.180 2711.330 1791.010 ;
        RECT 2716.510 1790.180 2716.850 1791.010 ;
        RECT 2721.365 1790.830 2721.655 1791.555 ;
        RECT 2721.825 1791.010 2727.170 1791.555 ;
        RECT 2727.345 1791.010 2732.690 1791.555 ;
        RECT 2723.410 1790.180 2723.750 1791.010 ;
        RECT 2728.930 1790.180 2729.270 1791.010 ;
        RECT 2732.865 1790.805 2734.075 1791.555 ;
        RECT 2733.555 1790.265 2734.075 1790.805 ;
        RECT 2376.695 1788.540 2376.865 1790.150 ;
        RECT 2391.955 1788.540 2392.125 1790.150 ;
        RECT 2407.215 1788.540 2407.385 1790.150 ;
        RECT 2422.475 1788.540 2422.645 1790.150 ;
        RECT 2437.735 1788.540 2437.905 1790.150 ;
        RECT 2376.635 1788.370 2376.865 1788.540 ;
        RECT 2391.895 1788.370 2392.125 1788.540 ;
        RECT 2407.155 1788.370 2407.385 1788.540 ;
        RECT 2422.415 1788.370 2422.645 1788.540 ;
        RECT 2437.675 1788.370 2437.905 1788.540 ;
        RECT 2376.635 1787.310 2376.805 1788.370 ;
        RECT 2391.895 1787.310 2392.065 1788.370 ;
        RECT 2407.155 1787.310 2407.325 1788.370 ;
        RECT 2422.415 1787.310 2422.585 1788.370 ;
        RECT 2437.675 1787.310 2437.845 1788.370 ;
        RECT 2695.605 1787.035 2696.125 1787.575 ;
        RECT 2695.605 1786.285 2696.815 1787.035 ;
        RECT 2697.425 1786.285 2697.755 1786.665 ;
        RECT 2699.725 1786.285 2700.035 1787.085 ;
        RECT 2701.790 1786.830 2702.130 1787.660 ;
        RECT 2705.725 1787.055 2706.935 1787.575 ;
        RECT 2700.205 1786.285 2705.550 1786.830 ;
        RECT 2705.725 1786.285 2708.315 1787.055 ;
        RECT 2708.485 1786.285 2708.775 1787.010 ;
        RECT 2710.530 1786.830 2710.870 1787.660 ;
        RECT 2716.050 1786.830 2716.390 1787.660 ;
        RECT 2721.570 1786.830 2721.910 1787.660 ;
        RECT 2727.090 1786.830 2727.430 1787.660 ;
        RECT 2731.025 1787.055 2731.775 1787.575 ;
        RECT 2708.945 1786.285 2714.290 1786.830 ;
        RECT 2714.465 1786.285 2719.810 1786.830 ;
        RECT 2719.985 1786.285 2725.330 1786.830 ;
        RECT 2725.505 1786.285 2730.850 1786.830 ;
        RECT 2731.025 1786.285 2732.695 1787.055 ;
        RECT 2733.555 1787.035 2734.075 1787.575 ;
        RECT 2732.865 1786.285 2734.075 1787.035 ;
        RECT 2695.520 1786.115 2734.160 1786.285 ;
        RECT 2523.330 1785.360 2523.670 1786.020 ;
        RECT 2695.605 1785.365 2696.815 1786.115 ;
        RECT 2697.725 1785.580 2698.235 1786.115 ;
        RECT 2700.195 1785.715 2700.525 1786.115 ;
        RECT 2701.125 1785.570 2706.470 1786.115 ;
        RECT 2706.645 1785.570 2711.990 1786.115 ;
        RECT 2712.165 1785.570 2717.510 1786.115 ;
        RECT 2522.130 1785.190 2523.935 1785.360 ;
        RECT 2695.605 1784.825 2696.125 1785.365 ;
        RECT 2702.710 1784.740 2703.050 1785.570 ;
        RECT 2708.230 1784.740 2708.570 1785.570 ;
        RECT 2713.750 1784.740 2714.090 1785.570 ;
        RECT 2717.685 1785.345 2721.195 1786.115 ;
        RECT 2721.365 1785.390 2721.655 1786.115 ;
        RECT 2721.825 1785.570 2727.170 1786.115 ;
        RECT 2727.345 1785.570 2732.690 1786.115 ;
        RECT 2717.685 1784.825 2719.335 1785.345 ;
        RECT 2723.410 1784.740 2723.750 1785.570 ;
        RECT 2728.930 1784.740 2729.270 1785.570 ;
        RECT 2732.865 1785.365 2734.075 1786.115 ;
        RECT 2733.555 1784.825 2734.075 1785.365 ;
        RECT 2372.045 1783.785 2372.215 1784.235 ;
        RECT 2373.365 1783.865 2373.735 1784.035 ;
        RECT 2373.365 1783.395 2373.535 1783.865 ;
        RECT 2387.305 1783.785 2387.475 1784.235 ;
        RECT 2388.625 1783.865 2388.995 1784.035 ;
        RECT 2388.625 1783.395 2388.795 1783.865 ;
        RECT 2402.565 1783.785 2402.735 1784.235 ;
        RECT 2403.885 1783.865 2404.255 1784.035 ;
        RECT 2403.885 1783.395 2404.055 1783.865 ;
        RECT 2417.825 1783.785 2417.995 1784.235 ;
        RECT 2419.145 1783.865 2419.515 1784.035 ;
        RECT 2419.145 1783.395 2419.315 1783.865 ;
        RECT 2433.085 1783.785 2433.255 1784.235 ;
        RECT 2434.405 1783.865 2434.775 1784.035 ;
        RECT 2434.405 1783.395 2434.575 1783.865 ;
        RECT 2372.765 1782.890 2372.935 1783.375 ;
        RECT 2373.245 1783.225 2373.535 1783.395 ;
        RECT 2372.765 1782.875 2373.040 1782.890 ;
        RECT 2374.685 1782.875 2374.855 1783.375 ;
        RECT 2375.645 1782.875 2375.815 1783.375 ;
        RECT 2376.520 1782.875 2376.715 1782.890 ;
        RECT 2377.565 1782.875 2377.735 1783.375 ;
        RECT 2378.525 1782.880 2378.695 1783.375 ;
        RECT 2378.370 1782.875 2378.695 1782.880 ;
        RECT 2379.465 1782.875 2379.635 1783.375 ;
        RECT 2388.025 1782.890 2388.195 1783.375 ;
        RECT 2388.505 1783.225 2388.795 1783.395 ;
        RECT 2380.040 1782.875 2380.235 1782.880 ;
        RECT 2388.025 1782.875 2388.300 1782.890 ;
        RECT 2389.945 1782.875 2390.115 1783.375 ;
        RECT 2390.905 1782.875 2391.075 1783.375 ;
        RECT 2391.780 1782.875 2391.975 1782.890 ;
        RECT 2392.825 1782.875 2392.995 1783.375 ;
        RECT 2393.785 1782.880 2393.955 1783.375 ;
        RECT 2393.630 1782.875 2393.955 1782.880 ;
        RECT 2394.725 1782.875 2394.895 1783.375 ;
        RECT 2403.285 1782.890 2403.455 1783.375 ;
        RECT 2403.765 1783.225 2404.055 1783.395 ;
        RECT 2395.300 1782.875 2395.495 1782.880 ;
        RECT 2403.285 1782.875 2403.560 1782.890 ;
        RECT 2405.205 1782.875 2405.375 1783.375 ;
        RECT 2406.165 1782.875 2406.335 1783.375 ;
        RECT 2407.040 1782.875 2407.235 1782.890 ;
        RECT 2408.085 1782.875 2408.255 1783.375 ;
        RECT 2409.045 1782.880 2409.215 1783.375 ;
        RECT 2408.890 1782.875 2409.215 1782.880 ;
        RECT 2409.985 1782.875 2410.155 1783.375 ;
        RECT 2418.545 1782.890 2418.715 1783.375 ;
        RECT 2419.025 1783.225 2419.315 1783.395 ;
        RECT 2410.560 1782.875 2410.755 1782.880 ;
        RECT 2418.545 1782.875 2418.820 1782.890 ;
        RECT 2420.465 1782.875 2420.635 1783.375 ;
        RECT 2421.425 1782.875 2421.595 1783.375 ;
        RECT 2422.300 1782.875 2422.495 1782.890 ;
        RECT 2423.345 1782.875 2423.515 1783.375 ;
        RECT 2424.305 1782.880 2424.475 1783.375 ;
        RECT 2424.150 1782.875 2424.475 1782.880 ;
        RECT 2425.245 1782.875 2425.415 1783.375 ;
        RECT 2433.805 1782.890 2433.975 1783.375 ;
        RECT 2434.285 1783.225 2434.575 1783.395 ;
        RECT 2425.820 1782.875 2426.015 1782.880 ;
        RECT 2433.805 1782.875 2434.080 1782.890 ;
        RECT 2435.725 1782.875 2435.895 1783.375 ;
        RECT 2436.685 1782.875 2436.855 1783.375 ;
        RECT 2437.560 1782.875 2437.755 1782.890 ;
        RECT 2438.605 1782.875 2438.775 1783.375 ;
        RECT 2439.565 1782.880 2439.735 1783.375 ;
        RECT 2439.410 1782.875 2439.735 1782.880 ;
        RECT 2440.505 1782.875 2440.675 1783.375 ;
        RECT 2441.080 1782.875 2441.275 1782.880 ;
        RECT 2371.495 1781.600 2380.235 1782.875 ;
        RECT 2381.295 1781.600 2381.465 1782.225 ;
        RECT 2384.040 1781.600 2384.210 1782.225 ;
        RECT 2385.025 1781.600 2385.195 1782.225 ;
        RECT 2386.755 1781.600 2395.495 1782.875 ;
        RECT 2396.555 1781.600 2396.725 1782.225 ;
        RECT 2399.300 1781.600 2399.470 1782.225 ;
        RECT 2400.285 1781.600 2400.455 1782.225 ;
        RECT 2402.015 1781.600 2410.755 1782.875 ;
        RECT 2411.815 1781.600 2411.985 1782.225 ;
        RECT 2414.560 1781.600 2414.730 1782.225 ;
        RECT 2415.545 1781.600 2415.715 1782.225 ;
        RECT 2417.275 1781.600 2426.015 1782.875 ;
        RECT 2427.075 1781.600 2427.245 1782.225 ;
        RECT 2429.820 1781.600 2429.990 1782.225 ;
        RECT 2430.805 1781.600 2430.975 1782.225 ;
        RECT 2432.535 1781.600 2441.275 1782.875 ;
        RECT 2442.335 1781.600 2442.505 1782.225 ;
        RECT 2445.080 1781.600 2445.250 1782.225 ;
        RECT 2446.065 1781.600 2446.235 1782.225 ;
        RECT 2343.000 1780.000 2447.045 1781.600 ;
        RECT 2695.605 1781.595 2696.125 1782.135 ;
        RECT 2695.605 1780.845 2696.815 1781.595 ;
        RECT 2699.950 1781.390 2700.290 1782.220 ;
        RECT 2703.885 1781.615 2705.535 1782.135 ;
        RECT 2697.425 1780.845 2697.755 1781.225 ;
        RECT 2698.365 1780.845 2703.710 1781.390 ;
        RECT 2703.885 1780.845 2707.395 1781.615 ;
        RECT 2708.485 1780.845 2708.775 1781.570 ;
        RECT 2710.530 1781.390 2710.870 1782.220 ;
        RECT 2716.050 1781.390 2716.390 1782.220 ;
        RECT 2721.570 1781.390 2721.910 1782.220 ;
        RECT 2727.090 1781.390 2727.430 1782.220 ;
        RECT 2731.025 1781.615 2731.775 1782.135 ;
        RECT 2708.945 1780.845 2714.290 1781.390 ;
        RECT 2714.465 1780.845 2719.810 1781.390 ;
        RECT 2719.985 1780.845 2725.330 1781.390 ;
        RECT 2725.505 1780.845 2730.850 1781.390 ;
        RECT 2731.025 1780.845 2732.695 1781.615 ;
        RECT 2733.555 1781.595 2734.075 1782.135 ;
        RECT 2732.865 1780.845 2734.075 1781.595 ;
        RECT 2695.520 1780.675 2734.160 1780.845 ;
        RECT 2523.330 1779.715 2523.670 1780.375 ;
        RECT 2695.605 1779.925 2696.815 1780.675 ;
        RECT 2696.985 1780.130 2702.330 1780.675 ;
        RECT 2702.505 1780.130 2707.850 1780.675 ;
        RECT 2708.025 1780.130 2713.370 1780.675 ;
        RECT 2713.545 1780.130 2718.890 1780.675 ;
        RECT 2522.130 1779.545 2523.935 1779.715 ;
        RECT 2695.605 1779.385 2696.125 1779.925 ;
        RECT 2698.570 1779.300 2698.910 1780.130 ;
        RECT 2704.090 1779.300 2704.430 1780.130 ;
        RECT 2709.610 1779.300 2709.950 1780.130 ;
        RECT 2715.130 1779.300 2715.470 1780.130 ;
        RECT 2719.065 1779.905 2720.735 1780.675 ;
        RECT 2721.365 1779.950 2721.655 1780.675 ;
        RECT 2721.825 1780.130 2727.170 1780.675 ;
        RECT 2727.345 1780.130 2732.690 1780.675 ;
        RECT 2719.065 1779.385 2719.815 1779.905 ;
        RECT 2723.410 1779.300 2723.750 1780.130 ;
        RECT 2728.930 1779.300 2729.270 1780.130 ;
        RECT 2732.865 1779.925 2734.075 1780.675 ;
        RECT 2733.555 1779.385 2734.075 1779.925 ;
        RECT 2695.605 1776.155 2696.125 1776.695 ;
        RECT 2695.605 1775.405 2696.815 1776.155 ;
        RECT 2699.950 1775.950 2700.290 1776.780 ;
        RECT 2703.885 1776.175 2705.535 1776.695 ;
        RECT 2697.425 1775.405 2697.755 1775.785 ;
        RECT 2698.365 1775.405 2703.710 1775.950 ;
        RECT 2703.885 1775.405 2707.395 1776.175 ;
        RECT 2708.485 1775.405 2708.775 1776.130 ;
        RECT 2710.530 1775.950 2710.870 1776.780 ;
        RECT 2716.050 1775.950 2716.390 1776.780 ;
        RECT 2721.570 1775.950 2721.910 1776.780 ;
        RECT 2727.090 1775.950 2727.430 1776.780 ;
        RECT 2731.025 1776.175 2731.775 1776.695 ;
        RECT 2708.945 1775.405 2714.290 1775.950 ;
        RECT 2714.465 1775.405 2719.810 1775.950 ;
        RECT 2719.985 1775.405 2725.330 1775.950 ;
        RECT 2725.505 1775.405 2730.850 1775.950 ;
        RECT 2731.025 1775.405 2732.695 1776.175 ;
        RECT 2733.555 1776.155 2734.075 1776.695 ;
        RECT 2732.865 1775.405 2734.075 1776.155 ;
        RECT 2695.520 1775.235 2734.160 1775.405 ;
        RECT 2695.605 1774.485 2696.815 1775.235 ;
        RECT 2696.985 1774.690 2702.330 1775.235 ;
        RECT 2702.505 1774.690 2707.850 1775.235 ;
        RECT 2708.025 1774.690 2713.370 1775.235 ;
        RECT 2713.545 1774.690 2718.890 1775.235 ;
        RECT 2695.605 1773.945 2696.125 1774.485 ;
        RECT 2698.570 1773.860 2698.910 1774.690 ;
        RECT 2704.090 1773.860 2704.430 1774.690 ;
        RECT 2709.610 1773.860 2709.950 1774.690 ;
        RECT 2715.130 1773.860 2715.470 1774.690 ;
        RECT 2719.065 1774.465 2720.735 1775.235 ;
        RECT 2721.365 1774.510 2721.655 1775.235 ;
        RECT 2721.825 1774.690 2727.170 1775.235 ;
        RECT 2727.345 1774.690 2732.690 1775.235 ;
        RECT 2719.065 1773.945 2719.815 1774.465 ;
        RECT 2723.410 1773.860 2723.750 1774.690 ;
        RECT 2728.930 1773.860 2729.270 1774.690 ;
        RECT 2732.865 1774.485 2734.075 1775.235 ;
        RECT 2733.555 1773.945 2734.075 1774.485 ;
        RECT 2695.605 1770.715 2696.125 1771.255 ;
        RECT 2695.605 1769.965 2696.815 1770.715 ;
        RECT 2701.330 1770.510 2701.670 1771.340 ;
        RECT 2705.265 1770.735 2706.475 1771.255 ;
        RECT 2697.425 1769.965 2697.755 1770.345 ;
        RECT 2698.805 1769.965 2699.135 1770.345 ;
        RECT 2699.745 1769.965 2705.090 1770.510 ;
        RECT 2705.265 1769.965 2707.855 1770.735 ;
        RECT 2708.485 1769.965 2708.775 1770.690 ;
        RECT 2710.530 1770.510 2710.870 1771.340 ;
        RECT 2716.050 1770.510 2716.390 1771.340 ;
        RECT 2719.985 1770.715 2720.505 1771.255 ;
        RECT 2708.945 1769.965 2714.290 1770.510 ;
        RECT 2714.465 1769.965 2719.810 1770.510 ;
        RECT 2719.985 1769.965 2721.195 1770.715 ;
        RECT 2721.365 1769.965 2721.655 1770.690 ;
        RECT 2723.410 1770.510 2723.750 1771.340 ;
        RECT 2728.930 1770.510 2729.270 1771.340 ;
        RECT 2733.555 1770.715 2734.075 1771.255 ;
        RECT 2721.825 1769.965 2727.170 1770.510 ;
        RECT 2727.345 1769.965 2732.690 1770.510 ;
        RECT 2732.865 1769.965 2734.075 1770.715 ;
        RECT 2695.520 1769.795 2734.160 1769.965 ;
        RECT 2523.330 1768.245 2523.670 1768.905 ;
        RECT 2522.130 1768.075 2523.935 1768.245 ;
        RECT 2410.920 1712.465 2444.085 1712.470 ;
        RECT 2394.335 1712.460 2444.085 1712.465 ;
        RECT 2343.000 1710.860 2444.085 1712.460 ;
        RECT 2358.415 1710.855 2361.165 1710.860 ;
        RECT 2361.645 1710.855 2365.170 1710.860 ;
        RECT 2358.585 1710.225 2358.755 1710.855 ;
        RECT 2361.815 1710.225 2361.985 1710.855 ;
        RECT 2362.770 1710.305 2362.940 1710.585 ;
        RECT 2362.770 1710.135 2363.000 1710.305 ;
        RECT 2362.830 1708.525 2363.000 1710.135 ;
        RECT 2364.880 1708.525 2365.170 1710.855 ;
        RECT 2365.450 1708.525 2365.730 1710.860 ;
        RECT 2366.010 1708.525 2366.290 1710.860 ;
        RECT 2366.570 1708.525 2366.850 1710.860 ;
        RECT 2367.130 1708.525 2367.410 1710.860 ;
        RECT 2367.690 1708.525 2367.970 1710.860 ;
        RECT 2368.250 1708.525 2368.530 1710.860 ;
        RECT 2368.810 1708.525 2369.090 1710.860 ;
        RECT 2369.370 1708.525 2369.650 1710.860 ;
        RECT 2369.930 1708.525 2370.210 1710.860 ;
        RECT 2370.490 1708.525 2370.770 1710.860 ;
        RECT 2371.050 1708.525 2371.330 1710.860 ;
        RECT 2371.610 1708.525 2371.785 1710.860 ;
        RECT 2373.040 1710.230 2373.210 1710.860 ;
        RECT 2375.785 1710.230 2375.955 1710.860 ;
        RECT 2376.775 1710.230 2376.945 1710.860 ;
        RECT 2378.230 1710.855 2381.755 1710.860 ;
        RECT 2378.400 1710.225 2378.570 1710.855 ;
        RECT 2379.355 1710.305 2379.525 1710.585 ;
        RECT 2379.355 1710.135 2379.585 1710.305 ;
        RECT 2379.415 1708.525 2379.585 1710.135 ;
        RECT 2381.465 1708.525 2381.755 1710.855 ;
        RECT 2382.035 1708.525 2382.315 1710.860 ;
        RECT 2382.595 1708.525 2382.875 1710.860 ;
        RECT 2383.155 1708.525 2383.435 1710.860 ;
        RECT 2383.715 1708.525 2383.995 1710.860 ;
        RECT 2384.275 1708.525 2384.555 1710.860 ;
        RECT 2384.835 1708.525 2385.115 1710.860 ;
        RECT 2385.395 1708.525 2385.675 1710.860 ;
        RECT 2385.955 1708.525 2386.235 1710.860 ;
        RECT 2386.515 1708.525 2386.795 1710.860 ;
        RECT 2387.075 1708.525 2387.355 1710.860 ;
        RECT 2387.635 1708.525 2387.915 1710.860 ;
        RECT 2388.195 1708.525 2388.370 1710.860 ;
        RECT 2389.625 1710.230 2389.795 1710.860 ;
        RECT 2392.370 1710.230 2392.540 1710.860 ;
        RECT 2393.360 1710.230 2393.530 1710.860 ;
        RECT 2394.985 1710.230 2395.155 1710.860 ;
        RECT 2395.940 1710.310 2396.110 1710.590 ;
        RECT 2395.940 1710.140 2396.170 1710.310 ;
        RECT 2396.000 1708.530 2396.170 1710.140 ;
        RECT 2398.050 1708.530 2398.340 1710.860 ;
        RECT 2398.620 1708.530 2398.900 1710.860 ;
        RECT 2399.180 1708.530 2399.460 1710.860 ;
        RECT 2399.740 1708.530 2400.020 1710.860 ;
        RECT 2400.300 1708.530 2400.580 1710.860 ;
        RECT 2400.860 1708.530 2401.140 1710.860 ;
        RECT 2401.420 1708.530 2401.700 1710.860 ;
        RECT 2401.980 1708.530 2402.260 1710.860 ;
        RECT 2402.540 1708.530 2402.820 1710.860 ;
        RECT 2403.100 1708.530 2403.380 1710.860 ;
        RECT 2403.660 1708.530 2403.940 1710.860 ;
        RECT 2404.220 1708.530 2404.500 1710.860 ;
        RECT 2404.780 1708.530 2404.955 1710.860 ;
        RECT 2406.210 1710.235 2406.380 1710.860 ;
        RECT 2408.955 1710.235 2409.125 1710.860 ;
        RECT 2409.945 1710.235 2410.115 1710.860 ;
        RECT 2411.570 1710.235 2411.740 1710.860 ;
        RECT 2412.525 1710.315 2412.695 1710.595 ;
        RECT 2412.525 1710.145 2412.755 1710.315 ;
        RECT 2412.585 1708.535 2412.755 1710.145 ;
        RECT 2414.635 1708.535 2414.925 1710.860 ;
        RECT 2415.205 1708.535 2415.485 1710.860 ;
        RECT 2415.765 1708.535 2416.045 1710.860 ;
        RECT 2416.325 1708.535 2416.605 1710.860 ;
        RECT 2416.885 1708.535 2417.165 1710.860 ;
        RECT 2417.445 1708.535 2417.725 1710.860 ;
        RECT 2418.005 1708.535 2418.285 1710.860 ;
        RECT 2418.565 1708.535 2418.845 1710.860 ;
        RECT 2419.125 1708.535 2419.405 1710.860 ;
        RECT 2419.685 1708.535 2419.965 1710.860 ;
        RECT 2420.245 1708.535 2420.525 1710.860 ;
        RECT 2420.805 1708.535 2421.085 1710.860 ;
        RECT 2421.365 1708.535 2421.540 1710.860 ;
        RECT 2422.795 1710.240 2422.965 1710.860 ;
        RECT 2425.540 1710.240 2425.710 1710.860 ;
        RECT 2426.530 1710.240 2426.700 1710.860 ;
        RECT 2428.150 1710.235 2428.320 1710.860 ;
        RECT 2429.105 1710.315 2429.275 1710.595 ;
        RECT 2429.105 1710.145 2429.335 1710.315 ;
        RECT 2429.165 1708.535 2429.335 1710.145 ;
        RECT 2431.215 1708.535 2431.505 1710.860 ;
        RECT 2431.785 1708.535 2432.065 1710.860 ;
        RECT 2432.345 1708.535 2432.625 1710.860 ;
        RECT 2432.905 1708.535 2433.185 1710.860 ;
        RECT 2433.465 1708.535 2433.745 1710.860 ;
        RECT 2434.025 1708.535 2434.305 1710.860 ;
        RECT 2434.585 1708.535 2434.865 1710.860 ;
        RECT 2435.145 1708.535 2435.425 1710.860 ;
        RECT 2435.705 1708.535 2435.985 1710.860 ;
        RECT 2436.265 1708.535 2436.545 1710.860 ;
        RECT 2436.825 1708.535 2437.105 1710.860 ;
        RECT 2437.385 1708.535 2437.665 1710.860 ;
        RECT 2437.945 1708.535 2438.120 1710.860 ;
        RECT 2439.375 1710.240 2439.545 1710.860 ;
        RECT 2442.120 1710.240 2442.290 1710.860 ;
        RECT 2443.110 1710.240 2443.280 1710.860 ;
        RECT 2362.770 1708.355 2363.000 1708.525 ;
        RECT 2364.740 1708.355 2371.785 1708.525 ;
        RECT 2379.355 1708.355 2379.585 1708.525 ;
        RECT 2381.325 1708.355 2388.370 1708.525 ;
        RECT 2395.940 1708.360 2396.170 1708.530 ;
        RECT 2397.910 1708.360 2404.955 1708.530 ;
        RECT 2412.525 1708.365 2412.755 1708.535 ;
        RECT 2414.495 1708.365 2421.540 1708.535 ;
        RECT 2429.105 1708.365 2429.335 1708.535 ;
        RECT 2431.075 1708.365 2438.120 1708.535 ;
        RECT 2362.770 1707.295 2362.940 1708.355 ;
        RECT 2366.150 1707.895 2366.400 1708.355 ;
        RECT 2368.220 1707.955 2368.550 1708.355 ;
        RECT 2370.310 1707.845 2370.760 1708.355 ;
        RECT 2366.300 1707.115 2366.640 1707.365 ;
        RECT 2368.520 1707.115 2368.850 1707.445 ;
        RECT 2379.355 1707.295 2379.525 1708.355 ;
        RECT 2382.735 1707.895 2382.985 1708.355 ;
        RECT 2384.805 1707.955 2385.135 1708.355 ;
        RECT 2386.895 1707.845 2387.345 1708.355 ;
        RECT 2382.885 1707.115 2383.225 1707.365 ;
        RECT 2385.105 1707.115 2385.435 1707.445 ;
        RECT 2395.940 1707.300 2396.110 1708.360 ;
        RECT 2399.320 1707.900 2399.570 1708.360 ;
        RECT 2401.390 1707.960 2401.720 1708.360 ;
        RECT 2403.480 1707.850 2403.930 1708.360 ;
        RECT 2399.470 1707.120 2399.810 1707.370 ;
        RECT 2401.690 1707.120 2402.020 1707.450 ;
        RECT 2412.525 1707.305 2412.695 1708.365 ;
        RECT 2415.905 1707.905 2416.155 1708.365 ;
        RECT 2417.975 1707.965 2418.305 1708.365 ;
        RECT 2420.065 1707.855 2420.515 1708.365 ;
        RECT 2416.055 1707.125 2416.395 1707.375 ;
        RECT 2418.275 1707.125 2418.605 1707.455 ;
        RECT 2429.105 1707.305 2429.275 1708.365 ;
        RECT 2432.485 1707.905 2432.735 1708.365 ;
        RECT 2434.555 1707.965 2434.885 1708.365 ;
        RECT 2436.645 1707.855 2437.095 1708.365 ;
        RECT 2432.635 1707.125 2432.975 1707.375 ;
        RECT 2434.855 1707.125 2435.185 1707.455 ;
        RECT 2364.660 1703.355 2364.915 1703.905 ;
        RECT 2364.660 1703.095 2364.920 1703.355 ;
        RECT 2367.250 1703.095 2367.580 1703.545 ;
        RECT 2369.630 1703.095 2369.880 1703.625 ;
        RECT 2370.500 1703.095 2370.740 1703.895 ;
        RECT 2371.410 1703.095 2371.680 1703.895 ;
        RECT 2381.245 1703.355 2381.500 1703.905 ;
        RECT 2381.245 1703.095 2381.505 1703.355 ;
        RECT 2383.835 1703.095 2384.165 1703.545 ;
        RECT 2386.215 1703.095 2386.465 1703.625 ;
        RECT 2387.085 1703.095 2387.325 1703.895 ;
        RECT 2387.995 1703.095 2388.265 1703.895 ;
        RECT 2397.830 1703.360 2398.085 1703.910 ;
        RECT 2397.830 1703.100 2398.090 1703.360 ;
        RECT 2400.420 1703.100 2400.750 1703.550 ;
        RECT 2402.800 1703.100 2403.050 1703.630 ;
        RECT 2403.670 1703.100 2403.910 1703.900 ;
        RECT 2404.580 1703.100 2404.850 1703.900 ;
        RECT 2414.415 1703.365 2414.670 1703.915 ;
        RECT 2414.415 1703.105 2414.675 1703.365 ;
        RECT 2417.005 1703.105 2417.335 1703.555 ;
        RECT 2419.385 1703.105 2419.635 1703.635 ;
        RECT 2420.255 1703.105 2420.495 1703.905 ;
        RECT 2421.165 1703.105 2421.435 1703.905 ;
        RECT 2430.995 1703.365 2431.250 1703.915 ;
        RECT 2430.995 1703.105 2431.255 1703.365 ;
        RECT 2433.585 1703.105 2433.915 1703.555 ;
        RECT 2435.965 1703.105 2436.215 1703.635 ;
        RECT 2436.835 1703.105 2437.075 1703.905 ;
        RECT 2437.745 1703.105 2438.015 1703.905 ;
        RECT 2364.580 1702.925 2371.970 1703.095 ;
        RECT 2381.165 1702.925 2388.555 1703.095 ;
        RECT 2397.750 1702.930 2405.140 1703.100 ;
        RECT 2414.335 1702.935 2421.725 1703.105 ;
        RECT 2430.915 1702.935 2438.305 1703.105 ;
        RECT 2364.625 1701.605 2364.920 1702.925 ;
        RECT 2365.210 1701.605 2365.500 1702.925 ;
        RECT 2365.790 1701.605 2366.080 1702.925 ;
        RECT 2366.370 1701.605 2366.660 1702.925 ;
        RECT 2366.950 1701.605 2367.240 1702.925 ;
        RECT 2367.530 1701.605 2367.815 1702.925 ;
        RECT 2368.105 1701.605 2368.395 1702.925 ;
        RECT 2368.685 1701.605 2368.975 1702.925 ;
        RECT 2369.265 1701.605 2369.555 1702.925 ;
        RECT 2369.845 1701.605 2370.130 1702.925 ;
        RECT 2370.420 1701.605 2370.710 1702.925 ;
        RECT 2371.000 1701.605 2371.290 1702.925 ;
        RECT 2371.580 1701.605 2371.970 1702.925 ;
        RECT 2364.625 1701.600 2371.970 1701.605 ;
        RECT 2373.040 1701.600 2373.210 1702.230 ;
        RECT 2375.785 1701.600 2375.955 1702.230 ;
        RECT 2376.775 1701.600 2376.945 1702.230 ;
        RECT 2381.210 1701.605 2381.505 1702.925 ;
        RECT 2381.795 1701.605 2382.085 1702.925 ;
        RECT 2382.375 1701.605 2382.665 1702.925 ;
        RECT 2382.955 1701.605 2383.245 1702.925 ;
        RECT 2383.535 1701.605 2383.825 1702.925 ;
        RECT 2384.115 1701.605 2384.400 1702.925 ;
        RECT 2384.690 1701.605 2384.980 1702.925 ;
        RECT 2385.270 1701.605 2385.560 1702.925 ;
        RECT 2385.850 1701.605 2386.140 1702.925 ;
        RECT 2386.430 1701.605 2386.715 1702.925 ;
        RECT 2387.005 1701.605 2387.295 1702.925 ;
        RECT 2387.585 1701.605 2387.875 1702.925 ;
        RECT 2388.165 1701.605 2388.555 1702.925 ;
        RECT 2381.210 1701.600 2388.555 1701.605 ;
        RECT 2389.625 1701.600 2389.795 1702.230 ;
        RECT 2392.370 1701.600 2392.540 1702.230 ;
        RECT 2393.360 1701.600 2393.530 1702.230 ;
        RECT 2397.795 1701.610 2398.090 1702.930 ;
        RECT 2398.380 1701.610 2398.670 1702.930 ;
        RECT 2398.960 1701.610 2399.250 1702.930 ;
        RECT 2399.540 1701.610 2399.830 1702.930 ;
        RECT 2400.120 1701.610 2400.410 1702.930 ;
        RECT 2400.700 1701.610 2400.985 1702.930 ;
        RECT 2401.275 1701.610 2401.565 1702.930 ;
        RECT 2401.855 1701.610 2402.145 1702.930 ;
        RECT 2402.435 1701.610 2402.725 1702.930 ;
        RECT 2403.015 1701.610 2403.300 1702.930 ;
        RECT 2403.590 1701.610 2403.880 1702.930 ;
        RECT 2404.170 1701.610 2404.460 1702.930 ;
        RECT 2404.750 1701.610 2405.140 1702.930 ;
        RECT 2397.795 1701.605 2405.140 1701.610 ;
        RECT 2406.210 1701.605 2406.380 1702.235 ;
        RECT 2408.955 1701.605 2409.125 1702.235 ;
        RECT 2409.945 1701.605 2410.115 1702.235 ;
        RECT 2414.380 1701.615 2414.675 1702.935 ;
        RECT 2414.965 1701.615 2415.255 1702.935 ;
        RECT 2415.545 1701.615 2415.835 1702.935 ;
        RECT 2416.125 1701.615 2416.415 1702.935 ;
        RECT 2416.705 1701.615 2416.995 1702.935 ;
        RECT 2417.285 1701.615 2417.570 1702.935 ;
        RECT 2417.860 1701.615 2418.150 1702.935 ;
        RECT 2418.440 1701.615 2418.730 1702.935 ;
        RECT 2419.020 1701.615 2419.310 1702.935 ;
        RECT 2419.600 1701.615 2419.885 1702.935 ;
        RECT 2420.175 1701.615 2420.465 1702.935 ;
        RECT 2420.755 1701.615 2421.045 1702.935 ;
        RECT 2421.335 1701.615 2421.725 1702.935 ;
        RECT 2414.380 1701.610 2421.725 1701.615 ;
        RECT 2422.795 1701.610 2422.965 1702.240 ;
        RECT 2425.540 1701.610 2425.710 1702.240 ;
        RECT 2426.530 1701.610 2426.700 1702.240 ;
        RECT 2430.960 1701.615 2431.255 1702.935 ;
        RECT 2431.545 1701.615 2431.835 1702.935 ;
        RECT 2432.125 1701.615 2432.415 1702.935 ;
        RECT 2432.705 1701.615 2432.995 1702.935 ;
        RECT 2433.285 1701.615 2433.575 1702.935 ;
        RECT 2433.865 1701.615 2434.150 1702.935 ;
        RECT 2434.440 1701.615 2434.730 1702.935 ;
        RECT 2435.020 1701.615 2435.310 1702.935 ;
        RECT 2435.600 1701.615 2435.890 1702.935 ;
        RECT 2436.180 1701.615 2436.465 1702.935 ;
        RECT 2436.755 1701.615 2437.045 1702.935 ;
        RECT 2437.335 1701.615 2437.625 1702.935 ;
        RECT 2437.915 1701.615 2438.305 1702.935 ;
        RECT 2430.960 1701.610 2438.305 1701.615 ;
        RECT 2439.375 1701.610 2439.545 1702.240 ;
        RECT 2442.120 1701.610 2442.290 1702.240 ;
        RECT 2443.110 1701.610 2443.280 1702.240 ;
        RECT 2410.920 1701.605 2444.085 1701.610 ;
        RECT 2394.335 1701.600 2444.085 1701.605 ;
        RECT 2343.000 1700.000 2444.085 1701.600 ;
        RECT 2695.520 1676.835 2734.160 1677.005 ;
        RECT 2695.605 1676.085 2696.815 1676.835 ;
        RECT 2697.455 1676.355 2697.730 1676.835 ;
        RECT 2698.315 1676.435 2698.650 1676.835 ;
        RECT 2699.265 1676.455 2699.595 1676.835 ;
        RECT 2700.645 1676.455 2700.975 1676.835 ;
        RECT 2701.585 1676.290 2706.930 1676.835 ;
        RECT 2695.605 1675.545 2696.125 1676.085 ;
        RECT 2703.170 1675.460 2703.510 1676.290 ;
        RECT 2707.105 1676.085 2708.315 1676.835 ;
        RECT 2708.485 1676.110 2708.775 1676.835 ;
        RECT 2709.420 1676.455 2709.750 1676.835 ;
        RECT 2707.105 1675.545 2707.625 1676.085 ;
        RECT 2710.350 1675.995 2710.610 1676.835 ;
        RECT 2710.785 1676.290 2716.130 1676.835 ;
        RECT 2712.370 1675.460 2712.710 1676.290 ;
        RECT 2716.305 1676.065 2719.815 1676.835 ;
        RECT 2719.985 1676.085 2721.195 1676.835 ;
        RECT 2721.365 1676.110 2721.655 1676.835 ;
        RECT 2721.830 1676.435 2722.165 1676.835 ;
        RECT 2722.750 1676.355 2723.025 1676.835 ;
        RECT 2723.665 1676.290 2729.010 1676.835 ;
        RECT 2716.305 1675.545 2717.955 1676.065 ;
        RECT 2719.985 1675.545 2720.505 1676.085 ;
        RECT 2725.250 1675.460 2725.590 1676.290 ;
        RECT 2729.185 1676.065 2730.855 1676.835 ;
        RECT 2731.925 1676.455 2732.255 1676.835 ;
        RECT 2732.865 1676.085 2734.075 1676.835 ;
        RECT 2729.185 1675.545 2729.935 1676.065 ;
        RECT 2733.555 1675.545 2734.075 1676.085 ;
        RECT 2695.605 1672.315 2696.125 1672.855 ;
        RECT 2695.605 1671.565 2696.815 1672.315 ;
        RECT 2699.950 1672.110 2700.290 1672.940 ;
        RECT 2703.885 1672.335 2705.535 1672.855 ;
        RECT 2697.425 1671.565 2697.755 1671.945 ;
        RECT 2698.365 1671.565 2703.710 1672.110 ;
        RECT 2703.885 1671.565 2707.395 1672.335 ;
        RECT 2708.485 1671.565 2708.775 1672.290 ;
        RECT 2710.530 1672.110 2710.870 1672.940 ;
        RECT 2716.050 1672.110 2716.390 1672.940 ;
        RECT 2721.570 1672.110 2721.910 1672.940 ;
        RECT 2727.090 1672.110 2727.430 1672.940 ;
        RECT 2731.025 1672.335 2731.775 1672.855 ;
        RECT 2708.945 1671.565 2714.290 1672.110 ;
        RECT 2714.465 1671.565 2719.810 1672.110 ;
        RECT 2719.985 1671.565 2725.330 1672.110 ;
        RECT 2725.505 1671.565 2730.850 1672.110 ;
        RECT 2731.025 1671.565 2732.695 1672.335 ;
        RECT 2733.555 1672.315 2734.075 1672.855 ;
        RECT 2732.865 1671.565 2734.075 1672.315 ;
        RECT 2695.520 1671.395 2734.160 1671.565 ;
        RECT 2695.605 1670.645 2696.815 1671.395 ;
        RECT 2696.985 1670.850 2702.330 1671.395 ;
        RECT 2702.505 1670.850 2707.850 1671.395 ;
        RECT 2708.025 1670.850 2713.370 1671.395 ;
        RECT 2713.545 1670.850 2718.890 1671.395 ;
        RECT 2695.605 1670.105 2696.125 1670.645 ;
        RECT 2698.570 1670.020 2698.910 1670.850 ;
        RECT 2704.090 1670.020 2704.430 1670.850 ;
        RECT 2709.610 1670.020 2709.950 1670.850 ;
        RECT 2715.130 1670.020 2715.470 1670.850 ;
        RECT 2719.065 1670.625 2720.735 1671.395 ;
        RECT 2721.365 1670.670 2721.655 1671.395 ;
        RECT 2721.825 1670.850 2727.170 1671.395 ;
        RECT 2727.345 1670.850 2732.690 1671.395 ;
        RECT 2719.065 1670.105 2719.815 1670.625 ;
        RECT 2723.410 1670.020 2723.750 1670.850 ;
        RECT 2728.930 1670.020 2729.270 1670.850 ;
        RECT 2732.865 1670.645 2734.075 1671.395 ;
        RECT 2733.555 1670.105 2734.075 1670.645 ;
        RECT 2695.605 1666.875 2696.125 1667.415 ;
        RECT 2695.605 1666.125 2696.815 1666.875 ;
        RECT 2698.570 1666.670 2698.910 1667.500 ;
        RECT 2704.090 1666.670 2704.430 1667.500 ;
        RECT 2696.985 1666.125 2702.330 1666.670 ;
        RECT 2702.505 1666.125 2707.850 1666.670 ;
        RECT 2708.485 1666.125 2708.775 1666.850 ;
        RECT 2710.530 1666.670 2710.870 1667.500 ;
        RECT 2716.050 1666.670 2716.390 1667.500 ;
        RECT 2721.570 1666.670 2721.910 1667.500 ;
        RECT 2727.090 1666.670 2727.430 1667.500 ;
        RECT 2731.025 1666.895 2731.775 1667.415 ;
        RECT 2708.945 1666.125 2714.290 1666.670 ;
        RECT 2714.465 1666.125 2719.810 1666.670 ;
        RECT 2719.985 1666.125 2725.330 1666.670 ;
        RECT 2725.505 1666.125 2730.850 1666.670 ;
        RECT 2731.025 1666.125 2732.695 1666.895 ;
        RECT 2733.555 1666.875 2734.075 1667.415 ;
        RECT 2732.865 1666.125 2734.075 1666.875 ;
        RECT 2695.520 1665.955 2734.160 1666.125 ;
        RECT 2695.605 1665.205 2696.815 1665.955 ;
        RECT 2697.425 1665.575 2697.755 1665.955 ;
        RECT 2698.365 1665.410 2703.710 1665.955 ;
        RECT 2703.885 1665.410 2709.230 1665.955 ;
        RECT 2709.405 1665.410 2714.750 1665.955 ;
        RECT 2714.925 1665.410 2720.270 1665.955 ;
        RECT 2695.605 1664.665 2696.125 1665.205 ;
        RECT 2699.950 1664.580 2700.290 1665.410 ;
        RECT 2705.470 1664.580 2705.810 1665.410 ;
        RECT 2710.990 1664.580 2711.330 1665.410 ;
        RECT 2716.510 1664.580 2716.850 1665.410 ;
        RECT 2721.365 1665.230 2721.655 1665.955 ;
        RECT 2721.825 1665.410 2727.170 1665.955 ;
        RECT 2727.345 1665.410 2732.690 1665.955 ;
        RECT 2723.410 1664.580 2723.750 1665.410 ;
        RECT 2728.930 1664.580 2729.270 1665.410 ;
        RECT 2732.865 1665.205 2734.075 1665.955 ;
        RECT 2733.555 1664.665 2734.075 1665.205 ;
        RECT 2695.605 1661.435 2696.125 1661.975 ;
        RECT 2695.605 1660.685 2696.815 1661.435 ;
        RECT 2698.570 1661.230 2698.910 1662.060 ;
        RECT 2704.090 1661.230 2704.430 1662.060 ;
        RECT 2696.985 1660.685 2702.330 1661.230 ;
        RECT 2702.505 1660.685 2707.850 1661.230 ;
        RECT 2708.485 1660.685 2708.775 1661.410 ;
        RECT 2710.530 1661.230 2710.870 1662.060 ;
        RECT 2716.050 1661.230 2716.390 1662.060 ;
        RECT 2721.570 1661.230 2721.910 1662.060 ;
        RECT 2727.090 1661.230 2727.430 1662.060 ;
        RECT 2731.025 1661.455 2731.775 1661.975 ;
        RECT 2708.945 1660.685 2714.290 1661.230 ;
        RECT 2714.465 1660.685 2719.810 1661.230 ;
        RECT 2719.985 1660.685 2725.330 1661.230 ;
        RECT 2725.505 1660.685 2730.850 1661.230 ;
        RECT 2731.025 1660.685 2732.695 1661.455 ;
        RECT 2733.555 1661.435 2734.075 1661.975 ;
        RECT 2732.865 1660.685 2734.075 1661.435 ;
        RECT 2695.520 1660.515 2734.160 1660.685 ;
        RECT 2695.605 1659.765 2696.815 1660.515 ;
        RECT 2697.415 1660.135 2697.745 1660.515 ;
        RECT 2699.700 1659.795 2699.990 1660.515 ;
        RECT 2702.050 1660.055 2702.220 1660.515 ;
        RECT 2702.910 1660.135 2703.240 1660.515 ;
        RECT 2705.795 1660.055 2705.965 1660.515 ;
        RECT 2706.645 1659.970 2711.990 1660.515 ;
        RECT 2712.165 1659.970 2717.510 1660.515 ;
        RECT 2695.605 1659.225 2696.125 1659.765 ;
        RECT 2708.230 1659.140 2708.570 1659.970 ;
        RECT 2713.750 1659.140 2714.090 1659.970 ;
        RECT 2717.685 1659.745 2721.195 1660.515 ;
        RECT 2721.365 1659.790 2721.655 1660.515 ;
        RECT 2721.825 1659.970 2727.170 1660.515 ;
        RECT 2727.345 1659.970 2732.690 1660.515 ;
        RECT 2717.685 1659.225 2719.335 1659.745 ;
        RECT 2723.410 1659.140 2723.750 1659.970 ;
        RECT 2728.930 1659.140 2729.270 1659.970 ;
        RECT 2732.865 1659.765 2734.075 1660.515 ;
        RECT 2733.555 1659.225 2734.075 1659.765 ;
        RECT 2695.605 1655.995 2696.125 1656.535 ;
        RECT 2695.605 1655.245 2696.815 1655.995 ;
        RECT 2699.950 1655.790 2700.290 1656.620 ;
        RECT 2703.885 1656.015 2705.535 1656.535 ;
        RECT 2697.425 1655.245 2697.755 1655.625 ;
        RECT 2698.365 1655.245 2703.710 1655.790 ;
        RECT 2703.885 1655.245 2707.395 1656.015 ;
        RECT 2708.485 1655.245 2708.775 1655.970 ;
        RECT 2710.530 1655.790 2710.870 1656.620 ;
        RECT 2716.050 1655.790 2716.390 1656.620 ;
        RECT 2721.570 1655.790 2721.910 1656.620 ;
        RECT 2727.090 1655.790 2727.430 1656.620 ;
        RECT 2731.025 1656.015 2731.775 1656.535 ;
        RECT 2708.945 1655.245 2714.290 1655.790 ;
        RECT 2714.465 1655.245 2719.810 1655.790 ;
        RECT 2719.985 1655.245 2725.330 1655.790 ;
        RECT 2725.505 1655.245 2730.850 1655.790 ;
        RECT 2731.025 1655.245 2732.695 1656.015 ;
        RECT 2733.555 1655.995 2734.075 1656.535 ;
        RECT 2732.865 1655.245 2734.075 1655.995 ;
        RECT 2695.520 1655.075 2734.160 1655.245 ;
        RECT 2695.605 1654.325 2696.815 1655.075 ;
        RECT 2697.415 1654.695 2697.745 1655.075 ;
        RECT 2699.700 1654.355 2699.990 1655.075 ;
        RECT 2702.050 1654.615 2702.220 1655.075 ;
        RECT 2702.910 1654.695 2703.240 1655.075 ;
        RECT 2705.795 1654.615 2705.965 1655.075 ;
        RECT 2706.645 1654.530 2711.990 1655.075 ;
        RECT 2712.165 1654.530 2717.510 1655.075 ;
        RECT 2695.605 1653.785 2696.125 1654.325 ;
        RECT 2708.230 1653.700 2708.570 1654.530 ;
        RECT 2713.750 1653.700 2714.090 1654.530 ;
        RECT 2717.685 1654.305 2721.195 1655.075 ;
        RECT 2721.365 1654.350 2721.655 1655.075 ;
        RECT 2721.825 1654.530 2727.170 1655.075 ;
        RECT 2727.345 1654.530 2732.690 1655.075 ;
        RECT 2717.685 1653.785 2719.335 1654.305 ;
        RECT 2723.410 1653.700 2723.750 1654.530 ;
        RECT 2728.930 1653.700 2729.270 1654.530 ;
        RECT 2732.865 1654.325 2734.075 1655.075 ;
        RECT 2733.555 1653.785 2734.075 1654.325 ;
        RECT 2695.605 1650.555 2696.125 1651.095 ;
        RECT 2698.365 1650.575 2699.575 1651.095 ;
        RECT 2705.725 1650.575 2706.935 1651.095 ;
        RECT 2695.605 1649.805 2696.815 1650.555 ;
        RECT 2697.425 1649.805 2697.755 1650.185 ;
        RECT 2698.365 1649.805 2700.955 1650.575 ;
        RECT 2702.015 1649.805 2702.345 1650.205 ;
        RECT 2704.305 1649.805 2704.815 1650.340 ;
        RECT 2705.725 1649.805 2708.315 1650.575 ;
        RECT 2708.485 1649.805 2708.775 1650.530 ;
        RECT 2710.530 1650.350 2710.870 1651.180 ;
        RECT 2716.050 1650.350 2716.390 1651.180 ;
        RECT 2721.570 1650.350 2721.910 1651.180 ;
        RECT 2727.090 1650.350 2727.430 1651.180 ;
        RECT 2731.025 1650.575 2731.775 1651.095 ;
        RECT 2708.945 1649.805 2714.290 1650.350 ;
        RECT 2714.465 1649.805 2719.810 1650.350 ;
        RECT 2719.985 1649.805 2725.330 1650.350 ;
        RECT 2725.505 1649.805 2730.850 1650.350 ;
        RECT 2731.025 1649.805 2732.695 1650.575 ;
        RECT 2733.555 1650.555 2734.075 1651.095 ;
        RECT 2732.865 1649.805 2734.075 1650.555 ;
        RECT 2695.520 1649.635 2734.160 1649.805 ;
        RECT 2695.605 1648.885 2696.815 1649.635 ;
        RECT 2696.985 1649.090 2702.330 1649.635 ;
        RECT 2702.505 1649.090 2707.850 1649.635 ;
        RECT 2708.025 1649.090 2713.370 1649.635 ;
        RECT 2713.545 1649.090 2718.890 1649.635 ;
        RECT 2695.605 1648.345 2696.125 1648.885 ;
        RECT 2698.570 1648.260 2698.910 1649.090 ;
        RECT 2704.090 1648.260 2704.430 1649.090 ;
        RECT 2709.610 1648.260 2709.950 1649.090 ;
        RECT 2715.130 1648.260 2715.470 1649.090 ;
        RECT 2719.065 1648.865 2720.735 1649.635 ;
        RECT 2721.365 1648.910 2721.655 1649.635 ;
        RECT 2721.825 1649.090 2727.170 1649.635 ;
        RECT 2727.345 1649.090 2732.690 1649.635 ;
        RECT 2719.065 1648.345 2719.815 1648.865 ;
        RECT 2723.410 1648.260 2723.750 1649.090 ;
        RECT 2728.930 1648.260 2729.270 1649.090 ;
        RECT 2732.865 1648.885 2734.075 1649.635 ;
        RECT 2733.555 1648.345 2734.075 1648.885 ;
        RECT 2695.605 1645.115 2696.125 1645.655 ;
        RECT 2695.605 1644.365 2696.815 1645.115 ;
        RECT 2699.950 1644.910 2700.290 1645.740 ;
        RECT 2703.885 1645.135 2705.535 1645.655 ;
        RECT 2697.425 1644.365 2697.755 1644.745 ;
        RECT 2698.365 1644.365 2703.710 1644.910 ;
        RECT 2703.885 1644.365 2707.395 1645.135 ;
        RECT 2708.485 1644.365 2708.775 1645.090 ;
        RECT 2710.530 1644.910 2710.870 1645.740 ;
        RECT 2716.050 1644.910 2716.390 1645.740 ;
        RECT 2721.570 1644.910 2721.910 1645.740 ;
        RECT 2727.090 1644.910 2727.430 1645.740 ;
        RECT 2731.025 1645.135 2731.775 1645.655 ;
        RECT 2708.945 1644.365 2714.290 1644.910 ;
        RECT 2714.465 1644.365 2719.810 1644.910 ;
        RECT 2719.985 1644.365 2725.330 1644.910 ;
        RECT 2725.505 1644.365 2730.850 1644.910 ;
        RECT 2731.025 1644.365 2732.695 1645.135 ;
        RECT 2733.555 1645.115 2734.075 1645.655 ;
        RECT 2732.865 1644.365 2734.075 1645.115 ;
        RECT 2695.520 1644.195 2734.160 1644.365 ;
        RECT 2695.605 1643.445 2696.815 1644.195 ;
        RECT 2696.985 1643.650 2702.330 1644.195 ;
        RECT 2702.505 1643.650 2707.850 1644.195 ;
        RECT 2708.025 1643.650 2713.370 1644.195 ;
        RECT 2713.545 1643.650 2718.890 1644.195 ;
        RECT 2695.605 1642.905 2696.125 1643.445 ;
        RECT 2698.570 1642.820 2698.910 1643.650 ;
        RECT 2704.090 1642.820 2704.430 1643.650 ;
        RECT 2709.610 1642.820 2709.950 1643.650 ;
        RECT 2715.130 1642.820 2715.470 1643.650 ;
        RECT 2719.065 1643.425 2720.735 1644.195 ;
        RECT 2721.365 1643.470 2721.655 1644.195 ;
        RECT 2721.825 1643.650 2727.170 1644.195 ;
        RECT 2727.345 1643.650 2732.690 1644.195 ;
        RECT 2719.065 1642.905 2719.815 1643.425 ;
        RECT 2723.410 1642.820 2723.750 1643.650 ;
        RECT 2728.930 1642.820 2729.270 1643.650 ;
        RECT 2732.865 1643.445 2734.075 1644.195 ;
        RECT 2733.555 1642.905 2734.075 1643.445 ;
        RECT 2695.605 1639.675 2696.125 1640.215 ;
        RECT 2696.985 1639.695 2698.635 1640.215 ;
        RECT 2695.605 1638.925 2696.815 1639.675 ;
        RECT 2696.985 1638.925 2700.495 1639.695 ;
        RECT 2701.605 1638.925 2701.845 1639.735 ;
        RECT 2702.515 1638.925 2702.785 1639.735 ;
        RECT 2704.550 1639.470 2704.890 1640.300 ;
        RECT 2702.965 1638.925 2708.310 1639.470 ;
        RECT 2708.485 1638.925 2708.775 1639.650 ;
        RECT 2710.530 1639.470 2710.870 1640.300 ;
        RECT 2716.050 1639.470 2716.390 1640.300 ;
        RECT 2721.570 1639.470 2721.910 1640.300 ;
        RECT 2727.090 1639.470 2727.430 1640.300 ;
        RECT 2731.025 1639.695 2731.775 1640.215 ;
        RECT 2708.945 1638.925 2714.290 1639.470 ;
        RECT 2714.465 1638.925 2719.810 1639.470 ;
        RECT 2719.985 1638.925 2725.330 1639.470 ;
        RECT 2725.505 1638.925 2730.850 1639.470 ;
        RECT 2731.025 1638.925 2732.695 1639.695 ;
        RECT 2733.555 1639.675 2734.075 1640.215 ;
        RECT 2732.865 1638.925 2734.075 1639.675 ;
        RECT 2695.520 1638.755 2734.160 1638.925 ;
        RECT 2695.605 1638.005 2696.815 1638.755 ;
        RECT 2697.425 1638.375 2697.755 1638.755 ;
        RECT 2695.605 1637.465 2696.125 1638.005 ;
        RECT 2698.365 1637.985 2701.875 1638.755 ;
        RECT 2702.055 1638.015 2702.385 1638.755 ;
        RECT 2703.090 1638.395 2703.420 1638.755 ;
        RECT 2698.365 1637.465 2700.015 1637.985 ;
        RECT 2704.785 1637.975 2705.080 1638.755 ;
        RECT 2705.265 1638.210 2710.610 1638.755 ;
        RECT 2710.785 1638.210 2716.130 1638.755 ;
        RECT 2706.850 1637.380 2707.190 1638.210 ;
        RECT 2712.370 1637.380 2712.710 1638.210 ;
        RECT 2716.305 1637.985 2719.815 1638.755 ;
        RECT 2719.985 1638.005 2721.195 1638.755 ;
        RECT 2721.365 1638.030 2721.655 1638.755 ;
        RECT 2721.825 1638.210 2727.170 1638.755 ;
        RECT 2727.345 1638.210 2732.690 1638.755 ;
        RECT 2716.305 1637.465 2717.955 1637.985 ;
        RECT 2719.985 1637.465 2720.505 1638.005 ;
        RECT 2723.410 1637.380 2723.750 1638.210 ;
        RECT 2728.930 1637.380 2729.270 1638.210 ;
        RECT 2732.865 1638.005 2734.075 1638.755 ;
        RECT 2733.555 1637.465 2734.075 1638.005 ;
        RECT 2695.605 1634.235 2696.125 1634.775 ;
        RECT 2695.605 1633.485 2696.815 1634.235 ;
        RECT 2698.570 1634.030 2698.910 1634.860 ;
        RECT 2704.090 1634.030 2704.430 1634.860 ;
        RECT 2696.985 1633.485 2702.330 1634.030 ;
        RECT 2702.505 1633.485 2707.850 1634.030 ;
        RECT 2708.485 1633.485 2708.775 1634.210 ;
        RECT 2710.530 1634.030 2710.870 1634.860 ;
        RECT 2716.050 1634.030 2716.390 1634.860 ;
        RECT 2721.570 1634.030 2721.910 1634.860 ;
        RECT 2708.945 1633.485 2714.290 1634.030 ;
        RECT 2714.465 1633.485 2719.810 1634.030 ;
        RECT 2719.985 1633.485 2725.330 1634.030 ;
        RECT 2725.515 1633.485 2725.845 1633.965 ;
        RECT 2726.355 1633.485 2726.685 1633.965 ;
        RECT 2727.195 1633.485 2727.525 1633.965 ;
        RECT 2728.035 1633.485 2728.365 1633.965 ;
        RECT 2728.875 1633.485 2729.205 1633.965 ;
        RECT 2729.715 1633.485 2730.045 1633.965 ;
        RECT 2730.555 1633.485 2730.885 1633.965 ;
        RECT 2731.395 1633.485 2731.725 1633.965 ;
        RECT 2732.235 1633.485 2732.565 1634.285 ;
        RECT 2733.555 1634.235 2734.075 1634.775 ;
        RECT 2732.865 1633.485 2734.075 1634.235 ;
        RECT 2695.520 1633.315 2734.160 1633.485 ;
        RECT 2695.605 1632.565 2696.815 1633.315 ;
        RECT 2697.425 1632.935 2697.755 1633.315 ;
        RECT 2698.365 1632.770 2703.710 1633.315 ;
        RECT 2703.885 1632.770 2709.230 1633.315 ;
        RECT 2709.405 1632.770 2714.750 1633.315 ;
        RECT 2714.925 1632.770 2720.270 1633.315 ;
        RECT 2695.605 1632.025 2696.125 1632.565 ;
        RECT 2699.950 1631.940 2700.290 1632.770 ;
        RECT 2705.470 1631.940 2705.810 1632.770 ;
        RECT 2710.990 1631.940 2711.330 1632.770 ;
        RECT 2716.510 1631.940 2716.850 1632.770 ;
        RECT 2721.365 1632.590 2721.655 1633.315 ;
        RECT 2721.825 1632.770 2727.170 1633.315 ;
        RECT 2727.345 1632.770 2732.690 1633.315 ;
        RECT 2723.410 1631.940 2723.750 1632.770 ;
        RECT 2728.930 1631.940 2729.270 1632.770 ;
        RECT 2732.865 1632.565 2734.075 1633.315 ;
        RECT 2733.555 1632.025 2734.075 1632.565 ;
        RECT 2695.605 1628.795 2696.125 1629.335 ;
        RECT 2695.605 1628.045 2696.815 1628.795 ;
        RECT 2698.570 1628.590 2698.910 1629.420 ;
        RECT 2704.090 1628.590 2704.430 1629.420 ;
        RECT 2696.985 1628.045 2702.330 1628.590 ;
        RECT 2702.505 1628.045 2707.850 1628.590 ;
        RECT 2708.485 1628.045 2708.775 1628.770 ;
        RECT 2710.530 1628.590 2710.870 1629.420 ;
        RECT 2716.050 1628.590 2716.390 1629.420 ;
        RECT 2721.570 1628.590 2721.910 1629.420 ;
        RECT 2727.090 1628.590 2727.430 1629.420 ;
        RECT 2731.025 1628.815 2731.775 1629.335 ;
        RECT 2708.945 1628.045 2714.290 1628.590 ;
        RECT 2714.465 1628.045 2719.810 1628.590 ;
        RECT 2719.985 1628.045 2725.330 1628.590 ;
        RECT 2725.505 1628.045 2730.850 1628.590 ;
        RECT 2731.025 1628.045 2732.695 1628.815 ;
        RECT 2733.555 1628.795 2734.075 1629.335 ;
        RECT 2732.865 1628.045 2734.075 1628.795 ;
        RECT 2695.520 1627.875 2734.160 1628.045 ;
        RECT 2695.605 1627.125 2696.815 1627.875 ;
        RECT 2697.715 1627.135 2698.045 1627.875 ;
        RECT 2698.555 1627.475 2698.885 1627.875 ;
        RECT 2699.745 1627.330 2705.090 1627.875 ;
        RECT 2705.265 1627.330 2710.610 1627.875 ;
        RECT 2710.785 1627.330 2716.130 1627.875 ;
        RECT 2695.605 1626.585 2696.125 1627.125 ;
        RECT 2701.330 1626.500 2701.670 1627.330 ;
        RECT 2706.850 1626.500 2707.190 1627.330 ;
        RECT 2712.370 1626.500 2712.710 1627.330 ;
        RECT 2716.305 1627.105 2719.815 1627.875 ;
        RECT 2719.985 1627.125 2721.195 1627.875 ;
        RECT 2721.365 1627.150 2721.655 1627.875 ;
        RECT 2721.825 1627.330 2727.170 1627.875 ;
        RECT 2727.345 1627.330 2732.690 1627.875 ;
        RECT 2716.305 1626.585 2717.955 1627.105 ;
        RECT 2719.985 1626.585 2720.505 1627.125 ;
        RECT 2723.410 1626.500 2723.750 1627.330 ;
        RECT 2728.930 1626.500 2729.270 1627.330 ;
        RECT 2732.865 1627.125 2734.075 1627.875 ;
        RECT 2733.555 1626.585 2734.075 1627.125 ;
        RECT 2882.265 1625.790 2882.605 1626.450 ;
        RECT 2881.575 1625.620 2883.380 1625.790 ;
        RECT 2523.330 1623.680 2523.670 1624.340 ;
        RECT 2522.130 1623.510 2523.935 1623.680 ;
        RECT 2695.605 1623.355 2696.125 1623.895 ;
        RECT 2695.605 1622.605 2696.815 1623.355 ;
        RECT 2699.950 1623.150 2700.290 1623.980 ;
        RECT 2703.885 1623.375 2705.535 1623.895 ;
        RECT 2697.425 1622.605 2697.755 1622.985 ;
        RECT 2698.365 1622.605 2703.710 1623.150 ;
        RECT 2703.885 1622.605 2707.395 1623.375 ;
        RECT 2708.485 1622.605 2708.775 1623.330 ;
        RECT 2710.530 1623.150 2710.870 1623.980 ;
        RECT 2716.050 1623.150 2716.390 1623.980 ;
        RECT 2721.570 1623.150 2721.910 1623.980 ;
        RECT 2727.090 1623.150 2727.430 1623.980 ;
        RECT 2731.025 1623.375 2731.775 1623.895 ;
        RECT 2708.945 1622.605 2714.290 1623.150 ;
        RECT 2714.465 1622.605 2719.810 1623.150 ;
        RECT 2719.985 1622.605 2725.330 1623.150 ;
        RECT 2725.505 1622.605 2730.850 1623.150 ;
        RECT 2731.025 1622.605 2732.695 1623.375 ;
        RECT 2733.555 1623.355 2734.075 1623.895 ;
        RECT 2732.865 1622.605 2734.075 1623.355 ;
        RECT 2695.520 1622.435 2734.160 1622.605 ;
        RECT 2695.605 1621.685 2696.815 1622.435 ;
        RECT 2697.725 1621.900 2698.235 1622.435 ;
        RECT 2700.195 1622.035 2700.525 1622.435 ;
        RECT 2701.210 1621.760 2701.450 1622.435 ;
        RECT 2702.840 1621.985 2703.170 1622.435 ;
        RECT 2704.090 1621.995 2704.405 1622.435 ;
        RECT 2704.805 1621.890 2710.150 1622.435 ;
        RECT 2710.325 1621.890 2715.670 1622.435 ;
        RECT 2715.845 1621.890 2721.190 1622.435 ;
        RECT 2695.605 1621.145 2696.125 1621.685 ;
        RECT 2706.390 1621.060 2706.730 1621.890 ;
        RECT 2711.910 1621.060 2712.250 1621.890 ;
        RECT 2717.430 1621.060 2717.770 1621.890 ;
        RECT 2721.365 1621.710 2721.655 1622.435 ;
        RECT 2721.825 1621.890 2727.170 1622.435 ;
        RECT 2727.345 1621.890 2732.690 1622.435 ;
        RECT 2723.410 1621.060 2723.750 1621.890 ;
        RECT 2728.930 1621.060 2729.270 1621.890 ;
        RECT 2732.865 1621.685 2734.075 1622.435 ;
        RECT 2733.555 1621.145 2734.075 1621.685 ;
        RECT 2523.330 1617.265 2523.670 1617.925 ;
        RECT 2695.605 1617.915 2696.125 1618.455 ;
        RECT 2522.130 1617.095 2523.935 1617.265 ;
        RECT 2695.605 1617.165 2696.815 1617.915 ;
        RECT 2696.985 1617.165 2697.245 1617.985 ;
        RECT 2701.790 1617.710 2702.130 1618.540 ;
        RECT 2705.725 1617.935 2706.935 1618.455 ;
        RECT 2699.275 1617.165 2699.605 1617.625 ;
        RECT 2700.205 1617.165 2705.550 1617.710 ;
        RECT 2705.725 1617.165 2708.315 1617.935 ;
        RECT 2708.485 1617.165 2708.775 1617.890 ;
        RECT 2710.530 1617.710 2710.870 1618.540 ;
        RECT 2716.050 1617.710 2716.390 1618.540 ;
        RECT 2721.570 1617.710 2721.910 1618.540 ;
        RECT 2727.090 1617.710 2727.430 1618.540 ;
        RECT 2731.025 1617.935 2731.775 1618.455 ;
        RECT 2708.945 1617.165 2714.290 1617.710 ;
        RECT 2714.465 1617.165 2719.810 1617.710 ;
        RECT 2719.985 1617.165 2725.330 1617.710 ;
        RECT 2725.505 1617.165 2730.850 1617.710 ;
        RECT 2731.025 1617.165 2732.695 1617.935 ;
        RECT 2733.555 1617.915 2734.075 1618.455 ;
        RECT 2732.865 1617.165 2734.075 1617.915 ;
        RECT 2695.520 1616.995 2734.160 1617.165 ;
        RECT 2695.605 1616.245 2696.815 1616.995 ;
        RECT 2697.425 1616.615 2697.755 1616.995 ;
        RECT 2698.365 1616.450 2703.710 1616.995 ;
        RECT 2703.885 1616.450 2709.230 1616.995 ;
        RECT 2709.405 1616.450 2714.750 1616.995 ;
        RECT 2714.925 1616.450 2720.270 1616.995 ;
        RECT 2695.605 1615.705 2696.125 1616.245 ;
        RECT 2699.950 1615.620 2700.290 1616.450 ;
        RECT 2705.470 1615.620 2705.810 1616.450 ;
        RECT 2710.990 1615.620 2711.330 1616.450 ;
        RECT 2716.510 1615.620 2716.850 1616.450 ;
        RECT 2721.365 1616.270 2721.655 1616.995 ;
        RECT 2721.825 1616.450 2727.170 1616.995 ;
        RECT 2727.345 1616.450 2732.690 1616.995 ;
        RECT 2723.410 1615.620 2723.750 1616.450 ;
        RECT 2728.930 1615.620 2729.270 1616.450 ;
        RECT 2732.865 1616.245 2734.075 1616.995 ;
        RECT 2733.555 1615.705 2734.075 1616.245 ;
        RECT 2695.605 1612.475 2696.125 1613.015 ;
        RECT 2696.985 1612.475 2697.505 1613.015 ;
        RECT 2395.235 1612.460 2412.475 1612.465 ;
        RECT 2343.045 1610.860 2446.915 1612.460 ;
        RECT 2695.605 1611.725 2696.815 1612.475 ;
        RECT 2696.985 1611.725 2698.195 1612.475 ;
        RECT 2698.365 1611.725 2698.705 1612.450 ;
        RECT 2703.630 1612.270 2703.970 1613.100 ;
        RECT 2701.035 1611.725 2701.365 1612.205 ;
        RECT 2702.045 1611.725 2707.390 1612.270 ;
        RECT 2708.485 1611.725 2708.775 1612.450 ;
        RECT 2710.530 1612.270 2710.870 1613.100 ;
        RECT 2716.050 1612.270 2716.390 1613.100 ;
        RECT 2721.570 1612.270 2721.910 1613.100 ;
        RECT 2727.090 1612.270 2727.430 1613.100 ;
        RECT 2731.025 1612.495 2731.775 1613.015 ;
        RECT 2708.945 1611.725 2714.290 1612.270 ;
        RECT 2714.465 1611.725 2719.810 1612.270 ;
        RECT 2719.985 1611.725 2725.330 1612.270 ;
        RECT 2725.505 1611.725 2730.850 1612.270 ;
        RECT 2731.025 1611.725 2732.695 1612.495 ;
        RECT 2733.555 1612.475 2734.075 1613.015 ;
        RECT 2732.865 1611.725 2734.075 1612.475 ;
        RECT 2695.520 1611.555 2734.160 1611.725 ;
        RECT 2358.215 1610.235 2358.385 1610.860 ;
        RECT 2361.625 1610.235 2361.795 1610.860 ;
        RECT 2362.580 1610.315 2362.750 1610.595 ;
        RECT 2362.580 1610.145 2362.810 1610.315 ;
        RECT 2362.640 1608.535 2362.810 1610.145 ;
        RECT 2362.580 1608.365 2362.810 1608.535 ;
        RECT 2364.585 1608.530 2364.910 1610.860 ;
        RECT 2365.235 1608.530 2365.560 1610.860 ;
        RECT 2365.885 1608.530 2366.210 1610.860 ;
        RECT 2366.535 1608.530 2366.860 1610.860 ;
        RECT 2367.185 1608.530 2367.510 1610.860 ;
        RECT 2367.835 1608.530 2368.160 1610.860 ;
        RECT 2368.485 1608.530 2368.810 1610.860 ;
        RECT 2369.135 1608.530 2369.460 1610.860 ;
        RECT 2369.785 1608.530 2370.110 1610.860 ;
        RECT 2370.435 1608.530 2370.760 1610.860 ;
        RECT 2371.085 1608.530 2371.410 1610.860 ;
        RECT 2371.735 1608.530 2371.945 1610.860 ;
        RECT 2373.310 1610.235 2373.480 1610.860 ;
        RECT 2376.055 1610.235 2376.225 1610.860 ;
        RECT 2377.045 1610.235 2377.215 1610.860 ;
        RECT 2378.845 1610.235 2379.015 1610.860 ;
        RECT 2379.800 1610.315 2379.970 1610.595 ;
        RECT 2379.800 1610.145 2380.030 1610.315 ;
        RECT 2379.860 1608.535 2380.030 1610.145 ;
        RECT 2362.580 1607.305 2362.750 1608.365 ;
        RECT 2364.585 1608.360 2371.945 1608.530 ;
        RECT 2379.800 1608.365 2380.030 1608.535 ;
        RECT 2381.805 1608.530 2382.130 1610.860 ;
        RECT 2382.455 1608.530 2382.780 1610.860 ;
        RECT 2383.105 1608.530 2383.430 1610.860 ;
        RECT 2383.755 1608.530 2384.080 1610.860 ;
        RECT 2384.405 1608.530 2384.730 1610.860 ;
        RECT 2385.055 1608.530 2385.380 1610.860 ;
        RECT 2385.705 1608.530 2386.030 1610.860 ;
        RECT 2386.355 1608.530 2386.680 1610.860 ;
        RECT 2387.005 1608.530 2387.330 1610.860 ;
        RECT 2387.655 1608.530 2387.980 1610.860 ;
        RECT 2388.305 1608.530 2388.630 1610.860 ;
        RECT 2388.955 1608.530 2389.165 1610.860 ;
        RECT 2390.530 1610.235 2390.700 1610.860 ;
        RECT 2393.275 1610.235 2393.445 1610.860 ;
        RECT 2394.265 1610.235 2394.435 1610.860 ;
        RECT 2396.065 1610.240 2396.235 1610.860 ;
        RECT 2397.020 1610.320 2397.190 1610.600 ;
        RECT 2397.020 1610.150 2397.250 1610.320 ;
        RECT 2397.080 1608.540 2397.250 1610.150 ;
        RECT 2365.130 1607.560 2365.440 1608.360 ;
        RECT 2365.140 1607.340 2365.475 1607.390 ;
        RECT 2367.060 1607.340 2367.230 1608.360 ;
        RECT 2367.430 1607.560 2367.740 1608.360 ;
        RECT 2369.710 1607.560 2370.020 1608.360 ;
        RECT 2371.090 1607.560 2371.400 1608.360 ;
        RECT 2367.440 1607.340 2367.775 1607.390 ;
        RECT 2364.670 1607.170 2365.475 1607.340 ;
        RECT 2367.050 1607.170 2367.775 1607.340 ;
        RECT 2379.800 1607.305 2379.970 1608.365 ;
        RECT 2381.805 1608.360 2389.165 1608.530 ;
        RECT 2397.020 1608.370 2397.250 1608.540 ;
        RECT 2399.025 1608.535 2399.350 1610.860 ;
        RECT 2399.675 1608.535 2400.000 1610.860 ;
        RECT 2400.325 1608.535 2400.650 1610.860 ;
        RECT 2400.975 1608.535 2401.300 1610.860 ;
        RECT 2401.625 1608.535 2401.950 1610.860 ;
        RECT 2402.275 1608.535 2402.600 1610.860 ;
        RECT 2402.925 1608.535 2403.250 1610.860 ;
        RECT 2403.575 1608.535 2403.900 1610.860 ;
        RECT 2404.225 1608.535 2404.550 1610.860 ;
        RECT 2404.875 1608.535 2405.200 1610.860 ;
        RECT 2405.525 1608.535 2405.850 1610.860 ;
        RECT 2406.175 1608.535 2406.385 1610.860 ;
        RECT 2407.750 1610.240 2407.920 1610.860 ;
        RECT 2410.495 1610.240 2410.665 1610.860 ;
        RECT 2411.485 1610.240 2411.655 1610.860 ;
        RECT 2413.285 1610.235 2413.455 1610.860 ;
        RECT 2414.240 1610.315 2414.410 1610.595 ;
        RECT 2414.240 1610.145 2414.470 1610.315 ;
        RECT 2414.300 1608.535 2414.470 1610.145 ;
        RECT 2382.350 1607.560 2382.660 1608.360 ;
        RECT 2382.360 1607.340 2382.695 1607.390 ;
        RECT 2384.280 1607.340 2384.450 1608.360 ;
        RECT 2384.650 1607.560 2384.960 1608.360 ;
        RECT 2386.930 1607.560 2387.240 1608.360 ;
        RECT 2388.310 1607.560 2388.620 1608.360 ;
        RECT 2384.660 1607.340 2384.995 1607.390 ;
        RECT 2381.890 1607.170 2382.695 1607.340 ;
        RECT 2384.270 1607.170 2384.995 1607.340 ;
        RECT 2397.020 1607.310 2397.190 1608.370 ;
        RECT 2399.025 1608.365 2406.385 1608.535 ;
        RECT 2414.240 1608.365 2414.470 1608.535 ;
        RECT 2416.245 1608.530 2416.570 1610.860 ;
        RECT 2416.895 1608.530 2417.220 1610.860 ;
        RECT 2417.545 1608.530 2417.870 1610.860 ;
        RECT 2418.195 1608.530 2418.520 1610.860 ;
        RECT 2418.845 1608.530 2419.170 1610.860 ;
        RECT 2419.495 1608.530 2419.820 1610.860 ;
        RECT 2420.145 1608.530 2420.470 1610.860 ;
        RECT 2420.795 1608.530 2421.120 1610.860 ;
        RECT 2421.445 1608.530 2421.770 1610.860 ;
        RECT 2422.095 1608.530 2422.420 1610.860 ;
        RECT 2422.745 1608.530 2423.070 1610.860 ;
        RECT 2423.395 1608.530 2423.605 1610.860 ;
        RECT 2424.970 1610.235 2425.140 1610.860 ;
        RECT 2427.715 1610.235 2427.885 1610.860 ;
        RECT 2428.705 1610.235 2428.875 1610.860 ;
        RECT 2430.505 1610.235 2430.675 1610.860 ;
        RECT 2431.460 1610.315 2431.630 1610.595 ;
        RECT 2431.460 1610.145 2431.690 1610.315 ;
        RECT 2431.520 1608.535 2431.690 1610.145 ;
        RECT 2399.570 1607.565 2399.880 1608.365 ;
        RECT 2399.580 1607.345 2399.915 1607.395 ;
        RECT 2401.500 1607.345 2401.670 1608.365 ;
        RECT 2401.870 1607.565 2402.180 1608.365 ;
        RECT 2404.150 1607.565 2404.460 1608.365 ;
        RECT 2405.530 1607.565 2405.840 1608.365 ;
        RECT 2401.880 1607.345 2402.215 1607.395 ;
        RECT 2399.110 1607.175 2399.915 1607.345 ;
        RECT 2401.490 1607.175 2402.215 1607.345 ;
        RECT 2414.240 1607.305 2414.410 1608.365 ;
        RECT 2416.245 1608.360 2423.605 1608.530 ;
        RECT 2431.460 1608.365 2431.690 1608.535 ;
        RECT 2433.465 1608.530 2433.790 1610.860 ;
        RECT 2434.115 1608.530 2434.440 1610.860 ;
        RECT 2434.765 1608.530 2435.090 1610.860 ;
        RECT 2435.415 1608.530 2435.740 1610.860 ;
        RECT 2436.065 1608.530 2436.390 1610.860 ;
        RECT 2436.715 1608.530 2437.040 1610.860 ;
        RECT 2437.365 1608.530 2437.690 1610.860 ;
        RECT 2438.015 1608.530 2438.340 1610.860 ;
        RECT 2438.665 1608.530 2438.990 1610.860 ;
        RECT 2439.315 1608.530 2439.640 1610.860 ;
        RECT 2439.965 1608.530 2440.290 1610.860 ;
        RECT 2440.615 1608.530 2440.825 1610.860 ;
        RECT 2442.190 1610.235 2442.360 1610.860 ;
        RECT 2444.935 1610.235 2445.105 1610.860 ;
        RECT 2445.925 1610.235 2446.095 1610.860 ;
        RECT 2695.605 1610.805 2696.815 1611.555 ;
        RECT 2695.605 1610.265 2696.125 1610.805 ;
        RECT 2697.905 1610.735 2698.165 1611.555 ;
        RECT 2699.275 1611.155 2699.605 1611.555 ;
        RECT 2700.115 1611.155 2700.490 1611.555 ;
        RECT 2702.760 1611.155 2703.090 1611.555 ;
        RECT 2703.885 1611.010 2709.230 1611.555 ;
        RECT 2709.405 1611.010 2714.750 1611.555 ;
        RECT 2714.925 1611.010 2720.270 1611.555 ;
        RECT 2705.470 1610.180 2705.810 1611.010 ;
        RECT 2710.990 1610.180 2711.330 1611.010 ;
        RECT 2716.510 1610.180 2716.850 1611.010 ;
        RECT 2721.365 1610.830 2721.655 1611.555 ;
        RECT 2721.825 1611.010 2727.170 1611.555 ;
        RECT 2727.345 1611.010 2732.690 1611.555 ;
        RECT 2723.410 1610.180 2723.750 1611.010 ;
        RECT 2728.930 1610.180 2729.270 1611.010 ;
        RECT 2732.865 1610.805 2734.075 1611.555 ;
        RECT 2733.555 1610.265 2734.075 1610.805 ;
        RECT 2416.790 1607.560 2417.100 1608.360 ;
        RECT 2416.800 1607.340 2417.135 1607.390 ;
        RECT 2418.720 1607.340 2418.890 1608.360 ;
        RECT 2419.090 1607.560 2419.400 1608.360 ;
        RECT 2421.370 1607.560 2421.680 1608.360 ;
        RECT 2422.750 1607.560 2423.060 1608.360 ;
        RECT 2419.100 1607.340 2419.435 1607.390 ;
        RECT 2365.140 1607.120 2365.475 1607.170 ;
        RECT 2367.440 1607.120 2367.775 1607.170 ;
        RECT 2382.360 1607.120 2382.695 1607.170 ;
        RECT 2384.660 1607.120 2384.995 1607.170 ;
        RECT 2399.580 1607.125 2399.915 1607.175 ;
        RECT 2401.880 1607.125 2402.215 1607.175 ;
        RECT 2416.330 1607.170 2417.135 1607.340 ;
        RECT 2418.710 1607.170 2419.435 1607.340 ;
        RECT 2431.460 1607.305 2431.630 1608.365 ;
        RECT 2433.465 1608.360 2440.825 1608.530 ;
        RECT 2434.010 1607.560 2434.320 1608.360 ;
        RECT 2434.020 1607.340 2434.355 1607.390 ;
        RECT 2435.940 1607.340 2436.110 1608.360 ;
        RECT 2436.310 1607.560 2436.620 1608.360 ;
        RECT 2438.590 1607.560 2438.900 1608.360 ;
        RECT 2439.970 1607.560 2440.280 1608.360 ;
        RECT 2436.320 1607.340 2436.655 1607.390 ;
        RECT 2433.550 1607.170 2434.355 1607.340 ;
        RECT 2435.930 1607.170 2436.655 1607.340 ;
        RECT 2416.800 1607.120 2417.135 1607.170 ;
        RECT 2419.100 1607.120 2419.435 1607.170 ;
        RECT 2434.020 1607.120 2434.355 1607.170 ;
        RECT 2436.320 1607.120 2436.655 1607.170 ;
        RECT 2695.605 1607.035 2696.125 1607.575 ;
        RECT 2695.605 1606.285 2696.815 1607.035 ;
        RECT 2697.425 1606.285 2697.755 1606.665 ;
        RECT 2699.725 1606.285 2700.035 1607.085 ;
        RECT 2701.790 1606.830 2702.130 1607.660 ;
        RECT 2705.725 1607.055 2706.935 1607.575 ;
        RECT 2700.205 1606.285 2705.550 1606.830 ;
        RECT 2705.725 1606.285 2708.315 1607.055 ;
        RECT 2708.485 1606.285 2708.775 1607.010 ;
        RECT 2710.530 1606.830 2710.870 1607.660 ;
        RECT 2716.050 1606.830 2716.390 1607.660 ;
        RECT 2721.570 1606.830 2721.910 1607.660 ;
        RECT 2727.090 1606.830 2727.430 1607.660 ;
        RECT 2731.025 1607.055 2731.775 1607.575 ;
        RECT 2708.945 1606.285 2714.290 1606.830 ;
        RECT 2714.465 1606.285 2719.810 1606.830 ;
        RECT 2719.985 1606.285 2725.330 1606.830 ;
        RECT 2725.505 1606.285 2730.850 1606.830 ;
        RECT 2731.025 1606.285 2732.695 1607.055 ;
        RECT 2733.555 1607.035 2734.075 1607.575 ;
        RECT 2732.865 1606.285 2734.075 1607.035 ;
        RECT 2695.520 1606.115 2734.160 1606.285 ;
        RECT 2695.605 1605.365 2696.815 1606.115 ;
        RECT 2697.725 1605.580 2698.235 1606.115 ;
        RECT 2700.195 1605.715 2700.525 1606.115 ;
        RECT 2701.125 1605.570 2706.470 1606.115 ;
        RECT 2706.645 1605.570 2711.990 1606.115 ;
        RECT 2712.165 1605.570 2717.510 1606.115 ;
        RECT 2695.605 1604.825 2696.125 1605.365 ;
        RECT 2702.710 1604.740 2703.050 1605.570 ;
        RECT 2708.230 1604.740 2708.570 1605.570 ;
        RECT 2713.750 1604.740 2714.090 1605.570 ;
        RECT 2717.685 1605.345 2721.195 1606.115 ;
        RECT 2721.365 1605.390 2721.655 1606.115 ;
        RECT 2721.825 1605.570 2727.170 1606.115 ;
        RECT 2727.345 1605.570 2732.690 1606.115 ;
        RECT 2717.685 1604.825 2719.335 1605.345 ;
        RECT 2723.410 1604.740 2723.750 1605.570 ;
        RECT 2728.930 1604.740 2729.270 1605.570 ;
        RECT 2732.865 1605.365 2734.075 1606.115 ;
        RECT 2733.555 1604.825 2734.075 1605.365 ;
        RECT 2364.730 1603.090 2364.940 1603.910 ;
        RECT 2365.610 1603.090 2365.840 1603.910 ;
        RECT 2366.060 1603.090 2366.330 1603.900 ;
        RECT 2367.000 1603.090 2367.240 1603.900 ;
        RECT 2367.450 1603.090 2367.690 1603.900 ;
        RECT 2368.360 1603.090 2368.630 1603.900 ;
        RECT 2368.810 1603.090 2369.100 1603.925 ;
        RECT 2370.640 1603.090 2370.970 1603.480 ;
        RECT 2371.480 1603.090 2371.810 1603.480 ;
        RECT 2381.950 1603.090 2382.160 1603.910 ;
        RECT 2382.830 1603.090 2383.060 1603.910 ;
        RECT 2383.280 1603.090 2383.550 1603.900 ;
        RECT 2384.220 1603.090 2384.460 1603.900 ;
        RECT 2384.670 1603.090 2384.910 1603.900 ;
        RECT 2385.580 1603.090 2385.850 1603.900 ;
        RECT 2386.030 1603.090 2386.320 1603.925 ;
        RECT 2387.860 1603.090 2388.190 1603.480 ;
        RECT 2388.700 1603.090 2389.030 1603.480 ;
        RECT 2399.170 1603.095 2399.380 1603.915 ;
        RECT 2400.050 1603.095 2400.280 1603.915 ;
        RECT 2400.500 1603.095 2400.770 1603.905 ;
        RECT 2401.440 1603.095 2401.680 1603.905 ;
        RECT 2401.890 1603.095 2402.130 1603.905 ;
        RECT 2402.800 1603.095 2403.070 1603.905 ;
        RECT 2403.250 1603.095 2403.540 1603.930 ;
        RECT 2405.080 1603.095 2405.410 1603.485 ;
        RECT 2405.920 1603.095 2406.250 1603.485 ;
        RECT 2364.580 1602.920 2372.325 1603.090 ;
        RECT 2364.580 1601.600 2364.925 1602.920 ;
        RECT 2365.270 1601.600 2365.600 1602.920 ;
        RECT 2365.945 1601.605 2366.290 1602.920 ;
        RECT 2366.635 1601.605 2366.980 1602.920 ;
        RECT 2367.325 1601.605 2367.670 1602.920 ;
        RECT 2368.015 1601.605 2368.360 1602.920 ;
        RECT 2368.705 1601.605 2369.050 1602.920 ;
        RECT 2369.395 1601.605 2369.740 1602.920 ;
        RECT 2370.085 1601.605 2370.430 1602.920 ;
        RECT 2370.775 1601.605 2371.120 1602.920 ;
        RECT 2371.465 1601.605 2371.810 1602.920 ;
        RECT 2372.155 1601.605 2372.325 1602.920 ;
        RECT 2381.800 1602.920 2389.545 1603.090 ;
        RECT 2365.945 1601.600 2372.325 1601.605 ;
        RECT 2373.310 1601.600 2373.480 1602.225 ;
        RECT 2376.055 1601.600 2376.225 1602.225 ;
        RECT 2377.040 1601.600 2377.210 1602.225 ;
        RECT 2381.800 1601.600 2382.145 1602.920 ;
        RECT 2382.490 1601.600 2382.820 1602.920 ;
        RECT 2383.165 1601.605 2383.510 1602.920 ;
        RECT 2383.855 1601.605 2384.200 1602.920 ;
        RECT 2384.545 1601.605 2384.890 1602.920 ;
        RECT 2385.235 1601.605 2385.580 1602.920 ;
        RECT 2385.925 1601.605 2386.270 1602.920 ;
        RECT 2386.615 1601.605 2386.960 1602.920 ;
        RECT 2387.305 1601.605 2387.650 1602.920 ;
        RECT 2387.995 1601.605 2388.340 1602.920 ;
        RECT 2388.685 1601.605 2389.030 1602.920 ;
        RECT 2389.375 1601.605 2389.545 1602.920 ;
        RECT 2399.020 1602.925 2406.765 1603.095 ;
        RECT 2416.390 1603.090 2416.600 1603.910 ;
        RECT 2417.270 1603.090 2417.500 1603.910 ;
        RECT 2417.720 1603.090 2417.990 1603.900 ;
        RECT 2418.660 1603.090 2418.900 1603.900 ;
        RECT 2419.110 1603.090 2419.350 1603.900 ;
        RECT 2420.020 1603.090 2420.290 1603.900 ;
        RECT 2420.470 1603.090 2420.760 1603.925 ;
        RECT 2422.300 1603.090 2422.630 1603.480 ;
        RECT 2423.140 1603.090 2423.470 1603.480 ;
        RECT 2433.610 1603.090 2433.820 1603.910 ;
        RECT 2434.490 1603.090 2434.720 1603.910 ;
        RECT 2434.940 1603.090 2435.210 1603.900 ;
        RECT 2435.880 1603.090 2436.120 1603.900 ;
        RECT 2436.330 1603.090 2436.570 1603.900 ;
        RECT 2437.240 1603.090 2437.510 1603.900 ;
        RECT 2437.690 1603.090 2437.980 1603.925 ;
        RECT 2439.520 1603.090 2439.850 1603.480 ;
        RECT 2440.360 1603.090 2440.690 1603.480 ;
        RECT 2383.165 1601.600 2389.545 1601.605 ;
        RECT 2390.530 1601.600 2390.700 1602.225 ;
        RECT 2393.275 1601.600 2393.445 1602.225 ;
        RECT 2394.260 1601.600 2394.430 1602.225 ;
        RECT 2399.020 1601.605 2399.365 1602.925 ;
        RECT 2399.710 1601.605 2400.040 1602.925 ;
        RECT 2400.385 1601.610 2400.730 1602.925 ;
        RECT 2401.075 1601.610 2401.420 1602.925 ;
        RECT 2401.765 1601.610 2402.110 1602.925 ;
        RECT 2402.455 1601.610 2402.800 1602.925 ;
        RECT 2403.145 1601.610 2403.490 1602.925 ;
        RECT 2403.835 1601.610 2404.180 1602.925 ;
        RECT 2404.525 1601.610 2404.870 1602.925 ;
        RECT 2405.215 1601.610 2405.560 1602.925 ;
        RECT 2405.905 1601.610 2406.250 1602.925 ;
        RECT 2406.595 1601.610 2406.765 1602.925 ;
        RECT 2416.240 1602.920 2423.985 1603.090 ;
        RECT 2400.385 1601.605 2406.765 1601.610 ;
        RECT 2407.750 1601.605 2407.920 1602.230 ;
        RECT 2410.495 1601.605 2410.665 1602.230 ;
        RECT 2411.480 1601.605 2411.650 1602.230 ;
        RECT 2395.235 1601.600 2412.475 1601.605 ;
        RECT 2416.240 1601.600 2416.585 1602.920 ;
        RECT 2416.930 1601.600 2417.260 1602.920 ;
        RECT 2417.605 1601.605 2417.950 1602.920 ;
        RECT 2418.295 1601.605 2418.640 1602.920 ;
        RECT 2418.985 1601.605 2419.330 1602.920 ;
        RECT 2419.675 1601.605 2420.020 1602.920 ;
        RECT 2420.365 1601.605 2420.710 1602.920 ;
        RECT 2421.055 1601.605 2421.400 1602.920 ;
        RECT 2421.745 1601.605 2422.090 1602.920 ;
        RECT 2422.435 1601.605 2422.780 1602.920 ;
        RECT 2423.125 1601.605 2423.470 1602.920 ;
        RECT 2423.815 1601.605 2423.985 1602.920 ;
        RECT 2433.460 1602.920 2441.205 1603.090 ;
        RECT 2417.605 1601.600 2423.985 1601.605 ;
        RECT 2424.970 1601.600 2425.140 1602.225 ;
        RECT 2427.715 1601.600 2427.885 1602.225 ;
        RECT 2428.700 1601.600 2428.870 1602.225 ;
        RECT 2433.460 1601.600 2433.805 1602.920 ;
        RECT 2434.150 1601.600 2434.480 1602.920 ;
        RECT 2434.825 1601.605 2435.170 1602.920 ;
        RECT 2435.515 1601.605 2435.860 1602.920 ;
        RECT 2436.205 1601.605 2436.550 1602.920 ;
        RECT 2436.895 1601.605 2437.240 1602.920 ;
        RECT 2437.585 1601.605 2437.930 1602.920 ;
        RECT 2438.275 1601.605 2438.620 1602.920 ;
        RECT 2438.965 1601.605 2439.310 1602.920 ;
        RECT 2439.655 1601.605 2440.000 1602.920 ;
        RECT 2440.345 1601.605 2440.690 1602.920 ;
        RECT 2441.035 1601.605 2441.205 1602.920 ;
        RECT 2434.825 1601.600 2441.205 1601.605 ;
        RECT 2442.190 1601.600 2442.360 1602.225 ;
        RECT 2444.935 1601.600 2445.105 1602.225 ;
        RECT 2445.920 1601.600 2446.090 1602.225 ;
        RECT 2343.045 1600.000 2446.915 1601.600 ;
        RECT 2695.605 1601.595 2696.125 1602.135 ;
        RECT 2695.605 1600.845 2696.815 1601.595 ;
        RECT 2699.950 1601.390 2700.290 1602.220 ;
        RECT 2703.885 1601.615 2705.535 1602.135 ;
        RECT 2697.425 1600.845 2697.755 1601.225 ;
        RECT 2698.365 1600.845 2703.710 1601.390 ;
        RECT 2703.885 1600.845 2707.395 1601.615 ;
        RECT 2708.485 1600.845 2708.775 1601.570 ;
        RECT 2710.530 1601.390 2710.870 1602.220 ;
        RECT 2716.050 1601.390 2716.390 1602.220 ;
        RECT 2721.570 1601.390 2721.910 1602.220 ;
        RECT 2727.090 1601.390 2727.430 1602.220 ;
        RECT 2731.025 1601.615 2731.775 1602.135 ;
        RECT 2708.945 1600.845 2714.290 1601.390 ;
        RECT 2714.465 1600.845 2719.810 1601.390 ;
        RECT 2719.985 1600.845 2725.330 1601.390 ;
        RECT 2725.505 1600.845 2730.850 1601.390 ;
        RECT 2731.025 1600.845 2732.695 1601.615 ;
        RECT 2733.555 1601.595 2734.075 1602.135 ;
        RECT 2732.865 1600.845 2734.075 1601.595 ;
        RECT 2695.520 1600.675 2734.160 1600.845 ;
        RECT 2695.605 1599.925 2696.815 1600.675 ;
        RECT 2696.985 1600.130 2702.330 1600.675 ;
        RECT 2702.505 1600.130 2707.850 1600.675 ;
        RECT 2708.025 1600.130 2713.370 1600.675 ;
        RECT 2713.545 1600.130 2718.890 1600.675 ;
        RECT 2695.605 1599.385 2696.125 1599.925 ;
        RECT 2698.570 1599.300 2698.910 1600.130 ;
        RECT 2704.090 1599.300 2704.430 1600.130 ;
        RECT 2709.610 1599.300 2709.950 1600.130 ;
        RECT 2715.130 1599.300 2715.470 1600.130 ;
        RECT 2719.065 1599.905 2720.735 1600.675 ;
        RECT 2721.365 1599.950 2721.655 1600.675 ;
        RECT 2721.825 1600.130 2727.170 1600.675 ;
        RECT 2727.345 1600.130 2732.690 1600.675 ;
        RECT 2719.065 1599.385 2719.815 1599.905 ;
        RECT 2723.410 1599.300 2723.750 1600.130 ;
        RECT 2728.930 1599.300 2729.270 1600.130 ;
        RECT 2732.865 1599.925 2734.075 1600.675 ;
        RECT 2733.555 1599.385 2734.075 1599.925 ;
        RECT 2695.605 1596.155 2696.125 1596.695 ;
        RECT 2695.605 1595.405 2696.815 1596.155 ;
        RECT 2699.950 1595.950 2700.290 1596.780 ;
        RECT 2703.885 1596.175 2705.535 1596.695 ;
        RECT 2697.425 1595.405 2697.755 1595.785 ;
        RECT 2698.365 1595.405 2703.710 1595.950 ;
        RECT 2703.885 1595.405 2707.395 1596.175 ;
        RECT 2708.485 1595.405 2708.775 1596.130 ;
        RECT 2710.530 1595.950 2710.870 1596.780 ;
        RECT 2716.050 1595.950 2716.390 1596.780 ;
        RECT 2721.570 1595.950 2721.910 1596.780 ;
        RECT 2727.090 1595.950 2727.430 1596.780 ;
        RECT 2731.025 1596.175 2731.775 1596.695 ;
        RECT 2708.945 1595.405 2714.290 1595.950 ;
        RECT 2714.465 1595.405 2719.810 1595.950 ;
        RECT 2719.985 1595.405 2725.330 1595.950 ;
        RECT 2725.505 1595.405 2730.850 1595.950 ;
        RECT 2731.025 1595.405 2732.695 1596.175 ;
        RECT 2733.555 1596.155 2734.075 1596.695 ;
        RECT 2732.865 1595.405 2734.075 1596.155 ;
        RECT 2695.520 1595.235 2734.160 1595.405 ;
        RECT 2695.605 1594.485 2696.815 1595.235 ;
        RECT 2696.985 1594.690 2702.330 1595.235 ;
        RECT 2702.505 1594.690 2707.850 1595.235 ;
        RECT 2708.025 1594.690 2713.370 1595.235 ;
        RECT 2713.545 1594.690 2718.890 1595.235 ;
        RECT 2695.605 1593.945 2696.125 1594.485 ;
        RECT 2698.570 1593.860 2698.910 1594.690 ;
        RECT 2704.090 1593.860 2704.430 1594.690 ;
        RECT 2709.610 1593.860 2709.950 1594.690 ;
        RECT 2715.130 1593.860 2715.470 1594.690 ;
        RECT 2719.065 1594.465 2720.735 1595.235 ;
        RECT 2721.365 1594.510 2721.655 1595.235 ;
        RECT 2721.825 1594.690 2727.170 1595.235 ;
        RECT 2727.345 1594.690 2732.690 1595.235 ;
        RECT 2719.065 1593.945 2719.815 1594.465 ;
        RECT 2723.410 1593.860 2723.750 1594.690 ;
        RECT 2728.930 1593.860 2729.270 1594.690 ;
        RECT 2732.865 1594.485 2734.075 1595.235 ;
        RECT 2733.555 1593.945 2734.075 1594.485 ;
        RECT 2695.605 1590.715 2696.125 1591.255 ;
        RECT 2695.605 1589.965 2696.815 1590.715 ;
        RECT 2701.330 1590.510 2701.670 1591.340 ;
        RECT 2705.265 1590.735 2706.475 1591.255 ;
        RECT 2697.425 1589.965 2697.755 1590.345 ;
        RECT 2698.805 1589.965 2699.135 1590.345 ;
        RECT 2699.745 1589.965 2705.090 1590.510 ;
        RECT 2705.265 1589.965 2707.855 1590.735 ;
        RECT 2708.485 1589.965 2708.775 1590.690 ;
        RECT 2710.530 1590.510 2710.870 1591.340 ;
        RECT 2716.050 1590.510 2716.390 1591.340 ;
        RECT 2719.985 1590.715 2720.505 1591.255 ;
        RECT 2708.945 1589.965 2714.290 1590.510 ;
        RECT 2714.465 1589.965 2719.810 1590.510 ;
        RECT 2719.985 1589.965 2721.195 1590.715 ;
        RECT 2721.365 1589.965 2721.655 1590.690 ;
        RECT 2723.410 1590.510 2723.750 1591.340 ;
        RECT 2728.930 1590.510 2729.270 1591.340 ;
        RECT 2733.555 1590.715 2734.075 1591.255 ;
        RECT 2721.825 1589.965 2727.170 1590.510 ;
        RECT 2727.345 1589.965 2732.690 1590.510 ;
        RECT 2732.865 1589.965 2734.075 1590.715 ;
        RECT 2695.520 1589.795 2734.160 1589.965 ;
        RECT 2523.330 1588.020 2523.670 1588.680 ;
        RECT 2522.130 1587.850 2523.935 1588.020 ;
        RECT 2523.330 1580.490 2523.670 1581.150 ;
        RECT 2522.130 1580.320 2523.935 1580.490 ;
        RECT 2523.330 1574.510 2523.670 1575.170 ;
        RECT 2522.130 1574.340 2523.935 1574.510 ;
        RECT 2523.330 1566.095 2523.670 1566.755 ;
        RECT 2522.130 1565.925 2523.935 1566.095 ;
        RECT 2343.000 1533.860 2442.425 1535.460 ;
        RECT 2358.215 1533.235 2358.385 1533.860 ;
        RECT 2366.795 1533.235 2366.965 1533.860 ;
        RECT 2367.750 1533.315 2367.920 1533.595 ;
        RECT 2367.750 1533.145 2367.980 1533.315 ;
        RECT 2372.410 1533.235 2372.580 1533.860 ;
        RECT 2375.155 1533.235 2375.325 1533.860 ;
        RECT 2376.150 1533.230 2376.320 1533.860 ;
        RECT 2383.120 1533.235 2383.290 1533.860 ;
        RECT 2384.075 1533.315 2384.245 1533.595 ;
        RECT 2384.075 1533.145 2384.305 1533.315 ;
        RECT 2388.735 1533.235 2388.905 1533.860 ;
        RECT 2391.480 1533.235 2391.650 1533.860 ;
        RECT 2392.475 1533.230 2392.645 1533.860 ;
        RECT 2399.445 1533.235 2399.615 1533.860 ;
        RECT 2400.400 1533.315 2400.570 1533.595 ;
        RECT 2400.400 1533.145 2400.630 1533.315 ;
        RECT 2405.060 1533.235 2405.230 1533.860 ;
        RECT 2407.805 1533.235 2407.975 1533.860 ;
        RECT 2408.800 1533.230 2408.970 1533.860 ;
        RECT 2415.770 1533.235 2415.940 1533.860 ;
        RECT 2416.725 1533.315 2416.895 1533.595 ;
        RECT 2416.725 1533.145 2416.955 1533.315 ;
        RECT 2421.385 1533.235 2421.555 1533.860 ;
        RECT 2424.130 1533.235 2424.300 1533.860 ;
        RECT 2425.125 1533.230 2425.295 1533.860 ;
        RECT 2432.095 1533.235 2432.265 1533.860 ;
        RECT 2433.050 1533.315 2433.220 1533.595 ;
        RECT 2433.050 1533.145 2433.280 1533.315 ;
        RECT 2437.710 1533.235 2437.880 1533.860 ;
        RECT 2440.455 1533.235 2440.625 1533.860 ;
        RECT 2441.450 1533.230 2441.620 1533.860 ;
        RECT 2367.810 1531.535 2367.980 1533.145 ;
        RECT 2384.135 1531.535 2384.305 1533.145 ;
        RECT 2400.460 1531.535 2400.630 1533.145 ;
        RECT 2416.785 1531.535 2416.955 1533.145 ;
        RECT 2433.110 1531.535 2433.280 1533.145 ;
        RECT 2367.750 1531.365 2367.980 1531.535 ;
        RECT 2384.075 1531.365 2384.305 1531.535 ;
        RECT 2400.400 1531.365 2400.630 1531.535 ;
        RECT 2416.725 1531.365 2416.955 1531.535 ;
        RECT 2433.050 1531.365 2433.280 1531.535 ;
        RECT 2367.750 1530.305 2367.920 1531.365 ;
        RECT 2384.075 1530.305 2384.245 1531.365 ;
        RECT 2400.400 1530.305 2400.570 1531.365 ;
        RECT 2416.725 1530.305 2416.895 1531.365 ;
        RECT 2433.050 1530.305 2433.220 1531.365 ;
        RECT 2368.665 1526.925 2368.835 1527.125 ;
        RECT 2370.625 1526.925 2370.795 1527.125 ;
        RECT 2384.990 1526.925 2385.160 1527.125 ;
        RECT 2386.950 1526.925 2387.120 1527.125 ;
        RECT 2401.315 1526.925 2401.485 1527.125 ;
        RECT 2403.275 1526.925 2403.445 1527.125 ;
        RECT 2417.640 1526.925 2417.810 1527.125 ;
        RECT 2419.600 1526.925 2419.770 1527.125 ;
        RECT 2433.965 1526.925 2434.135 1527.125 ;
        RECT 2435.925 1526.925 2436.095 1527.125 ;
        RECT 2368.345 1526.755 2368.835 1526.925 ;
        RECT 2370.305 1526.755 2370.795 1526.925 ;
        RECT 2384.670 1526.755 2385.160 1526.925 ;
        RECT 2386.630 1526.755 2387.120 1526.925 ;
        RECT 2400.995 1526.755 2401.485 1526.925 ;
        RECT 2402.955 1526.755 2403.445 1526.925 ;
        RECT 2417.320 1526.755 2417.810 1526.925 ;
        RECT 2419.280 1526.755 2419.770 1526.925 ;
        RECT 2433.645 1526.755 2434.135 1526.925 ;
        RECT 2435.605 1526.755 2436.095 1526.925 ;
        RECT 2361.865 1525.765 2362.035 1526.265 ;
        RECT 2362.825 1525.765 2362.995 1526.265 ;
        RECT 2363.785 1525.765 2363.955 1526.265 ;
        RECT 2364.305 1525.765 2364.475 1526.265 ;
        RECT 2365.265 1525.765 2365.435 1526.265 ;
        RECT 2367.705 1525.765 2367.875 1526.265 ;
        RECT 2369.665 1525.780 2369.835 1526.265 ;
        RECT 2369.485 1525.765 2369.835 1525.780 ;
        RECT 2378.190 1525.765 2378.360 1526.265 ;
        RECT 2379.150 1525.765 2379.320 1526.265 ;
        RECT 2380.110 1525.765 2380.280 1526.265 ;
        RECT 2380.630 1525.765 2380.800 1526.265 ;
        RECT 2381.590 1525.765 2381.760 1526.265 ;
        RECT 2384.030 1525.765 2384.200 1526.265 ;
        RECT 2385.990 1525.780 2386.160 1526.265 ;
        RECT 2385.810 1525.765 2386.160 1525.780 ;
        RECT 2394.515 1525.765 2394.685 1526.265 ;
        RECT 2395.475 1525.765 2395.645 1526.265 ;
        RECT 2396.435 1525.765 2396.605 1526.265 ;
        RECT 2396.955 1525.765 2397.125 1526.265 ;
        RECT 2397.915 1525.765 2398.085 1526.265 ;
        RECT 2400.355 1525.765 2400.525 1526.265 ;
        RECT 2402.315 1525.780 2402.485 1526.265 ;
        RECT 2402.135 1525.765 2402.485 1525.780 ;
        RECT 2410.840 1525.765 2411.010 1526.265 ;
        RECT 2411.800 1525.765 2411.970 1526.265 ;
        RECT 2412.760 1525.765 2412.930 1526.265 ;
        RECT 2413.280 1525.765 2413.450 1526.265 ;
        RECT 2414.240 1525.765 2414.410 1526.265 ;
        RECT 2416.680 1525.765 2416.850 1526.265 ;
        RECT 2418.640 1525.780 2418.810 1526.265 ;
        RECT 2418.460 1525.765 2418.810 1525.780 ;
        RECT 2427.165 1525.765 2427.335 1526.265 ;
        RECT 2428.125 1525.765 2428.295 1526.265 ;
        RECT 2429.085 1525.765 2429.255 1526.265 ;
        RECT 2429.605 1525.765 2429.775 1526.265 ;
        RECT 2430.565 1525.765 2430.735 1526.265 ;
        RECT 2433.005 1525.765 2433.175 1526.265 ;
        RECT 2434.965 1525.780 2435.135 1526.265 ;
        RECT 2434.785 1525.765 2435.135 1525.780 ;
        RECT 2361.535 1524.600 2371.350 1525.765 ;
        RECT 2372.410 1524.600 2372.580 1525.225 ;
        RECT 2375.155 1524.600 2375.325 1525.225 ;
        RECT 2376.145 1524.600 2376.315 1525.230 ;
        RECT 2377.860 1524.600 2387.675 1525.765 ;
        RECT 2388.735 1524.600 2388.905 1525.225 ;
        RECT 2391.480 1524.600 2391.650 1525.225 ;
        RECT 2392.470 1524.600 2392.640 1525.230 ;
        RECT 2394.185 1524.600 2404.000 1525.765 ;
        RECT 2405.060 1524.600 2405.230 1525.225 ;
        RECT 2407.805 1524.600 2407.975 1525.225 ;
        RECT 2408.795 1524.600 2408.965 1525.230 ;
        RECT 2410.510 1524.600 2420.325 1525.765 ;
        RECT 2421.385 1524.600 2421.555 1525.225 ;
        RECT 2424.130 1524.600 2424.300 1525.225 ;
        RECT 2425.120 1524.600 2425.290 1525.230 ;
        RECT 2426.835 1524.600 2436.650 1525.765 ;
        RECT 2437.710 1524.600 2437.880 1525.225 ;
        RECT 2440.455 1524.600 2440.625 1525.225 ;
        RECT 2441.445 1524.600 2441.615 1525.230 ;
        RECT 2343.000 1523.000 2442.420 1524.600 ;
        RECT 2695.520 1496.835 2734.160 1497.005 ;
        RECT 2695.605 1496.085 2696.815 1496.835 ;
        RECT 2697.455 1496.355 2697.730 1496.835 ;
        RECT 2698.315 1496.435 2698.650 1496.835 ;
        RECT 2699.265 1496.455 2699.595 1496.835 ;
        RECT 2700.645 1496.455 2700.975 1496.835 ;
        RECT 2701.585 1496.290 2706.930 1496.835 ;
        RECT 2695.605 1495.545 2696.125 1496.085 ;
        RECT 2703.170 1495.460 2703.510 1496.290 ;
        RECT 2707.105 1496.085 2708.315 1496.835 ;
        RECT 2708.485 1496.110 2708.775 1496.835 ;
        RECT 2709.420 1496.455 2709.750 1496.835 ;
        RECT 2707.105 1495.545 2707.625 1496.085 ;
        RECT 2710.350 1495.995 2710.610 1496.835 ;
        RECT 2710.785 1496.290 2716.130 1496.835 ;
        RECT 2712.370 1495.460 2712.710 1496.290 ;
        RECT 2716.305 1496.065 2719.815 1496.835 ;
        RECT 2719.985 1496.085 2721.195 1496.835 ;
        RECT 2721.365 1496.110 2721.655 1496.835 ;
        RECT 2721.830 1496.435 2722.165 1496.835 ;
        RECT 2722.750 1496.355 2723.025 1496.835 ;
        RECT 2723.665 1496.290 2729.010 1496.835 ;
        RECT 2716.305 1495.545 2717.955 1496.065 ;
        RECT 2719.985 1495.545 2720.505 1496.085 ;
        RECT 2725.250 1495.460 2725.590 1496.290 ;
        RECT 2729.185 1496.065 2730.855 1496.835 ;
        RECT 2731.925 1496.455 2732.255 1496.835 ;
        RECT 2732.865 1496.085 2734.075 1496.835 ;
        RECT 2729.185 1495.545 2729.935 1496.065 ;
        RECT 2733.555 1495.545 2734.075 1496.085 ;
        RECT 2695.605 1492.315 2696.125 1492.855 ;
        RECT 2695.605 1491.565 2696.815 1492.315 ;
        RECT 2699.950 1492.110 2700.290 1492.940 ;
        RECT 2703.885 1492.335 2705.535 1492.855 ;
        RECT 2697.425 1491.565 2697.755 1491.945 ;
        RECT 2698.365 1491.565 2703.710 1492.110 ;
        RECT 2703.885 1491.565 2707.395 1492.335 ;
        RECT 2708.485 1491.565 2708.775 1492.290 ;
        RECT 2710.530 1492.110 2710.870 1492.940 ;
        RECT 2716.050 1492.110 2716.390 1492.940 ;
        RECT 2721.570 1492.110 2721.910 1492.940 ;
        RECT 2727.090 1492.110 2727.430 1492.940 ;
        RECT 2731.025 1492.335 2731.775 1492.855 ;
        RECT 2708.945 1491.565 2714.290 1492.110 ;
        RECT 2714.465 1491.565 2719.810 1492.110 ;
        RECT 2719.985 1491.565 2725.330 1492.110 ;
        RECT 2725.505 1491.565 2730.850 1492.110 ;
        RECT 2731.025 1491.565 2732.695 1492.335 ;
        RECT 2733.555 1492.315 2734.075 1492.855 ;
        RECT 2732.865 1491.565 2734.075 1492.315 ;
        RECT 2695.520 1491.395 2734.160 1491.565 ;
        RECT 2695.605 1490.645 2696.815 1491.395 ;
        RECT 2696.985 1490.850 2702.330 1491.395 ;
        RECT 2702.505 1490.850 2707.850 1491.395 ;
        RECT 2708.025 1490.850 2713.370 1491.395 ;
        RECT 2713.545 1490.850 2718.890 1491.395 ;
        RECT 2695.605 1490.105 2696.125 1490.645 ;
        RECT 2698.570 1490.020 2698.910 1490.850 ;
        RECT 2704.090 1490.020 2704.430 1490.850 ;
        RECT 2709.610 1490.020 2709.950 1490.850 ;
        RECT 2715.130 1490.020 2715.470 1490.850 ;
        RECT 2719.065 1490.625 2720.735 1491.395 ;
        RECT 2721.365 1490.670 2721.655 1491.395 ;
        RECT 2721.825 1490.850 2727.170 1491.395 ;
        RECT 2727.345 1490.850 2732.690 1491.395 ;
        RECT 2719.065 1490.105 2719.815 1490.625 ;
        RECT 2723.410 1490.020 2723.750 1490.850 ;
        RECT 2728.930 1490.020 2729.270 1490.850 ;
        RECT 2732.865 1490.645 2734.075 1491.395 ;
        RECT 2733.555 1490.105 2734.075 1490.645 ;
        RECT 2695.605 1486.875 2696.125 1487.415 ;
        RECT 2695.605 1486.125 2696.815 1486.875 ;
        RECT 2698.570 1486.670 2698.910 1487.500 ;
        RECT 2704.090 1486.670 2704.430 1487.500 ;
        RECT 2696.985 1486.125 2702.330 1486.670 ;
        RECT 2702.505 1486.125 2707.850 1486.670 ;
        RECT 2708.485 1486.125 2708.775 1486.850 ;
        RECT 2710.530 1486.670 2710.870 1487.500 ;
        RECT 2716.050 1486.670 2716.390 1487.500 ;
        RECT 2721.570 1486.670 2721.910 1487.500 ;
        RECT 2727.090 1486.670 2727.430 1487.500 ;
        RECT 2731.025 1486.895 2731.775 1487.415 ;
        RECT 2708.945 1486.125 2714.290 1486.670 ;
        RECT 2714.465 1486.125 2719.810 1486.670 ;
        RECT 2719.985 1486.125 2725.330 1486.670 ;
        RECT 2725.505 1486.125 2730.850 1486.670 ;
        RECT 2731.025 1486.125 2732.695 1486.895 ;
        RECT 2733.555 1486.875 2734.075 1487.415 ;
        RECT 2732.865 1486.125 2734.075 1486.875 ;
        RECT 2695.520 1485.955 2734.160 1486.125 ;
        RECT 2695.605 1485.205 2696.815 1485.955 ;
        RECT 2697.425 1485.575 2697.755 1485.955 ;
        RECT 2698.365 1485.410 2703.710 1485.955 ;
        RECT 2703.885 1485.410 2709.230 1485.955 ;
        RECT 2709.405 1485.410 2714.750 1485.955 ;
        RECT 2714.925 1485.410 2720.270 1485.955 ;
        RECT 2695.605 1484.665 2696.125 1485.205 ;
        RECT 2699.950 1484.580 2700.290 1485.410 ;
        RECT 2705.470 1484.580 2705.810 1485.410 ;
        RECT 2710.990 1484.580 2711.330 1485.410 ;
        RECT 2716.510 1484.580 2716.850 1485.410 ;
        RECT 2721.365 1485.230 2721.655 1485.955 ;
        RECT 2721.825 1485.410 2727.170 1485.955 ;
        RECT 2727.345 1485.410 2732.690 1485.955 ;
        RECT 2723.410 1484.580 2723.750 1485.410 ;
        RECT 2728.930 1484.580 2729.270 1485.410 ;
        RECT 2732.865 1485.205 2734.075 1485.955 ;
        RECT 2733.555 1484.665 2734.075 1485.205 ;
        RECT 2695.605 1481.435 2696.125 1481.975 ;
        RECT 2695.605 1480.685 2696.815 1481.435 ;
        RECT 2698.570 1481.230 2698.910 1482.060 ;
        RECT 2704.090 1481.230 2704.430 1482.060 ;
        RECT 2696.985 1480.685 2702.330 1481.230 ;
        RECT 2702.505 1480.685 2707.850 1481.230 ;
        RECT 2708.485 1480.685 2708.775 1481.410 ;
        RECT 2710.530 1481.230 2710.870 1482.060 ;
        RECT 2716.050 1481.230 2716.390 1482.060 ;
        RECT 2721.570 1481.230 2721.910 1482.060 ;
        RECT 2727.090 1481.230 2727.430 1482.060 ;
        RECT 2731.025 1481.455 2731.775 1481.975 ;
        RECT 2708.945 1480.685 2714.290 1481.230 ;
        RECT 2714.465 1480.685 2719.810 1481.230 ;
        RECT 2719.985 1480.685 2725.330 1481.230 ;
        RECT 2725.505 1480.685 2730.850 1481.230 ;
        RECT 2731.025 1480.685 2732.695 1481.455 ;
        RECT 2733.555 1481.435 2734.075 1481.975 ;
        RECT 2732.865 1480.685 2734.075 1481.435 ;
        RECT 2695.520 1480.515 2734.160 1480.685 ;
        RECT 2695.605 1479.765 2696.815 1480.515 ;
        RECT 2697.415 1480.135 2697.745 1480.515 ;
        RECT 2699.700 1479.795 2699.990 1480.515 ;
        RECT 2702.050 1480.055 2702.220 1480.515 ;
        RECT 2702.910 1480.135 2703.240 1480.515 ;
        RECT 2705.795 1480.055 2705.965 1480.515 ;
        RECT 2706.645 1479.970 2711.990 1480.515 ;
        RECT 2712.165 1479.970 2717.510 1480.515 ;
        RECT 2695.605 1479.225 2696.125 1479.765 ;
        RECT 2708.230 1479.140 2708.570 1479.970 ;
        RECT 2713.750 1479.140 2714.090 1479.970 ;
        RECT 2717.685 1479.745 2721.195 1480.515 ;
        RECT 2721.365 1479.790 2721.655 1480.515 ;
        RECT 2721.825 1479.970 2727.170 1480.515 ;
        RECT 2727.345 1479.970 2732.690 1480.515 ;
        RECT 2717.685 1479.225 2719.335 1479.745 ;
        RECT 2723.410 1479.140 2723.750 1479.970 ;
        RECT 2728.930 1479.140 2729.270 1479.970 ;
        RECT 2732.865 1479.765 2734.075 1480.515 ;
        RECT 2733.555 1479.225 2734.075 1479.765 ;
        RECT 2695.605 1475.995 2696.125 1476.535 ;
        RECT 2695.605 1475.245 2696.815 1475.995 ;
        RECT 2699.950 1475.790 2700.290 1476.620 ;
        RECT 2703.885 1476.015 2705.535 1476.535 ;
        RECT 2697.425 1475.245 2697.755 1475.625 ;
        RECT 2698.365 1475.245 2703.710 1475.790 ;
        RECT 2703.885 1475.245 2707.395 1476.015 ;
        RECT 2708.485 1475.245 2708.775 1475.970 ;
        RECT 2710.530 1475.790 2710.870 1476.620 ;
        RECT 2716.050 1475.790 2716.390 1476.620 ;
        RECT 2721.570 1475.790 2721.910 1476.620 ;
        RECT 2727.090 1475.790 2727.430 1476.620 ;
        RECT 2731.025 1476.015 2731.775 1476.535 ;
        RECT 2708.945 1475.245 2714.290 1475.790 ;
        RECT 2714.465 1475.245 2719.810 1475.790 ;
        RECT 2719.985 1475.245 2725.330 1475.790 ;
        RECT 2725.505 1475.245 2730.850 1475.790 ;
        RECT 2731.025 1475.245 2732.695 1476.015 ;
        RECT 2733.555 1475.995 2734.075 1476.535 ;
        RECT 2732.865 1475.245 2734.075 1475.995 ;
        RECT 2695.520 1475.075 2734.160 1475.245 ;
        RECT 2695.605 1474.325 2696.815 1475.075 ;
        RECT 2697.415 1474.695 2697.745 1475.075 ;
        RECT 2699.700 1474.355 2699.990 1475.075 ;
        RECT 2702.050 1474.615 2702.220 1475.075 ;
        RECT 2702.910 1474.695 2703.240 1475.075 ;
        RECT 2705.795 1474.615 2705.965 1475.075 ;
        RECT 2706.645 1474.530 2711.990 1475.075 ;
        RECT 2712.165 1474.530 2717.510 1475.075 ;
        RECT 2695.605 1473.785 2696.125 1474.325 ;
        RECT 2708.230 1473.700 2708.570 1474.530 ;
        RECT 2713.750 1473.700 2714.090 1474.530 ;
        RECT 2717.685 1474.305 2721.195 1475.075 ;
        RECT 2721.365 1474.350 2721.655 1475.075 ;
        RECT 2721.825 1474.530 2727.170 1475.075 ;
        RECT 2727.345 1474.530 2732.690 1475.075 ;
        RECT 2717.685 1473.785 2719.335 1474.305 ;
        RECT 2723.410 1473.700 2723.750 1474.530 ;
        RECT 2728.930 1473.700 2729.270 1474.530 ;
        RECT 2732.865 1474.325 2734.075 1475.075 ;
        RECT 2733.555 1473.785 2734.075 1474.325 ;
        RECT 2695.605 1470.555 2696.125 1471.095 ;
        RECT 2698.365 1470.575 2699.575 1471.095 ;
        RECT 2705.725 1470.575 2706.935 1471.095 ;
        RECT 2695.605 1469.805 2696.815 1470.555 ;
        RECT 2697.425 1469.805 2697.755 1470.185 ;
        RECT 2698.365 1469.805 2700.955 1470.575 ;
        RECT 2702.015 1469.805 2702.345 1470.205 ;
        RECT 2704.305 1469.805 2704.815 1470.340 ;
        RECT 2705.725 1469.805 2708.315 1470.575 ;
        RECT 2708.485 1469.805 2708.775 1470.530 ;
        RECT 2710.530 1470.350 2710.870 1471.180 ;
        RECT 2716.050 1470.350 2716.390 1471.180 ;
        RECT 2721.570 1470.350 2721.910 1471.180 ;
        RECT 2727.090 1470.350 2727.430 1471.180 ;
        RECT 2731.025 1470.575 2731.775 1471.095 ;
        RECT 2708.945 1469.805 2714.290 1470.350 ;
        RECT 2714.465 1469.805 2719.810 1470.350 ;
        RECT 2719.985 1469.805 2725.330 1470.350 ;
        RECT 2725.505 1469.805 2730.850 1470.350 ;
        RECT 2731.025 1469.805 2732.695 1470.575 ;
        RECT 2733.555 1470.555 2734.075 1471.095 ;
        RECT 2732.865 1469.805 2734.075 1470.555 ;
        RECT 2695.520 1469.635 2734.160 1469.805 ;
        RECT 2695.605 1468.885 2696.815 1469.635 ;
        RECT 2696.985 1469.090 2702.330 1469.635 ;
        RECT 2702.505 1469.090 2707.850 1469.635 ;
        RECT 2708.025 1469.090 2713.370 1469.635 ;
        RECT 2713.545 1469.090 2718.890 1469.635 ;
        RECT 2695.605 1468.345 2696.125 1468.885 ;
        RECT 2698.570 1468.260 2698.910 1469.090 ;
        RECT 2704.090 1468.260 2704.430 1469.090 ;
        RECT 2709.610 1468.260 2709.950 1469.090 ;
        RECT 2715.130 1468.260 2715.470 1469.090 ;
        RECT 2719.065 1468.865 2720.735 1469.635 ;
        RECT 2721.365 1468.910 2721.655 1469.635 ;
        RECT 2721.825 1469.090 2727.170 1469.635 ;
        RECT 2727.345 1469.090 2732.690 1469.635 ;
        RECT 2719.065 1468.345 2719.815 1468.865 ;
        RECT 2723.410 1468.260 2723.750 1469.090 ;
        RECT 2728.930 1468.260 2729.270 1469.090 ;
        RECT 2732.865 1468.885 2734.075 1469.635 ;
        RECT 2733.555 1468.345 2734.075 1468.885 ;
        RECT 2695.605 1465.115 2696.125 1465.655 ;
        RECT 2695.605 1464.365 2696.815 1465.115 ;
        RECT 2699.950 1464.910 2700.290 1465.740 ;
        RECT 2703.885 1465.135 2705.535 1465.655 ;
        RECT 2697.425 1464.365 2697.755 1464.745 ;
        RECT 2698.365 1464.365 2703.710 1464.910 ;
        RECT 2703.885 1464.365 2707.395 1465.135 ;
        RECT 2708.485 1464.365 2708.775 1465.090 ;
        RECT 2710.530 1464.910 2710.870 1465.740 ;
        RECT 2716.050 1464.910 2716.390 1465.740 ;
        RECT 2721.570 1464.910 2721.910 1465.740 ;
        RECT 2727.090 1464.910 2727.430 1465.740 ;
        RECT 2731.025 1465.135 2731.775 1465.655 ;
        RECT 2708.945 1464.365 2714.290 1464.910 ;
        RECT 2714.465 1464.365 2719.810 1464.910 ;
        RECT 2719.985 1464.365 2725.330 1464.910 ;
        RECT 2725.505 1464.365 2730.850 1464.910 ;
        RECT 2731.025 1464.365 2732.695 1465.135 ;
        RECT 2733.555 1465.115 2734.075 1465.655 ;
        RECT 2732.865 1464.365 2734.075 1465.115 ;
        RECT 2695.520 1464.195 2734.160 1464.365 ;
        RECT 2695.605 1463.445 2696.815 1464.195 ;
        RECT 2696.985 1463.650 2702.330 1464.195 ;
        RECT 2702.505 1463.650 2707.850 1464.195 ;
        RECT 2708.025 1463.650 2713.370 1464.195 ;
        RECT 2713.545 1463.650 2718.890 1464.195 ;
        RECT 2695.605 1462.905 2696.125 1463.445 ;
        RECT 2698.570 1462.820 2698.910 1463.650 ;
        RECT 2704.090 1462.820 2704.430 1463.650 ;
        RECT 2709.610 1462.820 2709.950 1463.650 ;
        RECT 2715.130 1462.820 2715.470 1463.650 ;
        RECT 2719.065 1463.425 2720.735 1464.195 ;
        RECT 2721.365 1463.470 2721.655 1464.195 ;
        RECT 2721.825 1463.650 2727.170 1464.195 ;
        RECT 2727.345 1463.650 2732.690 1464.195 ;
        RECT 2719.065 1462.905 2719.815 1463.425 ;
        RECT 2723.410 1462.820 2723.750 1463.650 ;
        RECT 2728.930 1462.820 2729.270 1463.650 ;
        RECT 2732.865 1463.445 2734.075 1464.195 ;
        RECT 2733.555 1462.905 2734.075 1463.445 ;
        RECT 2695.605 1459.675 2696.125 1460.215 ;
        RECT 2696.985 1459.695 2698.635 1460.215 ;
        RECT 2695.605 1458.925 2696.815 1459.675 ;
        RECT 2696.985 1458.925 2700.495 1459.695 ;
        RECT 2701.605 1458.925 2701.845 1459.735 ;
        RECT 2702.515 1458.925 2702.785 1459.735 ;
        RECT 2704.550 1459.470 2704.890 1460.300 ;
        RECT 2702.965 1458.925 2708.310 1459.470 ;
        RECT 2708.485 1458.925 2708.775 1459.650 ;
        RECT 2710.530 1459.470 2710.870 1460.300 ;
        RECT 2716.050 1459.470 2716.390 1460.300 ;
        RECT 2721.570 1459.470 2721.910 1460.300 ;
        RECT 2727.090 1459.470 2727.430 1460.300 ;
        RECT 2731.025 1459.695 2731.775 1460.215 ;
        RECT 2708.945 1458.925 2714.290 1459.470 ;
        RECT 2714.465 1458.925 2719.810 1459.470 ;
        RECT 2719.985 1458.925 2725.330 1459.470 ;
        RECT 2725.505 1458.925 2730.850 1459.470 ;
        RECT 2731.025 1458.925 2732.695 1459.695 ;
        RECT 2733.555 1459.675 2734.075 1460.215 ;
        RECT 2732.865 1458.925 2734.075 1459.675 ;
        RECT 2695.520 1458.755 2734.160 1458.925 ;
        RECT 2695.605 1458.005 2696.815 1458.755 ;
        RECT 2697.425 1458.375 2697.755 1458.755 ;
        RECT 2695.605 1457.465 2696.125 1458.005 ;
        RECT 2698.365 1457.985 2701.875 1458.755 ;
        RECT 2702.055 1458.015 2702.385 1458.755 ;
        RECT 2703.090 1458.395 2703.420 1458.755 ;
        RECT 2698.365 1457.465 2700.015 1457.985 ;
        RECT 2704.785 1457.975 2705.080 1458.755 ;
        RECT 2705.265 1458.210 2710.610 1458.755 ;
        RECT 2710.785 1458.210 2716.130 1458.755 ;
        RECT 2706.850 1457.380 2707.190 1458.210 ;
        RECT 2712.370 1457.380 2712.710 1458.210 ;
        RECT 2716.305 1457.985 2719.815 1458.755 ;
        RECT 2719.985 1458.005 2721.195 1458.755 ;
        RECT 2721.365 1458.030 2721.655 1458.755 ;
        RECT 2721.825 1458.210 2727.170 1458.755 ;
        RECT 2727.345 1458.210 2732.690 1458.755 ;
        RECT 2716.305 1457.465 2717.955 1457.985 ;
        RECT 2719.985 1457.465 2720.505 1458.005 ;
        RECT 2723.410 1457.380 2723.750 1458.210 ;
        RECT 2728.930 1457.380 2729.270 1458.210 ;
        RECT 2732.865 1458.005 2734.075 1458.755 ;
        RECT 2733.555 1457.465 2734.075 1458.005 ;
        RECT 2695.605 1454.235 2696.125 1454.775 ;
        RECT 2695.605 1453.485 2696.815 1454.235 ;
        RECT 2698.570 1454.030 2698.910 1454.860 ;
        RECT 2704.090 1454.030 2704.430 1454.860 ;
        RECT 2696.985 1453.485 2702.330 1454.030 ;
        RECT 2702.505 1453.485 2707.850 1454.030 ;
        RECT 2708.485 1453.485 2708.775 1454.210 ;
        RECT 2710.530 1454.030 2710.870 1454.860 ;
        RECT 2716.050 1454.030 2716.390 1454.860 ;
        RECT 2721.570 1454.030 2721.910 1454.860 ;
        RECT 2708.945 1453.485 2714.290 1454.030 ;
        RECT 2714.465 1453.485 2719.810 1454.030 ;
        RECT 2719.985 1453.485 2725.330 1454.030 ;
        RECT 2725.515 1453.485 2725.845 1453.965 ;
        RECT 2726.355 1453.485 2726.685 1453.965 ;
        RECT 2727.195 1453.485 2727.525 1453.965 ;
        RECT 2728.035 1453.485 2728.365 1453.965 ;
        RECT 2728.875 1453.485 2729.205 1453.965 ;
        RECT 2729.715 1453.485 2730.045 1453.965 ;
        RECT 2730.555 1453.485 2730.885 1453.965 ;
        RECT 2731.395 1453.485 2731.725 1453.965 ;
        RECT 2732.235 1453.485 2732.565 1454.285 ;
        RECT 2733.555 1454.235 2734.075 1454.775 ;
        RECT 2732.865 1453.485 2734.075 1454.235 ;
        RECT 2695.520 1453.315 2734.160 1453.485 ;
        RECT 2695.605 1452.565 2696.815 1453.315 ;
        RECT 2697.425 1452.935 2697.755 1453.315 ;
        RECT 2698.365 1452.770 2703.710 1453.315 ;
        RECT 2703.885 1452.770 2709.230 1453.315 ;
        RECT 2709.405 1452.770 2714.750 1453.315 ;
        RECT 2714.925 1452.770 2720.270 1453.315 ;
        RECT 2695.605 1452.025 2696.125 1452.565 ;
        RECT 2699.950 1451.940 2700.290 1452.770 ;
        RECT 2705.470 1451.940 2705.810 1452.770 ;
        RECT 2710.990 1451.940 2711.330 1452.770 ;
        RECT 2716.510 1451.940 2716.850 1452.770 ;
        RECT 2721.365 1452.590 2721.655 1453.315 ;
        RECT 2721.825 1452.770 2727.170 1453.315 ;
        RECT 2727.345 1452.770 2732.690 1453.315 ;
        RECT 2723.410 1451.940 2723.750 1452.770 ;
        RECT 2728.930 1451.940 2729.270 1452.770 ;
        RECT 2732.865 1452.565 2734.075 1453.315 ;
        RECT 2733.555 1452.025 2734.075 1452.565 ;
        RECT 2695.605 1448.795 2696.125 1449.335 ;
        RECT 2695.605 1448.045 2696.815 1448.795 ;
        RECT 2698.570 1448.590 2698.910 1449.420 ;
        RECT 2704.090 1448.590 2704.430 1449.420 ;
        RECT 2696.985 1448.045 2702.330 1448.590 ;
        RECT 2702.505 1448.045 2707.850 1448.590 ;
        RECT 2708.485 1448.045 2708.775 1448.770 ;
        RECT 2710.530 1448.590 2710.870 1449.420 ;
        RECT 2716.050 1448.590 2716.390 1449.420 ;
        RECT 2721.570 1448.590 2721.910 1449.420 ;
        RECT 2727.090 1448.590 2727.430 1449.420 ;
        RECT 2731.025 1448.815 2731.775 1449.335 ;
        RECT 2708.945 1448.045 2714.290 1448.590 ;
        RECT 2714.465 1448.045 2719.810 1448.590 ;
        RECT 2719.985 1448.045 2725.330 1448.590 ;
        RECT 2725.505 1448.045 2730.850 1448.590 ;
        RECT 2731.025 1448.045 2732.695 1448.815 ;
        RECT 2733.555 1448.795 2734.075 1449.335 ;
        RECT 2732.865 1448.045 2734.075 1448.795 ;
        RECT 2695.520 1447.875 2734.160 1448.045 ;
        RECT 2695.605 1447.125 2696.815 1447.875 ;
        RECT 2697.715 1447.135 2698.045 1447.875 ;
        RECT 2698.555 1447.475 2698.885 1447.875 ;
        RECT 2699.745 1447.330 2705.090 1447.875 ;
        RECT 2705.265 1447.330 2710.610 1447.875 ;
        RECT 2710.785 1447.330 2716.130 1447.875 ;
        RECT 2695.605 1446.585 2696.125 1447.125 ;
        RECT 2701.330 1446.500 2701.670 1447.330 ;
        RECT 2706.850 1446.500 2707.190 1447.330 ;
        RECT 2712.370 1446.500 2712.710 1447.330 ;
        RECT 2716.305 1447.105 2719.815 1447.875 ;
        RECT 2719.985 1447.125 2721.195 1447.875 ;
        RECT 2721.365 1447.150 2721.655 1447.875 ;
        RECT 2721.825 1447.330 2727.170 1447.875 ;
        RECT 2727.345 1447.330 2732.690 1447.875 ;
        RECT 2716.305 1446.585 2717.955 1447.105 ;
        RECT 2719.985 1446.585 2720.505 1447.125 ;
        RECT 2723.410 1446.500 2723.750 1447.330 ;
        RECT 2728.930 1446.500 2729.270 1447.330 ;
        RECT 2732.865 1447.125 2734.075 1447.875 ;
        RECT 2733.555 1446.585 2734.075 1447.125 ;
        RECT 2695.605 1443.355 2696.125 1443.895 ;
        RECT 2695.605 1442.605 2696.815 1443.355 ;
        RECT 2699.950 1443.150 2700.290 1443.980 ;
        RECT 2703.885 1443.375 2705.535 1443.895 ;
        RECT 2697.425 1442.605 2697.755 1442.985 ;
        RECT 2698.365 1442.605 2703.710 1443.150 ;
        RECT 2703.885 1442.605 2707.395 1443.375 ;
        RECT 2708.485 1442.605 2708.775 1443.330 ;
        RECT 2710.530 1443.150 2710.870 1443.980 ;
        RECT 2716.050 1443.150 2716.390 1443.980 ;
        RECT 2721.570 1443.150 2721.910 1443.980 ;
        RECT 2727.090 1443.150 2727.430 1443.980 ;
        RECT 2731.025 1443.375 2731.775 1443.895 ;
        RECT 2708.945 1442.605 2714.290 1443.150 ;
        RECT 2714.465 1442.605 2719.810 1443.150 ;
        RECT 2719.985 1442.605 2725.330 1443.150 ;
        RECT 2725.505 1442.605 2730.850 1443.150 ;
        RECT 2731.025 1442.605 2732.695 1443.375 ;
        RECT 2733.555 1443.355 2734.075 1443.895 ;
        RECT 2732.865 1442.605 2734.075 1443.355 ;
        RECT 2695.520 1442.435 2734.160 1442.605 ;
        RECT 2695.605 1441.685 2696.815 1442.435 ;
        RECT 2697.725 1441.900 2698.235 1442.435 ;
        RECT 2700.195 1442.035 2700.525 1442.435 ;
        RECT 2701.210 1441.760 2701.450 1442.435 ;
        RECT 2702.840 1441.985 2703.170 1442.435 ;
        RECT 2704.090 1441.995 2704.405 1442.435 ;
        RECT 2704.805 1441.890 2710.150 1442.435 ;
        RECT 2710.325 1441.890 2715.670 1442.435 ;
        RECT 2715.845 1441.890 2721.190 1442.435 ;
        RECT 2695.605 1441.145 2696.125 1441.685 ;
        RECT 2706.390 1441.060 2706.730 1441.890 ;
        RECT 2711.910 1441.060 2712.250 1441.890 ;
        RECT 2717.430 1441.060 2717.770 1441.890 ;
        RECT 2721.365 1441.710 2721.655 1442.435 ;
        RECT 2721.825 1441.890 2727.170 1442.435 ;
        RECT 2727.345 1441.890 2732.690 1442.435 ;
        RECT 2723.410 1441.060 2723.750 1441.890 ;
        RECT 2728.930 1441.060 2729.270 1441.890 ;
        RECT 2732.865 1441.685 2734.075 1442.435 ;
        RECT 2733.555 1441.145 2734.075 1441.685 ;
        RECT 2695.605 1437.915 2696.125 1438.455 ;
        RECT 2343.000 1435.865 2453.600 1437.465 ;
        RECT 2695.605 1437.165 2696.815 1437.915 ;
        RECT 2696.985 1437.165 2697.245 1437.985 ;
        RECT 2701.790 1437.710 2702.130 1438.540 ;
        RECT 2705.725 1437.935 2706.935 1438.455 ;
        RECT 2699.275 1437.165 2699.605 1437.625 ;
        RECT 2700.205 1437.165 2705.550 1437.710 ;
        RECT 2705.725 1437.165 2708.315 1437.935 ;
        RECT 2708.485 1437.165 2708.775 1437.890 ;
        RECT 2710.530 1437.710 2710.870 1438.540 ;
        RECT 2716.050 1437.710 2716.390 1438.540 ;
        RECT 2721.570 1437.710 2721.910 1438.540 ;
        RECT 2727.090 1437.710 2727.430 1438.540 ;
        RECT 2731.025 1437.935 2731.775 1438.455 ;
        RECT 2708.945 1437.165 2714.290 1437.710 ;
        RECT 2714.465 1437.165 2719.810 1437.710 ;
        RECT 2719.985 1437.165 2725.330 1437.710 ;
        RECT 2725.505 1437.165 2730.850 1437.710 ;
        RECT 2731.025 1437.165 2732.695 1437.935 ;
        RECT 2733.555 1437.915 2734.075 1438.455 ;
        RECT 2732.865 1437.165 2734.075 1437.915 ;
        RECT 2523.330 1436.395 2523.670 1437.055 ;
        RECT 2695.520 1436.995 2734.160 1437.165 ;
        RECT 2522.130 1436.225 2523.935 1436.395 ;
        RECT 2695.605 1436.245 2696.815 1436.995 ;
        RECT 2697.425 1436.615 2697.755 1436.995 ;
        RECT 2698.365 1436.450 2703.710 1436.995 ;
        RECT 2703.885 1436.450 2709.230 1436.995 ;
        RECT 2709.405 1436.450 2714.750 1436.995 ;
        RECT 2714.925 1436.450 2720.270 1436.995 ;
        RECT 2358.215 1435.240 2358.385 1435.865 ;
        RECT 2369.030 1435.240 2369.200 1435.865 ;
        RECT 2369.985 1435.320 2370.155 1435.600 ;
        RECT 2369.985 1435.150 2370.215 1435.320 ;
        RECT 2374.645 1435.240 2374.815 1435.865 ;
        RECT 2377.390 1435.240 2377.560 1435.865 ;
        RECT 2378.385 1435.235 2378.555 1435.865 ;
        RECT 2387.590 1435.240 2387.760 1435.865 ;
        RECT 2388.545 1435.320 2388.715 1435.600 ;
        RECT 2388.545 1435.150 2388.775 1435.320 ;
        RECT 2393.205 1435.240 2393.375 1435.865 ;
        RECT 2395.950 1435.240 2396.120 1435.865 ;
        RECT 2396.945 1435.235 2397.115 1435.865 ;
        RECT 2406.150 1435.240 2406.320 1435.865 ;
        RECT 2407.105 1435.320 2407.275 1435.600 ;
        RECT 2407.105 1435.150 2407.335 1435.320 ;
        RECT 2411.765 1435.240 2411.935 1435.865 ;
        RECT 2414.510 1435.240 2414.680 1435.865 ;
        RECT 2415.505 1435.235 2415.675 1435.865 ;
        RECT 2424.710 1435.240 2424.880 1435.865 ;
        RECT 2425.665 1435.320 2425.835 1435.600 ;
        RECT 2425.665 1435.150 2425.895 1435.320 ;
        RECT 2430.325 1435.240 2430.495 1435.865 ;
        RECT 2433.070 1435.240 2433.240 1435.865 ;
        RECT 2434.065 1435.235 2434.235 1435.865 ;
        RECT 2443.270 1435.240 2443.440 1435.865 ;
        RECT 2444.225 1435.320 2444.395 1435.600 ;
        RECT 2444.225 1435.150 2444.455 1435.320 ;
        RECT 2448.885 1435.240 2449.055 1435.865 ;
        RECT 2451.630 1435.240 2451.800 1435.865 ;
        RECT 2452.625 1435.235 2452.795 1435.865 ;
        RECT 2695.605 1435.705 2696.125 1436.245 ;
        RECT 2699.950 1435.620 2700.290 1436.450 ;
        RECT 2705.470 1435.620 2705.810 1436.450 ;
        RECT 2710.990 1435.620 2711.330 1436.450 ;
        RECT 2716.510 1435.620 2716.850 1436.450 ;
        RECT 2721.365 1436.270 2721.655 1436.995 ;
        RECT 2721.825 1436.450 2727.170 1436.995 ;
        RECT 2727.345 1436.450 2732.690 1436.995 ;
        RECT 2723.410 1435.620 2723.750 1436.450 ;
        RECT 2728.930 1435.620 2729.270 1436.450 ;
        RECT 2732.865 1436.245 2734.075 1436.995 ;
        RECT 2733.555 1435.705 2734.075 1436.245 ;
        RECT 2370.045 1433.540 2370.215 1435.150 ;
        RECT 2388.605 1433.540 2388.775 1435.150 ;
        RECT 2407.165 1433.540 2407.335 1435.150 ;
        RECT 2425.725 1433.540 2425.895 1435.150 ;
        RECT 2444.285 1433.540 2444.455 1435.150 ;
        RECT 2369.985 1433.370 2370.215 1433.540 ;
        RECT 2388.545 1433.370 2388.775 1433.540 ;
        RECT 2407.105 1433.370 2407.335 1433.540 ;
        RECT 2425.665 1433.370 2425.895 1433.540 ;
        RECT 2444.225 1433.370 2444.455 1433.540 ;
        RECT 2369.985 1432.310 2370.155 1433.370 ;
        RECT 2388.545 1432.310 2388.715 1433.370 ;
        RECT 2407.105 1432.310 2407.275 1433.370 ;
        RECT 2425.665 1432.310 2425.835 1433.370 ;
        RECT 2444.225 1432.310 2444.395 1433.370 ;
        RECT 2695.605 1432.475 2696.125 1433.015 ;
        RECT 2696.985 1432.475 2697.505 1433.015 ;
        RECT 2695.605 1431.725 2696.815 1432.475 ;
        RECT 2696.985 1431.725 2698.195 1432.475 ;
        RECT 2698.365 1431.725 2698.705 1432.450 ;
        RECT 2703.630 1432.270 2703.970 1433.100 ;
        RECT 2701.035 1431.725 2701.365 1432.205 ;
        RECT 2702.045 1431.725 2707.390 1432.270 ;
        RECT 2708.485 1431.725 2708.775 1432.450 ;
        RECT 2710.530 1432.270 2710.870 1433.100 ;
        RECT 2716.050 1432.270 2716.390 1433.100 ;
        RECT 2721.570 1432.270 2721.910 1433.100 ;
        RECT 2727.090 1432.270 2727.430 1433.100 ;
        RECT 2731.025 1432.495 2731.775 1433.015 ;
        RECT 2708.945 1431.725 2714.290 1432.270 ;
        RECT 2714.465 1431.725 2719.810 1432.270 ;
        RECT 2719.985 1431.725 2725.330 1432.270 ;
        RECT 2725.505 1431.725 2730.850 1432.270 ;
        RECT 2731.025 1431.725 2732.695 1432.495 ;
        RECT 2733.555 1432.475 2734.075 1433.015 ;
        RECT 2732.865 1431.725 2734.075 1432.475 ;
        RECT 2695.520 1431.555 2734.160 1431.725 ;
        RECT 2695.605 1430.805 2696.815 1431.555 ;
        RECT 2523.330 1429.980 2523.670 1430.640 ;
        RECT 2695.605 1430.265 2696.125 1430.805 ;
        RECT 2697.905 1430.735 2698.165 1431.555 ;
        RECT 2699.275 1431.155 2699.605 1431.555 ;
        RECT 2700.115 1431.155 2700.490 1431.555 ;
        RECT 2702.760 1431.155 2703.090 1431.555 ;
        RECT 2703.885 1431.010 2709.230 1431.555 ;
        RECT 2709.405 1431.010 2714.750 1431.555 ;
        RECT 2714.925 1431.010 2720.270 1431.555 ;
        RECT 2705.470 1430.180 2705.810 1431.010 ;
        RECT 2710.990 1430.180 2711.330 1431.010 ;
        RECT 2716.510 1430.180 2716.850 1431.010 ;
        RECT 2721.365 1430.830 2721.655 1431.555 ;
        RECT 2721.825 1431.010 2727.170 1431.555 ;
        RECT 2727.345 1431.010 2732.690 1431.555 ;
        RECT 2723.410 1430.180 2723.750 1431.010 ;
        RECT 2728.930 1430.180 2729.270 1431.010 ;
        RECT 2732.865 1430.805 2734.075 1431.555 ;
        RECT 2733.555 1430.265 2734.075 1430.805 ;
        RECT 2522.130 1429.810 2523.935 1429.980 ;
        RECT 2363.190 1429.345 2363.480 1429.515 ;
        RECT 2381.750 1429.345 2382.040 1429.515 ;
        RECT 2400.310 1429.345 2400.600 1429.515 ;
        RECT 2418.870 1429.345 2419.160 1429.515 ;
        RECT 2437.430 1429.345 2437.720 1429.515 ;
        RECT 2363.190 1429.035 2363.360 1429.345 ;
        RECT 2362.990 1428.865 2363.360 1429.035 ;
        RECT 2365.030 1428.785 2365.200 1429.115 ;
        RECT 2381.750 1429.035 2381.920 1429.345 ;
        RECT 2381.550 1428.865 2381.920 1429.035 ;
        RECT 2383.590 1428.785 2383.760 1429.115 ;
        RECT 2400.310 1429.035 2400.480 1429.345 ;
        RECT 2400.110 1428.865 2400.480 1429.035 ;
        RECT 2402.150 1428.785 2402.320 1429.115 ;
        RECT 2418.870 1429.035 2419.040 1429.345 ;
        RECT 2418.670 1428.865 2419.040 1429.035 ;
        RECT 2420.710 1428.785 2420.880 1429.115 ;
        RECT 2437.430 1429.035 2437.600 1429.345 ;
        RECT 2437.230 1428.865 2437.600 1429.035 ;
        RECT 2439.270 1428.785 2439.440 1429.115 ;
        RECT 2362.350 1427.875 2362.520 1428.375 ;
        RECT 2363.830 1427.890 2364.000 1428.375 ;
        RECT 2363.830 1427.875 2364.090 1427.890 ;
        RECT 2365.750 1427.875 2365.920 1428.375 ;
        RECT 2366.195 1427.875 2366.390 1427.890 ;
        RECT 2367.230 1427.875 2367.400 1428.375 ;
        RECT 2368.190 1427.875 2368.360 1428.375 ;
        RECT 2369.190 1427.875 2369.360 1428.375 ;
        RECT 2370.150 1427.875 2370.320 1428.375 ;
        RECT 2370.670 1427.875 2370.840 1428.375 ;
        RECT 2371.630 1427.875 2371.800 1428.375 ;
        RECT 2372.590 1427.875 2372.760 1428.375 ;
        RECT 2373.395 1427.875 2373.585 1427.880 ;
        RECT 2380.910 1427.875 2381.080 1428.375 ;
        RECT 2382.390 1427.890 2382.560 1428.375 ;
        RECT 2382.390 1427.875 2382.650 1427.890 ;
        RECT 2384.310 1427.875 2384.480 1428.375 ;
        RECT 2384.755 1427.875 2384.950 1427.890 ;
        RECT 2385.790 1427.875 2385.960 1428.375 ;
        RECT 2386.750 1427.875 2386.920 1428.375 ;
        RECT 2387.750 1427.875 2387.920 1428.375 ;
        RECT 2388.710 1427.875 2388.880 1428.375 ;
        RECT 2389.230 1427.875 2389.400 1428.375 ;
        RECT 2390.190 1427.875 2390.360 1428.375 ;
        RECT 2391.150 1427.875 2391.320 1428.375 ;
        RECT 2391.955 1427.875 2392.145 1427.880 ;
        RECT 2399.470 1427.875 2399.640 1428.375 ;
        RECT 2400.950 1427.890 2401.120 1428.375 ;
        RECT 2400.950 1427.875 2401.210 1427.890 ;
        RECT 2402.870 1427.875 2403.040 1428.375 ;
        RECT 2403.315 1427.875 2403.510 1427.890 ;
        RECT 2404.350 1427.875 2404.520 1428.375 ;
        RECT 2405.310 1427.875 2405.480 1428.375 ;
        RECT 2406.310 1427.875 2406.480 1428.375 ;
        RECT 2407.270 1427.875 2407.440 1428.375 ;
        RECT 2407.790 1427.875 2407.960 1428.375 ;
        RECT 2408.750 1427.875 2408.920 1428.375 ;
        RECT 2409.710 1427.875 2409.880 1428.375 ;
        RECT 2410.515 1427.875 2410.705 1427.880 ;
        RECT 2418.030 1427.875 2418.200 1428.375 ;
        RECT 2419.510 1427.890 2419.680 1428.375 ;
        RECT 2419.510 1427.875 2419.770 1427.890 ;
        RECT 2421.430 1427.875 2421.600 1428.375 ;
        RECT 2421.875 1427.875 2422.070 1427.890 ;
        RECT 2422.910 1427.875 2423.080 1428.375 ;
        RECT 2423.870 1427.875 2424.040 1428.375 ;
        RECT 2424.870 1427.875 2425.040 1428.375 ;
        RECT 2425.830 1427.875 2426.000 1428.375 ;
        RECT 2426.350 1427.875 2426.520 1428.375 ;
        RECT 2427.310 1427.875 2427.480 1428.375 ;
        RECT 2428.270 1427.875 2428.440 1428.375 ;
        RECT 2429.075 1427.875 2429.265 1427.880 ;
        RECT 2436.590 1427.875 2436.760 1428.375 ;
        RECT 2438.070 1427.890 2438.240 1428.375 ;
        RECT 2438.070 1427.875 2438.330 1427.890 ;
        RECT 2439.990 1427.875 2440.160 1428.375 ;
        RECT 2440.435 1427.875 2440.630 1427.890 ;
        RECT 2441.470 1427.875 2441.640 1428.375 ;
        RECT 2442.430 1427.875 2442.600 1428.375 ;
        RECT 2443.430 1427.875 2443.600 1428.375 ;
        RECT 2444.390 1427.875 2444.560 1428.375 ;
        RECT 2444.910 1427.875 2445.080 1428.375 ;
        RECT 2445.870 1427.875 2446.040 1428.375 ;
        RECT 2446.830 1427.875 2447.000 1428.375 ;
        RECT 2447.635 1427.875 2447.825 1427.880 ;
        RECT 2361.540 1426.600 2373.585 1427.875 ;
        RECT 2374.645 1426.600 2374.815 1427.225 ;
        RECT 2377.390 1426.600 2377.560 1427.225 ;
        RECT 2378.380 1426.600 2378.550 1427.230 ;
        RECT 2380.100 1426.600 2392.145 1427.875 ;
        RECT 2393.205 1426.600 2393.375 1427.225 ;
        RECT 2395.950 1426.600 2396.120 1427.225 ;
        RECT 2396.940 1426.600 2397.110 1427.230 ;
        RECT 2398.660 1426.600 2410.705 1427.875 ;
        RECT 2411.765 1426.600 2411.935 1427.225 ;
        RECT 2414.510 1426.600 2414.680 1427.225 ;
        RECT 2415.500 1426.600 2415.670 1427.230 ;
        RECT 2417.220 1426.600 2429.265 1427.875 ;
        RECT 2430.325 1426.600 2430.495 1427.225 ;
        RECT 2433.070 1426.600 2433.240 1427.225 ;
        RECT 2434.060 1426.600 2434.230 1427.230 ;
        RECT 2435.780 1426.600 2447.825 1427.875 ;
        RECT 2448.885 1426.600 2449.055 1427.225 ;
        RECT 2451.630 1426.600 2451.800 1427.225 ;
        RECT 2452.620 1426.600 2452.790 1427.230 ;
        RECT 2695.605 1427.035 2696.125 1427.575 ;
        RECT 2343.000 1425.000 2453.595 1426.600 ;
        RECT 2695.605 1426.285 2696.815 1427.035 ;
        RECT 2697.425 1426.285 2697.755 1426.665 ;
        RECT 2699.725 1426.285 2700.035 1427.085 ;
        RECT 2701.790 1426.830 2702.130 1427.660 ;
        RECT 2705.725 1427.055 2706.935 1427.575 ;
        RECT 2700.205 1426.285 2705.550 1426.830 ;
        RECT 2705.725 1426.285 2708.315 1427.055 ;
        RECT 2708.485 1426.285 2708.775 1427.010 ;
        RECT 2710.530 1426.830 2710.870 1427.660 ;
        RECT 2716.050 1426.830 2716.390 1427.660 ;
        RECT 2721.570 1426.830 2721.910 1427.660 ;
        RECT 2727.090 1426.830 2727.430 1427.660 ;
        RECT 2731.025 1427.055 2731.775 1427.575 ;
        RECT 2708.945 1426.285 2714.290 1426.830 ;
        RECT 2714.465 1426.285 2719.810 1426.830 ;
        RECT 2719.985 1426.285 2725.330 1426.830 ;
        RECT 2725.505 1426.285 2730.850 1426.830 ;
        RECT 2731.025 1426.285 2732.695 1427.055 ;
        RECT 2733.555 1427.035 2734.075 1427.575 ;
        RECT 2732.865 1426.285 2734.075 1427.035 ;
        RECT 2695.520 1426.115 2734.160 1426.285 ;
        RECT 2695.605 1425.365 2696.815 1426.115 ;
        RECT 2697.725 1425.580 2698.235 1426.115 ;
        RECT 2700.195 1425.715 2700.525 1426.115 ;
        RECT 2701.125 1425.570 2706.470 1426.115 ;
        RECT 2706.645 1425.570 2711.990 1426.115 ;
        RECT 2712.165 1425.570 2717.510 1426.115 ;
        RECT 2695.605 1424.825 2696.125 1425.365 ;
        RECT 2702.710 1424.740 2703.050 1425.570 ;
        RECT 2708.230 1424.740 2708.570 1425.570 ;
        RECT 2713.750 1424.740 2714.090 1425.570 ;
        RECT 2717.685 1425.345 2721.195 1426.115 ;
        RECT 2721.365 1425.390 2721.655 1426.115 ;
        RECT 2721.825 1425.570 2727.170 1426.115 ;
        RECT 2727.345 1425.570 2732.690 1426.115 ;
        RECT 2717.685 1424.825 2719.335 1425.345 ;
        RECT 2723.410 1424.740 2723.750 1425.570 ;
        RECT 2728.930 1424.740 2729.270 1425.570 ;
        RECT 2732.865 1425.365 2734.075 1426.115 ;
        RECT 2733.555 1424.825 2734.075 1425.365 ;
        RECT 2695.605 1421.595 2696.125 1422.135 ;
        RECT 2695.605 1420.845 2696.815 1421.595 ;
        RECT 2699.950 1421.390 2700.290 1422.220 ;
        RECT 2703.885 1421.615 2705.535 1422.135 ;
        RECT 2697.425 1420.845 2697.755 1421.225 ;
        RECT 2698.365 1420.845 2703.710 1421.390 ;
        RECT 2703.885 1420.845 2707.395 1421.615 ;
        RECT 2708.485 1420.845 2708.775 1421.570 ;
        RECT 2710.530 1421.390 2710.870 1422.220 ;
        RECT 2716.050 1421.390 2716.390 1422.220 ;
        RECT 2721.570 1421.390 2721.910 1422.220 ;
        RECT 2727.090 1421.390 2727.430 1422.220 ;
        RECT 2731.025 1421.615 2731.775 1422.135 ;
        RECT 2708.945 1420.845 2714.290 1421.390 ;
        RECT 2714.465 1420.845 2719.810 1421.390 ;
        RECT 2719.985 1420.845 2725.330 1421.390 ;
        RECT 2725.505 1420.845 2730.850 1421.390 ;
        RECT 2731.025 1420.845 2732.695 1421.615 ;
        RECT 2733.555 1421.595 2734.075 1422.135 ;
        RECT 2732.865 1420.845 2734.075 1421.595 ;
        RECT 2695.520 1420.675 2734.160 1420.845 ;
        RECT 2695.605 1419.925 2696.815 1420.675 ;
        RECT 2696.985 1420.130 2702.330 1420.675 ;
        RECT 2702.505 1420.130 2707.850 1420.675 ;
        RECT 2708.025 1420.130 2713.370 1420.675 ;
        RECT 2713.545 1420.130 2718.890 1420.675 ;
        RECT 2695.605 1419.385 2696.125 1419.925 ;
        RECT 2698.570 1419.300 2698.910 1420.130 ;
        RECT 2704.090 1419.300 2704.430 1420.130 ;
        RECT 2709.610 1419.300 2709.950 1420.130 ;
        RECT 2715.130 1419.300 2715.470 1420.130 ;
        RECT 2719.065 1419.905 2720.735 1420.675 ;
        RECT 2721.365 1419.950 2721.655 1420.675 ;
        RECT 2721.825 1420.130 2727.170 1420.675 ;
        RECT 2727.345 1420.130 2732.690 1420.675 ;
        RECT 2719.065 1419.385 2719.815 1419.905 ;
        RECT 2723.410 1419.300 2723.750 1420.130 ;
        RECT 2728.930 1419.300 2729.270 1420.130 ;
        RECT 2732.865 1419.925 2734.075 1420.675 ;
        RECT 2733.555 1419.385 2734.075 1419.925 ;
        RECT 2523.330 1415.790 2523.670 1416.450 ;
        RECT 2695.605 1416.155 2696.125 1416.695 ;
        RECT 2522.130 1415.620 2523.935 1415.790 ;
        RECT 2695.605 1415.405 2696.815 1416.155 ;
        RECT 2699.950 1415.950 2700.290 1416.780 ;
        RECT 2703.885 1416.175 2705.535 1416.695 ;
        RECT 2697.425 1415.405 2697.755 1415.785 ;
        RECT 2698.365 1415.405 2703.710 1415.950 ;
        RECT 2703.885 1415.405 2707.395 1416.175 ;
        RECT 2708.485 1415.405 2708.775 1416.130 ;
        RECT 2710.530 1415.950 2710.870 1416.780 ;
        RECT 2716.050 1415.950 2716.390 1416.780 ;
        RECT 2721.570 1415.950 2721.910 1416.780 ;
        RECT 2727.090 1415.950 2727.430 1416.780 ;
        RECT 2731.025 1416.175 2731.775 1416.695 ;
        RECT 2708.945 1415.405 2714.290 1415.950 ;
        RECT 2714.465 1415.405 2719.810 1415.950 ;
        RECT 2719.985 1415.405 2725.330 1415.950 ;
        RECT 2725.505 1415.405 2730.850 1415.950 ;
        RECT 2731.025 1415.405 2732.695 1416.175 ;
        RECT 2733.555 1416.155 2734.075 1416.695 ;
        RECT 2732.865 1415.405 2734.075 1416.155 ;
        RECT 2695.520 1415.235 2734.160 1415.405 ;
        RECT 2695.605 1414.485 2696.815 1415.235 ;
        RECT 2696.985 1414.690 2702.330 1415.235 ;
        RECT 2702.505 1414.690 2707.850 1415.235 ;
        RECT 2708.025 1414.690 2713.370 1415.235 ;
        RECT 2713.545 1414.690 2718.890 1415.235 ;
        RECT 2695.605 1413.945 2696.125 1414.485 ;
        RECT 2698.570 1413.860 2698.910 1414.690 ;
        RECT 2704.090 1413.860 2704.430 1414.690 ;
        RECT 2709.610 1413.860 2709.950 1414.690 ;
        RECT 2715.130 1413.860 2715.470 1414.690 ;
        RECT 2719.065 1414.465 2720.735 1415.235 ;
        RECT 2721.365 1414.510 2721.655 1415.235 ;
        RECT 2721.825 1414.690 2727.170 1415.235 ;
        RECT 2727.345 1414.690 2732.690 1415.235 ;
        RECT 2719.065 1413.945 2719.815 1414.465 ;
        RECT 2723.410 1413.860 2723.750 1414.690 ;
        RECT 2728.930 1413.860 2729.270 1414.690 ;
        RECT 2732.865 1414.485 2734.075 1415.235 ;
        RECT 2733.555 1413.945 2734.075 1414.485 ;
        RECT 2695.605 1410.715 2696.125 1411.255 ;
        RECT 2695.605 1409.965 2696.815 1410.715 ;
        RECT 2701.330 1410.510 2701.670 1411.340 ;
        RECT 2705.265 1410.735 2706.475 1411.255 ;
        RECT 2697.425 1409.965 2697.755 1410.345 ;
        RECT 2698.805 1409.965 2699.135 1410.345 ;
        RECT 2699.745 1409.965 2705.090 1410.510 ;
        RECT 2705.265 1409.965 2707.855 1410.735 ;
        RECT 2708.485 1409.965 2708.775 1410.690 ;
        RECT 2710.530 1410.510 2710.870 1411.340 ;
        RECT 2716.050 1410.510 2716.390 1411.340 ;
        RECT 2719.985 1410.715 2720.505 1411.255 ;
        RECT 2708.945 1409.965 2714.290 1410.510 ;
        RECT 2714.465 1409.965 2719.810 1410.510 ;
        RECT 2719.985 1409.965 2721.195 1410.715 ;
        RECT 2721.365 1409.965 2721.655 1410.690 ;
        RECT 2723.410 1410.510 2723.750 1411.340 ;
        RECT 2728.930 1410.510 2729.270 1411.340 ;
        RECT 2733.555 1410.715 2734.075 1411.255 ;
        RECT 2721.825 1409.965 2727.170 1410.510 ;
        RECT 2727.345 1409.965 2732.690 1410.510 ;
        RECT 2732.865 1409.965 2734.075 1410.715 ;
        RECT 2695.520 1409.795 2734.160 1409.965 ;
        RECT 2523.330 1408.260 2523.670 1408.920 ;
        RECT 2522.130 1408.090 2523.935 1408.260 ;
        RECT 2523.330 1402.280 2523.670 1402.940 ;
        RECT 2522.130 1402.110 2523.935 1402.280 ;
        RECT 2523.330 1393.865 2523.670 1394.525 ;
        RECT 2522.130 1393.695 2523.935 1393.865 ;
        RECT 2882.265 1360.590 2882.605 1361.250 ;
        RECT 2881.575 1360.420 2883.380 1360.590 ;
        RECT 2343.000 1335.865 2447.095 1337.465 ;
        RECT 2368.215 1335.240 2368.385 1335.865 ;
        RECT 2375.730 1335.240 2375.900 1335.865 ;
        RECT 2376.685 1335.320 2376.855 1335.600 ;
        RECT 2376.685 1335.150 2376.915 1335.320 ;
        RECT 2381.345 1335.240 2381.515 1335.865 ;
        RECT 2384.090 1335.240 2384.260 1335.865 ;
        RECT 2385.080 1335.240 2385.250 1335.865 ;
        RECT 2390.990 1335.240 2391.160 1335.865 ;
        RECT 2391.945 1335.320 2392.115 1335.600 ;
        RECT 2391.945 1335.150 2392.175 1335.320 ;
        RECT 2396.605 1335.240 2396.775 1335.865 ;
        RECT 2399.350 1335.240 2399.520 1335.865 ;
        RECT 2400.340 1335.240 2400.510 1335.865 ;
        RECT 2406.250 1335.240 2406.420 1335.865 ;
        RECT 2407.205 1335.320 2407.375 1335.600 ;
        RECT 2407.205 1335.150 2407.435 1335.320 ;
        RECT 2411.865 1335.240 2412.035 1335.865 ;
        RECT 2414.610 1335.240 2414.780 1335.865 ;
        RECT 2415.600 1335.240 2415.770 1335.865 ;
        RECT 2421.510 1335.240 2421.680 1335.865 ;
        RECT 2422.465 1335.320 2422.635 1335.600 ;
        RECT 2422.465 1335.150 2422.695 1335.320 ;
        RECT 2427.125 1335.240 2427.295 1335.865 ;
        RECT 2429.870 1335.240 2430.040 1335.865 ;
        RECT 2430.860 1335.240 2431.030 1335.865 ;
        RECT 2436.770 1335.240 2436.940 1335.865 ;
        RECT 2437.725 1335.320 2437.895 1335.600 ;
        RECT 2437.725 1335.150 2437.955 1335.320 ;
        RECT 2442.385 1335.240 2442.555 1335.865 ;
        RECT 2445.130 1335.240 2445.300 1335.865 ;
        RECT 2446.120 1335.240 2446.290 1335.865 ;
        RECT 2376.745 1333.540 2376.915 1335.150 ;
        RECT 2392.005 1333.540 2392.175 1335.150 ;
        RECT 2407.265 1333.540 2407.435 1335.150 ;
        RECT 2422.525 1333.540 2422.695 1335.150 ;
        RECT 2437.785 1333.540 2437.955 1335.150 ;
        RECT 2376.685 1333.370 2376.915 1333.540 ;
        RECT 2391.945 1333.370 2392.175 1333.540 ;
        RECT 2407.205 1333.370 2407.435 1333.540 ;
        RECT 2422.465 1333.370 2422.695 1333.540 ;
        RECT 2437.725 1333.370 2437.955 1333.540 ;
        RECT 2376.685 1332.310 2376.855 1333.370 ;
        RECT 2391.945 1332.310 2392.115 1333.370 ;
        RECT 2407.205 1332.310 2407.375 1333.370 ;
        RECT 2422.465 1332.310 2422.635 1333.370 ;
        RECT 2437.725 1332.310 2437.895 1333.370 ;
        RECT 2372.095 1328.785 2372.265 1329.235 ;
        RECT 2373.415 1328.865 2373.785 1329.035 ;
        RECT 2373.415 1328.395 2373.585 1328.865 ;
        RECT 2387.355 1328.785 2387.525 1329.235 ;
        RECT 2388.675 1328.865 2389.045 1329.035 ;
        RECT 2388.675 1328.395 2388.845 1328.865 ;
        RECT 2402.615 1328.785 2402.785 1329.235 ;
        RECT 2403.935 1328.865 2404.305 1329.035 ;
        RECT 2403.935 1328.395 2404.105 1328.865 ;
        RECT 2417.875 1328.785 2418.045 1329.235 ;
        RECT 2419.195 1328.865 2419.565 1329.035 ;
        RECT 2419.195 1328.395 2419.365 1328.865 ;
        RECT 2433.135 1328.785 2433.305 1329.235 ;
        RECT 2434.455 1328.865 2434.825 1329.035 ;
        RECT 2434.455 1328.395 2434.625 1328.865 ;
        RECT 2372.815 1327.890 2372.985 1328.375 ;
        RECT 2373.295 1328.225 2373.585 1328.395 ;
        RECT 2372.815 1327.875 2373.090 1327.890 ;
        RECT 2374.735 1327.875 2374.905 1328.375 ;
        RECT 2375.695 1327.875 2375.865 1328.375 ;
        RECT 2376.570 1327.875 2376.765 1327.890 ;
        RECT 2377.615 1327.875 2377.785 1328.375 ;
        RECT 2378.575 1327.880 2378.745 1328.375 ;
        RECT 2378.420 1327.875 2378.745 1327.880 ;
        RECT 2379.515 1327.875 2379.685 1328.375 ;
        RECT 2388.075 1327.890 2388.245 1328.375 ;
        RECT 2388.555 1328.225 2388.845 1328.395 ;
        RECT 2380.090 1327.875 2380.285 1327.880 ;
        RECT 2388.075 1327.875 2388.350 1327.890 ;
        RECT 2389.995 1327.875 2390.165 1328.375 ;
        RECT 2390.955 1327.875 2391.125 1328.375 ;
        RECT 2391.830 1327.875 2392.025 1327.890 ;
        RECT 2392.875 1327.875 2393.045 1328.375 ;
        RECT 2393.835 1327.880 2394.005 1328.375 ;
        RECT 2393.680 1327.875 2394.005 1327.880 ;
        RECT 2394.775 1327.875 2394.945 1328.375 ;
        RECT 2403.335 1327.890 2403.505 1328.375 ;
        RECT 2403.815 1328.225 2404.105 1328.395 ;
        RECT 2395.350 1327.875 2395.545 1327.880 ;
        RECT 2403.335 1327.875 2403.610 1327.890 ;
        RECT 2405.255 1327.875 2405.425 1328.375 ;
        RECT 2406.215 1327.875 2406.385 1328.375 ;
        RECT 2407.090 1327.875 2407.285 1327.890 ;
        RECT 2408.135 1327.875 2408.305 1328.375 ;
        RECT 2409.095 1327.880 2409.265 1328.375 ;
        RECT 2408.940 1327.875 2409.265 1327.880 ;
        RECT 2410.035 1327.875 2410.205 1328.375 ;
        RECT 2418.595 1327.890 2418.765 1328.375 ;
        RECT 2419.075 1328.225 2419.365 1328.395 ;
        RECT 2410.610 1327.875 2410.805 1327.880 ;
        RECT 2418.595 1327.875 2418.870 1327.890 ;
        RECT 2420.515 1327.875 2420.685 1328.375 ;
        RECT 2421.475 1327.875 2421.645 1328.375 ;
        RECT 2422.350 1327.875 2422.545 1327.890 ;
        RECT 2423.395 1327.875 2423.565 1328.375 ;
        RECT 2424.355 1327.880 2424.525 1328.375 ;
        RECT 2424.200 1327.875 2424.525 1327.880 ;
        RECT 2425.295 1327.875 2425.465 1328.375 ;
        RECT 2433.855 1327.890 2434.025 1328.375 ;
        RECT 2434.335 1328.225 2434.625 1328.395 ;
        RECT 2425.870 1327.875 2426.065 1327.880 ;
        RECT 2433.855 1327.875 2434.130 1327.890 ;
        RECT 2435.775 1327.875 2435.945 1328.375 ;
        RECT 2436.735 1327.875 2436.905 1328.375 ;
        RECT 2437.610 1327.875 2437.805 1327.890 ;
        RECT 2438.655 1327.875 2438.825 1328.375 ;
        RECT 2439.615 1327.880 2439.785 1328.375 ;
        RECT 2439.460 1327.875 2439.785 1327.880 ;
        RECT 2440.555 1327.875 2440.725 1328.375 ;
        RECT 2441.130 1327.875 2441.325 1327.880 ;
        RECT 2371.545 1326.600 2380.285 1327.875 ;
        RECT 2381.345 1326.600 2381.515 1327.225 ;
        RECT 2384.090 1326.600 2384.260 1327.225 ;
        RECT 2385.075 1326.600 2385.245 1327.225 ;
        RECT 2386.805 1326.600 2395.545 1327.875 ;
        RECT 2396.605 1326.600 2396.775 1327.225 ;
        RECT 2399.350 1326.600 2399.520 1327.225 ;
        RECT 2400.335 1326.600 2400.505 1327.225 ;
        RECT 2402.065 1326.600 2410.805 1327.875 ;
        RECT 2411.865 1326.600 2412.035 1327.225 ;
        RECT 2414.610 1326.600 2414.780 1327.225 ;
        RECT 2415.595 1326.600 2415.765 1327.225 ;
        RECT 2417.325 1326.600 2426.065 1327.875 ;
        RECT 2427.125 1326.600 2427.295 1327.225 ;
        RECT 2429.870 1326.600 2430.040 1327.225 ;
        RECT 2430.855 1326.600 2431.025 1327.225 ;
        RECT 2432.585 1326.600 2441.325 1327.875 ;
        RECT 2442.385 1326.600 2442.555 1327.225 ;
        RECT 2445.130 1326.600 2445.300 1327.225 ;
        RECT 2446.115 1326.600 2446.285 1327.225 ;
        RECT 2343.000 1325.000 2447.095 1326.600 ;
        RECT 2882.265 1161.350 2882.605 1162.010 ;
        RECT 2881.575 1161.180 2883.380 1161.350 ;
      LAYER met1 ;
        RECT 1262.805 3512.595 1264.185 3512.630 ;
        RECT 1271.170 3512.595 1274.270 3513.715 ;
        RECT 1622.805 3513.045 1624.185 3513.080 ;
        RECT 1631.170 3513.045 1634.270 3514.165 ;
        RECT 1622.805 3512.925 1634.350 3513.045 ;
        RECT 1622.380 3512.755 1634.350 3512.925 ;
        RECT 1622.805 3512.600 1634.350 3512.755 ;
        RECT 1262.805 3512.150 1274.350 3512.595 ;
        RECT 1623.980 3512.565 1634.350 3512.600 ;
        RECT 1263.980 3512.115 1274.350 3512.150 ;
        RECT 1802.805 3511.125 1804.185 3511.160 ;
        RECT 1811.170 3511.125 1814.270 3512.245 ;
        RECT 1802.805 3511.005 1814.350 3511.125 ;
        RECT 1802.380 3510.835 1814.350 3511.005 ;
        RECT 1802.805 3510.680 1814.350 3510.835 ;
        RECT 1803.980 3510.645 1814.350 3510.680 ;
        RECT 2162.805 3510.765 2164.185 3510.800 ;
        RECT 2171.170 3510.765 2174.270 3511.885 ;
        RECT 2522.805 3511.450 2524.185 3511.485 ;
        RECT 2531.170 3511.450 2534.270 3512.570 ;
        RECT 2522.805 3511.330 2534.350 3511.450 ;
        RECT 2522.380 3511.160 2534.350 3511.330 ;
        RECT 2522.805 3511.005 2534.350 3511.160 ;
        RECT 2523.980 3510.970 2534.350 3511.005 ;
        RECT 2162.805 3510.645 2174.350 3510.765 ;
        RECT 2162.380 3510.475 2174.350 3510.645 ;
        RECT 2162.805 3510.320 2174.350 3510.475 ;
        RECT 2163.980 3510.285 2174.350 3510.320 ;
        RECT 2882.000 3485.590 2894.380 3485.745 ;
        RECT 2881.575 3485.420 2894.380 3485.590 ;
        RECT 2882.000 3485.265 2894.380 3485.420 ;
        RECT 2891.170 3484.010 2894.270 3485.265 ;
        RECT 2882.000 3219.710 2894.380 3219.865 ;
        RECT 2881.575 3219.540 2894.380 3219.710 ;
        RECT 2882.000 3219.385 2894.380 3219.540 ;
        RECT 2891.170 3218.130 2894.270 3219.385 ;
        RECT 2882.000 2954.510 2894.380 2954.665 ;
        RECT 2881.575 2954.340 2894.380 2954.510 ;
        RECT 2882.000 2954.185 2894.380 2954.340 ;
        RECT 2891.170 2952.930 2894.270 2954.185 ;
        RECT 2882.000 2688.630 2894.380 2688.785 ;
        RECT 2881.575 2688.460 2894.380 2688.630 ;
        RECT 2882.000 2688.305 2894.380 2688.460 ;
        RECT 2891.170 2687.050 2894.270 2688.305 ;
        RECT 2882.000 2422.750 2894.380 2422.905 ;
        RECT 2881.575 2422.580 2894.380 2422.750 ;
        RECT 2882.000 2422.425 2894.380 2422.580 ;
        RECT 2891.170 2421.170 2894.270 2422.425 ;
        RECT 2343.055 2255.855 2443.725 2257.455 ;
        RECT 2362.245 2253.805 2362.415 2255.855 ;
        RECT 2362.245 2253.775 2362.700 2253.805 ;
        RECT 2362.235 2253.605 2362.700 2253.775 ;
        RECT 2364.515 2253.685 2364.765 2255.855 ;
        RECT 2365.040 2253.685 2365.315 2255.855 ;
        RECT 2365.590 2253.685 2365.865 2255.855 ;
        RECT 2366.140 2253.685 2366.415 2255.855 ;
        RECT 2366.690 2253.685 2366.965 2255.855 ;
        RECT 2367.240 2253.685 2367.515 2255.855 ;
        RECT 2367.790 2253.685 2368.065 2255.855 ;
        RECT 2368.340 2253.685 2368.615 2255.855 ;
        RECT 2368.890 2253.685 2369.165 2255.855 ;
        RECT 2369.440 2253.685 2369.715 2255.855 ;
        RECT 2369.990 2253.685 2370.265 2255.855 ;
        RECT 2370.540 2253.685 2370.815 2255.855 ;
        RECT 2371.090 2253.685 2371.435 2255.855 ;
        RECT 2378.830 2253.805 2379.000 2255.855 ;
        RECT 2378.830 2253.775 2379.285 2253.805 ;
        RECT 2362.245 2253.600 2362.700 2253.605 ;
        RECT 2362.410 2253.575 2362.700 2253.600 ;
        RECT 2364.380 2253.325 2371.435 2253.685 ;
        RECT 2378.820 2253.605 2379.285 2253.775 ;
        RECT 2381.100 2253.685 2381.350 2255.855 ;
        RECT 2381.625 2253.685 2381.900 2255.855 ;
        RECT 2382.175 2253.685 2382.450 2255.855 ;
        RECT 2382.725 2253.685 2383.000 2255.855 ;
        RECT 2383.275 2253.685 2383.550 2255.855 ;
        RECT 2383.825 2253.685 2384.100 2255.855 ;
        RECT 2384.375 2253.685 2384.650 2255.855 ;
        RECT 2384.925 2253.685 2385.200 2255.855 ;
        RECT 2385.475 2253.685 2385.750 2255.855 ;
        RECT 2386.025 2253.685 2386.300 2255.855 ;
        RECT 2386.575 2253.685 2386.850 2255.855 ;
        RECT 2387.125 2253.685 2387.400 2255.855 ;
        RECT 2387.675 2253.685 2388.020 2255.855 ;
        RECT 2395.415 2253.805 2395.585 2255.855 ;
        RECT 2395.415 2253.775 2395.870 2253.805 ;
        RECT 2378.830 2253.600 2379.285 2253.605 ;
        RECT 2378.995 2253.575 2379.285 2253.600 ;
        RECT 2380.965 2253.325 2388.020 2253.685 ;
        RECT 2395.405 2253.605 2395.870 2253.775 ;
        RECT 2397.685 2253.685 2397.935 2255.855 ;
        RECT 2398.210 2253.685 2398.485 2255.855 ;
        RECT 2398.760 2253.685 2399.035 2255.855 ;
        RECT 2399.310 2253.685 2399.585 2255.855 ;
        RECT 2399.860 2253.685 2400.135 2255.855 ;
        RECT 2400.410 2253.685 2400.685 2255.855 ;
        RECT 2400.960 2253.685 2401.235 2255.855 ;
        RECT 2401.510 2253.685 2401.785 2255.855 ;
        RECT 2402.060 2253.685 2402.335 2255.855 ;
        RECT 2402.610 2253.685 2402.885 2255.855 ;
        RECT 2403.160 2253.685 2403.435 2255.855 ;
        RECT 2403.710 2253.685 2403.985 2255.855 ;
        RECT 2404.260 2253.685 2404.605 2255.855 ;
        RECT 2412.000 2253.805 2412.170 2255.855 ;
        RECT 2412.000 2253.775 2412.455 2253.805 ;
        RECT 2395.415 2253.600 2395.870 2253.605 ;
        RECT 2395.580 2253.575 2395.870 2253.600 ;
        RECT 2397.550 2253.325 2404.605 2253.685 ;
        RECT 2411.990 2253.605 2412.455 2253.775 ;
        RECT 2414.270 2253.685 2414.520 2255.855 ;
        RECT 2414.795 2253.685 2415.070 2255.855 ;
        RECT 2415.345 2253.685 2415.620 2255.855 ;
        RECT 2415.895 2253.685 2416.170 2255.855 ;
        RECT 2416.445 2253.685 2416.720 2255.855 ;
        RECT 2416.995 2253.685 2417.270 2255.855 ;
        RECT 2417.545 2253.685 2417.820 2255.855 ;
        RECT 2418.095 2253.685 2418.370 2255.855 ;
        RECT 2418.645 2253.685 2418.920 2255.855 ;
        RECT 2419.195 2253.685 2419.470 2255.855 ;
        RECT 2419.745 2253.685 2420.020 2255.855 ;
        RECT 2420.295 2253.685 2420.570 2255.855 ;
        RECT 2420.845 2253.685 2421.190 2255.855 ;
        RECT 2428.580 2253.805 2428.750 2255.855 ;
        RECT 2428.580 2253.775 2429.035 2253.805 ;
        RECT 2412.000 2253.600 2412.455 2253.605 ;
        RECT 2412.165 2253.575 2412.455 2253.600 ;
        RECT 2414.135 2253.325 2421.190 2253.685 ;
        RECT 2428.570 2253.605 2429.035 2253.775 ;
        RECT 2430.850 2253.685 2431.100 2255.855 ;
        RECT 2431.375 2253.685 2431.650 2255.855 ;
        RECT 2431.925 2253.685 2432.200 2255.855 ;
        RECT 2432.475 2253.685 2432.750 2255.855 ;
        RECT 2433.025 2253.685 2433.300 2255.855 ;
        RECT 2433.575 2253.685 2433.850 2255.855 ;
        RECT 2434.125 2253.685 2434.400 2255.855 ;
        RECT 2434.675 2253.685 2434.950 2255.855 ;
        RECT 2435.225 2253.685 2435.500 2255.855 ;
        RECT 2435.775 2253.685 2436.050 2255.855 ;
        RECT 2436.325 2253.685 2436.600 2255.855 ;
        RECT 2436.875 2253.685 2437.150 2255.855 ;
        RECT 2437.425 2253.685 2437.770 2255.855 ;
        RECT 2428.580 2253.600 2429.035 2253.605 ;
        RECT 2428.745 2253.575 2429.035 2253.600 ;
        RECT 2430.715 2253.325 2437.770 2253.685 ;
        RECT 2365.980 2252.945 2366.120 2253.325 ;
        RECT 2366.910 2252.945 2367.340 2253.045 ;
        RECT 2382.565 2252.945 2382.705 2253.325 ;
        RECT 2383.495 2252.945 2383.925 2253.045 ;
        RECT 2399.150 2252.945 2399.290 2253.325 ;
        RECT 2400.080 2252.945 2400.510 2253.045 ;
        RECT 2415.735 2252.945 2415.875 2253.325 ;
        RECT 2416.665 2252.945 2417.095 2253.045 ;
        RECT 2432.315 2252.945 2432.455 2253.325 ;
        RECT 2433.245 2252.945 2433.675 2253.045 ;
        RECT 2365.980 2252.805 2368.330 2252.945 ;
        RECT 2365.980 2252.365 2366.120 2252.805 ;
        RECT 2366.920 2252.775 2367.200 2252.805 ;
        RECT 2366.940 2252.745 2367.200 2252.775 ;
        RECT 2368.190 2252.365 2368.330 2252.805 ;
        RECT 2382.565 2252.805 2384.915 2252.945 ;
        RECT 2382.565 2252.365 2382.705 2252.805 ;
        RECT 2383.505 2252.775 2383.785 2252.805 ;
        RECT 2383.525 2252.745 2383.785 2252.775 ;
        RECT 2384.775 2252.365 2384.915 2252.805 ;
        RECT 2399.150 2252.805 2401.500 2252.945 ;
        RECT 2399.150 2252.365 2399.290 2252.805 ;
        RECT 2400.090 2252.775 2400.370 2252.805 ;
        RECT 2400.110 2252.745 2400.370 2252.775 ;
        RECT 2401.360 2252.365 2401.500 2252.805 ;
        RECT 2415.735 2252.805 2418.085 2252.945 ;
        RECT 2415.735 2252.365 2415.875 2252.805 ;
        RECT 2416.675 2252.775 2416.955 2252.805 ;
        RECT 2416.695 2252.745 2416.955 2252.775 ;
        RECT 2417.945 2252.365 2418.085 2252.805 ;
        RECT 2432.315 2252.805 2434.665 2252.945 ;
        RECT 2432.315 2252.365 2432.455 2252.805 ;
        RECT 2433.255 2252.775 2433.535 2252.805 ;
        RECT 2433.275 2252.745 2433.535 2252.775 ;
        RECT 2434.525 2252.365 2434.665 2252.805 ;
        RECT 2365.900 2252.135 2366.190 2252.365 ;
        RECT 2368.110 2252.135 2368.400 2252.365 ;
        RECT 2382.485 2252.135 2382.775 2252.365 ;
        RECT 2384.695 2252.135 2384.985 2252.365 ;
        RECT 2399.070 2252.135 2399.360 2252.365 ;
        RECT 2401.280 2252.135 2401.570 2252.365 ;
        RECT 2415.655 2252.135 2415.945 2252.365 ;
        RECT 2417.865 2252.135 2418.155 2252.365 ;
        RECT 2432.235 2252.135 2432.525 2252.365 ;
        RECT 2434.445 2252.135 2434.735 2252.365 ;
        RECT 2364.220 2247.765 2371.610 2248.125 ;
        RECT 2380.805 2247.765 2388.195 2248.125 ;
        RECT 2397.390 2247.765 2404.780 2248.125 ;
        RECT 2413.975 2247.765 2421.365 2248.125 ;
        RECT 2430.555 2247.765 2437.945 2248.125 ;
        RECT 2364.265 2246.600 2364.525 2247.765 ;
        RECT 2364.815 2246.600 2365.075 2247.765 ;
        RECT 2365.355 2246.600 2365.615 2247.765 ;
        RECT 2365.895 2246.600 2366.135 2247.765 ;
        RECT 2366.435 2246.600 2366.675 2247.765 ;
        RECT 2366.955 2246.600 2367.195 2247.765 ;
        RECT 2367.475 2246.600 2367.715 2247.765 ;
        RECT 2367.995 2246.600 2368.235 2247.765 ;
        RECT 2368.515 2246.600 2368.755 2247.765 ;
        RECT 2368.995 2246.600 2369.235 2247.765 ;
        RECT 2369.475 2246.600 2369.715 2247.765 ;
        RECT 2369.955 2246.600 2370.195 2247.765 ;
        RECT 2370.435 2246.600 2370.675 2247.765 ;
        RECT 2370.915 2246.600 2371.155 2247.765 ;
        RECT 2371.395 2246.600 2371.610 2247.765 ;
        RECT 2380.850 2246.600 2381.110 2247.765 ;
        RECT 2381.400 2246.600 2381.660 2247.765 ;
        RECT 2381.940 2246.600 2382.200 2247.765 ;
        RECT 2382.480 2246.600 2382.720 2247.765 ;
        RECT 2383.020 2246.600 2383.260 2247.765 ;
        RECT 2383.540 2246.600 2383.780 2247.765 ;
        RECT 2384.060 2246.600 2384.300 2247.765 ;
        RECT 2384.580 2246.600 2384.820 2247.765 ;
        RECT 2385.100 2246.600 2385.340 2247.765 ;
        RECT 2385.580 2246.600 2385.820 2247.765 ;
        RECT 2386.060 2246.600 2386.300 2247.765 ;
        RECT 2386.540 2246.600 2386.780 2247.765 ;
        RECT 2387.020 2246.600 2387.260 2247.765 ;
        RECT 2387.500 2246.600 2387.740 2247.765 ;
        RECT 2387.980 2246.600 2388.195 2247.765 ;
        RECT 2397.435 2246.600 2397.695 2247.765 ;
        RECT 2397.985 2246.600 2398.245 2247.765 ;
        RECT 2398.525 2246.600 2398.785 2247.765 ;
        RECT 2399.065 2246.600 2399.305 2247.765 ;
        RECT 2399.605 2246.600 2399.845 2247.765 ;
        RECT 2400.125 2246.600 2400.365 2247.765 ;
        RECT 2400.645 2246.600 2400.885 2247.765 ;
        RECT 2401.165 2246.600 2401.405 2247.765 ;
        RECT 2401.685 2246.600 2401.925 2247.765 ;
        RECT 2402.165 2246.600 2402.405 2247.765 ;
        RECT 2402.645 2246.600 2402.885 2247.765 ;
        RECT 2403.125 2246.600 2403.365 2247.765 ;
        RECT 2403.605 2246.600 2403.845 2247.765 ;
        RECT 2404.085 2246.600 2404.325 2247.765 ;
        RECT 2404.565 2246.600 2404.780 2247.765 ;
        RECT 2414.020 2246.600 2414.280 2247.765 ;
        RECT 2414.570 2246.600 2414.830 2247.765 ;
        RECT 2415.110 2246.600 2415.370 2247.765 ;
        RECT 2415.650 2246.600 2415.890 2247.765 ;
        RECT 2416.190 2246.600 2416.430 2247.765 ;
        RECT 2416.710 2246.600 2416.950 2247.765 ;
        RECT 2417.230 2246.600 2417.470 2247.765 ;
        RECT 2417.750 2246.600 2417.990 2247.765 ;
        RECT 2418.270 2246.600 2418.510 2247.765 ;
        RECT 2418.750 2246.600 2418.990 2247.765 ;
        RECT 2419.230 2246.600 2419.470 2247.765 ;
        RECT 2419.710 2246.600 2419.950 2247.765 ;
        RECT 2420.190 2246.600 2420.430 2247.765 ;
        RECT 2420.670 2246.600 2420.910 2247.765 ;
        RECT 2421.150 2246.600 2421.365 2247.765 ;
        RECT 2430.600 2246.600 2430.860 2247.765 ;
        RECT 2431.150 2246.600 2431.410 2247.765 ;
        RECT 2431.690 2246.600 2431.950 2247.765 ;
        RECT 2432.230 2246.600 2432.470 2247.765 ;
        RECT 2432.770 2246.600 2433.010 2247.765 ;
        RECT 2433.290 2246.600 2433.530 2247.765 ;
        RECT 2433.810 2246.600 2434.050 2247.765 ;
        RECT 2434.330 2246.600 2434.570 2247.765 ;
        RECT 2434.850 2246.600 2435.090 2247.765 ;
        RECT 2435.330 2246.600 2435.570 2247.765 ;
        RECT 2435.810 2246.600 2436.050 2247.765 ;
        RECT 2436.290 2246.600 2436.530 2247.765 ;
        RECT 2436.770 2246.600 2437.010 2247.765 ;
        RECT 2437.250 2246.600 2437.490 2247.765 ;
        RECT 2437.730 2246.600 2437.945 2247.765 ;
        RECT 2343.000 2245.000 2443.725 2246.600 ;
        RECT 2695.520 2216.680 2734.960 2217.160 ;
        RECT 2695.520 2211.240 2734.960 2211.720 ;
        RECT 2695.520 2205.800 2734.960 2206.280 ;
        RECT 2695.520 2200.360 2734.960 2200.840 ;
        RECT 2695.520 2194.920 2734.960 2195.400 ;
        RECT 2695.520 2189.480 2734.960 2189.960 ;
        RECT 2695.520 2184.040 2734.960 2184.520 ;
        RECT 2695.520 2178.600 2734.960 2179.080 ;
        RECT 2695.520 2173.160 2734.960 2173.640 ;
        RECT 2695.520 2167.720 2734.960 2168.200 ;
        RECT 2343.000 2163.860 2446.925 2165.460 ;
        RECT 2361.480 2163.855 2364.230 2163.860 ;
        RECT 2362.200 2161.775 2362.370 2163.855 ;
        RECT 2362.605 2161.775 2362.895 2161.805 ;
        RECT 2362.200 2161.595 2362.895 2161.775 ;
        RECT 2362.605 2161.575 2362.895 2161.595 ;
        RECT 2364.610 2161.685 2364.895 2163.860 ;
        RECT 2365.180 2161.685 2365.465 2163.860 ;
        RECT 2365.750 2161.685 2366.035 2163.860 ;
        RECT 2366.320 2161.685 2366.605 2163.860 ;
        RECT 2366.890 2161.685 2367.175 2163.860 ;
        RECT 2367.460 2161.685 2367.745 2163.860 ;
        RECT 2368.030 2161.685 2368.315 2163.860 ;
        RECT 2368.600 2161.685 2368.885 2163.860 ;
        RECT 2369.170 2161.685 2369.450 2163.860 ;
        RECT 2369.735 2161.685 2370.020 2163.860 ;
        RECT 2370.305 2161.685 2370.590 2163.860 ;
        RECT 2370.875 2161.685 2371.160 2163.860 ;
        RECT 2371.730 2161.685 2371.970 2163.860 ;
        RECT 2378.700 2163.855 2381.450 2163.860 ;
        RECT 2364.610 2161.330 2371.970 2161.685 ;
        RECT 2379.420 2161.775 2379.590 2163.855 ;
        RECT 2379.825 2161.775 2380.115 2161.805 ;
        RECT 2379.420 2161.595 2380.115 2161.775 ;
        RECT 2379.825 2161.575 2380.115 2161.595 ;
        RECT 2381.830 2161.685 2382.115 2163.860 ;
        RECT 2382.400 2161.685 2382.685 2163.860 ;
        RECT 2382.970 2161.685 2383.255 2163.860 ;
        RECT 2383.540 2161.685 2383.825 2163.860 ;
        RECT 2384.110 2161.685 2384.395 2163.860 ;
        RECT 2384.680 2161.685 2384.965 2163.860 ;
        RECT 2385.250 2161.685 2385.535 2163.860 ;
        RECT 2385.820 2161.685 2386.105 2163.860 ;
        RECT 2386.390 2161.685 2386.670 2163.860 ;
        RECT 2386.955 2161.685 2387.240 2163.860 ;
        RECT 2387.525 2161.685 2387.810 2163.860 ;
        RECT 2388.095 2161.685 2388.380 2163.860 ;
        RECT 2388.950 2161.685 2389.190 2163.860 ;
        RECT 2395.920 2163.855 2398.670 2163.860 ;
        RECT 2381.830 2161.330 2389.190 2161.685 ;
        RECT 2396.640 2161.775 2396.810 2163.855 ;
        RECT 2397.045 2161.775 2397.335 2161.805 ;
        RECT 2396.640 2161.595 2397.335 2161.775 ;
        RECT 2397.045 2161.575 2397.335 2161.595 ;
        RECT 2399.050 2161.685 2399.335 2163.860 ;
        RECT 2399.620 2161.685 2399.905 2163.860 ;
        RECT 2400.190 2161.685 2400.475 2163.860 ;
        RECT 2400.760 2161.685 2401.045 2163.860 ;
        RECT 2401.330 2161.685 2401.615 2163.860 ;
        RECT 2401.900 2161.685 2402.185 2163.860 ;
        RECT 2402.470 2161.685 2402.755 2163.860 ;
        RECT 2403.040 2161.685 2403.325 2163.860 ;
        RECT 2403.610 2161.685 2403.890 2163.860 ;
        RECT 2404.175 2161.685 2404.460 2163.860 ;
        RECT 2404.745 2161.685 2405.030 2163.860 ;
        RECT 2405.315 2161.685 2405.600 2163.860 ;
        RECT 2406.170 2161.685 2406.410 2163.860 ;
        RECT 2413.140 2163.855 2415.890 2163.860 ;
        RECT 2399.050 2161.330 2406.410 2161.685 ;
        RECT 2413.860 2161.775 2414.030 2163.855 ;
        RECT 2414.265 2161.775 2414.555 2161.805 ;
        RECT 2413.860 2161.595 2414.555 2161.775 ;
        RECT 2414.265 2161.575 2414.555 2161.595 ;
        RECT 2416.270 2161.685 2416.555 2163.860 ;
        RECT 2416.840 2161.685 2417.125 2163.860 ;
        RECT 2417.410 2161.685 2417.695 2163.860 ;
        RECT 2417.980 2161.685 2418.265 2163.860 ;
        RECT 2418.550 2161.685 2418.835 2163.860 ;
        RECT 2419.120 2161.685 2419.405 2163.860 ;
        RECT 2419.690 2161.685 2419.975 2163.860 ;
        RECT 2420.260 2161.685 2420.545 2163.860 ;
        RECT 2420.830 2161.685 2421.110 2163.860 ;
        RECT 2421.395 2161.685 2421.680 2163.860 ;
        RECT 2421.965 2161.685 2422.250 2163.860 ;
        RECT 2422.535 2161.685 2422.820 2163.860 ;
        RECT 2423.390 2161.685 2423.630 2163.860 ;
        RECT 2430.360 2163.855 2433.110 2163.860 ;
        RECT 2416.270 2161.330 2423.630 2161.685 ;
        RECT 2431.080 2161.775 2431.250 2163.855 ;
        RECT 2431.485 2161.775 2431.775 2161.805 ;
        RECT 2431.080 2161.595 2431.775 2161.775 ;
        RECT 2431.485 2161.575 2431.775 2161.595 ;
        RECT 2433.490 2161.685 2433.775 2163.860 ;
        RECT 2434.060 2161.685 2434.345 2163.860 ;
        RECT 2434.630 2161.685 2434.915 2163.860 ;
        RECT 2435.200 2161.685 2435.485 2163.860 ;
        RECT 2435.770 2161.685 2436.055 2163.860 ;
        RECT 2436.340 2161.685 2436.625 2163.860 ;
        RECT 2436.910 2161.685 2437.195 2163.860 ;
        RECT 2437.480 2161.685 2437.765 2163.860 ;
        RECT 2438.050 2161.685 2438.330 2163.860 ;
        RECT 2438.615 2161.685 2438.900 2163.860 ;
        RECT 2439.185 2161.685 2439.470 2163.860 ;
        RECT 2439.755 2161.685 2440.040 2163.860 ;
        RECT 2440.610 2161.685 2440.850 2163.860 ;
        RECT 2695.520 2162.280 2734.960 2162.760 ;
        RECT 2433.490 2161.330 2440.850 2161.685 ;
        RECT 2364.635 2160.325 2364.925 2160.370 ;
        RECT 2367.000 2160.325 2367.320 2160.385 ;
        RECT 2364.635 2160.185 2367.320 2160.325 ;
        RECT 2364.635 2160.140 2364.925 2160.185 ;
        RECT 2367.000 2160.125 2367.320 2160.185 ;
        RECT 2381.855 2160.325 2382.145 2160.370 ;
        RECT 2384.220 2160.325 2384.540 2160.385 ;
        RECT 2381.855 2160.185 2384.540 2160.325 ;
        RECT 2381.855 2160.140 2382.145 2160.185 ;
        RECT 2384.220 2160.125 2384.540 2160.185 ;
        RECT 2399.075 2160.325 2399.365 2160.370 ;
        RECT 2401.440 2160.325 2401.760 2160.385 ;
        RECT 2399.075 2160.185 2401.760 2160.325 ;
        RECT 2399.075 2160.140 2399.365 2160.185 ;
        RECT 2401.440 2160.125 2401.760 2160.185 ;
        RECT 2416.295 2160.325 2416.585 2160.370 ;
        RECT 2418.660 2160.325 2418.980 2160.385 ;
        RECT 2416.295 2160.185 2418.980 2160.325 ;
        RECT 2416.295 2160.140 2416.585 2160.185 ;
        RECT 2418.660 2160.125 2418.980 2160.185 ;
        RECT 2433.515 2160.325 2433.805 2160.370 ;
        RECT 2435.880 2160.325 2436.200 2160.385 ;
        RECT 2433.515 2160.185 2436.200 2160.325 ;
        RECT 2433.515 2160.140 2433.805 2160.185 ;
        RECT 2435.880 2160.125 2436.200 2160.185 ;
        RECT 2882.000 2157.550 2894.380 2157.705 ;
        RECT 2881.575 2157.380 2894.380 2157.550 ;
        RECT 2695.520 2156.840 2734.960 2157.320 ;
        RECT 2882.000 2157.225 2894.380 2157.380 ;
        RECT 2364.605 2155.765 2372.265 2156.120 ;
        RECT 2364.605 2154.605 2364.885 2155.765 ;
        RECT 2365.170 2154.605 2365.455 2155.765 ;
        RECT 2365.740 2154.605 2366.025 2155.765 ;
        RECT 2366.310 2154.605 2366.595 2155.765 ;
        RECT 2366.880 2154.605 2367.165 2155.765 ;
        RECT 2367.450 2154.605 2367.735 2155.765 ;
        RECT 2368.020 2154.605 2368.305 2155.765 ;
        RECT 2368.590 2154.605 2368.875 2155.765 ;
        RECT 2369.160 2154.605 2369.445 2155.765 ;
        RECT 2369.730 2154.605 2370.015 2155.765 ;
        RECT 2370.300 2154.605 2370.585 2155.765 ;
        RECT 2370.870 2154.605 2371.155 2155.765 ;
        RECT 2371.440 2154.605 2371.725 2155.765 ;
        RECT 2372.010 2154.605 2372.265 2155.765 ;
        RECT 2364.605 2154.600 2372.265 2154.605 ;
        RECT 2381.825 2155.765 2389.485 2156.120 ;
        RECT 2381.825 2154.605 2382.105 2155.765 ;
        RECT 2382.390 2154.605 2382.675 2155.765 ;
        RECT 2382.960 2154.605 2383.245 2155.765 ;
        RECT 2383.530 2154.605 2383.815 2155.765 ;
        RECT 2384.100 2154.605 2384.385 2155.765 ;
        RECT 2384.670 2154.605 2384.955 2155.765 ;
        RECT 2385.240 2154.605 2385.525 2155.765 ;
        RECT 2385.810 2154.605 2386.095 2155.765 ;
        RECT 2386.380 2154.605 2386.665 2155.765 ;
        RECT 2386.950 2154.605 2387.235 2155.765 ;
        RECT 2387.520 2154.605 2387.805 2155.765 ;
        RECT 2388.090 2154.605 2388.375 2155.765 ;
        RECT 2388.660 2154.605 2388.945 2155.765 ;
        RECT 2389.230 2154.605 2389.485 2155.765 ;
        RECT 2381.825 2154.600 2389.485 2154.605 ;
        RECT 2399.045 2155.765 2406.705 2156.120 ;
        RECT 2399.045 2154.605 2399.325 2155.765 ;
        RECT 2399.610 2154.605 2399.895 2155.765 ;
        RECT 2400.180 2154.605 2400.465 2155.765 ;
        RECT 2400.750 2154.605 2401.035 2155.765 ;
        RECT 2401.320 2154.605 2401.605 2155.765 ;
        RECT 2401.890 2154.605 2402.175 2155.765 ;
        RECT 2402.460 2154.605 2402.745 2155.765 ;
        RECT 2403.030 2154.605 2403.315 2155.765 ;
        RECT 2403.600 2154.605 2403.885 2155.765 ;
        RECT 2404.170 2154.605 2404.455 2155.765 ;
        RECT 2404.740 2154.605 2405.025 2155.765 ;
        RECT 2405.310 2154.605 2405.595 2155.765 ;
        RECT 2405.880 2154.605 2406.165 2155.765 ;
        RECT 2406.450 2154.605 2406.705 2155.765 ;
        RECT 2399.045 2154.600 2406.705 2154.605 ;
        RECT 2416.265 2155.765 2423.925 2156.120 ;
        RECT 2416.265 2154.605 2416.545 2155.765 ;
        RECT 2416.830 2154.605 2417.115 2155.765 ;
        RECT 2417.400 2154.605 2417.685 2155.765 ;
        RECT 2417.970 2154.605 2418.255 2155.765 ;
        RECT 2418.540 2154.605 2418.825 2155.765 ;
        RECT 2419.110 2154.605 2419.395 2155.765 ;
        RECT 2419.680 2154.605 2419.965 2155.765 ;
        RECT 2420.250 2154.605 2420.535 2155.765 ;
        RECT 2420.820 2154.605 2421.105 2155.765 ;
        RECT 2421.390 2154.605 2421.675 2155.765 ;
        RECT 2421.960 2154.605 2422.245 2155.765 ;
        RECT 2422.530 2154.605 2422.815 2155.765 ;
        RECT 2423.100 2154.605 2423.385 2155.765 ;
        RECT 2423.670 2154.605 2423.925 2155.765 ;
        RECT 2416.265 2154.600 2423.925 2154.605 ;
        RECT 2433.485 2155.765 2441.145 2156.120 ;
        RECT 2891.170 2155.970 2894.270 2157.225 ;
        RECT 2433.485 2154.605 2433.765 2155.765 ;
        RECT 2434.050 2154.605 2434.335 2155.765 ;
        RECT 2434.620 2154.605 2434.905 2155.765 ;
        RECT 2435.190 2154.605 2435.475 2155.765 ;
        RECT 2435.760 2154.605 2436.045 2155.765 ;
        RECT 2436.330 2154.605 2436.615 2155.765 ;
        RECT 2436.900 2154.605 2437.185 2155.765 ;
        RECT 2437.470 2154.605 2437.755 2155.765 ;
        RECT 2438.040 2154.605 2438.325 2155.765 ;
        RECT 2438.610 2154.605 2438.895 2155.765 ;
        RECT 2439.180 2154.605 2439.465 2155.765 ;
        RECT 2439.750 2154.605 2440.035 2155.765 ;
        RECT 2440.320 2154.605 2440.605 2155.765 ;
        RECT 2440.890 2154.605 2441.145 2155.765 ;
        RECT 2433.485 2154.600 2441.145 2154.605 ;
        RECT 2343.015 2153.000 2446.925 2154.600 ;
        RECT 2695.520 2151.400 2734.960 2151.880 ;
        RECT 2695.520 2145.960 2734.960 2146.440 ;
        RECT 2695.520 2140.520 2734.960 2141.000 ;
        RECT 2695.520 2135.080 2734.960 2135.560 ;
        RECT 2522.555 2134.040 2534.570 2134.195 ;
        RECT 2522.130 2133.870 2534.570 2134.040 ;
        RECT 2522.555 2133.715 2534.570 2133.870 ;
        RECT 2531.170 2132.595 2534.270 2133.715 ;
        RECT 2695.520 2129.640 2734.960 2130.120 ;
        RECT 2522.555 2126.510 2534.570 2126.665 ;
        RECT 2522.130 2126.340 2534.570 2126.510 ;
        RECT 2522.555 2126.185 2534.570 2126.340 ;
        RECT 2531.170 2125.065 2534.270 2126.185 ;
        RECT 2522.555 2120.530 2534.570 2120.685 ;
        RECT 2522.130 2120.360 2534.570 2120.530 ;
        RECT 2522.555 2120.205 2534.570 2120.360 ;
        RECT 2531.170 2119.085 2534.270 2120.205 ;
        RECT 2522.555 2114.585 2534.570 2114.740 ;
        RECT 2522.130 2114.415 2534.570 2114.585 ;
        RECT 2522.555 2114.260 2534.570 2114.415 ;
        RECT 2531.170 2113.140 2534.270 2114.260 ;
        RECT 2522.555 2108.940 2534.570 2109.095 ;
        RECT 2522.130 2108.770 2534.570 2108.940 ;
        RECT 2522.555 2108.615 2534.570 2108.770 ;
        RECT 2531.170 2107.495 2534.270 2108.615 ;
        RECT 2522.555 2102.935 2534.570 2103.090 ;
        RECT 2522.130 2102.765 2534.570 2102.935 ;
        RECT 2522.555 2102.610 2534.570 2102.765 ;
        RECT 2531.170 2101.490 2534.270 2102.610 ;
        RECT 2343.050 2058.860 2442.430 2060.460 ;
        RECT 2367.375 2056.785 2367.550 2058.860 ;
        RECT 2367.755 2056.785 2368.045 2056.815 ;
        RECT 2367.375 2056.600 2368.045 2056.785 ;
        RECT 2383.700 2056.785 2383.875 2058.860 ;
        RECT 2384.080 2056.785 2384.370 2056.815 ;
        RECT 2383.700 2056.600 2384.370 2056.785 ;
        RECT 2400.025 2056.785 2400.200 2058.860 ;
        RECT 2400.405 2056.785 2400.695 2056.815 ;
        RECT 2400.025 2056.600 2400.695 2056.785 ;
        RECT 2416.350 2056.785 2416.525 2058.860 ;
        RECT 2416.730 2056.785 2417.020 2056.815 ;
        RECT 2416.350 2056.600 2417.020 2056.785 ;
        RECT 2432.675 2056.785 2432.850 2058.860 ;
        RECT 2433.055 2056.785 2433.345 2056.815 ;
        RECT 2432.675 2056.600 2433.345 2056.785 ;
        RECT 2367.755 2056.585 2368.045 2056.600 ;
        RECT 2384.080 2056.585 2384.370 2056.600 ;
        RECT 2400.405 2056.585 2400.695 2056.600 ;
        RECT 2416.730 2056.585 2417.020 2056.600 ;
        RECT 2433.055 2056.585 2433.345 2056.600 ;
        RECT 2368.940 2052.350 2370.540 2052.365 ;
        RECT 2385.265 2052.350 2386.865 2052.365 ;
        RECT 2401.590 2052.350 2403.190 2052.365 ;
        RECT 2417.915 2052.350 2419.515 2052.365 ;
        RECT 2434.240 2052.350 2435.840 2052.365 ;
        RECT 2368.940 2052.285 2370.710 2052.350 ;
        RECT 2385.265 2052.285 2387.035 2052.350 ;
        RECT 2401.590 2052.285 2403.360 2052.350 ;
        RECT 2417.915 2052.285 2419.685 2052.350 ;
        RECT 2434.240 2052.285 2436.010 2052.350 ;
        RECT 2368.940 2052.265 2370.750 2052.285 ;
        RECT 2385.265 2052.265 2387.075 2052.285 ;
        RECT 2401.590 2052.265 2403.400 2052.285 ;
        RECT 2417.915 2052.265 2419.725 2052.285 ;
        RECT 2434.240 2052.265 2436.050 2052.285 ;
        RECT 2368.610 2052.240 2370.860 2052.265 ;
        RECT 2384.935 2052.240 2387.185 2052.265 ;
        RECT 2401.260 2052.240 2403.510 2052.265 ;
        RECT 2417.585 2052.240 2419.835 2052.265 ;
        RECT 2433.910 2052.240 2436.160 2052.265 ;
        RECT 2368.610 2052.225 2371.355 2052.240 ;
        RECT 2368.610 2052.085 2369.080 2052.225 ;
        RECT 2370.400 2052.085 2371.355 2052.225 ;
        RECT 2368.610 2052.035 2368.900 2052.085 ;
        RECT 2370.430 2052.055 2371.355 2052.085 ;
        RECT 2370.430 2052.035 2370.860 2052.055 ;
        RECT 2370.430 2052.025 2370.750 2052.035 ;
        RECT 2371.170 2050.905 2371.355 2052.055 ;
        RECT 2384.935 2052.225 2387.680 2052.240 ;
        RECT 2384.935 2052.085 2385.405 2052.225 ;
        RECT 2386.725 2052.085 2387.680 2052.225 ;
        RECT 2384.935 2052.035 2385.225 2052.085 ;
        RECT 2386.755 2052.055 2387.680 2052.085 ;
        RECT 2386.755 2052.035 2387.185 2052.055 ;
        RECT 2386.755 2052.025 2387.075 2052.035 ;
        RECT 2387.495 2050.905 2387.680 2052.055 ;
        RECT 2401.260 2052.225 2404.005 2052.240 ;
        RECT 2401.260 2052.085 2401.730 2052.225 ;
        RECT 2403.050 2052.085 2404.005 2052.225 ;
        RECT 2401.260 2052.035 2401.550 2052.085 ;
        RECT 2403.080 2052.055 2404.005 2052.085 ;
        RECT 2403.080 2052.035 2403.510 2052.055 ;
        RECT 2403.080 2052.025 2403.400 2052.035 ;
        RECT 2403.820 2050.905 2404.005 2052.055 ;
        RECT 2417.585 2052.225 2420.330 2052.240 ;
        RECT 2417.585 2052.085 2418.055 2052.225 ;
        RECT 2419.375 2052.085 2420.330 2052.225 ;
        RECT 2417.585 2052.035 2417.875 2052.085 ;
        RECT 2419.405 2052.055 2420.330 2052.085 ;
        RECT 2419.405 2052.035 2419.835 2052.055 ;
        RECT 2419.405 2052.025 2419.725 2052.035 ;
        RECT 2420.145 2050.905 2420.330 2052.055 ;
        RECT 2433.910 2052.225 2436.655 2052.240 ;
        RECT 2433.910 2052.085 2434.380 2052.225 ;
        RECT 2435.700 2052.085 2436.655 2052.225 ;
        RECT 2433.910 2052.035 2434.200 2052.085 ;
        RECT 2435.730 2052.055 2436.655 2052.085 ;
        RECT 2435.730 2052.035 2436.160 2052.055 ;
        RECT 2435.730 2052.025 2436.050 2052.035 ;
        RECT 2436.470 2050.905 2436.655 2052.055 ;
        RECT 2361.540 2049.600 2371.355 2050.905 ;
        RECT 2377.865 2049.600 2387.680 2050.905 ;
        RECT 2394.190 2049.600 2404.005 2050.905 ;
        RECT 2410.515 2049.600 2420.330 2050.905 ;
        RECT 2426.840 2049.600 2436.655 2050.905 ;
        RECT 2343.000 2048.000 2442.425 2049.600 ;
        RECT 2695.520 2036.680 2734.960 2037.160 ;
        RECT 2695.520 2031.240 2734.960 2031.720 ;
        RECT 2695.520 2025.800 2734.960 2026.280 ;
        RECT 2695.520 2020.360 2734.960 2020.840 ;
        RECT 2695.520 2014.920 2734.960 2015.400 ;
        RECT 2695.520 2009.480 2734.960 2009.960 ;
        RECT 2695.520 2004.040 2734.960 2004.520 ;
        RECT 2695.520 1998.600 2734.960 1999.080 ;
        RECT 2695.520 1993.160 2734.960 1993.640 ;
        RECT 2695.520 1987.720 2734.960 1988.200 ;
        RECT 2695.520 1982.280 2734.960 1982.760 ;
        RECT 2522.555 1981.785 2534.570 1981.940 ;
        RECT 2522.130 1981.615 2534.570 1981.785 ;
        RECT 2522.555 1981.460 2534.570 1981.615 ;
        RECT 2531.170 1980.340 2534.270 1981.460 ;
        RECT 2695.520 1976.840 2734.960 1977.320 ;
        RECT 2522.555 1974.255 2534.570 1974.410 ;
        RECT 2522.130 1974.085 2534.570 1974.255 ;
        RECT 2522.555 1973.930 2534.570 1974.085 ;
        RECT 2531.170 1972.810 2534.270 1973.930 ;
        RECT 2695.520 1971.400 2734.960 1971.880 ;
        RECT 2522.555 1968.275 2534.570 1968.430 ;
        RECT 2522.130 1968.105 2534.570 1968.275 ;
        RECT 2522.555 1967.950 2534.570 1968.105 ;
        RECT 2531.170 1966.830 2534.270 1967.950 ;
        RECT 2695.520 1965.960 2734.960 1966.440 ;
        RECT 2522.555 1962.330 2534.570 1962.485 ;
        RECT 2522.130 1962.160 2534.570 1962.330 ;
        RECT 2522.555 1962.005 2534.570 1962.160 ;
        RECT 2531.170 1960.885 2534.270 1962.005 ;
        RECT 2695.520 1960.520 2734.960 1961.000 ;
        RECT 2522.555 1956.685 2534.570 1956.840 ;
        RECT 2522.130 1956.515 2534.570 1956.685 ;
        RECT 2522.555 1956.360 2534.570 1956.515 ;
        RECT 2343.005 1953.865 2453.605 1955.465 ;
        RECT 2531.170 1955.240 2534.270 1956.360 ;
        RECT 2695.520 1955.080 2734.960 1955.560 ;
        RECT 2369.550 1951.790 2369.720 1953.865 ;
        RECT 2369.990 1951.790 2370.280 1951.820 ;
        RECT 2369.550 1951.605 2370.280 1951.790 ;
        RECT 2388.110 1951.790 2388.280 1953.865 ;
        RECT 2388.550 1951.790 2388.840 1951.820 ;
        RECT 2388.110 1951.605 2388.840 1951.790 ;
        RECT 2406.670 1951.790 2406.840 1953.865 ;
        RECT 2407.110 1951.790 2407.400 1951.820 ;
        RECT 2406.670 1951.605 2407.400 1951.790 ;
        RECT 2425.230 1951.790 2425.400 1953.865 ;
        RECT 2425.670 1951.790 2425.960 1951.820 ;
        RECT 2425.230 1951.605 2425.960 1951.790 ;
        RECT 2443.790 1951.790 2443.960 1953.865 ;
        RECT 2444.230 1951.790 2444.520 1951.820 ;
        RECT 2443.790 1951.605 2444.520 1951.790 ;
        RECT 2369.990 1951.590 2370.280 1951.605 ;
        RECT 2388.550 1951.590 2388.840 1951.605 ;
        RECT 2407.110 1951.590 2407.400 1951.605 ;
        RECT 2425.670 1951.590 2425.960 1951.605 ;
        RECT 2444.230 1951.590 2444.520 1951.605 ;
        RECT 2522.555 1950.680 2534.570 1950.835 ;
        RECT 2522.130 1950.510 2534.570 1950.680 ;
        RECT 2522.555 1950.355 2534.570 1950.510 ;
        RECT 2531.170 1949.235 2534.270 1950.355 ;
        RECT 2695.520 1949.640 2734.960 1950.120 ;
        RECT 2363.235 1947.305 2363.555 1947.565 ;
        RECT 2381.795 1947.305 2382.115 1947.565 ;
        RECT 2400.355 1947.305 2400.675 1947.565 ;
        RECT 2418.915 1947.305 2419.235 1947.565 ;
        RECT 2437.475 1947.305 2437.795 1947.565 ;
        RECT 2364.975 1946.805 2365.265 1947.035 ;
        RECT 2383.535 1946.805 2383.825 1947.035 ;
        RECT 2402.095 1946.805 2402.385 1947.035 ;
        RECT 2420.655 1946.805 2420.945 1947.035 ;
        RECT 2439.215 1946.805 2439.505 1947.035 ;
        RECT 2364.205 1946.665 2365.265 1946.805 ;
        RECT 2382.765 1946.665 2383.825 1946.805 ;
        RECT 2401.325 1946.665 2402.385 1946.805 ;
        RECT 2419.885 1946.665 2420.945 1946.805 ;
        RECT 2438.445 1946.665 2439.505 1946.805 ;
        RECT 2361.545 1944.600 2373.590 1945.905 ;
        RECT 2380.105 1944.600 2392.150 1945.905 ;
        RECT 2398.665 1944.600 2410.710 1945.905 ;
        RECT 2417.225 1944.600 2429.270 1945.905 ;
        RECT 2435.785 1944.600 2447.830 1945.905 ;
        RECT 2343.005 1943.000 2453.605 1944.600 ;
        RECT 2882.000 1891.670 2894.380 1891.825 ;
        RECT 2881.575 1891.500 2894.380 1891.670 ;
        RECT 2882.000 1891.345 2894.380 1891.500 ;
        RECT 2891.170 1890.090 2894.270 1891.345 ;
        RECT 2695.520 1856.680 2734.960 1857.160 ;
        RECT 2695.520 1851.240 2734.960 1851.720 ;
        RECT 2695.520 1845.800 2734.960 1846.280 ;
        RECT 2695.520 1840.360 2734.960 1840.840 ;
        RECT 2695.520 1834.920 2734.960 1835.400 ;
        RECT 2695.520 1829.480 2734.960 1829.960 ;
        RECT 2695.520 1824.040 2734.960 1824.520 ;
        RECT 2695.520 1818.600 2734.960 1819.080 ;
        RECT 2695.520 1813.160 2734.960 1813.640 ;
        RECT 2695.520 1807.720 2734.960 1808.200 ;
        RECT 2522.555 1804.815 2534.570 1804.970 ;
        RECT 2522.130 1804.645 2534.570 1804.815 ;
        RECT 2522.555 1804.490 2534.570 1804.645 ;
        RECT 2531.170 1803.370 2534.270 1804.490 ;
        RECT 2695.520 1802.280 2734.960 1802.760 ;
        RECT 2522.555 1797.285 2534.570 1797.440 ;
        RECT 2522.130 1797.115 2534.570 1797.285 ;
        RECT 2522.555 1796.960 2534.570 1797.115 ;
        RECT 2531.170 1795.840 2534.270 1796.960 ;
        RECT 2695.520 1796.840 2734.960 1797.320 ;
        RECT 2343.000 1790.865 2447.045 1792.465 ;
        RECT 2522.555 1791.305 2534.570 1791.460 ;
        RECT 2695.520 1791.400 2734.960 1791.880 ;
        RECT 2522.130 1791.135 2534.570 1791.305 ;
        RECT 2522.555 1790.980 2534.570 1791.135 ;
        RECT 2376.465 1788.820 2376.635 1790.865 ;
        RECT 2391.725 1788.820 2391.895 1790.865 ;
        RECT 2406.985 1788.820 2407.155 1790.865 ;
        RECT 2422.245 1788.820 2422.415 1790.865 ;
        RECT 2437.505 1788.820 2437.675 1790.865 ;
        RECT 2531.170 1789.860 2534.270 1790.980 ;
        RECT 2376.465 1788.790 2376.925 1788.820 ;
        RECT 2391.725 1788.790 2392.185 1788.820 ;
        RECT 2406.985 1788.790 2407.445 1788.820 ;
        RECT 2422.245 1788.790 2422.705 1788.820 ;
        RECT 2437.505 1788.790 2437.965 1788.820 ;
        RECT 2376.460 1788.620 2376.925 1788.790 ;
        RECT 2391.720 1788.620 2392.185 1788.790 ;
        RECT 2406.980 1788.620 2407.445 1788.790 ;
        RECT 2422.240 1788.620 2422.705 1788.790 ;
        RECT 2437.500 1788.620 2437.965 1788.790 ;
        RECT 2376.465 1788.605 2376.925 1788.620 ;
        RECT 2391.725 1788.605 2392.185 1788.620 ;
        RECT 2406.985 1788.605 2407.445 1788.620 ;
        RECT 2422.245 1788.605 2422.705 1788.620 ;
        RECT 2437.505 1788.605 2437.965 1788.620 ;
        RECT 2376.635 1788.590 2376.925 1788.605 ;
        RECT 2391.895 1788.590 2392.185 1788.605 ;
        RECT 2407.155 1788.590 2407.445 1788.605 ;
        RECT 2422.415 1788.590 2422.705 1788.605 ;
        RECT 2437.675 1788.590 2437.965 1788.605 ;
        RECT 2695.520 1785.960 2734.960 1786.440 ;
        RECT 2522.555 1785.360 2534.570 1785.515 ;
        RECT 2522.130 1785.190 2534.570 1785.360 ;
        RECT 2522.555 1785.035 2534.570 1785.190 ;
        RECT 2371.985 1784.035 2372.275 1784.265 ;
        RECT 2387.245 1784.035 2387.535 1784.265 ;
        RECT 2402.505 1784.035 2402.795 1784.265 ;
        RECT 2417.765 1784.035 2418.055 1784.265 ;
        RECT 2433.025 1784.035 2433.315 1784.265 ;
        RECT 2372.055 1783.805 2372.195 1784.035 ;
        RECT 2387.315 1783.805 2387.455 1784.035 ;
        RECT 2402.575 1783.805 2402.715 1784.035 ;
        RECT 2417.835 1783.805 2417.975 1784.035 ;
        RECT 2433.095 1783.805 2433.235 1784.035 ;
        RECT 2531.170 1783.915 2534.270 1785.035 ;
        RECT 2372.055 1783.665 2372.675 1783.805 ;
        RECT 2387.315 1783.665 2387.935 1783.805 ;
        RECT 2402.575 1783.665 2403.195 1783.805 ;
        RECT 2417.835 1783.665 2418.455 1783.805 ;
        RECT 2433.095 1783.665 2433.715 1783.805 ;
        RECT 2372.535 1783.505 2372.675 1783.665 ;
        RECT 2387.795 1783.505 2387.935 1783.665 ;
        RECT 2403.055 1783.505 2403.195 1783.665 ;
        RECT 2418.315 1783.505 2418.455 1783.665 ;
        RECT 2433.575 1783.505 2433.715 1783.665 ;
        RECT 2372.295 1783.445 2372.675 1783.505 ;
        RECT 2387.555 1783.445 2387.935 1783.505 ;
        RECT 2402.815 1783.445 2403.195 1783.505 ;
        RECT 2418.075 1783.445 2418.455 1783.505 ;
        RECT 2433.335 1783.445 2433.715 1783.505 ;
        RECT 2372.295 1783.385 2372.885 1783.445 ;
        RECT 2373.185 1783.385 2373.475 1783.425 ;
        RECT 2372.295 1783.245 2373.475 1783.385 ;
        RECT 2387.555 1783.385 2388.145 1783.445 ;
        RECT 2388.445 1783.385 2388.735 1783.425 ;
        RECT 2387.555 1783.245 2388.735 1783.385 ;
        RECT 2402.815 1783.385 2403.405 1783.445 ;
        RECT 2403.705 1783.385 2403.995 1783.425 ;
        RECT 2402.815 1783.245 2403.995 1783.385 ;
        RECT 2418.075 1783.385 2418.665 1783.445 ;
        RECT 2418.965 1783.385 2419.255 1783.425 ;
        RECT 2418.075 1783.245 2419.255 1783.385 ;
        RECT 2433.335 1783.385 2433.925 1783.445 ;
        RECT 2434.225 1783.385 2434.515 1783.425 ;
        RECT 2433.335 1783.245 2434.515 1783.385 ;
        RECT 2372.480 1783.185 2372.885 1783.245 ;
        RECT 2373.185 1783.195 2373.475 1783.245 ;
        RECT 2387.740 1783.185 2388.145 1783.245 ;
        RECT 2388.445 1783.195 2388.735 1783.245 ;
        RECT 2403.000 1783.185 2403.405 1783.245 ;
        RECT 2403.705 1783.195 2403.995 1783.245 ;
        RECT 2418.260 1783.185 2418.665 1783.245 ;
        RECT 2418.965 1783.195 2419.255 1783.245 ;
        RECT 2433.520 1783.185 2433.925 1783.245 ;
        RECT 2434.225 1783.195 2434.515 1783.245 ;
        RECT 2372.480 1782.915 2372.770 1783.185 ;
        RECT 2380.040 1782.915 2380.235 1782.920 ;
        RECT 2387.740 1782.915 2388.030 1783.185 ;
        RECT 2395.300 1782.915 2395.495 1782.920 ;
        RECT 2403.000 1782.915 2403.290 1783.185 ;
        RECT 2410.560 1782.915 2410.755 1782.920 ;
        RECT 2418.260 1782.915 2418.550 1783.185 ;
        RECT 2425.820 1782.915 2426.015 1782.920 ;
        RECT 2433.520 1782.915 2433.810 1783.185 ;
        RECT 2441.080 1782.915 2441.275 1782.920 ;
        RECT 2371.495 1781.600 2380.235 1782.915 ;
        RECT 2386.755 1781.600 2395.495 1782.915 ;
        RECT 2402.015 1781.600 2410.755 1782.915 ;
        RECT 2417.275 1781.600 2426.015 1782.915 ;
        RECT 2432.535 1781.600 2441.275 1782.915 ;
        RECT 2343.000 1780.000 2447.045 1781.600 ;
        RECT 2695.520 1780.520 2734.960 1781.000 ;
        RECT 2522.555 1779.715 2534.570 1779.870 ;
        RECT 2522.130 1779.545 2534.570 1779.715 ;
        RECT 2522.555 1779.390 2534.570 1779.545 ;
        RECT 2531.170 1778.270 2534.270 1779.390 ;
        RECT 2695.520 1775.080 2734.960 1775.560 ;
        RECT 2695.520 1769.640 2734.960 1770.120 ;
        RECT 2522.555 1768.245 2534.570 1768.400 ;
        RECT 2522.130 1768.075 2534.570 1768.245 ;
        RECT 2522.555 1767.920 2534.570 1768.075 ;
        RECT 2531.170 1766.800 2534.270 1767.920 ;
        RECT 2410.920 1712.465 2444.085 1712.470 ;
        RECT 2394.335 1712.460 2444.085 1712.465 ;
        RECT 2343.000 1710.860 2444.085 1712.460 ;
        RECT 2358.415 1710.855 2361.165 1710.860 ;
        RECT 2361.645 1710.855 2365.170 1710.860 ;
        RECT 2362.605 1710.850 2362.780 1710.855 ;
        RECT 2362.605 1708.805 2362.775 1710.850 ;
        RECT 2362.605 1708.775 2363.060 1708.805 ;
        RECT 2362.595 1708.605 2363.060 1708.775 ;
        RECT 2364.880 1708.685 2365.170 1710.855 ;
        RECT 2365.450 1708.685 2365.730 1710.860 ;
        RECT 2366.010 1708.685 2366.290 1710.860 ;
        RECT 2366.570 1708.685 2366.850 1710.860 ;
        RECT 2367.130 1708.685 2367.410 1710.860 ;
        RECT 2367.690 1708.685 2367.970 1710.860 ;
        RECT 2368.250 1708.685 2368.530 1710.860 ;
        RECT 2368.810 1708.685 2369.090 1710.860 ;
        RECT 2369.370 1708.685 2369.650 1710.860 ;
        RECT 2369.930 1708.685 2370.210 1710.860 ;
        RECT 2370.490 1708.685 2370.770 1710.860 ;
        RECT 2371.050 1708.685 2371.330 1710.860 ;
        RECT 2371.610 1708.685 2371.785 1710.860 ;
        RECT 2378.230 1710.855 2381.755 1710.860 ;
        RECT 2379.190 1710.850 2379.365 1710.855 ;
        RECT 2379.190 1708.805 2379.360 1710.850 ;
        RECT 2379.190 1708.775 2379.645 1708.805 ;
        RECT 2362.605 1708.600 2363.060 1708.605 ;
        RECT 2362.770 1708.575 2363.060 1708.600 ;
        RECT 2364.740 1708.325 2371.785 1708.685 ;
        RECT 2379.180 1708.605 2379.645 1708.775 ;
        RECT 2381.465 1708.685 2381.755 1710.855 ;
        RECT 2382.035 1708.685 2382.315 1710.860 ;
        RECT 2382.595 1708.685 2382.875 1710.860 ;
        RECT 2383.155 1708.685 2383.435 1710.860 ;
        RECT 2383.715 1708.685 2383.995 1710.860 ;
        RECT 2384.275 1708.685 2384.555 1710.860 ;
        RECT 2384.835 1708.685 2385.115 1710.860 ;
        RECT 2385.395 1708.685 2385.675 1710.860 ;
        RECT 2385.955 1708.685 2386.235 1710.860 ;
        RECT 2386.515 1708.685 2386.795 1710.860 ;
        RECT 2387.075 1708.685 2387.355 1710.860 ;
        RECT 2387.635 1708.685 2387.915 1710.860 ;
        RECT 2388.195 1708.685 2388.370 1710.860 ;
        RECT 2395.775 1710.855 2395.950 1710.860 ;
        RECT 2395.775 1708.810 2395.945 1710.855 ;
        RECT 2395.775 1708.780 2396.230 1708.810 ;
        RECT 2379.190 1708.600 2379.645 1708.605 ;
        RECT 2379.355 1708.575 2379.645 1708.600 ;
        RECT 2381.325 1708.325 2388.370 1708.685 ;
        RECT 2395.765 1708.610 2396.230 1708.780 ;
        RECT 2398.050 1708.690 2398.340 1710.860 ;
        RECT 2398.620 1708.690 2398.900 1710.860 ;
        RECT 2399.180 1708.690 2399.460 1710.860 ;
        RECT 2399.740 1708.690 2400.020 1710.860 ;
        RECT 2400.300 1708.690 2400.580 1710.860 ;
        RECT 2400.860 1708.690 2401.140 1710.860 ;
        RECT 2401.420 1708.690 2401.700 1710.860 ;
        RECT 2401.980 1708.690 2402.260 1710.860 ;
        RECT 2402.540 1708.690 2402.820 1710.860 ;
        RECT 2403.100 1708.690 2403.380 1710.860 ;
        RECT 2403.660 1708.690 2403.940 1710.860 ;
        RECT 2404.220 1708.690 2404.500 1710.860 ;
        RECT 2404.780 1708.690 2404.955 1710.860 ;
        RECT 2412.360 1708.815 2412.530 1710.860 ;
        RECT 2412.360 1708.785 2412.815 1708.815 ;
        RECT 2395.775 1708.605 2396.230 1708.610 ;
        RECT 2395.940 1708.580 2396.230 1708.605 ;
        RECT 2397.910 1708.330 2404.955 1708.690 ;
        RECT 2412.350 1708.615 2412.815 1708.785 ;
        RECT 2414.635 1708.695 2414.925 1710.860 ;
        RECT 2415.205 1708.695 2415.485 1710.860 ;
        RECT 2415.765 1708.695 2416.045 1710.860 ;
        RECT 2416.325 1708.695 2416.605 1710.860 ;
        RECT 2416.885 1708.695 2417.165 1710.860 ;
        RECT 2417.445 1708.695 2417.725 1710.860 ;
        RECT 2418.005 1708.695 2418.285 1710.860 ;
        RECT 2418.565 1708.695 2418.845 1710.860 ;
        RECT 2419.125 1708.695 2419.405 1710.860 ;
        RECT 2419.685 1708.695 2419.965 1710.860 ;
        RECT 2420.245 1708.695 2420.525 1710.860 ;
        RECT 2420.805 1708.695 2421.085 1710.860 ;
        RECT 2421.365 1708.695 2421.540 1710.860 ;
        RECT 2428.940 1708.815 2429.110 1710.860 ;
        RECT 2428.940 1708.785 2429.395 1708.815 ;
        RECT 2412.360 1708.610 2412.815 1708.615 ;
        RECT 2412.525 1708.585 2412.815 1708.610 ;
        RECT 2414.495 1708.335 2421.540 1708.695 ;
        RECT 2428.930 1708.615 2429.395 1708.785 ;
        RECT 2431.215 1708.695 2431.505 1710.860 ;
        RECT 2431.785 1708.695 2432.065 1710.860 ;
        RECT 2432.345 1708.695 2432.625 1710.860 ;
        RECT 2432.905 1708.695 2433.185 1710.860 ;
        RECT 2433.465 1708.695 2433.745 1710.860 ;
        RECT 2434.025 1708.695 2434.305 1710.860 ;
        RECT 2434.585 1708.695 2434.865 1710.860 ;
        RECT 2435.145 1708.695 2435.425 1710.860 ;
        RECT 2435.705 1708.695 2435.985 1710.860 ;
        RECT 2436.265 1708.695 2436.545 1710.860 ;
        RECT 2436.825 1708.695 2437.105 1710.860 ;
        RECT 2437.385 1708.695 2437.665 1710.860 ;
        RECT 2437.945 1708.695 2438.120 1710.860 ;
        RECT 2428.940 1708.610 2429.395 1708.615 ;
        RECT 2429.105 1708.585 2429.395 1708.610 ;
        RECT 2431.075 1708.335 2438.120 1708.695 ;
        RECT 2367.305 1708.045 2367.565 1708.325 ;
        RECT 2383.890 1708.045 2384.150 1708.325 ;
        RECT 2400.475 1708.050 2400.735 1708.330 ;
        RECT 2417.060 1708.055 2417.320 1708.335 ;
        RECT 2433.640 1708.055 2433.900 1708.335 ;
        RECT 2367.270 1707.945 2367.700 1708.045 ;
        RECT 2383.855 1707.945 2384.285 1708.045 ;
        RECT 2400.440 1707.950 2400.870 1708.050 ;
        RECT 2417.025 1707.955 2417.455 1708.055 ;
        RECT 2433.605 1707.955 2434.035 1708.055 ;
        RECT 2366.340 1707.805 2368.690 1707.945 ;
        RECT 2366.340 1707.365 2366.480 1707.805 ;
        RECT 2367.280 1707.775 2367.560 1707.805 ;
        RECT 2367.300 1707.745 2367.560 1707.775 ;
        RECT 2368.550 1707.365 2368.690 1707.805 ;
        RECT 2382.925 1707.805 2385.275 1707.945 ;
        RECT 2382.925 1707.365 2383.065 1707.805 ;
        RECT 2383.865 1707.775 2384.145 1707.805 ;
        RECT 2383.885 1707.745 2384.145 1707.775 ;
        RECT 2385.135 1707.365 2385.275 1707.805 ;
        RECT 2399.510 1707.810 2401.860 1707.950 ;
        RECT 2399.510 1707.370 2399.650 1707.810 ;
        RECT 2400.450 1707.780 2400.730 1707.810 ;
        RECT 2400.470 1707.750 2400.730 1707.780 ;
        RECT 2401.720 1707.370 2401.860 1707.810 ;
        RECT 2416.095 1707.815 2418.445 1707.955 ;
        RECT 2416.095 1707.375 2416.235 1707.815 ;
        RECT 2417.035 1707.785 2417.315 1707.815 ;
        RECT 2417.055 1707.755 2417.315 1707.785 ;
        RECT 2418.305 1707.375 2418.445 1707.815 ;
        RECT 2432.675 1707.815 2435.025 1707.955 ;
        RECT 2432.675 1707.375 2432.815 1707.815 ;
        RECT 2433.615 1707.785 2433.895 1707.815 ;
        RECT 2433.635 1707.755 2433.895 1707.785 ;
        RECT 2434.885 1707.375 2435.025 1707.815 ;
        RECT 2366.260 1707.135 2366.550 1707.365 ;
        RECT 2368.470 1707.135 2368.760 1707.365 ;
        RECT 2382.845 1707.135 2383.135 1707.365 ;
        RECT 2385.055 1707.135 2385.345 1707.365 ;
        RECT 2399.430 1707.140 2399.720 1707.370 ;
        RECT 2401.640 1707.140 2401.930 1707.370 ;
        RECT 2416.015 1707.145 2416.305 1707.375 ;
        RECT 2418.225 1707.145 2418.515 1707.375 ;
        RECT 2432.595 1707.145 2432.885 1707.375 ;
        RECT 2434.805 1707.145 2435.095 1707.375 ;
        RECT 2364.580 1702.765 2371.970 1703.125 ;
        RECT 2381.165 1702.765 2388.555 1703.125 ;
        RECT 2397.750 1702.770 2405.140 1703.130 ;
        RECT 2414.335 1702.775 2421.725 1703.135 ;
        RECT 2430.915 1702.775 2438.305 1703.135 ;
        RECT 2364.625 1701.605 2364.920 1702.765 ;
        RECT 2365.210 1701.605 2365.500 1702.765 ;
        RECT 2365.790 1701.605 2366.080 1702.765 ;
        RECT 2366.370 1701.605 2366.660 1702.765 ;
        RECT 2366.950 1701.605 2367.240 1702.765 ;
        RECT 2367.530 1701.605 2367.815 1702.765 ;
        RECT 2368.105 1701.605 2368.395 1702.765 ;
        RECT 2368.685 1701.605 2368.975 1702.765 ;
        RECT 2369.265 1701.605 2369.555 1702.765 ;
        RECT 2369.845 1701.605 2370.130 1702.765 ;
        RECT 2370.420 1701.605 2370.710 1702.765 ;
        RECT 2371.000 1701.605 2371.290 1702.765 ;
        RECT 2371.580 1701.605 2371.970 1702.765 ;
        RECT 2364.625 1701.600 2371.970 1701.605 ;
        RECT 2381.210 1701.605 2381.505 1702.765 ;
        RECT 2381.795 1701.605 2382.085 1702.765 ;
        RECT 2382.375 1701.605 2382.665 1702.765 ;
        RECT 2382.955 1701.605 2383.245 1702.765 ;
        RECT 2383.535 1701.605 2383.825 1702.765 ;
        RECT 2384.115 1701.605 2384.400 1702.765 ;
        RECT 2384.690 1701.605 2384.980 1702.765 ;
        RECT 2385.270 1701.605 2385.560 1702.765 ;
        RECT 2385.850 1701.605 2386.140 1702.765 ;
        RECT 2386.430 1701.605 2386.715 1702.765 ;
        RECT 2387.005 1701.605 2387.295 1702.765 ;
        RECT 2387.585 1701.605 2387.875 1702.765 ;
        RECT 2388.165 1701.605 2388.555 1702.765 ;
        RECT 2397.795 1701.610 2398.090 1702.770 ;
        RECT 2398.380 1701.610 2398.670 1702.770 ;
        RECT 2398.960 1701.610 2399.250 1702.770 ;
        RECT 2399.540 1701.610 2399.830 1702.770 ;
        RECT 2400.120 1701.610 2400.410 1702.770 ;
        RECT 2400.700 1701.610 2400.985 1702.770 ;
        RECT 2401.275 1701.610 2401.565 1702.770 ;
        RECT 2401.855 1701.610 2402.145 1702.770 ;
        RECT 2402.435 1701.610 2402.725 1702.770 ;
        RECT 2403.015 1701.610 2403.300 1702.770 ;
        RECT 2403.590 1701.610 2403.880 1702.770 ;
        RECT 2404.170 1701.610 2404.460 1702.770 ;
        RECT 2404.750 1701.610 2405.140 1702.770 ;
        RECT 2414.380 1701.615 2414.675 1702.775 ;
        RECT 2414.965 1701.615 2415.255 1702.775 ;
        RECT 2415.545 1701.615 2415.835 1702.775 ;
        RECT 2416.125 1701.615 2416.415 1702.775 ;
        RECT 2416.705 1701.615 2416.995 1702.775 ;
        RECT 2417.285 1701.615 2417.570 1702.775 ;
        RECT 2417.860 1701.615 2418.150 1702.775 ;
        RECT 2418.440 1701.615 2418.730 1702.775 ;
        RECT 2419.020 1701.615 2419.310 1702.775 ;
        RECT 2419.600 1701.615 2419.885 1702.775 ;
        RECT 2420.175 1701.615 2420.465 1702.775 ;
        RECT 2420.755 1701.615 2421.045 1702.775 ;
        RECT 2421.335 1701.615 2421.725 1702.775 ;
        RECT 2414.380 1701.610 2421.725 1701.615 ;
        RECT 2430.960 1701.615 2431.255 1702.775 ;
        RECT 2431.545 1701.615 2431.835 1702.775 ;
        RECT 2432.125 1701.615 2432.415 1702.775 ;
        RECT 2432.705 1701.615 2432.995 1702.775 ;
        RECT 2433.285 1701.615 2433.575 1702.775 ;
        RECT 2433.865 1701.615 2434.150 1702.775 ;
        RECT 2434.440 1701.615 2434.730 1702.775 ;
        RECT 2435.020 1701.615 2435.310 1702.775 ;
        RECT 2435.600 1701.615 2435.890 1702.775 ;
        RECT 2436.180 1701.615 2436.465 1702.775 ;
        RECT 2436.755 1701.615 2437.045 1702.775 ;
        RECT 2437.335 1701.615 2437.625 1702.775 ;
        RECT 2437.915 1701.615 2438.305 1702.775 ;
        RECT 2430.960 1701.610 2438.305 1701.615 ;
        RECT 2397.795 1701.605 2405.140 1701.610 ;
        RECT 2410.920 1701.605 2444.085 1701.610 ;
        RECT 2381.210 1701.600 2388.555 1701.605 ;
        RECT 2394.335 1701.600 2444.085 1701.605 ;
        RECT 2343.000 1700.000 2444.085 1701.600 ;
        RECT 2695.520 1676.680 2734.960 1677.160 ;
        RECT 2695.520 1671.240 2734.960 1671.720 ;
        RECT 2695.520 1665.800 2734.960 1666.280 ;
        RECT 2695.520 1660.360 2734.960 1660.840 ;
        RECT 2695.520 1654.920 2734.960 1655.400 ;
        RECT 2695.520 1649.480 2734.960 1649.960 ;
        RECT 2695.520 1644.040 2734.960 1644.520 ;
        RECT 2695.520 1638.600 2734.960 1639.080 ;
        RECT 2695.520 1633.160 2734.960 1633.640 ;
        RECT 2695.520 1627.720 2734.960 1628.200 ;
        RECT 2882.000 1625.790 2894.380 1625.945 ;
        RECT 2881.575 1625.620 2894.380 1625.790 ;
        RECT 2882.000 1625.465 2894.380 1625.620 ;
        RECT 2891.170 1624.210 2894.270 1625.465 ;
        RECT 2522.555 1623.680 2534.570 1623.835 ;
        RECT 2522.130 1623.510 2534.570 1623.680 ;
        RECT 2522.555 1623.355 2534.570 1623.510 ;
        RECT 2531.170 1622.235 2534.270 1623.355 ;
        RECT 2695.520 1622.280 2734.960 1622.760 ;
        RECT 2522.555 1617.265 2534.570 1617.420 ;
        RECT 2522.130 1617.095 2534.570 1617.265 ;
        RECT 2522.555 1616.940 2534.570 1617.095 ;
        RECT 2531.170 1615.820 2534.270 1616.940 ;
        RECT 2695.520 1616.840 2734.960 1617.320 ;
        RECT 2395.235 1612.460 2412.475 1612.465 ;
        RECT 2343.045 1610.860 2446.915 1612.460 ;
        RECT 2695.520 1611.400 2734.960 1611.880 ;
        RECT 2362.175 1608.785 2362.345 1610.860 ;
        RECT 2362.580 1608.785 2362.870 1608.815 ;
        RECT 2362.175 1608.600 2362.870 1608.785 ;
        RECT 2362.580 1608.585 2362.870 1608.600 ;
        RECT 2364.585 1608.685 2364.910 1610.860 ;
        RECT 2365.235 1608.685 2365.560 1610.860 ;
        RECT 2365.885 1608.685 2366.210 1610.860 ;
        RECT 2366.535 1608.685 2366.860 1610.860 ;
        RECT 2367.185 1608.685 2367.510 1610.860 ;
        RECT 2367.835 1608.685 2368.160 1610.860 ;
        RECT 2368.485 1608.685 2368.810 1610.860 ;
        RECT 2369.135 1608.685 2369.460 1610.860 ;
        RECT 2369.785 1608.685 2370.110 1610.860 ;
        RECT 2370.435 1608.685 2370.760 1610.860 ;
        RECT 2371.085 1608.685 2371.410 1610.860 ;
        RECT 2371.735 1608.685 2371.945 1610.860 ;
        RECT 2364.585 1608.330 2371.945 1608.685 ;
        RECT 2379.395 1608.785 2379.565 1610.860 ;
        RECT 2379.800 1608.785 2380.090 1608.815 ;
        RECT 2379.395 1608.600 2380.090 1608.785 ;
        RECT 2379.800 1608.585 2380.090 1608.600 ;
        RECT 2381.805 1608.685 2382.130 1610.860 ;
        RECT 2382.455 1608.685 2382.780 1610.860 ;
        RECT 2383.105 1608.685 2383.430 1610.860 ;
        RECT 2383.755 1608.685 2384.080 1610.860 ;
        RECT 2384.405 1608.685 2384.730 1610.860 ;
        RECT 2385.055 1608.685 2385.380 1610.860 ;
        RECT 2385.705 1608.685 2386.030 1610.860 ;
        RECT 2386.355 1608.685 2386.680 1610.860 ;
        RECT 2387.005 1608.685 2387.330 1610.860 ;
        RECT 2387.655 1608.685 2387.980 1610.860 ;
        RECT 2388.305 1608.685 2388.630 1610.860 ;
        RECT 2388.955 1608.685 2389.165 1610.860 ;
        RECT 2381.805 1608.330 2389.165 1608.685 ;
        RECT 2396.615 1608.790 2396.785 1610.860 ;
        RECT 2397.020 1608.790 2397.310 1608.820 ;
        RECT 2396.615 1608.605 2397.310 1608.790 ;
        RECT 2397.020 1608.590 2397.310 1608.605 ;
        RECT 2399.025 1608.690 2399.350 1610.860 ;
        RECT 2399.675 1608.690 2400.000 1610.860 ;
        RECT 2400.325 1608.690 2400.650 1610.860 ;
        RECT 2400.975 1608.690 2401.300 1610.860 ;
        RECT 2401.625 1608.690 2401.950 1610.860 ;
        RECT 2402.275 1608.690 2402.600 1610.860 ;
        RECT 2402.925 1608.690 2403.250 1610.860 ;
        RECT 2403.575 1608.690 2403.900 1610.860 ;
        RECT 2404.225 1608.690 2404.550 1610.860 ;
        RECT 2404.875 1608.690 2405.200 1610.860 ;
        RECT 2405.525 1608.690 2405.850 1610.860 ;
        RECT 2406.175 1608.690 2406.385 1610.860 ;
        RECT 2399.025 1608.335 2406.385 1608.690 ;
        RECT 2413.835 1608.785 2414.005 1610.860 ;
        RECT 2414.240 1608.785 2414.530 1608.815 ;
        RECT 2413.835 1608.600 2414.530 1608.785 ;
        RECT 2414.240 1608.585 2414.530 1608.600 ;
        RECT 2416.245 1608.685 2416.570 1610.860 ;
        RECT 2416.895 1608.685 2417.220 1610.860 ;
        RECT 2417.545 1608.685 2417.870 1610.860 ;
        RECT 2418.195 1608.685 2418.520 1610.860 ;
        RECT 2418.845 1608.685 2419.170 1610.860 ;
        RECT 2419.495 1608.685 2419.820 1610.860 ;
        RECT 2420.145 1608.685 2420.470 1610.860 ;
        RECT 2420.795 1608.685 2421.120 1610.860 ;
        RECT 2421.445 1608.685 2421.770 1610.860 ;
        RECT 2422.095 1608.685 2422.420 1610.860 ;
        RECT 2422.745 1608.685 2423.070 1610.860 ;
        RECT 2423.395 1608.685 2423.605 1610.860 ;
        RECT 2416.245 1608.330 2423.605 1608.685 ;
        RECT 2431.055 1608.785 2431.225 1610.860 ;
        RECT 2431.460 1608.785 2431.750 1608.815 ;
        RECT 2431.055 1608.600 2431.750 1608.785 ;
        RECT 2431.460 1608.585 2431.750 1608.600 ;
        RECT 2433.465 1608.685 2433.790 1610.860 ;
        RECT 2434.115 1608.685 2434.440 1610.860 ;
        RECT 2434.765 1608.685 2435.090 1610.860 ;
        RECT 2435.415 1608.685 2435.740 1610.860 ;
        RECT 2436.065 1608.685 2436.390 1610.860 ;
        RECT 2436.715 1608.685 2437.040 1610.860 ;
        RECT 2437.365 1608.685 2437.690 1610.860 ;
        RECT 2438.015 1608.685 2438.340 1610.860 ;
        RECT 2438.665 1608.685 2438.990 1610.860 ;
        RECT 2439.315 1608.685 2439.640 1610.860 ;
        RECT 2439.965 1608.685 2440.290 1610.860 ;
        RECT 2440.615 1608.685 2440.825 1610.860 ;
        RECT 2433.465 1608.330 2440.825 1608.685 ;
        RECT 2364.610 1607.325 2364.900 1607.370 ;
        RECT 2366.975 1607.325 2367.295 1607.385 ;
        RECT 2364.610 1607.185 2367.295 1607.325 ;
        RECT 2364.610 1607.140 2364.900 1607.185 ;
        RECT 2366.975 1607.125 2367.295 1607.185 ;
        RECT 2381.830 1607.325 2382.120 1607.370 ;
        RECT 2384.195 1607.325 2384.515 1607.385 ;
        RECT 2381.830 1607.185 2384.515 1607.325 ;
        RECT 2381.830 1607.140 2382.120 1607.185 ;
        RECT 2384.195 1607.125 2384.515 1607.185 ;
        RECT 2399.050 1607.330 2399.340 1607.375 ;
        RECT 2401.415 1607.330 2401.735 1607.390 ;
        RECT 2399.050 1607.190 2401.735 1607.330 ;
        RECT 2399.050 1607.145 2399.340 1607.190 ;
        RECT 2401.415 1607.130 2401.735 1607.190 ;
        RECT 2416.270 1607.325 2416.560 1607.370 ;
        RECT 2418.635 1607.325 2418.955 1607.385 ;
        RECT 2416.270 1607.185 2418.955 1607.325 ;
        RECT 2416.270 1607.140 2416.560 1607.185 ;
        RECT 2418.635 1607.125 2418.955 1607.185 ;
        RECT 2433.490 1607.325 2433.780 1607.370 ;
        RECT 2435.855 1607.325 2436.175 1607.385 ;
        RECT 2433.490 1607.185 2436.175 1607.325 ;
        RECT 2433.490 1607.140 2433.780 1607.185 ;
        RECT 2435.855 1607.125 2436.175 1607.185 ;
        RECT 2695.520 1605.960 2734.960 1606.440 ;
        RECT 2364.580 1602.765 2372.325 1603.120 ;
        RECT 2364.580 1601.600 2364.925 1602.765 ;
        RECT 2365.270 1601.600 2365.600 1602.765 ;
        RECT 2365.945 1601.605 2366.290 1602.765 ;
        RECT 2366.635 1601.605 2366.980 1602.765 ;
        RECT 2367.325 1601.605 2367.670 1602.765 ;
        RECT 2368.015 1601.605 2368.360 1602.765 ;
        RECT 2368.705 1601.605 2369.050 1602.765 ;
        RECT 2369.395 1601.605 2369.740 1602.765 ;
        RECT 2370.085 1601.605 2370.430 1602.765 ;
        RECT 2370.775 1601.605 2371.120 1602.765 ;
        RECT 2371.465 1601.605 2371.810 1602.765 ;
        RECT 2372.155 1601.605 2372.325 1602.765 ;
        RECT 2365.945 1601.600 2372.325 1601.605 ;
        RECT 2381.800 1602.765 2389.545 1603.120 ;
        RECT 2381.800 1601.600 2382.145 1602.765 ;
        RECT 2382.490 1601.600 2382.820 1602.765 ;
        RECT 2383.165 1601.605 2383.510 1602.765 ;
        RECT 2383.855 1601.605 2384.200 1602.765 ;
        RECT 2384.545 1601.605 2384.890 1602.765 ;
        RECT 2385.235 1601.605 2385.580 1602.765 ;
        RECT 2385.925 1601.605 2386.270 1602.765 ;
        RECT 2386.615 1601.605 2386.960 1602.765 ;
        RECT 2387.305 1601.605 2387.650 1602.765 ;
        RECT 2387.995 1601.605 2388.340 1602.765 ;
        RECT 2388.685 1601.605 2389.030 1602.765 ;
        RECT 2389.375 1601.605 2389.545 1602.765 ;
        RECT 2399.020 1602.770 2406.765 1603.125 ;
        RECT 2399.020 1601.605 2399.365 1602.770 ;
        RECT 2399.710 1601.605 2400.040 1602.770 ;
        RECT 2400.385 1601.610 2400.730 1602.770 ;
        RECT 2401.075 1601.610 2401.420 1602.770 ;
        RECT 2401.765 1601.610 2402.110 1602.770 ;
        RECT 2402.455 1601.610 2402.800 1602.770 ;
        RECT 2403.145 1601.610 2403.490 1602.770 ;
        RECT 2403.835 1601.610 2404.180 1602.770 ;
        RECT 2404.525 1601.610 2404.870 1602.770 ;
        RECT 2405.215 1601.610 2405.560 1602.770 ;
        RECT 2405.905 1601.610 2406.250 1602.770 ;
        RECT 2406.595 1601.610 2406.765 1602.770 ;
        RECT 2400.385 1601.605 2406.765 1601.610 ;
        RECT 2416.240 1602.765 2423.985 1603.120 ;
        RECT 2383.165 1601.600 2389.545 1601.605 ;
        RECT 2395.235 1601.600 2412.475 1601.605 ;
        RECT 2416.240 1601.600 2416.585 1602.765 ;
        RECT 2416.930 1601.600 2417.260 1602.765 ;
        RECT 2417.605 1601.605 2417.950 1602.765 ;
        RECT 2418.295 1601.605 2418.640 1602.765 ;
        RECT 2418.985 1601.605 2419.330 1602.765 ;
        RECT 2419.675 1601.605 2420.020 1602.765 ;
        RECT 2420.365 1601.605 2420.710 1602.765 ;
        RECT 2421.055 1601.605 2421.400 1602.765 ;
        RECT 2421.745 1601.605 2422.090 1602.765 ;
        RECT 2422.435 1601.605 2422.780 1602.765 ;
        RECT 2423.125 1601.605 2423.470 1602.765 ;
        RECT 2423.815 1601.605 2423.985 1602.765 ;
        RECT 2417.605 1601.600 2423.985 1601.605 ;
        RECT 2433.460 1602.765 2441.205 1603.120 ;
        RECT 2433.460 1601.600 2433.805 1602.765 ;
        RECT 2434.150 1601.600 2434.480 1602.765 ;
        RECT 2434.825 1601.605 2435.170 1602.765 ;
        RECT 2435.515 1601.605 2435.860 1602.765 ;
        RECT 2436.205 1601.605 2436.550 1602.765 ;
        RECT 2436.895 1601.605 2437.240 1602.765 ;
        RECT 2437.585 1601.605 2437.930 1602.765 ;
        RECT 2438.275 1601.605 2438.620 1602.765 ;
        RECT 2438.965 1601.605 2439.310 1602.765 ;
        RECT 2439.655 1601.605 2440.000 1602.765 ;
        RECT 2440.345 1601.605 2440.690 1602.765 ;
        RECT 2441.035 1601.605 2441.205 1602.765 ;
        RECT 2434.825 1601.600 2441.205 1601.605 ;
        RECT 2343.045 1600.000 2446.915 1601.600 ;
        RECT 2695.520 1600.520 2734.960 1601.000 ;
        RECT 2695.520 1595.080 2734.960 1595.560 ;
        RECT 2695.520 1589.640 2734.960 1590.120 ;
        RECT 2522.555 1588.020 2534.570 1588.175 ;
        RECT 2522.130 1587.850 2534.570 1588.020 ;
        RECT 2522.555 1587.695 2534.570 1587.850 ;
        RECT 2531.170 1586.575 2534.270 1587.695 ;
        RECT 2522.555 1580.490 2534.570 1580.645 ;
        RECT 2522.130 1580.320 2534.570 1580.490 ;
        RECT 2522.555 1580.165 2534.570 1580.320 ;
        RECT 2531.170 1579.045 2534.270 1580.165 ;
        RECT 2522.555 1574.510 2534.570 1574.665 ;
        RECT 2522.130 1574.340 2534.570 1574.510 ;
        RECT 2522.555 1574.185 2534.570 1574.340 ;
        RECT 2531.170 1573.065 2534.270 1574.185 ;
        RECT 2522.555 1566.095 2534.570 1566.250 ;
        RECT 2522.130 1565.925 2534.570 1566.095 ;
        RECT 2522.555 1565.770 2534.570 1565.925 ;
        RECT 2531.170 1564.650 2534.270 1565.770 ;
        RECT 2343.000 1533.860 2442.425 1535.460 ;
        RECT 2367.370 1531.785 2367.545 1533.860 ;
        RECT 2367.750 1531.785 2368.040 1531.815 ;
        RECT 2367.370 1531.600 2368.040 1531.785 ;
        RECT 2383.695 1531.785 2383.870 1533.860 ;
        RECT 2384.075 1531.785 2384.365 1531.815 ;
        RECT 2383.695 1531.600 2384.365 1531.785 ;
        RECT 2400.020 1531.785 2400.195 1533.860 ;
        RECT 2400.400 1531.785 2400.690 1531.815 ;
        RECT 2400.020 1531.600 2400.690 1531.785 ;
        RECT 2416.345 1531.785 2416.520 1533.860 ;
        RECT 2416.725 1531.785 2417.015 1531.815 ;
        RECT 2416.345 1531.600 2417.015 1531.785 ;
        RECT 2432.670 1531.785 2432.845 1533.860 ;
        RECT 2433.050 1531.785 2433.340 1531.815 ;
        RECT 2432.670 1531.600 2433.340 1531.785 ;
        RECT 2367.750 1531.585 2368.040 1531.600 ;
        RECT 2384.075 1531.585 2384.365 1531.600 ;
        RECT 2400.400 1531.585 2400.690 1531.600 ;
        RECT 2416.725 1531.585 2417.015 1531.600 ;
        RECT 2433.050 1531.585 2433.340 1531.600 ;
        RECT 2370.465 1527.255 2370.705 1527.350 ;
        RECT 2386.790 1527.255 2387.030 1527.350 ;
        RECT 2403.115 1527.255 2403.355 1527.350 ;
        RECT 2419.440 1527.255 2419.680 1527.350 ;
        RECT 2435.765 1527.255 2436.005 1527.350 ;
        RECT 2368.935 1527.240 2370.705 1527.255 ;
        RECT 2385.260 1527.240 2387.030 1527.255 ;
        RECT 2401.585 1527.240 2403.355 1527.255 ;
        RECT 2417.910 1527.240 2419.680 1527.255 ;
        RECT 2434.235 1527.240 2436.005 1527.255 ;
        RECT 2368.935 1527.155 2371.350 1527.240 ;
        RECT 2385.260 1527.155 2387.675 1527.240 ;
        RECT 2401.585 1527.155 2404.000 1527.240 ;
        RECT 2417.910 1527.155 2420.325 1527.240 ;
        RECT 2434.235 1527.155 2436.650 1527.240 ;
        RECT 2368.605 1527.115 2371.350 1527.155 ;
        RECT 2368.605 1526.975 2369.075 1527.115 ;
        RECT 2370.395 1527.055 2371.350 1527.115 ;
        RECT 2370.395 1526.975 2370.855 1527.055 ;
        RECT 2368.605 1526.925 2368.895 1526.975 ;
        RECT 2370.425 1526.925 2370.855 1526.975 ;
        RECT 2370.425 1526.915 2370.745 1526.925 ;
        RECT 2371.165 1525.880 2371.350 1527.055 ;
        RECT 2384.930 1527.115 2387.675 1527.155 ;
        RECT 2384.930 1526.975 2385.400 1527.115 ;
        RECT 2386.720 1527.055 2387.675 1527.115 ;
        RECT 2386.720 1526.975 2387.180 1527.055 ;
        RECT 2384.930 1526.925 2385.220 1526.975 ;
        RECT 2386.750 1526.925 2387.180 1526.975 ;
        RECT 2386.750 1526.915 2387.070 1526.925 ;
        RECT 2387.490 1525.880 2387.675 1527.055 ;
        RECT 2401.255 1527.115 2404.000 1527.155 ;
        RECT 2401.255 1526.975 2401.725 1527.115 ;
        RECT 2403.045 1527.055 2404.000 1527.115 ;
        RECT 2403.045 1526.975 2403.505 1527.055 ;
        RECT 2401.255 1526.925 2401.545 1526.975 ;
        RECT 2403.075 1526.925 2403.505 1526.975 ;
        RECT 2403.075 1526.915 2403.395 1526.925 ;
        RECT 2403.815 1525.880 2404.000 1527.055 ;
        RECT 2417.580 1527.115 2420.325 1527.155 ;
        RECT 2417.580 1526.975 2418.050 1527.115 ;
        RECT 2419.370 1527.055 2420.325 1527.115 ;
        RECT 2419.370 1526.975 2419.830 1527.055 ;
        RECT 2417.580 1526.925 2417.870 1526.975 ;
        RECT 2419.400 1526.925 2419.830 1526.975 ;
        RECT 2419.400 1526.915 2419.720 1526.925 ;
        RECT 2420.140 1525.880 2420.325 1527.055 ;
        RECT 2433.905 1527.115 2436.650 1527.155 ;
        RECT 2433.905 1526.975 2434.375 1527.115 ;
        RECT 2435.695 1527.055 2436.650 1527.115 ;
        RECT 2435.695 1526.975 2436.155 1527.055 ;
        RECT 2433.905 1526.925 2434.195 1526.975 ;
        RECT 2435.725 1526.925 2436.155 1526.975 ;
        RECT 2435.725 1526.915 2436.045 1526.925 ;
        RECT 2436.465 1525.880 2436.650 1527.055 ;
        RECT 2371.160 1525.860 2371.350 1525.880 ;
        RECT 2387.485 1525.860 2387.675 1525.880 ;
        RECT 2403.810 1525.860 2404.000 1525.880 ;
        RECT 2420.135 1525.860 2420.325 1525.880 ;
        RECT 2436.460 1525.860 2436.650 1525.880 ;
        RECT 2371.155 1525.795 2371.350 1525.860 ;
        RECT 2387.480 1525.795 2387.675 1525.860 ;
        RECT 2403.805 1525.795 2404.000 1525.860 ;
        RECT 2420.130 1525.795 2420.325 1525.860 ;
        RECT 2436.455 1525.795 2436.650 1525.860 ;
        RECT 2361.535 1524.600 2371.350 1525.795 ;
        RECT 2377.860 1524.600 2387.675 1525.795 ;
        RECT 2394.185 1524.600 2404.000 1525.795 ;
        RECT 2410.510 1524.600 2420.325 1525.795 ;
        RECT 2426.835 1524.600 2436.650 1525.795 ;
        RECT 2343.000 1523.000 2442.420 1524.600 ;
        RECT 2695.520 1496.680 2734.960 1497.160 ;
        RECT 2695.520 1491.240 2734.960 1491.720 ;
        RECT 2695.520 1485.800 2734.960 1486.280 ;
        RECT 2695.520 1480.360 2734.960 1480.840 ;
        RECT 2695.520 1474.920 2734.960 1475.400 ;
        RECT 2695.520 1469.480 2734.960 1469.960 ;
        RECT 2695.520 1464.040 2734.960 1464.520 ;
        RECT 2695.520 1458.600 2734.960 1459.080 ;
        RECT 2695.520 1453.160 2734.960 1453.640 ;
        RECT 2695.520 1447.720 2734.960 1448.200 ;
        RECT 2695.520 1442.280 2734.960 1442.760 ;
        RECT 2343.000 1435.865 2453.600 1437.465 ;
        RECT 2695.520 1436.840 2734.960 1437.320 ;
        RECT 2522.555 1436.395 2534.570 1436.550 ;
        RECT 2522.130 1436.225 2534.570 1436.395 ;
        RECT 2522.555 1436.070 2534.570 1436.225 ;
        RECT 2369.545 1433.790 2369.715 1435.865 ;
        RECT 2369.985 1433.790 2370.275 1433.820 ;
        RECT 2369.545 1433.605 2370.275 1433.790 ;
        RECT 2388.105 1433.790 2388.275 1435.865 ;
        RECT 2388.545 1433.790 2388.835 1433.820 ;
        RECT 2388.105 1433.605 2388.835 1433.790 ;
        RECT 2406.665 1433.790 2406.835 1435.865 ;
        RECT 2407.105 1433.790 2407.395 1433.820 ;
        RECT 2406.665 1433.605 2407.395 1433.790 ;
        RECT 2425.225 1433.790 2425.395 1435.865 ;
        RECT 2425.665 1433.790 2425.955 1433.820 ;
        RECT 2425.225 1433.605 2425.955 1433.790 ;
        RECT 2443.785 1433.790 2443.955 1435.865 ;
        RECT 2531.170 1434.950 2534.270 1436.070 ;
        RECT 2444.225 1433.790 2444.515 1433.820 ;
        RECT 2443.785 1433.605 2444.515 1433.790 ;
        RECT 2369.985 1433.590 2370.275 1433.605 ;
        RECT 2388.545 1433.590 2388.835 1433.605 ;
        RECT 2407.105 1433.590 2407.395 1433.605 ;
        RECT 2425.665 1433.590 2425.955 1433.605 ;
        RECT 2444.225 1433.590 2444.515 1433.605 ;
        RECT 2695.520 1431.400 2734.960 1431.880 ;
        RECT 2522.555 1429.980 2534.570 1430.135 ;
        RECT 2522.130 1429.810 2534.570 1429.980 ;
        RECT 2522.555 1429.655 2534.570 1429.810 ;
        RECT 2363.230 1429.305 2363.550 1429.565 ;
        RECT 2381.790 1429.305 2382.110 1429.565 ;
        RECT 2400.350 1429.305 2400.670 1429.565 ;
        RECT 2418.910 1429.305 2419.230 1429.565 ;
        RECT 2437.470 1429.305 2437.790 1429.565 ;
        RECT 2364.970 1428.805 2365.260 1429.035 ;
        RECT 2383.530 1428.805 2383.820 1429.035 ;
        RECT 2402.090 1428.805 2402.380 1429.035 ;
        RECT 2420.650 1428.805 2420.940 1429.035 ;
        RECT 2439.210 1428.805 2439.500 1429.035 ;
        RECT 2364.200 1428.665 2365.260 1428.805 ;
        RECT 2382.760 1428.665 2383.820 1428.805 ;
        RECT 2401.320 1428.665 2402.380 1428.805 ;
        RECT 2419.880 1428.665 2420.940 1428.805 ;
        RECT 2438.440 1428.665 2439.500 1428.805 ;
        RECT 2531.170 1428.535 2534.270 1429.655 ;
        RECT 2361.540 1427.880 2373.500 1427.905 ;
        RECT 2380.100 1427.880 2392.060 1427.905 ;
        RECT 2398.660 1427.880 2410.620 1427.905 ;
        RECT 2417.220 1427.880 2429.180 1427.905 ;
        RECT 2435.780 1427.880 2447.740 1427.905 ;
        RECT 2361.540 1426.600 2373.585 1427.880 ;
        RECT 2380.100 1426.600 2392.145 1427.880 ;
        RECT 2398.660 1426.600 2410.705 1427.880 ;
        RECT 2417.220 1426.600 2429.265 1427.880 ;
        RECT 2435.780 1426.600 2447.825 1427.880 ;
        RECT 2343.000 1425.000 2453.595 1426.600 ;
        RECT 2695.520 1425.960 2734.960 1426.440 ;
        RECT 2695.520 1420.520 2734.960 1421.000 ;
        RECT 2522.555 1415.790 2534.570 1415.945 ;
        RECT 2522.130 1415.620 2534.570 1415.790 ;
        RECT 2522.555 1415.465 2534.570 1415.620 ;
        RECT 2531.170 1414.345 2534.270 1415.465 ;
        RECT 2695.520 1415.080 2734.960 1415.560 ;
        RECT 2695.520 1409.640 2734.960 1410.120 ;
        RECT 2522.555 1408.260 2534.570 1408.415 ;
        RECT 2522.130 1408.090 2534.570 1408.260 ;
        RECT 2522.555 1407.935 2534.570 1408.090 ;
        RECT 2531.170 1406.815 2534.270 1407.935 ;
        RECT 2522.555 1402.280 2534.570 1402.435 ;
        RECT 2522.130 1402.110 2534.570 1402.280 ;
        RECT 2522.555 1401.955 2534.570 1402.110 ;
        RECT 2531.170 1400.835 2534.270 1401.955 ;
        RECT 2522.555 1393.865 2534.570 1394.020 ;
        RECT 2522.130 1393.695 2534.570 1393.865 ;
        RECT 2522.555 1393.540 2534.570 1393.695 ;
        RECT 2531.170 1392.420 2534.270 1393.540 ;
        RECT 2882.000 1360.590 2894.380 1360.745 ;
        RECT 2881.575 1360.420 2894.380 1360.590 ;
        RECT 2882.000 1360.265 2894.380 1360.420 ;
        RECT 2891.170 1359.010 2894.270 1360.265 ;
        RECT 2343.000 1335.865 2447.095 1337.465 ;
        RECT 2376.515 1333.820 2376.685 1335.865 ;
        RECT 2391.775 1333.820 2391.945 1335.865 ;
        RECT 2407.035 1333.820 2407.205 1335.865 ;
        RECT 2422.295 1333.820 2422.465 1335.865 ;
        RECT 2437.555 1333.820 2437.725 1335.865 ;
        RECT 2376.515 1333.790 2376.975 1333.820 ;
        RECT 2391.775 1333.790 2392.235 1333.820 ;
        RECT 2407.035 1333.790 2407.495 1333.820 ;
        RECT 2422.295 1333.790 2422.755 1333.820 ;
        RECT 2437.555 1333.790 2438.015 1333.820 ;
        RECT 2376.510 1333.620 2376.975 1333.790 ;
        RECT 2391.770 1333.620 2392.235 1333.790 ;
        RECT 2407.030 1333.620 2407.495 1333.790 ;
        RECT 2422.290 1333.620 2422.755 1333.790 ;
        RECT 2437.550 1333.620 2438.015 1333.790 ;
        RECT 2376.515 1333.605 2376.975 1333.620 ;
        RECT 2391.775 1333.605 2392.235 1333.620 ;
        RECT 2407.035 1333.605 2407.495 1333.620 ;
        RECT 2422.295 1333.605 2422.755 1333.620 ;
        RECT 2437.555 1333.605 2438.015 1333.620 ;
        RECT 2376.685 1333.590 2376.975 1333.605 ;
        RECT 2391.945 1333.590 2392.235 1333.605 ;
        RECT 2407.205 1333.590 2407.495 1333.605 ;
        RECT 2422.465 1333.590 2422.755 1333.605 ;
        RECT 2437.725 1333.590 2438.015 1333.605 ;
        RECT 2372.035 1329.035 2372.325 1329.265 ;
        RECT 2387.295 1329.035 2387.585 1329.265 ;
        RECT 2402.555 1329.035 2402.845 1329.265 ;
        RECT 2417.815 1329.035 2418.105 1329.265 ;
        RECT 2433.075 1329.035 2433.365 1329.265 ;
        RECT 2372.105 1328.805 2372.245 1329.035 ;
        RECT 2387.365 1328.805 2387.505 1329.035 ;
        RECT 2402.625 1328.805 2402.765 1329.035 ;
        RECT 2417.885 1328.805 2418.025 1329.035 ;
        RECT 2433.145 1328.805 2433.285 1329.035 ;
        RECT 2372.105 1328.665 2372.725 1328.805 ;
        RECT 2387.365 1328.665 2387.985 1328.805 ;
        RECT 2402.625 1328.665 2403.245 1328.805 ;
        RECT 2417.885 1328.665 2418.505 1328.805 ;
        RECT 2433.145 1328.665 2433.765 1328.805 ;
        RECT 2372.585 1328.505 2372.725 1328.665 ;
        RECT 2387.845 1328.505 2387.985 1328.665 ;
        RECT 2403.105 1328.505 2403.245 1328.665 ;
        RECT 2418.365 1328.505 2418.505 1328.665 ;
        RECT 2433.625 1328.505 2433.765 1328.665 ;
        RECT 2372.345 1328.445 2372.725 1328.505 ;
        RECT 2387.605 1328.445 2387.985 1328.505 ;
        RECT 2402.865 1328.445 2403.245 1328.505 ;
        RECT 2418.125 1328.445 2418.505 1328.505 ;
        RECT 2433.385 1328.445 2433.765 1328.505 ;
        RECT 2372.345 1328.385 2372.935 1328.445 ;
        RECT 2373.235 1328.385 2373.525 1328.425 ;
        RECT 2372.345 1328.245 2373.525 1328.385 ;
        RECT 2387.605 1328.385 2388.195 1328.445 ;
        RECT 2388.495 1328.385 2388.785 1328.425 ;
        RECT 2387.605 1328.245 2388.785 1328.385 ;
        RECT 2402.865 1328.385 2403.455 1328.445 ;
        RECT 2403.755 1328.385 2404.045 1328.425 ;
        RECT 2402.865 1328.245 2404.045 1328.385 ;
        RECT 2418.125 1328.385 2418.715 1328.445 ;
        RECT 2419.015 1328.385 2419.305 1328.425 ;
        RECT 2418.125 1328.245 2419.305 1328.385 ;
        RECT 2433.385 1328.385 2433.975 1328.445 ;
        RECT 2434.275 1328.385 2434.565 1328.425 ;
        RECT 2433.385 1328.245 2434.565 1328.385 ;
        RECT 2372.530 1328.185 2372.935 1328.245 ;
        RECT 2373.235 1328.195 2373.525 1328.245 ;
        RECT 2387.790 1328.185 2388.195 1328.245 ;
        RECT 2388.495 1328.195 2388.785 1328.245 ;
        RECT 2403.050 1328.185 2403.455 1328.245 ;
        RECT 2403.755 1328.195 2404.045 1328.245 ;
        RECT 2418.310 1328.185 2418.715 1328.245 ;
        RECT 2419.015 1328.195 2419.305 1328.245 ;
        RECT 2433.570 1328.185 2433.975 1328.245 ;
        RECT 2434.275 1328.195 2434.565 1328.245 ;
        RECT 2372.530 1327.915 2372.820 1328.185 ;
        RECT 2387.790 1327.915 2388.080 1328.185 ;
        RECT 2403.050 1327.915 2403.340 1328.185 ;
        RECT 2418.310 1327.915 2418.600 1328.185 ;
        RECT 2433.570 1327.915 2433.860 1328.185 ;
        RECT 2371.545 1326.600 2380.285 1327.915 ;
        RECT 2386.805 1326.600 2395.545 1327.915 ;
        RECT 2402.065 1326.600 2410.805 1327.915 ;
        RECT 2417.325 1326.600 2426.065 1327.915 ;
        RECT 2432.585 1326.600 2441.325 1327.915 ;
        RECT 2343.000 1325.000 2447.095 1326.600 ;
        RECT 2882.000 1161.350 2894.380 1161.505 ;
        RECT 2881.575 1161.180 2894.380 1161.350 ;
        RECT 2882.000 1161.025 2894.380 1161.180 ;
        RECT 2891.170 1159.770 2894.270 1161.025 ;
      LAYER met2 ;
        RECT 1271.310 3512.115 1274.130 3513.715 ;
        RECT 1631.310 3512.565 1634.130 3514.165 ;
        RECT 1811.310 3510.645 1814.130 3512.245 ;
        RECT 2171.310 3510.285 2174.130 3511.885 ;
        RECT 2531.310 3510.970 2534.130 3512.570 ;
        RECT 2891.310 3484.010 2894.130 3485.610 ;
        RECT 2891.310 3218.130 2894.130 3219.730 ;
        RECT 2891.310 2952.930 2894.130 2954.530 ;
        RECT 2891.310 2687.050 2894.130 2688.650 ;
        RECT 2891.310 2421.170 2894.130 2422.770 ;
        RECT 2351.310 2255.855 2354.130 2257.455 ;
        RECT 2366.920 2252.715 2367.200 2253.095 ;
        RECT 2383.505 2252.715 2383.785 2253.095 ;
        RECT 2400.090 2252.715 2400.370 2253.095 ;
        RECT 2416.675 2252.715 2416.955 2253.095 ;
        RECT 2433.255 2252.715 2433.535 2253.095 ;
        RECT 2351.310 2245.000 2354.130 2246.600 ;
        RECT 2704.410 2216.735 2705.950 2217.105 ;
        RECT 2714.070 2216.735 2715.610 2217.105 ;
        RECT 2723.730 2216.735 2725.270 2217.105 ;
        RECT 2733.390 2216.735 2734.930 2217.105 ;
        RECT 2704.410 2211.295 2705.950 2211.665 ;
        RECT 2714.070 2211.295 2715.610 2211.665 ;
        RECT 2723.730 2211.295 2725.270 2211.665 ;
        RECT 2733.390 2211.295 2734.930 2211.665 ;
        RECT 2704.410 2205.855 2705.950 2206.225 ;
        RECT 2714.070 2205.855 2715.610 2206.225 ;
        RECT 2723.730 2205.855 2725.270 2206.225 ;
        RECT 2733.390 2205.855 2734.930 2206.225 ;
        RECT 2704.410 2200.415 2705.950 2200.785 ;
        RECT 2714.070 2200.415 2715.610 2200.785 ;
        RECT 2723.730 2200.415 2725.270 2200.785 ;
        RECT 2733.390 2200.415 2734.930 2200.785 ;
        RECT 2704.410 2194.975 2705.950 2195.345 ;
        RECT 2714.070 2194.975 2715.610 2195.345 ;
        RECT 2723.730 2194.975 2725.270 2195.345 ;
        RECT 2733.390 2194.975 2734.930 2195.345 ;
        RECT 2704.410 2189.535 2705.950 2189.905 ;
        RECT 2714.070 2189.535 2715.610 2189.905 ;
        RECT 2723.730 2189.535 2725.270 2189.905 ;
        RECT 2733.390 2189.535 2734.930 2189.905 ;
        RECT 2704.410 2184.095 2705.950 2184.465 ;
        RECT 2714.070 2184.095 2715.610 2184.465 ;
        RECT 2723.730 2184.095 2725.270 2184.465 ;
        RECT 2733.390 2184.095 2734.930 2184.465 ;
        RECT 2704.410 2178.655 2705.950 2179.025 ;
        RECT 2714.070 2178.655 2715.610 2179.025 ;
        RECT 2723.730 2178.655 2725.270 2179.025 ;
        RECT 2733.390 2178.655 2734.930 2179.025 ;
        RECT 2704.410 2173.215 2705.950 2173.585 ;
        RECT 2714.070 2173.215 2715.610 2173.585 ;
        RECT 2723.730 2173.215 2725.270 2173.585 ;
        RECT 2733.390 2173.215 2734.930 2173.585 ;
        RECT 2704.410 2167.775 2705.950 2168.145 ;
        RECT 2714.070 2167.775 2715.610 2168.145 ;
        RECT 2723.730 2167.775 2725.270 2168.145 ;
        RECT 2733.390 2167.775 2734.930 2168.145 ;
        RECT 2351.310 2163.860 2354.130 2165.460 ;
        RECT 2704.410 2162.335 2705.950 2162.705 ;
        RECT 2714.070 2162.335 2715.610 2162.705 ;
        RECT 2723.730 2162.335 2725.270 2162.705 ;
        RECT 2733.390 2162.335 2734.930 2162.705 ;
        RECT 2367.020 2160.065 2367.300 2160.435 ;
        RECT 2384.240 2160.065 2384.520 2160.435 ;
        RECT 2401.460 2160.065 2401.740 2160.435 ;
        RECT 2418.680 2160.065 2418.960 2160.435 ;
        RECT 2435.900 2160.065 2436.180 2160.435 ;
        RECT 2704.410 2156.895 2705.950 2157.265 ;
        RECT 2714.070 2156.895 2715.610 2157.265 ;
        RECT 2723.730 2156.895 2725.270 2157.265 ;
        RECT 2733.390 2156.895 2734.930 2157.265 ;
        RECT 2891.310 2155.970 2894.130 2157.570 ;
        RECT 2351.310 2153.000 2354.130 2154.600 ;
        RECT 2704.410 2151.455 2705.950 2151.825 ;
        RECT 2714.070 2151.455 2715.610 2151.825 ;
        RECT 2723.730 2151.455 2725.270 2151.825 ;
        RECT 2733.390 2151.455 2734.930 2151.825 ;
        RECT 2704.410 2146.015 2705.950 2146.385 ;
        RECT 2714.070 2146.015 2715.610 2146.385 ;
        RECT 2723.730 2146.015 2725.270 2146.385 ;
        RECT 2733.390 2146.015 2734.930 2146.385 ;
        RECT 2704.410 2140.575 2705.950 2140.945 ;
        RECT 2714.070 2140.575 2715.610 2140.945 ;
        RECT 2723.730 2140.575 2725.270 2140.945 ;
        RECT 2733.390 2140.575 2734.930 2140.945 ;
        RECT 2704.410 2135.135 2705.950 2135.505 ;
        RECT 2714.070 2135.135 2715.610 2135.505 ;
        RECT 2723.730 2135.135 2725.270 2135.505 ;
        RECT 2733.390 2135.135 2734.930 2135.505 ;
        RECT 2531.310 2132.595 2534.130 2134.195 ;
        RECT 2704.410 2129.695 2705.950 2130.065 ;
        RECT 2714.070 2129.695 2715.610 2130.065 ;
        RECT 2723.730 2129.695 2725.270 2130.065 ;
        RECT 2733.390 2129.695 2734.930 2130.065 ;
        RECT 2531.310 2125.065 2534.130 2126.665 ;
        RECT 2531.310 2119.085 2534.130 2120.685 ;
        RECT 2531.310 2113.140 2534.130 2114.740 ;
        RECT 2531.310 2107.495 2534.130 2109.095 ;
        RECT 2531.310 2101.490 2534.130 2103.090 ;
        RECT 2351.310 2058.860 2354.130 2060.460 ;
        RECT 2370.450 2052.245 2370.730 2052.620 ;
        RECT 2386.775 2052.245 2387.055 2052.620 ;
        RECT 2403.100 2052.245 2403.380 2052.620 ;
        RECT 2419.425 2052.245 2419.705 2052.620 ;
        RECT 2435.750 2052.245 2436.030 2052.620 ;
        RECT 2370.460 2051.995 2370.720 2052.245 ;
        RECT 2386.785 2051.995 2387.045 2052.245 ;
        RECT 2403.110 2051.995 2403.370 2052.245 ;
        RECT 2419.435 2051.995 2419.695 2052.245 ;
        RECT 2435.760 2051.995 2436.020 2052.245 ;
        RECT 2351.310 2048.000 2354.130 2049.600 ;
        RECT 2704.410 2036.735 2705.950 2037.105 ;
        RECT 2714.070 2036.735 2715.610 2037.105 ;
        RECT 2723.730 2036.735 2725.270 2037.105 ;
        RECT 2733.390 2036.735 2734.930 2037.105 ;
        RECT 2704.410 2031.295 2705.950 2031.665 ;
        RECT 2714.070 2031.295 2715.610 2031.665 ;
        RECT 2723.730 2031.295 2725.270 2031.665 ;
        RECT 2733.390 2031.295 2734.930 2031.665 ;
        RECT 2704.410 2025.855 2705.950 2026.225 ;
        RECT 2714.070 2025.855 2715.610 2026.225 ;
        RECT 2723.730 2025.855 2725.270 2026.225 ;
        RECT 2733.390 2025.855 2734.930 2026.225 ;
        RECT 2704.410 2020.415 2705.950 2020.785 ;
        RECT 2714.070 2020.415 2715.610 2020.785 ;
        RECT 2723.730 2020.415 2725.270 2020.785 ;
        RECT 2733.390 2020.415 2734.930 2020.785 ;
        RECT 2704.410 2014.975 2705.950 2015.345 ;
        RECT 2714.070 2014.975 2715.610 2015.345 ;
        RECT 2723.730 2014.975 2725.270 2015.345 ;
        RECT 2733.390 2014.975 2734.930 2015.345 ;
        RECT 2704.410 2009.535 2705.950 2009.905 ;
        RECT 2714.070 2009.535 2715.610 2009.905 ;
        RECT 2723.730 2009.535 2725.270 2009.905 ;
        RECT 2733.390 2009.535 2734.930 2009.905 ;
        RECT 2704.410 2004.095 2705.950 2004.465 ;
        RECT 2714.070 2004.095 2715.610 2004.465 ;
        RECT 2723.730 2004.095 2725.270 2004.465 ;
        RECT 2733.390 2004.095 2734.930 2004.465 ;
        RECT 2704.410 1998.655 2705.950 1999.025 ;
        RECT 2714.070 1998.655 2715.610 1999.025 ;
        RECT 2723.730 1998.655 2725.270 1999.025 ;
        RECT 2733.390 1998.655 2734.930 1999.025 ;
        RECT 2704.410 1993.215 2705.950 1993.585 ;
        RECT 2714.070 1993.215 2715.610 1993.585 ;
        RECT 2723.730 1993.215 2725.270 1993.585 ;
        RECT 2733.390 1993.215 2734.930 1993.585 ;
        RECT 2704.410 1987.775 2705.950 1988.145 ;
        RECT 2714.070 1987.775 2715.610 1988.145 ;
        RECT 2723.730 1987.775 2725.270 1988.145 ;
        RECT 2733.390 1987.775 2734.930 1988.145 ;
        RECT 2704.410 1982.335 2705.950 1982.705 ;
        RECT 2714.070 1982.335 2715.610 1982.705 ;
        RECT 2723.730 1982.335 2725.270 1982.705 ;
        RECT 2733.390 1982.335 2734.930 1982.705 ;
        RECT 2531.310 1980.340 2534.130 1981.940 ;
        RECT 2704.410 1976.895 2705.950 1977.265 ;
        RECT 2714.070 1976.895 2715.610 1977.265 ;
        RECT 2723.730 1976.895 2725.270 1977.265 ;
        RECT 2733.390 1976.895 2734.930 1977.265 ;
        RECT 2531.310 1972.810 2534.130 1974.410 ;
        RECT 2704.410 1971.455 2705.950 1971.825 ;
        RECT 2714.070 1971.455 2715.610 1971.825 ;
        RECT 2723.730 1971.455 2725.270 1971.825 ;
        RECT 2733.390 1971.455 2734.930 1971.825 ;
        RECT 2531.310 1966.830 2534.130 1968.430 ;
        RECT 2704.410 1966.015 2705.950 1966.385 ;
        RECT 2714.070 1966.015 2715.610 1966.385 ;
        RECT 2723.730 1966.015 2725.270 1966.385 ;
        RECT 2733.390 1966.015 2734.930 1966.385 ;
        RECT 2531.310 1960.885 2534.130 1962.485 ;
        RECT 2704.410 1960.575 2705.950 1960.945 ;
        RECT 2714.070 1960.575 2715.610 1960.945 ;
        RECT 2723.730 1960.575 2725.270 1960.945 ;
        RECT 2733.390 1960.575 2734.930 1960.945 ;
        RECT 2351.310 1953.865 2354.130 1955.465 ;
        RECT 2531.310 1955.240 2534.130 1956.840 ;
        RECT 2704.410 1955.135 2705.950 1955.505 ;
        RECT 2714.070 1955.135 2715.610 1955.505 ;
        RECT 2723.730 1955.135 2725.270 1955.505 ;
        RECT 2733.390 1955.135 2734.930 1955.505 ;
        RECT 2531.310 1949.235 2534.130 1950.835 ;
        RECT 2704.410 1949.695 2705.950 1950.065 ;
        RECT 2714.070 1949.695 2715.610 1950.065 ;
        RECT 2723.730 1949.695 2725.270 1950.065 ;
        RECT 2733.390 1949.695 2734.930 1950.065 ;
        RECT 2363.265 1947.505 2363.525 1947.595 ;
        RECT 2381.825 1947.505 2382.085 1947.595 ;
        RECT 2400.385 1947.505 2400.645 1947.595 ;
        RECT 2418.945 1947.505 2419.205 1947.595 ;
        RECT 2437.505 1947.505 2437.765 1947.595 ;
        RECT 2363.205 1947.275 2363.525 1947.505 ;
        RECT 2381.765 1947.275 2382.085 1947.505 ;
        RECT 2400.325 1947.275 2400.645 1947.505 ;
        RECT 2418.885 1947.275 2419.205 1947.505 ;
        RECT 2437.445 1947.275 2437.765 1947.505 ;
        RECT 2363.205 1946.945 2363.345 1947.275 ;
        RECT 2363.515 1946.945 2363.795 1947.060 ;
        RECT 2364.985 1946.945 2365.245 1947.035 ;
        RECT 2363.205 1946.805 2365.245 1946.945 ;
        RECT 2381.765 1946.945 2381.905 1947.275 ;
        RECT 2382.075 1946.945 2382.355 1947.060 ;
        RECT 2383.545 1946.945 2383.805 1947.035 ;
        RECT 2381.765 1946.805 2383.805 1946.945 ;
        RECT 2400.325 1946.945 2400.465 1947.275 ;
        RECT 2400.635 1946.945 2400.915 1947.060 ;
        RECT 2402.105 1946.945 2402.365 1947.035 ;
        RECT 2400.325 1946.805 2402.365 1946.945 ;
        RECT 2418.885 1946.945 2419.025 1947.275 ;
        RECT 2419.195 1946.945 2419.475 1947.060 ;
        RECT 2420.665 1946.945 2420.925 1947.035 ;
        RECT 2418.885 1946.805 2420.925 1946.945 ;
        RECT 2437.445 1946.945 2437.585 1947.275 ;
        RECT 2437.755 1946.945 2438.035 1947.060 ;
        RECT 2439.225 1946.945 2439.485 1947.035 ;
        RECT 2437.445 1946.805 2439.485 1946.945 ;
        RECT 2363.515 1946.685 2363.795 1946.805 ;
        RECT 2364.985 1946.715 2365.245 1946.805 ;
        RECT 2382.075 1946.685 2382.355 1946.805 ;
        RECT 2383.545 1946.715 2383.805 1946.805 ;
        RECT 2400.635 1946.685 2400.915 1946.805 ;
        RECT 2402.105 1946.715 2402.365 1946.805 ;
        RECT 2419.195 1946.685 2419.475 1946.805 ;
        RECT 2420.665 1946.715 2420.925 1946.805 ;
        RECT 2437.755 1946.685 2438.035 1946.805 ;
        RECT 2439.225 1946.715 2439.485 1946.805 ;
        RECT 2363.615 1945.635 2363.785 1946.685 ;
        RECT 2382.175 1945.635 2382.345 1946.685 ;
        RECT 2400.735 1945.635 2400.905 1946.685 ;
        RECT 2419.295 1945.635 2419.465 1946.685 ;
        RECT 2437.855 1945.635 2438.025 1946.685 ;
        RECT 2363.590 1945.295 2363.930 1945.635 ;
        RECT 2382.150 1945.295 2382.490 1945.635 ;
        RECT 2400.710 1945.295 2401.050 1945.635 ;
        RECT 2419.270 1945.295 2419.610 1945.635 ;
        RECT 2437.830 1945.295 2438.170 1945.635 ;
        RECT 2351.310 1943.000 2354.130 1944.600 ;
        RECT 2891.310 1890.090 2894.130 1891.690 ;
        RECT 2704.410 1856.735 2705.950 1857.105 ;
        RECT 2714.070 1856.735 2715.610 1857.105 ;
        RECT 2723.730 1856.735 2725.270 1857.105 ;
        RECT 2733.390 1856.735 2734.930 1857.105 ;
        RECT 2704.410 1851.295 2705.950 1851.665 ;
        RECT 2714.070 1851.295 2715.610 1851.665 ;
        RECT 2723.730 1851.295 2725.270 1851.665 ;
        RECT 2733.390 1851.295 2734.930 1851.665 ;
        RECT 2704.410 1845.855 2705.950 1846.225 ;
        RECT 2714.070 1845.855 2715.610 1846.225 ;
        RECT 2723.730 1845.855 2725.270 1846.225 ;
        RECT 2733.390 1845.855 2734.930 1846.225 ;
        RECT 2704.410 1840.415 2705.950 1840.785 ;
        RECT 2714.070 1840.415 2715.610 1840.785 ;
        RECT 2723.730 1840.415 2725.270 1840.785 ;
        RECT 2733.390 1840.415 2734.930 1840.785 ;
        RECT 2704.410 1834.975 2705.950 1835.345 ;
        RECT 2714.070 1834.975 2715.610 1835.345 ;
        RECT 2723.730 1834.975 2725.270 1835.345 ;
        RECT 2733.390 1834.975 2734.930 1835.345 ;
        RECT 2704.410 1829.535 2705.950 1829.905 ;
        RECT 2714.070 1829.535 2715.610 1829.905 ;
        RECT 2723.730 1829.535 2725.270 1829.905 ;
        RECT 2733.390 1829.535 2734.930 1829.905 ;
        RECT 2704.410 1824.095 2705.950 1824.465 ;
        RECT 2714.070 1824.095 2715.610 1824.465 ;
        RECT 2723.730 1824.095 2725.270 1824.465 ;
        RECT 2733.390 1824.095 2734.930 1824.465 ;
        RECT 2704.410 1818.655 2705.950 1819.025 ;
        RECT 2714.070 1818.655 2715.610 1819.025 ;
        RECT 2723.730 1818.655 2725.270 1819.025 ;
        RECT 2733.390 1818.655 2734.930 1819.025 ;
        RECT 2704.410 1813.215 2705.950 1813.585 ;
        RECT 2714.070 1813.215 2715.610 1813.585 ;
        RECT 2723.730 1813.215 2725.270 1813.585 ;
        RECT 2733.390 1813.215 2734.930 1813.585 ;
        RECT 2704.410 1807.775 2705.950 1808.145 ;
        RECT 2714.070 1807.775 2715.610 1808.145 ;
        RECT 2723.730 1807.775 2725.270 1808.145 ;
        RECT 2733.390 1807.775 2734.930 1808.145 ;
        RECT 2531.310 1803.370 2534.130 1804.970 ;
        RECT 2704.410 1802.335 2705.950 1802.705 ;
        RECT 2714.070 1802.335 2715.610 1802.705 ;
        RECT 2723.730 1802.335 2725.270 1802.705 ;
        RECT 2733.390 1802.335 2734.930 1802.705 ;
        RECT 2531.310 1795.840 2534.130 1797.440 ;
        RECT 2704.410 1796.895 2705.950 1797.265 ;
        RECT 2714.070 1796.895 2715.610 1797.265 ;
        RECT 2723.730 1796.895 2725.270 1797.265 ;
        RECT 2733.390 1796.895 2734.930 1797.265 ;
        RECT 2351.310 1790.865 2354.130 1792.465 ;
        RECT 2531.310 1789.860 2534.130 1791.460 ;
        RECT 2704.410 1791.455 2705.950 1791.825 ;
        RECT 2714.070 1791.455 2715.610 1791.825 ;
        RECT 2723.730 1791.455 2725.270 1791.825 ;
        RECT 2733.390 1791.455 2734.930 1791.825 ;
        RECT 2704.410 1786.015 2705.950 1786.385 ;
        RECT 2714.070 1786.015 2715.610 1786.385 ;
        RECT 2723.730 1786.015 2725.270 1786.385 ;
        RECT 2733.390 1786.015 2734.930 1786.385 ;
        RECT 2531.310 1783.915 2534.130 1785.515 ;
        RECT 2372.465 1783.475 2372.745 1783.500 ;
        RECT 2387.725 1783.475 2388.005 1783.500 ;
        RECT 2402.985 1783.475 2403.265 1783.500 ;
        RECT 2418.245 1783.475 2418.525 1783.500 ;
        RECT 2433.505 1783.475 2433.785 1783.500 ;
        RECT 2372.465 1783.155 2372.855 1783.475 ;
        RECT 2387.725 1783.155 2388.115 1783.475 ;
        RECT 2402.985 1783.155 2403.375 1783.475 ;
        RECT 2418.245 1783.155 2418.635 1783.475 ;
        RECT 2433.505 1783.155 2433.895 1783.475 ;
        RECT 2372.465 1783.125 2372.745 1783.155 ;
        RECT 2387.725 1783.125 2388.005 1783.155 ;
        RECT 2402.985 1783.125 2403.265 1783.155 ;
        RECT 2418.245 1783.125 2418.525 1783.155 ;
        RECT 2433.505 1783.125 2433.785 1783.155 ;
        RECT 2351.310 1780.000 2354.130 1781.600 ;
        RECT 2704.410 1780.575 2705.950 1780.945 ;
        RECT 2714.070 1780.575 2715.610 1780.945 ;
        RECT 2723.730 1780.575 2725.270 1780.945 ;
        RECT 2733.390 1780.575 2734.930 1780.945 ;
        RECT 2531.310 1778.270 2534.130 1779.870 ;
        RECT 2704.410 1775.135 2705.950 1775.505 ;
        RECT 2714.070 1775.135 2715.610 1775.505 ;
        RECT 2723.730 1775.135 2725.270 1775.505 ;
        RECT 2733.390 1775.135 2734.930 1775.505 ;
        RECT 2704.410 1769.695 2705.950 1770.065 ;
        RECT 2714.070 1769.695 2715.610 1770.065 ;
        RECT 2723.730 1769.695 2725.270 1770.065 ;
        RECT 2733.390 1769.695 2734.930 1770.065 ;
        RECT 2531.310 1766.800 2534.130 1768.400 ;
        RECT 2351.310 1710.860 2354.130 1712.460 ;
        RECT 2367.280 1707.715 2367.560 1708.095 ;
        RECT 2383.865 1707.715 2384.145 1708.095 ;
        RECT 2400.450 1707.720 2400.730 1708.100 ;
        RECT 2417.035 1707.725 2417.315 1708.105 ;
        RECT 2433.615 1707.725 2433.895 1708.105 ;
        RECT 2351.310 1700.000 2354.130 1701.600 ;
        RECT 2704.410 1676.735 2705.950 1677.105 ;
        RECT 2714.070 1676.735 2715.610 1677.105 ;
        RECT 2723.730 1676.735 2725.270 1677.105 ;
        RECT 2733.390 1676.735 2734.930 1677.105 ;
        RECT 2704.410 1671.295 2705.950 1671.665 ;
        RECT 2714.070 1671.295 2715.610 1671.665 ;
        RECT 2723.730 1671.295 2725.270 1671.665 ;
        RECT 2733.390 1671.295 2734.930 1671.665 ;
        RECT 2704.410 1665.855 2705.950 1666.225 ;
        RECT 2714.070 1665.855 2715.610 1666.225 ;
        RECT 2723.730 1665.855 2725.270 1666.225 ;
        RECT 2733.390 1665.855 2734.930 1666.225 ;
        RECT 2704.410 1660.415 2705.950 1660.785 ;
        RECT 2714.070 1660.415 2715.610 1660.785 ;
        RECT 2723.730 1660.415 2725.270 1660.785 ;
        RECT 2733.390 1660.415 2734.930 1660.785 ;
        RECT 2704.410 1654.975 2705.950 1655.345 ;
        RECT 2714.070 1654.975 2715.610 1655.345 ;
        RECT 2723.730 1654.975 2725.270 1655.345 ;
        RECT 2733.390 1654.975 2734.930 1655.345 ;
        RECT 2704.410 1649.535 2705.950 1649.905 ;
        RECT 2714.070 1649.535 2715.610 1649.905 ;
        RECT 2723.730 1649.535 2725.270 1649.905 ;
        RECT 2733.390 1649.535 2734.930 1649.905 ;
        RECT 2704.410 1644.095 2705.950 1644.465 ;
        RECT 2714.070 1644.095 2715.610 1644.465 ;
        RECT 2723.730 1644.095 2725.270 1644.465 ;
        RECT 2733.390 1644.095 2734.930 1644.465 ;
        RECT 2704.410 1638.655 2705.950 1639.025 ;
        RECT 2714.070 1638.655 2715.610 1639.025 ;
        RECT 2723.730 1638.655 2725.270 1639.025 ;
        RECT 2733.390 1638.655 2734.930 1639.025 ;
        RECT 2704.410 1633.215 2705.950 1633.585 ;
        RECT 2714.070 1633.215 2715.610 1633.585 ;
        RECT 2723.730 1633.215 2725.270 1633.585 ;
        RECT 2733.390 1633.215 2734.930 1633.585 ;
        RECT 2704.410 1627.775 2705.950 1628.145 ;
        RECT 2714.070 1627.775 2715.610 1628.145 ;
        RECT 2723.730 1627.775 2725.270 1628.145 ;
        RECT 2733.390 1627.775 2734.930 1628.145 ;
        RECT 2891.310 1624.210 2894.130 1625.810 ;
        RECT 2531.310 1622.235 2534.130 1623.835 ;
        RECT 2704.410 1622.335 2705.950 1622.705 ;
        RECT 2714.070 1622.335 2715.610 1622.705 ;
        RECT 2723.730 1622.335 2725.270 1622.705 ;
        RECT 2733.390 1622.335 2734.930 1622.705 ;
        RECT 2531.310 1615.820 2534.130 1617.420 ;
        RECT 2704.410 1616.895 2705.950 1617.265 ;
        RECT 2714.070 1616.895 2715.610 1617.265 ;
        RECT 2723.730 1616.895 2725.270 1617.265 ;
        RECT 2733.390 1616.895 2734.930 1617.265 ;
        RECT 2351.310 1610.860 2354.130 1612.460 ;
        RECT 2704.410 1611.455 2705.950 1611.825 ;
        RECT 2714.070 1611.455 2715.610 1611.825 ;
        RECT 2723.730 1611.455 2725.270 1611.825 ;
        RECT 2733.390 1611.455 2734.930 1611.825 ;
        RECT 2366.995 1607.065 2367.275 1607.435 ;
        RECT 2384.215 1607.065 2384.495 1607.435 ;
        RECT 2401.435 1607.070 2401.715 1607.440 ;
        RECT 2418.655 1607.065 2418.935 1607.435 ;
        RECT 2435.875 1607.065 2436.155 1607.435 ;
        RECT 2704.410 1606.015 2705.950 1606.385 ;
        RECT 2714.070 1606.015 2715.610 1606.385 ;
        RECT 2723.730 1606.015 2725.270 1606.385 ;
        RECT 2733.390 1606.015 2734.930 1606.385 ;
        RECT 2351.310 1600.000 2354.130 1601.600 ;
        RECT 2704.410 1600.575 2705.950 1600.945 ;
        RECT 2714.070 1600.575 2715.610 1600.945 ;
        RECT 2723.730 1600.575 2725.270 1600.945 ;
        RECT 2733.390 1600.575 2734.930 1600.945 ;
        RECT 2704.410 1595.135 2705.950 1595.505 ;
        RECT 2714.070 1595.135 2715.610 1595.505 ;
        RECT 2723.730 1595.135 2725.270 1595.505 ;
        RECT 2733.390 1595.135 2734.930 1595.505 ;
        RECT 2704.410 1589.695 2705.950 1590.065 ;
        RECT 2714.070 1589.695 2715.610 1590.065 ;
        RECT 2723.730 1589.695 2725.270 1590.065 ;
        RECT 2733.390 1589.695 2734.930 1590.065 ;
        RECT 2531.310 1586.575 2534.130 1588.175 ;
        RECT 2531.310 1579.045 2534.130 1580.645 ;
        RECT 2531.310 1573.065 2534.130 1574.665 ;
        RECT 2531.310 1564.650 2534.130 1566.250 ;
        RECT 2351.310 1533.860 2354.130 1535.460 ;
        RECT 2370.445 1527.135 2370.725 1527.510 ;
        RECT 2386.770 1527.135 2387.050 1527.510 ;
        RECT 2403.095 1527.135 2403.375 1527.510 ;
        RECT 2419.420 1527.135 2419.700 1527.510 ;
        RECT 2435.745 1527.135 2436.025 1527.510 ;
        RECT 2370.455 1526.885 2370.715 1527.135 ;
        RECT 2386.780 1526.885 2387.040 1527.135 ;
        RECT 2403.105 1526.885 2403.365 1527.135 ;
        RECT 2419.430 1526.885 2419.690 1527.135 ;
        RECT 2435.755 1526.885 2436.015 1527.135 ;
        RECT 2351.310 1523.000 2354.130 1524.600 ;
        RECT 2704.410 1496.735 2705.950 1497.105 ;
        RECT 2714.070 1496.735 2715.610 1497.105 ;
        RECT 2723.730 1496.735 2725.270 1497.105 ;
        RECT 2733.390 1496.735 2734.930 1497.105 ;
        RECT 2704.410 1491.295 2705.950 1491.665 ;
        RECT 2714.070 1491.295 2715.610 1491.665 ;
        RECT 2723.730 1491.295 2725.270 1491.665 ;
        RECT 2733.390 1491.295 2734.930 1491.665 ;
        RECT 2704.410 1485.855 2705.950 1486.225 ;
        RECT 2714.070 1485.855 2715.610 1486.225 ;
        RECT 2723.730 1485.855 2725.270 1486.225 ;
        RECT 2733.390 1485.855 2734.930 1486.225 ;
        RECT 2704.410 1480.415 2705.950 1480.785 ;
        RECT 2714.070 1480.415 2715.610 1480.785 ;
        RECT 2723.730 1480.415 2725.270 1480.785 ;
        RECT 2733.390 1480.415 2734.930 1480.785 ;
        RECT 2704.410 1474.975 2705.950 1475.345 ;
        RECT 2714.070 1474.975 2715.610 1475.345 ;
        RECT 2723.730 1474.975 2725.270 1475.345 ;
        RECT 2733.390 1474.975 2734.930 1475.345 ;
        RECT 2704.410 1469.535 2705.950 1469.905 ;
        RECT 2714.070 1469.535 2715.610 1469.905 ;
        RECT 2723.730 1469.535 2725.270 1469.905 ;
        RECT 2733.390 1469.535 2734.930 1469.905 ;
        RECT 2704.410 1464.095 2705.950 1464.465 ;
        RECT 2714.070 1464.095 2715.610 1464.465 ;
        RECT 2723.730 1464.095 2725.270 1464.465 ;
        RECT 2733.390 1464.095 2734.930 1464.465 ;
        RECT 2704.410 1458.655 2705.950 1459.025 ;
        RECT 2714.070 1458.655 2715.610 1459.025 ;
        RECT 2723.730 1458.655 2725.270 1459.025 ;
        RECT 2733.390 1458.655 2734.930 1459.025 ;
        RECT 2704.410 1453.215 2705.950 1453.585 ;
        RECT 2714.070 1453.215 2715.610 1453.585 ;
        RECT 2723.730 1453.215 2725.270 1453.585 ;
        RECT 2733.390 1453.215 2734.930 1453.585 ;
        RECT 2704.410 1447.775 2705.950 1448.145 ;
        RECT 2714.070 1447.775 2715.610 1448.145 ;
        RECT 2723.730 1447.775 2725.270 1448.145 ;
        RECT 2733.390 1447.775 2734.930 1448.145 ;
        RECT 2704.410 1442.335 2705.950 1442.705 ;
        RECT 2714.070 1442.335 2715.610 1442.705 ;
        RECT 2723.730 1442.335 2725.270 1442.705 ;
        RECT 2733.390 1442.335 2734.930 1442.705 ;
        RECT 2351.310 1435.865 2354.130 1437.465 ;
        RECT 2704.410 1436.895 2705.950 1437.265 ;
        RECT 2714.070 1436.895 2715.610 1437.265 ;
        RECT 2723.730 1436.895 2725.270 1437.265 ;
        RECT 2733.390 1436.895 2734.930 1437.265 ;
        RECT 2531.310 1434.950 2534.130 1436.550 ;
        RECT 2704.410 1431.455 2705.950 1431.825 ;
        RECT 2714.070 1431.455 2715.610 1431.825 ;
        RECT 2723.730 1431.455 2725.270 1431.825 ;
        RECT 2733.390 1431.455 2734.930 1431.825 ;
        RECT 2363.260 1429.505 2363.520 1429.595 ;
        RECT 2381.820 1429.505 2382.080 1429.595 ;
        RECT 2400.380 1429.505 2400.640 1429.595 ;
        RECT 2418.940 1429.505 2419.200 1429.595 ;
        RECT 2437.500 1429.505 2437.760 1429.595 ;
        RECT 2363.200 1429.275 2363.520 1429.505 ;
        RECT 2381.760 1429.275 2382.080 1429.505 ;
        RECT 2400.320 1429.275 2400.640 1429.505 ;
        RECT 2418.880 1429.275 2419.200 1429.505 ;
        RECT 2437.440 1429.275 2437.760 1429.505 ;
        RECT 2363.200 1428.945 2363.340 1429.275 ;
        RECT 2363.510 1428.945 2363.790 1429.060 ;
        RECT 2364.980 1428.945 2365.240 1429.035 ;
        RECT 2363.200 1428.805 2365.240 1428.945 ;
        RECT 2381.760 1428.945 2381.900 1429.275 ;
        RECT 2382.070 1428.945 2382.350 1429.060 ;
        RECT 2383.540 1428.945 2383.800 1429.035 ;
        RECT 2381.760 1428.805 2383.800 1428.945 ;
        RECT 2400.320 1428.945 2400.460 1429.275 ;
        RECT 2400.630 1428.945 2400.910 1429.060 ;
        RECT 2402.100 1428.945 2402.360 1429.035 ;
        RECT 2400.320 1428.805 2402.360 1428.945 ;
        RECT 2418.880 1428.945 2419.020 1429.275 ;
        RECT 2419.190 1428.945 2419.470 1429.060 ;
        RECT 2420.660 1428.945 2420.920 1429.035 ;
        RECT 2418.880 1428.805 2420.920 1428.945 ;
        RECT 2437.440 1428.945 2437.580 1429.275 ;
        RECT 2437.750 1428.945 2438.030 1429.060 ;
        RECT 2439.220 1428.945 2439.480 1429.035 ;
        RECT 2437.440 1428.805 2439.480 1428.945 ;
        RECT 2363.510 1428.685 2363.790 1428.805 ;
        RECT 2364.980 1428.715 2365.240 1428.805 ;
        RECT 2382.070 1428.685 2382.350 1428.805 ;
        RECT 2383.540 1428.715 2383.800 1428.805 ;
        RECT 2400.630 1428.685 2400.910 1428.805 ;
        RECT 2402.100 1428.715 2402.360 1428.805 ;
        RECT 2419.190 1428.685 2419.470 1428.805 ;
        RECT 2420.660 1428.715 2420.920 1428.805 ;
        RECT 2437.750 1428.685 2438.030 1428.805 ;
        RECT 2439.220 1428.715 2439.480 1428.805 ;
        RECT 2363.610 1427.635 2363.780 1428.685 ;
        RECT 2382.170 1427.635 2382.340 1428.685 ;
        RECT 2400.730 1427.635 2400.900 1428.685 ;
        RECT 2419.290 1427.635 2419.460 1428.685 ;
        RECT 2437.850 1427.635 2438.020 1428.685 ;
        RECT 2531.310 1428.535 2534.130 1430.135 ;
        RECT 2363.585 1427.295 2363.925 1427.635 ;
        RECT 2382.145 1427.295 2382.485 1427.635 ;
        RECT 2400.705 1427.295 2401.045 1427.635 ;
        RECT 2419.265 1427.295 2419.605 1427.635 ;
        RECT 2437.825 1427.295 2438.165 1427.635 ;
        RECT 2351.310 1425.000 2354.130 1426.600 ;
        RECT 2704.410 1426.015 2705.950 1426.385 ;
        RECT 2714.070 1426.015 2715.610 1426.385 ;
        RECT 2723.730 1426.015 2725.270 1426.385 ;
        RECT 2733.390 1426.015 2734.930 1426.385 ;
        RECT 2704.410 1420.575 2705.950 1420.945 ;
        RECT 2714.070 1420.575 2715.610 1420.945 ;
        RECT 2723.730 1420.575 2725.270 1420.945 ;
        RECT 2733.390 1420.575 2734.930 1420.945 ;
        RECT 2531.310 1414.345 2534.130 1415.945 ;
        RECT 2704.410 1415.135 2705.950 1415.505 ;
        RECT 2714.070 1415.135 2715.610 1415.505 ;
        RECT 2723.730 1415.135 2725.270 1415.505 ;
        RECT 2733.390 1415.135 2734.930 1415.505 ;
        RECT 2704.410 1409.695 2705.950 1410.065 ;
        RECT 2714.070 1409.695 2715.610 1410.065 ;
        RECT 2723.730 1409.695 2725.270 1410.065 ;
        RECT 2733.390 1409.695 2734.930 1410.065 ;
        RECT 2531.310 1406.815 2534.130 1408.415 ;
        RECT 2531.310 1400.835 2534.130 1402.435 ;
        RECT 2531.310 1392.420 2534.130 1394.020 ;
        RECT 2891.310 1359.010 2894.130 1360.610 ;
        RECT 2351.310 1335.865 2354.130 1337.465 ;
        RECT 2372.515 1328.475 2372.795 1328.500 ;
        RECT 2387.775 1328.475 2388.055 1328.500 ;
        RECT 2403.035 1328.475 2403.315 1328.500 ;
        RECT 2418.295 1328.475 2418.575 1328.500 ;
        RECT 2433.555 1328.475 2433.835 1328.500 ;
        RECT 2372.515 1328.155 2372.905 1328.475 ;
        RECT 2387.775 1328.155 2388.165 1328.475 ;
        RECT 2403.035 1328.155 2403.425 1328.475 ;
        RECT 2418.295 1328.155 2418.685 1328.475 ;
        RECT 2433.555 1328.155 2433.945 1328.475 ;
        RECT 2372.515 1328.125 2372.795 1328.155 ;
        RECT 2387.775 1328.125 2388.055 1328.155 ;
        RECT 2403.035 1328.125 2403.315 1328.155 ;
        RECT 2418.295 1328.125 2418.575 1328.155 ;
        RECT 2433.555 1328.125 2433.835 1328.155 ;
        RECT 2351.310 1325.000 2354.130 1326.600 ;
        RECT 2891.310 1159.770 2894.130 1161.370 ;
      LAYER met3 ;
        RECT 1271.330 3512.150 1274.110 3513.680 ;
        RECT 1631.330 3512.600 1634.110 3514.130 ;
        RECT 1811.330 3510.680 1814.110 3512.210 ;
        RECT 2171.330 3510.320 2174.110 3511.850 ;
        RECT 2531.330 3511.005 2534.110 3512.535 ;
        RECT 2891.330 3484.045 2894.110 3485.575 ;
        RECT 2891.330 3218.165 2894.110 3219.695 ;
        RECT 2891.330 2952.965 2894.110 2954.495 ;
        RECT 2891.330 2687.085 2894.110 2688.615 ;
        RECT 2891.330 2421.205 2894.110 2422.735 ;
        RECT 2351.330 2255.890 2354.110 2257.420 ;
        RECT 2366.860 2253.095 2367.200 2253.195 ;
        RECT 2383.445 2253.095 2383.785 2253.195 ;
        RECT 2400.030 2253.095 2400.370 2253.195 ;
        RECT 2416.615 2253.095 2416.955 2253.195 ;
        RECT 2433.195 2253.095 2433.535 2253.195 ;
        RECT 2366.860 2253.085 2367.220 2253.095 ;
        RECT 2383.445 2253.085 2383.805 2253.095 ;
        RECT 2400.030 2253.085 2400.390 2253.095 ;
        RECT 2416.615 2253.085 2416.975 2253.095 ;
        RECT 2433.195 2253.085 2433.555 2253.095 ;
        RECT 2366.420 2253.065 2367.220 2253.085 ;
        RECT 2383.005 2253.065 2383.805 2253.085 ;
        RECT 2399.590 2253.065 2400.390 2253.085 ;
        RECT 2416.175 2253.065 2416.975 2253.085 ;
        RECT 2432.755 2253.065 2433.555 2253.085 ;
        RECT 2366.420 2252.785 2367.225 2253.065 ;
        RECT 2383.005 2252.785 2383.810 2253.065 ;
        RECT 2399.590 2252.785 2400.395 2253.065 ;
        RECT 2416.175 2252.785 2416.980 2253.065 ;
        RECT 2432.755 2252.785 2433.560 2253.065 ;
        RECT 2366.880 2252.755 2367.225 2252.785 ;
        RECT 2383.465 2252.755 2383.810 2252.785 ;
        RECT 2400.050 2252.755 2400.395 2252.785 ;
        RECT 2416.635 2252.755 2416.980 2252.785 ;
        RECT 2433.215 2252.755 2433.560 2252.785 ;
        RECT 2366.890 2252.725 2367.225 2252.755 ;
        RECT 2383.475 2252.725 2383.810 2252.755 ;
        RECT 2400.060 2252.725 2400.395 2252.755 ;
        RECT 2416.645 2252.725 2416.980 2252.755 ;
        RECT 2433.225 2252.725 2433.560 2252.755 ;
        RECT 2351.330 2245.035 2354.110 2246.565 ;
        RECT 2704.390 2216.755 2705.970 2217.085 ;
        RECT 2714.050 2216.755 2715.630 2217.085 ;
        RECT 2723.710 2216.755 2725.290 2217.085 ;
        RECT 2733.370 2216.755 2734.950 2217.085 ;
        RECT 2704.390 2211.315 2705.970 2211.645 ;
        RECT 2714.050 2211.315 2715.630 2211.645 ;
        RECT 2723.710 2211.315 2725.290 2211.645 ;
        RECT 2733.370 2211.315 2734.950 2211.645 ;
        RECT 2704.390 2205.875 2705.970 2206.205 ;
        RECT 2714.050 2205.875 2715.630 2206.205 ;
        RECT 2723.710 2205.875 2725.290 2206.205 ;
        RECT 2733.370 2205.875 2734.950 2206.205 ;
        RECT 2704.390 2200.435 2705.970 2200.765 ;
        RECT 2714.050 2200.435 2715.630 2200.765 ;
        RECT 2723.710 2200.435 2725.290 2200.765 ;
        RECT 2733.370 2200.435 2734.950 2200.765 ;
        RECT 2704.390 2194.995 2705.970 2195.325 ;
        RECT 2714.050 2194.995 2715.630 2195.325 ;
        RECT 2723.710 2194.995 2725.290 2195.325 ;
        RECT 2733.370 2194.995 2734.950 2195.325 ;
        RECT 2704.390 2189.555 2705.970 2189.885 ;
        RECT 2714.050 2189.555 2715.630 2189.885 ;
        RECT 2723.710 2189.555 2725.290 2189.885 ;
        RECT 2733.370 2189.555 2734.950 2189.885 ;
        RECT 2704.390 2184.115 2705.970 2184.445 ;
        RECT 2714.050 2184.115 2715.630 2184.445 ;
        RECT 2723.710 2184.115 2725.290 2184.445 ;
        RECT 2733.370 2184.115 2734.950 2184.445 ;
        RECT 2704.390 2178.675 2705.970 2179.005 ;
        RECT 2714.050 2178.675 2715.630 2179.005 ;
        RECT 2723.710 2178.675 2725.290 2179.005 ;
        RECT 2733.370 2178.675 2734.950 2179.005 ;
        RECT 2704.390 2173.235 2705.970 2173.565 ;
        RECT 2714.050 2173.235 2715.630 2173.565 ;
        RECT 2723.710 2173.235 2725.290 2173.565 ;
        RECT 2733.370 2173.235 2734.950 2173.565 ;
        RECT 2704.390 2167.795 2705.970 2168.125 ;
        RECT 2714.050 2167.795 2715.630 2168.125 ;
        RECT 2723.710 2167.795 2725.290 2168.125 ;
        RECT 2733.370 2167.795 2734.950 2168.125 ;
        RECT 2351.330 2163.895 2354.110 2165.425 ;
        RECT 2704.390 2162.355 2705.970 2162.685 ;
        RECT 2714.050 2162.355 2715.630 2162.685 ;
        RECT 2723.710 2162.355 2725.290 2162.685 ;
        RECT 2733.370 2162.355 2734.950 2162.685 ;
        RECT 2366.995 2160.400 2367.325 2160.415 ;
        RECT 2384.215 2160.400 2384.545 2160.415 ;
        RECT 2401.435 2160.400 2401.765 2160.415 ;
        RECT 2418.655 2160.400 2418.985 2160.415 ;
        RECT 2435.875 2160.400 2436.205 2160.415 ;
        RECT 2366.525 2160.100 2367.325 2160.400 ;
        RECT 2383.745 2160.100 2384.545 2160.400 ;
        RECT 2400.965 2160.100 2401.765 2160.400 ;
        RECT 2418.185 2160.100 2418.985 2160.400 ;
        RECT 2435.405 2160.100 2436.205 2160.400 ;
        RECT 2366.995 2160.085 2367.325 2160.100 ;
        RECT 2384.215 2160.085 2384.545 2160.100 ;
        RECT 2401.435 2160.085 2401.765 2160.100 ;
        RECT 2418.655 2160.085 2418.985 2160.100 ;
        RECT 2435.875 2160.085 2436.205 2160.100 ;
        RECT 2704.390 2156.915 2705.970 2157.245 ;
        RECT 2714.050 2156.915 2715.630 2157.245 ;
        RECT 2723.710 2156.915 2725.290 2157.245 ;
        RECT 2733.370 2156.915 2734.950 2157.245 ;
        RECT 2891.330 2156.005 2894.110 2157.535 ;
        RECT 2351.330 2153.035 2354.110 2154.565 ;
        RECT 2704.390 2151.475 2705.970 2151.805 ;
        RECT 2714.050 2151.475 2715.630 2151.805 ;
        RECT 2723.710 2151.475 2725.290 2151.805 ;
        RECT 2733.370 2151.475 2734.950 2151.805 ;
        RECT 2704.390 2146.035 2705.970 2146.365 ;
        RECT 2714.050 2146.035 2715.630 2146.365 ;
        RECT 2723.710 2146.035 2725.290 2146.365 ;
        RECT 2733.370 2146.035 2734.950 2146.365 ;
        RECT 2704.390 2140.595 2705.970 2140.925 ;
        RECT 2714.050 2140.595 2715.630 2140.925 ;
        RECT 2723.710 2140.595 2725.290 2140.925 ;
        RECT 2733.370 2140.595 2734.950 2140.925 ;
        RECT 2704.390 2135.155 2705.970 2135.485 ;
        RECT 2714.050 2135.155 2715.630 2135.485 ;
        RECT 2723.710 2135.155 2725.290 2135.485 ;
        RECT 2733.370 2135.155 2734.950 2135.485 ;
        RECT 2531.330 2132.630 2534.110 2134.160 ;
        RECT 2704.390 2129.715 2705.970 2130.045 ;
        RECT 2714.050 2129.715 2715.630 2130.045 ;
        RECT 2723.710 2129.715 2725.290 2130.045 ;
        RECT 2733.370 2129.715 2734.950 2130.045 ;
        RECT 2531.330 2125.100 2534.110 2126.630 ;
        RECT 2531.330 2119.120 2534.110 2120.650 ;
        RECT 2531.330 2113.175 2534.110 2114.705 ;
        RECT 2531.330 2107.530 2534.110 2109.060 ;
        RECT 2531.330 2101.525 2534.110 2103.055 ;
        RECT 2351.330 2058.895 2354.110 2060.425 ;
        RECT 2370.430 2052.595 2370.760 2052.995 ;
        RECT 2386.755 2052.595 2387.085 2052.995 ;
        RECT 2403.080 2052.595 2403.410 2052.995 ;
        RECT 2419.405 2052.595 2419.735 2052.995 ;
        RECT 2435.730 2052.595 2436.060 2052.995 ;
        RECT 2370.425 2052.265 2370.760 2052.595 ;
        RECT 2386.750 2052.265 2387.085 2052.595 ;
        RECT 2403.075 2052.265 2403.410 2052.595 ;
        RECT 2419.400 2052.265 2419.735 2052.595 ;
        RECT 2435.725 2052.265 2436.060 2052.595 ;
        RECT 2351.330 2048.035 2354.110 2049.565 ;
        RECT 2704.390 2036.755 2705.970 2037.085 ;
        RECT 2714.050 2036.755 2715.630 2037.085 ;
        RECT 2723.710 2036.755 2725.290 2037.085 ;
        RECT 2733.370 2036.755 2734.950 2037.085 ;
        RECT 2704.390 2031.315 2705.970 2031.645 ;
        RECT 2714.050 2031.315 2715.630 2031.645 ;
        RECT 2723.710 2031.315 2725.290 2031.645 ;
        RECT 2733.370 2031.315 2734.950 2031.645 ;
        RECT 2704.390 2025.875 2705.970 2026.205 ;
        RECT 2714.050 2025.875 2715.630 2026.205 ;
        RECT 2723.710 2025.875 2725.290 2026.205 ;
        RECT 2733.370 2025.875 2734.950 2026.205 ;
        RECT 2704.390 2020.435 2705.970 2020.765 ;
        RECT 2714.050 2020.435 2715.630 2020.765 ;
        RECT 2723.710 2020.435 2725.290 2020.765 ;
        RECT 2733.370 2020.435 2734.950 2020.765 ;
        RECT 2704.390 2014.995 2705.970 2015.325 ;
        RECT 2714.050 2014.995 2715.630 2015.325 ;
        RECT 2723.710 2014.995 2725.290 2015.325 ;
        RECT 2733.370 2014.995 2734.950 2015.325 ;
        RECT 2704.390 2009.555 2705.970 2009.885 ;
        RECT 2714.050 2009.555 2715.630 2009.885 ;
        RECT 2723.710 2009.555 2725.290 2009.885 ;
        RECT 2733.370 2009.555 2734.950 2009.885 ;
        RECT 2704.390 2004.115 2705.970 2004.445 ;
        RECT 2714.050 2004.115 2715.630 2004.445 ;
        RECT 2723.710 2004.115 2725.290 2004.445 ;
        RECT 2733.370 2004.115 2734.950 2004.445 ;
        RECT 2704.390 1998.675 2705.970 1999.005 ;
        RECT 2714.050 1998.675 2715.630 1999.005 ;
        RECT 2723.710 1998.675 2725.290 1999.005 ;
        RECT 2733.370 1998.675 2734.950 1999.005 ;
        RECT 2704.390 1993.235 2705.970 1993.565 ;
        RECT 2714.050 1993.235 2715.630 1993.565 ;
        RECT 2723.710 1993.235 2725.290 1993.565 ;
        RECT 2733.370 1993.235 2734.950 1993.565 ;
        RECT 2704.390 1987.795 2705.970 1988.125 ;
        RECT 2714.050 1987.795 2715.630 1988.125 ;
        RECT 2723.710 1987.795 2725.290 1988.125 ;
        RECT 2733.370 1987.795 2734.950 1988.125 ;
        RECT 2704.390 1982.355 2705.970 1982.685 ;
        RECT 2714.050 1982.355 2715.630 1982.685 ;
        RECT 2723.710 1982.355 2725.290 1982.685 ;
        RECT 2733.370 1982.355 2734.950 1982.685 ;
        RECT 2531.330 1980.375 2534.110 1981.905 ;
        RECT 2704.390 1976.915 2705.970 1977.245 ;
        RECT 2714.050 1976.915 2715.630 1977.245 ;
        RECT 2723.710 1976.915 2725.290 1977.245 ;
        RECT 2733.370 1976.915 2734.950 1977.245 ;
        RECT 2531.330 1972.845 2534.110 1974.375 ;
        RECT 2704.390 1971.475 2705.970 1971.805 ;
        RECT 2714.050 1971.475 2715.630 1971.805 ;
        RECT 2723.710 1971.475 2725.290 1971.805 ;
        RECT 2733.370 1971.475 2734.950 1971.805 ;
        RECT 2531.330 1966.865 2534.110 1968.395 ;
        RECT 2704.390 1966.035 2705.970 1966.365 ;
        RECT 2714.050 1966.035 2715.630 1966.365 ;
        RECT 2723.710 1966.035 2725.290 1966.365 ;
        RECT 2733.370 1966.035 2734.950 1966.365 ;
        RECT 2531.330 1960.920 2534.110 1962.450 ;
        RECT 2704.390 1960.595 2705.970 1960.925 ;
        RECT 2714.050 1960.595 2715.630 1960.925 ;
        RECT 2723.710 1960.595 2725.290 1960.925 ;
        RECT 2733.370 1960.595 2734.950 1960.925 ;
        RECT 2351.330 1953.900 2354.110 1955.430 ;
        RECT 2531.330 1955.275 2534.110 1956.805 ;
        RECT 2704.390 1955.155 2705.970 1955.485 ;
        RECT 2714.050 1955.155 2715.630 1955.485 ;
        RECT 2723.710 1955.155 2725.290 1955.485 ;
        RECT 2733.370 1955.155 2734.950 1955.485 ;
        RECT 2531.330 1949.270 2534.110 1950.800 ;
        RECT 2704.390 1949.715 2705.970 1950.045 ;
        RECT 2714.050 1949.715 2715.630 1950.045 ;
        RECT 2723.710 1949.715 2725.290 1950.045 ;
        RECT 2733.370 1949.715 2734.950 1950.045 ;
        RECT 2363.495 1947.035 2363.820 1947.040 ;
        RECT 2382.055 1947.035 2382.380 1947.040 ;
        RECT 2400.615 1947.035 2400.940 1947.040 ;
        RECT 2419.175 1947.035 2419.500 1947.040 ;
        RECT 2437.735 1947.035 2438.060 1947.040 ;
        RECT 2363.155 1946.705 2363.885 1947.035 ;
        RECT 2381.715 1946.705 2382.445 1947.035 ;
        RECT 2400.275 1946.705 2401.005 1947.035 ;
        RECT 2418.835 1946.705 2419.565 1947.035 ;
        RECT 2437.395 1946.705 2438.125 1947.035 ;
        RECT 2363.495 1946.700 2363.820 1946.705 ;
        RECT 2382.055 1946.700 2382.380 1946.705 ;
        RECT 2400.615 1946.700 2400.940 1946.705 ;
        RECT 2419.175 1946.700 2419.500 1946.705 ;
        RECT 2437.735 1946.700 2438.060 1946.705 ;
        RECT 2351.330 1943.035 2354.110 1944.565 ;
        RECT 2891.330 1890.125 2894.110 1891.655 ;
        RECT 2704.390 1856.755 2705.970 1857.085 ;
        RECT 2714.050 1856.755 2715.630 1857.085 ;
        RECT 2723.710 1856.755 2725.290 1857.085 ;
        RECT 2733.370 1856.755 2734.950 1857.085 ;
        RECT 2704.390 1851.315 2705.970 1851.645 ;
        RECT 2714.050 1851.315 2715.630 1851.645 ;
        RECT 2723.710 1851.315 2725.290 1851.645 ;
        RECT 2733.370 1851.315 2734.950 1851.645 ;
        RECT 2704.390 1845.875 2705.970 1846.205 ;
        RECT 2714.050 1845.875 2715.630 1846.205 ;
        RECT 2723.710 1845.875 2725.290 1846.205 ;
        RECT 2733.370 1845.875 2734.950 1846.205 ;
        RECT 2704.390 1840.435 2705.970 1840.765 ;
        RECT 2714.050 1840.435 2715.630 1840.765 ;
        RECT 2723.710 1840.435 2725.290 1840.765 ;
        RECT 2733.370 1840.435 2734.950 1840.765 ;
        RECT 2704.390 1834.995 2705.970 1835.325 ;
        RECT 2714.050 1834.995 2715.630 1835.325 ;
        RECT 2723.710 1834.995 2725.290 1835.325 ;
        RECT 2733.370 1834.995 2734.950 1835.325 ;
        RECT 2704.390 1829.555 2705.970 1829.885 ;
        RECT 2714.050 1829.555 2715.630 1829.885 ;
        RECT 2723.710 1829.555 2725.290 1829.885 ;
        RECT 2733.370 1829.555 2734.950 1829.885 ;
        RECT 2704.390 1824.115 2705.970 1824.445 ;
        RECT 2714.050 1824.115 2715.630 1824.445 ;
        RECT 2723.710 1824.115 2725.290 1824.445 ;
        RECT 2733.370 1824.115 2734.950 1824.445 ;
        RECT 2704.390 1818.675 2705.970 1819.005 ;
        RECT 2714.050 1818.675 2715.630 1819.005 ;
        RECT 2723.710 1818.675 2725.290 1819.005 ;
        RECT 2733.370 1818.675 2734.950 1819.005 ;
        RECT 2704.390 1813.235 2705.970 1813.565 ;
        RECT 2714.050 1813.235 2715.630 1813.565 ;
        RECT 2723.710 1813.235 2725.290 1813.565 ;
        RECT 2733.370 1813.235 2734.950 1813.565 ;
        RECT 2704.390 1807.795 2705.970 1808.125 ;
        RECT 2714.050 1807.795 2715.630 1808.125 ;
        RECT 2723.710 1807.795 2725.290 1808.125 ;
        RECT 2733.370 1807.795 2734.950 1808.125 ;
        RECT 2531.330 1803.405 2534.110 1804.935 ;
        RECT 2704.390 1802.355 2705.970 1802.685 ;
        RECT 2714.050 1802.355 2715.630 1802.685 ;
        RECT 2723.710 1802.355 2725.290 1802.685 ;
        RECT 2733.370 1802.355 2734.950 1802.685 ;
        RECT 2531.330 1795.875 2534.110 1797.405 ;
        RECT 2704.390 1796.915 2705.970 1797.245 ;
        RECT 2714.050 1796.915 2715.630 1797.245 ;
        RECT 2723.710 1796.915 2725.290 1797.245 ;
        RECT 2733.370 1796.915 2734.950 1797.245 ;
        RECT 2351.330 1790.900 2354.110 1792.430 ;
        RECT 2704.390 1791.475 2705.970 1791.805 ;
        RECT 2714.050 1791.475 2715.630 1791.805 ;
        RECT 2723.710 1791.475 2725.290 1791.805 ;
        RECT 2733.370 1791.475 2734.950 1791.805 ;
        RECT 2531.330 1789.895 2534.110 1791.425 ;
        RECT 2704.390 1786.035 2705.970 1786.365 ;
        RECT 2714.050 1786.035 2715.630 1786.365 ;
        RECT 2723.710 1786.035 2725.290 1786.365 ;
        RECT 2733.370 1786.035 2734.950 1786.365 ;
        RECT 2531.330 1783.950 2534.110 1785.480 ;
        RECT 2372.425 1783.475 2372.780 1783.480 ;
        RECT 2387.685 1783.475 2388.040 1783.480 ;
        RECT 2402.945 1783.475 2403.300 1783.480 ;
        RECT 2418.205 1783.475 2418.560 1783.480 ;
        RECT 2433.465 1783.475 2433.820 1783.480 ;
        RECT 2372.325 1783.145 2373.055 1783.475 ;
        RECT 2387.585 1783.145 2388.315 1783.475 ;
        RECT 2402.845 1783.145 2403.575 1783.475 ;
        RECT 2418.105 1783.145 2418.835 1783.475 ;
        RECT 2433.365 1783.145 2434.095 1783.475 ;
        RECT 2351.330 1780.035 2354.110 1781.565 ;
        RECT 2704.390 1780.595 2705.970 1780.925 ;
        RECT 2714.050 1780.595 2715.630 1780.925 ;
        RECT 2723.710 1780.595 2725.290 1780.925 ;
        RECT 2733.370 1780.595 2734.950 1780.925 ;
        RECT 2531.330 1778.305 2534.110 1779.835 ;
        RECT 2704.390 1775.155 2705.970 1775.485 ;
        RECT 2714.050 1775.155 2715.630 1775.485 ;
        RECT 2723.710 1775.155 2725.290 1775.485 ;
        RECT 2733.370 1775.155 2734.950 1775.485 ;
        RECT 2704.390 1769.715 2705.970 1770.045 ;
        RECT 2714.050 1769.715 2715.630 1770.045 ;
        RECT 2723.710 1769.715 2725.290 1770.045 ;
        RECT 2733.370 1769.715 2734.950 1770.045 ;
        RECT 2531.330 1766.835 2534.110 1768.365 ;
        RECT 2351.330 1710.895 2354.110 1712.425 ;
        RECT 2367.220 1708.095 2367.560 1708.195 ;
        RECT 2383.805 1708.095 2384.145 1708.195 ;
        RECT 2400.390 1708.100 2400.730 1708.200 ;
        RECT 2416.975 1708.105 2417.315 1708.205 ;
        RECT 2433.555 1708.105 2433.895 1708.205 ;
        RECT 2367.220 1708.085 2367.580 1708.095 ;
        RECT 2383.805 1708.085 2384.165 1708.095 ;
        RECT 2400.390 1708.090 2400.750 1708.100 ;
        RECT 2416.975 1708.095 2417.335 1708.105 ;
        RECT 2433.555 1708.095 2433.915 1708.105 ;
        RECT 2366.780 1708.065 2367.580 1708.085 ;
        RECT 2383.365 1708.065 2384.165 1708.085 ;
        RECT 2399.950 1708.070 2400.750 1708.090 ;
        RECT 2416.535 1708.075 2417.335 1708.095 ;
        RECT 2433.115 1708.075 2433.915 1708.095 ;
        RECT 2366.780 1707.785 2367.585 1708.065 ;
        RECT 2383.365 1707.785 2384.170 1708.065 ;
        RECT 2399.950 1707.790 2400.755 1708.070 ;
        RECT 2416.535 1707.795 2417.340 1708.075 ;
        RECT 2433.115 1707.795 2433.920 1708.075 ;
        RECT 2367.240 1707.755 2367.585 1707.785 ;
        RECT 2383.825 1707.755 2384.170 1707.785 ;
        RECT 2400.410 1707.760 2400.755 1707.790 ;
        RECT 2416.995 1707.765 2417.340 1707.795 ;
        RECT 2433.575 1707.765 2433.920 1707.795 ;
        RECT 2367.250 1707.725 2367.585 1707.755 ;
        RECT 2383.835 1707.725 2384.170 1707.755 ;
        RECT 2400.420 1707.730 2400.755 1707.760 ;
        RECT 2417.005 1707.735 2417.340 1707.765 ;
        RECT 2433.585 1707.735 2433.920 1707.765 ;
        RECT 2351.330 1700.035 2354.110 1701.565 ;
        RECT 2704.390 1676.755 2705.970 1677.085 ;
        RECT 2714.050 1676.755 2715.630 1677.085 ;
        RECT 2723.710 1676.755 2725.290 1677.085 ;
        RECT 2733.370 1676.755 2734.950 1677.085 ;
        RECT 2704.390 1671.315 2705.970 1671.645 ;
        RECT 2714.050 1671.315 2715.630 1671.645 ;
        RECT 2723.710 1671.315 2725.290 1671.645 ;
        RECT 2733.370 1671.315 2734.950 1671.645 ;
        RECT 2704.390 1665.875 2705.970 1666.205 ;
        RECT 2714.050 1665.875 2715.630 1666.205 ;
        RECT 2723.710 1665.875 2725.290 1666.205 ;
        RECT 2733.370 1665.875 2734.950 1666.205 ;
        RECT 2704.390 1660.435 2705.970 1660.765 ;
        RECT 2714.050 1660.435 2715.630 1660.765 ;
        RECT 2723.710 1660.435 2725.290 1660.765 ;
        RECT 2733.370 1660.435 2734.950 1660.765 ;
        RECT 2704.390 1654.995 2705.970 1655.325 ;
        RECT 2714.050 1654.995 2715.630 1655.325 ;
        RECT 2723.710 1654.995 2725.290 1655.325 ;
        RECT 2733.370 1654.995 2734.950 1655.325 ;
        RECT 2704.390 1649.555 2705.970 1649.885 ;
        RECT 2714.050 1649.555 2715.630 1649.885 ;
        RECT 2723.710 1649.555 2725.290 1649.885 ;
        RECT 2733.370 1649.555 2734.950 1649.885 ;
        RECT 2704.390 1644.115 2705.970 1644.445 ;
        RECT 2714.050 1644.115 2715.630 1644.445 ;
        RECT 2723.710 1644.115 2725.290 1644.445 ;
        RECT 2733.370 1644.115 2734.950 1644.445 ;
        RECT 2704.390 1638.675 2705.970 1639.005 ;
        RECT 2714.050 1638.675 2715.630 1639.005 ;
        RECT 2723.710 1638.675 2725.290 1639.005 ;
        RECT 2733.370 1638.675 2734.950 1639.005 ;
        RECT 2704.390 1633.235 2705.970 1633.565 ;
        RECT 2714.050 1633.235 2715.630 1633.565 ;
        RECT 2723.710 1633.235 2725.290 1633.565 ;
        RECT 2733.370 1633.235 2734.950 1633.565 ;
        RECT 2704.390 1627.795 2705.970 1628.125 ;
        RECT 2714.050 1627.795 2715.630 1628.125 ;
        RECT 2723.710 1627.795 2725.290 1628.125 ;
        RECT 2733.370 1627.795 2734.950 1628.125 ;
        RECT 2891.330 1624.245 2894.110 1625.775 ;
        RECT 2531.330 1622.270 2534.110 1623.800 ;
        RECT 2704.390 1622.355 2705.970 1622.685 ;
        RECT 2714.050 1622.355 2715.630 1622.685 ;
        RECT 2723.710 1622.355 2725.290 1622.685 ;
        RECT 2733.370 1622.355 2734.950 1622.685 ;
        RECT 2531.330 1615.855 2534.110 1617.385 ;
        RECT 2704.390 1616.915 2705.970 1617.245 ;
        RECT 2714.050 1616.915 2715.630 1617.245 ;
        RECT 2723.710 1616.915 2725.290 1617.245 ;
        RECT 2733.370 1616.915 2734.950 1617.245 ;
        RECT 2351.330 1610.895 2354.110 1612.425 ;
        RECT 2704.390 1611.475 2705.970 1611.805 ;
        RECT 2714.050 1611.475 2715.630 1611.805 ;
        RECT 2723.710 1611.475 2725.290 1611.805 ;
        RECT 2733.370 1611.475 2734.950 1611.805 ;
        RECT 2366.970 1607.400 2367.300 1607.415 ;
        RECT 2384.190 1607.400 2384.520 1607.415 ;
        RECT 2401.410 1607.405 2401.740 1607.420 ;
        RECT 2366.500 1607.100 2367.300 1607.400 ;
        RECT 2383.720 1607.100 2384.520 1607.400 ;
        RECT 2400.940 1607.105 2401.740 1607.405 ;
        RECT 2418.630 1607.400 2418.960 1607.415 ;
        RECT 2435.850 1607.400 2436.180 1607.415 ;
        RECT 2366.970 1607.085 2367.300 1607.100 ;
        RECT 2384.190 1607.085 2384.520 1607.100 ;
        RECT 2401.410 1607.090 2401.740 1607.105 ;
        RECT 2418.160 1607.100 2418.960 1607.400 ;
        RECT 2435.380 1607.100 2436.180 1607.400 ;
        RECT 2418.630 1607.085 2418.960 1607.100 ;
        RECT 2435.850 1607.085 2436.180 1607.100 ;
        RECT 2704.390 1606.035 2705.970 1606.365 ;
        RECT 2714.050 1606.035 2715.630 1606.365 ;
        RECT 2723.710 1606.035 2725.290 1606.365 ;
        RECT 2733.370 1606.035 2734.950 1606.365 ;
        RECT 2351.330 1600.035 2354.110 1601.565 ;
        RECT 2704.390 1600.595 2705.970 1600.925 ;
        RECT 2714.050 1600.595 2715.630 1600.925 ;
        RECT 2723.710 1600.595 2725.290 1600.925 ;
        RECT 2733.370 1600.595 2734.950 1600.925 ;
        RECT 2704.390 1595.155 2705.970 1595.485 ;
        RECT 2714.050 1595.155 2715.630 1595.485 ;
        RECT 2723.710 1595.155 2725.290 1595.485 ;
        RECT 2733.370 1595.155 2734.950 1595.485 ;
        RECT 2704.390 1589.715 2705.970 1590.045 ;
        RECT 2714.050 1589.715 2715.630 1590.045 ;
        RECT 2723.710 1589.715 2725.290 1590.045 ;
        RECT 2733.370 1589.715 2734.950 1590.045 ;
        RECT 2531.330 1586.610 2534.110 1588.140 ;
        RECT 2531.330 1579.080 2534.110 1580.610 ;
        RECT 2531.330 1573.100 2534.110 1574.630 ;
        RECT 2531.330 1564.685 2534.110 1566.215 ;
        RECT 2351.330 1533.895 2354.110 1535.425 ;
        RECT 2370.425 1527.485 2370.755 1527.885 ;
        RECT 2386.750 1527.485 2387.080 1527.885 ;
        RECT 2403.075 1527.485 2403.405 1527.885 ;
        RECT 2419.400 1527.485 2419.730 1527.885 ;
        RECT 2435.725 1527.485 2436.055 1527.885 ;
        RECT 2370.420 1527.155 2370.755 1527.485 ;
        RECT 2386.745 1527.155 2387.080 1527.485 ;
        RECT 2403.070 1527.155 2403.405 1527.485 ;
        RECT 2419.395 1527.155 2419.730 1527.485 ;
        RECT 2435.720 1527.155 2436.055 1527.485 ;
        RECT 2351.330 1523.035 2354.110 1524.565 ;
        RECT 2704.390 1496.755 2705.970 1497.085 ;
        RECT 2714.050 1496.755 2715.630 1497.085 ;
        RECT 2723.710 1496.755 2725.290 1497.085 ;
        RECT 2733.370 1496.755 2734.950 1497.085 ;
        RECT 2704.390 1491.315 2705.970 1491.645 ;
        RECT 2714.050 1491.315 2715.630 1491.645 ;
        RECT 2723.710 1491.315 2725.290 1491.645 ;
        RECT 2733.370 1491.315 2734.950 1491.645 ;
        RECT 2704.390 1485.875 2705.970 1486.205 ;
        RECT 2714.050 1485.875 2715.630 1486.205 ;
        RECT 2723.710 1485.875 2725.290 1486.205 ;
        RECT 2733.370 1485.875 2734.950 1486.205 ;
        RECT 2704.390 1480.435 2705.970 1480.765 ;
        RECT 2714.050 1480.435 2715.630 1480.765 ;
        RECT 2723.710 1480.435 2725.290 1480.765 ;
        RECT 2733.370 1480.435 2734.950 1480.765 ;
        RECT 2704.390 1474.995 2705.970 1475.325 ;
        RECT 2714.050 1474.995 2715.630 1475.325 ;
        RECT 2723.710 1474.995 2725.290 1475.325 ;
        RECT 2733.370 1474.995 2734.950 1475.325 ;
        RECT 2704.390 1469.555 2705.970 1469.885 ;
        RECT 2714.050 1469.555 2715.630 1469.885 ;
        RECT 2723.710 1469.555 2725.290 1469.885 ;
        RECT 2733.370 1469.555 2734.950 1469.885 ;
        RECT 2704.390 1464.115 2705.970 1464.445 ;
        RECT 2714.050 1464.115 2715.630 1464.445 ;
        RECT 2723.710 1464.115 2725.290 1464.445 ;
        RECT 2733.370 1464.115 2734.950 1464.445 ;
        RECT 2704.390 1458.675 2705.970 1459.005 ;
        RECT 2714.050 1458.675 2715.630 1459.005 ;
        RECT 2723.710 1458.675 2725.290 1459.005 ;
        RECT 2733.370 1458.675 2734.950 1459.005 ;
        RECT 2704.390 1453.235 2705.970 1453.565 ;
        RECT 2714.050 1453.235 2715.630 1453.565 ;
        RECT 2723.710 1453.235 2725.290 1453.565 ;
        RECT 2733.370 1453.235 2734.950 1453.565 ;
        RECT 2704.390 1447.795 2705.970 1448.125 ;
        RECT 2714.050 1447.795 2715.630 1448.125 ;
        RECT 2723.710 1447.795 2725.290 1448.125 ;
        RECT 2733.370 1447.795 2734.950 1448.125 ;
        RECT 2704.390 1442.355 2705.970 1442.685 ;
        RECT 2714.050 1442.355 2715.630 1442.685 ;
        RECT 2723.710 1442.355 2725.290 1442.685 ;
        RECT 2733.370 1442.355 2734.950 1442.685 ;
        RECT 2351.330 1435.900 2354.110 1437.430 ;
        RECT 2704.390 1436.915 2705.970 1437.245 ;
        RECT 2714.050 1436.915 2715.630 1437.245 ;
        RECT 2723.710 1436.915 2725.290 1437.245 ;
        RECT 2733.370 1436.915 2734.950 1437.245 ;
        RECT 2531.330 1434.985 2534.110 1436.515 ;
        RECT 2704.390 1431.475 2705.970 1431.805 ;
        RECT 2714.050 1431.475 2715.630 1431.805 ;
        RECT 2723.710 1431.475 2725.290 1431.805 ;
        RECT 2733.370 1431.475 2734.950 1431.805 ;
        RECT 2363.490 1429.035 2363.815 1429.040 ;
        RECT 2382.050 1429.035 2382.375 1429.040 ;
        RECT 2400.610 1429.035 2400.935 1429.040 ;
        RECT 2419.170 1429.035 2419.495 1429.040 ;
        RECT 2437.730 1429.035 2438.055 1429.040 ;
        RECT 2363.150 1428.705 2363.880 1429.035 ;
        RECT 2381.710 1428.705 2382.440 1429.035 ;
        RECT 2400.270 1428.705 2401.000 1429.035 ;
        RECT 2418.830 1428.705 2419.560 1429.035 ;
        RECT 2437.390 1428.705 2438.120 1429.035 ;
        RECT 2363.490 1428.700 2363.815 1428.705 ;
        RECT 2382.050 1428.700 2382.375 1428.705 ;
        RECT 2400.610 1428.700 2400.935 1428.705 ;
        RECT 2419.170 1428.700 2419.495 1428.705 ;
        RECT 2437.730 1428.700 2438.055 1428.705 ;
        RECT 2531.330 1428.570 2534.110 1430.100 ;
        RECT 2351.330 1425.035 2354.110 1426.565 ;
        RECT 2704.390 1426.035 2705.970 1426.365 ;
        RECT 2714.050 1426.035 2715.630 1426.365 ;
        RECT 2723.710 1426.035 2725.290 1426.365 ;
        RECT 2733.370 1426.035 2734.950 1426.365 ;
        RECT 2704.390 1420.595 2705.970 1420.925 ;
        RECT 2714.050 1420.595 2715.630 1420.925 ;
        RECT 2723.710 1420.595 2725.290 1420.925 ;
        RECT 2733.370 1420.595 2734.950 1420.925 ;
        RECT 2531.330 1414.380 2534.110 1415.910 ;
        RECT 2704.390 1415.155 2705.970 1415.485 ;
        RECT 2714.050 1415.155 2715.630 1415.485 ;
        RECT 2723.710 1415.155 2725.290 1415.485 ;
        RECT 2733.370 1415.155 2734.950 1415.485 ;
        RECT 2704.390 1409.715 2705.970 1410.045 ;
        RECT 2714.050 1409.715 2715.630 1410.045 ;
        RECT 2723.710 1409.715 2725.290 1410.045 ;
        RECT 2733.370 1409.715 2734.950 1410.045 ;
        RECT 2531.330 1406.850 2534.110 1408.380 ;
        RECT 2531.330 1400.870 2534.110 1402.400 ;
        RECT 2531.330 1392.455 2534.110 1393.985 ;
        RECT 2891.330 1359.045 2894.110 1360.575 ;
        RECT 2351.330 1335.900 2354.110 1337.430 ;
        RECT 2372.475 1328.475 2372.830 1328.480 ;
        RECT 2387.735 1328.475 2388.090 1328.480 ;
        RECT 2402.995 1328.475 2403.350 1328.480 ;
        RECT 2418.255 1328.475 2418.610 1328.480 ;
        RECT 2433.515 1328.475 2433.870 1328.480 ;
        RECT 2372.375 1328.145 2373.105 1328.475 ;
        RECT 2387.635 1328.145 2388.365 1328.475 ;
        RECT 2402.895 1328.145 2403.625 1328.475 ;
        RECT 2418.155 1328.145 2418.885 1328.475 ;
        RECT 2433.415 1328.145 2434.145 1328.475 ;
        RECT 2351.330 1325.035 2354.110 1326.565 ;
        RECT 2891.330 1159.805 2894.110 1161.335 ;
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
        RECT 11.170 -38.270 14.270 3557.950 ;
        RECT 191.170 -38.270 194.270 3557.950 ;
        RECT 371.170 -38.270 374.270 3557.950 ;
        RECT 551.170 -38.270 554.270 3557.950 ;
        RECT 731.170 -38.270 734.270 3557.950 ;
        RECT 911.170 -38.270 914.270 3557.950 ;
        RECT 1091.170 -38.270 1094.270 3557.950 ;
        RECT 1271.170 -38.270 1274.270 3557.950 ;
        RECT 1451.170 -38.270 1454.270 3557.950 ;
        RECT 1631.170 -38.270 1634.270 3557.950 ;
        RECT 1811.170 -38.270 1814.270 3557.950 ;
        RECT 1991.170 -38.270 1994.270 3557.950 ;
        RECT 2171.170 -38.270 2174.270 3557.950 ;
        RECT 2351.170 -38.270 2354.270 3557.950 ;
        RECT 2531.170 -38.270 2534.270 3557.950 ;
        RECT 2711.170 2227.860 2714.270 3557.950 ;
        RECT 2704.380 2129.640 2705.980 2217.160 ;
        RECT 2714.040 2129.640 2715.640 2217.160 ;
        RECT 2723.700 2129.640 2725.300 2217.160 ;
        RECT 2733.360 2129.640 2734.960 2217.160 ;
        RECT 2704.380 1949.640 2705.980 2037.160 ;
        RECT 2714.040 1949.640 2715.640 2037.160 ;
        RECT 2723.700 1949.640 2725.300 2037.160 ;
        RECT 2733.360 1949.640 2734.960 2037.160 ;
        RECT 2704.380 1769.640 2705.980 1857.160 ;
        RECT 2714.040 1769.640 2715.640 1857.160 ;
        RECT 2723.700 1769.640 2725.300 1857.160 ;
        RECT 2733.360 1769.640 2734.960 1857.160 ;
        RECT 2704.380 1589.640 2705.980 1677.160 ;
        RECT 2714.040 1589.640 2715.640 1677.160 ;
        RECT 2723.700 1589.640 2725.300 1677.160 ;
        RECT 2733.360 1589.640 2734.960 1677.160 ;
        RECT 2704.380 1409.640 2705.980 1497.160 ;
        RECT 2714.040 1409.640 2715.640 1497.160 ;
        RECT 2723.700 1409.640 2725.300 1497.160 ;
        RECT 2733.360 1409.640 2734.960 1497.160 ;
        RECT 2711.170 -38.270 2714.270 1398.940 ;
        RECT 2891.170 -38.270 2894.270 3557.950 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
        RECT -43.630 3436.530 2963.250 3439.630 ;
        RECT -43.630 3256.530 2963.250 3259.630 ;
        RECT -43.630 3076.530 2963.250 3079.630 ;
        RECT -43.630 2896.530 2963.250 2899.630 ;
        RECT -43.630 2716.530 2963.250 2719.630 ;
        RECT -43.630 2536.530 2963.250 2539.630 ;
        RECT -43.630 2356.530 2963.250 2359.630 ;
        RECT -43.630 2176.530 2963.250 2179.630 ;
        RECT -43.630 1996.530 2963.250 1999.630 ;
        RECT -43.630 1816.530 2963.250 1819.630 ;
        RECT -43.630 1636.530 2963.250 1639.630 ;
        RECT -43.630 1456.530 2963.250 1459.630 ;
        RECT -43.630 1276.530 2963.250 1279.630 ;
        RECT -43.630 1096.530 2963.250 1099.630 ;
        RECT -43.630 916.530 2963.250 919.630 ;
        RECT -43.630 736.530 2963.250 739.630 ;
        RECT -43.630 556.530 2963.250 559.630 ;
        RECT -43.630 376.530 2963.250 379.630 ;
        RECT -43.630 196.530 2963.250 199.630 ;
        RECT -43.630 16.530 2963.250 19.630 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
        RECT 23.570 -38.270 26.670 3557.950 ;
        RECT 203.570 -38.270 206.670 3557.950 ;
        RECT 383.570 -38.270 386.670 3557.950 ;
        RECT 563.570 -38.270 566.670 3557.950 ;
        RECT 743.570 -38.270 746.670 3557.950 ;
        RECT 923.570 -38.270 926.670 3557.950 ;
        RECT 1103.570 -38.270 1106.670 3557.950 ;
        RECT 1283.570 -38.270 1286.670 3557.950 ;
        RECT 1463.570 -38.270 1466.670 3557.950 ;
        RECT 1643.570 -38.270 1646.670 3557.950 ;
        RECT 1823.570 -38.270 1826.670 3557.950 ;
        RECT 2003.570 -38.270 2006.670 3557.950 ;
        RECT 2183.570 -38.270 2186.670 3557.950 ;
        RECT 2363.570 1795.300 2366.670 3557.950 ;
        RECT 2363.570 1340.300 2366.670 1773.075 ;
        RECT 2363.570 -38.270 2366.670 1318.075 ;
        RECT 2543.570 -38.270 2546.670 3557.950 ;
        RECT 2723.570 2227.860 2726.670 3557.950 ;
        RECT 2723.570 -38.270 2726.670 1398.940 ;
        RECT 2903.570 -38.270 2906.670 3557.950 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
        RECT -43.630 3448.930 2963.250 3452.030 ;
        RECT -43.630 3268.930 2963.250 3272.030 ;
        RECT -43.630 3088.930 2963.250 3092.030 ;
        RECT -43.630 2908.930 2963.250 2912.030 ;
        RECT -43.630 2728.930 2963.250 2732.030 ;
        RECT -43.630 2548.930 2963.250 2552.030 ;
        RECT -43.630 2368.930 2963.250 2372.030 ;
        RECT -43.630 2188.930 2963.250 2192.030 ;
        RECT -43.630 2008.930 2963.250 2012.030 ;
        RECT -43.630 1828.930 2963.250 1832.030 ;
        RECT -43.630 1648.930 2963.250 1652.030 ;
        RECT -43.630 1468.930 2963.250 1472.030 ;
        RECT -43.630 1288.930 2963.250 1292.030 ;
        RECT -43.630 1108.930 2963.250 1112.030 ;
        RECT -43.630 928.930 2963.250 932.030 ;
        RECT -43.630 748.930 2963.250 752.030 ;
        RECT -43.630 568.930 2963.250 572.030 ;
        RECT -43.630 388.930 2963.250 392.030 ;
        RECT -43.630 208.930 2963.250 212.030 ;
        RECT -43.630 28.930 2963.250 32.030 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER pwell ;
        RECT 1622.950 3512.755 1623.120 3512.925 ;
        RECT 1262.950 3512.305 1263.120 3512.475 ;
        RECT 2522.950 3511.160 2523.120 3511.330 ;
        RECT 1802.950 3510.835 1803.120 3511.005 ;
        RECT 2162.950 3510.475 2163.120 3510.645 ;
        RECT 2883.065 3485.420 2883.235 3485.590 ;
        RECT 2883.065 3219.540 2883.235 3219.710 ;
        RECT 2883.065 2954.340 2883.235 2954.510 ;
        RECT 2883.065 2688.460 2883.235 2688.630 ;
        RECT 2883.065 2422.580 2883.235 2422.750 ;
        RECT 2364.320 2253.335 2365.050 2253.745 ;
        RECT 2366.960 2253.495 2367.130 2253.525 ;
        RECT 2370.180 2253.495 2370.350 2253.525 ;
        RECT 2366.960 2253.335 2367.540 2253.495 ;
        RECT 2370.180 2253.385 2370.810 2253.495 ;
        RECT 2370.180 2253.335 2370.490 2253.385 ;
        RECT 2364.320 2253.145 2370.490 2253.335 ;
        RECT 2380.905 2253.335 2381.635 2253.745 ;
        RECT 2383.545 2253.495 2383.715 2253.525 ;
        RECT 2386.765 2253.495 2386.935 2253.525 ;
        RECT 2383.545 2253.335 2384.125 2253.495 ;
        RECT 2386.765 2253.385 2387.395 2253.495 ;
        RECT 2386.765 2253.335 2387.075 2253.385 ;
        RECT 2380.905 2253.145 2387.075 2253.335 ;
        RECT 2397.490 2253.335 2398.220 2253.745 ;
        RECT 2400.130 2253.495 2400.300 2253.525 ;
        RECT 2403.350 2253.495 2403.520 2253.525 ;
        RECT 2400.130 2253.335 2400.710 2253.495 ;
        RECT 2403.350 2253.385 2403.980 2253.495 ;
        RECT 2403.350 2253.335 2403.660 2253.385 ;
        RECT 2397.490 2253.145 2403.660 2253.335 ;
        RECT 2414.075 2253.335 2414.805 2253.745 ;
        RECT 2416.715 2253.495 2416.885 2253.525 ;
        RECT 2419.935 2253.495 2420.105 2253.525 ;
        RECT 2416.715 2253.335 2417.295 2253.495 ;
        RECT 2419.935 2253.385 2420.565 2253.495 ;
        RECT 2419.935 2253.335 2420.245 2253.385 ;
        RECT 2414.075 2253.145 2420.245 2253.335 ;
        RECT 2430.655 2253.335 2431.385 2253.745 ;
        RECT 2433.295 2253.495 2433.465 2253.525 ;
        RECT 2436.515 2253.495 2436.685 2253.525 ;
        RECT 2433.295 2253.335 2433.875 2253.495 ;
        RECT 2436.515 2253.385 2437.145 2253.495 ;
        RECT 2436.515 2253.335 2436.825 2253.385 ;
        RECT 2430.655 2253.145 2436.825 2253.335 ;
        RECT 2365.180 2252.515 2370.490 2253.145 ;
        RECT 2365.180 2252.425 2366.130 2252.515 ;
        RECT 2367.740 2252.425 2370.490 2252.515 ;
        RECT 2381.765 2252.515 2387.075 2253.145 ;
        RECT 2381.765 2252.425 2382.715 2252.515 ;
        RECT 2384.325 2252.425 2387.075 2252.515 ;
        RECT 2398.350 2252.515 2403.660 2253.145 ;
        RECT 2398.350 2252.425 2399.300 2252.515 ;
        RECT 2400.910 2252.425 2403.660 2252.515 ;
        RECT 2414.935 2252.515 2420.245 2253.145 ;
        RECT 2414.935 2252.425 2415.885 2252.515 ;
        RECT 2417.495 2252.425 2420.245 2252.515 ;
        RECT 2431.515 2252.515 2436.825 2253.145 ;
        RECT 2431.515 2252.425 2432.465 2252.515 ;
        RECT 2434.075 2252.425 2436.825 2252.515 ;
        RECT 2364.220 2248.815 2365.450 2249.015 ;
        RECT 2366.780 2248.815 2367.730 2249.015 ;
        RECT 2364.220 2248.790 2367.730 2248.815 ;
        RECT 2369.110 2248.790 2371.390 2249.015 ;
        RECT 2364.220 2248.305 2371.390 2248.790 ;
        RECT 2380.805 2248.815 2382.035 2249.015 ;
        RECT 2383.365 2248.815 2384.315 2249.015 ;
        RECT 2380.805 2248.790 2384.315 2248.815 ;
        RECT 2385.695 2248.790 2387.975 2249.015 ;
        RECT 2380.805 2248.305 2387.975 2248.790 ;
        RECT 2397.390 2248.815 2398.620 2249.015 ;
        RECT 2399.950 2248.815 2400.900 2249.015 ;
        RECT 2397.390 2248.790 2400.900 2248.815 ;
        RECT 2402.280 2248.790 2404.560 2249.015 ;
        RECT 2397.390 2248.305 2404.560 2248.790 ;
        RECT 2413.975 2248.815 2415.205 2249.015 ;
        RECT 2416.535 2248.815 2417.485 2249.015 ;
        RECT 2413.975 2248.790 2417.485 2248.815 ;
        RECT 2418.865 2248.790 2421.145 2249.015 ;
        RECT 2413.975 2248.305 2421.145 2248.790 ;
        RECT 2430.555 2248.815 2431.785 2249.015 ;
        RECT 2433.115 2248.815 2434.065 2249.015 ;
        RECT 2430.555 2248.790 2434.065 2248.815 ;
        RECT 2435.445 2248.790 2437.725 2249.015 ;
        RECT 2430.555 2248.305 2437.725 2248.790 ;
        RECT 2364.160 2248.135 2371.390 2248.305 ;
        RECT 2364.160 2247.705 2364.750 2248.135 ;
        RECT 2366.800 2248.110 2371.390 2248.135 ;
        RECT 2380.745 2248.135 2387.975 2248.305 ;
        RECT 2367.880 2247.925 2368.050 2248.105 ;
        RECT 2370.190 2248.095 2370.360 2248.105 ;
        RECT 2370.180 2248.085 2370.360 2248.095 ;
        RECT 2370.190 2247.925 2370.360 2248.085 ;
        RECT 2380.745 2247.705 2381.335 2248.135 ;
        RECT 2383.385 2248.110 2387.975 2248.135 ;
        RECT 2397.330 2248.135 2404.560 2248.305 ;
        RECT 2384.465 2247.925 2384.635 2248.105 ;
        RECT 2386.775 2248.095 2386.945 2248.105 ;
        RECT 2386.765 2248.085 2386.945 2248.095 ;
        RECT 2386.775 2247.925 2386.945 2248.085 ;
        RECT 2397.330 2247.705 2397.920 2248.135 ;
        RECT 2399.970 2248.110 2404.560 2248.135 ;
        RECT 2413.915 2248.135 2421.145 2248.305 ;
        RECT 2401.050 2247.925 2401.220 2248.105 ;
        RECT 2403.360 2248.095 2403.530 2248.105 ;
        RECT 2403.350 2248.085 2403.530 2248.095 ;
        RECT 2403.360 2247.925 2403.530 2248.085 ;
        RECT 2413.915 2247.705 2414.505 2248.135 ;
        RECT 2416.555 2248.110 2421.145 2248.135 ;
        RECT 2430.495 2248.135 2437.725 2248.305 ;
        RECT 2417.635 2247.925 2417.805 2248.105 ;
        RECT 2419.945 2248.095 2420.115 2248.105 ;
        RECT 2419.935 2248.085 2420.115 2248.095 ;
        RECT 2419.945 2247.925 2420.115 2248.085 ;
        RECT 2430.495 2247.705 2431.085 2248.135 ;
        RECT 2433.135 2248.110 2437.725 2248.135 ;
        RECT 2434.215 2247.925 2434.385 2248.105 ;
        RECT 2436.525 2248.095 2436.695 2248.105 ;
        RECT 2436.515 2248.085 2436.695 2248.095 ;
        RECT 2436.525 2247.925 2436.695 2248.085 ;
        RECT 2695.665 2216.815 2695.835 2217.005 ;
        RECT 2697.045 2216.815 2697.215 2217.005 ;
        RECT 2699.805 2216.815 2699.975 2217.005 ;
        RECT 2701.185 2216.815 2701.355 2217.005 ;
        RECT 2701.645 2216.815 2701.815 2217.005 ;
        RECT 2707.165 2216.815 2707.335 2217.005 ;
        RECT 2709.005 2216.815 2709.175 2217.005 ;
        RECT 2710.845 2216.815 2711.015 2217.005 ;
        RECT 2716.365 2216.815 2716.535 2217.005 ;
        RECT 2720.045 2216.815 2720.215 2217.005 ;
        RECT 2723.265 2216.815 2723.435 2217.005 ;
        RECT 2723.725 2216.815 2723.895 2217.005 ;
        RECT 2729.245 2216.815 2729.415 2217.005 ;
        RECT 2731.080 2216.865 2731.200 2216.975 ;
        RECT 2732.455 2216.815 2732.625 2217.005 ;
        RECT 2733.845 2216.815 2734.015 2217.005 ;
        RECT 2695.525 2216.005 2696.895 2216.815 ;
        RECT 2696.905 2216.135 2698.735 2216.815 ;
        RECT 2698.745 2216.035 2700.115 2216.815 ;
        RECT 2700.125 2216.035 2701.495 2216.815 ;
        RECT 2701.505 2216.005 2707.015 2216.815 ;
        RECT 2707.025 2216.005 2708.395 2216.815 ;
        RECT 2708.865 2216.135 2710.695 2216.815 ;
        RECT 2709.350 2215.905 2710.695 2216.135 ;
        RECT 2710.705 2216.005 2716.215 2216.815 ;
        RECT 2716.225 2216.005 2719.895 2216.815 ;
        RECT 2719.905 2216.005 2721.275 2216.815 ;
        RECT 2721.745 2216.135 2723.575 2216.815 ;
        RECT 2723.585 2216.005 2729.095 2216.815 ;
        RECT 2729.105 2216.005 2730.935 2216.815 ;
        RECT 2731.405 2216.035 2732.775 2216.815 ;
        RECT 2732.785 2216.005 2734.155 2216.815 ;
        RECT 2695.525 2211.585 2696.895 2212.395 ;
        RECT 2696.905 2211.585 2698.275 2212.365 ;
        RECT 2698.285 2211.585 2703.795 2212.395 ;
        RECT 2703.805 2211.585 2707.475 2212.395 ;
        RECT 2708.865 2211.585 2714.375 2212.395 ;
        RECT 2714.385 2211.585 2719.895 2212.395 ;
        RECT 2719.905 2211.585 2725.415 2212.395 ;
        RECT 2725.425 2211.585 2730.935 2212.395 ;
        RECT 2730.945 2211.585 2732.775 2212.395 ;
        RECT 2732.785 2211.585 2734.155 2212.395 ;
        RECT 2695.665 2211.375 2695.835 2211.585 ;
        RECT 2697.045 2211.375 2697.215 2211.585 ;
        RECT 2698.425 2211.395 2698.595 2211.585 ;
        RECT 2702.565 2211.375 2702.735 2211.565 ;
        RECT 2703.945 2211.395 2704.115 2211.585 ;
        RECT 2707.635 2211.430 2707.795 2211.540 ;
        RECT 2708.085 2211.375 2708.255 2211.565 ;
        RECT 2709.005 2211.395 2709.175 2211.585 ;
        RECT 2713.605 2211.375 2713.775 2211.565 ;
        RECT 2714.525 2211.395 2714.695 2211.585 ;
        RECT 2719.125 2211.375 2719.295 2211.565 ;
        RECT 2720.045 2211.395 2720.215 2211.585 ;
        RECT 2720.960 2211.425 2721.080 2211.535 ;
        RECT 2721.885 2211.375 2722.055 2211.565 ;
        RECT 2725.565 2211.395 2725.735 2211.585 ;
        RECT 2727.405 2211.375 2727.575 2211.565 ;
        RECT 2731.085 2211.395 2731.255 2211.585 ;
        RECT 2733.845 2211.375 2734.015 2211.585 ;
        RECT 2695.525 2210.565 2696.895 2211.375 ;
        RECT 2696.905 2210.565 2702.415 2211.375 ;
        RECT 2702.425 2210.565 2707.935 2211.375 ;
        RECT 2707.945 2210.565 2713.455 2211.375 ;
        RECT 2713.465 2210.565 2718.975 2211.375 ;
        RECT 2718.985 2210.565 2720.815 2211.375 ;
        RECT 2721.745 2210.565 2727.255 2211.375 ;
        RECT 2727.265 2210.565 2732.775 2211.375 ;
        RECT 2732.785 2210.565 2734.155 2211.375 ;
        RECT 2695.525 2206.145 2696.895 2206.955 ;
        RECT 2696.905 2206.145 2702.415 2206.955 ;
        RECT 2702.425 2206.145 2707.935 2206.955 ;
        RECT 2708.865 2206.145 2714.375 2206.955 ;
        RECT 2714.385 2206.145 2719.895 2206.955 ;
        RECT 2719.905 2206.145 2725.415 2206.955 ;
        RECT 2725.425 2206.145 2730.935 2206.955 ;
        RECT 2730.945 2206.145 2732.775 2206.955 ;
        RECT 2732.785 2206.145 2734.155 2206.955 ;
        RECT 2695.665 2205.935 2695.835 2206.145 ;
        RECT 2697.045 2205.935 2697.215 2206.145 ;
        RECT 2698.425 2205.935 2698.595 2206.125 ;
        RECT 2702.565 2205.955 2702.735 2206.145 ;
        RECT 2703.945 2205.935 2704.115 2206.125 ;
        RECT 2708.080 2205.985 2708.200 2206.095 ;
        RECT 2709.005 2205.955 2709.175 2206.145 ;
        RECT 2709.465 2205.935 2709.635 2206.125 ;
        RECT 2714.525 2205.955 2714.695 2206.145 ;
        RECT 2714.985 2205.935 2715.155 2206.125 ;
        RECT 2720.045 2205.955 2720.215 2206.145 ;
        RECT 2720.515 2205.980 2720.675 2206.090 ;
        RECT 2721.885 2205.935 2722.055 2206.125 ;
        RECT 2725.565 2205.955 2725.735 2206.145 ;
        RECT 2727.405 2205.935 2727.575 2206.125 ;
        RECT 2731.085 2205.955 2731.255 2206.145 ;
        RECT 2733.845 2205.935 2734.015 2206.145 ;
        RECT 2695.525 2205.125 2696.895 2205.935 ;
        RECT 2696.905 2205.155 2698.275 2205.935 ;
        RECT 2698.285 2205.125 2703.795 2205.935 ;
        RECT 2703.805 2205.125 2709.315 2205.935 ;
        RECT 2709.325 2205.125 2714.835 2205.935 ;
        RECT 2714.845 2205.125 2720.355 2205.935 ;
        RECT 2721.745 2205.125 2727.255 2205.935 ;
        RECT 2727.265 2205.125 2732.775 2205.935 ;
        RECT 2732.785 2205.125 2734.155 2205.935 ;
        RECT 2695.525 2200.705 2696.895 2201.515 ;
        RECT 2696.905 2200.705 2702.415 2201.515 ;
        RECT 2702.425 2200.705 2707.935 2201.515 ;
        RECT 2708.865 2200.705 2714.375 2201.515 ;
        RECT 2714.385 2200.705 2719.895 2201.515 ;
        RECT 2719.905 2200.705 2725.415 2201.515 ;
        RECT 2725.425 2200.705 2730.935 2201.515 ;
        RECT 2730.945 2200.705 2732.775 2201.515 ;
        RECT 2732.785 2200.705 2734.155 2201.515 ;
        RECT 2695.665 2200.495 2695.835 2200.705 ;
        RECT 2697.045 2200.495 2697.215 2200.705 ;
        RECT 2702.565 2200.515 2702.735 2200.705 ;
        RECT 2706.705 2200.495 2706.875 2200.685 ;
        RECT 2708.080 2200.545 2708.200 2200.655 ;
        RECT 2709.005 2200.515 2709.175 2200.705 ;
        RECT 2712.225 2200.495 2712.395 2200.685 ;
        RECT 2714.525 2200.515 2714.695 2200.705 ;
        RECT 2717.745 2200.495 2717.915 2200.685 ;
        RECT 2720.045 2200.515 2720.215 2200.705 ;
        RECT 2721.885 2200.495 2722.055 2200.685 ;
        RECT 2725.565 2200.515 2725.735 2200.705 ;
        RECT 2727.405 2200.495 2727.575 2200.685 ;
        RECT 2731.085 2200.515 2731.255 2200.705 ;
        RECT 2733.845 2200.495 2734.015 2200.705 ;
        RECT 2695.525 2199.685 2696.895 2200.495 ;
        RECT 2696.905 2200.325 2698.665 2200.495 ;
        RECT 2696.905 2200.280 2699.160 2200.325 ;
        RECT 2696.905 2200.245 2700.100 2200.280 ;
        RECT 2701.460 2200.245 2706.555 2200.495 ;
        RECT 2696.905 2199.815 2706.555 2200.245 ;
        RECT 2698.230 2199.645 2701.460 2199.815 ;
        RECT 2699.170 2199.600 2701.460 2199.645 ;
        RECT 2700.110 2199.565 2701.460 2199.600 ;
        RECT 2704.535 2199.585 2706.555 2199.815 ;
        RECT 2706.565 2199.685 2712.075 2200.495 ;
        RECT 2712.085 2199.685 2717.595 2200.495 ;
        RECT 2717.605 2199.685 2721.275 2200.495 ;
        RECT 2721.745 2199.685 2727.255 2200.495 ;
        RECT 2727.265 2199.685 2732.775 2200.495 ;
        RECT 2732.785 2199.685 2734.155 2200.495 ;
        RECT 2704.535 2199.565 2705.455 2199.585 ;
        RECT 2695.525 2195.265 2696.895 2196.075 ;
        RECT 2696.905 2195.265 2698.275 2196.045 ;
        RECT 2698.285 2195.265 2703.795 2196.075 ;
        RECT 2703.805 2195.265 2707.475 2196.075 ;
        RECT 2708.865 2195.265 2714.375 2196.075 ;
        RECT 2714.385 2195.265 2719.895 2196.075 ;
        RECT 2719.905 2195.265 2725.415 2196.075 ;
        RECT 2725.425 2195.265 2730.935 2196.075 ;
        RECT 2730.945 2195.265 2732.775 2196.075 ;
        RECT 2732.785 2195.265 2734.155 2196.075 ;
        RECT 2695.665 2195.055 2695.835 2195.265 ;
        RECT 2697.045 2195.055 2697.215 2195.265 ;
        RECT 2698.425 2195.075 2698.595 2195.265 ;
        RECT 2703.945 2195.075 2704.115 2195.265 ;
        RECT 2706.705 2195.055 2706.875 2195.245 ;
        RECT 2707.635 2195.110 2707.795 2195.220 ;
        RECT 2709.005 2195.075 2709.175 2195.265 ;
        RECT 2712.225 2195.055 2712.395 2195.245 ;
        RECT 2714.525 2195.075 2714.695 2195.265 ;
        RECT 2717.745 2195.055 2717.915 2195.245 ;
        RECT 2720.045 2195.075 2720.215 2195.265 ;
        RECT 2721.885 2195.055 2722.055 2195.245 ;
        RECT 2725.565 2195.075 2725.735 2195.265 ;
        RECT 2727.405 2195.055 2727.575 2195.245 ;
        RECT 2731.085 2195.075 2731.255 2195.265 ;
        RECT 2733.845 2195.055 2734.015 2195.265 ;
        RECT 2695.525 2194.245 2696.895 2195.055 ;
        RECT 2696.905 2194.885 2698.665 2195.055 ;
        RECT 2696.905 2194.840 2699.160 2194.885 ;
        RECT 2696.905 2194.805 2700.100 2194.840 ;
        RECT 2701.460 2194.805 2706.555 2195.055 ;
        RECT 2696.905 2194.375 2706.555 2194.805 ;
        RECT 2698.230 2194.205 2701.460 2194.375 ;
        RECT 2699.170 2194.160 2701.460 2194.205 ;
        RECT 2700.110 2194.125 2701.460 2194.160 ;
        RECT 2704.535 2194.145 2706.555 2194.375 ;
        RECT 2706.565 2194.245 2712.075 2195.055 ;
        RECT 2712.085 2194.245 2717.595 2195.055 ;
        RECT 2717.605 2194.245 2721.275 2195.055 ;
        RECT 2721.745 2194.245 2727.255 2195.055 ;
        RECT 2727.265 2194.245 2732.775 2195.055 ;
        RECT 2732.785 2194.245 2734.155 2195.055 ;
        RECT 2704.535 2194.125 2705.455 2194.145 ;
        RECT 2695.525 2189.825 2696.895 2190.635 ;
        RECT 2696.905 2189.825 2698.275 2190.605 ;
        RECT 2698.285 2189.825 2701.035 2190.635 ;
        RECT 2701.505 2190.505 2702.435 2190.735 ;
        RECT 2701.505 2189.825 2705.405 2190.505 ;
        RECT 2705.645 2189.825 2708.395 2190.635 ;
        RECT 2708.865 2189.825 2714.375 2190.635 ;
        RECT 2714.385 2189.825 2719.895 2190.635 ;
        RECT 2719.905 2189.825 2725.415 2190.635 ;
        RECT 2725.425 2189.825 2730.935 2190.635 ;
        RECT 2730.945 2189.825 2732.775 2190.635 ;
        RECT 2732.785 2189.825 2734.155 2190.635 ;
        RECT 2695.665 2189.615 2695.835 2189.825 ;
        RECT 2697.045 2189.615 2697.215 2189.825 ;
        RECT 2698.425 2189.635 2698.595 2189.825 ;
        RECT 2701.180 2189.665 2701.300 2189.775 ;
        RECT 2701.920 2189.635 2702.090 2189.825 ;
        RECT 2702.565 2189.615 2702.735 2189.805 ;
        RECT 2705.785 2189.635 2705.955 2189.825 ;
        RECT 2708.085 2189.615 2708.255 2189.805 ;
        RECT 2709.005 2189.635 2709.175 2189.825 ;
        RECT 2713.605 2189.615 2713.775 2189.805 ;
        RECT 2714.525 2189.635 2714.695 2189.825 ;
        RECT 2719.125 2189.615 2719.295 2189.805 ;
        RECT 2720.045 2189.635 2720.215 2189.825 ;
        RECT 2720.960 2189.665 2721.080 2189.775 ;
        RECT 2721.885 2189.615 2722.055 2189.805 ;
        RECT 2725.565 2189.635 2725.735 2189.825 ;
        RECT 2727.405 2189.615 2727.575 2189.805 ;
        RECT 2731.085 2189.635 2731.255 2189.825 ;
        RECT 2733.845 2189.615 2734.015 2189.825 ;
        RECT 2695.525 2188.805 2696.895 2189.615 ;
        RECT 2696.905 2188.805 2702.415 2189.615 ;
        RECT 2702.425 2188.805 2707.935 2189.615 ;
        RECT 2707.945 2188.805 2713.455 2189.615 ;
        RECT 2713.465 2188.805 2718.975 2189.615 ;
        RECT 2718.985 2188.805 2720.815 2189.615 ;
        RECT 2721.745 2188.805 2727.255 2189.615 ;
        RECT 2727.265 2188.805 2732.775 2189.615 ;
        RECT 2732.785 2188.805 2734.155 2189.615 ;
        RECT 2695.525 2184.385 2696.895 2185.195 ;
        RECT 2696.905 2184.385 2698.275 2185.165 ;
        RECT 2698.285 2184.385 2703.795 2185.195 ;
        RECT 2703.805 2184.385 2707.475 2185.195 ;
        RECT 2708.865 2184.385 2714.375 2185.195 ;
        RECT 2714.385 2184.385 2719.895 2185.195 ;
        RECT 2719.905 2184.385 2725.415 2185.195 ;
        RECT 2725.425 2184.385 2730.935 2185.195 ;
        RECT 2730.945 2184.385 2732.775 2185.195 ;
        RECT 2732.785 2184.385 2734.155 2185.195 ;
        RECT 2695.665 2184.175 2695.835 2184.385 ;
        RECT 2697.045 2184.175 2697.215 2184.385 ;
        RECT 2698.425 2184.195 2698.595 2184.385 ;
        RECT 2702.565 2184.175 2702.735 2184.365 ;
        RECT 2703.945 2184.195 2704.115 2184.385 ;
        RECT 2707.635 2184.230 2707.795 2184.340 ;
        RECT 2708.085 2184.175 2708.255 2184.365 ;
        RECT 2709.005 2184.195 2709.175 2184.385 ;
        RECT 2713.605 2184.175 2713.775 2184.365 ;
        RECT 2714.525 2184.195 2714.695 2184.385 ;
        RECT 2719.125 2184.175 2719.295 2184.365 ;
        RECT 2720.045 2184.195 2720.215 2184.385 ;
        RECT 2720.960 2184.225 2721.080 2184.335 ;
        RECT 2721.885 2184.175 2722.055 2184.365 ;
        RECT 2725.565 2184.195 2725.735 2184.385 ;
        RECT 2727.405 2184.175 2727.575 2184.365 ;
        RECT 2731.085 2184.195 2731.255 2184.385 ;
        RECT 2733.845 2184.175 2734.015 2184.385 ;
        RECT 2695.525 2183.365 2696.895 2184.175 ;
        RECT 2696.905 2183.365 2702.415 2184.175 ;
        RECT 2702.425 2183.365 2707.935 2184.175 ;
        RECT 2707.945 2183.365 2713.455 2184.175 ;
        RECT 2713.465 2183.365 2718.975 2184.175 ;
        RECT 2718.985 2183.365 2720.815 2184.175 ;
        RECT 2721.745 2183.365 2727.255 2184.175 ;
        RECT 2727.265 2183.365 2732.775 2184.175 ;
        RECT 2732.785 2183.365 2734.155 2184.175 ;
        RECT 2695.525 2178.945 2696.895 2179.755 ;
        RECT 2696.905 2178.945 2700.575 2179.755 ;
        RECT 2701.505 2178.945 2702.855 2179.855 ;
        RECT 2702.885 2178.945 2708.395 2179.755 ;
        RECT 2708.865 2178.945 2714.375 2179.755 ;
        RECT 2714.385 2178.945 2719.895 2179.755 ;
        RECT 2719.905 2178.945 2725.415 2179.755 ;
        RECT 2725.425 2178.945 2730.935 2179.755 ;
        RECT 2730.945 2178.945 2732.775 2179.755 ;
        RECT 2732.785 2178.945 2734.155 2179.755 ;
        RECT 2695.665 2178.735 2695.835 2178.945 ;
        RECT 2697.045 2178.735 2697.215 2178.945 ;
        RECT 2698.425 2178.735 2698.595 2178.925 ;
        RECT 2700.735 2178.790 2700.895 2178.900 ;
        RECT 2701.650 2178.755 2701.820 2178.945 ;
        RECT 2703.025 2178.755 2703.195 2178.945 ;
        RECT 2704.865 2178.735 2705.035 2178.925 ;
        RECT 2705.325 2178.735 2705.495 2178.925 ;
        RECT 2709.005 2178.755 2709.175 2178.945 ;
        RECT 2710.845 2178.735 2711.015 2178.925 ;
        RECT 2714.525 2178.755 2714.695 2178.945 ;
        RECT 2716.365 2178.735 2716.535 2178.925 ;
        RECT 2720.045 2178.735 2720.215 2178.945 ;
        RECT 2721.885 2178.735 2722.055 2178.925 ;
        RECT 2725.565 2178.755 2725.735 2178.945 ;
        RECT 2727.405 2178.735 2727.575 2178.925 ;
        RECT 2731.085 2178.755 2731.255 2178.945 ;
        RECT 2733.845 2178.735 2734.015 2178.945 ;
        RECT 2695.525 2177.925 2696.895 2178.735 ;
        RECT 2696.905 2177.955 2698.275 2178.735 ;
        RECT 2698.285 2177.925 2701.955 2178.735 ;
        RECT 2701.965 2177.825 2705.175 2178.735 ;
        RECT 2705.185 2177.925 2710.695 2178.735 ;
        RECT 2710.705 2177.925 2716.215 2178.735 ;
        RECT 2716.225 2177.925 2719.895 2178.735 ;
        RECT 2719.905 2177.925 2721.275 2178.735 ;
        RECT 2721.745 2177.925 2727.255 2178.735 ;
        RECT 2727.265 2177.925 2732.775 2178.735 ;
        RECT 2732.785 2177.925 2734.155 2178.735 ;
        RECT 2695.525 2173.505 2696.895 2174.315 ;
        RECT 2696.905 2173.505 2702.415 2174.315 ;
        RECT 2702.425 2173.505 2707.935 2174.315 ;
        RECT 2708.865 2173.505 2714.375 2174.315 ;
        RECT 2714.385 2173.505 2719.895 2174.315 ;
        RECT 2719.905 2173.505 2725.415 2174.315 ;
        RECT 2725.425 2173.505 2732.775 2174.415 ;
        RECT 2732.785 2173.505 2734.155 2174.315 ;
        RECT 2695.665 2173.295 2695.835 2173.505 ;
        RECT 2697.045 2173.295 2697.215 2173.505 ;
        RECT 2698.425 2173.295 2698.595 2173.485 ;
        RECT 2702.565 2173.315 2702.735 2173.505 ;
        RECT 2703.945 2173.295 2704.115 2173.485 ;
        RECT 2708.080 2173.345 2708.200 2173.455 ;
        RECT 2709.005 2173.315 2709.175 2173.505 ;
        RECT 2709.465 2173.295 2709.635 2173.485 ;
        RECT 2714.525 2173.315 2714.695 2173.505 ;
        RECT 2714.985 2173.295 2715.155 2173.485 ;
        RECT 2720.045 2173.315 2720.215 2173.505 ;
        RECT 2720.515 2173.340 2720.675 2173.450 ;
        RECT 2721.885 2173.295 2722.055 2173.485 ;
        RECT 2725.990 2173.315 2726.160 2173.505 ;
        RECT 2727.405 2173.295 2727.575 2173.485 ;
        RECT 2733.845 2173.295 2734.015 2173.505 ;
        RECT 2695.525 2172.485 2696.895 2173.295 ;
        RECT 2696.905 2172.515 2698.275 2173.295 ;
        RECT 2698.285 2172.485 2703.795 2173.295 ;
        RECT 2703.805 2172.485 2709.315 2173.295 ;
        RECT 2709.325 2172.485 2714.835 2173.295 ;
        RECT 2714.845 2172.485 2720.355 2173.295 ;
        RECT 2721.745 2172.485 2727.255 2173.295 ;
        RECT 2727.265 2172.485 2732.775 2173.295 ;
        RECT 2732.785 2172.485 2734.155 2173.295 ;
        RECT 2695.525 2168.065 2696.895 2168.875 ;
        RECT 2696.905 2168.065 2702.415 2168.875 ;
        RECT 2702.425 2168.065 2707.935 2168.875 ;
        RECT 2708.865 2168.065 2714.375 2168.875 ;
        RECT 2714.385 2168.065 2719.895 2168.875 ;
        RECT 2719.905 2168.065 2725.415 2168.875 ;
        RECT 2725.425 2168.065 2730.935 2168.875 ;
        RECT 2730.945 2168.065 2732.775 2168.875 ;
        RECT 2732.785 2168.065 2734.155 2168.875 ;
        RECT 2695.665 2167.855 2695.835 2168.065 ;
        RECT 2697.045 2167.875 2697.215 2168.065 ;
        RECT 2699.345 2167.875 2699.515 2168.045 ;
        RECT 2699.345 2167.855 2699.475 2167.875 ;
        RECT 2699.805 2167.855 2699.975 2168.045 ;
        RECT 2702.565 2167.875 2702.735 2168.065 ;
        RECT 2705.325 2167.855 2705.495 2168.045 ;
        RECT 2708.080 2167.905 2708.200 2168.015 ;
        RECT 2709.005 2167.875 2709.175 2168.065 ;
        RECT 2710.845 2167.855 2711.015 2168.045 ;
        RECT 2714.525 2167.875 2714.695 2168.065 ;
        RECT 2716.365 2167.855 2716.535 2168.045 ;
        RECT 2720.045 2167.855 2720.215 2168.065 ;
        RECT 2721.885 2167.855 2722.055 2168.045 ;
        RECT 2725.565 2167.875 2725.735 2168.065 ;
        RECT 2727.405 2167.855 2727.575 2168.045 ;
        RECT 2731.085 2167.875 2731.255 2168.065 ;
        RECT 2733.845 2167.855 2734.015 2168.065 ;
        RECT 2695.525 2167.045 2696.895 2167.855 ;
        RECT 2697.625 2167.625 2699.475 2167.855 ;
        RECT 2697.140 2166.945 2699.475 2167.625 ;
        RECT 2699.665 2167.045 2705.175 2167.855 ;
        RECT 2705.185 2167.045 2710.695 2167.855 ;
        RECT 2710.705 2167.045 2716.215 2167.855 ;
        RECT 2716.225 2167.045 2719.895 2167.855 ;
        RECT 2719.905 2167.045 2721.275 2167.855 ;
        RECT 2721.745 2167.045 2727.255 2167.855 ;
        RECT 2727.265 2167.045 2732.775 2167.855 ;
        RECT 2732.785 2167.045 2734.155 2167.855 ;
        RECT 2695.525 2162.625 2696.895 2163.435 ;
        RECT 2696.905 2162.625 2698.275 2163.405 ;
        RECT 2698.285 2162.625 2703.795 2163.435 ;
        RECT 2703.805 2162.625 2707.475 2163.435 ;
        RECT 2708.865 2162.625 2714.375 2163.435 ;
        RECT 2714.385 2162.625 2719.895 2163.435 ;
        RECT 2719.905 2162.625 2725.415 2163.435 ;
        RECT 2725.425 2162.625 2730.935 2163.435 ;
        RECT 2730.945 2162.625 2732.775 2163.435 ;
        RECT 2732.785 2162.625 2734.155 2163.435 ;
        RECT 2695.665 2162.415 2695.835 2162.625 ;
        RECT 2697.045 2162.435 2697.215 2162.625 ;
        RECT 2698.425 2162.435 2698.595 2162.625 ;
        RECT 2700.450 2162.415 2700.620 2162.605 ;
        RECT 2702.575 2162.415 2702.745 2162.585 ;
        RECT 2703.945 2162.435 2704.115 2162.625 ;
        RECT 2704.405 2162.415 2704.575 2162.605 ;
        RECT 2704.865 2162.415 2705.035 2162.605 ;
        RECT 2707.635 2162.470 2707.795 2162.580 ;
        RECT 2709.005 2162.435 2709.175 2162.625 ;
        RECT 2710.385 2162.415 2710.555 2162.605 ;
        RECT 2714.525 2162.435 2714.695 2162.625 ;
        RECT 2715.905 2162.415 2716.075 2162.605 ;
        RECT 2720.045 2162.435 2720.215 2162.625 ;
        RECT 2721.885 2162.415 2722.055 2162.605 ;
        RECT 2725.565 2162.435 2725.735 2162.625 ;
        RECT 2727.405 2162.415 2727.575 2162.605 ;
        RECT 2731.085 2162.435 2731.255 2162.625 ;
        RECT 2733.845 2162.415 2734.015 2162.625 ;
        RECT 2364.485 2161.530 2365.085 2161.745 ;
        RECT 2381.705 2161.530 2382.305 2161.745 ;
        RECT 2398.925 2161.530 2399.525 2161.745 ;
        RECT 2416.145 2161.530 2416.745 2161.745 ;
        RECT 2433.365 2161.530 2433.965 2161.745 ;
        RECT 2695.525 2161.605 2696.895 2162.415 ;
        RECT 2697.135 2161.735 2701.035 2162.415 ;
        RECT 2364.485 2161.340 2365.380 2161.530 ;
        RECT 2367.510 2161.495 2367.680 2161.530 ;
        RECT 2366.605 2161.385 2367.680 2161.495 ;
        RECT 2367.395 2161.340 2367.680 2161.385 ;
        RECT 2369.820 2161.340 2369.990 2161.530 ;
        RECT 2371.200 2161.500 2371.370 2161.530 ;
        RECT 2371.200 2161.390 2371.770 2161.500 ;
        RECT 2371.200 2161.340 2371.485 2161.390 ;
        RECT 2364.485 2161.145 2366.445 2161.340 ;
        RECT 2365.095 2160.430 2366.445 2161.145 ;
        RECT 2367.395 2160.430 2371.485 2161.340 ;
        RECT 2381.705 2161.340 2382.600 2161.530 ;
        RECT 2384.730 2161.495 2384.900 2161.530 ;
        RECT 2383.825 2161.385 2384.900 2161.495 ;
        RECT 2384.615 2161.340 2384.900 2161.385 ;
        RECT 2387.040 2161.340 2387.210 2161.530 ;
        RECT 2388.420 2161.500 2388.590 2161.530 ;
        RECT 2388.420 2161.390 2388.990 2161.500 ;
        RECT 2388.420 2161.340 2388.705 2161.390 ;
        RECT 2381.705 2161.145 2383.665 2161.340 ;
        RECT 2382.315 2160.430 2383.665 2161.145 ;
        RECT 2384.615 2160.430 2388.705 2161.340 ;
        RECT 2398.925 2161.340 2399.820 2161.530 ;
        RECT 2401.950 2161.495 2402.120 2161.530 ;
        RECT 2401.045 2161.385 2402.120 2161.495 ;
        RECT 2401.835 2161.340 2402.120 2161.385 ;
        RECT 2404.260 2161.340 2404.430 2161.530 ;
        RECT 2405.640 2161.500 2405.810 2161.530 ;
        RECT 2405.640 2161.390 2406.210 2161.500 ;
        RECT 2405.640 2161.340 2405.925 2161.390 ;
        RECT 2398.925 2161.145 2400.885 2161.340 ;
        RECT 2399.535 2160.430 2400.885 2161.145 ;
        RECT 2401.835 2160.430 2405.925 2161.340 ;
        RECT 2416.145 2161.340 2417.040 2161.530 ;
        RECT 2419.170 2161.495 2419.340 2161.530 ;
        RECT 2418.265 2161.385 2419.340 2161.495 ;
        RECT 2419.055 2161.340 2419.340 2161.385 ;
        RECT 2421.480 2161.340 2421.650 2161.530 ;
        RECT 2422.860 2161.500 2423.030 2161.530 ;
        RECT 2422.860 2161.390 2423.430 2161.500 ;
        RECT 2422.860 2161.340 2423.145 2161.390 ;
        RECT 2416.145 2161.145 2418.105 2161.340 ;
        RECT 2416.755 2160.430 2418.105 2161.145 ;
        RECT 2419.055 2160.430 2423.145 2161.340 ;
        RECT 2433.365 2161.340 2434.260 2161.530 ;
        RECT 2436.390 2161.495 2436.560 2161.530 ;
        RECT 2435.485 2161.385 2436.560 2161.495 ;
        RECT 2436.275 2161.340 2436.560 2161.385 ;
        RECT 2438.700 2161.340 2438.870 2161.530 ;
        RECT 2440.080 2161.500 2440.250 2161.530 ;
        RECT 2700.105 2161.505 2701.035 2161.735 ;
        RECT 2701.045 2161.505 2704.695 2162.415 ;
        RECT 2704.725 2161.605 2710.235 2162.415 ;
        RECT 2710.245 2161.605 2715.755 2162.415 ;
        RECT 2715.765 2161.605 2721.275 2162.415 ;
        RECT 2721.745 2161.605 2727.255 2162.415 ;
        RECT 2727.265 2161.605 2732.775 2162.415 ;
        RECT 2732.785 2161.605 2734.155 2162.415 ;
        RECT 2440.080 2161.390 2440.650 2161.500 ;
        RECT 2440.080 2161.340 2440.365 2161.390 ;
        RECT 2433.365 2161.145 2435.325 2161.340 ;
        RECT 2433.975 2160.430 2435.325 2161.145 ;
        RECT 2436.275 2160.430 2440.365 2161.340 ;
        RECT 2695.525 2157.185 2696.895 2157.995 ;
        RECT 2696.905 2157.895 2697.835 2158.095 ;
        RECT 2699.165 2157.895 2700.115 2158.095 ;
        RECT 2696.905 2157.415 2700.115 2157.895 ;
        RECT 2697.050 2157.215 2700.115 2157.415 ;
        RECT 2364.625 2156.305 2371.925 2157.020 ;
        RECT 2381.845 2156.305 2389.145 2157.020 ;
        RECT 2399.065 2156.305 2406.365 2157.020 ;
        RECT 2416.285 2156.305 2423.585 2157.020 ;
        RECT 2433.505 2156.305 2440.805 2157.020 ;
        RECT 2695.665 2156.975 2695.835 2157.185 ;
        RECT 2697.050 2157.165 2697.220 2157.215 ;
        RECT 2699.180 2157.185 2700.115 2157.215 ;
        RECT 2700.125 2157.185 2705.635 2157.995 ;
        RECT 2705.645 2157.185 2708.395 2157.995 ;
        RECT 2708.865 2157.185 2714.375 2157.995 ;
        RECT 2714.385 2157.185 2719.895 2157.995 ;
        RECT 2719.905 2157.185 2725.415 2157.995 ;
        RECT 2725.425 2157.185 2730.935 2157.995 ;
        RECT 2730.945 2157.185 2732.775 2157.995 ;
        RECT 2732.785 2157.185 2734.155 2157.995 ;
        RECT 2883.065 2157.380 2883.235 2157.550 ;
        RECT 2697.045 2156.995 2697.220 2157.165 ;
        RECT 2697.045 2156.975 2697.215 2156.995 ;
        RECT 2698.425 2156.975 2698.595 2157.165 ;
        RECT 2700.265 2156.995 2700.435 2157.185 ;
        RECT 2703.945 2156.975 2704.115 2157.165 ;
        RECT 2705.785 2156.995 2705.955 2157.185 ;
        RECT 2709.005 2156.995 2709.175 2157.185 ;
        RECT 2709.465 2156.975 2709.635 2157.165 ;
        RECT 2714.525 2156.995 2714.695 2157.185 ;
        RECT 2714.985 2156.975 2715.155 2157.165 ;
        RECT 2720.045 2156.995 2720.215 2157.185 ;
        RECT 2720.515 2157.020 2720.675 2157.130 ;
        RECT 2721.885 2156.975 2722.055 2157.165 ;
        RECT 2725.565 2156.995 2725.735 2157.185 ;
        RECT 2727.405 2156.975 2727.575 2157.165 ;
        RECT 2731.085 2156.995 2731.255 2157.185 ;
        RECT 2733.845 2156.975 2734.015 2157.185 ;
        RECT 2364.485 2156.110 2371.925 2156.305 ;
        RECT 2381.705 2156.110 2389.145 2156.305 ;
        RECT 2398.925 2156.110 2406.365 2156.305 ;
        RECT 2416.145 2156.110 2423.585 2156.305 ;
        RECT 2433.365 2156.110 2440.805 2156.305 ;
        RECT 2695.525 2156.165 2696.895 2156.975 ;
        RECT 2696.905 2156.195 2698.275 2156.975 ;
        RECT 2698.285 2156.165 2703.795 2156.975 ;
        RECT 2703.805 2156.165 2709.315 2156.975 ;
        RECT 2709.325 2156.165 2714.835 2156.975 ;
        RECT 2714.845 2156.165 2720.355 2156.975 ;
        RECT 2721.745 2156.165 2727.255 2156.975 ;
        RECT 2727.265 2156.165 2732.775 2156.975 ;
        RECT 2732.785 2156.165 2734.155 2156.975 ;
        RECT 2364.485 2155.920 2365.845 2156.110 ;
        RECT 2367.050 2155.920 2367.690 2156.110 ;
        RECT 2371.655 2155.920 2371.825 2156.110 ;
        RECT 2381.705 2155.920 2383.065 2156.110 ;
        RECT 2384.270 2155.920 2384.910 2156.110 ;
        RECT 2388.875 2155.920 2389.045 2156.110 ;
        RECT 2398.925 2155.920 2400.285 2156.110 ;
        RECT 2401.490 2155.920 2402.130 2156.110 ;
        RECT 2406.095 2155.920 2406.265 2156.110 ;
        RECT 2416.145 2155.920 2417.505 2156.110 ;
        RECT 2418.710 2155.920 2419.350 2156.110 ;
        RECT 2423.315 2155.920 2423.485 2156.110 ;
        RECT 2433.365 2155.920 2434.725 2156.110 ;
        RECT 2435.930 2155.920 2436.570 2156.110 ;
        RECT 2440.535 2155.920 2440.705 2156.110 ;
        RECT 2364.485 2155.705 2365.085 2155.920 ;
        RECT 2381.705 2155.705 2382.305 2155.920 ;
        RECT 2398.925 2155.705 2399.525 2155.920 ;
        RECT 2416.145 2155.705 2416.745 2155.920 ;
        RECT 2433.365 2155.705 2433.965 2155.920 ;
        RECT 2695.525 2151.745 2696.895 2152.555 ;
        RECT 2696.905 2151.745 2698.275 2152.555 ;
        RECT 2698.285 2151.745 2701.955 2152.655 ;
        RECT 2701.965 2151.745 2707.475 2152.555 ;
        RECT 2708.865 2151.745 2714.375 2152.555 ;
        RECT 2714.385 2151.745 2719.895 2152.555 ;
        RECT 2719.905 2151.745 2725.415 2152.555 ;
        RECT 2725.425 2151.745 2730.935 2152.555 ;
        RECT 2730.945 2151.745 2732.775 2152.555 ;
        RECT 2732.785 2151.745 2734.155 2152.555 ;
        RECT 2695.665 2151.535 2695.835 2151.745 ;
        RECT 2697.045 2151.555 2697.215 2151.745 ;
        RECT 2695.525 2150.725 2696.895 2151.535 ;
        RECT 2697.965 2151.505 2698.135 2151.725 ;
        RECT 2701.640 2151.555 2701.810 2151.745 ;
        RECT 2702.105 2151.555 2702.275 2151.745 ;
        RECT 2703.485 2151.535 2703.655 2151.725 ;
        RECT 2703.945 2151.535 2704.115 2151.725 ;
        RECT 2707.635 2151.590 2707.795 2151.700 ;
        RECT 2709.005 2151.555 2709.175 2151.745 ;
        RECT 2709.465 2151.535 2709.635 2151.725 ;
        RECT 2714.525 2151.555 2714.695 2151.745 ;
        RECT 2714.985 2151.535 2715.155 2151.725 ;
        RECT 2720.045 2151.555 2720.215 2151.745 ;
        RECT 2720.515 2151.580 2720.675 2151.690 ;
        RECT 2721.885 2151.535 2722.055 2151.725 ;
        RECT 2725.565 2151.555 2725.735 2151.745 ;
        RECT 2727.405 2151.535 2727.575 2151.725 ;
        RECT 2731.085 2151.555 2731.255 2151.745 ;
        RECT 2733.845 2151.535 2734.015 2151.745 ;
        RECT 2700.090 2151.505 2701.035 2151.535 ;
        RECT 2697.965 2151.305 2701.035 2151.505 ;
        RECT 2697.825 2150.825 2701.035 2151.305 ;
        RECT 2697.825 2150.625 2698.755 2150.825 ;
        RECT 2700.090 2150.625 2701.035 2150.825 ;
        RECT 2701.275 2151.305 2703.655 2151.535 ;
        RECT 2701.275 2150.625 2703.665 2151.305 ;
        RECT 2703.805 2150.725 2709.315 2151.535 ;
        RECT 2709.325 2150.725 2714.835 2151.535 ;
        RECT 2714.845 2150.725 2720.355 2151.535 ;
        RECT 2721.745 2150.725 2727.255 2151.535 ;
        RECT 2727.265 2150.725 2732.775 2151.535 ;
        RECT 2732.785 2150.725 2734.155 2151.535 ;
        RECT 2695.525 2146.305 2696.895 2147.115 ;
        RECT 2696.905 2146.305 2698.275 2147.085 ;
        RECT 2698.745 2146.305 2700.095 2147.215 ;
        RECT 2700.125 2146.305 2705.635 2147.115 ;
        RECT 2705.645 2146.305 2708.395 2147.115 ;
        RECT 2708.865 2146.305 2714.375 2147.115 ;
        RECT 2714.385 2146.305 2719.895 2147.115 ;
        RECT 2719.905 2146.305 2725.415 2147.115 ;
        RECT 2725.425 2146.305 2730.935 2147.115 ;
        RECT 2730.945 2146.305 2732.775 2147.115 ;
        RECT 2732.785 2146.305 2734.155 2147.115 ;
        RECT 2695.665 2146.095 2695.835 2146.305 ;
        RECT 2697.045 2146.115 2697.215 2146.305 ;
        RECT 2698.420 2146.145 2698.540 2146.255 ;
        RECT 2699.810 2146.115 2699.980 2146.305 ;
        RECT 2700.265 2146.115 2700.435 2146.305 ;
        RECT 2700.450 2146.095 2700.620 2146.285 ;
        RECT 2701.185 2146.095 2701.355 2146.285 ;
        RECT 2705.785 2146.115 2705.955 2146.305 ;
        RECT 2706.705 2146.095 2706.875 2146.285 ;
        RECT 2709.005 2146.115 2709.175 2146.305 ;
        RECT 2712.225 2146.095 2712.395 2146.285 ;
        RECT 2714.525 2146.115 2714.695 2146.305 ;
        RECT 2717.745 2146.095 2717.915 2146.285 ;
        RECT 2720.045 2146.115 2720.215 2146.305 ;
        RECT 2721.885 2146.095 2722.055 2146.285 ;
        RECT 2725.565 2146.115 2725.735 2146.305 ;
        RECT 2727.405 2146.095 2727.575 2146.285 ;
        RECT 2731.085 2146.115 2731.255 2146.305 ;
        RECT 2733.845 2146.095 2734.015 2146.305 ;
        RECT 2695.525 2145.285 2696.895 2146.095 ;
        RECT 2697.135 2145.415 2701.035 2146.095 ;
        RECT 2700.105 2145.185 2701.035 2145.415 ;
        RECT 2701.045 2145.285 2706.555 2146.095 ;
        RECT 2706.565 2145.285 2712.075 2146.095 ;
        RECT 2712.085 2145.285 2717.595 2146.095 ;
        RECT 2717.605 2145.285 2721.275 2146.095 ;
        RECT 2721.745 2145.285 2727.255 2146.095 ;
        RECT 2727.265 2145.285 2732.775 2146.095 ;
        RECT 2732.785 2145.285 2734.155 2146.095 ;
        RECT 2695.525 2140.865 2696.895 2141.675 ;
        RECT 2696.905 2140.865 2698.275 2141.645 ;
        RECT 2698.285 2140.865 2703.795 2141.675 ;
        RECT 2703.805 2140.865 2707.475 2141.675 ;
        RECT 2708.865 2140.865 2714.375 2141.675 ;
        RECT 2714.385 2140.865 2719.895 2141.675 ;
        RECT 2719.905 2140.865 2725.415 2141.675 ;
        RECT 2725.425 2140.865 2730.935 2141.675 ;
        RECT 2730.945 2140.865 2732.775 2141.675 ;
        RECT 2732.785 2140.865 2734.155 2141.675 ;
        RECT 2695.665 2140.655 2695.835 2140.865 ;
        RECT 2697.045 2140.655 2697.215 2140.865 ;
        RECT 2698.425 2140.675 2698.595 2140.865 ;
        RECT 2702.565 2140.655 2702.735 2140.845 ;
        RECT 2703.945 2140.675 2704.115 2140.865 ;
        RECT 2707.635 2140.710 2707.795 2140.820 ;
        RECT 2708.085 2140.655 2708.255 2140.845 ;
        RECT 2709.005 2140.675 2709.175 2140.865 ;
        RECT 2713.605 2140.655 2713.775 2140.845 ;
        RECT 2714.525 2140.675 2714.695 2140.865 ;
        RECT 2719.125 2140.655 2719.295 2140.845 ;
        RECT 2720.045 2140.675 2720.215 2140.865 ;
        RECT 2720.960 2140.705 2721.080 2140.815 ;
        RECT 2721.885 2140.655 2722.055 2140.845 ;
        RECT 2725.565 2140.675 2725.735 2140.865 ;
        RECT 2727.405 2140.655 2727.575 2140.845 ;
        RECT 2731.085 2140.675 2731.255 2140.865 ;
        RECT 2733.845 2140.655 2734.015 2140.865 ;
        RECT 2695.525 2139.845 2696.895 2140.655 ;
        RECT 2696.905 2139.845 2702.415 2140.655 ;
        RECT 2702.425 2139.845 2707.935 2140.655 ;
        RECT 2707.945 2139.845 2713.455 2140.655 ;
        RECT 2713.465 2139.845 2718.975 2140.655 ;
        RECT 2718.985 2139.845 2720.815 2140.655 ;
        RECT 2721.745 2139.845 2727.255 2140.655 ;
        RECT 2727.265 2139.845 2732.775 2140.655 ;
        RECT 2732.785 2139.845 2734.155 2140.655 ;
        RECT 2695.525 2135.425 2696.895 2136.235 ;
        RECT 2696.905 2135.425 2698.275 2136.205 ;
        RECT 2698.285 2135.425 2703.795 2136.235 ;
        RECT 2703.805 2135.425 2707.475 2136.235 ;
        RECT 2708.865 2135.425 2714.375 2136.235 ;
        RECT 2714.385 2135.425 2719.895 2136.235 ;
        RECT 2719.905 2135.425 2725.415 2136.235 ;
        RECT 2725.425 2135.425 2730.935 2136.235 ;
        RECT 2730.945 2135.425 2732.775 2136.235 ;
        RECT 2732.785 2135.425 2734.155 2136.235 ;
        RECT 2695.665 2135.215 2695.835 2135.425 ;
        RECT 2697.045 2135.215 2697.215 2135.425 ;
        RECT 2698.425 2135.235 2698.595 2135.425 ;
        RECT 2702.565 2135.215 2702.735 2135.405 ;
        RECT 2703.945 2135.235 2704.115 2135.425 ;
        RECT 2707.635 2135.270 2707.795 2135.380 ;
        RECT 2708.085 2135.215 2708.255 2135.405 ;
        RECT 2709.005 2135.235 2709.175 2135.425 ;
        RECT 2713.605 2135.215 2713.775 2135.405 ;
        RECT 2714.525 2135.235 2714.695 2135.425 ;
        RECT 2719.125 2135.215 2719.295 2135.405 ;
        RECT 2720.045 2135.235 2720.215 2135.425 ;
        RECT 2720.960 2135.265 2721.080 2135.375 ;
        RECT 2721.885 2135.215 2722.055 2135.405 ;
        RECT 2725.565 2135.235 2725.735 2135.425 ;
        RECT 2727.405 2135.215 2727.575 2135.405 ;
        RECT 2731.085 2135.235 2731.255 2135.425 ;
        RECT 2733.845 2135.215 2734.015 2135.425 ;
        RECT 2695.525 2134.405 2696.895 2135.215 ;
        RECT 2696.905 2134.405 2702.415 2135.215 ;
        RECT 2702.425 2134.405 2707.935 2135.215 ;
        RECT 2707.945 2134.405 2713.455 2135.215 ;
        RECT 2713.465 2134.405 2718.975 2135.215 ;
        RECT 2718.985 2134.405 2720.815 2135.215 ;
        RECT 2721.745 2134.405 2727.255 2135.215 ;
        RECT 2727.265 2134.405 2732.775 2135.215 ;
        RECT 2732.785 2134.405 2734.155 2135.215 ;
        RECT 2522.700 2133.870 2522.870 2134.040 ;
        RECT 2695.525 2129.985 2696.895 2130.795 ;
        RECT 2696.905 2129.985 2698.275 2130.765 ;
        RECT 2698.285 2129.985 2699.655 2130.765 ;
        RECT 2699.665 2129.985 2705.175 2130.795 ;
        RECT 2705.185 2129.985 2707.935 2130.795 ;
        RECT 2708.865 2129.985 2714.375 2130.795 ;
        RECT 2714.385 2129.985 2719.895 2130.795 ;
        RECT 2719.905 2129.985 2721.275 2130.795 ;
        RECT 2721.745 2129.985 2727.255 2130.795 ;
        RECT 2727.265 2129.985 2732.775 2130.795 ;
        RECT 2732.785 2129.985 2734.155 2130.795 ;
        RECT 2695.665 2129.795 2695.835 2129.985 ;
        RECT 2697.045 2129.795 2697.215 2129.985 ;
        RECT 2698.425 2129.795 2698.595 2129.985 ;
        RECT 2699.805 2129.795 2699.975 2129.985 ;
        RECT 2705.325 2129.795 2705.495 2129.985 ;
        RECT 2708.080 2129.825 2708.200 2129.935 ;
        RECT 2709.005 2129.795 2709.175 2129.985 ;
        RECT 2714.525 2129.795 2714.695 2129.985 ;
        RECT 2720.045 2129.795 2720.215 2129.985 ;
        RECT 2721.885 2129.795 2722.055 2129.985 ;
        RECT 2727.405 2129.795 2727.575 2129.985 ;
        RECT 2733.845 2129.795 2734.015 2129.985 ;
        RECT 2522.700 2126.340 2522.870 2126.510 ;
        RECT 2522.700 2120.360 2522.870 2120.530 ;
        RECT 2522.700 2114.415 2522.870 2114.585 ;
        RECT 2522.700 2108.770 2522.870 2108.940 ;
        RECT 2522.700 2102.765 2522.870 2102.935 ;
        RECT 2361.700 2050.735 2361.870 2050.875 ;
        RECT 2361.680 2050.715 2361.870 2050.735 ;
        RECT 2364.140 2050.715 2364.310 2050.875 ;
        RECT 2366.580 2050.715 2366.750 2050.875 ;
        RECT 2369.020 2050.735 2369.190 2050.875 ;
        RECT 2378.025 2050.735 2378.195 2050.875 ;
        RECT 2369.020 2050.715 2369.210 2050.735 ;
        RECT 2361.680 2050.705 2361.850 2050.715 ;
        RECT 2369.040 2050.705 2369.210 2050.715 ;
        RECT 2378.005 2050.715 2378.195 2050.735 ;
        RECT 2380.465 2050.715 2380.635 2050.875 ;
        RECT 2382.905 2050.715 2383.075 2050.875 ;
        RECT 2385.345 2050.735 2385.515 2050.875 ;
        RECT 2394.350 2050.735 2394.520 2050.875 ;
        RECT 2385.345 2050.715 2385.535 2050.735 ;
        RECT 2378.005 2050.705 2378.175 2050.715 ;
        RECT 2385.365 2050.705 2385.535 2050.715 ;
        RECT 2394.330 2050.715 2394.520 2050.735 ;
        RECT 2396.790 2050.715 2396.960 2050.875 ;
        RECT 2399.230 2050.715 2399.400 2050.875 ;
        RECT 2401.670 2050.735 2401.840 2050.875 ;
        RECT 2410.675 2050.735 2410.845 2050.875 ;
        RECT 2401.670 2050.715 2401.860 2050.735 ;
        RECT 2394.330 2050.705 2394.500 2050.715 ;
        RECT 2401.690 2050.705 2401.860 2050.715 ;
        RECT 2410.655 2050.715 2410.845 2050.735 ;
        RECT 2413.115 2050.715 2413.285 2050.875 ;
        RECT 2415.555 2050.715 2415.725 2050.875 ;
        RECT 2417.995 2050.735 2418.165 2050.875 ;
        RECT 2427.000 2050.735 2427.170 2050.875 ;
        RECT 2417.995 2050.715 2418.185 2050.735 ;
        RECT 2410.655 2050.705 2410.825 2050.715 ;
        RECT 2418.015 2050.705 2418.185 2050.715 ;
        RECT 2426.980 2050.715 2427.170 2050.735 ;
        RECT 2429.440 2050.715 2429.610 2050.875 ;
        RECT 2431.880 2050.715 2432.050 2050.875 ;
        RECT 2434.320 2050.735 2434.490 2050.875 ;
        RECT 2434.320 2050.715 2434.510 2050.735 ;
        RECT 2426.980 2050.705 2427.150 2050.715 ;
        RECT 2434.340 2050.705 2434.510 2050.715 ;
        RECT 2695.665 2036.815 2695.835 2037.005 ;
        RECT 2697.045 2036.815 2697.215 2037.005 ;
        RECT 2699.805 2036.815 2699.975 2037.005 ;
        RECT 2701.185 2036.815 2701.355 2037.005 ;
        RECT 2701.645 2036.815 2701.815 2037.005 ;
        RECT 2707.165 2036.815 2707.335 2037.005 ;
        RECT 2709.005 2036.815 2709.175 2037.005 ;
        RECT 2710.845 2036.815 2711.015 2037.005 ;
        RECT 2716.365 2036.815 2716.535 2037.005 ;
        RECT 2720.045 2036.815 2720.215 2037.005 ;
        RECT 2723.265 2036.815 2723.435 2037.005 ;
        RECT 2723.725 2036.815 2723.895 2037.005 ;
        RECT 2729.245 2036.815 2729.415 2037.005 ;
        RECT 2731.080 2036.865 2731.200 2036.975 ;
        RECT 2732.455 2036.815 2732.625 2037.005 ;
        RECT 2733.845 2036.815 2734.015 2037.005 ;
        RECT 2695.525 2036.005 2696.895 2036.815 ;
        RECT 2696.905 2036.135 2698.735 2036.815 ;
        RECT 2698.745 2036.035 2700.115 2036.815 ;
        RECT 2700.125 2036.035 2701.495 2036.815 ;
        RECT 2701.505 2036.005 2707.015 2036.815 ;
        RECT 2707.025 2036.005 2708.395 2036.815 ;
        RECT 2708.865 2036.135 2710.695 2036.815 ;
        RECT 2709.350 2035.905 2710.695 2036.135 ;
        RECT 2710.705 2036.005 2716.215 2036.815 ;
        RECT 2716.225 2036.005 2719.895 2036.815 ;
        RECT 2719.905 2036.005 2721.275 2036.815 ;
        RECT 2721.745 2036.135 2723.575 2036.815 ;
        RECT 2723.585 2036.005 2729.095 2036.815 ;
        RECT 2729.105 2036.005 2730.935 2036.815 ;
        RECT 2731.405 2036.035 2732.775 2036.815 ;
        RECT 2732.785 2036.005 2734.155 2036.815 ;
        RECT 2695.525 2031.585 2696.895 2032.395 ;
        RECT 2696.905 2031.585 2698.275 2032.365 ;
        RECT 2698.285 2031.585 2703.795 2032.395 ;
        RECT 2703.805 2031.585 2707.475 2032.395 ;
        RECT 2708.865 2031.585 2714.375 2032.395 ;
        RECT 2714.385 2031.585 2719.895 2032.395 ;
        RECT 2719.905 2031.585 2725.415 2032.395 ;
        RECT 2725.425 2031.585 2730.935 2032.395 ;
        RECT 2730.945 2031.585 2732.775 2032.395 ;
        RECT 2732.785 2031.585 2734.155 2032.395 ;
        RECT 2695.665 2031.375 2695.835 2031.585 ;
        RECT 2697.045 2031.375 2697.215 2031.585 ;
        RECT 2698.425 2031.395 2698.595 2031.585 ;
        RECT 2702.565 2031.375 2702.735 2031.565 ;
        RECT 2703.945 2031.395 2704.115 2031.585 ;
        RECT 2707.635 2031.430 2707.795 2031.540 ;
        RECT 2708.085 2031.375 2708.255 2031.565 ;
        RECT 2709.005 2031.395 2709.175 2031.585 ;
        RECT 2713.605 2031.375 2713.775 2031.565 ;
        RECT 2714.525 2031.395 2714.695 2031.585 ;
        RECT 2719.125 2031.375 2719.295 2031.565 ;
        RECT 2720.045 2031.395 2720.215 2031.585 ;
        RECT 2720.960 2031.425 2721.080 2031.535 ;
        RECT 2721.885 2031.375 2722.055 2031.565 ;
        RECT 2725.565 2031.395 2725.735 2031.585 ;
        RECT 2727.405 2031.375 2727.575 2031.565 ;
        RECT 2731.085 2031.395 2731.255 2031.585 ;
        RECT 2733.845 2031.375 2734.015 2031.585 ;
        RECT 2695.525 2030.565 2696.895 2031.375 ;
        RECT 2696.905 2030.565 2702.415 2031.375 ;
        RECT 2702.425 2030.565 2707.935 2031.375 ;
        RECT 2707.945 2030.565 2713.455 2031.375 ;
        RECT 2713.465 2030.565 2718.975 2031.375 ;
        RECT 2718.985 2030.565 2720.815 2031.375 ;
        RECT 2721.745 2030.565 2727.255 2031.375 ;
        RECT 2727.265 2030.565 2732.775 2031.375 ;
        RECT 2732.785 2030.565 2734.155 2031.375 ;
        RECT 2695.525 2026.145 2696.895 2026.955 ;
        RECT 2696.905 2026.145 2702.415 2026.955 ;
        RECT 2702.425 2026.145 2707.935 2026.955 ;
        RECT 2708.865 2026.145 2714.375 2026.955 ;
        RECT 2714.385 2026.145 2719.895 2026.955 ;
        RECT 2719.905 2026.145 2725.415 2026.955 ;
        RECT 2725.425 2026.145 2730.935 2026.955 ;
        RECT 2730.945 2026.145 2732.775 2026.955 ;
        RECT 2732.785 2026.145 2734.155 2026.955 ;
        RECT 2695.665 2025.935 2695.835 2026.145 ;
        RECT 2697.045 2025.935 2697.215 2026.145 ;
        RECT 2698.425 2025.935 2698.595 2026.125 ;
        RECT 2702.565 2025.955 2702.735 2026.145 ;
        RECT 2703.945 2025.935 2704.115 2026.125 ;
        RECT 2708.080 2025.985 2708.200 2026.095 ;
        RECT 2709.005 2025.955 2709.175 2026.145 ;
        RECT 2709.465 2025.935 2709.635 2026.125 ;
        RECT 2714.525 2025.955 2714.695 2026.145 ;
        RECT 2714.985 2025.935 2715.155 2026.125 ;
        RECT 2720.045 2025.955 2720.215 2026.145 ;
        RECT 2720.515 2025.980 2720.675 2026.090 ;
        RECT 2721.885 2025.935 2722.055 2026.125 ;
        RECT 2725.565 2025.955 2725.735 2026.145 ;
        RECT 2727.405 2025.935 2727.575 2026.125 ;
        RECT 2731.085 2025.955 2731.255 2026.145 ;
        RECT 2733.845 2025.935 2734.015 2026.145 ;
        RECT 2695.525 2025.125 2696.895 2025.935 ;
        RECT 2696.905 2025.155 2698.275 2025.935 ;
        RECT 2698.285 2025.125 2703.795 2025.935 ;
        RECT 2703.805 2025.125 2709.315 2025.935 ;
        RECT 2709.325 2025.125 2714.835 2025.935 ;
        RECT 2714.845 2025.125 2720.355 2025.935 ;
        RECT 2721.745 2025.125 2727.255 2025.935 ;
        RECT 2727.265 2025.125 2732.775 2025.935 ;
        RECT 2732.785 2025.125 2734.155 2025.935 ;
        RECT 2695.525 2020.705 2696.895 2021.515 ;
        RECT 2696.905 2020.705 2702.415 2021.515 ;
        RECT 2702.425 2020.705 2707.935 2021.515 ;
        RECT 2708.865 2020.705 2714.375 2021.515 ;
        RECT 2714.385 2020.705 2719.895 2021.515 ;
        RECT 2719.905 2020.705 2725.415 2021.515 ;
        RECT 2725.425 2020.705 2730.935 2021.515 ;
        RECT 2730.945 2020.705 2732.775 2021.515 ;
        RECT 2732.785 2020.705 2734.155 2021.515 ;
        RECT 2695.665 2020.495 2695.835 2020.705 ;
        RECT 2697.045 2020.495 2697.215 2020.705 ;
        RECT 2702.565 2020.515 2702.735 2020.705 ;
        RECT 2706.705 2020.495 2706.875 2020.685 ;
        RECT 2708.080 2020.545 2708.200 2020.655 ;
        RECT 2709.005 2020.515 2709.175 2020.705 ;
        RECT 2712.225 2020.495 2712.395 2020.685 ;
        RECT 2714.525 2020.515 2714.695 2020.705 ;
        RECT 2717.745 2020.495 2717.915 2020.685 ;
        RECT 2720.045 2020.515 2720.215 2020.705 ;
        RECT 2721.885 2020.495 2722.055 2020.685 ;
        RECT 2725.565 2020.515 2725.735 2020.705 ;
        RECT 2727.405 2020.495 2727.575 2020.685 ;
        RECT 2731.085 2020.515 2731.255 2020.705 ;
        RECT 2733.845 2020.495 2734.015 2020.705 ;
        RECT 2695.525 2019.685 2696.895 2020.495 ;
        RECT 2696.905 2020.325 2698.665 2020.495 ;
        RECT 2696.905 2020.280 2699.160 2020.325 ;
        RECT 2696.905 2020.245 2700.100 2020.280 ;
        RECT 2701.460 2020.245 2706.555 2020.495 ;
        RECT 2696.905 2019.815 2706.555 2020.245 ;
        RECT 2698.230 2019.645 2701.460 2019.815 ;
        RECT 2699.170 2019.600 2701.460 2019.645 ;
        RECT 2700.110 2019.565 2701.460 2019.600 ;
        RECT 2704.535 2019.585 2706.555 2019.815 ;
        RECT 2706.565 2019.685 2712.075 2020.495 ;
        RECT 2712.085 2019.685 2717.595 2020.495 ;
        RECT 2717.605 2019.685 2721.275 2020.495 ;
        RECT 2721.745 2019.685 2727.255 2020.495 ;
        RECT 2727.265 2019.685 2732.775 2020.495 ;
        RECT 2732.785 2019.685 2734.155 2020.495 ;
        RECT 2704.535 2019.565 2705.455 2019.585 ;
        RECT 2695.525 2015.265 2696.895 2016.075 ;
        RECT 2696.905 2015.265 2698.275 2016.045 ;
        RECT 2698.285 2015.265 2703.795 2016.075 ;
        RECT 2703.805 2015.265 2707.475 2016.075 ;
        RECT 2708.865 2015.265 2714.375 2016.075 ;
        RECT 2714.385 2015.265 2719.895 2016.075 ;
        RECT 2719.905 2015.265 2725.415 2016.075 ;
        RECT 2725.425 2015.265 2730.935 2016.075 ;
        RECT 2730.945 2015.265 2732.775 2016.075 ;
        RECT 2732.785 2015.265 2734.155 2016.075 ;
        RECT 2695.665 2015.055 2695.835 2015.265 ;
        RECT 2697.045 2015.055 2697.215 2015.265 ;
        RECT 2698.425 2015.075 2698.595 2015.265 ;
        RECT 2703.945 2015.075 2704.115 2015.265 ;
        RECT 2706.705 2015.055 2706.875 2015.245 ;
        RECT 2707.635 2015.110 2707.795 2015.220 ;
        RECT 2709.005 2015.075 2709.175 2015.265 ;
        RECT 2712.225 2015.055 2712.395 2015.245 ;
        RECT 2714.525 2015.075 2714.695 2015.265 ;
        RECT 2717.745 2015.055 2717.915 2015.245 ;
        RECT 2720.045 2015.075 2720.215 2015.265 ;
        RECT 2721.885 2015.055 2722.055 2015.245 ;
        RECT 2725.565 2015.075 2725.735 2015.265 ;
        RECT 2727.405 2015.055 2727.575 2015.245 ;
        RECT 2731.085 2015.075 2731.255 2015.265 ;
        RECT 2733.845 2015.055 2734.015 2015.265 ;
        RECT 2695.525 2014.245 2696.895 2015.055 ;
        RECT 2696.905 2014.885 2698.665 2015.055 ;
        RECT 2696.905 2014.840 2699.160 2014.885 ;
        RECT 2696.905 2014.805 2700.100 2014.840 ;
        RECT 2701.460 2014.805 2706.555 2015.055 ;
        RECT 2696.905 2014.375 2706.555 2014.805 ;
        RECT 2698.230 2014.205 2701.460 2014.375 ;
        RECT 2699.170 2014.160 2701.460 2014.205 ;
        RECT 2700.110 2014.125 2701.460 2014.160 ;
        RECT 2704.535 2014.145 2706.555 2014.375 ;
        RECT 2706.565 2014.245 2712.075 2015.055 ;
        RECT 2712.085 2014.245 2717.595 2015.055 ;
        RECT 2717.605 2014.245 2721.275 2015.055 ;
        RECT 2721.745 2014.245 2727.255 2015.055 ;
        RECT 2727.265 2014.245 2732.775 2015.055 ;
        RECT 2732.785 2014.245 2734.155 2015.055 ;
        RECT 2704.535 2014.125 2705.455 2014.145 ;
        RECT 2695.525 2009.825 2696.895 2010.635 ;
        RECT 2696.905 2009.825 2698.275 2010.605 ;
        RECT 2698.285 2009.825 2701.035 2010.635 ;
        RECT 2701.505 2010.505 2702.435 2010.735 ;
        RECT 2701.505 2009.825 2705.405 2010.505 ;
        RECT 2705.645 2009.825 2708.395 2010.635 ;
        RECT 2708.865 2009.825 2714.375 2010.635 ;
        RECT 2714.385 2009.825 2719.895 2010.635 ;
        RECT 2719.905 2009.825 2725.415 2010.635 ;
        RECT 2725.425 2009.825 2730.935 2010.635 ;
        RECT 2730.945 2009.825 2732.775 2010.635 ;
        RECT 2732.785 2009.825 2734.155 2010.635 ;
        RECT 2695.665 2009.615 2695.835 2009.825 ;
        RECT 2697.045 2009.615 2697.215 2009.825 ;
        RECT 2698.425 2009.635 2698.595 2009.825 ;
        RECT 2701.180 2009.665 2701.300 2009.775 ;
        RECT 2701.920 2009.635 2702.090 2009.825 ;
        RECT 2702.565 2009.615 2702.735 2009.805 ;
        RECT 2705.785 2009.635 2705.955 2009.825 ;
        RECT 2708.085 2009.615 2708.255 2009.805 ;
        RECT 2709.005 2009.635 2709.175 2009.825 ;
        RECT 2713.605 2009.615 2713.775 2009.805 ;
        RECT 2714.525 2009.635 2714.695 2009.825 ;
        RECT 2719.125 2009.615 2719.295 2009.805 ;
        RECT 2720.045 2009.635 2720.215 2009.825 ;
        RECT 2720.960 2009.665 2721.080 2009.775 ;
        RECT 2721.885 2009.615 2722.055 2009.805 ;
        RECT 2725.565 2009.635 2725.735 2009.825 ;
        RECT 2727.405 2009.615 2727.575 2009.805 ;
        RECT 2731.085 2009.635 2731.255 2009.825 ;
        RECT 2733.845 2009.615 2734.015 2009.825 ;
        RECT 2695.525 2008.805 2696.895 2009.615 ;
        RECT 2696.905 2008.805 2702.415 2009.615 ;
        RECT 2702.425 2008.805 2707.935 2009.615 ;
        RECT 2707.945 2008.805 2713.455 2009.615 ;
        RECT 2713.465 2008.805 2718.975 2009.615 ;
        RECT 2718.985 2008.805 2720.815 2009.615 ;
        RECT 2721.745 2008.805 2727.255 2009.615 ;
        RECT 2727.265 2008.805 2732.775 2009.615 ;
        RECT 2732.785 2008.805 2734.155 2009.615 ;
        RECT 2695.525 2004.385 2696.895 2005.195 ;
        RECT 2696.905 2004.385 2698.275 2005.165 ;
        RECT 2698.285 2004.385 2703.795 2005.195 ;
        RECT 2703.805 2004.385 2707.475 2005.195 ;
        RECT 2708.865 2004.385 2714.375 2005.195 ;
        RECT 2714.385 2004.385 2719.895 2005.195 ;
        RECT 2719.905 2004.385 2725.415 2005.195 ;
        RECT 2725.425 2004.385 2730.935 2005.195 ;
        RECT 2730.945 2004.385 2732.775 2005.195 ;
        RECT 2732.785 2004.385 2734.155 2005.195 ;
        RECT 2695.665 2004.175 2695.835 2004.385 ;
        RECT 2697.045 2004.175 2697.215 2004.385 ;
        RECT 2698.425 2004.195 2698.595 2004.385 ;
        RECT 2702.565 2004.175 2702.735 2004.365 ;
        RECT 2703.945 2004.195 2704.115 2004.385 ;
        RECT 2707.635 2004.230 2707.795 2004.340 ;
        RECT 2708.085 2004.175 2708.255 2004.365 ;
        RECT 2709.005 2004.195 2709.175 2004.385 ;
        RECT 2713.605 2004.175 2713.775 2004.365 ;
        RECT 2714.525 2004.195 2714.695 2004.385 ;
        RECT 2719.125 2004.175 2719.295 2004.365 ;
        RECT 2720.045 2004.195 2720.215 2004.385 ;
        RECT 2720.960 2004.225 2721.080 2004.335 ;
        RECT 2721.885 2004.175 2722.055 2004.365 ;
        RECT 2725.565 2004.195 2725.735 2004.385 ;
        RECT 2727.405 2004.175 2727.575 2004.365 ;
        RECT 2731.085 2004.195 2731.255 2004.385 ;
        RECT 2733.845 2004.175 2734.015 2004.385 ;
        RECT 2695.525 2003.365 2696.895 2004.175 ;
        RECT 2696.905 2003.365 2702.415 2004.175 ;
        RECT 2702.425 2003.365 2707.935 2004.175 ;
        RECT 2707.945 2003.365 2713.455 2004.175 ;
        RECT 2713.465 2003.365 2718.975 2004.175 ;
        RECT 2718.985 2003.365 2720.815 2004.175 ;
        RECT 2721.745 2003.365 2727.255 2004.175 ;
        RECT 2727.265 2003.365 2732.775 2004.175 ;
        RECT 2732.785 2003.365 2734.155 2004.175 ;
        RECT 2695.525 1998.945 2696.895 1999.755 ;
        RECT 2696.905 1998.945 2700.575 1999.755 ;
        RECT 2701.505 1998.945 2702.855 1999.855 ;
        RECT 2702.885 1998.945 2708.395 1999.755 ;
        RECT 2708.865 1998.945 2714.375 1999.755 ;
        RECT 2714.385 1998.945 2719.895 1999.755 ;
        RECT 2719.905 1998.945 2725.415 1999.755 ;
        RECT 2725.425 1998.945 2730.935 1999.755 ;
        RECT 2730.945 1998.945 2732.775 1999.755 ;
        RECT 2732.785 1998.945 2734.155 1999.755 ;
        RECT 2695.665 1998.735 2695.835 1998.945 ;
        RECT 2697.045 1998.735 2697.215 1998.945 ;
        RECT 2698.425 1998.735 2698.595 1998.925 ;
        RECT 2700.735 1998.790 2700.895 1998.900 ;
        RECT 2701.650 1998.755 2701.820 1998.945 ;
        RECT 2703.025 1998.755 2703.195 1998.945 ;
        RECT 2704.865 1998.735 2705.035 1998.925 ;
        RECT 2705.325 1998.735 2705.495 1998.925 ;
        RECT 2709.005 1998.755 2709.175 1998.945 ;
        RECT 2710.845 1998.735 2711.015 1998.925 ;
        RECT 2714.525 1998.755 2714.695 1998.945 ;
        RECT 2716.365 1998.735 2716.535 1998.925 ;
        RECT 2720.045 1998.735 2720.215 1998.945 ;
        RECT 2721.885 1998.735 2722.055 1998.925 ;
        RECT 2725.565 1998.755 2725.735 1998.945 ;
        RECT 2727.405 1998.735 2727.575 1998.925 ;
        RECT 2731.085 1998.755 2731.255 1998.945 ;
        RECT 2733.845 1998.735 2734.015 1998.945 ;
        RECT 2695.525 1997.925 2696.895 1998.735 ;
        RECT 2696.905 1997.955 2698.275 1998.735 ;
        RECT 2698.285 1997.925 2701.955 1998.735 ;
        RECT 2701.965 1997.825 2705.175 1998.735 ;
        RECT 2705.185 1997.925 2710.695 1998.735 ;
        RECT 2710.705 1997.925 2716.215 1998.735 ;
        RECT 2716.225 1997.925 2719.895 1998.735 ;
        RECT 2719.905 1997.925 2721.275 1998.735 ;
        RECT 2721.745 1997.925 2727.255 1998.735 ;
        RECT 2727.265 1997.925 2732.775 1998.735 ;
        RECT 2732.785 1997.925 2734.155 1998.735 ;
        RECT 2695.525 1993.505 2696.895 1994.315 ;
        RECT 2696.905 1993.505 2702.415 1994.315 ;
        RECT 2702.425 1993.505 2707.935 1994.315 ;
        RECT 2708.865 1993.505 2714.375 1994.315 ;
        RECT 2714.385 1993.505 2719.895 1994.315 ;
        RECT 2719.905 1993.505 2725.415 1994.315 ;
        RECT 2725.425 1993.505 2732.775 1994.415 ;
        RECT 2732.785 1993.505 2734.155 1994.315 ;
        RECT 2695.665 1993.295 2695.835 1993.505 ;
        RECT 2697.045 1993.295 2697.215 1993.505 ;
        RECT 2698.425 1993.295 2698.595 1993.485 ;
        RECT 2702.565 1993.315 2702.735 1993.505 ;
        RECT 2703.945 1993.295 2704.115 1993.485 ;
        RECT 2708.080 1993.345 2708.200 1993.455 ;
        RECT 2709.005 1993.315 2709.175 1993.505 ;
        RECT 2709.465 1993.295 2709.635 1993.485 ;
        RECT 2714.525 1993.315 2714.695 1993.505 ;
        RECT 2714.985 1993.295 2715.155 1993.485 ;
        RECT 2720.045 1993.315 2720.215 1993.505 ;
        RECT 2720.515 1993.340 2720.675 1993.450 ;
        RECT 2721.885 1993.295 2722.055 1993.485 ;
        RECT 2725.990 1993.315 2726.160 1993.505 ;
        RECT 2727.405 1993.295 2727.575 1993.485 ;
        RECT 2733.845 1993.295 2734.015 1993.505 ;
        RECT 2695.525 1992.485 2696.895 1993.295 ;
        RECT 2696.905 1992.515 2698.275 1993.295 ;
        RECT 2698.285 1992.485 2703.795 1993.295 ;
        RECT 2703.805 1992.485 2709.315 1993.295 ;
        RECT 2709.325 1992.485 2714.835 1993.295 ;
        RECT 2714.845 1992.485 2720.355 1993.295 ;
        RECT 2721.745 1992.485 2727.255 1993.295 ;
        RECT 2727.265 1992.485 2732.775 1993.295 ;
        RECT 2732.785 1992.485 2734.155 1993.295 ;
        RECT 2695.525 1988.065 2696.895 1988.875 ;
        RECT 2696.905 1988.065 2702.415 1988.875 ;
        RECT 2702.425 1988.065 2707.935 1988.875 ;
        RECT 2708.865 1988.065 2714.375 1988.875 ;
        RECT 2714.385 1988.065 2719.895 1988.875 ;
        RECT 2719.905 1988.065 2725.415 1988.875 ;
        RECT 2725.425 1988.065 2730.935 1988.875 ;
        RECT 2730.945 1988.065 2732.775 1988.875 ;
        RECT 2732.785 1988.065 2734.155 1988.875 ;
        RECT 2695.665 1987.855 2695.835 1988.065 ;
        RECT 2697.045 1987.875 2697.215 1988.065 ;
        RECT 2699.345 1987.875 2699.515 1988.045 ;
        RECT 2699.345 1987.855 2699.475 1987.875 ;
        RECT 2699.805 1987.855 2699.975 1988.045 ;
        RECT 2702.565 1987.875 2702.735 1988.065 ;
        RECT 2705.325 1987.855 2705.495 1988.045 ;
        RECT 2708.080 1987.905 2708.200 1988.015 ;
        RECT 2709.005 1987.875 2709.175 1988.065 ;
        RECT 2710.845 1987.855 2711.015 1988.045 ;
        RECT 2714.525 1987.875 2714.695 1988.065 ;
        RECT 2716.365 1987.855 2716.535 1988.045 ;
        RECT 2720.045 1987.855 2720.215 1988.065 ;
        RECT 2721.885 1987.855 2722.055 1988.045 ;
        RECT 2725.565 1987.875 2725.735 1988.065 ;
        RECT 2727.405 1987.855 2727.575 1988.045 ;
        RECT 2731.085 1987.875 2731.255 1988.065 ;
        RECT 2733.845 1987.855 2734.015 1988.065 ;
        RECT 2695.525 1987.045 2696.895 1987.855 ;
        RECT 2697.625 1987.625 2699.475 1987.855 ;
        RECT 2697.140 1986.945 2699.475 1987.625 ;
        RECT 2699.665 1987.045 2705.175 1987.855 ;
        RECT 2705.185 1987.045 2710.695 1987.855 ;
        RECT 2710.705 1987.045 2716.215 1987.855 ;
        RECT 2716.225 1987.045 2719.895 1987.855 ;
        RECT 2719.905 1987.045 2721.275 1987.855 ;
        RECT 2721.745 1987.045 2727.255 1987.855 ;
        RECT 2727.265 1987.045 2732.775 1987.855 ;
        RECT 2732.785 1987.045 2734.155 1987.855 ;
        RECT 2695.525 1982.625 2696.895 1983.435 ;
        RECT 2696.905 1982.625 2698.275 1983.405 ;
        RECT 2698.285 1982.625 2703.795 1983.435 ;
        RECT 2703.805 1982.625 2707.475 1983.435 ;
        RECT 2708.865 1982.625 2714.375 1983.435 ;
        RECT 2714.385 1982.625 2719.895 1983.435 ;
        RECT 2719.905 1982.625 2725.415 1983.435 ;
        RECT 2725.425 1982.625 2730.935 1983.435 ;
        RECT 2730.945 1982.625 2732.775 1983.435 ;
        RECT 2732.785 1982.625 2734.155 1983.435 ;
        RECT 2695.665 1982.415 2695.835 1982.625 ;
        RECT 2697.045 1982.435 2697.215 1982.625 ;
        RECT 2698.425 1982.435 2698.595 1982.625 ;
        RECT 2700.450 1982.415 2700.620 1982.605 ;
        RECT 2702.575 1982.415 2702.745 1982.585 ;
        RECT 2703.945 1982.435 2704.115 1982.625 ;
        RECT 2704.405 1982.415 2704.575 1982.605 ;
        RECT 2704.865 1982.415 2705.035 1982.605 ;
        RECT 2707.635 1982.470 2707.795 1982.580 ;
        RECT 2709.005 1982.435 2709.175 1982.625 ;
        RECT 2710.385 1982.415 2710.555 1982.605 ;
        RECT 2714.525 1982.435 2714.695 1982.625 ;
        RECT 2715.905 1982.415 2716.075 1982.605 ;
        RECT 2720.045 1982.435 2720.215 1982.625 ;
        RECT 2721.885 1982.415 2722.055 1982.605 ;
        RECT 2725.565 1982.435 2725.735 1982.625 ;
        RECT 2727.405 1982.415 2727.575 1982.605 ;
        RECT 2731.085 1982.435 2731.255 1982.625 ;
        RECT 2733.845 1982.415 2734.015 1982.625 ;
        RECT 2522.700 1981.615 2522.870 1981.785 ;
        RECT 2695.525 1981.605 2696.895 1982.415 ;
        RECT 2697.135 1981.735 2701.035 1982.415 ;
        RECT 2700.105 1981.505 2701.035 1981.735 ;
        RECT 2701.045 1981.505 2704.695 1982.415 ;
        RECT 2704.725 1981.605 2710.235 1982.415 ;
        RECT 2710.245 1981.605 2715.755 1982.415 ;
        RECT 2715.765 1981.605 2721.275 1982.415 ;
        RECT 2721.745 1981.605 2727.255 1982.415 ;
        RECT 2727.265 1981.605 2732.775 1982.415 ;
        RECT 2732.785 1981.605 2734.155 1982.415 ;
        RECT 2695.525 1977.185 2696.895 1977.995 ;
        RECT 2696.905 1977.895 2697.835 1978.095 ;
        RECT 2699.165 1977.895 2700.115 1978.095 ;
        RECT 2696.905 1977.415 2700.115 1977.895 ;
        RECT 2697.050 1977.215 2700.115 1977.415 ;
        RECT 2695.665 1976.975 2695.835 1977.185 ;
        RECT 2697.050 1977.165 2697.220 1977.215 ;
        RECT 2699.180 1977.185 2700.115 1977.215 ;
        RECT 2700.125 1977.185 2705.635 1977.995 ;
        RECT 2705.645 1977.185 2708.395 1977.995 ;
        RECT 2708.865 1977.185 2714.375 1977.995 ;
        RECT 2714.385 1977.185 2719.895 1977.995 ;
        RECT 2719.905 1977.185 2725.415 1977.995 ;
        RECT 2725.425 1977.185 2730.935 1977.995 ;
        RECT 2730.945 1977.185 2732.775 1977.995 ;
        RECT 2732.785 1977.185 2734.155 1977.995 ;
        RECT 2697.045 1976.995 2697.220 1977.165 ;
        RECT 2697.045 1976.975 2697.215 1976.995 ;
        RECT 2698.425 1976.975 2698.595 1977.165 ;
        RECT 2700.265 1976.995 2700.435 1977.185 ;
        RECT 2703.945 1976.975 2704.115 1977.165 ;
        RECT 2705.785 1976.995 2705.955 1977.185 ;
        RECT 2709.005 1976.995 2709.175 1977.185 ;
        RECT 2709.465 1976.975 2709.635 1977.165 ;
        RECT 2714.525 1976.995 2714.695 1977.185 ;
        RECT 2714.985 1976.975 2715.155 1977.165 ;
        RECT 2720.045 1976.995 2720.215 1977.185 ;
        RECT 2720.515 1977.020 2720.675 1977.130 ;
        RECT 2721.885 1976.975 2722.055 1977.165 ;
        RECT 2725.565 1976.995 2725.735 1977.185 ;
        RECT 2727.405 1976.975 2727.575 1977.165 ;
        RECT 2731.085 1976.995 2731.255 1977.185 ;
        RECT 2733.845 1976.975 2734.015 1977.185 ;
        RECT 2695.525 1976.165 2696.895 1976.975 ;
        RECT 2696.905 1976.195 2698.275 1976.975 ;
        RECT 2698.285 1976.165 2703.795 1976.975 ;
        RECT 2703.805 1976.165 2709.315 1976.975 ;
        RECT 2709.325 1976.165 2714.835 1976.975 ;
        RECT 2714.845 1976.165 2720.355 1976.975 ;
        RECT 2721.745 1976.165 2727.255 1976.975 ;
        RECT 2727.265 1976.165 2732.775 1976.975 ;
        RECT 2732.785 1976.165 2734.155 1976.975 ;
        RECT 2522.700 1974.085 2522.870 1974.255 ;
        RECT 2695.525 1971.745 2696.895 1972.555 ;
        RECT 2696.905 1971.745 2698.275 1972.555 ;
        RECT 2698.285 1971.745 2701.955 1972.655 ;
        RECT 2701.965 1971.745 2707.475 1972.555 ;
        RECT 2708.865 1971.745 2714.375 1972.555 ;
        RECT 2714.385 1971.745 2719.895 1972.555 ;
        RECT 2719.905 1971.745 2725.415 1972.555 ;
        RECT 2725.425 1971.745 2730.935 1972.555 ;
        RECT 2730.945 1971.745 2732.775 1972.555 ;
        RECT 2732.785 1971.745 2734.155 1972.555 ;
        RECT 2695.665 1971.535 2695.835 1971.745 ;
        RECT 2697.045 1971.555 2697.215 1971.745 ;
        RECT 2695.525 1970.725 2696.895 1971.535 ;
        RECT 2697.965 1971.505 2698.135 1971.725 ;
        RECT 2701.640 1971.555 2701.810 1971.745 ;
        RECT 2702.105 1971.555 2702.275 1971.745 ;
        RECT 2703.485 1971.535 2703.655 1971.725 ;
        RECT 2703.945 1971.535 2704.115 1971.725 ;
        RECT 2707.635 1971.590 2707.795 1971.700 ;
        RECT 2709.005 1971.555 2709.175 1971.745 ;
        RECT 2709.465 1971.535 2709.635 1971.725 ;
        RECT 2714.525 1971.555 2714.695 1971.745 ;
        RECT 2714.985 1971.535 2715.155 1971.725 ;
        RECT 2720.045 1971.555 2720.215 1971.745 ;
        RECT 2720.515 1971.580 2720.675 1971.690 ;
        RECT 2721.885 1971.535 2722.055 1971.725 ;
        RECT 2725.565 1971.555 2725.735 1971.745 ;
        RECT 2727.405 1971.535 2727.575 1971.725 ;
        RECT 2731.085 1971.555 2731.255 1971.745 ;
        RECT 2733.845 1971.535 2734.015 1971.745 ;
        RECT 2700.090 1971.505 2701.035 1971.535 ;
        RECT 2697.965 1971.305 2701.035 1971.505 ;
        RECT 2697.825 1970.825 2701.035 1971.305 ;
        RECT 2697.825 1970.625 2698.755 1970.825 ;
        RECT 2700.090 1970.625 2701.035 1970.825 ;
        RECT 2701.275 1971.305 2703.655 1971.535 ;
        RECT 2701.275 1970.625 2703.665 1971.305 ;
        RECT 2703.805 1970.725 2709.315 1971.535 ;
        RECT 2709.325 1970.725 2714.835 1971.535 ;
        RECT 2714.845 1970.725 2720.355 1971.535 ;
        RECT 2721.745 1970.725 2727.255 1971.535 ;
        RECT 2727.265 1970.725 2732.775 1971.535 ;
        RECT 2732.785 1970.725 2734.155 1971.535 ;
        RECT 2522.700 1968.105 2522.870 1968.275 ;
        RECT 2695.525 1966.305 2696.895 1967.115 ;
        RECT 2696.905 1966.305 2698.275 1967.085 ;
        RECT 2698.745 1966.305 2700.095 1967.215 ;
        RECT 2700.125 1966.305 2705.635 1967.115 ;
        RECT 2705.645 1966.305 2708.395 1967.115 ;
        RECT 2708.865 1966.305 2714.375 1967.115 ;
        RECT 2714.385 1966.305 2719.895 1967.115 ;
        RECT 2719.905 1966.305 2725.415 1967.115 ;
        RECT 2725.425 1966.305 2730.935 1967.115 ;
        RECT 2730.945 1966.305 2732.775 1967.115 ;
        RECT 2732.785 1966.305 2734.155 1967.115 ;
        RECT 2695.665 1966.095 2695.835 1966.305 ;
        RECT 2697.045 1966.115 2697.215 1966.305 ;
        RECT 2698.420 1966.145 2698.540 1966.255 ;
        RECT 2699.810 1966.115 2699.980 1966.305 ;
        RECT 2700.265 1966.115 2700.435 1966.305 ;
        RECT 2700.450 1966.095 2700.620 1966.285 ;
        RECT 2701.185 1966.095 2701.355 1966.285 ;
        RECT 2705.785 1966.115 2705.955 1966.305 ;
        RECT 2706.705 1966.095 2706.875 1966.285 ;
        RECT 2709.005 1966.115 2709.175 1966.305 ;
        RECT 2712.225 1966.095 2712.395 1966.285 ;
        RECT 2714.525 1966.115 2714.695 1966.305 ;
        RECT 2717.745 1966.095 2717.915 1966.285 ;
        RECT 2720.045 1966.115 2720.215 1966.305 ;
        RECT 2721.885 1966.095 2722.055 1966.285 ;
        RECT 2725.565 1966.115 2725.735 1966.305 ;
        RECT 2727.405 1966.095 2727.575 1966.285 ;
        RECT 2731.085 1966.115 2731.255 1966.305 ;
        RECT 2733.845 1966.095 2734.015 1966.305 ;
        RECT 2695.525 1965.285 2696.895 1966.095 ;
        RECT 2697.135 1965.415 2701.035 1966.095 ;
        RECT 2700.105 1965.185 2701.035 1965.415 ;
        RECT 2701.045 1965.285 2706.555 1966.095 ;
        RECT 2706.565 1965.285 2712.075 1966.095 ;
        RECT 2712.085 1965.285 2717.595 1966.095 ;
        RECT 2717.605 1965.285 2721.275 1966.095 ;
        RECT 2721.745 1965.285 2727.255 1966.095 ;
        RECT 2727.265 1965.285 2732.775 1966.095 ;
        RECT 2732.785 1965.285 2734.155 1966.095 ;
        RECT 2522.700 1962.160 2522.870 1962.330 ;
        RECT 2695.525 1960.865 2696.895 1961.675 ;
        RECT 2696.905 1960.865 2698.275 1961.645 ;
        RECT 2698.285 1960.865 2703.795 1961.675 ;
        RECT 2703.805 1960.865 2707.475 1961.675 ;
        RECT 2708.865 1960.865 2714.375 1961.675 ;
        RECT 2714.385 1960.865 2719.895 1961.675 ;
        RECT 2719.905 1960.865 2725.415 1961.675 ;
        RECT 2725.425 1960.865 2730.935 1961.675 ;
        RECT 2730.945 1960.865 2732.775 1961.675 ;
        RECT 2732.785 1960.865 2734.155 1961.675 ;
        RECT 2695.665 1960.655 2695.835 1960.865 ;
        RECT 2697.045 1960.655 2697.215 1960.865 ;
        RECT 2698.425 1960.675 2698.595 1960.865 ;
        RECT 2702.565 1960.655 2702.735 1960.845 ;
        RECT 2703.945 1960.675 2704.115 1960.865 ;
        RECT 2707.635 1960.710 2707.795 1960.820 ;
        RECT 2708.085 1960.655 2708.255 1960.845 ;
        RECT 2709.005 1960.675 2709.175 1960.865 ;
        RECT 2713.605 1960.655 2713.775 1960.845 ;
        RECT 2714.525 1960.675 2714.695 1960.865 ;
        RECT 2719.125 1960.655 2719.295 1960.845 ;
        RECT 2720.045 1960.675 2720.215 1960.865 ;
        RECT 2720.960 1960.705 2721.080 1960.815 ;
        RECT 2721.885 1960.655 2722.055 1960.845 ;
        RECT 2725.565 1960.675 2725.735 1960.865 ;
        RECT 2727.405 1960.655 2727.575 1960.845 ;
        RECT 2731.085 1960.675 2731.255 1960.865 ;
        RECT 2733.845 1960.655 2734.015 1960.865 ;
        RECT 2695.525 1959.845 2696.895 1960.655 ;
        RECT 2696.905 1959.845 2702.415 1960.655 ;
        RECT 2702.425 1959.845 2707.935 1960.655 ;
        RECT 2707.945 1959.845 2713.455 1960.655 ;
        RECT 2713.465 1959.845 2718.975 1960.655 ;
        RECT 2718.985 1959.845 2720.815 1960.655 ;
        RECT 2721.745 1959.845 2727.255 1960.655 ;
        RECT 2727.265 1959.845 2732.775 1960.655 ;
        RECT 2732.785 1959.845 2734.155 1960.655 ;
        RECT 2522.700 1956.515 2522.870 1956.685 ;
        RECT 2695.525 1955.425 2696.895 1956.235 ;
        RECT 2696.905 1955.425 2698.275 1956.205 ;
        RECT 2698.285 1955.425 2703.795 1956.235 ;
        RECT 2703.805 1955.425 2707.475 1956.235 ;
        RECT 2708.865 1955.425 2714.375 1956.235 ;
        RECT 2714.385 1955.425 2719.895 1956.235 ;
        RECT 2719.905 1955.425 2725.415 1956.235 ;
        RECT 2725.425 1955.425 2730.935 1956.235 ;
        RECT 2730.945 1955.425 2732.775 1956.235 ;
        RECT 2732.785 1955.425 2734.155 1956.235 ;
        RECT 2695.665 1955.215 2695.835 1955.425 ;
        RECT 2697.045 1955.215 2697.215 1955.425 ;
        RECT 2698.425 1955.235 2698.595 1955.425 ;
        RECT 2702.565 1955.215 2702.735 1955.405 ;
        RECT 2703.945 1955.235 2704.115 1955.425 ;
        RECT 2707.635 1955.270 2707.795 1955.380 ;
        RECT 2708.085 1955.215 2708.255 1955.405 ;
        RECT 2709.005 1955.235 2709.175 1955.425 ;
        RECT 2713.605 1955.215 2713.775 1955.405 ;
        RECT 2714.525 1955.235 2714.695 1955.425 ;
        RECT 2719.125 1955.215 2719.295 1955.405 ;
        RECT 2720.045 1955.235 2720.215 1955.425 ;
        RECT 2720.960 1955.265 2721.080 1955.375 ;
        RECT 2721.885 1955.215 2722.055 1955.405 ;
        RECT 2725.565 1955.235 2725.735 1955.425 ;
        RECT 2727.405 1955.215 2727.575 1955.405 ;
        RECT 2731.085 1955.235 2731.255 1955.425 ;
        RECT 2733.845 1955.215 2734.015 1955.425 ;
        RECT 2695.525 1954.405 2696.895 1955.215 ;
        RECT 2696.905 1954.405 2702.415 1955.215 ;
        RECT 2702.425 1954.405 2707.935 1955.215 ;
        RECT 2707.945 1954.405 2713.455 1955.215 ;
        RECT 2713.465 1954.405 2718.975 1955.215 ;
        RECT 2718.985 1954.405 2720.815 1955.215 ;
        RECT 2721.745 1954.405 2727.255 1955.215 ;
        RECT 2727.265 1954.405 2732.775 1955.215 ;
        RECT 2732.785 1954.405 2734.155 1955.215 ;
        RECT 2522.700 1950.510 2522.870 1950.680 ;
        RECT 2695.525 1949.985 2696.895 1950.795 ;
        RECT 2696.905 1949.985 2698.275 1950.765 ;
        RECT 2698.285 1949.985 2699.655 1950.765 ;
        RECT 2699.665 1949.985 2705.175 1950.795 ;
        RECT 2705.185 1949.985 2707.935 1950.795 ;
        RECT 2708.865 1949.985 2714.375 1950.795 ;
        RECT 2714.385 1949.985 2719.895 1950.795 ;
        RECT 2719.905 1949.985 2721.275 1950.795 ;
        RECT 2721.745 1949.985 2727.255 1950.795 ;
        RECT 2727.265 1949.985 2732.775 1950.795 ;
        RECT 2732.785 1949.985 2734.155 1950.795 ;
        RECT 2695.665 1949.795 2695.835 1949.985 ;
        RECT 2697.045 1949.795 2697.215 1949.985 ;
        RECT 2698.425 1949.795 2698.595 1949.985 ;
        RECT 2699.805 1949.795 2699.975 1949.985 ;
        RECT 2705.325 1949.795 2705.495 1949.985 ;
        RECT 2708.080 1949.825 2708.200 1949.935 ;
        RECT 2709.005 1949.795 2709.175 1949.985 ;
        RECT 2714.525 1949.795 2714.695 1949.985 ;
        RECT 2720.045 1949.795 2720.215 1949.985 ;
        RECT 2721.885 1949.795 2722.055 1949.985 ;
        RECT 2727.405 1949.795 2727.575 1949.985 ;
        RECT 2733.845 1949.795 2734.015 1949.985 ;
        RECT 2361.705 1945.735 2361.875 1945.875 ;
        RECT 2361.685 1945.715 2361.875 1945.735 ;
        RECT 2361.685 1945.705 2361.855 1945.715 ;
        RECT 2363.665 1945.705 2363.835 1945.875 ;
        RECT 2366.105 1945.705 2366.275 1945.875 ;
        RECT 2368.545 1945.705 2368.715 1945.875 ;
        RECT 2370.505 1945.705 2370.675 1945.875 ;
        RECT 2380.265 1945.735 2380.435 1945.875 ;
        RECT 2380.245 1945.715 2380.435 1945.735 ;
        RECT 2380.245 1945.705 2380.415 1945.715 ;
        RECT 2382.225 1945.705 2382.395 1945.875 ;
        RECT 2384.665 1945.705 2384.835 1945.875 ;
        RECT 2387.105 1945.705 2387.275 1945.875 ;
        RECT 2389.065 1945.705 2389.235 1945.875 ;
        RECT 2398.825 1945.735 2398.995 1945.875 ;
        RECT 2398.805 1945.715 2398.995 1945.735 ;
        RECT 2398.805 1945.705 2398.975 1945.715 ;
        RECT 2400.785 1945.705 2400.955 1945.875 ;
        RECT 2403.225 1945.705 2403.395 1945.875 ;
        RECT 2405.665 1945.705 2405.835 1945.875 ;
        RECT 2407.625 1945.705 2407.795 1945.875 ;
        RECT 2417.385 1945.735 2417.555 1945.875 ;
        RECT 2417.365 1945.715 2417.555 1945.735 ;
        RECT 2417.365 1945.705 2417.535 1945.715 ;
        RECT 2419.345 1945.705 2419.515 1945.875 ;
        RECT 2421.785 1945.705 2421.955 1945.875 ;
        RECT 2424.225 1945.705 2424.395 1945.875 ;
        RECT 2426.185 1945.705 2426.355 1945.875 ;
        RECT 2435.945 1945.735 2436.115 1945.875 ;
        RECT 2435.925 1945.715 2436.115 1945.735 ;
        RECT 2435.925 1945.705 2436.095 1945.715 ;
        RECT 2437.905 1945.705 2438.075 1945.875 ;
        RECT 2440.345 1945.705 2440.515 1945.875 ;
        RECT 2442.785 1945.705 2442.955 1945.875 ;
        RECT 2444.745 1945.705 2444.915 1945.875 ;
        RECT 2883.065 1891.500 2883.235 1891.670 ;
        RECT 2695.665 1856.815 2695.835 1857.005 ;
        RECT 2697.045 1856.815 2697.215 1857.005 ;
        RECT 2699.805 1856.815 2699.975 1857.005 ;
        RECT 2701.185 1856.815 2701.355 1857.005 ;
        RECT 2701.645 1856.815 2701.815 1857.005 ;
        RECT 2707.165 1856.815 2707.335 1857.005 ;
        RECT 2709.005 1856.815 2709.175 1857.005 ;
        RECT 2710.845 1856.815 2711.015 1857.005 ;
        RECT 2716.365 1856.815 2716.535 1857.005 ;
        RECT 2720.045 1856.815 2720.215 1857.005 ;
        RECT 2723.265 1856.815 2723.435 1857.005 ;
        RECT 2723.725 1856.815 2723.895 1857.005 ;
        RECT 2729.245 1856.815 2729.415 1857.005 ;
        RECT 2731.080 1856.865 2731.200 1856.975 ;
        RECT 2732.455 1856.815 2732.625 1857.005 ;
        RECT 2733.845 1856.815 2734.015 1857.005 ;
        RECT 2695.525 1856.005 2696.895 1856.815 ;
        RECT 2696.905 1856.135 2698.735 1856.815 ;
        RECT 2698.745 1856.035 2700.115 1856.815 ;
        RECT 2700.125 1856.035 2701.495 1856.815 ;
        RECT 2701.505 1856.005 2707.015 1856.815 ;
        RECT 2707.025 1856.005 2708.395 1856.815 ;
        RECT 2708.865 1856.135 2710.695 1856.815 ;
        RECT 2709.350 1855.905 2710.695 1856.135 ;
        RECT 2710.705 1856.005 2716.215 1856.815 ;
        RECT 2716.225 1856.005 2719.895 1856.815 ;
        RECT 2719.905 1856.005 2721.275 1856.815 ;
        RECT 2721.745 1856.135 2723.575 1856.815 ;
        RECT 2723.585 1856.005 2729.095 1856.815 ;
        RECT 2729.105 1856.005 2730.935 1856.815 ;
        RECT 2731.405 1856.035 2732.775 1856.815 ;
        RECT 2732.785 1856.005 2734.155 1856.815 ;
        RECT 2695.525 1851.585 2696.895 1852.395 ;
        RECT 2696.905 1851.585 2698.275 1852.365 ;
        RECT 2698.285 1851.585 2703.795 1852.395 ;
        RECT 2703.805 1851.585 2707.475 1852.395 ;
        RECT 2708.865 1851.585 2714.375 1852.395 ;
        RECT 2714.385 1851.585 2719.895 1852.395 ;
        RECT 2719.905 1851.585 2725.415 1852.395 ;
        RECT 2725.425 1851.585 2730.935 1852.395 ;
        RECT 2730.945 1851.585 2732.775 1852.395 ;
        RECT 2732.785 1851.585 2734.155 1852.395 ;
        RECT 2695.665 1851.375 2695.835 1851.585 ;
        RECT 2697.045 1851.375 2697.215 1851.585 ;
        RECT 2698.425 1851.395 2698.595 1851.585 ;
        RECT 2702.565 1851.375 2702.735 1851.565 ;
        RECT 2703.945 1851.395 2704.115 1851.585 ;
        RECT 2707.635 1851.430 2707.795 1851.540 ;
        RECT 2708.085 1851.375 2708.255 1851.565 ;
        RECT 2709.005 1851.395 2709.175 1851.585 ;
        RECT 2713.605 1851.375 2713.775 1851.565 ;
        RECT 2714.525 1851.395 2714.695 1851.585 ;
        RECT 2719.125 1851.375 2719.295 1851.565 ;
        RECT 2720.045 1851.395 2720.215 1851.585 ;
        RECT 2720.960 1851.425 2721.080 1851.535 ;
        RECT 2721.885 1851.375 2722.055 1851.565 ;
        RECT 2725.565 1851.395 2725.735 1851.585 ;
        RECT 2727.405 1851.375 2727.575 1851.565 ;
        RECT 2731.085 1851.395 2731.255 1851.585 ;
        RECT 2733.845 1851.375 2734.015 1851.585 ;
        RECT 2695.525 1850.565 2696.895 1851.375 ;
        RECT 2696.905 1850.565 2702.415 1851.375 ;
        RECT 2702.425 1850.565 2707.935 1851.375 ;
        RECT 2707.945 1850.565 2713.455 1851.375 ;
        RECT 2713.465 1850.565 2718.975 1851.375 ;
        RECT 2718.985 1850.565 2720.815 1851.375 ;
        RECT 2721.745 1850.565 2727.255 1851.375 ;
        RECT 2727.265 1850.565 2732.775 1851.375 ;
        RECT 2732.785 1850.565 2734.155 1851.375 ;
        RECT 2695.525 1846.145 2696.895 1846.955 ;
        RECT 2696.905 1846.145 2702.415 1846.955 ;
        RECT 2702.425 1846.145 2707.935 1846.955 ;
        RECT 2708.865 1846.145 2714.375 1846.955 ;
        RECT 2714.385 1846.145 2719.895 1846.955 ;
        RECT 2719.905 1846.145 2725.415 1846.955 ;
        RECT 2725.425 1846.145 2730.935 1846.955 ;
        RECT 2730.945 1846.145 2732.775 1846.955 ;
        RECT 2732.785 1846.145 2734.155 1846.955 ;
        RECT 2695.665 1845.935 2695.835 1846.145 ;
        RECT 2697.045 1845.935 2697.215 1846.145 ;
        RECT 2698.425 1845.935 2698.595 1846.125 ;
        RECT 2702.565 1845.955 2702.735 1846.145 ;
        RECT 2703.945 1845.935 2704.115 1846.125 ;
        RECT 2708.080 1845.985 2708.200 1846.095 ;
        RECT 2709.005 1845.955 2709.175 1846.145 ;
        RECT 2709.465 1845.935 2709.635 1846.125 ;
        RECT 2714.525 1845.955 2714.695 1846.145 ;
        RECT 2714.985 1845.935 2715.155 1846.125 ;
        RECT 2720.045 1845.955 2720.215 1846.145 ;
        RECT 2720.515 1845.980 2720.675 1846.090 ;
        RECT 2721.885 1845.935 2722.055 1846.125 ;
        RECT 2725.565 1845.955 2725.735 1846.145 ;
        RECT 2727.405 1845.935 2727.575 1846.125 ;
        RECT 2731.085 1845.955 2731.255 1846.145 ;
        RECT 2733.845 1845.935 2734.015 1846.145 ;
        RECT 2695.525 1845.125 2696.895 1845.935 ;
        RECT 2696.905 1845.155 2698.275 1845.935 ;
        RECT 2698.285 1845.125 2703.795 1845.935 ;
        RECT 2703.805 1845.125 2709.315 1845.935 ;
        RECT 2709.325 1845.125 2714.835 1845.935 ;
        RECT 2714.845 1845.125 2720.355 1845.935 ;
        RECT 2721.745 1845.125 2727.255 1845.935 ;
        RECT 2727.265 1845.125 2732.775 1845.935 ;
        RECT 2732.785 1845.125 2734.155 1845.935 ;
        RECT 2695.525 1840.705 2696.895 1841.515 ;
        RECT 2696.905 1840.705 2702.415 1841.515 ;
        RECT 2702.425 1840.705 2707.935 1841.515 ;
        RECT 2708.865 1840.705 2714.375 1841.515 ;
        RECT 2714.385 1840.705 2719.895 1841.515 ;
        RECT 2719.905 1840.705 2725.415 1841.515 ;
        RECT 2725.425 1840.705 2730.935 1841.515 ;
        RECT 2730.945 1840.705 2732.775 1841.515 ;
        RECT 2732.785 1840.705 2734.155 1841.515 ;
        RECT 2695.665 1840.495 2695.835 1840.705 ;
        RECT 2697.045 1840.495 2697.215 1840.705 ;
        RECT 2702.565 1840.515 2702.735 1840.705 ;
        RECT 2706.705 1840.495 2706.875 1840.685 ;
        RECT 2708.080 1840.545 2708.200 1840.655 ;
        RECT 2709.005 1840.515 2709.175 1840.705 ;
        RECT 2712.225 1840.495 2712.395 1840.685 ;
        RECT 2714.525 1840.515 2714.695 1840.705 ;
        RECT 2717.745 1840.495 2717.915 1840.685 ;
        RECT 2720.045 1840.515 2720.215 1840.705 ;
        RECT 2721.885 1840.495 2722.055 1840.685 ;
        RECT 2725.565 1840.515 2725.735 1840.705 ;
        RECT 2727.405 1840.495 2727.575 1840.685 ;
        RECT 2731.085 1840.515 2731.255 1840.705 ;
        RECT 2733.845 1840.495 2734.015 1840.705 ;
        RECT 2695.525 1839.685 2696.895 1840.495 ;
        RECT 2696.905 1840.325 2698.665 1840.495 ;
        RECT 2696.905 1840.280 2699.160 1840.325 ;
        RECT 2696.905 1840.245 2700.100 1840.280 ;
        RECT 2701.460 1840.245 2706.555 1840.495 ;
        RECT 2696.905 1839.815 2706.555 1840.245 ;
        RECT 2698.230 1839.645 2701.460 1839.815 ;
        RECT 2699.170 1839.600 2701.460 1839.645 ;
        RECT 2700.110 1839.565 2701.460 1839.600 ;
        RECT 2704.535 1839.585 2706.555 1839.815 ;
        RECT 2706.565 1839.685 2712.075 1840.495 ;
        RECT 2712.085 1839.685 2717.595 1840.495 ;
        RECT 2717.605 1839.685 2721.275 1840.495 ;
        RECT 2721.745 1839.685 2727.255 1840.495 ;
        RECT 2727.265 1839.685 2732.775 1840.495 ;
        RECT 2732.785 1839.685 2734.155 1840.495 ;
        RECT 2704.535 1839.565 2705.455 1839.585 ;
        RECT 2695.525 1835.265 2696.895 1836.075 ;
        RECT 2696.905 1835.265 2698.275 1836.045 ;
        RECT 2698.285 1835.265 2703.795 1836.075 ;
        RECT 2703.805 1835.265 2707.475 1836.075 ;
        RECT 2708.865 1835.265 2714.375 1836.075 ;
        RECT 2714.385 1835.265 2719.895 1836.075 ;
        RECT 2719.905 1835.265 2725.415 1836.075 ;
        RECT 2725.425 1835.265 2730.935 1836.075 ;
        RECT 2730.945 1835.265 2732.775 1836.075 ;
        RECT 2732.785 1835.265 2734.155 1836.075 ;
        RECT 2695.665 1835.055 2695.835 1835.265 ;
        RECT 2697.045 1835.055 2697.215 1835.265 ;
        RECT 2698.425 1835.075 2698.595 1835.265 ;
        RECT 2703.945 1835.075 2704.115 1835.265 ;
        RECT 2706.705 1835.055 2706.875 1835.245 ;
        RECT 2707.635 1835.110 2707.795 1835.220 ;
        RECT 2709.005 1835.075 2709.175 1835.265 ;
        RECT 2712.225 1835.055 2712.395 1835.245 ;
        RECT 2714.525 1835.075 2714.695 1835.265 ;
        RECT 2717.745 1835.055 2717.915 1835.245 ;
        RECT 2720.045 1835.075 2720.215 1835.265 ;
        RECT 2721.885 1835.055 2722.055 1835.245 ;
        RECT 2725.565 1835.075 2725.735 1835.265 ;
        RECT 2727.405 1835.055 2727.575 1835.245 ;
        RECT 2731.085 1835.075 2731.255 1835.265 ;
        RECT 2733.845 1835.055 2734.015 1835.265 ;
        RECT 2695.525 1834.245 2696.895 1835.055 ;
        RECT 2696.905 1834.885 2698.665 1835.055 ;
        RECT 2696.905 1834.840 2699.160 1834.885 ;
        RECT 2696.905 1834.805 2700.100 1834.840 ;
        RECT 2701.460 1834.805 2706.555 1835.055 ;
        RECT 2696.905 1834.375 2706.555 1834.805 ;
        RECT 2698.230 1834.205 2701.460 1834.375 ;
        RECT 2699.170 1834.160 2701.460 1834.205 ;
        RECT 2700.110 1834.125 2701.460 1834.160 ;
        RECT 2704.535 1834.145 2706.555 1834.375 ;
        RECT 2706.565 1834.245 2712.075 1835.055 ;
        RECT 2712.085 1834.245 2717.595 1835.055 ;
        RECT 2717.605 1834.245 2721.275 1835.055 ;
        RECT 2721.745 1834.245 2727.255 1835.055 ;
        RECT 2727.265 1834.245 2732.775 1835.055 ;
        RECT 2732.785 1834.245 2734.155 1835.055 ;
        RECT 2704.535 1834.125 2705.455 1834.145 ;
        RECT 2695.525 1829.825 2696.895 1830.635 ;
        RECT 2696.905 1829.825 2698.275 1830.605 ;
        RECT 2698.285 1829.825 2701.035 1830.635 ;
        RECT 2701.505 1830.505 2702.435 1830.735 ;
        RECT 2701.505 1829.825 2705.405 1830.505 ;
        RECT 2705.645 1829.825 2708.395 1830.635 ;
        RECT 2708.865 1829.825 2714.375 1830.635 ;
        RECT 2714.385 1829.825 2719.895 1830.635 ;
        RECT 2719.905 1829.825 2725.415 1830.635 ;
        RECT 2725.425 1829.825 2730.935 1830.635 ;
        RECT 2730.945 1829.825 2732.775 1830.635 ;
        RECT 2732.785 1829.825 2734.155 1830.635 ;
        RECT 2695.665 1829.615 2695.835 1829.825 ;
        RECT 2697.045 1829.615 2697.215 1829.825 ;
        RECT 2698.425 1829.635 2698.595 1829.825 ;
        RECT 2701.180 1829.665 2701.300 1829.775 ;
        RECT 2701.920 1829.635 2702.090 1829.825 ;
        RECT 2702.565 1829.615 2702.735 1829.805 ;
        RECT 2705.785 1829.635 2705.955 1829.825 ;
        RECT 2708.085 1829.615 2708.255 1829.805 ;
        RECT 2709.005 1829.635 2709.175 1829.825 ;
        RECT 2713.605 1829.615 2713.775 1829.805 ;
        RECT 2714.525 1829.635 2714.695 1829.825 ;
        RECT 2719.125 1829.615 2719.295 1829.805 ;
        RECT 2720.045 1829.635 2720.215 1829.825 ;
        RECT 2720.960 1829.665 2721.080 1829.775 ;
        RECT 2721.885 1829.615 2722.055 1829.805 ;
        RECT 2725.565 1829.635 2725.735 1829.825 ;
        RECT 2727.405 1829.615 2727.575 1829.805 ;
        RECT 2731.085 1829.635 2731.255 1829.825 ;
        RECT 2733.845 1829.615 2734.015 1829.825 ;
        RECT 2695.525 1828.805 2696.895 1829.615 ;
        RECT 2696.905 1828.805 2702.415 1829.615 ;
        RECT 2702.425 1828.805 2707.935 1829.615 ;
        RECT 2707.945 1828.805 2713.455 1829.615 ;
        RECT 2713.465 1828.805 2718.975 1829.615 ;
        RECT 2718.985 1828.805 2720.815 1829.615 ;
        RECT 2721.745 1828.805 2727.255 1829.615 ;
        RECT 2727.265 1828.805 2732.775 1829.615 ;
        RECT 2732.785 1828.805 2734.155 1829.615 ;
        RECT 2695.525 1824.385 2696.895 1825.195 ;
        RECT 2696.905 1824.385 2698.275 1825.165 ;
        RECT 2698.285 1824.385 2703.795 1825.195 ;
        RECT 2703.805 1824.385 2707.475 1825.195 ;
        RECT 2708.865 1824.385 2714.375 1825.195 ;
        RECT 2714.385 1824.385 2719.895 1825.195 ;
        RECT 2719.905 1824.385 2725.415 1825.195 ;
        RECT 2725.425 1824.385 2730.935 1825.195 ;
        RECT 2730.945 1824.385 2732.775 1825.195 ;
        RECT 2732.785 1824.385 2734.155 1825.195 ;
        RECT 2695.665 1824.175 2695.835 1824.385 ;
        RECT 2697.045 1824.175 2697.215 1824.385 ;
        RECT 2698.425 1824.195 2698.595 1824.385 ;
        RECT 2702.565 1824.175 2702.735 1824.365 ;
        RECT 2703.945 1824.195 2704.115 1824.385 ;
        RECT 2707.635 1824.230 2707.795 1824.340 ;
        RECT 2708.085 1824.175 2708.255 1824.365 ;
        RECT 2709.005 1824.195 2709.175 1824.385 ;
        RECT 2713.605 1824.175 2713.775 1824.365 ;
        RECT 2714.525 1824.195 2714.695 1824.385 ;
        RECT 2719.125 1824.175 2719.295 1824.365 ;
        RECT 2720.045 1824.195 2720.215 1824.385 ;
        RECT 2720.960 1824.225 2721.080 1824.335 ;
        RECT 2721.885 1824.175 2722.055 1824.365 ;
        RECT 2725.565 1824.195 2725.735 1824.385 ;
        RECT 2727.405 1824.175 2727.575 1824.365 ;
        RECT 2731.085 1824.195 2731.255 1824.385 ;
        RECT 2733.845 1824.175 2734.015 1824.385 ;
        RECT 2695.525 1823.365 2696.895 1824.175 ;
        RECT 2696.905 1823.365 2702.415 1824.175 ;
        RECT 2702.425 1823.365 2707.935 1824.175 ;
        RECT 2707.945 1823.365 2713.455 1824.175 ;
        RECT 2713.465 1823.365 2718.975 1824.175 ;
        RECT 2718.985 1823.365 2720.815 1824.175 ;
        RECT 2721.745 1823.365 2727.255 1824.175 ;
        RECT 2727.265 1823.365 2732.775 1824.175 ;
        RECT 2732.785 1823.365 2734.155 1824.175 ;
        RECT 2695.525 1818.945 2696.895 1819.755 ;
        RECT 2696.905 1818.945 2700.575 1819.755 ;
        RECT 2701.505 1818.945 2702.855 1819.855 ;
        RECT 2702.885 1818.945 2708.395 1819.755 ;
        RECT 2708.865 1818.945 2714.375 1819.755 ;
        RECT 2714.385 1818.945 2719.895 1819.755 ;
        RECT 2719.905 1818.945 2725.415 1819.755 ;
        RECT 2725.425 1818.945 2730.935 1819.755 ;
        RECT 2730.945 1818.945 2732.775 1819.755 ;
        RECT 2732.785 1818.945 2734.155 1819.755 ;
        RECT 2695.665 1818.735 2695.835 1818.945 ;
        RECT 2697.045 1818.735 2697.215 1818.945 ;
        RECT 2698.425 1818.735 2698.595 1818.925 ;
        RECT 2700.735 1818.790 2700.895 1818.900 ;
        RECT 2701.650 1818.755 2701.820 1818.945 ;
        RECT 2703.025 1818.755 2703.195 1818.945 ;
        RECT 2704.865 1818.735 2705.035 1818.925 ;
        RECT 2705.325 1818.735 2705.495 1818.925 ;
        RECT 2709.005 1818.755 2709.175 1818.945 ;
        RECT 2710.845 1818.735 2711.015 1818.925 ;
        RECT 2714.525 1818.755 2714.695 1818.945 ;
        RECT 2716.365 1818.735 2716.535 1818.925 ;
        RECT 2720.045 1818.735 2720.215 1818.945 ;
        RECT 2721.885 1818.735 2722.055 1818.925 ;
        RECT 2725.565 1818.755 2725.735 1818.945 ;
        RECT 2727.405 1818.735 2727.575 1818.925 ;
        RECT 2731.085 1818.755 2731.255 1818.945 ;
        RECT 2733.845 1818.735 2734.015 1818.945 ;
        RECT 2695.525 1817.925 2696.895 1818.735 ;
        RECT 2696.905 1817.955 2698.275 1818.735 ;
        RECT 2698.285 1817.925 2701.955 1818.735 ;
        RECT 2701.965 1817.825 2705.175 1818.735 ;
        RECT 2705.185 1817.925 2710.695 1818.735 ;
        RECT 2710.705 1817.925 2716.215 1818.735 ;
        RECT 2716.225 1817.925 2719.895 1818.735 ;
        RECT 2719.905 1817.925 2721.275 1818.735 ;
        RECT 2721.745 1817.925 2727.255 1818.735 ;
        RECT 2727.265 1817.925 2732.775 1818.735 ;
        RECT 2732.785 1817.925 2734.155 1818.735 ;
        RECT 2695.525 1813.505 2696.895 1814.315 ;
        RECT 2696.905 1813.505 2702.415 1814.315 ;
        RECT 2702.425 1813.505 2707.935 1814.315 ;
        RECT 2708.865 1813.505 2714.375 1814.315 ;
        RECT 2714.385 1813.505 2719.895 1814.315 ;
        RECT 2719.905 1813.505 2725.415 1814.315 ;
        RECT 2725.425 1813.505 2732.775 1814.415 ;
        RECT 2732.785 1813.505 2734.155 1814.315 ;
        RECT 2695.665 1813.295 2695.835 1813.505 ;
        RECT 2697.045 1813.295 2697.215 1813.505 ;
        RECT 2698.425 1813.295 2698.595 1813.485 ;
        RECT 2702.565 1813.315 2702.735 1813.505 ;
        RECT 2703.945 1813.295 2704.115 1813.485 ;
        RECT 2708.080 1813.345 2708.200 1813.455 ;
        RECT 2709.005 1813.315 2709.175 1813.505 ;
        RECT 2709.465 1813.295 2709.635 1813.485 ;
        RECT 2714.525 1813.315 2714.695 1813.505 ;
        RECT 2714.985 1813.295 2715.155 1813.485 ;
        RECT 2720.045 1813.315 2720.215 1813.505 ;
        RECT 2720.515 1813.340 2720.675 1813.450 ;
        RECT 2721.885 1813.295 2722.055 1813.485 ;
        RECT 2725.990 1813.315 2726.160 1813.505 ;
        RECT 2727.405 1813.295 2727.575 1813.485 ;
        RECT 2733.845 1813.295 2734.015 1813.505 ;
        RECT 2695.525 1812.485 2696.895 1813.295 ;
        RECT 2696.905 1812.515 2698.275 1813.295 ;
        RECT 2698.285 1812.485 2703.795 1813.295 ;
        RECT 2703.805 1812.485 2709.315 1813.295 ;
        RECT 2709.325 1812.485 2714.835 1813.295 ;
        RECT 2714.845 1812.485 2720.355 1813.295 ;
        RECT 2721.745 1812.485 2727.255 1813.295 ;
        RECT 2727.265 1812.485 2732.775 1813.295 ;
        RECT 2732.785 1812.485 2734.155 1813.295 ;
        RECT 2695.525 1808.065 2696.895 1808.875 ;
        RECT 2696.905 1808.065 2702.415 1808.875 ;
        RECT 2702.425 1808.065 2707.935 1808.875 ;
        RECT 2708.865 1808.065 2714.375 1808.875 ;
        RECT 2714.385 1808.065 2719.895 1808.875 ;
        RECT 2719.905 1808.065 2725.415 1808.875 ;
        RECT 2725.425 1808.065 2730.935 1808.875 ;
        RECT 2730.945 1808.065 2732.775 1808.875 ;
        RECT 2732.785 1808.065 2734.155 1808.875 ;
        RECT 2695.665 1807.855 2695.835 1808.065 ;
        RECT 2697.045 1807.875 2697.215 1808.065 ;
        RECT 2699.345 1807.875 2699.515 1808.045 ;
        RECT 2699.345 1807.855 2699.475 1807.875 ;
        RECT 2699.805 1807.855 2699.975 1808.045 ;
        RECT 2702.565 1807.875 2702.735 1808.065 ;
        RECT 2705.325 1807.855 2705.495 1808.045 ;
        RECT 2708.080 1807.905 2708.200 1808.015 ;
        RECT 2709.005 1807.875 2709.175 1808.065 ;
        RECT 2710.845 1807.855 2711.015 1808.045 ;
        RECT 2714.525 1807.875 2714.695 1808.065 ;
        RECT 2716.365 1807.855 2716.535 1808.045 ;
        RECT 2720.045 1807.855 2720.215 1808.065 ;
        RECT 2721.885 1807.855 2722.055 1808.045 ;
        RECT 2725.565 1807.875 2725.735 1808.065 ;
        RECT 2727.405 1807.855 2727.575 1808.045 ;
        RECT 2731.085 1807.875 2731.255 1808.065 ;
        RECT 2733.845 1807.855 2734.015 1808.065 ;
        RECT 2695.525 1807.045 2696.895 1807.855 ;
        RECT 2697.625 1807.625 2699.475 1807.855 ;
        RECT 2697.140 1806.945 2699.475 1807.625 ;
        RECT 2699.665 1807.045 2705.175 1807.855 ;
        RECT 2705.185 1807.045 2710.695 1807.855 ;
        RECT 2710.705 1807.045 2716.215 1807.855 ;
        RECT 2716.225 1807.045 2719.895 1807.855 ;
        RECT 2719.905 1807.045 2721.275 1807.855 ;
        RECT 2721.745 1807.045 2727.255 1807.855 ;
        RECT 2727.265 1807.045 2732.775 1807.855 ;
        RECT 2732.785 1807.045 2734.155 1807.855 ;
        RECT 2522.700 1804.645 2522.870 1804.815 ;
        RECT 2695.525 1802.625 2696.895 1803.435 ;
        RECT 2696.905 1802.625 2698.275 1803.405 ;
        RECT 2698.285 1802.625 2703.795 1803.435 ;
        RECT 2703.805 1802.625 2707.475 1803.435 ;
        RECT 2708.865 1802.625 2714.375 1803.435 ;
        RECT 2714.385 1802.625 2719.895 1803.435 ;
        RECT 2719.905 1802.625 2725.415 1803.435 ;
        RECT 2725.425 1802.625 2730.935 1803.435 ;
        RECT 2730.945 1802.625 2732.775 1803.435 ;
        RECT 2732.785 1802.625 2734.155 1803.435 ;
        RECT 2695.665 1802.415 2695.835 1802.625 ;
        RECT 2697.045 1802.435 2697.215 1802.625 ;
        RECT 2698.425 1802.435 2698.595 1802.625 ;
        RECT 2700.450 1802.415 2700.620 1802.605 ;
        RECT 2702.575 1802.415 2702.745 1802.585 ;
        RECT 2703.945 1802.435 2704.115 1802.625 ;
        RECT 2704.405 1802.415 2704.575 1802.605 ;
        RECT 2704.865 1802.415 2705.035 1802.605 ;
        RECT 2707.635 1802.470 2707.795 1802.580 ;
        RECT 2709.005 1802.435 2709.175 1802.625 ;
        RECT 2710.385 1802.415 2710.555 1802.605 ;
        RECT 2714.525 1802.435 2714.695 1802.625 ;
        RECT 2715.905 1802.415 2716.075 1802.605 ;
        RECT 2720.045 1802.435 2720.215 1802.625 ;
        RECT 2721.885 1802.415 2722.055 1802.605 ;
        RECT 2725.565 1802.435 2725.735 1802.625 ;
        RECT 2727.405 1802.415 2727.575 1802.605 ;
        RECT 2731.085 1802.435 2731.255 1802.625 ;
        RECT 2733.845 1802.415 2734.015 1802.625 ;
        RECT 2695.525 1801.605 2696.895 1802.415 ;
        RECT 2697.135 1801.735 2701.035 1802.415 ;
        RECT 2700.105 1801.505 2701.035 1801.735 ;
        RECT 2701.045 1801.505 2704.695 1802.415 ;
        RECT 2704.725 1801.605 2710.235 1802.415 ;
        RECT 2710.245 1801.605 2715.755 1802.415 ;
        RECT 2715.765 1801.605 2721.275 1802.415 ;
        RECT 2721.745 1801.605 2727.255 1802.415 ;
        RECT 2727.265 1801.605 2732.775 1802.415 ;
        RECT 2732.785 1801.605 2734.155 1802.415 ;
        RECT 2522.700 1797.115 2522.870 1797.285 ;
        RECT 2695.525 1797.185 2696.895 1797.995 ;
        RECT 2696.905 1797.895 2697.835 1798.095 ;
        RECT 2699.165 1797.895 2700.115 1798.095 ;
        RECT 2696.905 1797.415 2700.115 1797.895 ;
        RECT 2697.050 1797.215 2700.115 1797.415 ;
        RECT 2695.665 1796.975 2695.835 1797.185 ;
        RECT 2697.050 1797.165 2697.220 1797.215 ;
        RECT 2699.180 1797.185 2700.115 1797.215 ;
        RECT 2700.125 1797.185 2705.635 1797.995 ;
        RECT 2705.645 1797.185 2708.395 1797.995 ;
        RECT 2708.865 1797.185 2714.375 1797.995 ;
        RECT 2714.385 1797.185 2719.895 1797.995 ;
        RECT 2719.905 1797.185 2725.415 1797.995 ;
        RECT 2725.425 1797.185 2730.935 1797.995 ;
        RECT 2730.945 1797.185 2732.775 1797.995 ;
        RECT 2732.785 1797.185 2734.155 1797.995 ;
        RECT 2697.045 1796.995 2697.220 1797.165 ;
        RECT 2697.045 1796.975 2697.215 1796.995 ;
        RECT 2698.425 1796.975 2698.595 1797.165 ;
        RECT 2700.265 1796.995 2700.435 1797.185 ;
        RECT 2703.945 1796.975 2704.115 1797.165 ;
        RECT 2705.785 1796.995 2705.955 1797.185 ;
        RECT 2709.005 1796.995 2709.175 1797.185 ;
        RECT 2709.465 1796.975 2709.635 1797.165 ;
        RECT 2714.525 1796.995 2714.695 1797.185 ;
        RECT 2714.985 1796.975 2715.155 1797.165 ;
        RECT 2720.045 1796.995 2720.215 1797.185 ;
        RECT 2720.515 1797.020 2720.675 1797.130 ;
        RECT 2721.885 1796.975 2722.055 1797.165 ;
        RECT 2725.565 1796.995 2725.735 1797.185 ;
        RECT 2727.405 1796.975 2727.575 1797.165 ;
        RECT 2731.085 1796.995 2731.255 1797.185 ;
        RECT 2733.845 1796.975 2734.015 1797.185 ;
        RECT 2695.525 1796.165 2696.895 1796.975 ;
        RECT 2696.905 1796.195 2698.275 1796.975 ;
        RECT 2698.285 1796.165 2703.795 1796.975 ;
        RECT 2703.805 1796.165 2709.315 1796.975 ;
        RECT 2709.325 1796.165 2714.835 1796.975 ;
        RECT 2714.845 1796.165 2720.355 1796.975 ;
        RECT 2721.745 1796.165 2727.255 1796.975 ;
        RECT 2727.265 1796.165 2732.775 1796.975 ;
        RECT 2732.785 1796.165 2734.155 1796.975 ;
        RECT 2695.525 1791.745 2696.895 1792.555 ;
        RECT 2696.905 1791.745 2698.275 1792.555 ;
        RECT 2698.285 1791.745 2701.955 1792.655 ;
        RECT 2701.965 1791.745 2707.475 1792.555 ;
        RECT 2708.865 1791.745 2714.375 1792.555 ;
        RECT 2714.385 1791.745 2719.895 1792.555 ;
        RECT 2719.905 1791.745 2725.415 1792.555 ;
        RECT 2725.425 1791.745 2730.935 1792.555 ;
        RECT 2730.945 1791.745 2732.775 1792.555 ;
        RECT 2732.785 1791.745 2734.155 1792.555 ;
        RECT 2695.665 1791.535 2695.835 1791.745 ;
        RECT 2697.045 1791.555 2697.215 1791.745 ;
        RECT 2522.700 1791.135 2522.870 1791.305 ;
        RECT 2695.525 1790.725 2696.895 1791.535 ;
        RECT 2697.965 1791.505 2698.135 1791.725 ;
        RECT 2701.640 1791.555 2701.810 1791.745 ;
        RECT 2702.105 1791.555 2702.275 1791.745 ;
        RECT 2703.485 1791.535 2703.655 1791.725 ;
        RECT 2703.945 1791.535 2704.115 1791.725 ;
        RECT 2707.635 1791.590 2707.795 1791.700 ;
        RECT 2709.005 1791.555 2709.175 1791.745 ;
        RECT 2709.465 1791.535 2709.635 1791.725 ;
        RECT 2714.525 1791.555 2714.695 1791.745 ;
        RECT 2714.985 1791.535 2715.155 1791.725 ;
        RECT 2720.045 1791.555 2720.215 1791.745 ;
        RECT 2720.515 1791.580 2720.675 1791.690 ;
        RECT 2721.885 1791.535 2722.055 1791.725 ;
        RECT 2725.565 1791.555 2725.735 1791.745 ;
        RECT 2727.405 1791.535 2727.575 1791.725 ;
        RECT 2731.085 1791.555 2731.255 1791.745 ;
        RECT 2733.845 1791.535 2734.015 1791.745 ;
        RECT 2700.090 1791.505 2701.035 1791.535 ;
        RECT 2697.965 1791.305 2701.035 1791.505 ;
        RECT 2697.825 1790.825 2701.035 1791.305 ;
        RECT 2697.825 1790.625 2698.755 1790.825 ;
        RECT 2700.090 1790.625 2701.035 1790.825 ;
        RECT 2701.275 1791.305 2703.655 1791.535 ;
        RECT 2701.275 1790.625 2703.665 1791.305 ;
        RECT 2703.805 1790.725 2709.315 1791.535 ;
        RECT 2709.325 1790.725 2714.835 1791.535 ;
        RECT 2714.845 1790.725 2720.355 1791.535 ;
        RECT 2721.745 1790.725 2727.255 1791.535 ;
        RECT 2727.265 1790.725 2732.775 1791.535 ;
        RECT 2732.785 1790.725 2734.155 1791.535 ;
        RECT 2695.525 1786.305 2696.895 1787.115 ;
        RECT 2696.905 1786.305 2698.275 1787.085 ;
        RECT 2698.745 1786.305 2700.095 1787.215 ;
        RECT 2700.125 1786.305 2705.635 1787.115 ;
        RECT 2705.645 1786.305 2708.395 1787.115 ;
        RECT 2708.865 1786.305 2714.375 1787.115 ;
        RECT 2714.385 1786.305 2719.895 1787.115 ;
        RECT 2719.905 1786.305 2725.415 1787.115 ;
        RECT 2725.425 1786.305 2730.935 1787.115 ;
        RECT 2730.945 1786.305 2732.775 1787.115 ;
        RECT 2732.785 1786.305 2734.155 1787.115 ;
        RECT 2695.665 1786.095 2695.835 1786.305 ;
        RECT 2697.045 1786.115 2697.215 1786.305 ;
        RECT 2698.420 1786.145 2698.540 1786.255 ;
        RECT 2699.810 1786.115 2699.980 1786.305 ;
        RECT 2700.265 1786.115 2700.435 1786.305 ;
        RECT 2700.450 1786.095 2700.620 1786.285 ;
        RECT 2701.185 1786.095 2701.355 1786.285 ;
        RECT 2705.785 1786.115 2705.955 1786.305 ;
        RECT 2706.705 1786.095 2706.875 1786.285 ;
        RECT 2709.005 1786.115 2709.175 1786.305 ;
        RECT 2712.225 1786.095 2712.395 1786.285 ;
        RECT 2714.525 1786.115 2714.695 1786.305 ;
        RECT 2717.745 1786.095 2717.915 1786.285 ;
        RECT 2720.045 1786.115 2720.215 1786.305 ;
        RECT 2721.885 1786.095 2722.055 1786.285 ;
        RECT 2725.565 1786.115 2725.735 1786.305 ;
        RECT 2727.405 1786.095 2727.575 1786.285 ;
        RECT 2731.085 1786.115 2731.255 1786.305 ;
        RECT 2733.845 1786.095 2734.015 1786.305 ;
        RECT 2522.700 1785.190 2522.870 1785.360 ;
        RECT 2695.525 1785.285 2696.895 1786.095 ;
        RECT 2697.135 1785.415 2701.035 1786.095 ;
        RECT 2700.105 1785.185 2701.035 1785.415 ;
        RECT 2701.045 1785.285 2706.555 1786.095 ;
        RECT 2706.565 1785.285 2712.075 1786.095 ;
        RECT 2712.085 1785.285 2717.595 1786.095 ;
        RECT 2717.605 1785.285 2721.275 1786.095 ;
        RECT 2721.745 1785.285 2727.255 1786.095 ;
        RECT 2727.265 1785.285 2732.775 1786.095 ;
        RECT 2732.785 1785.285 2734.155 1786.095 ;
        RECT 2371.875 1782.715 2372.045 1782.875 ;
        RECT 2387.135 1782.715 2387.305 1782.875 ;
        RECT 2402.395 1782.715 2402.565 1782.875 ;
        RECT 2417.655 1782.715 2417.825 1782.875 ;
        RECT 2432.915 1782.715 2433.085 1782.875 ;
        RECT 2695.525 1780.865 2696.895 1781.675 ;
        RECT 2696.905 1780.865 2698.275 1781.645 ;
        RECT 2698.285 1780.865 2703.795 1781.675 ;
        RECT 2703.805 1780.865 2707.475 1781.675 ;
        RECT 2708.865 1780.865 2714.375 1781.675 ;
        RECT 2714.385 1780.865 2719.895 1781.675 ;
        RECT 2719.905 1780.865 2725.415 1781.675 ;
        RECT 2725.425 1780.865 2730.935 1781.675 ;
        RECT 2730.945 1780.865 2732.775 1781.675 ;
        RECT 2732.785 1780.865 2734.155 1781.675 ;
        RECT 2695.665 1780.655 2695.835 1780.865 ;
        RECT 2697.045 1780.655 2697.215 1780.865 ;
        RECT 2698.425 1780.675 2698.595 1780.865 ;
        RECT 2702.565 1780.655 2702.735 1780.845 ;
        RECT 2703.945 1780.675 2704.115 1780.865 ;
        RECT 2707.635 1780.710 2707.795 1780.820 ;
        RECT 2708.085 1780.655 2708.255 1780.845 ;
        RECT 2709.005 1780.675 2709.175 1780.865 ;
        RECT 2713.605 1780.655 2713.775 1780.845 ;
        RECT 2714.525 1780.675 2714.695 1780.865 ;
        RECT 2719.125 1780.655 2719.295 1780.845 ;
        RECT 2720.045 1780.675 2720.215 1780.865 ;
        RECT 2720.960 1780.705 2721.080 1780.815 ;
        RECT 2721.885 1780.655 2722.055 1780.845 ;
        RECT 2725.565 1780.675 2725.735 1780.865 ;
        RECT 2727.405 1780.655 2727.575 1780.845 ;
        RECT 2731.085 1780.675 2731.255 1780.865 ;
        RECT 2733.845 1780.655 2734.015 1780.865 ;
        RECT 2695.525 1779.845 2696.895 1780.655 ;
        RECT 2696.905 1779.845 2702.415 1780.655 ;
        RECT 2702.425 1779.845 2707.935 1780.655 ;
        RECT 2707.945 1779.845 2713.455 1780.655 ;
        RECT 2713.465 1779.845 2718.975 1780.655 ;
        RECT 2718.985 1779.845 2720.815 1780.655 ;
        RECT 2721.745 1779.845 2727.255 1780.655 ;
        RECT 2727.265 1779.845 2732.775 1780.655 ;
        RECT 2732.785 1779.845 2734.155 1780.655 ;
        RECT 2522.700 1779.545 2522.870 1779.715 ;
        RECT 2695.525 1775.425 2696.895 1776.235 ;
        RECT 2696.905 1775.425 2698.275 1776.205 ;
        RECT 2698.285 1775.425 2703.795 1776.235 ;
        RECT 2703.805 1775.425 2707.475 1776.235 ;
        RECT 2708.865 1775.425 2714.375 1776.235 ;
        RECT 2714.385 1775.425 2719.895 1776.235 ;
        RECT 2719.905 1775.425 2725.415 1776.235 ;
        RECT 2725.425 1775.425 2730.935 1776.235 ;
        RECT 2730.945 1775.425 2732.775 1776.235 ;
        RECT 2732.785 1775.425 2734.155 1776.235 ;
        RECT 2695.665 1775.215 2695.835 1775.425 ;
        RECT 2697.045 1775.215 2697.215 1775.425 ;
        RECT 2698.425 1775.235 2698.595 1775.425 ;
        RECT 2702.565 1775.215 2702.735 1775.405 ;
        RECT 2703.945 1775.235 2704.115 1775.425 ;
        RECT 2707.635 1775.270 2707.795 1775.380 ;
        RECT 2708.085 1775.215 2708.255 1775.405 ;
        RECT 2709.005 1775.235 2709.175 1775.425 ;
        RECT 2713.605 1775.215 2713.775 1775.405 ;
        RECT 2714.525 1775.235 2714.695 1775.425 ;
        RECT 2719.125 1775.215 2719.295 1775.405 ;
        RECT 2720.045 1775.235 2720.215 1775.425 ;
        RECT 2720.960 1775.265 2721.080 1775.375 ;
        RECT 2721.885 1775.215 2722.055 1775.405 ;
        RECT 2725.565 1775.235 2725.735 1775.425 ;
        RECT 2727.405 1775.215 2727.575 1775.405 ;
        RECT 2731.085 1775.235 2731.255 1775.425 ;
        RECT 2733.845 1775.215 2734.015 1775.425 ;
        RECT 2695.525 1774.405 2696.895 1775.215 ;
        RECT 2696.905 1774.405 2702.415 1775.215 ;
        RECT 2702.425 1774.405 2707.935 1775.215 ;
        RECT 2707.945 1774.405 2713.455 1775.215 ;
        RECT 2713.465 1774.405 2718.975 1775.215 ;
        RECT 2718.985 1774.405 2720.815 1775.215 ;
        RECT 2721.745 1774.405 2727.255 1775.215 ;
        RECT 2727.265 1774.405 2732.775 1775.215 ;
        RECT 2732.785 1774.405 2734.155 1775.215 ;
        RECT 2695.525 1769.985 2696.895 1770.795 ;
        RECT 2696.905 1769.985 2698.275 1770.765 ;
        RECT 2698.285 1769.985 2699.655 1770.765 ;
        RECT 2699.665 1769.985 2705.175 1770.795 ;
        RECT 2705.185 1769.985 2707.935 1770.795 ;
        RECT 2708.865 1769.985 2714.375 1770.795 ;
        RECT 2714.385 1769.985 2719.895 1770.795 ;
        RECT 2719.905 1769.985 2721.275 1770.795 ;
        RECT 2721.745 1769.985 2727.255 1770.795 ;
        RECT 2727.265 1769.985 2732.775 1770.795 ;
        RECT 2732.785 1769.985 2734.155 1770.795 ;
        RECT 2695.665 1769.795 2695.835 1769.985 ;
        RECT 2697.045 1769.795 2697.215 1769.985 ;
        RECT 2698.425 1769.795 2698.595 1769.985 ;
        RECT 2699.805 1769.795 2699.975 1769.985 ;
        RECT 2705.325 1769.795 2705.495 1769.985 ;
        RECT 2708.080 1769.825 2708.200 1769.935 ;
        RECT 2709.005 1769.795 2709.175 1769.985 ;
        RECT 2714.525 1769.795 2714.695 1769.985 ;
        RECT 2720.045 1769.795 2720.215 1769.985 ;
        RECT 2721.885 1769.795 2722.055 1769.985 ;
        RECT 2727.405 1769.795 2727.575 1769.985 ;
        RECT 2733.845 1769.795 2734.015 1769.985 ;
        RECT 2522.700 1768.075 2522.870 1768.245 ;
        RECT 2364.680 1708.335 2365.410 1708.745 ;
        RECT 2367.320 1708.495 2367.490 1708.525 ;
        RECT 2370.540 1708.495 2370.710 1708.525 ;
        RECT 2367.320 1708.335 2367.900 1708.495 ;
        RECT 2370.540 1708.385 2371.170 1708.495 ;
        RECT 2370.540 1708.335 2370.850 1708.385 ;
        RECT 2364.680 1708.145 2370.850 1708.335 ;
        RECT 2381.265 1708.335 2381.995 1708.745 ;
        RECT 2383.905 1708.495 2384.075 1708.525 ;
        RECT 2387.125 1708.495 2387.295 1708.525 ;
        RECT 2383.905 1708.335 2384.485 1708.495 ;
        RECT 2387.125 1708.385 2387.755 1708.495 ;
        RECT 2387.125 1708.335 2387.435 1708.385 ;
        RECT 2381.265 1708.145 2387.435 1708.335 ;
        RECT 2397.850 1708.340 2398.580 1708.750 ;
        RECT 2400.490 1708.500 2400.660 1708.530 ;
        RECT 2403.710 1708.500 2403.880 1708.530 ;
        RECT 2400.490 1708.340 2401.070 1708.500 ;
        RECT 2403.710 1708.390 2404.340 1708.500 ;
        RECT 2403.710 1708.340 2404.020 1708.390 ;
        RECT 2397.850 1708.150 2404.020 1708.340 ;
        RECT 2414.435 1708.345 2415.165 1708.755 ;
        RECT 2417.075 1708.505 2417.245 1708.535 ;
        RECT 2420.295 1708.505 2420.465 1708.535 ;
        RECT 2417.075 1708.345 2417.655 1708.505 ;
        RECT 2420.295 1708.395 2420.925 1708.505 ;
        RECT 2420.295 1708.345 2420.605 1708.395 ;
        RECT 2414.435 1708.155 2420.605 1708.345 ;
        RECT 2431.015 1708.345 2431.745 1708.755 ;
        RECT 2433.655 1708.505 2433.825 1708.535 ;
        RECT 2436.875 1708.505 2437.045 1708.535 ;
        RECT 2433.655 1708.345 2434.235 1708.505 ;
        RECT 2436.875 1708.395 2437.505 1708.505 ;
        RECT 2436.875 1708.345 2437.185 1708.395 ;
        RECT 2431.015 1708.155 2437.185 1708.345 ;
        RECT 2365.540 1707.515 2370.850 1708.145 ;
        RECT 2365.540 1707.425 2366.490 1707.515 ;
        RECT 2368.100 1707.425 2370.850 1707.515 ;
        RECT 2382.125 1707.515 2387.435 1708.145 ;
        RECT 2382.125 1707.425 2383.075 1707.515 ;
        RECT 2384.685 1707.425 2387.435 1707.515 ;
        RECT 2398.710 1707.520 2404.020 1708.150 ;
        RECT 2398.710 1707.430 2399.660 1707.520 ;
        RECT 2401.270 1707.430 2404.020 1707.520 ;
        RECT 2415.295 1707.525 2420.605 1708.155 ;
        RECT 2415.295 1707.435 2416.245 1707.525 ;
        RECT 2417.855 1707.435 2420.605 1707.525 ;
        RECT 2431.875 1707.525 2437.185 1708.155 ;
        RECT 2431.875 1707.435 2432.825 1707.525 ;
        RECT 2434.435 1707.435 2437.185 1707.525 ;
        RECT 2364.580 1703.815 2365.810 1704.015 ;
        RECT 2367.140 1703.815 2368.090 1704.015 ;
        RECT 2364.580 1703.790 2368.090 1703.815 ;
        RECT 2369.470 1703.790 2371.750 1704.015 ;
        RECT 2364.580 1703.305 2371.750 1703.790 ;
        RECT 2381.165 1703.815 2382.395 1704.015 ;
        RECT 2383.725 1703.815 2384.675 1704.015 ;
        RECT 2381.165 1703.790 2384.675 1703.815 ;
        RECT 2386.055 1703.790 2388.335 1704.015 ;
        RECT 2381.165 1703.305 2388.335 1703.790 ;
        RECT 2397.750 1703.820 2398.980 1704.020 ;
        RECT 2400.310 1703.820 2401.260 1704.020 ;
        RECT 2397.750 1703.795 2401.260 1703.820 ;
        RECT 2402.640 1703.795 2404.920 1704.020 ;
        RECT 2397.750 1703.310 2404.920 1703.795 ;
        RECT 2414.335 1703.825 2415.565 1704.025 ;
        RECT 2416.895 1703.825 2417.845 1704.025 ;
        RECT 2414.335 1703.800 2417.845 1703.825 ;
        RECT 2419.225 1703.800 2421.505 1704.025 ;
        RECT 2414.335 1703.315 2421.505 1703.800 ;
        RECT 2430.915 1703.825 2432.145 1704.025 ;
        RECT 2433.475 1703.825 2434.425 1704.025 ;
        RECT 2430.915 1703.800 2434.425 1703.825 ;
        RECT 2435.805 1703.800 2438.085 1704.025 ;
        RECT 2430.915 1703.315 2438.085 1703.800 ;
        RECT 2364.520 1703.135 2371.750 1703.305 ;
        RECT 2364.520 1702.705 2365.110 1703.135 ;
        RECT 2367.160 1703.110 2371.750 1703.135 ;
        RECT 2381.105 1703.135 2388.335 1703.305 ;
        RECT 2368.240 1702.925 2368.410 1703.105 ;
        RECT 2370.550 1703.095 2370.720 1703.105 ;
        RECT 2370.540 1703.085 2370.720 1703.095 ;
        RECT 2370.550 1702.925 2370.720 1703.085 ;
        RECT 2381.105 1702.705 2381.695 1703.135 ;
        RECT 2383.745 1703.110 2388.335 1703.135 ;
        RECT 2397.690 1703.140 2404.920 1703.310 ;
        RECT 2384.825 1702.925 2384.995 1703.105 ;
        RECT 2387.135 1703.095 2387.305 1703.105 ;
        RECT 2387.125 1703.085 2387.305 1703.095 ;
        RECT 2387.135 1702.925 2387.305 1703.085 ;
        RECT 2397.690 1702.710 2398.280 1703.140 ;
        RECT 2400.330 1703.115 2404.920 1703.140 ;
        RECT 2414.275 1703.145 2421.505 1703.315 ;
        RECT 2401.410 1702.930 2401.580 1703.110 ;
        RECT 2403.720 1703.100 2403.890 1703.110 ;
        RECT 2403.710 1703.090 2403.890 1703.100 ;
        RECT 2403.720 1702.930 2403.890 1703.090 ;
        RECT 2414.275 1702.715 2414.865 1703.145 ;
        RECT 2416.915 1703.120 2421.505 1703.145 ;
        RECT 2430.855 1703.145 2438.085 1703.315 ;
        RECT 2417.995 1702.935 2418.165 1703.115 ;
        RECT 2420.305 1703.105 2420.475 1703.115 ;
        RECT 2420.295 1703.095 2420.475 1703.105 ;
        RECT 2420.305 1702.935 2420.475 1703.095 ;
        RECT 2430.855 1702.715 2431.445 1703.145 ;
        RECT 2433.495 1703.120 2438.085 1703.145 ;
        RECT 2434.575 1702.935 2434.745 1703.115 ;
        RECT 2436.885 1703.105 2437.055 1703.115 ;
        RECT 2436.875 1703.095 2437.055 1703.105 ;
        RECT 2436.885 1702.935 2437.055 1703.095 ;
        RECT 2695.665 1676.815 2695.835 1677.005 ;
        RECT 2697.045 1676.815 2697.215 1677.005 ;
        RECT 2699.805 1676.815 2699.975 1677.005 ;
        RECT 2701.185 1676.815 2701.355 1677.005 ;
        RECT 2701.645 1676.815 2701.815 1677.005 ;
        RECT 2707.165 1676.815 2707.335 1677.005 ;
        RECT 2709.005 1676.815 2709.175 1677.005 ;
        RECT 2710.845 1676.815 2711.015 1677.005 ;
        RECT 2716.365 1676.815 2716.535 1677.005 ;
        RECT 2720.045 1676.815 2720.215 1677.005 ;
        RECT 2723.265 1676.815 2723.435 1677.005 ;
        RECT 2723.725 1676.815 2723.895 1677.005 ;
        RECT 2729.245 1676.815 2729.415 1677.005 ;
        RECT 2731.080 1676.865 2731.200 1676.975 ;
        RECT 2732.455 1676.815 2732.625 1677.005 ;
        RECT 2733.845 1676.815 2734.015 1677.005 ;
        RECT 2695.525 1676.005 2696.895 1676.815 ;
        RECT 2696.905 1676.135 2698.735 1676.815 ;
        RECT 2698.745 1676.035 2700.115 1676.815 ;
        RECT 2700.125 1676.035 2701.495 1676.815 ;
        RECT 2701.505 1676.005 2707.015 1676.815 ;
        RECT 2707.025 1676.005 2708.395 1676.815 ;
        RECT 2708.865 1676.135 2710.695 1676.815 ;
        RECT 2709.350 1675.905 2710.695 1676.135 ;
        RECT 2710.705 1676.005 2716.215 1676.815 ;
        RECT 2716.225 1676.005 2719.895 1676.815 ;
        RECT 2719.905 1676.005 2721.275 1676.815 ;
        RECT 2721.745 1676.135 2723.575 1676.815 ;
        RECT 2723.585 1676.005 2729.095 1676.815 ;
        RECT 2729.105 1676.005 2730.935 1676.815 ;
        RECT 2731.405 1676.035 2732.775 1676.815 ;
        RECT 2732.785 1676.005 2734.155 1676.815 ;
        RECT 2695.525 1671.585 2696.895 1672.395 ;
        RECT 2696.905 1671.585 2698.275 1672.365 ;
        RECT 2698.285 1671.585 2703.795 1672.395 ;
        RECT 2703.805 1671.585 2707.475 1672.395 ;
        RECT 2708.865 1671.585 2714.375 1672.395 ;
        RECT 2714.385 1671.585 2719.895 1672.395 ;
        RECT 2719.905 1671.585 2725.415 1672.395 ;
        RECT 2725.425 1671.585 2730.935 1672.395 ;
        RECT 2730.945 1671.585 2732.775 1672.395 ;
        RECT 2732.785 1671.585 2734.155 1672.395 ;
        RECT 2695.665 1671.375 2695.835 1671.585 ;
        RECT 2697.045 1671.375 2697.215 1671.585 ;
        RECT 2698.425 1671.395 2698.595 1671.585 ;
        RECT 2702.565 1671.375 2702.735 1671.565 ;
        RECT 2703.945 1671.395 2704.115 1671.585 ;
        RECT 2707.635 1671.430 2707.795 1671.540 ;
        RECT 2708.085 1671.375 2708.255 1671.565 ;
        RECT 2709.005 1671.395 2709.175 1671.585 ;
        RECT 2713.605 1671.375 2713.775 1671.565 ;
        RECT 2714.525 1671.395 2714.695 1671.585 ;
        RECT 2719.125 1671.375 2719.295 1671.565 ;
        RECT 2720.045 1671.395 2720.215 1671.585 ;
        RECT 2720.960 1671.425 2721.080 1671.535 ;
        RECT 2721.885 1671.375 2722.055 1671.565 ;
        RECT 2725.565 1671.395 2725.735 1671.585 ;
        RECT 2727.405 1671.375 2727.575 1671.565 ;
        RECT 2731.085 1671.395 2731.255 1671.585 ;
        RECT 2733.845 1671.375 2734.015 1671.585 ;
        RECT 2695.525 1670.565 2696.895 1671.375 ;
        RECT 2696.905 1670.565 2702.415 1671.375 ;
        RECT 2702.425 1670.565 2707.935 1671.375 ;
        RECT 2707.945 1670.565 2713.455 1671.375 ;
        RECT 2713.465 1670.565 2718.975 1671.375 ;
        RECT 2718.985 1670.565 2720.815 1671.375 ;
        RECT 2721.745 1670.565 2727.255 1671.375 ;
        RECT 2727.265 1670.565 2732.775 1671.375 ;
        RECT 2732.785 1670.565 2734.155 1671.375 ;
        RECT 2695.525 1666.145 2696.895 1666.955 ;
        RECT 2696.905 1666.145 2702.415 1666.955 ;
        RECT 2702.425 1666.145 2707.935 1666.955 ;
        RECT 2708.865 1666.145 2714.375 1666.955 ;
        RECT 2714.385 1666.145 2719.895 1666.955 ;
        RECT 2719.905 1666.145 2725.415 1666.955 ;
        RECT 2725.425 1666.145 2730.935 1666.955 ;
        RECT 2730.945 1666.145 2732.775 1666.955 ;
        RECT 2732.785 1666.145 2734.155 1666.955 ;
        RECT 2695.665 1665.935 2695.835 1666.145 ;
        RECT 2697.045 1665.935 2697.215 1666.145 ;
        RECT 2698.425 1665.935 2698.595 1666.125 ;
        RECT 2702.565 1665.955 2702.735 1666.145 ;
        RECT 2703.945 1665.935 2704.115 1666.125 ;
        RECT 2708.080 1665.985 2708.200 1666.095 ;
        RECT 2709.005 1665.955 2709.175 1666.145 ;
        RECT 2709.465 1665.935 2709.635 1666.125 ;
        RECT 2714.525 1665.955 2714.695 1666.145 ;
        RECT 2714.985 1665.935 2715.155 1666.125 ;
        RECT 2720.045 1665.955 2720.215 1666.145 ;
        RECT 2720.515 1665.980 2720.675 1666.090 ;
        RECT 2721.885 1665.935 2722.055 1666.125 ;
        RECT 2725.565 1665.955 2725.735 1666.145 ;
        RECT 2727.405 1665.935 2727.575 1666.125 ;
        RECT 2731.085 1665.955 2731.255 1666.145 ;
        RECT 2733.845 1665.935 2734.015 1666.145 ;
        RECT 2695.525 1665.125 2696.895 1665.935 ;
        RECT 2696.905 1665.155 2698.275 1665.935 ;
        RECT 2698.285 1665.125 2703.795 1665.935 ;
        RECT 2703.805 1665.125 2709.315 1665.935 ;
        RECT 2709.325 1665.125 2714.835 1665.935 ;
        RECT 2714.845 1665.125 2720.355 1665.935 ;
        RECT 2721.745 1665.125 2727.255 1665.935 ;
        RECT 2727.265 1665.125 2732.775 1665.935 ;
        RECT 2732.785 1665.125 2734.155 1665.935 ;
        RECT 2695.525 1660.705 2696.895 1661.515 ;
        RECT 2696.905 1660.705 2702.415 1661.515 ;
        RECT 2702.425 1660.705 2707.935 1661.515 ;
        RECT 2708.865 1660.705 2714.375 1661.515 ;
        RECT 2714.385 1660.705 2719.895 1661.515 ;
        RECT 2719.905 1660.705 2725.415 1661.515 ;
        RECT 2725.425 1660.705 2730.935 1661.515 ;
        RECT 2730.945 1660.705 2732.775 1661.515 ;
        RECT 2732.785 1660.705 2734.155 1661.515 ;
        RECT 2695.665 1660.495 2695.835 1660.705 ;
        RECT 2697.045 1660.495 2697.215 1660.705 ;
        RECT 2702.565 1660.515 2702.735 1660.705 ;
        RECT 2706.705 1660.495 2706.875 1660.685 ;
        RECT 2708.080 1660.545 2708.200 1660.655 ;
        RECT 2709.005 1660.515 2709.175 1660.705 ;
        RECT 2712.225 1660.495 2712.395 1660.685 ;
        RECT 2714.525 1660.515 2714.695 1660.705 ;
        RECT 2717.745 1660.495 2717.915 1660.685 ;
        RECT 2720.045 1660.515 2720.215 1660.705 ;
        RECT 2721.885 1660.495 2722.055 1660.685 ;
        RECT 2725.565 1660.515 2725.735 1660.705 ;
        RECT 2727.405 1660.495 2727.575 1660.685 ;
        RECT 2731.085 1660.515 2731.255 1660.705 ;
        RECT 2733.845 1660.495 2734.015 1660.705 ;
        RECT 2695.525 1659.685 2696.895 1660.495 ;
        RECT 2696.905 1660.325 2698.665 1660.495 ;
        RECT 2696.905 1660.280 2699.160 1660.325 ;
        RECT 2696.905 1660.245 2700.100 1660.280 ;
        RECT 2701.460 1660.245 2706.555 1660.495 ;
        RECT 2696.905 1659.815 2706.555 1660.245 ;
        RECT 2698.230 1659.645 2701.460 1659.815 ;
        RECT 2699.170 1659.600 2701.460 1659.645 ;
        RECT 2700.110 1659.565 2701.460 1659.600 ;
        RECT 2704.535 1659.585 2706.555 1659.815 ;
        RECT 2706.565 1659.685 2712.075 1660.495 ;
        RECT 2712.085 1659.685 2717.595 1660.495 ;
        RECT 2717.605 1659.685 2721.275 1660.495 ;
        RECT 2721.745 1659.685 2727.255 1660.495 ;
        RECT 2727.265 1659.685 2732.775 1660.495 ;
        RECT 2732.785 1659.685 2734.155 1660.495 ;
        RECT 2704.535 1659.565 2705.455 1659.585 ;
        RECT 2695.525 1655.265 2696.895 1656.075 ;
        RECT 2696.905 1655.265 2698.275 1656.045 ;
        RECT 2698.285 1655.265 2703.795 1656.075 ;
        RECT 2703.805 1655.265 2707.475 1656.075 ;
        RECT 2708.865 1655.265 2714.375 1656.075 ;
        RECT 2714.385 1655.265 2719.895 1656.075 ;
        RECT 2719.905 1655.265 2725.415 1656.075 ;
        RECT 2725.425 1655.265 2730.935 1656.075 ;
        RECT 2730.945 1655.265 2732.775 1656.075 ;
        RECT 2732.785 1655.265 2734.155 1656.075 ;
        RECT 2695.665 1655.055 2695.835 1655.265 ;
        RECT 2697.045 1655.055 2697.215 1655.265 ;
        RECT 2698.425 1655.075 2698.595 1655.265 ;
        RECT 2703.945 1655.075 2704.115 1655.265 ;
        RECT 2706.705 1655.055 2706.875 1655.245 ;
        RECT 2707.635 1655.110 2707.795 1655.220 ;
        RECT 2709.005 1655.075 2709.175 1655.265 ;
        RECT 2712.225 1655.055 2712.395 1655.245 ;
        RECT 2714.525 1655.075 2714.695 1655.265 ;
        RECT 2717.745 1655.055 2717.915 1655.245 ;
        RECT 2720.045 1655.075 2720.215 1655.265 ;
        RECT 2721.885 1655.055 2722.055 1655.245 ;
        RECT 2725.565 1655.075 2725.735 1655.265 ;
        RECT 2727.405 1655.055 2727.575 1655.245 ;
        RECT 2731.085 1655.075 2731.255 1655.265 ;
        RECT 2733.845 1655.055 2734.015 1655.265 ;
        RECT 2695.525 1654.245 2696.895 1655.055 ;
        RECT 2696.905 1654.885 2698.665 1655.055 ;
        RECT 2696.905 1654.840 2699.160 1654.885 ;
        RECT 2696.905 1654.805 2700.100 1654.840 ;
        RECT 2701.460 1654.805 2706.555 1655.055 ;
        RECT 2696.905 1654.375 2706.555 1654.805 ;
        RECT 2698.230 1654.205 2701.460 1654.375 ;
        RECT 2699.170 1654.160 2701.460 1654.205 ;
        RECT 2700.110 1654.125 2701.460 1654.160 ;
        RECT 2704.535 1654.145 2706.555 1654.375 ;
        RECT 2706.565 1654.245 2712.075 1655.055 ;
        RECT 2712.085 1654.245 2717.595 1655.055 ;
        RECT 2717.605 1654.245 2721.275 1655.055 ;
        RECT 2721.745 1654.245 2727.255 1655.055 ;
        RECT 2727.265 1654.245 2732.775 1655.055 ;
        RECT 2732.785 1654.245 2734.155 1655.055 ;
        RECT 2704.535 1654.125 2705.455 1654.145 ;
        RECT 2695.525 1649.825 2696.895 1650.635 ;
        RECT 2696.905 1649.825 2698.275 1650.605 ;
        RECT 2698.285 1649.825 2701.035 1650.635 ;
        RECT 2701.505 1650.505 2702.435 1650.735 ;
        RECT 2701.505 1649.825 2705.405 1650.505 ;
        RECT 2705.645 1649.825 2708.395 1650.635 ;
        RECT 2708.865 1649.825 2714.375 1650.635 ;
        RECT 2714.385 1649.825 2719.895 1650.635 ;
        RECT 2719.905 1649.825 2725.415 1650.635 ;
        RECT 2725.425 1649.825 2730.935 1650.635 ;
        RECT 2730.945 1649.825 2732.775 1650.635 ;
        RECT 2732.785 1649.825 2734.155 1650.635 ;
        RECT 2695.665 1649.615 2695.835 1649.825 ;
        RECT 2697.045 1649.615 2697.215 1649.825 ;
        RECT 2698.425 1649.635 2698.595 1649.825 ;
        RECT 2701.180 1649.665 2701.300 1649.775 ;
        RECT 2701.920 1649.635 2702.090 1649.825 ;
        RECT 2702.565 1649.615 2702.735 1649.805 ;
        RECT 2705.785 1649.635 2705.955 1649.825 ;
        RECT 2708.085 1649.615 2708.255 1649.805 ;
        RECT 2709.005 1649.635 2709.175 1649.825 ;
        RECT 2713.605 1649.615 2713.775 1649.805 ;
        RECT 2714.525 1649.635 2714.695 1649.825 ;
        RECT 2719.125 1649.615 2719.295 1649.805 ;
        RECT 2720.045 1649.635 2720.215 1649.825 ;
        RECT 2720.960 1649.665 2721.080 1649.775 ;
        RECT 2721.885 1649.615 2722.055 1649.805 ;
        RECT 2725.565 1649.635 2725.735 1649.825 ;
        RECT 2727.405 1649.615 2727.575 1649.805 ;
        RECT 2731.085 1649.635 2731.255 1649.825 ;
        RECT 2733.845 1649.615 2734.015 1649.825 ;
        RECT 2695.525 1648.805 2696.895 1649.615 ;
        RECT 2696.905 1648.805 2702.415 1649.615 ;
        RECT 2702.425 1648.805 2707.935 1649.615 ;
        RECT 2707.945 1648.805 2713.455 1649.615 ;
        RECT 2713.465 1648.805 2718.975 1649.615 ;
        RECT 2718.985 1648.805 2720.815 1649.615 ;
        RECT 2721.745 1648.805 2727.255 1649.615 ;
        RECT 2727.265 1648.805 2732.775 1649.615 ;
        RECT 2732.785 1648.805 2734.155 1649.615 ;
        RECT 2695.525 1644.385 2696.895 1645.195 ;
        RECT 2696.905 1644.385 2698.275 1645.165 ;
        RECT 2698.285 1644.385 2703.795 1645.195 ;
        RECT 2703.805 1644.385 2707.475 1645.195 ;
        RECT 2708.865 1644.385 2714.375 1645.195 ;
        RECT 2714.385 1644.385 2719.895 1645.195 ;
        RECT 2719.905 1644.385 2725.415 1645.195 ;
        RECT 2725.425 1644.385 2730.935 1645.195 ;
        RECT 2730.945 1644.385 2732.775 1645.195 ;
        RECT 2732.785 1644.385 2734.155 1645.195 ;
        RECT 2695.665 1644.175 2695.835 1644.385 ;
        RECT 2697.045 1644.175 2697.215 1644.385 ;
        RECT 2698.425 1644.195 2698.595 1644.385 ;
        RECT 2702.565 1644.175 2702.735 1644.365 ;
        RECT 2703.945 1644.195 2704.115 1644.385 ;
        RECT 2707.635 1644.230 2707.795 1644.340 ;
        RECT 2708.085 1644.175 2708.255 1644.365 ;
        RECT 2709.005 1644.195 2709.175 1644.385 ;
        RECT 2713.605 1644.175 2713.775 1644.365 ;
        RECT 2714.525 1644.195 2714.695 1644.385 ;
        RECT 2719.125 1644.175 2719.295 1644.365 ;
        RECT 2720.045 1644.195 2720.215 1644.385 ;
        RECT 2720.960 1644.225 2721.080 1644.335 ;
        RECT 2721.885 1644.175 2722.055 1644.365 ;
        RECT 2725.565 1644.195 2725.735 1644.385 ;
        RECT 2727.405 1644.175 2727.575 1644.365 ;
        RECT 2731.085 1644.195 2731.255 1644.385 ;
        RECT 2733.845 1644.175 2734.015 1644.385 ;
        RECT 2695.525 1643.365 2696.895 1644.175 ;
        RECT 2696.905 1643.365 2702.415 1644.175 ;
        RECT 2702.425 1643.365 2707.935 1644.175 ;
        RECT 2707.945 1643.365 2713.455 1644.175 ;
        RECT 2713.465 1643.365 2718.975 1644.175 ;
        RECT 2718.985 1643.365 2720.815 1644.175 ;
        RECT 2721.745 1643.365 2727.255 1644.175 ;
        RECT 2727.265 1643.365 2732.775 1644.175 ;
        RECT 2732.785 1643.365 2734.155 1644.175 ;
        RECT 2695.525 1638.945 2696.895 1639.755 ;
        RECT 2696.905 1638.945 2700.575 1639.755 ;
        RECT 2701.505 1638.945 2702.855 1639.855 ;
        RECT 2702.885 1638.945 2708.395 1639.755 ;
        RECT 2708.865 1638.945 2714.375 1639.755 ;
        RECT 2714.385 1638.945 2719.895 1639.755 ;
        RECT 2719.905 1638.945 2725.415 1639.755 ;
        RECT 2725.425 1638.945 2730.935 1639.755 ;
        RECT 2730.945 1638.945 2732.775 1639.755 ;
        RECT 2732.785 1638.945 2734.155 1639.755 ;
        RECT 2695.665 1638.735 2695.835 1638.945 ;
        RECT 2697.045 1638.735 2697.215 1638.945 ;
        RECT 2698.425 1638.735 2698.595 1638.925 ;
        RECT 2700.735 1638.790 2700.895 1638.900 ;
        RECT 2701.650 1638.755 2701.820 1638.945 ;
        RECT 2703.025 1638.755 2703.195 1638.945 ;
        RECT 2704.865 1638.735 2705.035 1638.925 ;
        RECT 2705.325 1638.735 2705.495 1638.925 ;
        RECT 2709.005 1638.755 2709.175 1638.945 ;
        RECT 2710.845 1638.735 2711.015 1638.925 ;
        RECT 2714.525 1638.755 2714.695 1638.945 ;
        RECT 2716.365 1638.735 2716.535 1638.925 ;
        RECT 2720.045 1638.735 2720.215 1638.945 ;
        RECT 2721.885 1638.735 2722.055 1638.925 ;
        RECT 2725.565 1638.755 2725.735 1638.945 ;
        RECT 2727.405 1638.735 2727.575 1638.925 ;
        RECT 2731.085 1638.755 2731.255 1638.945 ;
        RECT 2733.845 1638.735 2734.015 1638.945 ;
        RECT 2695.525 1637.925 2696.895 1638.735 ;
        RECT 2696.905 1637.955 2698.275 1638.735 ;
        RECT 2698.285 1637.925 2701.955 1638.735 ;
        RECT 2701.965 1637.825 2705.175 1638.735 ;
        RECT 2705.185 1637.925 2710.695 1638.735 ;
        RECT 2710.705 1637.925 2716.215 1638.735 ;
        RECT 2716.225 1637.925 2719.895 1638.735 ;
        RECT 2719.905 1637.925 2721.275 1638.735 ;
        RECT 2721.745 1637.925 2727.255 1638.735 ;
        RECT 2727.265 1637.925 2732.775 1638.735 ;
        RECT 2732.785 1637.925 2734.155 1638.735 ;
        RECT 2695.525 1633.505 2696.895 1634.315 ;
        RECT 2696.905 1633.505 2702.415 1634.315 ;
        RECT 2702.425 1633.505 2707.935 1634.315 ;
        RECT 2708.865 1633.505 2714.375 1634.315 ;
        RECT 2714.385 1633.505 2719.895 1634.315 ;
        RECT 2719.905 1633.505 2725.415 1634.315 ;
        RECT 2725.425 1633.505 2732.775 1634.415 ;
        RECT 2732.785 1633.505 2734.155 1634.315 ;
        RECT 2695.665 1633.295 2695.835 1633.505 ;
        RECT 2697.045 1633.295 2697.215 1633.505 ;
        RECT 2698.425 1633.295 2698.595 1633.485 ;
        RECT 2702.565 1633.315 2702.735 1633.505 ;
        RECT 2703.945 1633.295 2704.115 1633.485 ;
        RECT 2708.080 1633.345 2708.200 1633.455 ;
        RECT 2709.005 1633.315 2709.175 1633.505 ;
        RECT 2709.465 1633.295 2709.635 1633.485 ;
        RECT 2714.525 1633.315 2714.695 1633.505 ;
        RECT 2714.985 1633.295 2715.155 1633.485 ;
        RECT 2720.045 1633.315 2720.215 1633.505 ;
        RECT 2720.515 1633.340 2720.675 1633.450 ;
        RECT 2721.885 1633.295 2722.055 1633.485 ;
        RECT 2725.990 1633.315 2726.160 1633.505 ;
        RECT 2727.405 1633.295 2727.575 1633.485 ;
        RECT 2733.845 1633.295 2734.015 1633.505 ;
        RECT 2695.525 1632.485 2696.895 1633.295 ;
        RECT 2696.905 1632.515 2698.275 1633.295 ;
        RECT 2698.285 1632.485 2703.795 1633.295 ;
        RECT 2703.805 1632.485 2709.315 1633.295 ;
        RECT 2709.325 1632.485 2714.835 1633.295 ;
        RECT 2714.845 1632.485 2720.355 1633.295 ;
        RECT 2721.745 1632.485 2727.255 1633.295 ;
        RECT 2727.265 1632.485 2732.775 1633.295 ;
        RECT 2732.785 1632.485 2734.155 1633.295 ;
        RECT 2695.525 1628.065 2696.895 1628.875 ;
        RECT 2696.905 1628.065 2702.415 1628.875 ;
        RECT 2702.425 1628.065 2707.935 1628.875 ;
        RECT 2708.865 1628.065 2714.375 1628.875 ;
        RECT 2714.385 1628.065 2719.895 1628.875 ;
        RECT 2719.905 1628.065 2725.415 1628.875 ;
        RECT 2725.425 1628.065 2730.935 1628.875 ;
        RECT 2730.945 1628.065 2732.775 1628.875 ;
        RECT 2732.785 1628.065 2734.155 1628.875 ;
        RECT 2695.665 1627.855 2695.835 1628.065 ;
        RECT 2697.045 1627.875 2697.215 1628.065 ;
        RECT 2699.345 1627.875 2699.515 1628.045 ;
        RECT 2699.345 1627.855 2699.475 1627.875 ;
        RECT 2699.805 1627.855 2699.975 1628.045 ;
        RECT 2702.565 1627.875 2702.735 1628.065 ;
        RECT 2705.325 1627.855 2705.495 1628.045 ;
        RECT 2708.080 1627.905 2708.200 1628.015 ;
        RECT 2709.005 1627.875 2709.175 1628.065 ;
        RECT 2710.845 1627.855 2711.015 1628.045 ;
        RECT 2714.525 1627.875 2714.695 1628.065 ;
        RECT 2716.365 1627.855 2716.535 1628.045 ;
        RECT 2720.045 1627.855 2720.215 1628.065 ;
        RECT 2721.885 1627.855 2722.055 1628.045 ;
        RECT 2725.565 1627.875 2725.735 1628.065 ;
        RECT 2727.405 1627.855 2727.575 1628.045 ;
        RECT 2731.085 1627.875 2731.255 1628.065 ;
        RECT 2733.845 1627.855 2734.015 1628.065 ;
        RECT 2695.525 1627.045 2696.895 1627.855 ;
        RECT 2697.625 1627.625 2699.475 1627.855 ;
        RECT 2697.140 1626.945 2699.475 1627.625 ;
        RECT 2699.665 1627.045 2705.175 1627.855 ;
        RECT 2705.185 1627.045 2710.695 1627.855 ;
        RECT 2710.705 1627.045 2716.215 1627.855 ;
        RECT 2716.225 1627.045 2719.895 1627.855 ;
        RECT 2719.905 1627.045 2721.275 1627.855 ;
        RECT 2721.745 1627.045 2727.255 1627.855 ;
        RECT 2727.265 1627.045 2732.775 1627.855 ;
        RECT 2732.785 1627.045 2734.155 1627.855 ;
        RECT 2883.065 1625.620 2883.235 1625.790 ;
        RECT 2522.700 1623.510 2522.870 1623.680 ;
        RECT 2695.525 1622.625 2696.895 1623.435 ;
        RECT 2696.905 1622.625 2698.275 1623.405 ;
        RECT 2698.285 1622.625 2703.795 1623.435 ;
        RECT 2703.805 1622.625 2707.475 1623.435 ;
        RECT 2708.865 1622.625 2714.375 1623.435 ;
        RECT 2714.385 1622.625 2719.895 1623.435 ;
        RECT 2719.905 1622.625 2725.415 1623.435 ;
        RECT 2725.425 1622.625 2730.935 1623.435 ;
        RECT 2730.945 1622.625 2732.775 1623.435 ;
        RECT 2732.785 1622.625 2734.155 1623.435 ;
        RECT 2695.665 1622.415 2695.835 1622.625 ;
        RECT 2697.045 1622.435 2697.215 1622.625 ;
        RECT 2698.425 1622.435 2698.595 1622.625 ;
        RECT 2700.450 1622.415 2700.620 1622.605 ;
        RECT 2702.575 1622.415 2702.745 1622.585 ;
        RECT 2703.945 1622.435 2704.115 1622.625 ;
        RECT 2704.405 1622.415 2704.575 1622.605 ;
        RECT 2704.865 1622.415 2705.035 1622.605 ;
        RECT 2707.635 1622.470 2707.795 1622.580 ;
        RECT 2709.005 1622.435 2709.175 1622.625 ;
        RECT 2710.385 1622.415 2710.555 1622.605 ;
        RECT 2714.525 1622.435 2714.695 1622.625 ;
        RECT 2715.905 1622.415 2716.075 1622.605 ;
        RECT 2720.045 1622.435 2720.215 1622.625 ;
        RECT 2721.885 1622.415 2722.055 1622.605 ;
        RECT 2725.565 1622.435 2725.735 1622.625 ;
        RECT 2727.405 1622.415 2727.575 1622.605 ;
        RECT 2731.085 1622.435 2731.255 1622.625 ;
        RECT 2733.845 1622.415 2734.015 1622.625 ;
        RECT 2695.525 1621.605 2696.895 1622.415 ;
        RECT 2697.135 1621.735 2701.035 1622.415 ;
        RECT 2700.105 1621.505 2701.035 1621.735 ;
        RECT 2701.045 1621.505 2704.695 1622.415 ;
        RECT 2704.725 1621.605 2710.235 1622.415 ;
        RECT 2710.245 1621.605 2715.755 1622.415 ;
        RECT 2715.765 1621.605 2721.275 1622.415 ;
        RECT 2721.745 1621.605 2727.255 1622.415 ;
        RECT 2727.265 1621.605 2732.775 1622.415 ;
        RECT 2732.785 1621.605 2734.155 1622.415 ;
        RECT 2522.700 1617.095 2522.870 1617.265 ;
        RECT 2695.525 1617.185 2696.895 1617.995 ;
        RECT 2696.905 1617.895 2697.835 1618.095 ;
        RECT 2699.165 1617.895 2700.115 1618.095 ;
        RECT 2696.905 1617.415 2700.115 1617.895 ;
        RECT 2697.050 1617.215 2700.115 1617.415 ;
        RECT 2695.665 1616.975 2695.835 1617.185 ;
        RECT 2697.050 1617.165 2697.220 1617.215 ;
        RECT 2699.180 1617.185 2700.115 1617.215 ;
        RECT 2700.125 1617.185 2705.635 1617.995 ;
        RECT 2705.645 1617.185 2708.395 1617.995 ;
        RECT 2708.865 1617.185 2714.375 1617.995 ;
        RECT 2714.385 1617.185 2719.895 1617.995 ;
        RECT 2719.905 1617.185 2725.415 1617.995 ;
        RECT 2725.425 1617.185 2730.935 1617.995 ;
        RECT 2730.945 1617.185 2732.775 1617.995 ;
        RECT 2732.785 1617.185 2734.155 1617.995 ;
        RECT 2697.045 1616.995 2697.220 1617.165 ;
        RECT 2697.045 1616.975 2697.215 1616.995 ;
        RECT 2698.425 1616.975 2698.595 1617.165 ;
        RECT 2700.265 1616.995 2700.435 1617.185 ;
        RECT 2703.945 1616.975 2704.115 1617.165 ;
        RECT 2705.785 1616.995 2705.955 1617.185 ;
        RECT 2709.005 1616.995 2709.175 1617.185 ;
        RECT 2709.465 1616.975 2709.635 1617.165 ;
        RECT 2714.525 1616.995 2714.695 1617.185 ;
        RECT 2714.985 1616.975 2715.155 1617.165 ;
        RECT 2720.045 1616.995 2720.215 1617.185 ;
        RECT 2720.515 1617.020 2720.675 1617.130 ;
        RECT 2721.885 1616.975 2722.055 1617.165 ;
        RECT 2725.565 1616.995 2725.735 1617.185 ;
        RECT 2727.405 1616.975 2727.575 1617.165 ;
        RECT 2731.085 1616.995 2731.255 1617.185 ;
        RECT 2733.845 1616.975 2734.015 1617.185 ;
        RECT 2695.525 1616.165 2696.895 1616.975 ;
        RECT 2696.905 1616.195 2698.275 1616.975 ;
        RECT 2698.285 1616.165 2703.795 1616.975 ;
        RECT 2703.805 1616.165 2709.315 1616.975 ;
        RECT 2709.325 1616.165 2714.835 1616.975 ;
        RECT 2714.845 1616.165 2720.355 1616.975 ;
        RECT 2721.745 1616.165 2727.255 1616.975 ;
        RECT 2727.265 1616.165 2732.775 1616.975 ;
        RECT 2732.785 1616.165 2734.155 1616.975 ;
        RECT 2695.525 1611.745 2696.895 1612.555 ;
        RECT 2696.905 1611.745 2698.275 1612.555 ;
        RECT 2698.285 1611.745 2701.955 1612.655 ;
        RECT 2701.965 1611.745 2707.475 1612.555 ;
        RECT 2708.865 1611.745 2714.375 1612.555 ;
        RECT 2714.385 1611.745 2719.895 1612.555 ;
        RECT 2719.905 1611.745 2725.415 1612.555 ;
        RECT 2725.425 1611.745 2730.935 1612.555 ;
        RECT 2730.945 1611.745 2732.775 1612.555 ;
        RECT 2732.785 1611.745 2734.155 1612.555 ;
        RECT 2695.665 1611.535 2695.835 1611.745 ;
        RECT 2697.045 1611.555 2697.215 1611.745 ;
        RECT 2695.525 1610.725 2696.895 1611.535 ;
        RECT 2697.965 1611.505 2698.135 1611.725 ;
        RECT 2701.640 1611.555 2701.810 1611.745 ;
        RECT 2702.105 1611.555 2702.275 1611.745 ;
        RECT 2703.485 1611.535 2703.655 1611.725 ;
        RECT 2703.945 1611.535 2704.115 1611.725 ;
        RECT 2707.635 1611.590 2707.795 1611.700 ;
        RECT 2709.005 1611.555 2709.175 1611.745 ;
        RECT 2709.465 1611.535 2709.635 1611.725 ;
        RECT 2714.525 1611.555 2714.695 1611.745 ;
        RECT 2714.985 1611.535 2715.155 1611.725 ;
        RECT 2720.045 1611.555 2720.215 1611.745 ;
        RECT 2720.515 1611.580 2720.675 1611.690 ;
        RECT 2721.885 1611.535 2722.055 1611.725 ;
        RECT 2725.565 1611.555 2725.735 1611.745 ;
        RECT 2727.405 1611.535 2727.575 1611.725 ;
        RECT 2731.085 1611.555 2731.255 1611.745 ;
        RECT 2733.845 1611.535 2734.015 1611.745 ;
        RECT 2700.090 1611.505 2701.035 1611.535 ;
        RECT 2697.965 1611.305 2701.035 1611.505 ;
        RECT 2697.825 1610.825 2701.035 1611.305 ;
        RECT 2697.825 1610.625 2698.755 1610.825 ;
        RECT 2700.090 1610.625 2701.035 1610.825 ;
        RECT 2701.275 1611.305 2703.655 1611.535 ;
        RECT 2701.275 1610.625 2703.665 1611.305 ;
        RECT 2703.805 1610.725 2709.315 1611.535 ;
        RECT 2709.325 1610.725 2714.835 1611.535 ;
        RECT 2714.845 1610.725 2720.355 1611.535 ;
        RECT 2721.745 1610.725 2727.255 1611.535 ;
        RECT 2727.265 1610.725 2732.775 1611.535 ;
        RECT 2732.785 1610.725 2734.155 1611.535 ;
        RECT 2364.460 1608.530 2365.060 1608.745 ;
        RECT 2381.680 1608.530 2382.280 1608.745 ;
        RECT 2398.900 1608.535 2399.500 1608.750 ;
        RECT 2364.460 1608.340 2365.355 1608.530 ;
        RECT 2367.485 1608.495 2367.655 1608.530 ;
        RECT 2366.580 1608.385 2367.655 1608.495 ;
        RECT 2367.370 1608.340 2367.655 1608.385 ;
        RECT 2369.795 1608.340 2369.965 1608.530 ;
        RECT 2371.175 1608.500 2371.345 1608.530 ;
        RECT 2371.175 1608.390 2371.745 1608.500 ;
        RECT 2371.175 1608.340 2371.460 1608.390 ;
        RECT 2364.460 1608.145 2366.420 1608.340 ;
        RECT 2365.070 1607.430 2366.420 1608.145 ;
        RECT 2367.370 1607.430 2371.460 1608.340 ;
        RECT 2381.680 1608.340 2382.575 1608.530 ;
        RECT 2384.705 1608.495 2384.875 1608.530 ;
        RECT 2383.800 1608.385 2384.875 1608.495 ;
        RECT 2384.590 1608.340 2384.875 1608.385 ;
        RECT 2387.015 1608.340 2387.185 1608.530 ;
        RECT 2388.395 1608.500 2388.565 1608.530 ;
        RECT 2388.395 1608.390 2388.965 1608.500 ;
        RECT 2388.395 1608.340 2388.680 1608.390 ;
        RECT 2381.680 1608.145 2383.640 1608.340 ;
        RECT 2382.290 1607.430 2383.640 1608.145 ;
        RECT 2384.590 1607.430 2388.680 1608.340 ;
        RECT 2398.900 1608.345 2399.795 1608.535 ;
        RECT 2401.925 1608.500 2402.095 1608.535 ;
        RECT 2401.020 1608.390 2402.095 1608.500 ;
        RECT 2401.810 1608.345 2402.095 1608.390 ;
        RECT 2404.235 1608.345 2404.405 1608.535 ;
        RECT 2405.615 1608.505 2405.785 1608.535 ;
        RECT 2416.120 1608.530 2416.720 1608.745 ;
        RECT 2433.340 1608.530 2433.940 1608.745 ;
        RECT 2405.615 1608.395 2406.185 1608.505 ;
        RECT 2405.615 1608.345 2405.900 1608.395 ;
        RECT 2398.900 1608.150 2400.860 1608.345 ;
        RECT 2399.510 1607.435 2400.860 1608.150 ;
        RECT 2401.810 1607.435 2405.900 1608.345 ;
        RECT 2416.120 1608.340 2417.015 1608.530 ;
        RECT 2419.145 1608.495 2419.315 1608.530 ;
        RECT 2418.240 1608.385 2419.315 1608.495 ;
        RECT 2419.030 1608.340 2419.315 1608.385 ;
        RECT 2421.455 1608.340 2421.625 1608.530 ;
        RECT 2422.835 1608.500 2423.005 1608.530 ;
        RECT 2422.835 1608.390 2423.405 1608.500 ;
        RECT 2422.835 1608.340 2423.120 1608.390 ;
        RECT 2416.120 1608.145 2418.080 1608.340 ;
        RECT 2416.730 1607.430 2418.080 1608.145 ;
        RECT 2419.030 1607.430 2423.120 1608.340 ;
        RECT 2433.340 1608.340 2434.235 1608.530 ;
        RECT 2436.365 1608.495 2436.535 1608.530 ;
        RECT 2435.460 1608.385 2436.535 1608.495 ;
        RECT 2436.250 1608.340 2436.535 1608.385 ;
        RECT 2438.675 1608.340 2438.845 1608.530 ;
        RECT 2440.055 1608.500 2440.225 1608.530 ;
        RECT 2440.055 1608.390 2440.625 1608.500 ;
        RECT 2440.055 1608.340 2440.340 1608.390 ;
        RECT 2433.340 1608.145 2435.300 1608.340 ;
        RECT 2433.950 1607.430 2435.300 1608.145 ;
        RECT 2436.250 1607.430 2440.340 1608.340 ;
        RECT 2695.525 1606.305 2696.895 1607.115 ;
        RECT 2696.905 1606.305 2698.275 1607.085 ;
        RECT 2698.745 1606.305 2700.095 1607.215 ;
        RECT 2700.125 1606.305 2705.635 1607.115 ;
        RECT 2705.645 1606.305 2708.395 1607.115 ;
        RECT 2708.865 1606.305 2714.375 1607.115 ;
        RECT 2714.385 1606.305 2719.895 1607.115 ;
        RECT 2719.905 1606.305 2725.415 1607.115 ;
        RECT 2725.425 1606.305 2730.935 1607.115 ;
        RECT 2730.945 1606.305 2732.775 1607.115 ;
        RECT 2732.785 1606.305 2734.155 1607.115 ;
        RECT 2695.665 1606.095 2695.835 1606.305 ;
        RECT 2697.045 1606.115 2697.215 1606.305 ;
        RECT 2698.420 1606.145 2698.540 1606.255 ;
        RECT 2699.810 1606.115 2699.980 1606.305 ;
        RECT 2700.265 1606.115 2700.435 1606.305 ;
        RECT 2700.450 1606.095 2700.620 1606.285 ;
        RECT 2701.185 1606.095 2701.355 1606.285 ;
        RECT 2705.785 1606.115 2705.955 1606.305 ;
        RECT 2706.705 1606.095 2706.875 1606.285 ;
        RECT 2709.005 1606.115 2709.175 1606.305 ;
        RECT 2712.225 1606.095 2712.395 1606.285 ;
        RECT 2714.525 1606.115 2714.695 1606.305 ;
        RECT 2717.745 1606.095 2717.915 1606.285 ;
        RECT 2720.045 1606.115 2720.215 1606.305 ;
        RECT 2721.885 1606.095 2722.055 1606.285 ;
        RECT 2725.565 1606.115 2725.735 1606.305 ;
        RECT 2727.405 1606.095 2727.575 1606.285 ;
        RECT 2731.085 1606.115 2731.255 1606.305 ;
        RECT 2733.845 1606.095 2734.015 1606.305 ;
        RECT 2695.525 1605.285 2696.895 1606.095 ;
        RECT 2697.135 1605.415 2701.035 1606.095 ;
        RECT 2700.105 1605.185 2701.035 1605.415 ;
        RECT 2701.045 1605.285 2706.555 1606.095 ;
        RECT 2706.565 1605.285 2712.075 1606.095 ;
        RECT 2712.085 1605.285 2717.595 1606.095 ;
        RECT 2717.605 1605.285 2721.275 1606.095 ;
        RECT 2721.745 1605.285 2727.255 1606.095 ;
        RECT 2727.265 1605.285 2732.775 1606.095 ;
        RECT 2732.785 1605.285 2734.155 1606.095 ;
        RECT 2364.600 1603.305 2371.900 1604.020 ;
        RECT 2381.820 1603.305 2389.120 1604.020 ;
        RECT 2399.040 1603.310 2406.340 1604.025 ;
        RECT 2364.460 1603.110 2371.900 1603.305 ;
        RECT 2381.680 1603.110 2389.120 1603.305 ;
        RECT 2398.900 1603.115 2406.340 1603.310 ;
        RECT 2416.260 1603.305 2423.560 1604.020 ;
        RECT 2433.480 1603.305 2440.780 1604.020 ;
        RECT 2364.460 1602.920 2365.820 1603.110 ;
        RECT 2367.025 1602.920 2367.665 1603.110 ;
        RECT 2371.630 1602.920 2371.800 1603.110 ;
        RECT 2381.680 1602.920 2383.040 1603.110 ;
        RECT 2384.245 1602.920 2384.885 1603.110 ;
        RECT 2388.850 1602.920 2389.020 1603.110 ;
        RECT 2398.900 1602.925 2400.260 1603.115 ;
        RECT 2401.465 1602.925 2402.105 1603.115 ;
        RECT 2406.070 1602.925 2406.240 1603.115 ;
        RECT 2416.120 1603.110 2423.560 1603.305 ;
        RECT 2433.340 1603.110 2440.780 1603.305 ;
        RECT 2364.460 1602.705 2365.060 1602.920 ;
        RECT 2381.680 1602.705 2382.280 1602.920 ;
        RECT 2398.900 1602.710 2399.500 1602.925 ;
        RECT 2416.120 1602.920 2417.480 1603.110 ;
        RECT 2418.685 1602.920 2419.325 1603.110 ;
        RECT 2423.290 1602.920 2423.460 1603.110 ;
        RECT 2433.340 1602.920 2434.700 1603.110 ;
        RECT 2435.905 1602.920 2436.545 1603.110 ;
        RECT 2440.510 1602.920 2440.680 1603.110 ;
        RECT 2416.120 1602.705 2416.720 1602.920 ;
        RECT 2433.340 1602.705 2433.940 1602.920 ;
        RECT 2695.525 1600.865 2696.895 1601.675 ;
        RECT 2696.905 1600.865 2698.275 1601.645 ;
        RECT 2698.285 1600.865 2703.795 1601.675 ;
        RECT 2703.805 1600.865 2707.475 1601.675 ;
        RECT 2708.865 1600.865 2714.375 1601.675 ;
        RECT 2714.385 1600.865 2719.895 1601.675 ;
        RECT 2719.905 1600.865 2725.415 1601.675 ;
        RECT 2725.425 1600.865 2730.935 1601.675 ;
        RECT 2730.945 1600.865 2732.775 1601.675 ;
        RECT 2732.785 1600.865 2734.155 1601.675 ;
        RECT 2695.665 1600.655 2695.835 1600.865 ;
        RECT 2697.045 1600.655 2697.215 1600.865 ;
        RECT 2698.425 1600.675 2698.595 1600.865 ;
        RECT 2702.565 1600.655 2702.735 1600.845 ;
        RECT 2703.945 1600.675 2704.115 1600.865 ;
        RECT 2707.635 1600.710 2707.795 1600.820 ;
        RECT 2708.085 1600.655 2708.255 1600.845 ;
        RECT 2709.005 1600.675 2709.175 1600.865 ;
        RECT 2713.605 1600.655 2713.775 1600.845 ;
        RECT 2714.525 1600.675 2714.695 1600.865 ;
        RECT 2719.125 1600.655 2719.295 1600.845 ;
        RECT 2720.045 1600.675 2720.215 1600.865 ;
        RECT 2720.960 1600.705 2721.080 1600.815 ;
        RECT 2721.885 1600.655 2722.055 1600.845 ;
        RECT 2725.565 1600.675 2725.735 1600.865 ;
        RECT 2727.405 1600.655 2727.575 1600.845 ;
        RECT 2731.085 1600.675 2731.255 1600.865 ;
        RECT 2733.845 1600.655 2734.015 1600.865 ;
        RECT 2695.525 1599.845 2696.895 1600.655 ;
        RECT 2696.905 1599.845 2702.415 1600.655 ;
        RECT 2702.425 1599.845 2707.935 1600.655 ;
        RECT 2707.945 1599.845 2713.455 1600.655 ;
        RECT 2713.465 1599.845 2718.975 1600.655 ;
        RECT 2718.985 1599.845 2720.815 1600.655 ;
        RECT 2721.745 1599.845 2727.255 1600.655 ;
        RECT 2727.265 1599.845 2732.775 1600.655 ;
        RECT 2732.785 1599.845 2734.155 1600.655 ;
        RECT 2695.525 1595.425 2696.895 1596.235 ;
        RECT 2696.905 1595.425 2698.275 1596.205 ;
        RECT 2698.285 1595.425 2703.795 1596.235 ;
        RECT 2703.805 1595.425 2707.475 1596.235 ;
        RECT 2708.865 1595.425 2714.375 1596.235 ;
        RECT 2714.385 1595.425 2719.895 1596.235 ;
        RECT 2719.905 1595.425 2725.415 1596.235 ;
        RECT 2725.425 1595.425 2730.935 1596.235 ;
        RECT 2730.945 1595.425 2732.775 1596.235 ;
        RECT 2732.785 1595.425 2734.155 1596.235 ;
        RECT 2695.665 1595.215 2695.835 1595.425 ;
        RECT 2697.045 1595.215 2697.215 1595.425 ;
        RECT 2698.425 1595.235 2698.595 1595.425 ;
        RECT 2702.565 1595.215 2702.735 1595.405 ;
        RECT 2703.945 1595.235 2704.115 1595.425 ;
        RECT 2707.635 1595.270 2707.795 1595.380 ;
        RECT 2708.085 1595.215 2708.255 1595.405 ;
        RECT 2709.005 1595.235 2709.175 1595.425 ;
        RECT 2713.605 1595.215 2713.775 1595.405 ;
        RECT 2714.525 1595.235 2714.695 1595.425 ;
        RECT 2719.125 1595.215 2719.295 1595.405 ;
        RECT 2720.045 1595.235 2720.215 1595.425 ;
        RECT 2720.960 1595.265 2721.080 1595.375 ;
        RECT 2721.885 1595.215 2722.055 1595.405 ;
        RECT 2725.565 1595.235 2725.735 1595.425 ;
        RECT 2727.405 1595.215 2727.575 1595.405 ;
        RECT 2731.085 1595.235 2731.255 1595.425 ;
        RECT 2733.845 1595.215 2734.015 1595.425 ;
        RECT 2695.525 1594.405 2696.895 1595.215 ;
        RECT 2696.905 1594.405 2702.415 1595.215 ;
        RECT 2702.425 1594.405 2707.935 1595.215 ;
        RECT 2707.945 1594.405 2713.455 1595.215 ;
        RECT 2713.465 1594.405 2718.975 1595.215 ;
        RECT 2718.985 1594.405 2720.815 1595.215 ;
        RECT 2721.745 1594.405 2727.255 1595.215 ;
        RECT 2727.265 1594.405 2732.775 1595.215 ;
        RECT 2732.785 1594.405 2734.155 1595.215 ;
        RECT 2695.525 1589.985 2696.895 1590.795 ;
        RECT 2696.905 1589.985 2698.275 1590.765 ;
        RECT 2698.285 1589.985 2699.655 1590.765 ;
        RECT 2699.665 1589.985 2705.175 1590.795 ;
        RECT 2705.185 1589.985 2707.935 1590.795 ;
        RECT 2708.865 1589.985 2714.375 1590.795 ;
        RECT 2714.385 1589.985 2719.895 1590.795 ;
        RECT 2719.905 1589.985 2721.275 1590.795 ;
        RECT 2721.745 1589.985 2727.255 1590.795 ;
        RECT 2727.265 1589.985 2732.775 1590.795 ;
        RECT 2732.785 1589.985 2734.155 1590.795 ;
        RECT 2695.665 1589.795 2695.835 1589.985 ;
        RECT 2697.045 1589.795 2697.215 1589.985 ;
        RECT 2698.425 1589.795 2698.595 1589.985 ;
        RECT 2699.805 1589.795 2699.975 1589.985 ;
        RECT 2705.325 1589.795 2705.495 1589.985 ;
        RECT 2708.080 1589.825 2708.200 1589.935 ;
        RECT 2709.005 1589.795 2709.175 1589.985 ;
        RECT 2714.525 1589.795 2714.695 1589.985 ;
        RECT 2720.045 1589.795 2720.215 1589.985 ;
        RECT 2721.885 1589.795 2722.055 1589.985 ;
        RECT 2727.405 1589.795 2727.575 1589.985 ;
        RECT 2733.845 1589.795 2734.015 1589.985 ;
        RECT 2522.700 1587.850 2522.870 1588.020 ;
        RECT 2522.700 1580.320 2522.870 1580.490 ;
        RECT 2522.700 1574.340 2522.870 1574.510 ;
        RECT 2522.700 1565.925 2522.870 1566.095 ;
        RECT 2361.695 1525.625 2361.865 1525.765 ;
        RECT 2361.675 1525.605 2361.865 1525.625 ;
        RECT 2364.135 1525.605 2364.305 1525.765 ;
        RECT 2366.575 1525.605 2366.745 1525.765 ;
        RECT 2369.015 1525.625 2369.185 1525.765 ;
        RECT 2378.020 1525.625 2378.190 1525.765 ;
        RECT 2369.015 1525.605 2369.205 1525.625 ;
        RECT 2361.675 1525.595 2361.845 1525.605 ;
        RECT 2369.035 1525.595 2369.205 1525.605 ;
        RECT 2378.000 1525.605 2378.190 1525.625 ;
        RECT 2380.460 1525.605 2380.630 1525.765 ;
        RECT 2382.900 1525.605 2383.070 1525.765 ;
        RECT 2385.340 1525.625 2385.510 1525.765 ;
        RECT 2394.345 1525.625 2394.515 1525.765 ;
        RECT 2385.340 1525.605 2385.530 1525.625 ;
        RECT 2378.000 1525.595 2378.170 1525.605 ;
        RECT 2385.360 1525.595 2385.530 1525.605 ;
        RECT 2394.325 1525.605 2394.515 1525.625 ;
        RECT 2396.785 1525.605 2396.955 1525.765 ;
        RECT 2399.225 1525.605 2399.395 1525.765 ;
        RECT 2401.665 1525.625 2401.835 1525.765 ;
        RECT 2410.670 1525.625 2410.840 1525.765 ;
        RECT 2401.665 1525.605 2401.855 1525.625 ;
        RECT 2394.325 1525.595 2394.495 1525.605 ;
        RECT 2401.685 1525.595 2401.855 1525.605 ;
        RECT 2410.650 1525.605 2410.840 1525.625 ;
        RECT 2413.110 1525.605 2413.280 1525.765 ;
        RECT 2415.550 1525.605 2415.720 1525.765 ;
        RECT 2417.990 1525.625 2418.160 1525.765 ;
        RECT 2426.995 1525.625 2427.165 1525.765 ;
        RECT 2417.990 1525.605 2418.180 1525.625 ;
        RECT 2410.650 1525.595 2410.820 1525.605 ;
        RECT 2418.010 1525.595 2418.180 1525.605 ;
        RECT 2426.975 1525.605 2427.165 1525.625 ;
        RECT 2429.435 1525.605 2429.605 1525.765 ;
        RECT 2431.875 1525.605 2432.045 1525.765 ;
        RECT 2434.315 1525.625 2434.485 1525.765 ;
        RECT 2434.315 1525.605 2434.505 1525.625 ;
        RECT 2426.975 1525.595 2427.145 1525.605 ;
        RECT 2434.335 1525.595 2434.505 1525.605 ;
        RECT 2695.665 1496.815 2695.835 1497.005 ;
        RECT 2697.045 1496.815 2697.215 1497.005 ;
        RECT 2699.805 1496.815 2699.975 1497.005 ;
        RECT 2701.185 1496.815 2701.355 1497.005 ;
        RECT 2701.645 1496.815 2701.815 1497.005 ;
        RECT 2707.165 1496.815 2707.335 1497.005 ;
        RECT 2709.005 1496.815 2709.175 1497.005 ;
        RECT 2710.845 1496.815 2711.015 1497.005 ;
        RECT 2716.365 1496.815 2716.535 1497.005 ;
        RECT 2720.045 1496.815 2720.215 1497.005 ;
        RECT 2723.265 1496.815 2723.435 1497.005 ;
        RECT 2723.725 1496.815 2723.895 1497.005 ;
        RECT 2729.245 1496.815 2729.415 1497.005 ;
        RECT 2731.080 1496.865 2731.200 1496.975 ;
        RECT 2732.455 1496.815 2732.625 1497.005 ;
        RECT 2733.845 1496.815 2734.015 1497.005 ;
        RECT 2695.525 1496.005 2696.895 1496.815 ;
        RECT 2696.905 1496.135 2698.735 1496.815 ;
        RECT 2698.745 1496.035 2700.115 1496.815 ;
        RECT 2700.125 1496.035 2701.495 1496.815 ;
        RECT 2701.505 1496.005 2707.015 1496.815 ;
        RECT 2707.025 1496.005 2708.395 1496.815 ;
        RECT 2708.865 1496.135 2710.695 1496.815 ;
        RECT 2709.350 1495.905 2710.695 1496.135 ;
        RECT 2710.705 1496.005 2716.215 1496.815 ;
        RECT 2716.225 1496.005 2719.895 1496.815 ;
        RECT 2719.905 1496.005 2721.275 1496.815 ;
        RECT 2721.745 1496.135 2723.575 1496.815 ;
        RECT 2723.585 1496.005 2729.095 1496.815 ;
        RECT 2729.105 1496.005 2730.935 1496.815 ;
        RECT 2731.405 1496.035 2732.775 1496.815 ;
        RECT 2732.785 1496.005 2734.155 1496.815 ;
        RECT 2695.525 1491.585 2696.895 1492.395 ;
        RECT 2696.905 1491.585 2698.275 1492.365 ;
        RECT 2698.285 1491.585 2703.795 1492.395 ;
        RECT 2703.805 1491.585 2707.475 1492.395 ;
        RECT 2708.865 1491.585 2714.375 1492.395 ;
        RECT 2714.385 1491.585 2719.895 1492.395 ;
        RECT 2719.905 1491.585 2725.415 1492.395 ;
        RECT 2725.425 1491.585 2730.935 1492.395 ;
        RECT 2730.945 1491.585 2732.775 1492.395 ;
        RECT 2732.785 1491.585 2734.155 1492.395 ;
        RECT 2695.665 1491.375 2695.835 1491.585 ;
        RECT 2697.045 1491.375 2697.215 1491.585 ;
        RECT 2698.425 1491.395 2698.595 1491.585 ;
        RECT 2702.565 1491.375 2702.735 1491.565 ;
        RECT 2703.945 1491.395 2704.115 1491.585 ;
        RECT 2707.635 1491.430 2707.795 1491.540 ;
        RECT 2708.085 1491.375 2708.255 1491.565 ;
        RECT 2709.005 1491.395 2709.175 1491.585 ;
        RECT 2713.605 1491.375 2713.775 1491.565 ;
        RECT 2714.525 1491.395 2714.695 1491.585 ;
        RECT 2719.125 1491.375 2719.295 1491.565 ;
        RECT 2720.045 1491.395 2720.215 1491.585 ;
        RECT 2720.960 1491.425 2721.080 1491.535 ;
        RECT 2721.885 1491.375 2722.055 1491.565 ;
        RECT 2725.565 1491.395 2725.735 1491.585 ;
        RECT 2727.405 1491.375 2727.575 1491.565 ;
        RECT 2731.085 1491.395 2731.255 1491.585 ;
        RECT 2733.845 1491.375 2734.015 1491.585 ;
        RECT 2695.525 1490.565 2696.895 1491.375 ;
        RECT 2696.905 1490.565 2702.415 1491.375 ;
        RECT 2702.425 1490.565 2707.935 1491.375 ;
        RECT 2707.945 1490.565 2713.455 1491.375 ;
        RECT 2713.465 1490.565 2718.975 1491.375 ;
        RECT 2718.985 1490.565 2720.815 1491.375 ;
        RECT 2721.745 1490.565 2727.255 1491.375 ;
        RECT 2727.265 1490.565 2732.775 1491.375 ;
        RECT 2732.785 1490.565 2734.155 1491.375 ;
        RECT 2695.525 1486.145 2696.895 1486.955 ;
        RECT 2696.905 1486.145 2702.415 1486.955 ;
        RECT 2702.425 1486.145 2707.935 1486.955 ;
        RECT 2708.865 1486.145 2714.375 1486.955 ;
        RECT 2714.385 1486.145 2719.895 1486.955 ;
        RECT 2719.905 1486.145 2725.415 1486.955 ;
        RECT 2725.425 1486.145 2730.935 1486.955 ;
        RECT 2730.945 1486.145 2732.775 1486.955 ;
        RECT 2732.785 1486.145 2734.155 1486.955 ;
        RECT 2695.665 1485.935 2695.835 1486.145 ;
        RECT 2697.045 1485.935 2697.215 1486.145 ;
        RECT 2698.425 1485.935 2698.595 1486.125 ;
        RECT 2702.565 1485.955 2702.735 1486.145 ;
        RECT 2703.945 1485.935 2704.115 1486.125 ;
        RECT 2708.080 1485.985 2708.200 1486.095 ;
        RECT 2709.005 1485.955 2709.175 1486.145 ;
        RECT 2709.465 1485.935 2709.635 1486.125 ;
        RECT 2714.525 1485.955 2714.695 1486.145 ;
        RECT 2714.985 1485.935 2715.155 1486.125 ;
        RECT 2720.045 1485.955 2720.215 1486.145 ;
        RECT 2720.515 1485.980 2720.675 1486.090 ;
        RECT 2721.885 1485.935 2722.055 1486.125 ;
        RECT 2725.565 1485.955 2725.735 1486.145 ;
        RECT 2727.405 1485.935 2727.575 1486.125 ;
        RECT 2731.085 1485.955 2731.255 1486.145 ;
        RECT 2733.845 1485.935 2734.015 1486.145 ;
        RECT 2695.525 1485.125 2696.895 1485.935 ;
        RECT 2696.905 1485.155 2698.275 1485.935 ;
        RECT 2698.285 1485.125 2703.795 1485.935 ;
        RECT 2703.805 1485.125 2709.315 1485.935 ;
        RECT 2709.325 1485.125 2714.835 1485.935 ;
        RECT 2714.845 1485.125 2720.355 1485.935 ;
        RECT 2721.745 1485.125 2727.255 1485.935 ;
        RECT 2727.265 1485.125 2732.775 1485.935 ;
        RECT 2732.785 1485.125 2734.155 1485.935 ;
        RECT 2695.525 1480.705 2696.895 1481.515 ;
        RECT 2696.905 1480.705 2702.415 1481.515 ;
        RECT 2702.425 1480.705 2707.935 1481.515 ;
        RECT 2708.865 1480.705 2714.375 1481.515 ;
        RECT 2714.385 1480.705 2719.895 1481.515 ;
        RECT 2719.905 1480.705 2725.415 1481.515 ;
        RECT 2725.425 1480.705 2730.935 1481.515 ;
        RECT 2730.945 1480.705 2732.775 1481.515 ;
        RECT 2732.785 1480.705 2734.155 1481.515 ;
        RECT 2695.665 1480.495 2695.835 1480.705 ;
        RECT 2697.045 1480.495 2697.215 1480.705 ;
        RECT 2702.565 1480.515 2702.735 1480.705 ;
        RECT 2706.705 1480.495 2706.875 1480.685 ;
        RECT 2708.080 1480.545 2708.200 1480.655 ;
        RECT 2709.005 1480.515 2709.175 1480.705 ;
        RECT 2712.225 1480.495 2712.395 1480.685 ;
        RECT 2714.525 1480.515 2714.695 1480.705 ;
        RECT 2717.745 1480.495 2717.915 1480.685 ;
        RECT 2720.045 1480.515 2720.215 1480.705 ;
        RECT 2721.885 1480.495 2722.055 1480.685 ;
        RECT 2725.565 1480.515 2725.735 1480.705 ;
        RECT 2727.405 1480.495 2727.575 1480.685 ;
        RECT 2731.085 1480.515 2731.255 1480.705 ;
        RECT 2733.845 1480.495 2734.015 1480.705 ;
        RECT 2695.525 1479.685 2696.895 1480.495 ;
        RECT 2696.905 1480.325 2698.665 1480.495 ;
        RECT 2696.905 1480.280 2699.160 1480.325 ;
        RECT 2696.905 1480.245 2700.100 1480.280 ;
        RECT 2701.460 1480.245 2706.555 1480.495 ;
        RECT 2696.905 1479.815 2706.555 1480.245 ;
        RECT 2698.230 1479.645 2701.460 1479.815 ;
        RECT 2699.170 1479.600 2701.460 1479.645 ;
        RECT 2700.110 1479.565 2701.460 1479.600 ;
        RECT 2704.535 1479.585 2706.555 1479.815 ;
        RECT 2706.565 1479.685 2712.075 1480.495 ;
        RECT 2712.085 1479.685 2717.595 1480.495 ;
        RECT 2717.605 1479.685 2721.275 1480.495 ;
        RECT 2721.745 1479.685 2727.255 1480.495 ;
        RECT 2727.265 1479.685 2732.775 1480.495 ;
        RECT 2732.785 1479.685 2734.155 1480.495 ;
        RECT 2704.535 1479.565 2705.455 1479.585 ;
        RECT 2695.525 1475.265 2696.895 1476.075 ;
        RECT 2696.905 1475.265 2698.275 1476.045 ;
        RECT 2698.285 1475.265 2703.795 1476.075 ;
        RECT 2703.805 1475.265 2707.475 1476.075 ;
        RECT 2708.865 1475.265 2714.375 1476.075 ;
        RECT 2714.385 1475.265 2719.895 1476.075 ;
        RECT 2719.905 1475.265 2725.415 1476.075 ;
        RECT 2725.425 1475.265 2730.935 1476.075 ;
        RECT 2730.945 1475.265 2732.775 1476.075 ;
        RECT 2732.785 1475.265 2734.155 1476.075 ;
        RECT 2695.665 1475.055 2695.835 1475.265 ;
        RECT 2697.045 1475.055 2697.215 1475.265 ;
        RECT 2698.425 1475.075 2698.595 1475.265 ;
        RECT 2703.945 1475.075 2704.115 1475.265 ;
        RECT 2706.705 1475.055 2706.875 1475.245 ;
        RECT 2707.635 1475.110 2707.795 1475.220 ;
        RECT 2709.005 1475.075 2709.175 1475.265 ;
        RECT 2712.225 1475.055 2712.395 1475.245 ;
        RECT 2714.525 1475.075 2714.695 1475.265 ;
        RECT 2717.745 1475.055 2717.915 1475.245 ;
        RECT 2720.045 1475.075 2720.215 1475.265 ;
        RECT 2721.885 1475.055 2722.055 1475.245 ;
        RECT 2725.565 1475.075 2725.735 1475.265 ;
        RECT 2727.405 1475.055 2727.575 1475.245 ;
        RECT 2731.085 1475.075 2731.255 1475.265 ;
        RECT 2733.845 1475.055 2734.015 1475.265 ;
        RECT 2695.525 1474.245 2696.895 1475.055 ;
        RECT 2696.905 1474.885 2698.665 1475.055 ;
        RECT 2696.905 1474.840 2699.160 1474.885 ;
        RECT 2696.905 1474.805 2700.100 1474.840 ;
        RECT 2701.460 1474.805 2706.555 1475.055 ;
        RECT 2696.905 1474.375 2706.555 1474.805 ;
        RECT 2698.230 1474.205 2701.460 1474.375 ;
        RECT 2699.170 1474.160 2701.460 1474.205 ;
        RECT 2700.110 1474.125 2701.460 1474.160 ;
        RECT 2704.535 1474.145 2706.555 1474.375 ;
        RECT 2706.565 1474.245 2712.075 1475.055 ;
        RECT 2712.085 1474.245 2717.595 1475.055 ;
        RECT 2717.605 1474.245 2721.275 1475.055 ;
        RECT 2721.745 1474.245 2727.255 1475.055 ;
        RECT 2727.265 1474.245 2732.775 1475.055 ;
        RECT 2732.785 1474.245 2734.155 1475.055 ;
        RECT 2704.535 1474.125 2705.455 1474.145 ;
        RECT 2695.525 1469.825 2696.895 1470.635 ;
        RECT 2696.905 1469.825 2698.275 1470.605 ;
        RECT 2698.285 1469.825 2701.035 1470.635 ;
        RECT 2701.505 1470.505 2702.435 1470.735 ;
        RECT 2701.505 1469.825 2705.405 1470.505 ;
        RECT 2705.645 1469.825 2708.395 1470.635 ;
        RECT 2708.865 1469.825 2714.375 1470.635 ;
        RECT 2714.385 1469.825 2719.895 1470.635 ;
        RECT 2719.905 1469.825 2725.415 1470.635 ;
        RECT 2725.425 1469.825 2730.935 1470.635 ;
        RECT 2730.945 1469.825 2732.775 1470.635 ;
        RECT 2732.785 1469.825 2734.155 1470.635 ;
        RECT 2695.665 1469.615 2695.835 1469.825 ;
        RECT 2697.045 1469.615 2697.215 1469.825 ;
        RECT 2698.425 1469.635 2698.595 1469.825 ;
        RECT 2701.180 1469.665 2701.300 1469.775 ;
        RECT 2701.920 1469.635 2702.090 1469.825 ;
        RECT 2702.565 1469.615 2702.735 1469.805 ;
        RECT 2705.785 1469.635 2705.955 1469.825 ;
        RECT 2708.085 1469.615 2708.255 1469.805 ;
        RECT 2709.005 1469.635 2709.175 1469.825 ;
        RECT 2713.605 1469.615 2713.775 1469.805 ;
        RECT 2714.525 1469.635 2714.695 1469.825 ;
        RECT 2719.125 1469.615 2719.295 1469.805 ;
        RECT 2720.045 1469.635 2720.215 1469.825 ;
        RECT 2720.960 1469.665 2721.080 1469.775 ;
        RECT 2721.885 1469.615 2722.055 1469.805 ;
        RECT 2725.565 1469.635 2725.735 1469.825 ;
        RECT 2727.405 1469.615 2727.575 1469.805 ;
        RECT 2731.085 1469.635 2731.255 1469.825 ;
        RECT 2733.845 1469.615 2734.015 1469.825 ;
        RECT 2695.525 1468.805 2696.895 1469.615 ;
        RECT 2696.905 1468.805 2702.415 1469.615 ;
        RECT 2702.425 1468.805 2707.935 1469.615 ;
        RECT 2707.945 1468.805 2713.455 1469.615 ;
        RECT 2713.465 1468.805 2718.975 1469.615 ;
        RECT 2718.985 1468.805 2720.815 1469.615 ;
        RECT 2721.745 1468.805 2727.255 1469.615 ;
        RECT 2727.265 1468.805 2732.775 1469.615 ;
        RECT 2732.785 1468.805 2734.155 1469.615 ;
        RECT 2695.525 1464.385 2696.895 1465.195 ;
        RECT 2696.905 1464.385 2698.275 1465.165 ;
        RECT 2698.285 1464.385 2703.795 1465.195 ;
        RECT 2703.805 1464.385 2707.475 1465.195 ;
        RECT 2708.865 1464.385 2714.375 1465.195 ;
        RECT 2714.385 1464.385 2719.895 1465.195 ;
        RECT 2719.905 1464.385 2725.415 1465.195 ;
        RECT 2725.425 1464.385 2730.935 1465.195 ;
        RECT 2730.945 1464.385 2732.775 1465.195 ;
        RECT 2732.785 1464.385 2734.155 1465.195 ;
        RECT 2695.665 1464.175 2695.835 1464.385 ;
        RECT 2697.045 1464.175 2697.215 1464.385 ;
        RECT 2698.425 1464.195 2698.595 1464.385 ;
        RECT 2702.565 1464.175 2702.735 1464.365 ;
        RECT 2703.945 1464.195 2704.115 1464.385 ;
        RECT 2707.635 1464.230 2707.795 1464.340 ;
        RECT 2708.085 1464.175 2708.255 1464.365 ;
        RECT 2709.005 1464.195 2709.175 1464.385 ;
        RECT 2713.605 1464.175 2713.775 1464.365 ;
        RECT 2714.525 1464.195 2714.695 1464.385 ;
        RECT 2719.125 1464.175 2719.295 1464.365 ;
        RECT 2720.045 1464.195 2720.215 1464.385 ;
        RECT 2720.960 1464.225 2721.080 1464.335 ;
        RECT 2721.885 1464.175 2722.055 1464.365 ;
        RECT 2725.565 1464.195 2725.735 1464.385 ;
        RECT 2727.405 1464.175 2727.575 1464.365 ;
        RECT 2731.085 1464.195 2731.255 1464.385 ;
        RECT 2733.845 1464.175 2734.015 1464.385 ;
        RECT 2695.525 1463.365 2696.895 1464.175 ;
        RECT 2696.905 1463.365 2702.415 1464.175 ;
        RECT 2702.425 1463.365 2707.935 1464.175 ;
        RECT 2707.945 1463.365 2713.455 1464.175 ;
        RECT 2713.465 1463.365 2718.975 1464.175 ;
        RECT 2718.985 1463.365 2720.815 1464.175 ;
        RECT 2721.745 1463.365 2727.255 1464.175 ;
        RECT 2727.265 1463.365 2732.775 1464.175 ;
        RECT 2732.785 1463.365 2734.155 1464.175 ;
        RECT 2695.525 1458.945 2696.895 1459.755 ;
        RECT 2696.905 1458.945 2700.575 1459.755 ;
        RECT 2701.505 1458.945 2702.855 1459.855 ;
        RECT 2702.885 1458.945 2708.395 1459.755 ;
        RECT 2708.865 1458.945 2714.375 1459.755 ;
        RECT 2714.385 1458.945 2719.895 1459.755 ;
        RECT 2719.905 1458.945 2725.415 1459.755 ;
        RECT 2725.425 1458.945 2730.935 1459.755 ;
        RECT 2730.945 1458.945 2732.775 1459.755 ;
        RECT 2732.785 1458.945 2734.155 1459.755 ;
        RECT 2695.665 1458.735 2695.835 1458.945 ;
        RECT 2697.045 1458.735 2697.215 1458.945 ;
        RECT 2698.425 1458.735 2698.595 1458.925 ;
        RECT 2700.735 1458.790 2700.895 1458.900 ;
        RECT 2701.650 1458.755 2701.820 1458.945 ;
        RECT 2703.025 1458.755 2703.195 1458.945 ;
        RECT 2704.865 1458.735 2705.035 1458.925 ;
        RECT 2705.325 1458.735 2705.495 1458.925 ;
        RECT 2709.005 1458.755 2709.175 1458.945 ;
        RECT 2710.845 1458.735 2711.015 1458.925 ;
        RECT 2714.525 1458.755 2714.695 1458.945 ;
        RECT 2716.365 1458.735 2716.535 1458.925 ;
        RECT 2720.045 1458.735 2720.215 1458.945 ;
        RECT 2721.885 1458.735 2722.055 1458.925 ;
        RECT 2725.565 1458.755 2725.735 1458.945 ;
        RECT 2727.405 1458.735 2727.575 1458.925 ;
        RECT 2731.085 1458.755 2731.255 1458.945 ;
        RECT 2733.845 1458.735 2734.015 1458.945 ;
        RECT 2695.525 1457.925 2696.895 1458.735 ;
        RECT 2696.905 1457.955 2698.275 1458.735 ;
        RECT 2698.285 1457.925 2701.955 1458.735 ;
        RECT 2701.965 1457.825 2705.175 1458.735 ;
        RECT 2705.185 1457.925 2710.695 1458.735 ;
        RECT 2710.705 1457.925 2716.215 1458.735 ;
        RECT 2716.225 1457.925 2719.895 1458.735 ;
        RECT 2719.905 1457.925 2721.275 1458.735 ;
        RECT 2721.745 1457.925 2727.255 1458.735 ;
        RECT 2727.265 1457.925 2732.775 1458.735 ;
        RECT 2732.785 1457.925 2734.155 1458.735 ;
        RECT 2695.525 1453.505 2696.895 1454.315 ;
        RECT 2696.905 1453.505 2702.415 1454.315 ;
        RECT 2702.425 1453.505 2707.935 1454.315 ;
        RECT 2708.865 1453.505 2714.375 1454.315 ;
        RECT 2714.385 1453.505 2719.895 1454.315 ;
        RECT 2719.905 1453.505 2725.415 1454.315 ;
        RECT 2725.425 1453.505 2732.775 1454.415 ;
        RECT 2732.785 1453.505 2734.155 1454.315 ;
        RECT 2695.665 1453.295 2695.835 1453.505 ;
        RECT 2697.045 1453.295 2697.215 1453.505 ;
        RECT 2698.425 1453.295 2698.595 1453.485 ;
        RECT 2702.565 1453.315 2702.735 1453.505 ;
        RECT 2703.945 1453.295 2704.115 1453.485 ;
        RECT 2708.080 1453.345 2708.200 1453.455 ;
        RECT 2709.005 1453.315 2709.175 1453.505 ;
        RECT 2709.465 1453.295 2709.635 1453.485 ;
        RECT 2714.525 1453.315 2714.695 1453.505 ;
        RECT 2714.985 1453.295 2715.155 1453.485 ;
        RECT 2720.045 1453.315 2720.215 1453.505 ;
        RECT 2720.515 1453.340 2720.675 1453.450 ;
        RECT 2721.885 1453.295 2722.055 1453.485 ;
        RECT 2725.990 1453.315 2726.160 1453.505 ;
        RECT 2727.405 1453.295 2727.575 1453.485 ;
        RECT 2733.845 1453.295 2734.015 1453.505 ;
        RECT 2695.525 1452.485 2696.895 1453.295 ;
        RECT 2696.905 1452.515 2698.275 1453.295 ;
        RECT 2698.285 1452.485 2703.795 1453.295 ;
        RECT 2703.805 1452.485 2709.315 1453.295 ;
        RECT 2709.325 1452.485 2714.835 1453.295 ;
        RECT 2714.845 1452.485 2720.355 1453.295 ;
        RECT 2721.745 1452.485 2727.255 1453.295 ;
        RECT 2727.265 1452.485 2732.775 1453.295 ;
        RECT 2732.785 1452.485 2734.155 1453.295 ;
        RECT 2695.525 1448.065 2696.895 1448.875 ;
        RECT 2696.905 1448.065 2702.415 1448.875 ;
        RECT 2702.425 1448.065 2707.935 1448.875 ;
        RECT 2708.865 1448.065 2714.375 1448.875 ;
        RECT 2714.385 1448.065 2719.895 1448.875 ;
        RECT 2719.905 1448.065 2725.415 1448.875 ;
        RECT 2725.425 1448.065 2730.935 1448.875 ;
        RECT 2730.945 1448.065 2732.775 1448.875 ;
        RECT 2732.785 1448.065 2734.155 1448.875 ;
        RECT 2695.665 1447.855 2695.835 1448.065 ;
        RECT 2697.045 1447.875 2697.215 1448.065 ;
        RECT 2699.345 1447.875 2699.515 1448.045 ;
        RECT 2699.345 1447.855 2699.475 1447.875 ;
        RECT 2699.805 1447.855 2699.975 1448.045 ;
        RECT 2702.565 1447.875 2702.735 1448.065 ;
        RECT 2705.325 1447.855 2705.495 1448.045 ;
        RECT 2708.080 1447.905 2708.200 1448.015 ;
        RECT 2709.005 1447.875 2709.175 1448.065 ;
        RECT 2710.845 1447.855 2711.015 1448.045 ;
        RECT 2714.525 1447.875 2714.695 1448.065 ;
        RECT 2716.365 1447.855 2716.535 1448.045 ;
        RECT 2720.045 1447.855 2720.215 1448.065 ;
        RECT 2721.885 1447.855 2722.055 1448.045 ;
        RECT 2725.565 1447.875 2725.735 1448.065 ;
        RECT 2727.405 1447.855 2727.575 1448.045 ;
        RECT 2731.085 1447.875 2731.255 1448.065 ;
        RECT 2733.845 1447.855 2734.015 1448.065 ;
        RECT 2695.525 1447.045 2696.895 1447.855 ;
        RECT 2697.625 1447.625 2699.475 1447.855 ;
        RECT 2697.140 1446.945 2699.475 1447.625 ;
        RECT 2699.665 1447.045 2705.175 1447.855 ;
        RECT 2705.185 1447.045 2710.695 1447.855 ;
        RECT 2710.705 1447.045 2716.215 1447.855 ;
        RECT 2716.225 1447.045 2719.895 1447.855 ;
        RECT 2719.905 1447.045 2721.275 1447.855 ;
        RECT 2721.745 1447.045 2727.255 1447.855 ;
        RECT 2727.265 1447.045 2732.775 1447.855 ;
        RECT 2732.785 1447.045 2734.155 1447.855 ;
        RECT 2695.525 1442.625 2696.895 1443.435 ;
        RECT 2696.905 1442.625 2698.275 1443.405 ;
        RECT 2698.285 1442.625 2703.795 1443.435 ;
        RECT 2703.805 1442.625 2707.475 1443.435 ;
        RECT 2708.865 1442.625 2714.375 1443.435 ;
        RECT 2714.385 1442.625 2719.895 1443.435 ;
        RECT 2719.905 1442.625 2725.415 1443.435 ;
        RECT 2725.425 1442.625 2730.935 1443.435 ;
        RECT 2730.945 1442.625 2732.775 1443.435 ;
        RECT 2732.785 1442.625 2734.155 1443.435 ;
        RECT 2695.665 1442.415 2695.835 1442.625 ;
        RECT 2697.045 1442.435 2697.215 1442.625 ;
        RECT 2698.425 1442.435 2698.595 1442.625 ;
        RECT 2700.450 1442.415 2700.620 1442.605 ;
        RECT 2702.575 1442.415 2702.745 1442.585 ;
        RECT 2703.945 1442.435 2704.115 1442.625 ;
        RECT 2704.405 1442.415 2704.575 1442.605 ;
        RECT 2704.865 1442.415 2705.035 1442.605 ;
        RECT 2707.635 1442.470 2707.795 1442.580 ;
        RECT 2709.005 1442.435 2709.175 1442.625 ;
        RECT 2710.385 1442.415 2710.555 1442.605 ;
        RECT 2714.525 1442.435 2714.695 1442.625 ;
        RECT 2715.905 1442.415 2716.075 1442.605 ;
        RECT 2720.045 1442.435 2720.215 1442.625 ;
        RECT 2721.885 1442.415 2722.055 1442.605 ;
        RECT 2725.565 1442.435 2725.735 1442.625 ;
        RECT 2727.405 1442.415 2727.575 1442.605 ;
        RECT 2731.085 1442.435 2731.255 1442.625 ;
        RECT 2733.845 1442.415 2734.015 1442.625 ;
        RECT 2695.525 1441.605 2696.895 1442.415 ;
        RECT 2697.135 1441.735 2701.035 1442.415 ;
        RECT 2700.105 1441.505 2701.035 1441.735 ;
        RECT 2701.045 1441.505 2704.695 1442.415 ;
        RECT 2704.725 1441.605 2710.235 1442.415 ;
        RECT 2710.245 1441.605 2715.755 1442.415 ;
        RECT 2715.765 1441.605 2721.275 1442.415 ;
        RECT 2721.745 1441.605 2727.255 1442.415 ;
        RECT 2727.265 1441.605 2732.775 1442.415 ;
        RECT 2732.785 1441.605 2734.155 1442.415 ;
        RECT 2695.525 1437.185 2696.895 1437.995 ;
        RECT 2696.905 1437.895 2697.835 1438.095 ;
        RECT 2699.165 1437.895 2700.115 1438.095 ;
        RECT 2696.905 1437.415 2700.115 1437.895 ;
        RECT 2697.050 1437.215 2700.115 1437.415 ;
        RECT 2695.665 1436.975 2695.835 1437.185 ;
        RECT 2697.050 1437.165 2697.220 1437.215 ;
        RECT 2699.180 1437.185 2700.115 1437.215 ;
        RECT 2700.125 1437.185 2705.635 1437.995 ;
        RECT 2705.645 1437.185 2708.395 1437.995 ;
        RECT 2708.865 1437.185 2714.375 1437.995 ;
        RECT 2714.385 1437.185 2719.895 1437.995 ;
        RECT 2719.905 1437.185 2725.415 1437.995 ;
        RECT 2725.425 1437.185 2730.935 1437.995 ;
        RECT 2730.945 1437.185 2732.775 1437.995 ;
        RECT 2732.785 1437.185 2734.155 1437.995 ;
        RECT 2697.045 1436.995 2697.220 1437.165 ;
        RECT 2697.045 1436.975 2697.215 1436.995 ;
        RECT 2698.425 1436.975 2698.595 1437.165 ;
        RECT 2700.265 1436.995 2700.435 1437.185 ;
        RECT 2703.945 1436.975 2704.115 1437.165 ;
        RECT 2705.785 1436.995 2705.955 1437.185 ;
        RECT 2709.005 1436.995 2709.175 1437.185 ;
        RECT 2709.465 1436.975 2709.635 1437.165 ;
        RECT 2714.525 1436.995 2714.695 1437.185 ;
        RECT 2714.985 1436.975 2715.155 1437.165 ;
        RECT 2720.045 1436.995 2720.215 1437.185 ;
        RECT 2720.515 1437.020 2720.675 1437.130 ;
        RECT 2721.885 1436.975 2722.055 1437.165 ;
        RECT 2725.565 1436.995 2725.735 1437.185 ;
        RECT 2727.405 1436.975 2727.575 1437.165 ;
        RECT 2731.085 1436.995 2731.255 1437.185 ;
        RECT 2733.845 1436.975 2734.015 1437.185 ;
        RECT 2522.700 1436.225 2522.870 1436.395 ;
        RECT 2695.525 1436.165 2696.895 1436.975 ;
        RECT 2696.905 1436.195 2698.275 1436.975 ;
        RECT 2698.285 1436.165 2703.795 1436.975 ;
        RECT 2703.805 1436.165 2709.315 1436.975 ;
        RECT 2709.325 1436.165 2714.835 1436.975 ;
        RECT 2714.845 1436.165 2720.355 1436.975 ;
        RECT 2721.745 1436.165 2727.255 1436.975 ;
        RECT 2727.265 1436.165 2732.775 1436.975 ;
        RECT 2732.785 1436.165 2734.155 1436.975 ;
        RECT 2695.525 1431.745 2696.895 1432.555 ;
        RECT 2696.905 1431.745 2698.275 1432.555 ;
        RECT 2698.285 1431.745 2701.955 1432.655 ;
        RECT 2701.965 1431.745 2707.475 1432.555 ;
        RECT 2708.865 1431.745 2714.375 1432.555 ;
        RECT 2714.385 1431.745 2719.895 1432.555 ;
        RECT 2719.905 1431.745 2725.415 1432.555 ;
        RECT 2725.425 1431.745 2730.935 1432.555 ;
        RECT 2730.945 1431.745 2732.775 1432.555 ;
        RECT 2732.785 1431.745 2734.155 1432.555 ;
        RECT 2695.665 1431.535 2695.835 1431.745 ;
        RECT 2697.045 1431.555 2697.215 1431.745 ;
        RECT 2695.525 1430.725 2696.895 1431.535 ;
        RECT 2697.965 1431.505 2698.135 1431.725 ;
        RECT 2701.640 1431.555 2701.810 1431.745 ;
        RECT 2702.105 1431.555 2702.275 1431.745 ;
        RECT 2703.485 1431.535 2703.655 1431.725 ;
        RECT 2703.945 1431.535 2704.115 1431.725 ;
        RECT 2707.635 1431.590 2707.795 1431.700 ;
        RECT 2709.005 1431.555 2709.175 1431.745 ;
        RECT 2709.465 1431.535 2709.635 1431.725 ;
        RECT 2714.525 1431.555 2714.695 1431.745 ;
        RECT 2714.985 1431.535 2715.155 1431.725 ;
        RECT 2720.045 1431.555 2720.215 1431.745 ;
        RECT 2720.515 1431.580 2720.675 1431.690 ;
        RECT 2721.885 1431.535 2722.055 1431.725 ;
        RECT 2725.565 1431.555 2725.735 1431.745 ;
        RECT 2727.405 1431.535 2727.575 1431.725 ;
        RECT 2731.085 1431.555 2731.255 1431.745 ;
        RECT 2733.845 1431.535 2734.015 1431.745 ;
        RECT 2700.090 1431.505 2701.035 1431.535 ;
        RECT 2697.965 1431.305 2701.035 1431.505 ;
        RECT 2697.825 1430.825 2701.035 1431.305 ;
        RECT 2697.825 1430.625 2698.755 1430.825 ;
        RECT 2700.090 1430.625 2701.035 1430.825 ;
        RECT 2701.275 1431.305 2703.655 1431.535 ;
        RECT 2701.275 1430.625 2703.665 1431.305 ;
        RECT 2703.805 1430.725 2709.315 1431.535 ;
        RECT 2709.325 1430.725 2714.835 1431.535 ;
        RECT 2714.845 1430.725 2720.355 1431.535 ;
        RECT 2721.745 1430.725 2727.255 1431.535 ;
        RECT 2727.265 1430.725 2732.775 1431.535 ;
        RECT 2732.785 1430.725 2734.155 1431.535 ;
        RECT 2522.700 1429.810 2522.870 1429.980 ;
        RECT 2361.700 1427.735 2361.870 1427.875 ;
        RECT 2361.680 1427.715 2361.870 1427.735 ;
        RECT 2361.680 1427.705 2361.850 1427.715 ;
        RECT 2363.660 1427.705 2363.830 1427.875 ;
        RECT 2366.100 1427.705 2366.270 1427.875 ;
        RECT 2368.540 1427.705 2368.710 1427.875 ;
        RECT 2370.500 1427.705 2370.670 1427.875 ;
        RECT 2380.260 1427.735 2380.430 1427.875 ;
        RECT 2380.240 1427.715 2380.430 1427.735 ;
        RECT 2380.240 1427.705 2380.410 1427.715 ;
        RECT 2382.220 1427.705 2382.390 1427.875 ;
        RECT 2384.660 1427.705 2384.830 1427.875 ;
        RECT 2387.100 1427.705 2387.270 1427.875 ;
        RECT 2389.060 1427.705 2389.230 1427.875 ;
        RECT 2398.820 1427.735 2398.990 1427.875 ;
        RECT 2398.800 1427.715 2398.990 1427.735 ;
        RECT 2398.800 1427.705 2398.970 1427.715 ;
        RECT 2400.780 1427.705 2400.950 1427.875 ;
        RECT 2403.220 1427.705 2403.390 1427.875 ;
        RECT 2405.660 1427.705 2405.830 1427.875 ;
        RECT 2407.620 1427.705 2407.790 1427.875 ;
        RECT 2417.380 1427.735 2417.550 1427.875 ;
        RECT 2417.360 1427.715 2417.550 1427.735 ;
        RECT 2417.360 1427.705 2417.530 1427.715 ;
        RECT 2419.340 1427.705 2419.510 1427.875 ;
        RECT 2421.780 1427.705 2421.950 1427.875 ;
        RECT 2424.220 1427.705 2424.390 1427.875 ;
        RECT 2426.180 1427.705 2426.350 1427.875 ;
        RECT 2435.940 1427.735 2436.110 1427.875 ;
        RECT 2435.920 1427.715 2436.110 1427.735 ;
        RECT 2435.920 1427.705 2436.090 1427.715 ;
        RECT 2437.900 1427.705 2438.070 1427.875 ;
        RECT 2440.340 1427.705 2440.510 1427.875 ;
        RECT 2442.780 1427.705 2442.950 1427.875 ;
        RECT 2444.740 1427.705 2444.910 1427.875 ;
        RECT 2695.525 1426.305 2696.895 1427.115 ;
        RECT 2696.905 1426.305 2698.275 1427.085 ;
        RECT 2698.745 1426.305 2700.095 1427.215 ;
        RECT 2700.125 1426.305 2705.635 1427.115 ;
        RECT 2705.645 1426.305 2708.395 1427.115 ;
        RECT 2708.865 1426.305 2714.375 1427.115 ;
        RECT 2714.385 1426.305 2719.895 1427.115 ;
        RECT 2719.905 1426.305 2725.415 1427.115 ;
        RECT 2725.425 1426.305 2730.935 1427.115 ;
        RECT 2730.945 1426.305 2732.775 1427.115 ;
        RECT 2732.785 1426.305 2734.155 1427.115 ;
        RECT 2695.665 1426.095 2695.835 1426.305 ;
        RECT 2697.045 1426.115 2697.215 1426.305 ;
        RECT 2698.420 1426.145 2698.540 1426.255 ;
        RECT 2699.810 1426.115 2699.980 1426.305 ;
        RECT 2700.265 1426.115 2700.435 1426.305 ;
        RECT 2700.450 1426.095 2700.620 1426.285 ;
        RECT 2701.185 1426.095 2701.355 1426.285 ;
        RECT 2705.785 1426.115 2705.955 1426.305 ;
        RECT 2706.705 1426.095 2706.875 1426.285 ;
        RECT 2709.005 1426.115 2709.175 1426.305 ;
        RECT 2712.225 1426.095 2712.395 1426.285 ;
        RECT 2714.525 1426.115 2714.695 1426.305 ;
        RECT 2717.745 1426.095 2717.915 1426.285 ;
        RECT 2720.045 1426.115 2720.215 1426.305 ;
        RECT 2721.885 1426.095 2722.055 1426.285 ;
        RECT 2725.565 1426.115 2725.735 1426.305 ;
        RECT 2727.405 1426.095 2727.575 1426.285 ;
        RECT 2731.085 1426.115 2731.255 1426.305 ;
        RECT 2733.845 1426.095 2734.015 1426.305 ;
        RECT 2695.525 1425.285 2696.895 1426.095 ;
        RECT 2697.135 1425.415 2701.035 1426.095 ;
        RECT 2700.105 1425.185 2701.035 1425.415 ;
        RECT 2701.045 1425.285 2706.555 1426.095 ;
        RECT 2706.565 1425.285 2712.075 1426.095 ;
        RECT 2712.085 1425.285 2717.595 1426.095 ;
        RECT 2717.605 1425.285 2721.275 1426.095 ;
        RECT 2721.745 1425.285 2727.255 1426.095 ;
        RECT 2727.265 1425.285 2732.775 1426.095 ;
        RECT 2732.785 1425.285 2734.155 1426.095 ;
        RECT 2695.525 1420.865 2696.895 1421.675 ;
        RECT 2696.905 1420.865 2698.275 1421.645 ;
        RECT 2698.285 1420.865 2703.795 1421.675 ;
        RECT 2703.805 1420.865 2707.475 1421.675 ;
        RECT 2708.865 1420.865 2714.375 1421.675 ;
        RECT 2714.385 1420.865 2719.895 1421.675 ;
        RECT 2719.905 1420.865 2725.415 1421.675 ;
        RECT 2725.425 1420.865 2730.935 1421.675 ;
        RECT 2730.945 1420.865 2732.775 1421.675 ;
        RECT 2732.785 1420.865 2734.155 1421.675 ;
        RECT 2695.665 1420.655 2695.835 1420.865 ;
        RECT 2697.045 1420.655 2697.215 1420.865 ;
        RECT 2698.425 1420.675 2698.595 1420.865 ;
        RECT 2702.565 1420.655 2702.735 1420.845 ;
        RECT 2703.945 1420.675 2704.115 1420.865 ;
        RECT 2707.635 1420.710 2707.795 1420.820 ;
        RECT 2708.085 1420.655 2708.255 1420.845 ;
        RECT 2709.005 1420.675 2709.175 1420.865 ;
        RECT 2713.605 1420.655 2713.775 1420.845 ;
        RECT 2714.525 1420.675 2714.695 1420.865 ;
        RECT 2719.125 1420.655 2719.295 1420.845 ;
        RECT 2720.045 1420.675 2720.215 1420.865 ;
        RECT 2720.960 1420.705 2721.080 1420.815 ;
        RECT 2721.885 1420.655 2722.055 1420.845 ;
        RECT 2725.565 1420.675 2725.735 1420.865 ;
        RECT 2727.405 1420.655 2727.575 1420.845 ;
        RECT 2731.085 1420.675 2731.255 1420.865 ;
        RECT 2733.845 1420.655 2734.015 1420.865 ;
        RECT 2695.525 1419.845 2696.895 1420.655 ;
        RECT 2696.905 1419.845 2702.415 1420.655 ;
        RECT 2702.425 1419.845 2707.935 1420.655 ;
        RECT 2707.945 1419.845 2713.455 1420.655 ;
        RECT 2713.465 1419.845 2718.975 1420.655 ;
        RECT 2718.985 1419.845 2720.815 1420.655 ;
        RECT 2721.745 1419.845 2727.255 1420.655 ;
        RECT 2727.265 1419.845 2732.775 1420.655 ;
        RECT 2732.785 1419.845 2734.155 1420.655 ;
        RECT 2522.700 1415.620 2522.870 1415.790 ;
        RECT 2695.525 1415.425 2696.895 1416.235 ;
        RECT 2696.905 1415.425 2698.275 1416.205 ;
        RECT 2698.285 1415.425 2703.795 1416.235 ;
        RECT 2703.805 1415.425 2707.475 1416.235 ;
        RECT 2708.865 1415.425 2714.375 1416.235 ;
        RECT 2714.385 1415.425 2719.895 1416.235 ;
        RECT 2719.905 1415.425 2725.415 1416.235 ;
        RECT 2725.425 1415.425 2730.935 1416.235 ;
        RECT 2730.945 1415.425 2732.775 1416.235 ;
        RECT 2732.785 1415.425 2734.155 1416.235 ;
        RECT 2695.665 1415.215 2695.835 1415.425 ;
        RECT 2697.045 1415.215 2697.215 1415.425 ;
        RECT 2698.425 1415.235 2698.595 1415.425 ;
        RECT 2702.565 1415.215 2702.735 1415.405 ;
        RECT 2703.945 1415.235 2704.115 1415.425 ;
        RECT 2707.635 1415.270 2707.795 1415.380 ;
        RECT 2708.085 1415.215 2708.255 1415.405 ;
        RECT 2709.005 1415.235 2709.175 1415.425 ;
        RECT 2713.605 1415.215 2713.775 1415.405 ;
        RECT 2714.525 1415.235 2714.695 1415.425 ;
        RECT 2719.125 1415.215 2719.295 1415.405 ;
        RECT 2720.045 1415.235 2720.215 1415.425 ;
        RECT 2720.960 1415.265 2721.080 1415.375 ;
        RECT 2721.885 1415.215 2722.055 1415.405 ;
        RECT 2725.565 1415.235 2725.735 1415.425 ;
        RECT 2727.405 1415.215 2727.575 1415.405 ;
        RECT 2731.085 1415.235 2731.255 1415.425 ;
        RECT 2733.845 1415.215 2734.015 1415.425 ;
        RECT 2695.525 1414.405 2696.895 1415.215 ;
        RECT 2696.905 1414.405 2702.415 1415.215 ;
        RECT 2702.425 1414.405 2707.935 1415.215 ;
        RECT 2707.945 1414.405 2713.455 1415.215 ;
        RECT 2713.465 1414.405 2718.975 1415.215 ;
        RECT 2718.985 1414.405 2720.815 1415.215 ;
        RECT 2721.745 1414.405 2727.255 1415.215 ;
        RECT 2727.265 1414.405 2732.775 1415.215 ;
        RECT 2732.785 1414.405 2734.155 1415.215 ;
        RECT 2695.525 1409.985 2696.895 1410.795 ;
        RECT 2696.905 1409.985 2698.275 1410.765 ;
        RECT 2698.285 1409.985 2699.655 1410.765 ;
        RECT 2699.665 1409.985 2705.175 1410.795 ;
        RECT 2705.185 1409.985 2707.935 1410.795 ;
        RECT 2708.865 1409.985 2714.375 1410.795 ;
        RECT 2714.385 1409.985 2719.895 1410.795 ;
        RECT 2719.905 1409.985 2721.275 1410.795 ;
        RECT 2721.745 1409.985 2727.255 1410.795 ;
        RECT 2727.265 1409.985 2732.775 1410.795 ;
        RECT 2732.785 1409.985 2734.155 1410.795 ;
        RECT 2695.665 1409.795 2695.835 1409.985 ;
        RECT 2697.045 1409.795 2697.215 1409.985 ;
        RECT 2698.425 1409.795 2698.595 1409.985 ;
        RECT 2699.805 1409.795 2699.975 1409.985 ;
        RECT 2705.325 1409.795 2705.495 1409.985 ;
        RECT 2708.080 1409.825 2708.200 1409.935 ;
        RECT 2709.005 1409.795 2709.175 1409.985 ;
        RECT 2714.525 1409.795 2714.695 1409.985 ;
        RECT 2720.045 1409.795 2720.215 1409.985 ;
        RECT 2721.885 1409.795 2722.055 1409.985 ;
        RECT 2727.405 1409.795 2727.575 1409.985 ;
        RECT 2733.845 1409.795 2734.015 1409.985 ;
        RECT 2522.700 1408.090 2522.870 1408.260 ;
        RECT 2522.700 1402.110 2522.870 1402.280 ;
        RECT 2522.700 1393.695 2522.870 1393.865 ;
        RECT 2883.065 1360.420 2883.235 1360.590 ;
        RECT 2371.925 1327.715 2372.095 1327.875 ;
        RECT 2387.185 1327.715 2387.355 1327.875 ;
        RECT 2402.445 1327.715 2402.615 1327.875 ;
        RECT 2417.705 1327.715 2417.875 1327.875 ;
        RECT 2432.965 1327.715 2433.135 1327.875 ;
        RECT 2883.065 1161.180 2883.235 1161.350 ;
      LAYER li1 ;
        RECT 1262.890 3510.650 1263.410 3512.135 ;
        RECT 1622.890 3511.100 1623.410 3512.585 ;
        RECT 1802.890 3509.180 1803.410 3510.665 ;
        RECT 2162.890 3508.820 2163.410 3510.305 ;
        RECT 2522.890 3509.505 2523.410 3510.990 ;
        RECT 2882.085 3486.420 2882.605 3487.970 ;
        RECT 2882.085 3220.540 2882.605 3222.090 ;
        RECT 2882.085 2955.340 2882.605 2956.890 ;
        RECT 2882.085 2689.460 2882.605 2691.010 ;
        RECT 2882.085 2423.580 2882.605 2425.130 ;
        RECT 2358.655 2255.095 2358.830 2255.585 ;
        RECT 2359.180 2255.305 2359.350 2255.585 ;
        RECT 2359.180 2255.135 2359.410 2255.305 ;
        RECT 2358.655 2254.925 2358.825 2255.095 ;
        RECT 2358.655 2254.595 2359.065 2254.925 ;
        RECT 2358.655 2254.085 2358.825 2254.595 ;
        RECT 2358.655 2253.755 2359.065 2254.085 ;
        RECT 2358.655 2253.555 2358.825 2253.755 ;
        RECT 2358.655 2252.295 2358.830 2253.555 ;
        RECT 2359.240 2253.525 2359.410 2255.135 ;
        RECT 2359.610 2255.075 2359.785 2255.585 ;
        RECT 2361.885 2255.095 2362.060 2255.585 ;
        RECT 2361.885 2254.925 2362.055 2255.095 ;
        RECT 2362.840 2255.075 2363.015 2255.585 ;
        RECT 2363.270 2255.035 2363.445 2255.585 ;
        RECT 2373.110 2255.100 2373.285 2255.590 ;
        RECT 2373.635 2255.310 2373.805 2255.590 ;
        RECT 2373.635 2255.140 2373.865 2255.310 ;
        RECT 2361.885 2254.595 2362.295 2254.925 ;
        RECT 2359.180 2253.355 2359.410 2253.525 ;
        RECT 2359.610 2253.555 2359.780 2254.505 ;
        RECT 2361.885 2254.085 2362.055 2254.595 ;
        RECT 2361.885 2253.755 2362.295 2254.085 ;
        RECT 2361.885 2253.555 2362.055 2253.755 ;
        RECT 2362.840 2253.555 2363.010 2254.505 ;
        RECT 2359.180 2252.295 2359.350 2253.355 ;
        RECT 2359.610 2252.295 2359.785 2253.555 ;
        RECT 2361.885 2252.295 2362.060 2253.555 ;
        RECT 2362.840 2252.295 2363.015 2253.555 ;
        RECT 2363.270 2253.435 2363.440 2255.035 ;
        RECT 2373.110 2254.930 2373.280 2255.100 ;
        RECT 2373.110 2254.600 2373.520 2254.930 ;
        RECT 2373.110 2254.090 2373.280 2254.600 ;
        RECT 2373.110 2253.760 2373.520 2254.090 ;
        RECT 2373.110 2253.560 2373.280 2253.760 ;
        RECT 2363.270 2252.295 2363.445 2253.435 ;
        RECT 2365.060 2252.895 2365.620 2253.185 ;
        RECT 2366.660 2253.055 2366.920 2253.085 ;
        RECT 2365.060 2251.525 2365.310 2252.895 ;
        RECT 2366.660 2252.725 2366.990 2253.055 ;
        RECT 2368.370 2252.935 2369.680 2253.185 ;
        RECT 2368.370 2252.785 2368.550 2252.935 ;
        RECT 2365.600 2252.535 2366.990 2252.725 ;
        RECT 2367.820 2252.615 2368.550 2252.785 ;
        RECT 2365.600 2252.445 2365.770 2252.535 ;
        RECT 2365.480 2252.115 2365.770 2252.445 ;
        RECT 2366.500 2252.115 2367.180 2252.365 ;
        RECT 2365.600 2251.865 2365.770 2252.115 ;
        RECT 2365.600 2251.695 2366.545 2251.865 ;
        RECT 2366.910 2251.755 2367.180 2252.115 ;
        RECT 2367.820 2251.945 2367.990 2252.615 ;
        RECT 2368.800 2252.365 2369.010 2252.765 ;
        RECT 2368.660 2252.165 2369.010 2252.365 ;
        RECT 2369.260 2252.365 2369.510 2252.765 ;
        RECT 2369.260 2252.165 2369.730 2252.365 ;
        RECT 2369.920 2252.165 2370.370 2252.675 ;
        RECT 2373.110 2252.300 2373.285 2253.560 ;
        RECT 2373.695 2253.530 2373.865 2255.140 ;
        RECT 2374.065 2255.080 2374.240 2255.590 ;
        RECT 2374.495 2255.040 2374.670 2255.590 ;
        RECT 2375.860 2255.080 2376.030 2255.590 ;
        RECT 2376.850 2255.080 2377.020 2255.590 ;
        RECT 2378.470 2255.095 2378.645 2255.585 ;
        RECT 2373.635 2253.360 2373.865 2253.530 ;
        RECT 2374.065 2253.560 2374.235 2254.510 ;
        RECT 2373.635 2252.300 2373.805 2253.360 ;
        RECT 2374.065 2252.300 2374.240 2253.560 ;
        RECT 2374.495 2253.440 2374.665 2255.040 ;
        RECT 2378.470 2254.925 2378.640 2255.095 ;
        RECT 2379.425 2255.075 2379.600 2255.585 ;
        RECT 2379.855 2255.035 2380.030 2255.585 ;
        RECT 2389.695 2255.100 2389.870 2255.590 ;
        RECT 2390.220 2255.310 2390.390 2255.590 ;
        RECT 2390.220 2255.140 2390.450 2255.310 ;
        RECT 2378.470 2254.595 2378.880 2254.925 ;
        RECT 2375.035 2254.475 2375.265 2254.570 ;
        RECT 2375.035 2254.420 2375.655 2254.475 ;
        RECT 2375.035 2254.305 2375.955 2254.420 ;
        RECT 2375.485 2254.250 2375.955 2254.305 ;
        RECT 2376.475 2254.250 2376.945 2254.420 ;
        RECT 2375.485 2253.560 2375.655 2254.250 ;
        RECT 2375.855 2253.770 2376.025 2253.880 ;
        RECT 2376.475 2253.770 2376.645 2254.250 ;
        RECT 2378.470 2254.085 2378.640 2254.595 ;
        RECT 2375.855 2253.600 2376.645 2253.770 ;
        RECT 2374.495 2252.300 2374.670 2253.440 ;
        RECT 2375.855 2252.300 2376.030 2253.600 ;
        RECT 2376.475 2253.560 2376.645 2253.600 ;
        RECT 2376.845 2253.445 2377.015 2253.880 ;
        RECT 2378.470 2253.755 2378.880 2254.085 ;
        RECT 2378.470 2253.555 2378.640 2253.755 ;
        RECT 2379.425 2253.555 2379.595 2254.505 ;
        RECT 2376.845 2252.300 2377.020 2253.445 ;
        RECT 2378.470 2252.295 2378.645 2253.555 ;
        RECT 2379.425 2252.295 2379.600 2253.555 ;
        RECT 2379.855 2253.435 2380.025 2255.035 ;
        RECT 2389.695 2254.930 2389.865 2255.100 ;
        RECT 2389.695 2254.600 2390.105 2254.930 ;
        RECT 2389.695 2254.090 2389.865 2254.600 ;
        RECT 2389.695 2253.760 2390.105 2254.090 ;
        RECT 2389.695 2253.560 2389.865 2253.760 ;
        RECT 2379.855 2252.295 2380.030 2253.435 ;
        RECT 2381.645 2252.895 2382.205 2253.185 ;
        RECT 2383.245 2253.055 2383.505 2253.085 ;
        RECT 2368.660 2251.945 2370.400 2251.995 ;
        RECT 2367.820 2251.815 2370.400 2251.945 ;
        RECT 2367.820 2251.775 2368.880 2251.815 ;
        RECT 2365.060 2250.975 2365.520 2251.525 ;
        RECT 2366.240 2250.975 2366.545 2251.695 ;
        RECT 2369.020 2251.605 2369.900 2251.645 ;
        RECT 2368.370 2251.405 2369.900 2251.605 ;
        RECT 2368.370 2251.275 2368.540 2251.405 ;
        RECT 2369.290 2251.355 2369.900 2251.405 ;
        RECT 2369.670 2251.315 2369.900 2251.355 ;
        RECT 2370.070 2251.315 2370.400 2251.815 ;
        RECT 2381.645 2251.525 2381.895 2252.895 ;
        RECT 2383.245 2252.725 2383.575 2253.055 ;
        RECT 2384.955 2252.935 2386.265 2253.185 ;
        RECT 2384.955 2252.785 2385.135 2252.935 ;
        RECT 2382.185 2252.535 2383.575 2252.725 ;
        RECT 2384.405 2252.615 2385.135 2252.785 ;
        RECT 2382.185 2252.445 2382.355 2252.535 ;
        RECT 2382.065 2252.115 2382.355 2252.445 ;
        RECT 2383.085 2252.115 2383.765 2252.365 ;
        RECT 2382.185 2251.865 2382.355 2252.115 ;
        RECT 2382.185 2251.695 2383.130 2251.865 ;
        RECT 2383.495 2251.755 2383.765 2252.115 ;
        RECT 2384.405 2251.945 2384.575 2252.615 ;
        RECT 2385.385 2252.365 2385.595 2252.765 ;
        RECT 2385.245 2252.165 2385.595 2252.365 ;
        RECT 2385.845 2252.365 2386.095 2252.765 ;
        RECT 2385.845 2252.165 2386.315 2252.365 ;
        RECT 2386.505 2252.165 2386.955 2252.675 ;
        RECT 2389.695 2252.300 2389.870 2253.560 ;
        RECT 2390.280 2253.530 2390.450 2255.140 ;
        RECT 2390.650 2255.080 2390.825 2255.590 ;
        RECT 2391.080 2255.040 2391.255 2255.590 ;
        RECT 2392.445 2255.080 2392.615 2255.590 ;
        RECT 2393.435 2255.080 2393.605 2255.590 ;
        RECT 2395.055 2255.095 2395.230 2255.585 ;
        RECT 2390.220 2253.360 2390.450 2253.530 ;
        RECT 2390.650 2253.560 2390.820 2254.510 ;
        RECT 2390.220 2252.300 2390.390 2253.360 ;
        RECT 2390.650 2252.300 2390.825 2253.560 ;
        RECT 2391.080 2253.440 2391.250 2255.040 ;
        RECT 2395.055 2254.925 2395.225 2255.095 ;
        RECT 2396.010 2255.075 2396.185 2255.585 ;
        RECT 2396.440 2255.035 2396.615 2255.585 ;
        RECT 2406.280 2255.100 2406.455 2255.590 ;
        RECT 2406.805 2255.310 2406.975 2255.590 ;
        RECT 2406.805 2255.140 2407.035 2255.310 ;
        RECT 2395.055 2254.595 2395.465 2254.925 ;
        RECT 2391.620 2254.475 2391.850 2254.570 ;
        RECT 2391.620 2254.420 2392.240 2254.475 ;
        RECT 2391.620 2254.305 2392.540 2254.420 ;
        RECT 2392.070 2254.250 2392.540 2254.305 ;
        RECT 2393.060 2254.250 2393.530 2254.420 ;
        RECT 2392.070 2253.560 2392.240 2254.250 ;
        RECT 2392.440 2253.770 2392.610 2253.880 ;
        RECT 2393.060 2253.770 2393.230 2254.250 ;
        RECT 2395.055 2254.085 2395.225 2254.595 ;
        RECT 2392.440 2253.600 2393.230 2253.770 ;
        RECT 2391.080 2252.300 2391.255 2253.440 ;
        RECT 2392.440 2252.300 2392.615 2253.600 ;
        RECT 2393.060 2253.560 2393.230 2253.600 ;
        RECT 2393.430 2253.445 2393.600 2253.880 ;
        RECT 2395.055 2253.755 2395.465 2254.085 ;
        RECT 2395.055 2253.555 2395.225 2253.755 ;
        RECT 2396.010 2253.555 2396.180 2254.505 ;
        RECT 2393.430 2252.300 2393.605 2253.445 ;
        RECT 2395.055 2252.295 2395.230 2253.555 ;
        RECT 2396.010 2252.295 2396.185 2253.555 ;
        RECT 2396.440 2253.435 2396.610 2255.035 ;
        RECT 2406.280 2254.930 2406.450 2255.100 ;
        RECT 2406.280 2254.600 2406.690 2254.930 ;
        RECT 2406.280 2254.090 2406.450 2254.600 ;
        RECT 2406.280 2253.760 2406.690 2254.090 ;
        RECT 2406.280 2253.560 2406.450 2253.760 ;
        RECT 2396.440 2252.295 2396.615 2253.435 ;
        RECT 2398.230 2252.895 2398.790 2253.185 ;
        RECT 2399.830 2253.055 2400.090 2253.085 ;
        RECT 2385.245 2251.945 2386.985 2251.995 ;
        RECT 2384.405 2251.815 2386.985 2251.945 ;
        RECT 2384.405 2251.775 2385.465 2251.815 ;
        RECT 2369.230 2251.145 2369.560 2251.185 ;
        RECT 2370.070 2251.145 2370.890 2251.315 ;
        RECT 2369.230 2250.975 2370.400 2251.145 ;
        RECT 2381.645 2250.975 2382.105 2251.525 ;
        RECT 2382.825 2250.975 2383.130 2251.695 ;
        RECT 2385.605 2251.605 2386.485 2251.645 ;
        RECT 2384.955 2251.405 2386.485 2251.605 ;
        RECT 2384.955 2251.275 2385.125 2251.405 ;
        RECT 2385.875 2251.355 2386.485 2251.405 ;
        RECT 2386.255 2251.315 2386.485 2251.355 ;
        RECT 2386.655 2251.315 2386.985 2251.815 ;
        RECT 2398.230 2251.525 2398.480 2252.895 ;
        RECT 2399.830 2252.725 2400.160 2253.055 ;
        RECT 2401.540 2252.935 2402.850 2253.185 ;
        RECT 2401.540 2252.785 2401.720 2252.935 ;
        RECT 2398.770 2252.535 2400.160 2252.725 ;
        RECT 2400.990 2252.615 2401.720 2252.785 ;
        RECT 2398.770 2252.445 2398.940 2252.535 ;
        RECT 2398.650 2252.115 2398.940 2252.445 ;
        RECT 2399.670 2252.115 2400.350 2252.365 ;
        RECT 2398.770 2251.865 2398.940 2252.115 ;
        RECT 2398.770 2251.695 2399.715 2251.865 ;
        RECT 2400.080 2251.755 2400.350 2252.115 ;
        RECT 2400.990 2251.945 2401.160 2252.615 ;
        RECT 2401.970 2252.365 2402.180 2252.765 ;
        RECT 2401.830 2252.165 2402.180 2252.365 ;
        RECT 2402.430 2252.365 2402.680 2252.765 ;
        RECT 2402.430 2252.165 2402.900 2252.365 ;
        RECT 2403.090 2252.165 2403.540 2252.675 ;
        RECT 2406.280 2252.300 2406.455 2253.560 ;
        RECT 2406.865 2253.530 2407.035 2255.140 ;
        RECT 2407.235 2255.080 2407.410 2255.590 ;
        RECT 2407.665 2255.040 2407.840 2255.590 ;
        RECT 2409.030 2255.080 2409.200 2255.590 ;
        RECT 2410.020 2255.080 2410.190 2255.590 ;
        RECT 2411.640 2255.095 2411.815 2255.585 ;
        RECT 2406.805 2253.360 2407.035 2253.530 ;
        RECT 2407.235 2253.560 2407.405 2254.510 ;
        RECT 2406.805 2252.300 2406.975 2253.360 ;
        RECT 2407.235 2252.300 2407.410 2253.560 ;
        RECT 2407.665 2253.440 2407.835 2255.040 ;
        RECT 2411.640 2254.925 2411.810 2255.095 ;
        RECT 2412.595 2255.075 2412.770 2255.585 ;
        RECT 2413.025 2255.035 2413.200 2255.585 ;
        RECT 2422.865 2255.100 2423.040 2255.590 ;
        RECT 2423.390 2255.310 2423.560 2255.590 ;
        RECT 2423.390 2255.140 2423.620 2255.310 ;
        RECT 2411.640 2254.595 2412.050 2254.925 ;
        RECT 2408.205 2254.475 2408.435 2254.570 ;
        RECT 2408.205 2254.420 2408.825 2254.475 ;
        RECT 2408.205 2254.305 2409.125 2254.420 ;
        RECT 2408.655 2254.250 2409.125 2254.305 ;
        RECT 2409.645 2254.250 2410.115 2254.420 ;
        RECT 2408.655 2253.560 2408.825 2254.250 ;
        RECT 2409.025 2253.770 2409.195 2253.880 ;
        RECT 2409.645 2253.770 2409.815 2254.250 ;
        RECT 2411.640 2254.085 2411.810 2254.595 ;
        RECT 2409.025 2253.600 2409.815 2253.770 ;
        RECT 2407.665 2252.300 2407.840 2253.440 ;
        RECT 2409.025 2252.300 2409.200 2253.600 ;
        RECT 2409.645 2253.560 2409.815 2253.600 ;
        RECT 2410.015 2253.445 2410.185 2253.880 ;
        RECT 2411.640 2253.755 2412.050 2254.085 ;
        RECT 2411.640 2253.555 2411.810 2253.755 ;
        RECT 2412.595 2253.555 2412.765 2254.505 ;
        RECT 2410.015 2252.300 2410.190 2253.445 ;
        RECT 2411.640 2252.295 2411.815 2253.555 ;
        RECT 2412.595 2252.295 2412.770 2253.555 ;
        RECT 2413.025 2253.435 2413.195 2255.035 ;
        RECT 2422.865 2254.930 2423.035 2255.100 ;
        RECT 2422.865 2254.600 2423.275 2254.930 ;
        RECT 2422.865 2254.090 2423.035 2254.600 ;
        RECT 2422.865 2253.760 2423.275 2254.090 ;
        RECT 2422.865 2253.560 2423.035 2253.760 ;
        RECT 2413.025 2252.295 2413.200 2253.435 ;
        RECT 2414.815 2252.895 2415.375 2253.185 ;
        RECT 2416.415 2253.055 2416.675 2253.085 ;
        RECT 2401.830 2251.945 2403.570 2251.995 ;
        RECT 2400.990 2251.815 2403.570 2251.945 ;
        RECT 2400.990 2251.775 2402.050 2251.815 ;
        RECT 2385.815 2251.145 2386.145 2251.185 ;
        RECT 2386.655 2251.145 2387.475 2251.315 ;
        RECT 2385.815 2250.975 2386.985 2251.145 ;
        RECT 2398.230 2250.975 2398.690 2251.525 ;
        RECT 2399.410 2250.975 2399.715 2251.695 ;
        RECT 2402.190 2251.605 2403.070 2251.645 ;
        RECT 2401.540 2251.405 2403.070 2251.605 ;
        RECT 2401.540 2251.275 2401.710 2251.405 ;
        RECT 2402.460 2251.355 2403.070 2251.405 ;
        RECT 2402.840 2251.315 2403.070 2251.355 ;
        RECT 2403.240 2251.315 2403.570 2251.815 ;
        RECT 2414.815 2251.525 2415.065 2252.895 ;
        RECT 2416.415 2252.725 2416.745 2253.055 ;
        RECT 2418.125 2252.935 2419.435 2253.185 ;
        RECT 2418.125 2252.785 2418.305 2252.935 ;
        RECT 2415.355 2252.535 2416.745 2252.725 ;
        RECT 2417.575 2252.615 2418.305 2252.785 ;
        RECT 2415.355 2252.445 2415.525 2252.535 ;
        RECT 2415.235 2252.115 2415.525 2252.445 ;
        RECT 2416.255 2252.115 2416.935 2252.365 ;
        RECT 2415.355 2251.865 2415.525 2252.115 ;
        RECT 2415.355 2251.695 2416.300 2251.865 ;
        RECT 2416.665 2251.755 2416.935 2252.115 ;
        RECT 2417.575 2251.945 2417.745 2252.615 ;
        RECT 2418.555 2252.365 2418.765 2252.765 ;
        RECT 2418.415 2252.165 2418.765 2252.365 ;
        RECT 2419.015 2252.365 2419.265 2252.765 ;
        RECT 2419.015 2252.165 2419.485 2252.365 ;
        RECT 2419.675 2252.165 2420.125 2252.675 ;
        RECT 2422.865 2252.300 2423.040 2253.560 ;
        RECT 2423.450 2253.530 2423.620 2255.140 ;
        RECT 2423.820 2255.080 2423.995 2255.590 ;
        RECT 2424.250 2255.040 2424.425 2255.590 ;
        RECT 2425.615 2255.080 2425.785 2255.590 ;
        RECT 2426.605 2255.080 2426.775 2255.590 ;
        RECT 2428.220 2255.095 2428.395 2255.585 ;
        RECT 2423.390 2253.360 2423.620 2253.530 ;
        RECT 2423.820 2253.560 2423.990 2254.510 ;
        RECT 2423.390 2252.300 2423.560 2253.360 ;
        RECT 2423.820 2252.300 2423.995 2253.560 ;
        RECT 2424.250 2253.440 2424.420 2255.040 ;
        RECT 2428.220 2254.925 2428.390 2255.095 ;
        RECT 2429.175 2255.075 2429.350 2255.585 ;
        RECT 2429.605 2255.035 2429.780 2255.585 ;
        RECT 2439.445 2255.100 2439.620 2255.590 ;
        RECT 2439.970 2255.310 2440.140 2255.590 ;
        RECT 2439.970 2255.140 2440.200 2255.310 ;
        RECT 2428.220 2254.595 2428.630 2254.925 ;
        RECT 2424.790 2254.475 2425.020 2254.570 ;
        RECT 2424.790 2254.420 2425.410 2254.475 ;
        RECT 2424.790 2254.305 2425.710 2254.420 ;
        RECT 2425.240 2254.250 2425.710 2254.305 ;
        RECT 2426.230 2254.250 2426.700 2254.420 ;
        RECT 2425.240 2253.560 2425.410 2254.250 ;
        RECT 2425.610 2253.770 2425.780 2253.880 ;
        RECT 2426.230 2253.770 2426.400 2254.250 ;
        RECT 2428.220 2254.085 2428.390 2254.595 ;
        RECT 2425.610 2253.600 2426.400 2253.770 ;
        RECT 2424.250 2252.300 2424.425 2253.440 ;
        RECT 2425.610 2252.300 2425.785 2253.600 ;
        RECT 2426.230 2253.560 2426.400 2253.600 ;
        RECT 2426.600 2253.445 2426.770 2253.880 ;
        RECT 2428.220 2253.755 2428.630 2254.085 ;
        RECT 2428.220 2253.555 2428.390 2253.755 ;
        RECT 2429.175 2253.555 2429.345 2254.505 ;
        RECT 2426.600 2252.300 2426.775 2253.445 ;
        RECT 2428.220 2252.295 2428.395 2253.555 ;
        RECT 2429.175 2252.295 2429.350 2253.555 ;
        RECT 2429.605 2253.435 2429.775 2255.035 ;
        RECT 2439.445 2254.930 2439.615 2255.100 ;
        RECT 2439.445 2254.600 2439.855 2254.930 ;
        RECT 2439.445 2254.090 2439.615 2254.600 ;
        RECT 2439.445 2253.760 2439.855 2254.090 ;
        RECT 2439.445 2253.560 2439.615 2253.760 ;
        RECT 2429.605 2252.295 2429.780 2253.435 ;
        RECT 2431.395 2252.895 2431.955 2253.185 ;
        RECT 2432.995 2253.055 2433.255 2253.085 ;
        RECT 2418.415 2251.945 2420.155 2251.995 ;
        RECT 2417.575 2251.815 2420.155 2251.945 ;
        RECT 2417.575 2251.775 2418.635 2251.815 ;
        RECT 2402.400 2251.145 2402.730 2251.185 ;
        RECT 2403.240 2251.145 2404.060 2251.315 ;
        RECT 2402.400 2250.975 2403.570 2251.145 ;
        RECT 2414.815 2250.975 2415.275 2251.525 ;
        RECT 2415.995 2250.975 2416.300 2251.695 ;
        RECT 2418.775 2251.605 2419.655 2251.645 ;
        RECT 2418.125 2251.405 2419.655 2251.605 ;
        RECT 2418.125 2251.275 2418.295 2251.405 ;
        RECT 2419.045 2251.355 2419.655 2251.405 ;
        RECT 2419.425 2251.315 2419.655 2251.355 ;
        RECT 2419.825 2251.315 2420.155 2251.815 ;
        RECT 2431.395 2251.525 2431.645 2252.895 ;
        RECT 2432.995 2252.725 2433.325 2253.055 ;
        RECT 2434.705 2252.935 2436.015 2253.185 ;
        RECT 2434.705 2252.785 2434.885 2252.935 ;
        RECT 2431.935 2252.535 2433.325 2252.725 ;
        RECT 2434.155 2252.615 2434.885 2252.785 ;
        RECT 2431.935 2252.445 2432.105 2252.535 ;
        RECT 2431.815 2252.115 2432.105 2252.445 ;
        RECT 2432.835 2252.115 2433.515 2252.365 ;
        RECT 2431.935 2251.865 2432.105 2252.115 ;
        RECT 2431.935 2251.695 2432.880 2251.865 ;
        RECT 2433.245 2251.755 2433.515 2252.115 ;
        RECT 2434.155 2251.945 2434.325 2252.615 ;
        RECT 2435.135 2252.365 2435.345 2252.765 ;
        RECT 2434.995 2252.165 2435.345 2252.365 ;
        RECT 2435.595 2252.365 2435.845 2252.765 ;
        RECT 2435.595 2252.165 2436.065 2252.365 ;
        RECT 2436.255 2252.165 2436.705 2252.675 ;
        RECT 2439.445 2252.300 2439.620 2253.560 ;
        RECT 2440.030 2253.530 2440.200 2255.140 ;
        RECT 2440.400 2255.080 2440.575 2255.590 ;
        RECT 2440.830 2255.040 2441.005 2255.590 ;
        RECT 2442.195 2255.080 2442.365 2255.590 ;
        RECT 2443.185 2255.080 2443.355 2255.590 ;
        RECT 2439.970 2253.360 2440.200 2253.530 ;
        RECT 2440.400 2253.560 2440.570 2254.510 ;
        RECT 2439.970 2252.300 2440.140 2253.360 ;
        RECT 2440.400 2252.300 2440.575 2253.560 ;
        RECT 2440.830 2253.440 2441.000 2255.040 ;
        RECT 2441.370 2254.475 2441.600 2254.570 ;
        RECT 2441.370 2254.420 2441.990 2254.475 ;
        RECT 2441.370 2254.305 2442.290 2254.420 ;
        RECT 2441.820 2254.250 2442.290 2254.305 ;
        RECT 2442.810 2254.250 2443.280 2254.420 ;
        RECT 2441.820 2253.560 2441.990 2254.250 ;
        RECT 2442.190 2253.770 2442.360 2253.880 ;
        RECT 2442.810 2253.770 2442.980 2254.250 ;
        RECT 2442.190 2253.600 2442.980 2253.770 ;
        RECT 2440.830 2252.300 2441.005 2253.440 ;
        RECT 2442.190 2252.300 2442.365 2253.600 ;
        RECT 2442.810 2253.560 2442.980 2253.600 ;
        RECT 2443.180 2253.445 2443.350 2253.880 ;
        RECT 2443.180 2252.300 2443.355 2253.445 ;
        RECT 2434.995 2251.945 2436.735 2251.995 ;
        RECT 2434.155 2251.815 2436.735 2251.945 ;
        RECT 2434.155 2251.775 2435.215 2251.815 ;
        RECT 2418.985 2251.145 2419.315 2251.185 ;
        RECT 2419.825 2251.145 2420.645 2251.315 ;
        RECT 2418.985 2250.975 2420.155 2251.145 ;
        RECT 2431.395 2250.975 2431.855 2251.525 ;
        RECT 2432.575 2250.975 2432.880 2251.695 ;
        RECT 2435.355 2251.605 2436.235 2251.645 ;
        RECT 2434.705 2251.405 2436.235 2251.605 ;
        RECT 2434.705 2251.275 2434.875 2251.405 ;
        RECT 2435.625 2251.355 2436.235 2251.405 ;
        RECT 2436.005 2251.315 2436.235 2251.355 ;
        RECT 2436.405 2251.315 2436.735 2251.815 ;
        RECT 2435.565 2251.145 2435.895 2251.185 ;
        RECT 2436.405 2251.145 2437.225 2251.315 ;
        RECT 2435.565 2250.975 2436.735 2251.145 ;
        RECT 2364.815 2250.125 2364.985 2250.465 ;
        RECT 2366.310 2250.125 2366.780 2250.465 ;
        RECT 2364.810 2250.065 2364.985 2250.125 ;
        RECT 2364.300 2249.075 2364.640 2249.955 ;
        RECT 2364.810 2249.245 2364.980 2250.065 ;
        RECT 2365.520 2249.595 2365.770 2249.965 ;
        RECT 2366.490 2249.595 2367.210 2249.895 ;
        RECT 2367.380 2249.765 2367.650 2250.465 ;
        RECT 2368.600 2250.125 2369.080 2250.465 ;
        RECT 2365.520 2249.425 2367.310 2249.595 ;
        RECT 2364.810 2248.995 2365.910 2249.245 ;
        RECT 2364.810 2248.905 2365.060 2248.995 ;
        RECT 2364.760 2248.485 2365.060 2248.905 ;
        RECT 2366.080 2248.575 2366.330 2249.425 ;
        RECT 2365.540 2248.305 2366.330 2248.575 ;
        RECT 2366.500 2248.725 2366.910 2249.245 ;
        RECT 2367.080 2248.995 2367.310 2249.425 ;
        RECT 2367.480 2248.735 2367.650 2249.765 ;
        RECT 2367.820 2249.365 2368.080 2249.815 ;
        RECT 2368.750 2249.635 2369.510 2249.885 ;
        RECT 2369.680 2249.765 2369.950 2250.465 ;
        RECT 2368.740 2249.605 2369.510 2249.635 ;
        RECT 2368.720 2249.595 2369.510 2249.605 ;
        RECT 2368.720 2249.575 2369.610 2249.595 ;
        RECT 2368.700 2249.565 2369.610 2249.575 ;
        RECT 2368.680 2249.555 2369.610 2249.565 ;
        RECT 2368.650 2249.545 2369.610 2249.555 ;
        RECT 2368.580 2249.515 2369.610 2249.545 ;
        RECT 2368.560 2249.485 2369.610 2249.515 ;
        RECT 2368.540 2249.455 2369.610 2249.485 ;
        RECT 2368.510 2249.425 2369.610 2249.455 ;
        RECT 2368.480 2249.395 2369.610 2249.425 ;
        RECT 2368.450 2249.385 2369.610 2249.395 ;
        RECT 2368.450 2249.375 2368.810 2249.385 ;
        RECT 2368.450 2249.365 2368.800 2249.375 ;
        RECT 2367.820 2249.355 2368.780 2249.365 ;
        RECT 2367.820 2249.345 2368.770 2249.355 ;
        RECT 2367.820 2249.325 2368.750 2249.345 ;
        RECT 2367.820 2249.315 2368.740 2249.325 ;
        RECT 2367.820 2249.195 2368.710 2249.315 ;
        RECT 2366.500 2248.305 2366.700 2248.725 ;
        RECT 2367.390 2248.265 2367.650 2248.735 ;
        RECT 2367.820 2248.635 2368.370 2249.025 ;
        RECT 2368.540 2248.465 2368.710 2249.195 ;
        RECT 2367.820 2248.295 2368.710 2248.465 ;
        RECT 2368.880 2248.795 2369.210 2249.215 ;
        RECT 2369.380 2248.995 2369.610 2249.385 ;
        RECT 2369.780 2249.275 2369.950 2249.765 ;
        RECT 2370.130 2249.665 2370.460 2250.455 ;
        RECT 2370.130 2249.495 2370.810 2249.665 ;
        RECT 2370.120 2249.275 2370.470 2249.325 ;
        RECT 2369.780 2249.105 2370.470 2249.275 ;
        RECT 2368.880 2248.305 2369.100 2248.795 ;
        RECT 2369.780 2248.735 2369.950 2249.105 ;
        RECT 2370.120 2249.075 2370.470 2249.105 ;
        RECT 2370.640 2248.895 2370.810 2249.495 ;
        RECT 2370.980 2249.075 2371.330 2249.325 ;
        RECT 2373.110 2248.900 2373.285 2250.160 ;
        RECT 2373.635 2249.100 2373.805 2250.160 ;
        RECT 2373.635 2248.930 2373.865 2249.100 ;
        RECT 2369.690 2248.265 2369.950 2248.735 ;
        RECT 2370.550 2248.265 2370.880 2248.895 ;
        RECT 2373.110 2248.700 2373.280 2248.900 ;
        RECT 2373.110 2248.370 2373.520 2248.700 ;
        RECT 2373.110 2247.860 2373.280 2248.370 ;
        RECT 2373.110 2247.530 2373.520 2247.860 ;
        RECT 2373.110 2247.360 2373.280 2247.530 ;
        RECT 2373.110 2246.870 2373.285 2247.360 ;
        RECT 2373.695 2247.320 2373.865 2248.930 ;
        RECT 2374.065 2248.900 2374.240 2250.160 ;
        RECT 2374.495 2249.020 2374.670 2250.160 ;
        RECT 2374.065 2247.950 2374.235 2248.900 ;
        RECT 2374.495 2247.420 2374.665 2249.020 ;
        RECT 2375.855 2249.015 2376.030 2250.160 ;
        RECT 2376.845 2249.015 2377.020 2250.160 ;
        RECT 2381.400 2250.125 2381.570 2250.465 ;
        RECT 2382.895 2250.125 2383.365 2250.465 ;
        RECT 2381.395 2250.065 2381.570 2250.125 ;
        RECT 2380.885 2249.075 2381.225 2249.955 ;
        RECT 2381.395 2249.245 2381.565 2250.065 ;
        RECT 2382.105 2249.595 2382.355 2249.965 ;
        RECT 2383.075 2249.595 2383.795 2249.895 ;
        RECT 2383.965 2249.765 2384.235 2250.465 ;
        RECT 2385.185 2250.125 2385.665 2250.465 ;
        RECT 2382.105 2249.425 2383.895 2249.595 ;
        RECT 2375.485 2248.210 2375.655 2248.900 ;
        RECT 2375.855 2248.750 2376.025 2249.015 ;
        RECT 2376.475 2248.750 2376.645 2248.900 ;
        RECT 2375.855 2248.580 2376.645 2248.750 ;
        RECT 2376.845 2248.580 2377.015 2249.015 ;
        RECT 2381.395 2248.995 2382.495 2249.245 ;
        RECT 2381.395 2248.905 2381.645 2248.995 ;
        RECT 2376.475 2248.210 2376.645 2248.580 ;
        RECT 2381.345 2248.485 2381.645 2248.905 ;
        RECT 2382.665 2248.575 2382.915 2249.425 ;
        RECT 2382.125 2248.305 2382.915 2248.575 ;
        RECT 2383.085 2248.725 2383.495 2249.245 ;
        RECT 2383.665 2248.995 2383.895 2249.425 ;
        RECT 2384.065 2248.735 2384.235 2249.765 ;
        RECT 2384.405 2249.365 2384.665 2249.815 ;
        RECT 2385.335 2249.635 2386.095 2249.885 ;
        RECT 2386.265 2249.765 2386.535 2250.465 ;
        RECT 2385.325 2249.605 2386.095 2249.635 ;
        RECT 2385.305 2249.595 2386.095 2249.605 ;
        RECT 2385.305 2249.575 2386.195 2249.595 ;
        RECT 2385.285 2249.565 2386.195 2249.575 ;
        RECT 2385.265 2249.555 2386.195 2249.565 ;
        RECT 2385.235 2249.545 2386.195 2249.555 ;
        RECT 2385.165 2249.515 2386.195 2249.545 ;
        RECT 2385.145 2249.485 2386.195 2249.515 ;
        RECT 2385.125 2249.455 2386.195 2249.485 ;
        RECT 2385.095 2249.425 2386.195 2249.455 ;
        RECT 2385.065 2249.395 2386.195 2249.425 ;
        RECT 2385.035 2249.385 2386.195 2249.395 ;
        RECT 2385.035 2249.375 2385.395 2249.385 ;
        RECT 2385.035 2249.365 2385.385 2249.375 ;
        RECT 2384.405 2249.355 2385.365 2249.365 ;
        RECT 2384.405 2249.345 2385.355 2249.355 ;
        RECT 2384.405 2249.325 2385.335 2249.345 ;
        RECT 2384.405 2249.315 2385.325 2249.325 ;
        RECT 2384.405 2249.195 2385.295 2249.315 ;
        RECT 2383.085 2248.305 2383.285 2248.725 ;
        RECT 2383.975 2248.265 2384.235 2248.735 ;
        RECT 2384.405 2248.635 2384.955 2249.025 ;
        RECT 2385.125 2248.465 2385.295 2249.195 ;
        RECT 2384.405 2248.295 2385.295 2248.465 ;
        RECT 2385.465 2248.795 2385.795 2249.215 ;
        RECT 2385.965 2248.995 2386.195 2249.385 ;
        RECT 2386.365 2249.275 2386.535 2249.765 ;
        RECT 2386.715 2249.665 2387.045 2250.455 ;
        RECT 2386.715 2249.495 2387.395 2249.665 ;
        RECT 2386.705 2249.275 2387.055 2249.325 ;
        RECT 2386.365 2249.105 2387.055 2249.275 ;
        RECT 2385.465 2248.305 2385.685 2248.795 ;
        RECT 2386.365 2248.735 2386.535 2249.105 ;
        RECT 2386.705 2249.075 2387.055 2249.105 ;
        RECT 2387.225 2248.895 2387.395 2249.495 ;
        RECT 2387.565 2249.075 2387.915 2249.325 ;
        RECT 2389.695 2248.900 2389.870 2250.160 ;
        RECT 2390.220 2249.100 2390.390 2250.160 ;
        RECT 2390.220 2248.930 2390.450 2249.100 ;
        RECT 2386.275 2248.265 2386.535 2248.735 ;
        RECT 2387.135 2248.265 2387.465 2248.895 ;
        RECT 2389.695 2248.700 2389.865 2248.900 ;
        RECT 2389.695 2248.370 2390.105 2248.700 ;
        RECT 2375.035 2248.040 2375.955 2248.210 ;
        RECT 2376.475 2248.040 2376.945 2248.210 ;
        RECT 2375.035 2247.890 2375.265 2248.040 ;
        RECT 2389.695 2247.860 2389.865 2248.370 ;
        RECT 2389.695 2247.530 2390.105 2247.860 ;
        RECT 2373.635 2247.150 2373.865 2247.320 ;
        RECT 2373.635 2246.870 2373.805 2247.150 ;
        RECT 2374.065 2246.870 2374.240 2247.380 ;
        RECT 2374.495 2246.870 2374.670 2247.420 ;
        RECT 2375.860 2246.870 2376.030 2247.380 ;
        RECT 2376.850 2246.870 2377.020 2247.380 ;
        RECT 2389.695 2247.360 2389.865 2247.530 ;
        RECT 2389.695 2246.870 2389.870 2247.360 ;
        RECT 2390.280 2247.320 2390.450 2248.930 ;
        RECT 2390.650 2248.900 2390.825 2250.160 ;
        RECT 2391.080 2249.020 2391.255 2250.160 ;
        RECT 2390.650 2247.950 2390.820 2248.900 ;
        RECT 2391.080 2247.420 2391.250 2249.020 ;
        RECT 2392.440 2249.015 2392.615 2250.160 ;
        RECT 2393.430 2249.015 2393.605 2250.160 ;
        RECT 2397.985 2250.125 2398.155 2250.465 ;
        RECT 2399.480 2250.125 2399.950 2250.465 ;
        RECT 2397.980 2250.065 2398.155 2250.125 ;
        RECT 2397.470 2249.075 2397.810 2249.955 ;
        RECT 2397.980 2249.245 2398.150 2250.065 ;
        RECT 2398.690 2249.595 2398.940 2249.965 ;
        RECT 2399.660 2249.595 2400.380 2249.895 ;
        RECT 2400.550 2249.765 2400.820 2250.465 ;
        RECT 2401.770 2250.125 2402.250 2250.465 ;
        RECT 2398.690 2249.425 2400.480 2249.595 ;
        RECT 2392.070 2248.210 2392.240 2248.900 ;
        RECT 2392.440 2248.750 2392.610 2249.015 ;
        RECT 2393.060 2248.750 2393.230 2248.900 ;
        RECT 2392.440 2248.580 2393.230 2248.750 ;
        RECT 2393.430 2248.580 2393.600 2249.015 ;
        RECT 2397.980 2248.995 2399.080 2249.245 ;
        RECT 2397.980 2248.905 2398.230 2248.995 ;
        RECT 2393.060 2248.210 2393.230 2248.580 ;
        RECT 2397.930 2248.485 2398.230 2248.905 ;
        RECT 2399.250 2248.575 2399.500 2249.425 ;
        RECT 2398.710 2248.305 2399.500 2248.575 ;
        RECT 2399.670 2248.725 2400.080 2249.245 ;
        RECT 2400.250 2248.995 2400.480 2249.425 ;
        RECT 2400.650 2248.735 2400.820 2249.765 ;
        RECT 2400.990 2249.365 2401.250 2249.815 ;
        RECT 2401.920 2249.635 2402.680 2249.885 ;
        RECT 2402.850 2249.765 2403.120 2250.465 ;
        RECT 2401.910 2249.605 2402.680 2249.635 ;
        RECT 2401.890 2249.595 2402.680 2249.605 ;
        RECT 2401.890 2249.575 2402.780 2249.595 ;
        RECT 2401.870 2249.565 2402.780 2249.575 ;
        RECT 2401.850 2249.555 2402.780 2249.565 ;
        RECT 2401.820 2249.545 2402.780 2249.555 ;
        RECT 2401.750 2249.515 2402.780 2249.545 ;
        RECT 2401.730 2249.485 2402.780 2249.515 ;
        RECT 2401.710 2249.455 2402.780 2249.485 ;
        RECT 2401.680 2249.425 2402.780 2249.455 ;
        RECT 2401.650 2249.395 2402.780 2249.425 ;
        RECT 2401.620 2249.385 2402.780 2249.395 ;
        RECT 2401.620 2249.375 2401.980 2249.385 ;
        RECT 2401.620 2249.365 2401.970 2249.375 ;
        RECT 2400.990 2249.355 2401.950 2249.365 ;
        RECT 2400.990 2249.345 2401.940 2249.355 ;
        RECT 2400.990 2249.325 2401.920 2249.345 ;
        RECT 2400.990 2249.315 2401.910 2249.325 ;
        RECT 2400.990 2249.195 2401.880 2249.315 ;
        RECT 2399.670 2248.305 2399.870 2248.725 ;
        RECT 2400.560 2248.265 2400.820 2248.735 ;
        RECT 2400.990 2248.635 2401.540 2249.025 ;
        RECT 2401.710 2248.465 2401.880 2249.195 ;
        RECT 2400.990 2248.295 2401.880 2248.465 ;
        RECT 2402.050 2248.795 2402.380 2249.215 ;
        RECT 2402.550 2248.995 2402.780 2249.385 ;
        RECT 2402.950 2249.275 2403.120 2249.765 ;
        RECT 2403.300 2249.665 2403.630 2250.455 ;
        RECT 2403.300 2249.495 2403.980 2249.665 ;
        RECT 2403.290 2249.275 2403.640 2249.325 ;
        RECT 2402.950 2249.105 2403.640 2249.275 ;
        RECT 2402.050 2248.305 2402.270 2248.795 ;
        RECT 2402.950 2248.735 2403.120 2249.105 ;
        RECT 2403.290 2249.075 2403.640 2249.105 ;
        RECT 2403.810 2248.895 2403.980 2249.495 ;
        RECT 2404.150 2249.075 2404.500 2249.325 ;
        RECT 2406.280 2248.900 2406.455 2250.160 ;
        RECT 2406.805 2249.100 2406.975 2250.160 ;
        RECT 2406.805 2248.930 2407.035 2249.100 ;
        RECT 2402.860 2248.265 2403.120 2248.735 ;
        RECT 2403.720 2248.265 2404.050 2248.895 ;
        RECT 2406.280 2248.700 2406.450 2248.900 ;
        RECT 2406.280 2248.370 2406.690 2248.700 ;
        RECT 2391.620 2248.040 2392.540 2248.210 ;
        RECT 2393.060 2248.040 2393.530 2248.210 ;
        RECT 2391.620 2247.890 2391.850 2248.040 ;
        RECT 2406.280 2247.860 2406.450 2248.370 ;
        RECT 2406.280 2247.530 2406.690 2247.860 ;
        RECT 2390.220 2247.150 2390.450 2247.320 ;
        RECT 2390.220 2246.870 2390.390 2247.150 ;
        RECT 2390.650 2246.870 2390.825 2247.380 ;
        RECT 2391.080 2246.870 2391.255 2247.420 ;
        RECT 2392.445 2246.870 2392.615 2247.380 ;
        RECT 2393.435 2246.870 2393.605 2247.380 ;
        RECT 2406.280 2247.360 2406.450 2247.530 ;
        RECT 2406.280 2246.870 2406.455 2247.360 ;
        RECT 2406.865 2247.320 2407.035 2248.930 ;
        RECT 2407.235 2248.900 2407.410 2250.160 ;
        RECT 2407.665 2249.020 2407.840 2250.160 ;
        RECT 2407.235 2247.950 2407.405 2248.900 ;
        RECT 2407.665 2247.420 2407.835 2249.020 ;
        RECT 2409.025 2249.015 2409.200 2250.160 ;
        RECT 2410.015 2249.015 2410.190 2250.160 ;
        RECT 2414.570 2250.125 2414.740 2250.465 ;
        RECT 2416.065 2250.125 2416.535 2250.465 ;
        RECT 2414.565 2250.065 2414.740 2250.125 ;
        RECT 2414.055 2249.075 2414.395 2249.955 ;
        RECT 2414.565 2249.245 2414.735 2250.065 ;
        RECT 2415.275 2249.595 2415.525 2249.965 ;
        RECT 2416.245 2249.595 2416.965 2249.895 ;
        RECT 2417.135 2249.765 2417.405 2250.465 ;
        RECT 2418.355 2250.125 2418.835 2250.465 ;
        RECT 2415.275 2249.425 2417.065 2249.595 ;
        RECT 2408.655 2248.210 2408.825 2248.900 ;
        RECT 2409.025 2248.750 2409.195 2249.015 ;
        RECT 2409.645 2248.750 2409.815 2248.900 ;
        RECT 2409.025 2248.580 2409.815 2248.750 ;
        RECT 2410.015 2248.580 2410.185 2249.015 ;
        RECT 2414.565 2248.995 2415.665 2249.245 ;
        RECT 2414.565 2248.905 2414.815 2248.995 ;
        RECT 2409.645 2248.210 2409.815 2248.580 ;
        RECT 2414.515 2248.485 2414.815 2248.905 ;
        RECT 2415.835 2248.575 2416.085 2249.425 ;
        RECT 2415.295 2248.305 2416.085 2248.575 ;
        RECT 2416.255 2248.725 2416.665 2249.245 ;
        RECT 2416.835 2248.995 2417.065 2249.425 ;
        RECT 2417.235 2248.735 2417.405 2249.765 ;
        RECT 2417.575 2249.365 2417.835 2249.815 ;
        RECT 2418.505 2249.635 2419.265 2249.885 ;
        RECT 2419.435 2249.765 2419.705 2250.465 ;
        RECT 2418.495 2249.605 2419.265 2249.635 ;
        RECT 2418.475 2249.595 2419.265 2249.605 ;
        RECT 2418.475 2249.575 2419.365 2249.595 ;
        RECT 2418.455 2249.565 2419.365 2249.575 ;
        RECT 2418.435 2249.555 2419.365 2249.565 ;
        RECT 2418.405 2249.545 2419.365 2249.555 ;
        RECT 2418.335 2249.515 2419.365 2249.545 ;
        RECT 2418.315 2249.485 2419.365 2249.515 ;
        RECT 2418.295 2249.455 2419.365 2249.485 ;
        RECT 2418.265 2249.425 2419.365 2249.455 ;
        RECT 2418.235 2249.395 2419.365 2249.425 ;
        RECT 2418.205 2249.385 2419.365 2249.395 ;
        RECT 2418.205 2249.375 2418.565 2249.385 ;
        RECT 2418.205 2249.365 2418.555 2249.375 ;
        RECT 2417.575 2249.355 2418.535 2249.365 ;
        RECT 2417.575 2249.345 2418.525 2249.355 ;
        RECT 2417.575 2249.325 2418.505 2249.345 ;
        RECT 2417.575 2249.315 2418.495 2249.325 ;
        RECT 2417.575 2249.195 2418.465 2249.315 ;
        RECT 2416.255 2248.305 2416.455 2248.725 ;
        RECT 2417.145 2248.265 2417.405 2248.735 ;
        RECT 2417.575 2248.635 2418.125 2249.025 ;
        RECT 2418.295 2248.465 2418.465 2249.195 ;
        RECT 2417.575 2248.295 2418.465 2248.465 ;
        RECT 2418.635 2248.795 2418.965 2249.215 ;
        RECT 2419.135 2248.995 2419.365 2249.385 ;
        RECT 2419.535 2249.275 2419.705 2249.765 ;
        RECT 2419.885 2249.665 2420.215 2250.455 ;
        RECT 2419.885 2249.495 2420.565 2249.665 ;
        RECT 2419.875 2249.275 2420.225 2249.325 ;
        RECT 2419.535 2249.105 2420.225 2249.275 ;
        RECT 2418.635 2248.305 2418.855 2248.795 ;
        RECT 2419.535 2248.735 2419.705 2249.105 ;
        RECT 2419.875 2249.075 2420.225 2249.105 ;
        RECT 2420.395 2248.895 2420.565 2249.495 ;
        RECT 2420.735 2249.075 2421.085 2249.325 ;
        RECT 2422.865 2248.900 2423.040 2250.160 ;
        RECT 2423.390 2249.100 2423.560 2250.160 ;
        RECT 2423.390 2248.930 2423.620 2249.100 ;
        RECT 2419.445 2248.265 2419.705 2248.735 ;
        RECT 2420.305 2248.265 2420.635 2248.895 ;
        RECT 2422.865 2248.700 2423.035 2248.900 ;
        RECT 2422.865 2248.370 2423.275 2248.700 ;
        RECT 2408.205 2248.040 2409.125 2248.210 ;
        RECT 2409.645 2248.040 2410.115 2248.210 ;
        RECT 2408.205 2247.890 2408.435 2248.040 ;
        RECT 2422.865 2247.860 2423.035 2248.370 ;
        RECT 2422.865 2247.530 2423.275 2247.860 ;
        RECT 2406.805 2247.150 2407.035 2247.320 ;
        RECT 2406.805 2246.870 2406.975 2247.150 ;
        RECT 2407.235 2246.870 2407.410 2247.380 ;
        RECT 2407.665 2246.870 2407.840 2247.420 ;
        RECT 2409.030 2246.870 2409.200 2247.380 ;
        RECT 2410.020 2246.870 2410.190 2247.380 ;
        RECT 2422.865 2247.360 2423.035 2247.530 ;
        RECT 2422.865 2246.870 2423.040 2247.360 ;
        RECT 2423.450 2247.320 2423.620 2248.930 ;
        RECT 2423.820 2248.900 2423.995 2250.160 ;
        RECT 2424.250 2249.020 2424.425 2250.160 ;
        RECT 2423.820 2247.950 2423.990 2248.900 ;
        RECT 2424.250 2247.420 2424.420 2249.020 ;
        RECT 2425.610 2249.015 2425.785 2250.160 ;
        RECT 2426.600 2249.015 2426.775 2250.160 ;
        RECT 2431.150 2250.125 2431.320 2250.465 ;
        RECT 2432.645 2250.125 2433.115 2250.465 ;
        RECT 2431.145 2250.065 2431.320 2250.125 ;
        RECT 2430.635 2249.075 2430.975 2249.955 ;
        RECT 2431.145 2249.245 2431.315 2250.065 ;
        RECT 2431.855 2249.595 2432.105 2249.965 ;
        RECT 2432.825 2249.595 2433.545 2249.895 ;
        RECT 2433.715 2249.765 2433.985 2250.465 ;
        RECT 2434.935 2250.125 2435.415 2250.465 ;
        RECT 2431.855 2249.425 2433.645 2249.595 ;
        RECT 2425.240 2248.210 2425.410 2248.900 ;
        RECT 2425.610 2248.750 2425.780 2249.015 ;
        RECT 2426.230 2248.750 2426.400 2248.900 ;
        RECT 2425.610 2248.580 2426.400 2248.750 ;
        RECT 2426.600 2248.580 2426.770 2249.015 ;
        RECT 2431.145 2248.995 2432.245 2249.245 ;
        RECT 2431.145 2248.905 2431.395 2248.995 ;
        RECT 2426.230 2248.210 2426.400 2248.580 ;
        RECT 2431.095 2248.485 2431.395 2248.905 ;
        RECT 2432.415 2248.575 2432.665 2249.425 ;
        RECT 2431.875 2248.305 2432.665 2248.575 ;
        RECT 2432.835 2248.725 2433.245 2249.245 ;
        RECT 2433.415 2248.995 2433.645 2249.425 ;
        RECT 2433.815 2248.735 2433.985 2249.765 ;
        RECT 2434.155 2249.365 2434.415 2249.815 ;
        RECT 2435.085 2249.635 2435.845 2249.885 ;
        RECT 2436.015 2249.765 2436.285 2250.465 ;
        RECT 2435.075 2249.605 2435.845 2249.635 ;
        RECT 2435.055 2249.595 2435.845 2249.605 ;
        RECT 2435.055 2249.575 2435.945 2249.595 ;
        RECT 2435.035 2249.565 2435.945 2249.575 ;
        RECT 2435.015 2249.555 2435.945 2249.565 ;
        RECT 2434.985 2249.545 2435.945 2249.555 ;
        RECT 2434.915 2249.515 2435.945 2249.545 ;
        RECT 2434.895 2249.485 2435.945 2249.515 ;
        RECT 2434.875 2249.455 2435.945 2249.485 ;
        RECT 2434.845 2249.425 2435.945 2249.455 ;
        RECT 2434.815 2249.395 2435.945 2249.425 ;
        RECT 2434.785 2249.385 2435.945 2249.395 ;
        RECT 2434.785 2249.375 2435.145 2249.385 ;
        RECT 2434.785 2249.365 2435.135 2249.375 ;
        RECT 2434.155 2249.355 2435.115 2249.365 ;
        RECT 2434.155 2249.345 2435.105 2249.355 ;
        RECT 2434.155 2249.325 2435.085 2249.345 ;
        RECT 2434.155 2249.315 2435.075 2249.325 ;
        RECT 2434.155 2249.195 2435.045 2249.315 ;
        RECT 2432.835 2248.305 2433.035 2248.725 ;
        RECT 2433.725 2248.265 2433.985 2248.735 ;
        RECT 2434.155 2248.635 2434.705 2249.025 ;
        RECT 2434.875 2248.465 2435.045 2249.195 ;
        RECT 2434.155 2248.295 2435.045 2248.465 ;
        RECT 2435.215 2248.795 2435.545 2249.215 ;
        RECT 2435.715 2248.995 2435.945 2249.385 ;
        RECT 2436.115 2249.275 2436.285 2249.765 ;
        RECT 2436.465 2249.665 2436.795 2250.455 ;
        RECT 2436.465 2249.495 2437.145 2249.665 ;
        RECT 2436.455 2249.275 2436.805 2249.325 ;
        RECT 2436.115 2249.105 2436.805 2249.275 ;
        RECT 2435.215 2248.305 2435.435 2248.795 ;
        RECT 2436.115 2248.735 2436.285 2249.105 ;
        RECT 2436.455 2249.075 2436.805 2249.105 ;
        RECT 2436.975 2248.895 2437.145 2249.495 ;
        RECT 2437.315 2249.075 2437.665 2249.325 ;
        RECT 2439.445 2248.900 2439.620 2250.160 ;
        RECT 2439.970 2249.100 2440.140 2250.160 ;
        RECT 2439.970 2248.930 2440.200 2249.100 ;
        RECT 2436.025 2248.265 2436.285 2248.735 ;
        RECT 2436.885 2248.265 2437.215 2248.895 ;
        RECT 2439.445 2248.700 2439.615 2248.900 ;
        RECT 2439.445 2248.370 2439.855 2248.700 ;
        RECT 2424.790 2248.040 2425.710 2248.210 ;
        RECT 2426.230 2248.040 2426.700 2248.210 ;
        RECT 2424.790 2247.890 2425.020 2248.040 ;
        RECT 2439.445 2247.860 2439.615 2248.370 ;
        RECT 2439.445 2247.530 2439.855 2247.860 ;
        RECT 2423.390 2247.150 2423.620 2247.320 ;
        RECT 2423.390 2246.870 2423.560 2247.150 ;
        RECT 2423.820 2246.870 2423.995 2247.380 ;
        RECT 2424.250 2246.870 2424.425 2247.420 ;
        RECT 2425.615 2246.870 2425.785 2247.380 ;
        RECT 2426.605 2246.870 2426.775 2247.380 ;
        RECT 2439.445 2247.360 2439.615 2247.530 ;
        RECT 2439.445 2246.870 2439.620 2247.360 ;
        RECT 2440.030 2247.320 2440.200 2248.930 ;
        RECT 2440.400 2248.900 2440.575 2250.160 ;
        RECT 2440.830 2249.020 2441.005 2250.160 ;
        RECT 2440.400 2247.950 2440.570 2248.900 ;
        RECT 2440.830 2247.420 2441.000 2249.020 ;
        RECT 2442.190 2249.015 2442.365 2250.160 ;
        RECT 2443.180 2249.015 2443.355 2250.160 ;
        RECT 2441.820 2248.210 2441.990 2248.900 ;
        RECT 2442.190 2248.750 2442.360 2249.015 ;
        RECT 2442.810 2248.750 2442.980 2248.900 ;
        RECT 2442.190 2248.580 2442.980 2248.750 ;
        RECT 2443.180 2248.580 2443.350 2249.015 ;
        RECT 2442.810 2248.210 2442.980 2248.580 ;
        RECT 2441.370 2248.040 2442.290 2248.210 ;
        RECT 2442.810 2248.040 2443.280 2248.210 ;
        RECT 2441.370 2247.890 2441.600 2248.040 ;
        RECT 2439.970 2247.150 2440.200 2247.320 ;
        RECT 2439.970 2246.870 2440.140 2247.150 ;
        RECT 2440.400 2246.870 2440.575 2247.380 ;
        RECT 2440.830 2246.870 2441.005 2247.420 ;
        RECT 2442.195 2246.870 2442.365 2247.380 ;
        RECT 2443.185 2246.870 2443.355 2247.380 ;
        RECT 2696.985 2216.335 2697.245 2216.665 ;
        RECT 2696.985 2215.425 2697.155 2216.335 ;
        RECT 2697.940 2216.265 2698.145 2216.665 ;
        RECT 2697.940 2216.095 2698.625 2216.265 ;
        RECT 2697.865 2215.425 2698.115 2215.925 ;
        RECT 2696.985 2215.255 2698.115 2215.425 ;
        RECT 2696.985 2214.485 2697.255 2215.255 ;
        RECT 2698.285 2215.065 2698.625 2216.095 ;
        RECT 2697.960 2214.890 2698.625 2215.065 ;
        RECT 2698.825 2216.160 2699.085 2216.665 ;
        RECT 2699.775 2216.285 2699.945 2216.665 ;
        RECT 2698.825 2215.360 2698.995 2216.160 ;
        RECT 2699.280 2216.115 2699.945 2216.285 ;
        RECT 2700.205 2216.160 2700.465 2216.665 ;
        RECT 2701.155 2216.285 2701.325 2216.665 ;
        RECT 2699.280 2215.860 2699.450 2216.115 ;
        RECT 2699.165 2215.530 2699.450 2215.860 ;
        RECT 2699.685 2215.565 2700.015 2215.935 ;
        RECT 2699.280 2215.385 2699.450 2215.530 ;
        RECT 2697.960 2214.485 2698.145 2214.890 ;
        RECT 2698.825 2214.455 2699.095 2215.360 ;
        RECT 2699.280 2215.215 2699.945 2215.385 ;
        RECT 2699.775 2214.455 2699.945 2215.215 ;
        RECT 2700.205 2215.360 2700.375 2216.160 ;
        RECT 2700.660 2216.115 2701.325 2216.285 ;
        RECT 2709.035 2216.285 2709.205 2216.665 ;
        RECT 2709.035 2216.115 2709.750 2216.285 ;
        RECT 2700.660 2215.860 2700.830 2216.115 ;
        RECT 2700.545 2215.530 2700.830 2215.860 ;
        RECT 2701.065 2215.565 2701.395 2215.935 ;
        RECT 2709.580 2215.925 2709.750 2216.115 ;
        RECT 2709.920 2216.090 2710.175 2216.665 ;
        RECT 2722.335 2216.265 2722.540 2216.665 ;
        RECT 2723.235 2216.335 2723.495 2216.665 ;
        RECT 2709.580 2215.595 2709.835 2215.925 ;
        RECT 2700.660 2215.385 2700.830 2215.530 ;
        RECT 2709.580 2215.385 2709.750 2215.595 ;
        RECT 2700.205 2214.455 2700.475 2215.360 ;
        RECT 2700.660 2215.215 2701.325 2215.385 ;
        RECT 2701.155 2214.455 2701.325 2215.215 ;
        RECT 2709.035 2215.215 2709.750 2215.385 ;
        RECT 2710.005 2215.360 2710.175 2216.090 ;
        RECT 2709.035 2214.455 2709.205 2215.215 ;
        RECT 2709.920 2214.455 2710.175 2215.360 ;
        RECT 2721.855 2216.095 2722.540 2216.265 ;
        RECT 2721.855 2215.065 2722.195 2216.095 ;
        RECT 2722.365 2215.425 2722.615 2215.925 ;
        RECT 2723.325 2215.425 2723.495 2216.335 ;
        RECT 2722.365 2215.255 2723.495 2215.425 ;
        RECT 2721.855 2214.890 2722.520 2215.065 ;
        RECT 2722.335 2214.485 2722.520 2214.890 ;
        RECT 2723.225 2214.485 2723.495 2215.255 ;
        RECT 2731.485 2216.160 2731.745 2216.665 ;
        RECT 2732.435 2216.285 2732.605 2216.665 ;
        RECT 2731.485 2215.360 2731.665 2216.160 ;
        RECT 2731.940 2216.115 2732.605 2216.285 ;
        RECT 2731.940 2215.860 2732.110 2216.115 ;
        RECT 2731.835 2215.530 2732.110 2215.860 ;
        RECT 2731.940 2215.385 2732.110 2215.530 ;
        RECT 2731.485 2214.455 2731.755 2215.360 ;
        RECT 2731.940 2215.215 2732.615 2215.385 ;
        RECT 2732.435 2214.455 2732.615 2215.215 ;
        RECT 2697.075 2213.185 2697.245 2213.945 ;
        RECT 2697.075 2213.015 2697.740 2213.185 ;
        RECT 2697.925 2213.040 2698.195 2213.945 ;
        RECT 2697.570 2212.870 2697.740 2213.015 ;
        RECT 2697.005 2212.465 2697.335 2212.835 ;
        RECT 2697.570 2212.540 2697.855 2212.870 ;
        RECT 2697.570 2212.285 2697.740 2212.540 ;
        RECT 2697.075 2212.115 2697.740 2212.285 ;
        RECT 2698.025 2212.240 2698.195 2213.040 ;
        RECT 2697.075 2211.735 2697.245 2212.115 ;
        RECT 2697.935 2211.735 2698.195 2212.240 ;
        RECT 2697.075 2205.405 2697.245 2205.785 ;
        RECT 2697.075 2205.235 2697.740 2205.405 ;
        RECT 2697.935 2205.280 2698.195 2205.785 ;
        RECT 2697.005 2204.685 2697.335 2205.055 ;
        RECT 2697.570 2204.980 2697.740 2205.235 ;
        RECT 2697.570 2204.650 2697.855 2204.980 ;
        RECT 2697.570 2204.505 2697.740 2204.650 ;
        RECT 2697.075 2204.335 2697.740 2204.505 ;
        RECT 2698.025 2204.480 2698.195 2205.280 ;
        RECT 2697.075 2203.575 2697.245 2204.335 ;
        RECT 2697.925 2203.575 2698.195 2204.480 ;
        RECT 2697.075 2199.965 2697.245 2200.340 ;
        RECT 2697.915 2200.175 2698.990 2200.345 ;
        RECT 2697.915 2199.965 2698.085 2200.175 ;
        RECT 2697.075 2199.795 2698.085 2199.965 ;
        RECT 2698.310 2199.835 2698.650 2200.005 ;
        RECT 2698.820 2199.840 2698.990 2200.175 ;
        RECT 2700.280 2200.175 2701.880 2200.345 ;
        RECT 2698.310 2199.665 2698.600 2199.835 ;
        RECT 2697.050 2199.495 2697.395 2199.605 ;
        RECT 2697.045 2199.325 2697.395 2199.495 ;
        RECT 2697.050 2198.985 2697.395 2199.325 ;
        RECT 2697.705 2198.985 2698.140 2199.605 ;
        RECT 2698.310 2199.145 2698.480 2199.665 ;
        RECT 2699.160 2199.495 2699.520 2200.170 ;
        RECT 2700.280 2199.805 2700.450 2200.175 ;
        RECT 2701.525 2200.135 2701.880 2200.175 ;
        RECT 2700.620 2199.755 2700.950 2200.005 ;
        RECT 2700.635 2199.680 2700.950 2199.755 ;
        RECT 2701.120 2199.885 2701.290 2200.005 ;
        RECT 2702.395 2199.885 2702.640 2200.305 ;
        RECT 2703.410 2199.945 2703.585 2200.275 ;
        RECT 2703.930 2200.185 2704.100 2200.345 ;
        RECT 2703.930 2200.015 2704.460 2200.185 ;
        RECT 2704.630 2200.175 2705.625 2200.345 ;
        RECT 2704.630 2200.015 2704.800 2200.175 ;
        RECT 2701.120 2199.715 2702.640 2199.885 ;
        RECT 2698.980 2199.315 2699.520 2199.495 ;
        RECT 2699.160 2199.205 2699.520 2199.315 ;
        RECT 2698.310 2198.975 2698.945 2199.145 ;
        RECT 2699.160 2198.975 2699.965 2199.205 ;
        RECT 2697.075 2198.635 2698.605 2198.805 ;
        RECT 2697.075 2198.135 2697.245 2198.635 ;
        RECT 2698.435 2198.475 2698.605 2198.635 ;
        RECT 2698.775 2198.645 2698.945 2198.975 ;
        RECT 2698.775 2198.475 2699.105 2198.645 ;
        RECT 2697.915 2198.305 2698.085 2198.465 ;
        RECT 2699.275 2198.305 2699.445 2198.805 ;
        RECT 2697.915 2198.135 2699.445 2198.305 ;
        RECT 2699.615 2198.135 2699.965 2198.975 ;
        RECT 2700.165 2198.605 2700.465 2199.605 ;
        RECT 2700.635 2199.155 2700.805 2199.680 ;
        RECT 2701.120 2199.675 2701.290 2199.715 ;
        RECT 2700.975 2199.495 2701.305 2199.505 ;
        RECT 2700.975 2199.335 2701.360 2199.495 ;
        RECT 2701.190 2199.325 2701.360 2199.335 ;
        RECT 2701.700 2199.155 2701.945 2199.545 ;
        RECT 2700.635 2198.985 2701.395 2199.155 ;
        RECT 2701.645 2198.985 2701.945 2199.155 ;
        RECT 2700.725 2198.305 2700.895 2198.815 ;
        RECT 2701.065 2198.475 2701.395 2198.985 ;
        RECT 2701.700 2198.925 2701.945 2198.985 ;
        RECT 2702.150 2198.925 2702.480 2199.545 ;
        RECT 2702.955 2198.925 2703.245 2199.605 ;
        RECT 2703.415 2199.495 2703.585 2199.945 ;
        RECT 2703.880 2199.665 2704.120 2199.835 ;
        RECT 2703.415 2199.325 2703.705 2199.495 ;
        RECT 2701.565 2198.515 2702.630 2198.685 ;
        RECT 2701.565 2198.305 2701.735 2198.515 ;
        RECT 2700.725 2198.135 2701.735 2198.305 ;
        RECT 2702.460 2198.135 2702.630 2198.515 ;
        RECT 2703.415 2198.465 2703.585 2199.325 ;
        RECT 2703.400 2198.135 2703.585 2198.465 ;
        RECT 2703.880 2198.465 2704.050 2199.665 ;
        RECT 2704.290 2198.845 2704.460 2200.015 ;
        RECT 2705.110 2199.835 2705.285 2200.005 ;
        RECT 2704.870 2199.675 2705.285 2199.835 ;
        RECT 2705.455 2199.885 2705.625 2200.175 ;
        RECT 2705.455 2199.715 2706.025 2199.885 ;
        RECT 2704.870 2199.665 2705.280 2199.675 ;
        RECT 2705.090 2199.325 2705.545 2199.495 ;
        RECT 2705.855 2198.935 2706.025 2199.715 ;
        RECT 2704.290 2198.615 2705.075 2198.845 ;
        RECT 2704.745 2198.475 2705.075 2198.615 ;
        RECT 2705.375 2198.765 2706.025 2198.935 ;
        RECT 2703.880 2198.135 2704.090 2198.465 ;
        RECT 2704.260 2198.305 2704.590 2198.345 ;
        RECT 2705.375 2198.305 2705.545 2198.765 ;
        RECT 2704.260 2198.135 2705.545 2198.305 ;
        RECT 2706.215 2198.135 2706.475 2200.345 ;
        RECT 2697.075 2196.865 2697.245 2197.625 ;
        RECT 2697.075 2196.695 2697.740 2196.865 ;
        RECT 2697.925 2196.720 2698.195 2197.625 ;
        RECT 2697.570 2196.550 2697.740 2196.695 ;
        RECT 2697.005 2196.145 2697.335 2196.515 ;
        RECT 2697.570 2196.220 2697.855 2196.550 ;
        RECT 2697.570 2195.965 2697.740 2196.220 ;
        RECT 2697.075 2195.795 2697.740 2195.965 ;
        RECT 2698.025 2195.920 2698.195 2196.720 ;
        RECT 2697.075 2195.415 2697.245 2195.795 ;
        RECT 2697.935 2195.415 2698.195 2195.920 ;
        RECT 2697.075 2194.525 2697.245 2194.900 ;
        RECT 2697.915 2194.735 2698.990 2194.905 ;
        RECT 2697.915 2194.525 2698.085 2194.735 ;
        RECT 2697.075 2194.355 2698.085 2194.525 ;
        RECT 2698.310 2194.395 2698.650 2194.565 ;
        RECT 2698.820 2194.400 2698.990 2194.735 ;
        RECT 2700.280 2194.735 2701.880 2194.905 ;
        RECT 2698.310 2194.225 2698.600 2194.395 ;
        RECT 2697.050 2194.055 2697.395 2194.165 ;
        RECT 2697.045 2193.885 2697.395 2194.055 ;
        RECT 2697.050 2193.545 2697.395 2193.885 ;
        RECT 2697.705 2193.545 2698.140 2194.165 ;
        RECT 2698.310 2193.705 2698.480 2194.225 ;
        RECT 2699.160 2194.055 2699.520 2194.730 ;
        RECT 2700.280 2194.365 2700.450 2194.735 ;
        RECT 2701.525 2194.695 2701.880 2194.735 ;
        RECT 2700.620 2194.315 2700.950 2194.565 ;
        RECT 2700.635 2194.240 2700.950 2194.315 ;
        RECT 2701.120 2194.445 2701.290 2194.565 ;
        RECT 2702.395 2194.445 2702.640 2194.865 ;
        RECT 2703.410 2194.505 2703.585 2194.835 ;
        RECT 2703.930 2194.745 2704.100 2194.905 ;
        RECT 2703.930 2194.575 2704.460 2194.745 ;
        RECT 2704.630 2194.735 2705.625 2194.905 ;
        RECT 2704.630 2194.575 2704.800 2194.735 ;
        RECT 2701.120 2194.275 2702.640 2194.445 ;
        RECT 2698.980 2193.875 2699.520 2194.055 ;
        RECT 2699.160 2193.765 2699.520 2193.875 ;
        RECT 2698.310 2193.535 2698.945 2193.705 ;
        RECT 2699.160 2193.535 2699.965 2193.765 ;
        RECT 2697.075 2193.195 2698.605 2193.365 ;
        RECT 2697.075 2192.695 2697.245 2193.195 ;
        RECT 2698.435 2193.035 2698.605 2193.195 ;
        RECT 2698.775 2193.205 2698.945 2193.535 ;
        RECT 2698.775 2193.035 2699.105 2193.205 ;
        RECT 2697.915 2192.865 2698.085 2193.025 ;
        RECT 2699.275 2192.865 2699.445 2193.365 ;
        RECT 2697.915 2192.695 2699.445 2192.865 ;
        RECT 2699.615 2192.695 2699.965 2193.535 ;
        RECT 2700.165 2193.165 2700.465 2194.165 ;
        RECT 2700.635 2193.715 2700.805 2194.240 ;
        RECT 2701.120 2194.235 2701.290 2194.275 ;
        RECT 2700.975 2194.055 2701.305 2194.065 ;
        RECT 2700.975 2193.895 2701.360 2194.055 ;
        RECT 2701.190 2193.885 2701.360 2193.895 ;
        RECT 2701.700 2193.715 2701.945 2194.105 ;
        RECT 2700.635 2193.545 2701.395 2193.715 ;
        RECT 2701.645 2193.545 2701.945 2193.715 ;
        RECT 2700.725 2192.865 2700.895 2193.375 ;
        RECT 2701.065 2193.035 2701.395 2193.545 ;
        RECT 2701.700 2193.485 2701.945 2193.545 ;
        RECT 2702.150 2193.485 2702.480 2194.105 ;
        RECT 2702.955 2193.485 2703.245 2194.165 ;
        RECT 2703.415 2194.055 2703.585 2194.505 ;
        RECT 2703.880 2194.225 2704.120 2194.395 ;
        RECT 2703.415 2193.885 2703.705 2194.055 ;
        RECT 2701.565 2193.075 2702.630 2193.245 ;
        RECT 2701.565 2192.865 2701.735 2193.075 ;
        RECT 2700.725 2192.695 2701.735 2192.865 ;
        RECT 2702.460 2192.695 2702.630 2193.075 ;
        RECT 2703.415 2193.025 2703.585 2193.885 ;
        RECT 2703.400 2192.695 2703.585 2193.025 ;
        RECT 2703.880 2193.025 2704.050 2194.225 ;
        RECT 2704.290 2193.405 2704.460 2194.575 ;
        RECT 2705.110 2194.395 2705.285 2194.565 ;
        RECT 2704.870 2194.235 2705.285 2194.395 ;
        RECT 2705.455 2194.445 2705.625 2194.735 ;
        RECT 2705.455 2194.275 2706.025 2194.445 ;
        RECT 2704.870 2194.225 2705.280 2194.235 ;
        RECT 2705.090 2193.885 2705.545 2194.055 ;
        RECT 2705.855 2193.495 2706.025 2194.275 ;
        RECT 2704.290 2193.175 2705.075 2193.405 ;
        RECT 2704.745 2193.035 2705.075 2193.175 ;
        RECT 2705.375 2193.325 2706.025 2193.495 ;
        RECT 2703.880 2192.695 2704.090 2193.025 ;
        RECT 2704.260 2192.865 2704.590 2192.905 ;
        RECT 2705.375 2192.865 2705.545 2193.325 ;
        RECT 2704.260 2192.695 2705.545 2192.865 ;
        RECT 2706.215 2192.695 2706.475 2194.905 ;
        RECT 2697.075 2191.425 2697.245 2192.185 ;
        RECT 2697.075 2191.255 2697.740 2191.425 ;
        RECT 2697.925 2191.280 2698.195 2192.185 ;
        RECT 2697.570 2191.110 2697.740 2191.255 ;
        RECT 2697.005 2190.705 2697.335 2191.075 ;
        RECT 2697.570 2190.780 2697.855 2191.110 ;
        RECT 2697.570 2190.525 2697.740 2190.780 ;
        RECT 2697.075 2190.355 2697.740 2190.525 ;
        RECT 2698.025 2190.480 2698.195 2191.280 ;
        RECT 2697.075 2189.975 2697.245 2190.355 ;
        RECT 2697.935 2189.975 2698.195 2190.480 ;
        RECT 2701.590 2191.215 2701.925 2192.185 ;
        RECT 2702.435 2192.015 2704.465 2192.185 ;
        RECT 2701.590 2190.545 2701.760 2191.215 ;
        RECT 2702.435 2191.045 2702.605 2192.015 ;
        RECT 2701.930 2190.715 2702.185 2191.045 ;
        RECT 2702.410 2190.715 2702.605 2191.045 ;
        RECT 2702.775 2191.675 2703.900 2191.845 ;
        RECT 2702.015 2190.545 2702.185 2190.715 ;
        RECT 2702.775 2190.545 2702.945 2191.675 ;
        RECT 2701.590 2189.975 2701.845 2190.545 ;
        RECT 2702.015 2190.375 2702.945 2190.545 ;
        RECT 2703.115 2191.335 2704.125 2191.505 ;
        RECT 2703.115 2190.535 2703.285 2191.335 ;
        RECT 2703.490 2190.655 2703.765 2191.135 ;
        RECT 2703.485 2190.485 2703.765 2190.655 ;
        RECT 2702.770 2190.340 2702.945 2190.375 ;
        RECT 2702.770 2189.975 2703.300 2190.340 ;
        RECT 2703.490 2189.975 2703.765 2190.485 ;
        RECT 2703.935 2189.975 2704.125 2191.335 ;
        RECT 2704.295 2191.350 2704.465 2192.015 ;
        RECT 2705.040 2191.595 2705.555 2192.005 ;
        RECT 2704.295 2191.160 2705.045 2191.350 ;
        RECT 2705.215 2190.785 2705.555 2191.595 ;
        RECT 2704.325 2190.615 2705.555 2190.785 ;
        RECT 2705.035 2190.010 2705.280 2190.615 ;
        RECT 2697.075 2185.985 2697.245 2186.745 ;
        RECT 2697.075 2185.815 2697.740 2185.985 ;
        RECT 2697.925 2185.840 2698.195 2186.745 ;
        RECT 2697.570 2185.670 2697.740 2185.815 ;
        RECT 2697.005 2185.265 2697.335 2185.635 ;
        RECT 2697.570 2185.340 2697.855 2185.670 ;
        RECT 2697.570 2185.085 2697.740 2185.340 ;
        RECT 2697.075 2184.915 2697.740 2185.085 ;
        RECT 2698.025 2185.040 2698.195 2185.840 ;
        RECT 2697.075 2184.535 2697.245 2184.915 ;
        RECT 2697.935 2184.535 2698.195 2185.040 ;
        RECT 2701.595 2180.505 2701.925 2181.290 ;
        RECT 2701.595 2180.335 2702.275 2180.505 ;
        RECT 2701.585 2179.915 2701.935 2180.165 ;
        RECT 2702.105 2179.735 2702.275 2180.335 ;
        RECT 2702.445 2179.915 2702.795 2180.165 ;
        RECT 2702.015 2179.095 2702.345 2179.735 ;
        RECT 2697.075 2178.205 2697.245 2178.585 ;
        RECT 2697.075 2178.035 2697.740 2178.205 ;
        RECT 2697.935 2178.080 2698.195 2178.585 ;
        RECT 2697.005 2177.485 2697.335 2177.855 ;
        RECT 2697.570 2177.780 2697.740 2178.035 ;
        RECT 2697.570 2177.450 2697.855 2177.780 ;
        RECT 2697.570 2177.305 2697.740 2177.450 ;
        RECT 2697.075 2177.135 2697.740 2177.305 ;
        RECT 2698.025 2177.280 2698.195 2178.080 ;
        RECT 2702.565 2178.225 2702.885 2178.585 ;
        RECT 2703.880 2178.225 2704.225 2178.585 ;
        RECT 2702.565 2178.055 2704.225 2178.225 ;
        RECT 2697.075 2176.375 2697.245 2177.135 ;
        RECT 2697.925 2176.375 2698.195 2177.280 ;
        RECT 2702.105 2177.215 2702.380 2177.845 ;
        RECT 2702.090 2176.555 2702.395 2177.045 ;
        RECT 2702.565 2176.725 2702.865 2178.055 ;
        RECT 2703.245 2177.595 2703.575 2177.765 ;
        RECT 2703.250 2177.345 2703.575 2177.595 ;
        RECT 2703.755 2177.515 2704.365 2177.845 ;
        RECT 2704.535 2177.345 2705.035 2177.805 ;
        RECT 2703.250 2177.165 2705.035 2177.345 ;
        RECT 2703.035 2176.815 2705.070 2176.985 ;
        RECT 2703.035 2176.555 2703.365 2176.815 ;
        RECT 2702.090 2176.375 2703.365 2176.555 ;
        RECT 2703.960 2176.735 2705.070 2176.815 ;
        RECT 2703.960 2176.375 2704.130 2176.735 ;
        RECT 2704.810 2176.375 2705.070 2176.735 ;
        RECT 2725.935 2175.015 2726.265 2175.865 ;
        RECT 2726.775 2175.015 2727.105 2175.865 ;
        RECT 2725.935 2174.845 2727.435 2175.015 ;
        RECT 2725.555 2174.475 2727.080 2174.675 ;
        RECT 2727.260 2174.645 2727.435 2174.845 ;
        RECT 2727.260 2174.475 2729.885 2174.645 ;
        RECT 2727.260 2174.305 2727.435 2174.475 ;
        RECT 2726.015 2174.135 2727.435 2174.305 ;
        RECT 2726.015 2173.655 2726.185 2174.135 ;
        RECT 2726.855 2173.660 2727.025 2174.135 ;
        RECT 2697.075 2172.765 2697.245 2173.145 ;
        RECT 2697.075 2172.595 2697.740 2172.765 ;
        RECT 2697.935 2172.640 2698.195 2173.145 ;
        RECT 2697.005 2172.045 2697.335 2172.415 ;
        RECT 2697.570 2172.340 2697.740 2172.595 ;
        RECT 2697.570 2172.010 2697.855 2172.340 ;
        RECT 2697.570 2171.865 2697.740 2172.010 ;
        RECT 2697.075 2171.695 2697.740 2171.865 ;
        RECT 2698.025 2171.840 2698.195 2172.640 ;
        RECT 2697.075 2170.935 2697.245 2171.695 ;
        RECT 2697.925 2170.935 2698.195 2171.840 ;
        RECT 2697.310 2167.305 2697.480 2167.555 ;
        RECT 2696.985 2167.135 2697.480 2167.305 ;
        RECT 2698.215 2167.305 2698.385 2167.650 ;
        RECT 2699.055 2167.305 2699.575 2167.705 ;
        RECT 2698.215 2167.135 2699.575 2167.305 ;
        RECT 2696.985 2166.175 2697.155 2167.135 ;
        RECT 2697.325 2166.345 2697.675 2166.965 ;
        RECT 2697.845 2166.345 2698.185 2166.965 ;
        RECT 2698.355 2166.345 2698.595 2166.965 ;
        RECT 2698.775 2166.715 2699.235 2166.885 ;
        RECT 2698.775 2166.175 2698.945 2166.715 ;
        RECT 2699.405 2166.515 2699.575 2167.135 ;
        RECT 2696.985 2166.005 2698.945 2166.175 ;
        RECT 2699.115 2165.505 2699.575 2166.515 ;
        RECT 2697.075 2164.225 2697.245 2164.985 ;
        RECT 2697.075 2164.055 2697.740 2164.225 ;
        RECT 2697.925 2164.080 2698.195 2164.985 ;
        RECT 2697.570 2163.910 2697.740 2164.055 ;
        RECT 2358.670 2163.105 2358.845 2163.595 ;
        RECT 2359.195 2163.315 2359.365 2163.595 ;
        RECT 2359.195 2163.145 2359.425 2163.315 ;
        RECT 2358.670 2162.935 2358.840 2163.105 ;
        RECT 2358.670 2162.605 2359.080 2162.935 ;
        RECT 2358.670 2162.095 2358.840 2162.605 ;
        RECT 2358.670 2161.765 2359.080 2162.095 ;
        RECT 2358.670 2161.565 2358.840 2161.765 ;
        RECT 2358.670 2160.305 2358.845 2161.565 ;
        RECT 2359.255 2161.535 2359.425 2163.145 ;
        RECT 2359.625 2163.085 2359.800 2163.595 ;
        RECT 2362.080 2163.095 2362.255 2163.585 ;
        RECT 2362.080 2162.925 2362.250 2163.095 ;
        RECT 2363.035 2163.075 2363.210 2163.585 ;
        RECT 2363.465 2163.035 2363.640 2163.585 ;
        RECT 2373.765 2163.105 2373.940 2163.595 ;
        RECT 2374.290 2163.315 2374.460 2163.595 ;
        RECT 2374.290 2163.145 2374.520 2163.315 ;
        RECT 2362.080 2162.595 2362.490 2162.925 ;
        RECT 2359.195 2161.365 2359.425 2161.535 ;
        RECT 2359.625 2161.565 2359.795 2162.515 ;
        RECT 2362.080 2162.085 2362.250 2162.595 ;
        RECT 2362.080 2161.755 2362.490 2162.085 ;
        RECT 2359.195 2160.305 2359.365 2161.365 ;
        RECT 2359.625 2160.305 2359.800 2161.565 ;
        RECT 2362.080 2161.555 2362.250 2161.755 ;
        RECT 2363.035 2161.555 2363.205 2162.505 ;
        RECT 2362.080 2160.295 2362.255 2161.555 ;
        RECT 2363.035 2160.295 2363.210 2161.555 ;
        RECT 2363.465 2161.435 2363.635 2163.035 ;
        RECT 2373.765 2162.935 2373.935 2163.105 ;
        RECT 2373.765 2162.605 2374.175 2162.935 ;
        RECT 2373.765 2162.095 2373.935 2162.605 ;
        RECT 2373.765 2161.765 2374.175 2162.095 ;
        RECT 2373.765 2161.565 2373.935 2161.765 ;
        RECT 2363.465 2160.295 2363.640 2161.435 ;
        RECT 2365.670 2160.560 2366.365 2161.190 ;
        RECT 2365.670 2159.960 2365.840 2160.560 ;
        RECT 2366.010 2160.340 2366.345 2160.370 ;
        RECT 2366.735 2160.340 2366.905 2161.020 ;
        RECT 2366.010 2160.170 2366.905 2160.340 ;
        RECT 2367.970 2160.560 2368.665 2161.190 ;
        RECT 2368.835 2160.560 2369.530 2161.190 ;
        RECT 2370.215 2160.560 2370.910 2161.190 ;
        RECT 2366.010 2160.120 2366.345 2160.170 ;
        RECT 2367.970 2159.960 2368.140 2160.560 ;
        RECT 2368.310 2160.340 2368.645 2160.370 ;
        RECT 2368.855 2160.340 2369.190 2160.370 ;
        RECT 2368.310 2160.170 2369.190 2160.340 ;
        RECT 2368.310 2160.120 2368.645 2160.170 ;
        RECT 2368.855 2160.120 2369.190 2160.170 ;
        RECT 2369.360 2159.960 2369.530 2160.560 ;
        RECT 2369.700 2160.120 2370.035 2160.390 ;
        RECT 2370.235 2160.120 2370.570 2160.370 ;
        RECT 2370.740 2159.960 2370.910 2160.560 ;
        RECT 2371.080 2160.120 2371.415 2160.390 ;
        RECT 2373.765 2160.305 2373.940 2161.565 ;
        RECT 2374.350 2161.535 2374.520 2163.145 ;
        RECT 2374.720 2163.085 2374.895 2163.595 ;
        RECT 2375.150 2163.045 2375.325 2163.595 ;
        RECT 2376.515 2163.085 2376.685 2163.595 ;
        RECT 2377.505 2163.085 2377.675 2163.595 ;
        RECT 2379.300 2163.095 2379.475 2163.585 ;
        RECT 2374.290 2161.365 2374.520 2161.535 ;
        RECT 2374.720 2161.565 2374.890 2162.515 ;
        RECT 2374.290 2160.305 2374.460 2161.365 ;
        RECT 2374.720 2160.305 2374.895 2161.565 ;
        RECT 2375.150 2161.445 2375.320 2163.045 ;
        RECT 2379.300 2162.925 2379.470 2163.095 ;
        RECT 2380.255 2163.075 2380.430 2163.585 ;
        RECT 2380.685 2163.035 2380.860 2163.585 ;
        RECT 2390.985 2163.105 2391.160 2163.595 ;
        RECT 2391.510 2163.315 2391.680 2163.595 ;
        RECT 2391.510 2163.145 2391.740 2163.315 ;
        RECT 2376.080 2162.425 2376.310 2162.610 ;
        RECT 2379.300 2162.595 2379.710 2162.925 ;
        RECT 2376.080 2162.380 2376.610 2162.425 ;
        RECT 2376.140 2162.255 2376.610 2162.380 ;
        RECT 2377.130 2162.255 2377.600 2162.425 ;
        RECT 2376.140 2161.565 2376.310 2162.255 ;
        RECT 2376.510 2161.780 2376.680 2161.885 ;
        RECT 2377.130 2161.780 2377.300 2162.255 ;
        RECT 2379.300 2162.085 2379.470 2162.595 ;
        RECT 2376.510 2161.605 2377.300 2161.780 ;
        RECT 2375.150 2160.305 2375.325 2161.445 ;
        RECT 2376.510 2160.305 2376.685 2161.605 ;
        RECT 2377.130 2161.565 2377.300 2161.605 ;
        RECT 2377.500 2161.450 2377.670 2161.885 ;
        RECT 2379.300 2161.755 2379.710 2162.085 ;
        RECT 2379.300 2161.555 2379.470 2161.755 ;
        RECT 2380.255 2161.555 2380.425 2162.505 ;
        RECT 2377.500 2160.305 2377.675 2161.450 ;
        RECT 2379.300 2160.295 2379.475 2161.555 ;
        RECT 2380.255 2160.295 2380.430 2161.555 ;
        RECT 2380.685 2161.435 2380.855 2163.035 ;
        RECT 2390.985 2162.935 2391.155 2163.105 ;
        RECT 2390.985 2162.605 2391.395 2162.935 ;
        RECT 2390.985 2162.095 2391.155 2162.605 ;
        RECT 2390.985 2161.765 2391.395 2162.095 ;
        RECT 2390.985 2161.565 2391.155 2161.765 ;
        RECT 2380.685 2160.295 2380.860 2161.435 ;
        RECT 2382.890 2160.560 2383.585 2161.190 ;
        RECT 2382.890 2159.960 2383.060 2160.560 ;
        RECT 2383.230 2160.340 2383.565 2160.370 ;
        RECT 2383.955 2160.340 2384.125 2161.020 ;
        RECT 2383.230 2160.170 2384.125 2160.340 ;
        RECT 2385.190 2160.560 2385.885 2161.190 ;
        RECT 2386.055 2160.560 2386.750 2161.190 ;
        RECT 2387.435 2160.560 2388.130 2161.190 ;
        RECT 2383.230 2160.120 2383.565 2160.170 ;
        RECT 2385.190 2159.960 2385.360 2160.560 ;
        RECT 2385.530 2160.340 2385.865 2160.370 ;
        RECT 2386.075 2160.340 2386.410 2160.370 ;
        RECT 2385.530 2160.170 2386.410 2160.340 ;
        RECT 2385.530 2160.120 2385.865 2160.170 ;
        RECT 2386.075 2160.120 2386.410 2160.170 ;
        RECT 2386.580 2159.960 2386.750 2160.560 ;
        RECT 2386.920 2160.120 2387.255 2160.390 ;
        RECT 2387.455 2160.120 2387.790 2160.370 ;
        RECT 2387.960 2159.960 2388.130 2160.560 ;
        RECT 2388.300 2160.120 2388.635 2160.390 ;
        RECT 2390.985 2160.305 2391.160 2161.565 ;
        RECT 2391.570 2161.535 2391.740 2163.145 ;
        RECT 2391.940 2163.085 2392.115 2163.595 ;
        RECT 2392.370 2163.045 2392.545 2163.595 ;
        RECT 2393.735 2163.085 2393.905 2163.595 ;
        RECT 2394.725 2163.085 2394.895 2163.595 ;
        RECT 2396.520 2163.095 2396.695 2163.585 ;
        RECT 2391.510 2161.365 2391.740 2161.535 ;
        RECT 2391.940 2161.565 2392.110 2162.515 ;
        RECT 2391.510 2160.305 2391.680 2161.365 ;
        RECT 2391.940 2160.305 2392.115 2161.565 ;
        RECT 2392.370 2161.445 2392.540 2163.045 ;
        RECT 2396.520 2162.925 2396.690 2163.095 ;
        RECT 2397.475 2163.075 2397.650 2163.585 ;
        RECT 2397.905 2163.035 2398.080 2163.585 ;
        RECT 2408.205 2163.105 2408.380 2163.595 ;
        RECT 2408.730 2163.315 2408.900 2163.595 ;
        RECT 2408.730 2163.145 2408.960 2163.315 ;
        RECT 2393.300 2162.425 2393.530 2162.610 ;
        RECT 2396.520 2162.595 2396.930 2162.925 ;
        RECT 2393.300 2162.380 2393.830 2162.425 ;
        RECT 2393.360 2162.255 2393.830 2162.380 ;
        RECT 2394.350 2162.255 2394.820 2162.425 ;
        RECT 2393.360 2161.565 2393.530 2162.255 ;
        RECT 2393.730 2161.780 2393.900 2161.885 ;
        RECT 2394.350 2161.780 2394.520 2162.255 ;
        RECT 2396.520 2162.085 2396.690 2162.595 ;
        RECT 2393.730 2161.605 2394.520 2161.780 ;
        RECT 2392.370 2160.305 2392.545 2161.445 ;
        RECT 2393.730 2160.305 2393.905 2161.605 ;
        RECT 2394.350 2161.565 2394.520 2161.605 ;
        RECT 2394.720 2161.450 2394.890 2161.885 ;
        RECT 2396.520 2161.755 2396.930 2162.085 ;
        RECT 2396.520 2161.555 2396.690 2161.755 ;
        RECT 2397.475 2161.555 2397.645 2162.505 ;
        RECT 2394.720 2160.305 2394.895 2161.450 ;
        RECT 2396.520 2160.295 2396.695 2161.555 ;
        RECT 2397.475 2160.295 2397.650 2161.555 ;
        RECT 2397.905 2161.435 2398.075 2163.035 ;
        RECT 2408.205 2162.935 2408.375 2163.105 ;
        RECT 2408.205 2162.605 2408.615 2162.935 ;
        RECT 2408.205 2162.095 2408.375 2162.605 ;
        RECT 2408.205 2161.765 2408.615 2162.095 ;
        RECT 2408.205 2161.565 2408.375 2161.765 ;
        RECT 2397.905 2160.295 2398.080 2161.435 ;
        RECT 2400.110 2160.560 2400.805 2161.190 ;
        RECT 2400.110 2159.960 2400.280 2160.560 ;
        RECT 2400.450 2160.340 2400.785 2160.370 ;
        RECT 2401.175 2160.340 2401.345 2161.020 ;
        RECT 2400.450 2160.170 2401.345 2160.340 ;
        RECT 2402.410 2160.560 2403.105 2161.190 ;
        RECT 2403.275 2160.560 2403.970 2161.190 ;
        RECT 2404.655 2160.560 2405.350 2161.190 ;
        RECT 2400.450 2160.120 2400.785 2160.170 ;
        RECT 2402.410 2159.960 2402.580 2160.560 ;
        RECT 2402.750 2160.340 2403.085 2160.370 ;
        RECT 2403.295 2160.340 2403.630 2160.370 ;
        RECT 2402.750 2160.170 2403.630 2160.340 ;
        RECT 2402.750 2160.120 2403.085 2160.170 ;
        RECT 2403.295 2160.120 2403.630 2160.170 ;
        RECT 2403.800 2159.960 2403.970 2160.560 ;
        RECT 2404.140 2160.120 2404.475 2160.390 ;
        RECT 2404.675 2160.120 2405.010 2160.370 ;
        RECT 2405.180 2159.960 2405.350 2160.560 ;
        RECT 2405.520 2160.120 2405.855 2160.390 ;
        RECT 2408.205 2160.305 2408.380 2161.565 ;
        RECT 2408.790 2161.535 2408.960 2163.145 ;
        RECT 2409.160 2163.085 2409.335 2163.595 ;
        RECT 2409.590 2163.045 2409.765 2163.595 ;
        RECT 2410.955 2163.085 2411.125 2163.595 ;
        RECT 2411.945 2163.085 2412.115 2163.595 ;
        RECT 2413.740 2163.095 2413.915 2163.585 ;
        RECT 2408.730 2161.365 2408.960 2161.535 ;
        RECT 2409.160 2161.565 2409.330 2162.515 ;
        RECT 2408.730 2160.305 2408.900 2161.365 ;
        RECT 2409.160 2160.305 2409.335 2161.565 ;
        RECT 2409.590 2161.445 2409.760 2163.045 ;
        RECT 2413.740 2162.925 2413.910 2163.095 ;
        RECT 2414.695 2163.075 2414.870 2163.585 ;
        RECT 2415.125 2163.035 2415.300 2163.585 ;
        RECT 2425.425 2163.105 2425.600 2163.595 ;
        RECT 2425.950 2163.315 2426.120 2163.595 ;
        RECT 2425.950 2163.145 2426.180 2163.315 ;
        RECT 2410.520 2162.425 2410.750 2162.610 ;
        RECT 2413.740 2162.595 2414.150 2162.925 ;
        RECT 2410.520 2162.380 2411.050 2162.425 ;
        RECT 2410.580 2162.255 2411.050 2162.380 ;
        RECT 2411.570 2162.255 2412.040 2162.425 ;
        RECT 2410.580 2161.565 2410.750 2162.255 ;
        RECT 2410.950 2161.780 2411.120 2161.885 ;
        RECT 2411.570 2161.780 2411.740 2162.255 ;
        RECT 2413.740 2162.085 2413.910 2162.595 ;
        RECT 2410.950 2161.605 2411.740 2161.780 ;
        RECT 2409.590 2160.305 2409.765 2161.445 ;
        RECT 2410.950 2160.305 2411.125 2161.605 ;
        RECT 2411.570 2161.565 2411.740 2161.605 ;
        RECT 2411.940 2161.450 2412.110 2161.885 ;
        RECT 2413.740 2161.755 2414.150 2162.085 ;
        RECT 2413.740 2161.555 2413.910 2161.755 ;
        RECT 2414.695 2161.555 2414.865 2162.505 ;
        RECT 2411.940 2160.305 2412.115 2161.450 ;
        RECT 2413.740 2160.295 2413.915 2161.555 ;
        RECT 2414.695 2160.295 2414.870 2161.555 ;
        RECT 2415.125 2161.435 2415.295 2163.035 ;
        RECT 2425.425 2162.935 2425.595 2163.105 ;
        RECT 2425.425 2162.605 2425.835 2162.935 ;
        RECT 2425.425 2162.095 2425.595 2162.605 ;
        RECT 2425.425 2161.765 2425.835 2162.095 ;
        RECT 2425.425 2161.565 2425.595 2161.765 ;
        RECT 2415.125 2160.295 2415.300 2161.435 ;
        RECT 2417.330 2160.560 2418.025 2161.190 ;
        RECT 2417.330 2159.960 2417.500 2160.560 ;
        RECT 2417.670 2160.340 2418.005 2160.370 ;
        RECT 2418.395 2160.340 2418.565 2161.020 ;
        RECT 2417.670 2160.170 2418.565 2160.340 ;
        RECT 2419.630 2160.560 2420.325 2161.190 ;
        RECT 2420.495 2160.560 2421.190 2161.190 ;
        RECT 2421.875 2160.560 2422.570 2161.190 ;
        RECT 2417.670 2160.120 2418.005 2160.170 ;
        RECT 2419.630 2159.960 2419.800 2160.560 ;
        RECT 2419.970 2160.340 2420.305 2160.370 ;
        RECT 2420.515 2160.340 2420.850 2160.370 ;
        RECT 2419.970 2160.170 2420.850 2160.340 ;
        RECT 2419.970 2160.120 2420.305 2160.170 ;
        RECT 2420.515 2160.120 2420.850 2160.170 ;
        RECT 2421.020 2159.960 2421.190 2160.560 ;
        RECT 2421.360 2160.120 2421.695 2160.390 ;
        RECT 2421.895 2160.120 2422.230 2160.370 ;
        RECT 2422.400 2159.960 2422.570 2160.560 ;
        RECT 2422.740 2160.120 2423.075 2160.390 ;
        RECT 2425.425 2160.305 2425.600 2161.565 ;
        RECT 2426.010 2161.535 2426.180 2163.145 ;
        RECT 2426.380 2163.085 2426.555 2163.595 ;
        RECT 2426.810 2163.045 2426.985 2163.595 ;
        RECT 2428.175 2163.085 2428.345 2163.595 ;
        RECT 2429.165 2163.085 2429.335 2163.595 ;
        RECT 2430.960 2163.095 2431.135 2163.585 ;
        RECT 2425.950 2161.365 2426.180 2161.535 ;
        RECT 2426.380 2161.565 2426.550 2162.515 ;
        RECT 2425.950 2160.305 2426.120 2161.365 ;
        RECT 2426.380 2160.305 2426.555 2161.565 ;
        RECT 2426.810 2161.445 2426.980 2163.045 ;
        RECT 2430.960 2162.925 2431.130 2163.095 ;
        RECT 2431.915 2163.075 2432.090 2163.585 ;
        RECT 2432.345 2163.035 2432.520 2163.585 ;
        RECT 2442.645 2163.105 2442.820 2163.595 ;
        RECT 2443.170 2163.315 2443.340 2163.595 ;
        RECT 2443.170 2163.145 2443.400 2163.315 ;
        RECT 2427.740 2162.425 2427.970 2162.610 ;
        RECT 2430.960 2162.595 2431.370 2162.925 ;
        RECT 2427.740 2162.380 2428.270 2162.425 ;
        RECT 2427.800 2162.255 2428.270 2162.380 ;
        RECT 2428.790 2162.255 2429.260 2162.425 ;
        RECT 2427.800 2161.565 2427.970 2162.255 ;
        RECT 2428.170 2161.780 2428.340 2161.885 ;
        RECT 2428.790 2161.780 2428.960 2162.255 ;
        RECT 2430.960 2162.085 2431.130 2162.595 ;
        RECT 2428.170 2161.605 2428.960 2161.780 ;
        RECT 2426.810 2160.305 2426.985 2161.445 ;
        RECT 2428.170 2160.305 2428.345 2161.605 ;
        RECT 2428.790 2161.565 2428.960 2161.605 ;
        RECT 2429.160 2161.450 2429.330 2161.885 ;
        RECT 2430.960 2161.755 2431.370 2162.085 ;
        RECT 2430.960 2161.555 2431.130 2161.755 ;
        RECT 2431.915 2161.555 2432.085 2162.505 ;
        RECT 2429.160 2160.305 2429.335 2161.450 ;
        RECT 2430.960 2160.295 2431.135 2161.555 ;
        RECT 2431.915 2160.295 2432.090 2161.555 ;
        RECT 2432.345 2161.435 2432.515 2163.035 ;
        RECT 2442.645 2162.935 2442.815 2163.105 ;
        RECT 2442.645 2162.605 2443.055 2162.935 ;
        RECT 2442.645 2162.095 2442.815 2162.605 ;
        RECT 2442.645 2161.765 2443.055 2162.095 ;
        RECT 2442.645 2161.565 2442.815 2161.765 ;
        RECT 2432.345 2160.295 2432.520 2161.435 ;
        RECT 2434.550 2160.560 2435.245 2161.190 ;
        RECT 2434.550 2159.960 2434.720 2160.560 ;
        RECT 2434.890 2160.340 2435.225 2160.370 ;
        RECT 2435.615 2160.340 2435.785 2161.020 ;
        RECT 2434.890 2160.170 2435.785 2160.340 ;
        RECT 2436.850 2160.560 2437.545 2161.190 ;
        RECT 2437.715 2160.560 2438.410 2161.190 ;
        RECT 2439.095 2160.560 2439.790 2161.190 ;
        RECT 2434.890 2160.120 2435.225 2160.170 ;
        RECT 2436.850 2159.960 2437.020 2160.560 ;
        RECT 2437.190 2160.340 2437.525 2160.370 ;
        RECT 2437.735 2160.340 2438.070 2160.370 ;
        RECT 2437.190 2160.170 2438.070 2160.340 ;
        RECT 2437.190 2160.120 2437.525 2160.170 ;
        RECT 2437.735 2160.120 2438.070 2160.170 ;
        RECT 2438.240 2159.960 2438.410 2160.560 ;
        RECT 2438.580 2160.120 2438.915 2160.390 ;
        RECT 2439.115 2160.120 2439.450 2160.370 ;
        RECT 2439.620 2159.960 2439.790 2160.560 ;
        RECT 2439.960 2160.120 2440.295 2160.390 ;
        RECT 2442.645 2160.305 2442.820 2161.565 ;
        RECT 2443.230 2161.535 2443.400 2163.145 ;
        RECT 2443.600 2163.085 2443.775 2163.595 ;
        RECT 2444.030 2163.045 2444.205 2163.595 ;
        RECT 2445.395 2163.085 2445.565 2163.595 ;
        RECT 2446.385 2163.085 2446.555 2163.595 ;
        RECT 2697.005 2163.505 2697.335 2163.875 ;
        RECT 2697.570 2163.580 2697.855 2163.910 ;
        RECT 2697.570 2163.325 2697.740 2163.580 ;
        RECT 2697.075 2163.155 2697.740 2163.325 ;
        RECT 2698.025 2163.280 2698.195 2164.080 ;
        RECT 2443.170 2161.365 2443.400 2161.535 ;
        RECT 2443.600 2161.565 2443.770 2162.515 ;
        RECT 2443.170 2160.305 2443.340 2161.365 ;
        RECT 2443.600 2160.305 2443.775 2161.565 ;
        RECT 2444.030 2161.445 2444.200 2163.045 ;
        RECT 2697.075 2162.775 2697.245 2163.155 ;
        RECT 2697.935 2162.775 2698.195 2163.280 ;
        RECT 2444.960 2162.425 2445.190 2162.610 ;
        RECT 2444.960 2162.380 2445.490 2162.425 ;
        RECT 2445.020 2162.255 2445.490 2162.380 ;
        RECT 2446.010 2162.255 2446.480 2162.425 ;
        RECT 2445.020 2161.565 2445.190 2162.255 ;
        RECT 2445.390 2161.780 2445.560 2161.885 ;
        RECT 2446.010 2161.780 2446.180 2162.255 ;
        RECT 2445.390 2161.605 2446.180 2161.780 ;
        RECT 2444.030 2160.305 2444.205 2161.445 ;
        RECT 2445.390 2160.305 2445.565 2161.605 ;
        RECT 2446.010 2161.565 2446.180 2161.605 ;
        RECT 2446.380 2161.450 2446.550 2161.885 ;
        RECT 2697.260 2161.625 2697.505 2162.230 ;
        RECT 2696.985 2161.455 2698.215 2161.625 ;
        RECT 2446.380 2160.305 2446.555 2161.450 ;
        RECT 2696.985 2160.645 2697.325 2161.455 ;
        RECT 2697.495 2160.890 2698.245 2161.080 ;
        RECT 2696.985 2160.235 2697.500 2160.645 ;
        RECT 2698.075 2160.225 2698.245 2160.890 ;
        RECT 2698.415 2160.905 2698.605 2162.265 ;
        RECT 2698.775 2162.095 2699.050 2162.265 ;
        RECT 2698.775 2161.925 2699.055 2162.095 ;
        RECT 2698.775 2161.105 2699.050 2161.925 ;
        RECT 2699.240 2161.900 2699.770 2162.265 ;
        RECT 2699.595 2161.865 2699.770 2161.900 ;
        RECT 2699.255 2160.905 2699.425 2161.705 ;
        RECT 2698.415 2160.735 2699.425 2160.905 ;
        RECT 2699.595 2161.695 2700.525 2161.865 ;
        RECT 2700.695 2161.695 2700.950 2162.265 ;
        RECT 2699.595 2160.565 2699.765 2161.695 ;
        RECT 2700.355 2161.525 2700.525 2161.695 ;
        RECT 2698.640 2160.395 2699.765 2160.565 ;
        RECT 2699.935 2161.195 2700.130 2161.525 ;
        RECT 2700.355 2161.195 2700.610 2161.525 ;
        RECT 2699.935 2160.225 2700.105 2161.195 ;
        RECT 2700.780 2161.025 2700.950 2161.695 ;
        RECT 2701.630 2161.500 2701.815 2162.170 ;
        RECT 2702.300 2161.815 2702.630 2162.215 ;
        RECT 2703.345 2161.820 2703.675 2162.260 ;
        RECT 2703.345 2161.815 2704.575 2161.820 ;
        RECT 2702.300 2161.705 2704.575 2161.815 ;
        RECT 2702.420 2161.640 2704.575 2161.705 ;
        RECT 2701.180 2161.230 2701.815 2161.500 ;
        RECT 2701.995 2161.120 2702.280 2161.525 ;
        RECT 2702.450 2161.120 2702.780 2161.470 ;
        RECT 2698.075 2160.055 2700.105 2160.225 ;
        RECT 2700.615 2160.055 2700.950 2161.025 ;
        RECT 2701.215 2160.770 2702.325 2160.940 ;
        RECT 2701.215 2160.060 2701.410 2160.770 ;
        RECT 2702.095 2160.060 2702.325 2160.770 ;
        RECT 2702.505 2160.065 2702.780 2161.120 ;
        RECT 2702.950 2160.065 2703.285 2161.470 ;
        RECT 2703.485 2160.065 2703.935 2161.470 ;
        RECT 2704.190 2160.060 2704.575 2161.640 ;
        RECT 2365.605 2158.980 2365.935 2159.960 ;
        RECT 2367.905 2158.980 2368.235 2159.960 ;
        RECT 2369.265 2158.980 2369.595 2159.960 ;
        RECT 2370.645 2158.980 2370.975 2159.960 ;
        RECT 2382.825 2158.980 2383.155 2159.960 ;
        RECT 2385.125 2158.980 2385.455 2159.960 ;
        RECT 2386.485 2158.980 2386.815 2159.960 ;
        RECT 2387.865 2158.980 2388.195 2159.960 ;
        RECT 2400.045 2158.980 2400.375 2159.960 ;
        RECT 2402.345 2158.980 2402.675 2159.960 ;
        RECT 2403.705 2158.980 2404.035 2159.960 ;
        RECT 2405.085 2158.980 2405.415 2159.960 ;
        RECT 2417.265 2158.980 2417.595 2159.960 ;
        RECT 2419.565 2158.980 2419.895 2159.960 ;
        RECT 2420.925 2158.980 2421.255 2159.960 ;
        RECT 2422.305 2158.980 2422.635 2159.960 ;
        RECT 2434.485 2158.980 2434.815 2159.960 ;
        RECT 2436.785 2158.980 2437.115 2159.960 ;
        RECT 2438.145 2158.980 2438.475 2159.960 ;
        RECT 2439.525 2158.980 2439.855 2159.960 ;
        RECT 2365.135 2157.490 2365.465 2158.470 ;
        RECT 2366.945 2157.670 2367.275 2158.455 ;
        RECT 2366.595 2157.500 2367.275 2157.670 ;
        RECT 2367.465 2157.670 2367.795 2158.455 ;
        RECT 2367.465 2157.500 2368.145 2157.670 ;
        RECT 2365.135 2156.890 2365.385 2157.490 ;
        RECT 2365.555 2157.280 2365.885 2157.330 ;
        RECT 2366.075 2157.280 2366.425 2157.330 ;
        RECT 2365.555 2157.110 2366.425 2157.280 ;
        RECT 2365.555 2157.080 2365.885 2157.110 ;
        RECT 2366.075 2157.080 2366.425 2157.110 ;
        RECT 2366.595 2156.900 2366.765 2157.500 ;
        RECT 2366.935 2157.080 2367.285 2157.330 ;
        RECT 2367.455 2157.080 2367.805 2157.330 ;
        RECT 2367.975 2156.900 2368.145 2157.500 ;
        RECT 2368.835 2157.620 2369.155 2158.470 ;
        RECT 2369.335 2157.960 2369.735 2158.470 ;
        RECT 2370.245 2157.960 2370.575 2158.470 ;
        RECT 2369.335 2157.790 2370.575 2157.960 ;
        RECT 2371.155 2157.620 2371.325 2158.300 ;
        RECT 2371.505 2157.790 2371.885 2158.470 ;
        RECT 2368.835 2157.540 2369.285 2157.620 ;
        RECT 2368.835 2157.370 2369.465 2157.540 ;
        RECT 2368.315 2157.080 2368.665 2157.330 ;
        RECT 2365.135 2156.260 2365.465 2156.890 ;
        RECT 2366.525 2156.260 2366.855 2156.900 ;
        RECT 2367.885 2156.260 2368.215 2156.900 ;
        RECT 2369.295 2156.490 2369.465 2157.370 ;
        RECT 2370.240 2157.450 2371.545 2157.620 ;
        RECT 2369.635 2156.830 2369.865 2157.330 ;
        RECT 2370.240 2157.250 2370.410 2157.450 ;
        RECT 2370.035 2157.080 2370.410 2157.250 ;
        RECT 2370.580 2157.080 2371.130 2157.280 ;
        RECT 2371.300 2157.000 2371.545 2157.450 ;
        RECT 2371.715 2156.830 2371.885 2157.790 ;
        RECT 2369.635 2156.660 2371.885 2156.830 ;
        RECT 2373.765 2156.895 2373.940 2158.155 ;
        RECT 2374.290 2157.095 2374.460 2158.155 ;
        RECT 2374.290 2156.925 2374.520 2157.095 ;
        RECT 2373.765 2156.695 2373.935 2156.895 ;
        RECT 2369.295 2156.320 2370.250 2156.490 ;
        RECT 2371.165 2156.340 2371.335 2156.660 ;
        RECT 2373.765 2156.365 2374.175 2156.695 ;
        RECT 2373.765 2155.855 2373.935 2156.365 ;
        RECT 2373.765 2155.525 2374.175 2155.855 ;
        RECT 2373.765 2155.355 2373.935 2155.525 ;
        RECT 2373.765 2154.865 2373.940 2155.355 ;
        RECT 2374.350 2155.315 2374.520 2156.925 ;
        RECT 2374.720 2156.895 2374.895 2158.155 ;
        RECT 2375.150 2157.015 2375.325 2158.155 ;
        RECT 2374.720 2155.945 2374.890 2156.895 ;
        RECT 2375.150 2155.415 2375.320 2157.015 ;
        RECT 2376.510 2157.010 2376.685 2158.155 ;
        RECT 2377.495 2157.010 2377.670 2158.155 ;
        RECT 2382.355 2157.490 2382.685 2158.470 ;
        RECT 2384.165 2157.670 2384.495 2158.455 ;
        RECT 2383.815 2157.500 2384.495 2157.670 ;
        RECT 2384.685 2157.670 2385.015 2158.455 ;
        RECT 2384.685 2157.500 2385.365 2157.670 ;
        RECT 2376.140 2156.205 2376.310 2156.895 ;
        RECT 2376.510 2156.805 2376.680 2157.010 ;
        RECT 2377.125 2156.805 2377.295 2156.895 ;
        RECT 2376.510 2156.625 2377.295 2156.805 ;
        RECT 2376.510 2156.575 2376.680 2156.625 ;
        RECT 2377.125 2156.205 2377.295 2156.625 ;
        RECT 2377.495 2156.575 2377.665 2157.010 ;
        RECT 2382.355 2156.890 2382.605 2157.490 ;
        RECT 2382.775 2157.280 2383.105 2157.330 ;
        RECT 2383.295 2157.280 2383.645 2157.330 ;
        RECT 2382.775 2157.110 2383.645 2157.280 ;
        RECT 2382.775 2157.080 2383.105 2157.110 ;
        RECT 2383.295 2157.080 2383.645 2157.110 ;
        RECT 2383.815 2156.900 2383.985 2157.500 ;
        RECT 2384.155 2157.080 2384.505 2157.330 ;
        RECT 2384.675 2157.080 2385.025 2157.330 ;
        RECT 2385.195 2156.900 2385.365 2157.500 ;
        RECT 2386.055 2157.620 2386.375 2158.470 ;
        RECT 2386.555 2157.960 2386.955 2158.470 ;
        RECT 2387.465 2157.960 2387.795 2158.470 ;
        RECT 2386.555 2157.790 2387.795 2157.960 ;
        RECT 2388.375 2157.620 2388.545 2158.300 ;
        RECT 2388.725 2157.790 2389.105 2158.470 ;
        RECT 2386.055 2157.540 2386.505 2157.620 ;
        RECT 2386.055 2157.370 2386.685 2157.540 ;
        RECT 2385.535 2157.080 2385.885 2157.330 ;
        RECT 2382.355 2156.260 2382.685 2156.890 ;
        RECT 2383.745 2156.260 2384.075 2156.900 ;
        RECT 2385.105 2156.260 2385.435 2156.900 ;
        RECT 2386.515 2156.490 2386.685 2157.370 ;
        RECT 2387.460 2157.450 2388.765 2157.620 ;
        RECT 2386.855 2156.830 2387.085 2157.330 ;
        RECT 2387.460 2157.250 2387.630 2157.450 ;
        RECT 2387.255 2157.080 2387.630 2157.250 ;
        RECT 2387.800 2157.080 2388.350 2157.280 ;
        RECT 2388.520 2157.000 2388.765 2157.450 ;
        RECT 2388.935 2156.830 2389.105 2157.790 ;
        RECT 2386.855 2156.660 2389.105 2156.830 ;
        RECT 2390.985 2156.895 2391.160 2158.155 ;
        RECT 2391.510 2157.095 2391.680 2158.155 ;
        RECT 2391.510 2156.925 2391.740 2157.095 ;
        RECT 2390.985 2156.695 2391.155 2156.895 ;
        RECT 2386.515 2156.320 2387.470 2156.490 ;
        RECT 2388.385 2156.340 2388.555 2156.660 ;
        RECT 2390.985 2156.365 2391.395 2156.695 ;
        RECT 2376.140 2156.175 2376.610 2156.205 ;
        RECT 2376.095 2156.035 2376.610 2156.175 ;
        RECT 2377.125 2156.035 2377.595 2156.205 ;
        RECT 2376.095 2155.945 2376.325 2156.035 ;
        RECT 2390.985 2155.855 2391.155 2156.365 ;
        RECT 2390.985 2155.525 2391.395 2155.855 ;
        RECT 2374.290 2155.145 2374.520 2155.315 ;
        RECT 2374.290 2154.865 2374.460 2155.145 ;
        RECT 2374.720 2154.865 2374.895 2155.375 ;
        RECT 2375.150 2154.865 2375.325 2155.415 ;
        RECT 2376.515 2154.865 2376.685 2155.375 ;
        RECT 2377.500 2154.865 2377.670 2155.375 ;
        RECT 2390.985 2155.355 2391.155 2155.525 ;
        RECT 2390.985 2154.865 2391.160 2155.355 ;
        RECT 2391.570 2155.315 2391.740 2156.925 ;
        RECT 2391.940 2156.895 2392.115 2158.155 ;
        RECT 2392.370 2157.015 2392.545 2158.155 ;
        RECT 2391.940 2155.945 2392.110 2156.895 ;
        RECT 2392.370 2155.415 2392.540 2157.015 ;
        RECT 2393.730 2157.010 2393.905 2158.155 ;
        RECT 2394.715 2157.010 2394.890 2158.155 ;
        RECT 2399.575 2157.490 2399.905 2158.470 ;
        RECT 2401.385 2157.670 2401.715 2158.455 ;
        RECT 2401.035 2157.500 2401.715 2157.670 ;
        RECT 2401.905 2157.670 2402.235 2158.455 ;
        RECT 2401.905 2157.500 2402.585 2157.670 ;
        RECT 2393.360 2156.205 2393.530 2156.895 ;
        RECT 2393.730 2156.805 2393.900 2157.010 ;
        RECT 2394.345 2156.805 2394.515 2156.895 ;
        RECT 2393.730 2156.625 2394.515 2156.805 ;
        RECT 2393.730 2156.575 2393.900 2156.625 ;
        RECT 2394.345 2156.205 2394.515 2156.625 ;
        RECT 2394.715 2156.575 2394.885 2157.010 ;
        RECT 2399.575 2156.890 2399.825 2157.490 ;
        RECT 2399.995 2157.280 2400.325 2157.330 ;
        RECT 2400.515 2157.280 2400.865 2157.330 ;
        RECT 2399.995 2157.110 2400.865 2157.280 ;
        RECT 2399.995 2157.080 2400.325 2157.110 ;
        RECT 2400.515 2157.080 2400.865 2157.110 ;
        RECT 2401.035 2156.900 2401.205 2157.500 ;
        RECT 2401.375 2157.080 2401.725 2157.330 ;
        RECT 2401.895 2157.080 2402.245 2157.330 ;
        RECT 2402.415 2156.900 2402.585 2157.500 ;
        RECT 2403.275 2157.620 2403.595 2158.470 ;
        RECT 2403.775 2157.960 2404.175 2158.470 ;
        RECT 2404.685 2157.960 2405.015 2158.470 ;
        RECT 2403.775 2157.790 2405.015 2157.960 ;
        RECT 2405.595 2157.620 2405.765 2158.300 ;
        RECT 2405.945 2157.790 2406.325 2158.470 ;
        RECT 2403.275 2157.540 2403.725 2157.620 ;
        RECT 2403.275 2157.370 2403.905 2157.540 ;
        RECT 2402.755 2157.080 2403.105 2157.330 ;
        RECT 2399.575 2156.260 2399.905 2156.890 ;
        RECT 2400.965 2156.260 2401.295 2156.900 ;
        RECT 2402.325 2156.260 2402.655 2156.900 ;
        RECT 2403.735 2156.490 2403.905 2157.370 ;
        RECT 2404.680 2157.450 2405.985 2157.620 ;
        RECT 2404.075 2156.830 2404.305 2157.330 ;
        RECT 2404.680 2157.250 2404.850 2157.450 ;
        RECT 2404.475 2157.080 2404.850 2157.250 ;
        RECT 2405.020 2157.080 2405.570 2157.280 ;
        RECT 2405.740 2157.000 2405.985 2157.450 ;
        RECT 2406.155 2156.830 2406.325 2157.790 ;
        RECT 2404.075 2156.660 2406.325 2156.830 ;
        RECT 2408.205 2156.895 2408.380 2158.155 ;
        RECT 2408.730 2157.095 2408.900 2158.155 ;
        RECT 2408.730 2156.925 2408.960 2157.095 ;
        RECT 2408.205 2156.695 2408.375 2156.895 ;
        RECT 2403.735 2156.320 2404.690 2156.490 ;
        RECT 2405.605 2156.340 2405.775 2156.660 ;
        RECT 2408.205 2156.365 2408.615 2156.695 ;
        RECT 2393.360 2156.175 2393.830 2156.205 ;
        RECT 2393.315 2156.035 2393.830 2156.175 ;
        RECT 2394.345 2156.035 2394.815 2156.205 ;
        RECT 2393.315 2155.945 2393.545 2156.035 ;
        RECT 2408.205 2155.855 2408.375 2156.365 ;
        RECT 2408.205 2155.525 2408.615 2155.855 ;
        RECT 2391.510 2155.145 2391.740 2155.315 ;
        RECT 2391.510 2154.865 2391.680 2155.145 ;
        RECT 2391.940 2154.865 2392.115 2155.375 ;
        RECT 2392.370 2154.865 2392.545 2155.415 ;
        RECT 2393.735 2154.865 2393.905 2155.375 ;
        RECT 2394.720 2154.865 2394.890 2155.375 ;
        RECT 2408.205 2155.355 2408.375 2155.525 ;
        RECT 2408.205 2154.865 2408.380 2155.355 ;
        RECT 2408.790 2155.315 2408.960 2156.925 ;
        RECT 2409.160 2156.895 2409.335 2158.155 ;
        RECT 2409.590 2157.015 2409.765 2158.155 ;
        RECT 2409.160 2155.945 2409.330 2156.895 ;
        RECT 2409.590 2155.415 2409.760 2157.015 ;
        RECT 2410.950 2157.010 2411.125 2158.155 ;
        RECT 2411.935 2157.010 2412.110 2158.155 ;
        RECT 2416.795 2157.490 2417.125 2158.470 ;
        RECT 2418.605 2157.670 2418.935 2158.455 ;
        RECT 2418.255 2157.500 2418.935 2157.670 ;
        RECT 2419.125 2157.670 2419.455 2158.455 ;
        RECT 2419.125 2157.500 2419.805 2157.670 ;
        RECT 2410.580 2156.205 2410.750 2156.895 ;
        RECT 2410.950 2156.805 2411.120 2157.010 ;
        RECT 2411.565 2156.805 2411.735 2156.895 ;
        RECT 2410.950 2156.625 2411.735 2156.805 ;
        RECT 2410.950 2156.575 2411.120 2156.625 ;
        RECT 2411.565 2156.205 2411.735 2156.625 ;
        RECT 2411.935 2156.575 2412.105 2157.010 ;
        RECT 2416.795 2156.890 2417.045 2157.490 ;
        RECT 2417.215 2157.280 2417.545 2157.330 ;
        RECT 2417.735 2157.280 2418.085 2157.330 ;
        RECT 2417.215 2157.110 2418.085 2157.280 ;
        RECT 2417.215 2157.080 2417.545 2157.110 ;
        RECT 2417.735 2157.080 2418.085 2157.110 ;
        RECT 2418.255 2156.900 2418.425 2157.500 ;
        RECT 2418.595 2157.080 2418.945 2157.330 ;
        RECT 2419.115 2157.080 2419.465 2157.330 ;
        RECT 2419.635 2156.900 2419.805 2157.500 ;
        RECT 2420.495 2157.620 2420.815 2158.470 ;
        RECT 2420.995 2157.960 2421.395 2158.470 ;
        RECT 2421.905 2157.960 2422.235 2158.470 ;
        RECT 2420.995 2157.790 2422.235 2157.960 ;
        RECT 2422.815 2157.620 2422.985 2158.300 ;
        RECT 2423.165 2157.790 2423.545 2158.470 ;
        RECT 2420.495 2157.540 2420.945 2157.620 ;
        RECT 2420.495 2157.370 2421.125 2157.540 ;
        RECT 2419.975 2157.080 2420.325 2157.330 ;
        RECT 2416.795 2156.260 2417.125 2156.890 ;
        RECT 2418.185 2156.260 2418.515 2156.900 ;
        RECT 2419.545 2156.260 2419.875 2156.900 ;
        RECT 2420.955 2156.490 2421.125 2157.370 ;
        RECT 2421.900 2157.450 2423.205 2157.620 ;
        RECT 2421.295 2156.830 2421.525 2157.330 ;
        RECT 2421.900 2157.250 2422.070 2157.450 ;
        RECT 2421.695 2157.080 2422.070 2157.250 ;
        RECT 2422.240 2157.080 2422.790 2157.280 ;
        RECT 2422.960 2157.000 2423.205 2157.450 ;
        RECT 2423.375 2156.830 2423.545 2157.790 ;
        RECT 2421.295 2156.660 2423.545 2156.830 ;
        RECT 2425.425 2156.895 2425.600 2158.155 ;
        RECT 2425.950 2157.095 2426.120 2158.155 ;
        RECT 2425.950 2156.925 2426.180 2157.095 ;
        RECT 2425.425 2156.695 2425.595 2156.895 ;
        RECT 2420.955 2156.320 2421.910 2156.490 ;
        RECT 2422.825 2156.340 2422.995 2156.660 ;
        RECT 2425.425 2156.365 2425.835 2156.695 ;
        RECT 2410.580 2156.175 2411.050 2156.205 ;
        RECT 2410.535 2156.035 2411.050 2156.175 ;
        RECT 2411.565 2156.035 2412.035 2156.205 ;
        RECT 2410.535 2155.945 2410.765 2156.035 ;
        RECT 2425.425 2155.855 2425.595 2156.365 ;
        RECT 2425.425 2155.525 2425.835 2155.855 ;
        RECT 2408.730 2155.145 2408.960 2155.315 ;
        RECT 2408.730 2154.865 2408.900 2155.145 ;
        RECT 2409.160 2154.865 2409.335 2155.375 ;
        RECT 2409.590 2154.865 2409.765 2155.415 ;
        RECT 2410.955 2154.865 2411.125 2155.375 ;
        RECT 2411.940 2154.865 2412.110 2155.375 ;
        RECT 2425.425 2155.355 2425.595 2155.525 ;
        RECT 2425.425 2154.865 2425.600 2155.355 ;
        RECT 2426.010 2155.315 2426.180 2156.925 ;
        RECT 2426.380 2156.895 2426.555 2158.155 ;
        RECT 2426.810 2157.015 2426.985 2158.155 ;
        RECT 2426.380 2155.945 2426.550 2156.895 ;
        RECT 2426.810 2155.415 2426.980 2157.015 ;
        RECT 2428.170 2157.010 2428.345 2158.155 ;
        RECT 2429.155 2157.010 2429.330 2158.155 ;
        RECT 2434.015 2157.490 2434.345 2158.470 ;
        RECT 2435.825 2157.670 2436.155 2158.455 ;
        RECT 2435.475 2157.500 2436.155 2157.670 ;
        RECT 2436.345 2157.670 2436.675 2158.455 ;
        RECT 2436.345 2157.500 2437.025 2157.670 ;
        RECT 2427.800 2156.205 2427.970 2156.895 ;
        RECT 2428.170 2156.805 2428.340 2157.010 ;
        RECT 2428.785 2156.805 2428.955 2156.895 ;
        RECT 2428.170 2156.625 2428.955 2156.805 ;
        RECT 2428.170 2156.575 2428.340 2156.625 ;
        RECT 2428.785 2156.205 2428.955 2156.625 ;
        RECT 2429.155 2156.575 2429.325 2157.010 ;
        RECT 2434.015 2156.890 2434.265 2157.490 ;
        RECT 2434.435 2157.280 2434.765 2157.330 ;
        RECT 2434.955 2157.280 2435.305 2157.330 ;
        RECT 2434.435 2157.110 2435.305 2157.280 ;
        RECT 2434.435 2157.080 2434.765 2157.110 ;
        RECT 2434.955 2157.080 2435.305 2157.110 ;
        RECT 2435.475 2156.900 2435.645 2157.500 ;
        RECT 2435.815 2157.080 2436.165 2157.330 ;
        RECT 2436.335 2157.080 2436.685 2157.330 ;
        RECT 2436.855 2156.900 2437.025 2157.500 ;
        RECT 2437.715 2157.620 2438.035 2158.470 ;
        RECT 2438.215 2157.960 2438.615 2158.470 ;
        RECT 2439.125 2157.960 2439.455 2158.470 ;
        RECT 2438.215 2157.790 2439.455 2157.960 ;
        RECT 2440.035 2157.620 2440.205 2158.300 ;
        RECT 2440.385 2157.790 2440.765 2158.470 ;
        RECT 2696.985 2158.155 2697.325 2159.035 ;
        RECT 2697.495 2158.325 2697.665 2159.545 ;
        RECT 2698.690 2159.205 2699.165 2159.545 ;
        RECT 2697.905 2158.675 2698.155 2159.040 ;
        RECT 2698.875 2158.675 2699.590 2158.970 ;
        RECT 2699.760 2158.845 2700.035 2159.545 ;
        RECT 2697.905 2158.505 2699.695 2158.675 ;
        RECT 2437.715 2157.540 2438.165 2157.620 ;
        RECT 2437.715 2157.370 2438.345 2157.540 ;
        RECT 2437.195 2157.080 2437.545 2157.330 ;
        RECT 2434.015 2156.260 2434.345 2156.890 ;
        RECT 2435.405 2156.260 2435.735 2156.900 ;
        RECT 2436.765 2156.260 2437.095 2156.900 ;
        RECT 2438.175 2156.490 2438.345 2157.370 ;
        RECT 2439.120 2157.450 2440.425 2157.620 ;
        RECT 2438.515 2156.830 2438.745 2157.330 ;
        RECT 2439.120 2157.250 2439.290 2157.450 ;
        RECT 2438.915 2157.080 2439.290 2157.250 ;
        RECT 2439.460 2157.080 2440.010 2157.280 ;
        RECT 2440.180 2157.000 2440.425 2157.450 ;
        RECT 2440.595 2156.830 2440.765 2157.790 ;
        RECT 2438.515 2156.660 2440.765 2156.830 ;
        RECT 2442.645 2156.895 2442.820 2158.155 ;
        RECT 2443.170 2157.095 2443.340 2158.155 ;
        RECT 2443.170 2156.925 2443.400 2157.095 ;
        RECT 2442.645 2156.695 2442.815 2156.895 ;
        RECT 2438.175 2156.320 2439.130 2156.490 ;
        RECT 2440.045 2156.340 2440.215 2156.660 ;
        RECT 2442.645 2156.365 2443.055 2156.695 ;
        RECT 2427.800 2156.175 2428.270 2156.205 ;
        RECT 2427.755 2156.035 2428.270 2156.175 ;
        RECT 2428.785 2156.035 2429.255 2156.205 ;
        RECT 2427.755 2155.945 2427.985 2156.035 ;
        RECT 2442.645 2155.855 2442.815 2156.365 ;
        RECT 2442.645 2155.525 2443.055 2155.855 ;
        RECT 2425.950 2155.145 2426.180 2155.315 ;
        RECT 2425.950 2154.865 2426.120 2155.145 ;
        RECT 2426.380 2154.865 2426.555 2155.375 ;
        RECT 2426.810 2154.865 2426.985 2155.415 ;
        RECT 2428.175 2154.865 2428.345 2155.375 ;
        RECT 2429.160 2154.865 2429.330 2155.375 ;
        RECT 2442.645 2155.355 2442.815 2155.525 ;
        RECT 2442.645 2154.865 2442.820 2155.355 ;
        RECT 2443.230 2155.315 2443.400 2156.925 ;
        RECT 2443.600 2156.895 2443.775 2158.155 ;
        RECT 2444.030 2157.015 2444.205 2158.155 ;
        RECT 2443.600 2155.945 2443.770 2156.895 ;
        RECT 2444.030 2155.415 2444.200 2157.015 ;
        RECT 2445.390 2157.010 2445.565 2158.155 ;
        RECT 2446.375 2157.010 2446.550 2158.155 ;
        RECT 2697.495 2158.075 2698.290 2158.325 ;
        RECT 2697.495 2157.985 2697.745 2158.075 ;
        RECT 2697.415 2157.565 2697.745 2157.985 ;
        RECT 2698.460 2157.650 2698.715 2158.505 ;
        RECT 2697.925 2157.385 2698.715 2157.650 ;
        RECT 2698.885 2157.805 2699.295 2158.325 ;
        RECT 2699.465 2158.075 2699.695 2158.505 ;
        RECT 2699.865 2157.815 2700.035 2158.845 ;
        RECT 2882.085 2158.380 2882.605 2159.930 ;
        RECT 2698.885 2157.385 2699.085 2157.805 ;
        RECT 2699.775 2157.335 2700.035 2157.815 ;
        RECT 2445.020 2156.205 2445.190 2156.895 ;
        RECT 2445.390 2156.805 2445.560 2157.010 ;
        RECT 2446.005 2156.805 2446.175 2156.895 ;
        RECT 2445.390 2156.625 2446.175 2156.805 ;
        RECT 2445.390 2156.575 2445.560 2156.625 ;
        RECT 2446.005 2156.205 2446.175 2156.625 ;
        RECT 2446.375 2156.575 2446.545 2157.010 ;
        RECT 2697.075 2156.445 2697.245 2156.825 ;
        RECT 2697.075 2156.275 2697.740 2156.445 ;
        RECT 2697.935 2156.320 2698.195 2156.825 ;
        RECT 2445.020 2156.175 2445.490 2156.205 ;
        RECT 2444.975 2156.035 2445.490 2156.175 ;
        RECT 2446.005 2156.035 2446.475 2156.205 ;
        RECT 2444.975 2155.945 2445.205 2156.035 ;
        RECT 2697.005 2155.725 2697.335 2156.095 ;
        RECT 2697.570 2156.020 2697.740 2156.275 ;
        RECT 2697.570 2155.690 2697.855 2156.020 ;
        RECT 2697.570 2155.545 2697.740 2155.690 ;
        RECT 2443.170 2155.145 2443.400 2155.315 ;
        RECT 2443.170 2154.865 2443.340 2155.145 ;
        RECT 2443.600 2154.865 2443.775 2155.375 ;
        RECT 2444.030 2154.865 2444.205 2155.415 ;
        RECT 2697.075 2155.375 2697.740 2155.545 ;
        RECT 2698.025 2155.520 2698.195 2156.320 ;
        RECT 2445.395 2154.865 2445.565 2155.375 ;
        RECT 2446.380 2154.865 2446.550 2155.375 ;
        RECT 2697.075 2154.615 2697.245 2155.375 ;
        RECT 2697.925 2154.615 2698.195 2155.520 ;
        RECT 2698.455 2153.605 2698.625 2154.105 ;
        RECT 2699.415 2153.605 2699.585 2154.105 ;
        RECT 2700.255 2153.605 2700.425 2154.105 ;
        RECT 2698.455 2153.435 2700.425 2153.605 ;
        RECT 2700.595 2153.635 2700.925 2154.065 ;
        RECT 2701.535 2153.805 2701.875 2154.065 ;
        RECT 2700.595 2153.465 2701.445 2153.635 ;
        RECT 2698.390 2152.635 2698.645 2153.265 ;
        RECT 2698.875 2152.635 2699.255 2153.265 ;
        RECT 2700.125 2153.255 2700.425 2153.260 ;
        RECT 2700.125 2153.085 2700.435 2153.255 ;
        RECT 2700.125 2152.965 2700.425 2153.085 ;
        RECT 2698.875 2152.035 2699.080 2152.635 ;
        RECT 2699.515 2152.240 2699.735 2152.965 ;
        RECT 2700.045 2152.635 2700.425 2152.965 ;
        RECT 2700.625 2152.715 2700.955 2153.275 ;
        RECT 2701.275 2152.545 2701.445 2153.465 ;
        RECT 2700.625 2152.450 2701.445 2152.545 ;
        RECT 2700.430 2152.375 2701.445 2152.450 ;
        RECT 2699.310 2152.055 2700.260 2152.240 ;
        RECT 2700.430 2151.940 2700.845 2152.375 ;
        RECT 2701.615 2152.200 2701.875 2153.805 ;
        RECT 2701.535 2151.940 2701.875 2152.200 ;
        RECT 2698.335 2150.735 2698.665 2151.155 ;
        RECT 2698.845 2150.985 2699.105 2151.385 ;
        RECT 2699.775 2150.985 2699.945 2151.335 ;
        RECT 2698.845 2150.815 2700.510 2150.985 ;
        RECT 2700.680 2150.880 2700.955 2151.225 ;
        RECT 2698.415 2150.645 2698.665 2150.735 ;
        RECT 2700.340 2150.645 2700.510 2150.815 ;
        RECT 2697.910 2150.315 2698.245 2150.565 ;
        RECT 2698.415 2150.315 2699.130 2150.645 ;
        RECT 2699.345 2150.315 2700.170 2150.645 ;
        RECT 2700.340 2150.315 2700.615 2150.645 ;
        RECT 2698.415 2149.755 2698.585 2150.315 ;
        RECT 2698.845 2149.855 2699.175 2150.145 ;
        RECT 2699.345 2150.025 2699.590 2150.315 ;
        RECT 2700.340 2150.145 2700.510 2150.315 ;
        RECT 2700.785 2150.145 2700.955 2150.880 ;
        RECT 2699.850 2149.975 2700.510 2150.145 ;
        RECT 2699.850 2149.855 2700.020 2149.975 ;
        RECT 2698.845 2149.685 2700.020 2149.855 ;
        RECT 2698.405 2149.185 2700.020 2149.515 ;
        RECT 2700.680 2149.175 2700.955 2150.145 ;
        RECT 2701.125 2151.155 2701.715 2151.385 ;
        RECT 2701.125 2150.145 2701.415 2151.155 ;
        RECT 2703.290 2150.985 2703.715 2151.195 ;
        RECT 2701.585 2150.815 2703.715 2150.985 ;
        RECT 2701.585 2150.315 2701.755 2150.815 ;
        RECT 2702.045 2150.315 2702.375 2150.645 ;
        RECT 2702.565 2150.315 2702.835 2150.645 ;
        RECT 2703.025 2150.315 2703.375 2150.645 ;
        RECT 2701.125 2149.975 2702.670 2150.145 ;
        RECT 2703.545 2150.045 2703.715 2150.815 ;
        RECT 2701.125 2149.175 2701.715 2149.975 ;
        RECT 2702.340 2149.175 2702.670 2149.975 ;
        RECT 2703.290 2149.715 2703.715 2150.045 ;
        RECT 2697.075 2147.905 2697.245 2148.665 ;
        RECT 2697.075 2147.735 2697.740 2147.905 ;
        RECT 2697.925 2147.760 2698.195 2148.665 ;
        RECT 2697.570 2147.590 2697.740 2147.735 ;
        RECT 2697.005 2147.185 2697.335 2147.555 ;
        RECT 2697.570 2147.260 2697.855 2147.590 ;
        RECT 2697.570 2147.005 2697.740 2147.260 ;
        RECT 2697.075 2146.835 2697.740 2147.005 ;
        RECT 2698.025 2146.960 2698.195 2147.760 ;
        RECT 2699.255 2147.685 2699.585 2148.665 ;
        RECT 2698.845 2147.275 2699.180 2147.525 ;
        RECT 2699.350 2147.085 2699.520 2147.685 ;
        RECT 2699.690 2147.255 2700.025 2147.525 ;
        RECT 2697.075 2146.455 2697.245 2146.835 ;
        RECT 2697.935 2146.455 2698.195 2146.960 ;
        RECT 2698.825 2146.455 2699.520 2147.085 ;
        RECT 2697.260 2145.305 2697.505 2145.910 ;
        RECT 2696.985 2145.135 2698.215 2145.305 ;
        RECT 2696.985 2144.325 2697.325 2145.135 ;
        RECT 2697.495 2144.570 2698.245 2144.760 ;
        RECT 2696.985 2143.915 2697.500 2144.325 ;
        RECT 2698.075 2143.905 2698.245 2144.570 ;
        RECT 2698.415 2144.585 2698.605 2145.945 ;
        RECT 2698.775 2145.095 2699.050 2145.945 ;
        RECT 2699.240 2145.580 2699.770 2145.945 ;
        RECT 2699.595 2145.545 2699.770 2145.580 ;
        RECT 2698.775 2144.925 2699.055 2145.095 ;
        RECT 2698.775 2144.785 2699.050 2144.925 ;
        RECT 2699.255 2144.585 2699.425 2145.385 ;
        RECT 2698.415 2144.415 2699.425 2144.585 ;
        RECT 2699.595 2145.375 2700.525 2145.545 ;
        RECT 2700.695 2145.375 2700.950 2145.945 ;
        RECT 2699.595 2144.245 2699.765 2145.375 ;
        RECT 2700.355 2145.205 2700.525 2145.375 ;
        RECT 2698.640 2144.075 2699.765 2144.245 ;
        RECT 2699.935 2144.875 2700.130 2145.205 ;
        RECT 2700.355 2144.875 2700.610 2145.205 ;
        RECT 2699.935 2143.905 2700.105 2144.875 ;
        RECT 2700.780 2144.705 2700.950 2145.375 ;
        RECT 2698.075 2143.735 2700.105 2143.905 ;
        RECT 2700.615 2143.735 2700.950 2144.705 ;
        RECT 2697.075 2142.465 2697.245 2143.225 ;
        RECT 2697.075 2142.295 2697.740 2142.465 ;
        RECT 2697.925 2142.320 2698.195 2143.225 ;
        RECT 2697.570 2142.150 2697.740 2142.295 ;
        RECT 2697.005 2141.745 2697.335 2142.115 ;
        RECT 2697.570 2141.820 2697.855 2142.150 ;
        RECT 2697.570 2141.565 2697.740 2141.820 ;
        RECT 2697.075 2141.395 2697.740 2141.565 ;
        RECT 2698.025 2141.520 2698.195 2142.320 ;
        RECT 2697.075 2141.015 2697.245 2141.395 ;
        RECT 2697.935 2141.015 2698.195 2141.520 ;
        RECT 2697.075 2137.025 2697.245 2137.785 ;
        RECT 2697.075 2136.855 2697.740 2137.025 ;
        RECT 2697.925 2136.880 2698.195 2137.785 ;
        RECT 2697.570 2136.710 2697.740 2136.855 ;
        RECT 2522.640 2134.210 2523.160 2135.695 ;
        RECT 2523.330 2134.870 2523.850 2136.420 ;
        RECT 2697.005 2136.305 2697.335 2136.675 ;
        RECT 2697.570 2136.380 2697.855 2136.710 ;
        RECT 2697.570 2136.125 2697.740 2136.380 ;
        RECT 2697.075 2135.955 2697.740 2136.125 ;
        RECT 2698.025 2136.080 2698.195 2136.880 ;
        RECT 2697.075 2135.575 2697.245 2135.955 ;
        RECT 2697.935 2135.575 2698.195 2136.080 ;
        RECT 2697.075 2131.585 2697.245 2132.345 ;
        RECT 2697.075 2131.415 2697.740 2131.585 ;
        RECT 2697.925 2131.440 2698.195 2132.345 ;
        RECT 2697.570 2131.270 2697.740 2131.415 ;
        RECT 2697.005 2130.865 2697.335 2131.235 ;
        RECT 2697.570 2130.940 2697.855 2131.270 ;
        RECT 2697.570 2130.685 2697.740 2130.940 ;
        RECT 2697.075 2130.515 2697.740 2130.685 ;
        RECT 2698.025 2130.640 2698.195 2131.440 ;
        RECT 2698.455 2131.585 2698.625 2132.345 ;
        RECT 2698.455 2131.415 2699.120 2131.585 ;
        RECT 2699.305 2131.440 2699.575 2132.345 ;
        RECT 2698.950 2131.270 2699.120 2131.415 ;
        RECT 2698.385 2130.865 2698.715 2131.235 ;
        RECT 2698.950 2130.940 2699.235 2131.270 ;
        RECT 2698.950 2130.685 2699.120 2130.940 ;
        RECT 2697.075 2130.135 2697.245 2130.515 ;
        RECT 2697.935 2130.135 2698.195 2130.640 ;
        RECT 2698.455 2130.515 2699.120 2130.685 ;
        RECT 2699.405 2130.640 2699.575 2131.440 ;
        RECT 2698.455 2130.135 2698.625 2130.515 ;
        RECT 2699.315 2130.135 2699.575 2130.640 ;
        RECT 2522.640 2126.680 2523.160 2128.165 ;
        RECT 2523.330 2127.340 2523.850 2128.890 ;
        RECT 2522.640 2120.700 2523.160 2122.185 ;
        RECT 2523.330 2121.360 2523.850 2122.910 ;
        RECT 2522.640 2114.755 2523.160 2116.240 ;
        RECT 2523.330 2115.415 2523.850 2116.965 ;
        RECT 2522.640 2109.110 2523.160 2110.595 ;
        RECT 2523.330 2109.770 2523.850 2111.320 ;
        RECT 2522.640 2103.105 2523.160 2104.590 ;
        RECT 2523.330 2103.765 2523.850 2105.315 ;
        RECT 2358.650 2058.105 2358.825 2058.595 ;
        RECT 2359.175 2058.315 2359.345 2058.595 ;
        RECT 2359.175 2058.145 2359.405 2058.315 ;
        RECT 2358.650 2057.935 2358.820 2058.105 ;
        RECT 2358.650 2057.605 2359.060 2057.935 ;
        RECT 2358.650 2057.095 2358.820 2057.605 ;
        RECT 2358.650 2056.765 2359.060 2057.095 ;
        RECT 2358.650 2056.565 2358.820 2056.765 ;
        RECT 2358.650 2055.305 2358.825 2056.565 ;
        RECT 2359.235 2056.535 2359.405 2058.145 ;
        RECT 2359.605 2058.085 2359.780 2058.595 ;
        RECT 2367.230 2058.105 2367.405 2058.595 ;
        RECT 2367.230 2057.935 2367.400 2058.105 ;
        RECT 2368.185 2058.085 2368.360 2058.595 ;
        RECT 2368.615 2058.045 2368.790 2058.595 ;
        RECT 2372.845 2058.105 2373.020 2058.595 ;
        RECT 2373.370 2058.315 2373.540 2058.595 ;
        RECT 2373.370 2058.145 2373.600 2058.315 ;
        RECT 2367.230 2057.605 2367.640 2057.935 ;
        RECT 2359.175 2056.365 2359.405 2056.535 ;
        RECT 2359.605 2056.565 2359.775 2057.515 ;
        RECT 2367.230 2057.095 2367.400 2057.605 ;
        RECT 2367.230 2056.765 2367.640 2057.095 ;
        RECT 2367.230 2056.565 2367.400 2056.765 ;
        RECT 2368.185 2056.565 2368.355 2057.515 ;
        RECT 2359.175 2055.305 2359.345 2056.365 ;
        RECT 2359.605 2055.305 2359.780 2056.565 ;
        RECT 2367.230 2055.305 2367.405 2056.565 ;
        RECT 2368.185 2055.305 2368.360 2056.565 ;
        RECT 2368.615 2056.445 2368.785 2058.045 ;
        RECT 2372.845 2057.935 2373.015 2058.105 ;
        RECT 2372.845 2057.605 2373.255 2057.935 ;
        RECT 2372.845 2057.095 2373.015 2057.605 ;
        RECT 2372.845 2056.765 2373.255 2057.095 ;
        RECT 2372.845 2056.565 2373.015 2056.765 ;
        RECT 2368.615 2055.305 2368.790 2056.445 ;
        RECT 2372.845 2055.305 2373.020 2056.565 ;
        RECT 2373.430 2056.535 2373.600 2058.145 ;
        RECT 2373.800 2058.085 2373.975 2058.595 ;
        RECT 2374.230 2058.045 2374.405 2058.595 ;
        RECT 2375.595 2058.085 2375.765 2058.595 ;
        RECT 2376.590 2058.080 2376.760 2058.590 ;
        RECT 2383.555 2058.105 2383.730 2058.595 ;
        RECT 2373.370 2056.365 2373.600 2056.535 ;
        RECT 2373.800 2056.565 2373.970 2057.515 ;
        RECT 2373.370 2055.305 2373.540 2056.365 ;
        RECT 2373.800 2055.305 2373.975 2056.565 ;
        RECT 2374.230 2056.445 2374.400 2058.045 ;
        RECT 2383.555 2057.935 2383.725 2058.105 ;
        RECT 2384.510 2058.085 2384.685 2058.595 ;
        RECT 2384.940 2058.045 2385.115 2058.595 ;
        RECT 2389.170 2058.105 2389.345 2058.595 ;
        RECT 2389.695 2058.315 2389.865 2058.595 ;
        RECT 2389.695 2058.145 2389.925 2058.315 ;
        RECT 2383.555 2057.605 2383.965 2057.935 ;
        RECT 2374.770 2057.425 2375.000 2057.575 ;
        RECT 2374.770 2057.255 2375.690 2057.425 ;
        RECT 2375.220 2056.565 2375.390 2057.255 ;
        RECT 2376.215 2057.250 2376.685 2057.420 ;
        RECT 2375.590 2056.775 2375.760 2056.885 ;
        RECT 2376.215 2056.775 2376.385 2057.250 ;
        RECT 2383.555 2057.095 2383.725 2057.605 ;
        RECT 2375.590 2056.605 2376.385 2056.775 ;
        RECT 2374.230 2055.305 2374.405 2056.445 ;
        RECT 2375.590 2055.305 2375.765 2056.605 ;
        RECT 2376.215 2056.560 2376.385 2056.605 ;
        RECT 2376.585 2056.445 2376.755 2056.880 ;
        RECT 2383.555 2056.765 2383.965 2057.095 ;
        RECT 2383.555 2056.565 2383.725 2056.765 ;
        RECT 2384.510 2056.565 2384.680 2057.515 ;
        RECT 2376.585 2055.300 2376.760 2056.445 ;
        RECT 2383.555 2055.305 2383.730 2056.565 ;
        RECT 2384.510 2055.305 2384.685 2056.565 ;
        RECT 2384.940 2056.445 2385.110 2058.045 ;
        RECT 2389.170 2057.935 2389.340 2058.105 ;
        RECT 2389.170 2057.605 2389.580 2057.935 ;
        RECT 2389.170 2057.095 2389.340 2057.605 ;
        RECT 2389.170 2056.765 2389.580 2057.095 ;
        RECT 2389.170 2056.565 2389.340 2056.765 ;
        RECT 2384.940 2055.305 2385.115 2056.445 ;
        RECT 2389.170 2055.305 2389.345 2056.565 ;
        RECT 2389.755 2056.535 2389.925 2058.145 ;
        RECT 2390.125 2058.085 2390.300 2058.595 ;
        RECT 2390.555 2058.045 2390.730 2058.595 ;
        RECT 2391.920 2058.085 2392.090 2058.595 ;
        RECT 2392.915 2058.080 2393.085 2058.590 ;
        RECT 2399.880 2058.105 2400.055 2058.595 ;
        RECT 2389.695 2056.365 2389.925 2056.535 ;
        RECT 2390.125 2056.565 2390.295 2057.515 ;
        RECT 2389.695 2055.305 2389.865 2056.365 ;
        RECT 2390.125 2055.305 2390.300 2056.565 ;
        RECT 2390.555 2056.445 2390.725 2058.045 ;
        RECT 2399.880 2057.935 2400.050 2058.105 ;
        RECT 2400.835 2058.085 2401.010 2058.595 ;
        RECT 2401.265 2058.045 2401.440 2058.595 ;
        RECT 2405.495 2058.105 2405.670 2058.595 ;
        RECT 2406.020 2058.315 2406.190 2058.595 ;
        RECT 2406.020 2058.145 2406.250 2058.315 ;
        RECT 2399.880 2057.605 2400.290 2057.935 ;
        RECT 2391.095 2057.425 2391.325 2057.575 ;
        RECT 2391.095 2057.255 2392.015 2057.425 ;
        RECT 2391.545 2056.565 2391.715 2057.255 ;
        RECT 2392.540 2057.250 2393.010 2057.420 ;
        RECT 2391.915 2056.775 2392.085 2056.885 ;
        RECT 2392.540 2056.775 2392.710 2057.250 ;
        RECT 2399.880 2057.095 2400.050 2057.605 ;
        RECT 2391.915 2056.605 2392.710 2056.775 ;
        RECT 2390.555 2055.305 2390.730 2056.445 ;
        RECT 2391.915 2055.305 2392.090 2056.605 ;
        RECT 2392.540 2056.560 2392.710 2056.605 ;
        RECT 2392.910 2056.445 2393.080 2056.880 ;
        RECT 2399.880 2056.765 2400.290 2057.095 ;
        RECT 2399.880 2056.565 2400.050 2056.765 ;
        RECT 2400.835 2056.565 2401.005 2057.515 ;
        RECT 2392.910 2055.300 2393.085 2056.445 ;
        RECT 2399.880 2055.305 2400.055 2056.565 ;
        RECT 2400.835 2055.305 2401.010 2056.565 ;
        RECT 2401.265 2056.445 2401.435 2058.045 ;
        RECT 2405.495 2057.935 2405.665 2058.105 ;
        RECT 2405.495 2057.605 2405.905 2057.935 ;
        RECT 2405.495 2057.095 2405.665 2057.605 ;
        RECT 2405.495 2056.765 2405.905 2057.095 ;
        RECT 2405.495 2056.565 2405.665 2056.765 ;
        RECT 2401.265 2055.305 2401.440 2056.445 ;
        RECT 2405.495 2055.305 2405.670 2056.565 ;
        RECT 2406.080 2056.535 2406.250 2058.145 ;
        RECT 2406.450 2058.085 2406.625 2058.595 ;
        RECT 2406.880 2058.045 2407.055 2058.595 ;
        RECT 2408.245 2058.085 2408.415 2058.595 ;
        RECT 2409.240 2058.080 2409.410 2058.590 ;
        RECT 2416.205 2058.105 2416.380 2058.595 ;
        RECT 2406.020 2056.365 2406.250 2056.535 ;
        RECT 2406.450 2056.565 2406.620 2057.515 ;
        RECT 2406.020 2055.305 2406.190 2056.365 ;
        RECT 2406.450 2055.305 2406.625 2056.565 ;
        RECT 2406.880 2056.445 2407.050 2058.045 ;
        RECT 2416.205 2057.935 2416.375 2058.105 ;
        RECT 2417.160 2058.085 2417.335 2058.595 ;
        RECT 2417.590 2058.045 2417.765 2058.595 ;
        RECT 2421.820 2058.105 2421.995 2058.595 ;
        RECT 2422.345 2058.315 2422.515 2058.595 ;
        RECT 2422.345 2058.145 2422.575 2058.315 ;
        RECT 2416.205 2057.605 2416.615 2057.935 ;
        RECT 2407.420 2057.425 2407.650 2057.575 ;
        RECT 2407.420 2057.255 2408.340 2057.425 ;
        RECT 2407.870 2056.565 2408.040 2057.255 ;
        RECT 2408.865 2057.250 2409.335 2057.420 ;
        RECT 2408.240 2056.775 2408.410 2056.885 ;
        RECT 2408.865 2056.775 2409.035 2057.250 ;
        RECT 2416.205 2057.095 2416.375 2057.605 ;
        RECT 2408.240 2056.605 2409.035 2056.775 ;
        RECT 2406.880 2055.305 2407.055 2056.445 ;
        RECT 2408.240 2055.305 2408.415 2056.605 ;
        RECT 2408.865 2056.560 2409.035 2056.605 ;
        RECT 2409.235 2056.445 2409.405 2056.880 ;
        RECT 2416.205 2056.765 2416.615 2057.095 ;
        RECT 2416.205 2056.565 2416.375 2056.765 ;
        RECT 2417.160 2056.565 2417.330 2057.515 ;
        RECT 2409.235 2055.300 2409.410 2056.445 ;
        RECT 2416.205 2055.305 2416.380 2056.565 ;
        RECT 2417.160 2055.305 2417.335 2056.565 ;
        RECT 2417.590 2056.445 2417.760 2058.045 ;
        RECT 2421.820 2057.935 2421.990 2058.105 ;
        RECT 2421.820 2057.605 2422.230 2057.935 ;
        RECT 2421.820 2057.095 2421.990 2057.605 ;
        RECT 2421.820 2056.765 2422.230 2057.095 ;
        RECT 2421.820 2056.565 2421.990 2056.765 ;
        RECT 2417.590 2055.305 2417.765 2056.445 ;
        RECT 2421.820 2055.305 2421.995 2056.565 ;
        RECT 2422.405 2056.535 2422.575 2058.145 ;
        RECT 2422.775 2058.085 2422.950 2058.595 ;
        RECT 2423.205 2058.045 2423.380 2058.595 ;
        RECT 2424.570 2058.085 2424.740 2058.595 ;
        RECT 2425.565 2058.080 2425.735 2058.590 ;
        RECT 2432.530 2058.105 2432.705 2058.595 ;
        RECT 2422.345 2056.365 2422.575 2056.535 ;
        RECT 2422.775 2056.565 2422.945 2057.515 ;
        RECT 2422.345 2055.305 2422.515 2056.365 ;
        RECT 2422.775 2055.305 2422.950 2056.565 ;
        RECT 2423.205 2056.445 2423.375 2058.045 ;
        RECT 2432.530 2057.935 2432.700 2058.105 ;
        RECT 2433.485 2058.085 2433.660 2058.595 ;
        RECT 2433.915 2058.045 2434.090 2058.595 ;
        RECT 2438.145 2058.105 2438.320 2058.595 ;
        RECT 2438.670 2058.315 2438.840 2058.595 ;
        RECT 2438.670 2058.145 2438.900 2058.315 ;
        RECT 2432.530 2057.605 2432.940 2057.935 ;
        RECT 2423.745 2057.425 2423.975 2057.575 ;
        RECT 2423.745 2057.255 2424.665 2057.425 ;
        RECT 2424.195 2056.565 2424.365 2057.255 ;
        RECT 2425.190 2057.250 2425.660 2057.420 ;
        RECT 2424.565 2056.775 2424.735 2056.885 ;
        RECT 2425.190 2056.775 2425.360 2057.250 ;
        RECT 2432.530 2057.095 2432.700 2057.605 ;
        RECT 2424.565 2056.605 2425.360 2056.775 ;
        RECT 2423.205 2055.305 2423.380 2056.445 ;
        RECT 2424.565 2055.305 2424.740 2056.605 ;
        RECT 2425.190 2056.560 2425.360 2056.605 ;
        RECT 2425.560 2056.445 2425.730 2056.880 ;
        RECT 2432.530 2056.765 2432.940 2057.095 ;
        RECT 2432.530 2056.565 2432.700 2056.765 ;
        RECT 2433.485 2056.565 2433.655 2057.515 ;
        RECT 2425.560 2055.300 2425.735 2056.445 ;
        RECT 2432.530 2055.305 2432.705 2056.565 ;
        RECT 2433.485 2055.305 2433.660 2056.565 ;
        RECT 2433.915 2056.445 2434.085 2058.045 ;
        RECT 2438.145 2057.935 2438.315 2058.105 ;
        RECT 2438.145 2057.605 2438.555 2057.935 ;
        RECT 2438.145 2057.095 2438.315 2057.605 ;
        RECT 2438.145 2056.765 2438.555 2057.095 ;
        RECT 2438.145 2056.565 2438.315 2056.765 ;
        RECT 2433.915 2055.305 2434.090 2056.445 ;
        RECT 2438.145 2055.305 2438.320 2056.565 ;
        RECT 2438.730 2056.535 2438.900 2058.145 ;
        RECT 2439.100 2058.085 2439.275 2058.595 ;
        RECT 2439.530 2058.045 2439.705 2058.595 ;
        RECT 2440.895 2058.085 2441.065 2058.595 ;
        RECT 2441.890 2058.080 2442.060 2058.590 ;
        RECT 2438.670 2056.365 2438.900 2056.535 ;
        RECT 2439.100 2056.565 2439.270 2057.515 ;
        RECT 2438.670 2055.305 2438.840 2056.365 ;
        RECT 2439.100 2055.305 2439.275 2056.565 ;
        RECT 2439.530 2056.445 2439.700 2058.045 ;
        RECT 2440.070 2057.425 2440.300 2057.575 ;
        RECT 2440.070 2057.255 2440.990 2057.425 ;
        RECT 2440.520 2056.565 2440.690 2057.255 ;
        RECT 2441.515 2057.250 2441.985 2057.420 ;
        RECT 2440.890 2056.775 2441.060 2056.885 ;
        RECT 2441.515 2056.775 2441.685 2057.250 ;
        RECT 2440.890 2056.605 2441.685 2056.775 ;
        RECT 2439.530 2055.305 2439.705 2056.445 ;
        RECT 2440.890 2055.305 2441.065 2056.605 ;
        RECT 2441.515 2056.560 2441.685 2056.605 ;
        RECT 2441.885 2056.445 2442.055 2056.880 ;
        RECT 2441.885 2055.300 2442.060 2056.445 ;
        RECT 2362.230 2052.905 2362.520 2053.075 ;
        RECT 2361.870 2052.345 2362.040 2052.765 ;
        RECT 2362.230 2052.035 2362.400 2052.905 ;
        RECT 2363.550 2052.625 2363.960 2052.795 ;
        RECT 2362.030 2051.865 2362.400 2052.035 ;
        RECT 2362.590 2052.345 2363.240 2052.515 ;
        RECT 2363.790 2052.435 2363.960 2052.625 ;
        RECT 2364.310 2052.345 2364.480 2052.765 ;
        RECT 2364.670 2052.625 2364.960 2052.795 ;
        RECT 2362.590 2051.785 2362.760 2052.345 ;
        RECT 2363.070 2051.785 2363.240 2052.115 ;
        RECT 2364.670 2052.035 2364.840 2052.625 ;
        RECT 2365.750 2052.435 2365.920 2052.795 ;
        RECT 2368.190 2052.775 2368.360 2053.105 ;
        RECT 2369.190 2052.775 2369.360 2053.105 ;
        RECT 2366.670 2052.605 2367.960 2052.685 ;
        RECT 2368.590 2052.605 2368.920 2052.685 ;
        RECT 2366.670 2052.515 2368.920 2052.605 ;
        RECT 2370.070 2052.515 2370.400 2052.685 ;
        RECT 2367.710 2052.435 2368.840 2052.515 ;
        RECT 2369.310 2052.345 2370.320 2052.515 ;
        RECT 2363.470 2051.865 2363.960 2052.035 ;
        RECT 2364.470 2051.865 2364.840 2052.035 ;
        RECT 2363.790 2051.785 2363.960 2051.865 ;
        RECT 2365.030 2051.785 2365.200 2052.115 ;
        RECT 2365.510 2051.785 2365.680 2052.235 ;
        RECT 2365.910 2051.865 2367.240 2052.035 ;
        RECT 2366.990 2051.785 2367.160 2051.865 ;
        RECT 2367.470 2051.785 2367.640 2052.115 ;
        RECT 2367.950 2051.785 2368.120 2052.235 ;
        RECT 2369.310 2052.115 2369.480 2052.345 ;
        RECT 2369.310 2051.865 2369.600 2052.115 ;
        RECT 2369.430 2051.785 2369.600 2051.865 ;
        RECT 2369.910 2051.785 2370.080 2052.115 ;
        RECT 2372.845 2051.895 2373.020 2053.155 ;
        RECT 2373.370 2052.095 2373.540 2053.155 ;
        RECT 2373.370 2051.925 2373.600 2052.095 ;
        RECT 2372.845 2051.695 2373.015 2051.895 ;
        RECT 2365.990 2051.635 2366.160 2051.675 ;
        RECT 2365.990 2051.465 2366.480 2051.635 ;
        RECT 2368.430 2051.505 2368.840 2051.675 ;
        RECT 2362.350 2051.045 2362.520 2051.395 ;
        RECT 2363.310 2051.045 2363.480 2051.395 ;
        RECT 2364.790 2051.045 2364.960 2051.395 ;
        RECT 2366.750 2051.045 2366.920 2051.395 ;
        RECT 2368.670 2051.045 2368.840 2051.505 ;
        RECT 2369.190 2051.045 2369.360 2051.395 ;
        RECT 2370.150 2051.295 2370.320 2051.395 ;
        RECT 2372.845 2051.365 2373.255 2051.695 ;
        RECT 2370.150 2051.125 2370.880 2051.295 ;
        RECT 2372.845 2050.855 2373.015 2051.365 ;
        RECT 2372.845 2050.525 2373.255 2050.855 ;
        RECT 2372.845 2050.355 2373.015 2050.525 ;
        RECT 2372.845 2049.865 2373.020 2050.355 ;
        RECT 2373.430 2050.315 2373.600 2051.925 ;
        RECT 2373.800 2051.895 2373.975 2053.155 ;
        RECT 2374.230 2052.015 2374.405 2053.155 ;
        RECT 2373.800 2050.945 2373.970 2051.895 ;
        RECT 2374.230 2050.415 2374.400 2052.015 ;
        RECT 2375.590 2052.010 2375.765 2053.155 ;
        RECT 2376.580 2052.015 2376.755 2053.160 ;
        RECT 2378.555 2052.905 2378.845 2053.075 ;
        RECT 2378.195 2052.345 2378.365 2052.765 ;
        RECT 2378.555 2052.035 2378.725 2052.905 ;
        RECT 2379.875 2052.625 2380.285 2052.795 ;
        RECT 2375.220 2051.205 2375.390 2051.895 ;
        RECT 2375.590 2051.795 2375.760 2052.010 ;
        RECT 2376.210 2051.795 2376.380 2051.900 ;
        RECT 2375.590 2051.625 2376.380 2051.795 ;
        RECT 2375.590 2051.575 2375.760 2051.625 ;
        RECT 2376.210 2051.210 2376.380 2051.625 ;
        RECT 2376.580 2051.580 2376.750 2052.015 ;
        RECT 2378.355 2051.865 2378.725 2052.035 ;
        RECT 2378.915 2052.345 2379.565 2052.515 ;
        RECT 2380.115 2052.435 2380.285 2052.625 ;
        RECT 2380.635 2052.345 2380.805 2052.765 ;
        RECT 2380.995 2052.625 2381.285 2052.795 ;
        RECT 2378.915 2051.785 2379.085 2052.345 ;
        RECT 2379.395 2051.785 2379.565 2052.115 ;
        RECT 2380.995 2052.035 2381.165 2052.625 ;
        RECT 2382.075 2052.435 2382.245 2052.795 ;
        RECT 2384.515 2052.775 2384.685 2053.105 ;
        RECT 2385.515 2052.775 2385.685 2053.105 ;
        RECT 2382.995 2052.605 2384.285 2052.685 ;
        RECT 2384.915 2052.605 2385.245 2052.685 ;
        RECT 2382.995 2052.515 2385.245 2052.605 ;
        RECT 2386.395 2052.515 2386.725 2052.685 ;
        RECT 2384.035 2052.435 2385.165 2052.515 ;
        RECT 2385.635 2052.345 2386.645 2052.515 ;
        RECT 2379.795 2051.865 2380.285 2052.035 ;
        RECT 2380.795 2051.865 2381.165 2052.035 ;
        RECT 2380.115 2051.785 2380.285 2051.865 ;
        RECT 2381.355 2051.785 2381.525 2052.115 ;
        RECT 2381.835 2051.785 2382.005 2052.235 ;
        RECT 2382.235 2051.865 2383.565 2052.035 ;
        RECT 2383.315 2051.785 2383.485 2051.865 ;
        RECT 2383.795 2051.785 2383.965 2052.115 ;
        RECT 2384.275 2051.785 2384.445 2052.235 ;
        RECT 2385.635 2052.115 2385.805 2052.345 ;
        RECT 2385.635 2051.865 2385.925 2052.115 ;
        RECT 2385.755 2051.785 2385.925 2051.865 ;
        RECT 2386.235 2051.785 2386.405 2052.115 ;
        RECT 2389.170 2051.895 2389.345 2053.155 ;
        RECT 2389.695 2052.095 2389.865 2053.155 ;
        RECT 2389.695 2051.925 2389.925 2052.095 ;
        RECT 2389.170 2051.695 2389.340 2051.895 ;
        RECT 2382.315 2051.635 2382.485 2051.675 ;
        RECT 2382.315 2051.465 2382.805 2051.635 ;
        RECT 2384.755 2051.505 2385.165 2051.675 ;
        RECT 2374.770 2051.035 2375.690 2051.205 ;
        RECT 2376.210 2051.040 2376.680 2051.210 ;
        RECT 2378.675 2051.045 2378.845 2051.395 ;
        RECT 2379.635 2051.045 2379.805 2051.395 ;
        RECT 2381.115 2051.045 2381.285 2051.395 ;
        RECT 2383.075 2051.045 2383.245 2051.395 ;
        RECT 2384.995 2051.045 2385.165 2051.505 ;
        RECT 2385.515 2051.045 2385.685 2051.395 ;
        RECT 2386.475 2051.295 2386.645 2051.395 ;
        RECT 2389.170 2051.365 2389.580 2051.695 ;
        RECT 2386.475 2051.125 2387.205 2051.295 ;
        RECT 2374.770 2050.885 2375.000 2051.035 ;
        RECT 2389.170 2050.855 2389.340 2051.365 ;
        RECT 2389.170 2050.525 2389.580 2050.855 ;
        RECT 2373.370 2050.145 2373.600 2050.315 ;
        RECT 2373.370 2049.865 2373.540 2050.145 ;
        RECT 2373.800 2049.865 2373.975 2050.375 ;
        RECT 2374.230 2049.865 2374.405 2050.415 ;
        RECT 2375.595 2049.865 2375.765 2050.375 ;
        RECT 2376.585 2049.870 2376.755 2050.380 ;
        RECT 2389.170 2050.355 2389.340 2050.525 ;
        RECT 2389.170 2049.865 2389.345 2050.355 ;
        RECT 2389.755 2050.315 2389.925 2051.925 ;
        RECT 2390.125 2051.895 2390.300 2053.155 ;
        RECT 2390.555 2052.015 2390.730 2053.155 ;
        RECT 2390.125 2050.945 2390.295 2051.895 ;
        RECT 2390.555 2050.415 2390.725 2052.015 ;
        RECT 2391.915 2052.010 2392.090 2053.155 ;
        RECT 2392.905 2052.015 2393.080 2053.160 ;
        RECT 2394.880 2052.905 2395.170 2053.075 ;
        RECT 2394.520 2052.345 2394.690 2052.765 ;
        RECT 2394.880 2052.035 2395.050 2052.905 ;
        RECT 2396.200 2052.625 2396.610 2052.795 ;
        RECT 2391.545 2051.205 2391.715 2051.895 ;
        RECT 2391.915 2051.795 2392.085 2052.010 ;
        RECT 2392.535 2051.795 2392.705 2051.900 ;
        RECT 2391.915 2051.625 2392.705 2051.795 ;
        RECT 2391.915 2051.575 2392.085 2051.625 ;
        RECT 2392.535 2051.210 2392.705 2051.625 ;
        RECT 2392.905 2051.580 2393.075 2052.015 ;
        RECT 2394.680 2051.865 2395.050 2052.035 ;
        RECT 2395.240 2052.345 2395.890 2052.515 ;
        RECT 2396.440 2052.435 2396.610 2052.625 ;
        RECT 2396.960 2052.345 2397.130 2052.765 ;
        RECT 2397.320 2052.625 2397.610 2052.795 ;
        RECT 2395.240 2051.785 2395.410 2052.345 ;
        RECT 2395.720 2051.785 2395.890 2052.115 ;
        RECT 2397.320 2052.035 2397.490 2052.625 ;
        RECT 2398.400 2052.435 2398.570 2052.795 ;
        RECT 2400.840 2052.775 2401.010 2053.105 ;
        RECT 2401.840 2052.775 2402.010 2053.105 ;
        RECT 2399.320 2052.605 2400.610 2052.685 ;
        RECT 2401.240 2052.605 2401.570 2052.685 ;
        RECT 2399.320 2052.515 2401.570 2052.605 ;
        RECT 2402.720 2052.515 2403.050 2052.685 ;
        RECT 2400.360 2052.435 2401.490 2052.515 ;
        RECT 2401.960 2052.345 2402.970 2052.515 ;
        RECT 2396.120 2051.865 2396.610 2052.035 ;
        RECT 2397.120 2051.865 2397.490 2052.035 ;
        RECT 2396.440 2051.785 2396.610 2051.865 ;
        RECT 2397.680 2051.785 2397.850 2052.115 ;
        RECT 2398.160 2051.785 2398.330 2052.235 ;
        RECT 2398.560 2051.865 2399.890 2052.035 ;
        RECT 2399.640 2051.785 2399.810 2051.865 ;
        RECT 2400.120 2051.785 2400.290 2052.115 ;
        RECT 2400.600 2051.785 2400.770 2052.235 ;
        RECT 2401.960 2052.115 2402.130 2052.345 ;
        RECT 2401.960 2051.865 2402.250 2052.115 ;
        RECT 2402.080 2051.785 2402.250 2051.865 ;
        RECT 2402.560 2051.785 2402.730 2052.115 ;
        RECT 2405.495 2051.895 2405.670 2053.155 ;
        RECT 2406.020 2052.095 2406.190 2053.155 ;
        RECT 2406.020 2051.925 2406.250 2052.095 ;
        RECT 2405.495 2051.695 2405.665 2051.895 ;
        RECT 2398.640 2051.635 2398.810 2051.675 ;
        RECT 2398.640 2051.465 2399.130 2051.635 ;
        RECT 2401.080 2051.505 2401.490 2051.675 ;
        RECT 2391.095 2051.035 2392.015 2051.205 ;
        RECT 2392.535 2051.040 2393.005 2051.210 ;
        RECT 2395.000 2051.045 2395.170 2051.395 ;
        RECT 2395.960 2051.045 2396.130 2051.395 ;
        RECT 2397.440 2051.045 2397.610 2051.395 ;
        RECT 2399.400 2051.045 2399.570 2051.395 ;
        RECT 2401.320 2051.045 2401.490 2051.505 ;
        RECT 2401.840 2051.045 2402.010 2051.395 ;
        RECT 2402.800 2051.295 2402.970 2051.395 ;
        RECT 2405.495 2051.365 2405.905 2051.695 ;
        RECT 2402.800 2051.125 2403.530 2051.295 ;
        RECT 2391.095 2050.885 2391.325 2051.035 ;
        RECT 2405.495 2050.855 2405.665 2051.365 ;
        RECT 2405.495 2050.525 2405.905 2050.855 ;
        RECT 2389.695 2050.145 2389.925 2050.315 ;
        RECT 2389.695 2049.865 2389.865 2050.145 ;
        RECT 2390.125 2049.865 2390.300 2050.375 ;
        RECT 2390.555 2049.865 2390.730 2050.415 ;
        RECT 2391.920 2049.865 2392.090 2050.375 ;
        RECT 2392.910 2049.870 2393.080 2050.380 ;
        RECT 2405.495 2050.355 2405.665 2050.525 ;
        RECT 2405.495 2049.865 2405.670 2050.355 ;
        RECT 2406.080 2050.315 2406.250 2051.925 ;
        RECT 2406.450 2051.895 2406.625 2053.155 ;
        RECT 2406.880 2052.015 2407.055 2053.155 ;
        RECT 2406.450 2050.945 2406.620 2051.895 ;
        RECT 2406.880 2050.415 2407.050 2052.015 ;
        RECT 2408.240 2052.010 2408.415 2053.155 ;
        RECT 2409.230 2052.015 2409.405 2053.160 ;
        RECT 2411.205 2052.905 2411.495 2053.075 ;
        RECT 2410.845 2052.345 2411.015 2052.765 ;
        RECT 2411.205 2052.035 2411.375 2052.905 ;
        RECT 2412.525 2052.625 2412.935 2052.795 ;
        RECT 2407.870 2051.205 2408.040 2051.895 ;
        RECT 2408.240 2051.795 2408.410 2052.010 ;
        RECT 2408.860 2051.795 2409.030 2051.900 ;
        RECT 2408.240 2051.625 2409.030 2051.795 ;
        RECT 2408.240 2051.575 2408.410 2051.625 ;
        RECT 2408.860 2051.210 2409.030 2051.625 ;
        RECT 2409.230 2051.580 2409.400 2052.015 ;
        RECT 2411.005 2051.865 2411.375 2052.035 ;
        RECT 2411.565 2052.345 2412.215 2052.515 ;
        RECT 2412.765 2052.435 2412.935 2052.625 ;
        RECT 2413.285 2052.345 2413.455 2052.765 ;
        RECT 2413.645 2052.625 2413.935 2052.795 ;
        RECT 2411.565 2051.785 2411.735 2052.345 ;
        RECT 2412.045 2051.785 2412.215 2052.115 ;
        RECT 2413.645 2052.035 2413.815 2052.625 ;
        RECT 2414.725 2052.435 2414.895 2052.795 ;
        RECT 2417.165 2052.775 2417.335 2053.105 ;
        RECT 2418.165 2052.775 2418.335 2053.105 ;
        RECT 2415.645 2052.605 2416.935 2052.685 ;
        RECT 2417.565 2052.605 2417.895 2052.685 ;
        RECT 2415.645 2052.515 2417.895 2052.605 ;
        RECT 2419.045 2052.515 2419.375 2052.685 ;
        RECT 2416.685 2052.435 2417.815 2052.515 ;
        RECT 2418.285 2052.345 2419.295 2052.515 ;
        RECT 2412.445 2051.865 2412.935 2052.035 ;
        RECT 2413.445 2051.865 2413.815 2052.035 ;
        RECT 2412.765 2051.785 2412.935 2051.865 ;
        RECT 2414.005 2051.785 2414.175 2052.115 ;
        RECT 2414.485 2051.785 2414.655 2052.235 ;
        RECT 2414.885 2051.865 2416.215 2052.035 ;
        RECT 2415.965 2051.785 2416.135 2051.865 ;
        RECT 2416.445 2051.785 2416.615 2052.115 ;
        RECT 2416.925 2051.785 2417.095 2052.235 ;
        RECT 2418.285 2052.115 2418.455 2052.345 ;
        RECT 2418.285 2051.865 2418.575 2052.115 ;
        RECT 2418.405 2051.785 2418.575 2051.865 ;
        RECT 2418.885 2051.785 2419.055 2052.115 ;
        RECT 2421.820 2051.895 2421.995 2053.155 ;
        RECT 2422.345 2052.095 2422.515 2053.155 ;
        RECT 2422.345 2051.925 2422.575 2052.095 ;
        RECT 2421.820 2051.695 2421.990 2051.895 ;
        RECT 2414.965 2051.635 2415.135 2051.675 ;
        RECT 2414.965 2051.465 2415.455 2051.635 ;
        RECT 2417.405 2051.505 2417.815 2051.675 ;
        RECT 2407.420 2051.035 2408.340 2051.205 ;
        RECT 2408.860 2051.040 2409.330 2051.210 ;
        RECT 2411.325 2051.045 2411.495 2051.395 ;
        RECT 2412.285 2051.045 2412.455 2051.395 ;
        RECT 2413.765 2051.045 2413.935 2051.395 ;
        RECT 2415.725 2051.045 2415.895 2051.395 ;
        RECT 2417.645 2051.045 2417.815 2051.505 ;
        RECT 2418.165 2051.045 2418.335 2051.395 ;
        RECT 2419.125 2051.295 2419.295 2051.395 ;
        RECT 2421.820 2051.365 2422.230 2051.695 ;
        RECT 2419.125 2051.125 2419.855 2051.295 ;
        RECT 2407.420 2050.885 2407.650 2051.035 ;
        RECT 2421.820 2050.855 2421.990 2051.365 ;
        RECT 2421.820 2050.525 2422.230 2050.855 ;
        RECT 2406.020 2050.145 2406.250 2050.315 ;
        RECT 2406.020 2049.865 2406.190 2050.145 ;
        RECT 2406.450 2049.865 2406.625 2050.375 ;
        RECT 2406.880 2049.865 2407.055 2050.415 ;
        RECT 2408.245 2049.865 2408.415 2050.375 ;
        RECT 2409.235 2049.870 2409.405 2050.380 ;
        RECT 2421.820 2050.355 2421.990 2050.525 ;
        RECT 2421.820 2049.865 2421.995 2050.355 ;
        RECT 2422.405 2050.315 2422.575 2051.925 ;
        RECT 2422.775 2051.895 2422.950 2053.155 ;
        RECT 2423.205 2052.015 2423.380 2053.155 ;
        RECT 2422.775 2050.945 2422.945 2051.895 ;
        RECT 2423.205 2050.415 2423.375 2052.015 ;
        RECT 2424.565 2052.010 2424.740 2053.155 ;
        RECT 2425.555 2052.015 2425.730 2053.160 ;
        RECT 2427.530 2052.905 2427.820 2053.075 ;
        RECT 2427.170 2052.345 2427.340 2052.765 ;
        RECT 2427.530 2052.035 2427.700 2052.905 ;
        RECT 2428.850 2052.625 2429.260 2052.795 ;
        RECT 2424.195 2051.205 2424.365 2051.895 ;
        RECT 2424.565 2051.795 2424.735 2052.010 ;
        RECT 2425.185 2051.795 2425.355 2051.900 ;
        RECT 2424.565 2051.625 2425.355 2051.795 ;
        RECT 2424.565 2051.575 2424.735 2051.625 ;
        RECT 2425.185 2051.210 2425.355 2051.625 ;
        RECT 2425.555 2051.580 2425.725 2052.015 ;
        RECT 2427.330 2051.865 2427.700 2052.035 ;
        RECT 2427.890 2052.345 2428.540 2052.515 ;
        RECT 2429.090 2052.435 2429.260 2052.625 ;
        RECT 2429.610 2052.345 2429.780 2052.765 ;
        RECT 2429.970 2052.625 2430.260 2052.795 ;
        RECT 2427.890 2051.785 2428.060 2052.345 ;
        RECT 2428.370 2051.785 2428.540 2052.115 ;
        RECT 2429.970 2052.035 2430.140 2052.625 ;
        RECT 2431.050 2052.435 2431.220 2052.795 ;
        RECT 2433.490 2052.775 2433.660 2053.105 ;
        RECT 2434.490 2052.775 2434.660 2053.105 ;
        RECT 2431.970 2052.605 2433.260 2052.685 ;
        RECT 2433.890 2052.605 2434.220 2052.685 ;
        RECT 2431.970 2052.515 2434.220 2052.605 ;
        RECT 2435.370 2052.515 2435.700 2052.685 ;
        RECT 2433.010 2052.435 2434.140 2052.515 ;
        RECT 2434.610 2052.345 2435.620 2052.515 ;
        RECT 2428.770 2051.865 2429.260 2052.035 ;
        RECT 2429.770 2051.865 2430.140 2052.035 ;
        RECT 2429.090 2051.785 2429.260 2051.865 ;
        RECT 2430.330 2051.785 2430.500 2052.115 ;
        RECT 2430.810 2051.785 2430.980 2052.235 ;
        RECT 2431.210 2051.865 2432.540 2052.035 ;
        RECT 2432.290 2051.785 2432.460 2051.865 ;
        RECT 2432.770 2051.785 2432.940 2052.115 ;
        RECT 2433.250 2051.785 2433.420 2052.235 ;
        RECT 2434.610 2052.115 2434.780 2052.345 ;
        RECT 2434.610 2051.865 2434.900 2052.115 ;
        RECT 2434.730 2051.785 2434.900 2051.865 ;
        RECT 2435.210 2051.785 2435.380 2052.115 ;
        RECT 2438.145 2051.895 2438.320 2053.155 ;
        RECT 2438.670 2052.095 2438.840 2053.155 ;
        RECT 2438.670 2051.925 2438.900 2052.095 ;
        RECT 2438.145 2051.695 2438.315 2051.895 ;
        RECT 2431.290 2051.635 2431.460 2051.675 ;
        RECT 2431.290 2051.465 2431.780 2051.635 ;
        RECT 2433.730 2051.505 2434.140 2051.675 ;
        RECT 2423.745 2051.035 2424.665 2051.205 ;
        RECT 2425.185 2051.040 2425.655 2051.210 ;
        RECT 2427.650 2051.045 2427.820 2051.395 ;
        RECT 2428.610 2051.045 2428.780 2051.395 ;
        RECT 2430.090 2051.045 2430.260 2051.395 ;
        RECT 2432.050 2051.045 2432.220 2051.395 ;
        RECT 2433.970 2051.045 2434.140 2051.505 ;
        RECT 2434.490 2051.045 2434.660 2051.395 ;
        RECT 2435.450 2051.295 2435.620 2051.395 ;
        RECT 2438.145 2051.365 2438.555 2051.695 ;
        RECT 2435.450 2051.125 2436.180 2051.295 ;
        RECT 2423.745 2050.885 2423.975 2051.035 ;
        RECT 2438.145 2050.855 2438.315 2051.365 ;
        RECT 2438.145 2050.525 2438.555 2050.855 ;
        RECT 2422.345 2050.145 2422.575 2050.315 ;
        RECT 2422.345 2049.865 2422.515 2050.145 ;
        RECT 2422.775 2049.865 2422.950 2050.375 ;
        RECT 2423.205 2049.865 2423.380 2050.415 ;
        RECT 2424.570 2049.865 2424.740 2050.375 ;
        RECT 2425.560 2049.870 2425.730 2050.380 ;
        RECT 2438.145 2050.355 2438.315 2050.525 ;
        RECT 2438.145 2049.865 2438.320 2050.355 ;
        RECT 2438.730 2050.315 2438.900 2051.925 ;
        RECT 2439.100 2051.895 2439.275 2053.155 ;
        RECT 2439.530 2052.015 2439.705 2053.155 ;
        RECT 2439.100 2050.945 2439.270 2051.895 ;
        RECT 2439.530 2050.415 2439.700 2052.015 ;
        RECT 2440.890 2052.010 2441.065 2053.155 ;
        RECT 2441.880 2052.015 2442.055 2053.160 ;
        RECT 2440.520 2051.205 2440.690 2051.895 ;
        RECT 2440.890 2051.795 2441.060 2052.010 ;
        RECT 2441.510 2051.795 2441.680 2051.900 ;
        RECT 2440.890 2051.625 2441.680 2051.795 ;
        RECT 2440.890 2051.575 2441.060 2051.625 ;
        RECT 2441.510 2051.210 2441.680 2051.625 ;
        RECT 2441.880 2051.580 2442.050 2052.015 ;
        RECT 2440.070 2051.035 2440.990 2051.205 ;
        RECT 2441.510 2051.040 2441.980 2051.210 ;
        RECT 2440.070 2050.885 2440.300 2051.035 ;
        RECT 2438.670 2050.145 2438.900 2050.315 ;
        RECT 2438.670 2049.865 2438.840 2050.145 ;
        RECT 2439.100 2049.865 2439.275 2050.375 ;
        RECT 2439.530 2049.865 2439.705 2050.415 ;
        RECT 2440.895 2049.865 2441.065 2050.375 ;
        RECT 2441.885 2049.870 2442.055 2050.380 ;
        RECT 2696.985 2036.335 2697.245 2036.665 ;
        RECT 2696.985 2035.425 2697.155 2036.335 ;
        RECT 2697.940 2036.265 2698.145 2036.665 ;
        RECT 2697.940 2036.095 2698.625 2036.265 ;
        RECT 2697.865 2035.425 2698.115 2035.925 ;
        RECT 2696.985 2035.255 2698.115 2035.425 ;
        RECT 2696.985 2034.485 2697.255 2035.255 ;
        RECT 2698.285 2035.065 2698.625 2036.095 ;
        RECT 2697.960 2034.890 2698.625 2035.065 ;
        RECT 2698.825 2036.160 2699.085 2036.665 ;
        RECT 2699.775 2036.285 2699.945 2036.665 ;
        RECT 2698.825 2035.360 2698.995 2036.160 ;
        RECT 2699.280 2036.115 2699.945 2036.285 ;
        RECT 2700.205 2036.160 2700.465 2036.665 ;
        RECT 2701.155 2036.285 2701.325 2036.665 ;
        RECT 2699.280 2035.860 2699.450 2036.115 ;
        RECT 2699.165 2035.530 2699.450 2035.860 ;
        RECT 2699.685 2035.565 2700.015 2035.935 ;
        RECT 2699.280 2035.385 2699.450 2035.530 ;
        RECT 2697.960 2034.485 2698.145 2034.890 ;
        RECT 2698.825 2034.455 2699.095 2035.360 ;
        RECT 2699.280 2035.215 2699.945 2035.385 ;
        RECT 2699.775 2034.455 2699.945 2035.215 ;
        RECT 2700.205 2035.360 2700.375 2036.160 ;
        RECT 2700.660 2036.115 2701.325 2036.285 ;
        RECT 2709.035 2036.285 2709.205 2036.665 ;
        RECT 2709.035 2036.115 2709.750 2036.285 ;
        RECT 2700.660 2035.860 2700.830 2036.115 ;
        RECT 2700.545 2035.530 2700.830 2035.860 ;
        RECT 2701.065 2035.565 2701.395 2035.935 ;
        RECT 2709.580 2035.925 2709.750 2036.115 ;
        RECT 2709.920 2036.090 2710.175 2036.665 ;
        RECT 2722.335 2036.265 2722.540 2036.665 ;
        RECT 2723.235 2036.335 2723.495 2036.665 ;
        RECT 2709.580 2035.595 2709.835 2035.925 ;
        RECT 2700.660 2035.385 2700.830 2035.530 ;
        RECT 2709.580 2035.385 2709.750 2035.595 ;
        RECT 2700.205 2034.455 2700.475 2035.360 ;
        RECT 2700.660 2035.215 2701.325 2035.385 ;
        RECT 2701.155 2034.455 2701.325 2035.215 ;
        RECT 2709.035 2035.215 2709.750 2035.385 ;
        RECT 2710.005 2035.360 2710.175 2036.090 ;
        RECT 2709.035 2034.455 2709.205 2035.215 ;
        RECT 2709.920 2034.455 2710.175 2035.360 ;
        RECT 2721.855 2036.095 2722.540 2036.265 ;
        RECT 2721.855 2035.065 2722.195 2036.095 ;
        RECT 2722.365 2035.425 2722.615 2035.925 ;
        RECT 2723.325 2035.425 2723.495 2036.335 ;
        RECT 2722.365 2035.255 2723.495 2035.425 ;
        RECT 2721.855 2034.890 2722.520 2035.065 ;
        RECT 2722.335 2034.485 2722.520 2034.890 ;
        RECT 2723.225 2034.485 2723.495 2035.255 ;
        RECT 2731.485 2036.160 2731.745 2036.665 ;
        RECT 2732.435 2036.285 2732.605 2036.665 ;
        RECT 2731.485 2035.360 2731.665 2036.160 ;
        RECT 2731.940 2036.115 2732.605 2036.285 ;
        RECT 2731.940 2035.860 2732.110 2036.115 ;
        RECT 2731.835 2035.530 2732.110 2035.860 ;
        RECT 2731.940 2035.385 2732.110 2035.530 ;
        RECT 2731.485 2034.455 2731.755 2035.360 ;
        RECT 2731.940 2035.215 2732.615 2035.385 ;
        RECT 2732.435 2034.455 2732.615 2035.215 ;
        RECT 2697.075 2033.185 2697.245 2033.945 ;
        RECT 2697.075 2033.015 2697.740 2033.185 ;
        RECT 2697.925 2033.040 2698.195 2033.945 ;
        RECT 2697.570 2032.870 2697.740 2033.015 ;
        RECT 2697.005 2032.465 2697.335 2032.835 ;
        RECT 2697.570 2032.540 2697.855 2032.870 ;
        RECT 2697.570 2032.285 2697.740 2032.540 ;
        RECT 2697.075 2032.115 2697.740 2032.285 ;
        RECT 2698.025 2032.240 2698.195 2033.040 ;
        RECT 2697.075 2031.735 2697.245 2032.115 ;
        RECT 2697.935 2031.735 2698.195 2032.240 ;
        RECT 2697.075 2025.405 2697.245 2025.785 ;
        RECT 2697.075 2025.235 2697.740 2025.405 ;
        RECT 2697.935 2025.280 2698.195 2025.785 ;
        RECT 2697.005 2024.685 2697.335 2025.055 ;
        RECT 2697.570 2024.980 2697.740 2025.235 ;
        RECT 2697.570 2024.650 2697.855 2024.980 ;
        RECT 2697.570 2024.505 2697.740 2024.650 ;
        RECT 2697.075 2024.335 2697.740 2024.505 ;
        RECT 2698.025 2024.480 2698.195 2025.280 ;
        RECT 2697.075 2023.575 2697.245 2024.335 ;
        RECT 2697.925 2023.575 2698.195 2024.480 ;
        RECT 2697.075 2019.965 2697.245 2020.340 ;
        RECT 2697.915 2020.175 2698.990 2020.345 ;
        RECT 2697.915 2019.965 2698.085 2020.175 ;
        RECT 2697.075 2019.795 2698.085 2019.965 ;
        RECT 2698.310 2019.835 2698.650 2020.005 ;
        RECT 2698.820 2019.840 2698.990 2020.175 ;
        RECT 2700.280 2020.175 2701.880 2020.345 ;
        RECT 2698.310 2019.665 2698.600 2019.835 ;
        RECT 2697.050 2019.495 2697.395 2019.605 ;
        RECT 2697.045 2019.325 2697.395 2019.495 ;
        RECT 2697.050 2018.985 2697.395 2019.325 ;
        RECT 2697.705 2018.985 2698.140 2019.605 ;
        RECT 2698.310 2019.145 2698.480 2019.665 ;
        RECT 2699.160 2019.495 2699.520 2020.170 ;
        RECT 2700.280 2019.805 2700.450 2020.175 ;
        RECT 2701.525 2020.135 2701.880 2020.175 ;
        RECT 2700.620 2019.755 2700.950 2020.005 ;
        RECT 2700.635 2019.680 2700.950 2019.755 ;
        RECT 2701.120 2019.885 2701.290 2020.005 ;
        RECT 2702.395 2019.885 2702.640 2020.305 ;
        RECT 2703.410 2019.945 2703.585 2020.275 ;
        RECT 2703.930 2020.185 2704.100 2020.345 ;
        RECT 2703.930 2020.015 2704.460 2020.185 ;
        RECT 2704.630 2020.175 2705.625 2020.345 ;
        RECT 2704.630 2020.015 2704.800 2020.175 ;
        RECT 2701.120 2019.715 2702.640 2019.885 ;
        RECT 2698.980 2019.315 2699.520 2019.495 ;
        RECT 2699.160 2019.205 2699.520 2019.315 ;
        RECT 2698.310 2018.975 2698.945 2019.145 ;
        RECT 2699.160 2018.975 2699.965 2019.205 ;
        RECT 2697.075 2018.635 2698.605 2018.805 ;
        RECT 2697.075 2018.135 2697.245 2018.635 ;
        RECT 2698.435 2018.475 2698.605 2018.635 ;
        RECT 2698.775 2018.645 2698.945 2018.975 ;
        RECT 2698.775 2018.475 2699.105 2018.645 ;
        RECT 2697.915 2018.305 2698.085 2018.465 ;
        RECT 2699.275 2018.305 2699.445 2018.805 ;
        RECT 2697.915 2018.135 2699.445 2018.305 ;
        RECT 2699.615 2018.135 2699.965 2018.975 ;
        RECT 2700.165 2018.605 2700.465 2019.605 ;
        RECT 2700.635 2019.155 2700.805 2019.680 ;
        RECT 2701.120 2019.675 2701.290 2019.715 ;
        RECT 2700.975 2019.495 2701.305 2019.505 ;
        RECT 2700.975 2019.335 2701.360 2019.495 ;
        RECT 2701.190 2019.325 2701.360 2019.335 ;
        RECT 2701.700 2019.155 2701.945 2019.545 ;
        RECT 2700.635 2018.985 2701.395 2019.155 ;
        RECT 2701.645 2018.985 2701.945 2019.155 ;
        RECT 2700.725 2018.305 2700.895 2018.815 ;
        RECT 2701.065 2018.475 2701.395 2018.985 ;
        RECT 2701.700 2018.925 2701.945 2018.985 ;
        RECT 2702.150 2018.925 2702.480 2019.545 ;
        RECT 2702.955 2018.925 2703.245 2019.605 ;
        RECT 2703.415 2019.495 2703.585 2019.945 ;
        RECT 2703.880 2019.665 2704.120 2019.835 ;
        RECT 2703.415 2019.325 2703.705 2019.495 ;
        RECT 2701.565 2018.515 2702.630 2018.685 ;
        RECT 2701.565 2018.305 2701.735 2018.515 ;
        RECT 2700.725 2018.135 2701.735 2018.305 ;
        RECT 2702.460 2018.135 2702.630 2018.515 ;
        RECT 2703.415 2018.465 2703.585 2019.325 ;
        RECT 2703.400 2018.135 2703.585 2018.465 ;
        RECT 2703.880 2018.465 2704.050 2019.665 ;
        RECT 2704.290 2018.845 2704.460 2020.015 ;
        RECT 2705.110 2019.835 2705.285 2020.005 ;
        RECT 2704.870 2019.675 2705.285 2019.835 ;
        RECT 2705.455 2019.885 2705.625 2020.175 ;
        RECT 2705.455 2019.715 2706.025 2019.885 ;
        RECT 2704.870 2019.665 2705.280 2019.675 ;
        RECT 2705.090 2019.325 2705.545 2019.495 ;
        RECT 2705.855 2018.935 2706.025 2019.715 ;
        RECT 2704.290 2018.615 2705.075 2018.845 ;
        RECT 2704.745 2018.475 2705.075 2018.615 ;
        RECT 2705.375 2018.765 2706.025 2018.935 ;
        RECT 2703.880 2018.135 2704.090 2018.465 ;
        RECT 2704.260 2018.305 2704.590 2018.345 ;
        RECT 2705.375 2018.305 2705.545 2018.765 ;
        RECT 2704.260 2018.135 2705.545 2018.305 ;
        RECT 2706.215 2018.135 2706.475 2020.345 ;
        RECT 2697.075 2016.865 2697.245 2017.625 ;
        RECT 2697.075 2016.695 2697.740 2016.865 ;
        RECT 2697.925 2016.720 2698.195 2017.625 ;
        RECT 2697.570 2016.550 2697.740 2016.695 ;
        RECT 2697.005 2016.145 2697.335 2016.515 ;
        RECT 2697.570 2016.220 2697.855 2016.550 ;
        RECT 2697.570 2015.965 2697.740 2016.220 ;
        RECT 2697.075 2015.795 2697.740 2015.965 ;
        RECT 2698.025 2015.920 2698.195 2016.720 ;
        RECT 2697.075 2015.415 2697.245 2015.795 ;
        RECT 2697.935 2015.415 2698.195 2015.920 ;
        RECT 2697.075 2014.525 2697.245 2014.900 ;
        RECT 2697.915 2014.735 2698.990 2014.905 ;
        RECT 2697.915 2014.525 2698.085 2014.735 ;
        RECT 2697.075 2014.355 2698.085 2014.525 ;
        RECT 2698.310 2014.395 2698.650 2014.565 ;
        RECT 2698.820 2014.400 2698.990 2014.735 ;
        RECT 2700.280 2014.735 2701.880 2014.905 ;
        RECT 2698.310 2014.225 2698.600 2014.395 ;
        RECT 2697.050 2014.055 2697.395 2014.165 ;
        RECT 2697.045 2013.885 2697.395 2014.055 ;
        RECT 2697.050 2013.545 2697.395 2013.885 ;
        RECT 2697.705 2013.545 2698.140 2014.165 ;
        RECT 2698.310 2013.705 2698.480 2014.225 ;
        RECT 2699.160 2014.055 2699.520 2014.730 ;
        RECT 2700.280 2014.365 2700.450 2014.735 ;
        RECT 2701.525 2014.695 2701.880 2014.735 ;
        RECT 2700.620 2014.315 2700.950 2014.565 ;
        RECT 2700.635 2014.240 2700.950 2014.315 ;
        RECT 2701.120 2014.445 2701.290 2014.565 ;
        RECT 2702.395 2014.445 2702.640 2014.865 ;
        RECT 2703.410 2014.505 2703.585 2014.835 ;
        RECT 2703.930 2014.745 2704.100 2014.905 ;
        RECT 2703.930 2014.575 2704.460 2014.745 ;
        RECT 2704.630 2014.735 2705.625 2014.905 ;
        RECT 2704.630 2014.575 2704.800 2014.735 ;
        RECT 2701.120 2014.275 2702.640 2014.445 ;
        RECT 2698.980 2013.875 2699.520 2014.055 ;
        RECT 2699.160 2013.765 2699.520 2013.875 ;
        RECT 2698.310 2013.535 2698.945 2013.705 ;
        RECT 2699.160 2013.535 2699.965 2013.765 ;
        RECT 2697.075 2013.195 2698.605 2013.365 ;
        RECT 2697.075 2012.695 2697.245 2013.195 ;
        RECT 2698.435 2013.035 2698.605 2013.195 ;
        RECT 2698.775 2013.205 2698.945 2013.535 ;
        RECT 2698.775 2013.035 2699.105 2013.205 ;
        RECT 2697.915 2012.865 2698.085 2013.025 ;
        RECT 2699.275 2012.865 2699.445 2013.365 ;
        RECT 2697.915 2012.695 2699.445 2012.865 ;
        RECT 2699.615 2012.695 2699.965 2013.535 ;
        RECT 2700.165 2013.165 2700.465 2014.165 ;
        RECT 2700.635 2013.715 2700.805 2014.240 ;
        RECT 2701.120 2014.235 2701.290 2014.275 ;
        RECT 2700.975 2014.055 2701.305 2014.065 ;
        RECT 2700.975 2013.895 2701.360 2014.055 ;
        RECT 2701.190 2013.885 2701.360 2013.895 ;
        RECT 2701.700 2013.715 2701.945 2014.105 ;
        RECT 2700.635 2013.545 2701.395 2013.715 ;
        RECT 2701.645 2013.545 2701.945 2013.715 ;
        RECT 2700.725 2012.865 2700.895 2013.375 ;
        RECT 2701.065 2013.035 2701.395 2013.545 ;
        RECT 2701.700 2013.485 2701.945 2013.545 ;
        RECT 2702.150 2013.485 2702.480 2014.105 ;
        RECT 2702.955 2013.485 2703.245 2014.165 ;
        RECT 2703.415 2014.055 2703.585 2014.505 ;
        RECT 2703.880 2014.225 2704.120 2014.395 ;
        RECT 2703.415 2013.885 2703.705 2014.055 ;
        RECT 2701.565 2013.075 2702.630 2013.245 ;
        RECT 2701.565 2012.865 2701.735 2013.075 ;
        RECT 2700.725 2012.695 2701.735 2012.865 ;
        RECT 2702.460 2012.695 2702.630 2013.075 ;
        RECT 2703.415 2013.025 2703.585 2013.885 ;
        RECT 2703.400 2012.695 2703.585 2013.025 ;
        RECT 2703.880 2013.025 2704.050 2014.225 ;
        RECT 2704.290 2013.405 2704.460 2014.575 ;
        RECT 2705.110 2014.395 2705.285 2014.565 ;
        RECT 2704.870 2014.235 2705.285 2014.395 ;
        RECT 2705.455 2014.445 2705.625 2014.735 ;
        RECT 2705.455 2014.275 2706.025 2014.445 ;
        RECT 2704.870 2014.225 2705.280 2014.235 ;
        RECT 2705.090 2013.885 2705.545 2014.055 ;
        RECT 2705.855 2013.495 2706.025 2014.275 ;
        RECT 2704.290 2013.175 2705.075 2013.405 ;
        RECT 2704.745 2013.035 2705.075 2013.175 ;
        RECT 2705.375 2013.325 2706.025 2013.495 ;
        RECT 2703.880 2012.695 2704.090 2013.025 ;
        RECT 2704.260 2012.865 2704.590 2012.905 ;
        RECT 2705.375 2012.865 2705.545 2013.325 ;
        RECT 2704.260 2012.695 2705.545 2012.865 ;
        RECT 2706.215 2012.695 2706.475 2014.905 ;
        RECT 2697.075 2011.425 2697.245 2012.185 ;
        RECT 2697.075 2011.255 2697.740 2011.425 ;
        RECT 2697.925 2011.280 2698.195 2012.185 ;
        RECT 2697.570 2011.110 2697.740 2011.255 ;
        RECT 2697.005 2010.705 2697.335 2011.075 ;
        RECT 2697.570 2010.780 2697.855 2011.110 ;
        RECT 2697.570 2010.525 2697.740 2010.780 ;
        RECT 2697.075 2010.355 2697.740 2010.525 ;
        RECT 2698.025 2010.480 2698.195 2011.280 ;
        RECT 2697.075 2009.975 2697.245 2010.355 ;
        RECT 2697.935 2009.975 2698.195 2010.480 ;
        RECT 2701.590 2011.215 2701.925 2012.185 ;
        RECT 2702.435 2012.015 2704.465 2012.185 ;
        RECT 2701.590 2010.545 2701.760 2011.215 ;
        RECT 2702.435 2011.045 2702.605 2012.015 ;
        RECT 2701.930 2010.715 2702.185 2011.045 ;
        RECT 2702.410 2010.715 2702.605 2011.045 ;
        RECT 2702.775 2011.675 2703.900 2011.845 ;
        RECT 2702.015 2010.545 2702.185 2010.715 ;
        RECT 2702.775 2010.545 2702.945 2011.675 ;
        RECT 2701.590 2009.975 2701.845 2010.545 ;
        RECT 2702.015 2010.375 2702.945 2010.545 ;
        RECT 2703.115 2011.335 2704.125 2011.505 ;
        RECT 2703.115 2010.535 2703.285 2011.335 ;
        RECT 2703.490 2010.655 2703.765 2011.135 ;
        RECT 2703.485 2010.485 2703.765 2010.655 ;
        RECT 2702.770 2010.340 2702.945 2010.375 ;
        RECT 2702.770 2009.975 2703.300 2010.340 ;
        RECT 2703.490 2009.975 2703.765 2010.485 ;
        RECT 2703.935 2009.975 2704.125 2011.335 ;
        RECT 2704.295 2011.350 2704.465 2012.015 ;
        RECT 2705.040 2011.595 2705.555 2012.005 ;
        RECT 2704.295 2011.160 2705.045 2011.350 ;
        RECT 2705.215 2010.785 2705.555 2011.595 ;
        RECT 2704.325 2010.615 2705.555 2010.785 ;
        RECT 2705.035 2010.010 2705.280 2010.615 ;
        RECT 2697.075 2005.985 2697.245 2006.745 ;
        RECT 2697.075 2005.815 2697.740 2005.985 ;
        RECT 2697.925 2005.840 2698.195 2006.745 ;
        RECT 2697.570 2005.670 2697.740 2005.815 ;
        RECT 2697.005 2005.265 2697.335 2005.635 ;
        RECT 2697.570 2005.340 2697.855 2005.670 ;
        RECT 2697.570 2005.085 2697.740 2005.340 ;
        RECT 2697.075 2004.915 2697.740 2005.085 ;
        RECT 2698.025 2005.040 2698.195 2005.840 ;
        RECT 2697.075 2004.535 2697.245 2004.915 ;
        RECT 2697.935 2004.535 2698.195 2005.040 ;
        RECT 2701.595 2000.505 2701.925 2001.290 ;
        RECT 2701.595 2000.335 2702.275 2000.505 ;
        RECT 2701.585 1999.915 2701.935 2000.165 ;
        RECT 2702.105 1999.735 2702.275 2000.335 ;
        RECT 2702.445 1999.915 2702.795 2000.165 ;
        RECT 2702.015 1999.095 2702.345 1999.735 ;
        RECT 2697.075 1998.205 2697.245 1998.585 ;
        RECT 2697.075 1998.035 2697.740 1998.205 ;
        RECT 2697.935 1998.080 2698.195 1998.585 ;
        RECT 2697.005 1997.485 2697.335 1997.855 ;
        RECT 2697.570 1997.780 2697.740 1998.035 ;
        RECT 2697.570 1997.450 2697.855 1997.780 ;
        RECT 2697.570 1997.305 2697.740 1997.450 ;
        RECT 2697.075 1997.135 2697.740 1997.305 ;
        RECT 2698.025 1997.280 2698.195 1998.080 ;
        RECT 2702.565 1998.225 2702.885 1998.585 ;
        RECT 2703.880 1998.225 2704.225 1998.585 ;
        RECT 2702.565 1998.055 2704.225 1998.225 ;
        RECT 2697.075 1996.375 2697.245 1997.135 ;
        RECT 2697.925 1996.375 2698.195 1997.280 ;
        RECT 2702.105 1997.215 2702.380 1997.845 ;
        RECT 2702.090 1996.555 2702.395 1997.045 ;
        RECT 2702.565 1996.725 2702.865 1998.055 ;
        RECT 2703.245 1997.595 2703.575 1997.765 ;
        RECT 2703.250 1997.345 2703.575 1997.595 ;
        RECT 2703.755 1997.515 2704.365 1997.845 ;
        RECT 2704.535 1997.345 2705.035 1997.805 ;
        RECT 2703.250 1997.165 2705.035 1997.345 ;
        RECT 2703.035 1996.815 2705.070 1996.985 ;
        RECT 2703.035 1996.555 2703.365 1996.815 ;
        RECT 2702.090 1996.375 2703.365 1996.555 ;
        RECT 2703.960 1996.735 2705.070 1996.815 ;
        RECT 2703.960 1996.375 2704.130 1996.735 ;
        RECT 2704.810 1996.375 2705.070 1996.735 ;
        RECT 2725.935 1995.015 2726.265 1995.865 ;
        RECT 2726.775 1995.015 2727.105 1995.865 ;
        RECT 2725.935 1994.845 2727.435 1995.015 ;
        RECT 2725.555 1994.475 2727.080 1994.675 ;
        RECT 2727.260 1994.645 2727.435 1994.845 ;
        RECT 2727.260 1994.475 2729.885 1994.645 ;
        RECT 2727.260 1994.305 2727.435 1994.475 ;
        RECT 2726.015 1994.135 2727.435 1994.305 ;
        RECT 2726.015 1993.655 2726.185 1994.135 ;
        RECT 2726.855 1993.660 2727.025 1994.135 ;
        RECT 2697.075 1992.765 2697.245 1993.145 ;
        RECT 2697.075 1992.595 2697.740 1992.765 ;
        RECT 2697.935 1992.640 2698.195 1993.145 ;
        RECT 2697.005 1992.045 2697.335 1992.415 ;
        RECT 2697.570 1992.340 2697.740 1992.595 ;
        RECT 2697.570 1992.010 2697.855 1992.340 ;
        RECT 2697.570 1991.865 2697.740 1992.010 ;
        RECT 2697.075 1991.695 2697.740 1991.865 ;
        RECT 2698.025 1991.840 2698.195 1992.640 ;
        RECT 2697.075 1990.935 2697.245 1991.695 ;
        RECT 2697.925 1990.935 2698.195 1991.840 ;
        RECT 2697.310 1987.305 2697.480 1987.555 ;
        RECT 2696.985 1987.135 2697.480 1987.305 ;
        RECT 2698.215 1987.305 2698.385 1987.650 ;
        RECT 2699.055 1987.305 2699.575 1987.705 ;
        RECT 2698.215 1987.135 2699.575 1987.305 ;
        RECT 2696.985 1986.175 2697.155 1987.135 ;
        RECT 2697.325 1986.345 2697.675 1986.965 ;
        RECT 2697.845 1986.345 2698.185 1986.965 ;
        RECT 2698.355 1986.345 2698.595 1986.965 ;
        RECT 2698.775 1986.715 2699.235 1986.885 ;
        RECT 2698.775 1986.175 2698.945 1986.715 ;
        RECT 2699.405 1986.515 2699.575 1987.135 ;
        RECT 2696.985 1986.005 2698.945 1986.175 ;
        RECT 2699.115 1985.505 2699.575 1986.515 ;
        RECT 2697.075 1984.225 2697.245 1984.985 ;
        RECT 2522.640 1981.955 2523.160 1983.440 ;
        RECT 2523.330 1982.615 2523.850 1984.165 ;
        RECT 2697.075 1984.055 2697.740 1984.225 ;
        RECT 2697.925 1984.080 2698.195 1984.985 ;
        RECT 2697.570 1983.910 2697.740 1984.055 ;
        RECT 2697.005 1983.505 2697.335 1983.875 ;
        RECT 2697.570 1983.580 2697.855 1983.910 ;
        RECT 2697.570 1983.325 2697.740 1983.580 ;
        RECT 2697.075 1983.155 2697.740 1983.325 ;
        RECT 2698.025 1983.280 2698.195 1984.080 ;
        RECT 2697.075 1982.775 2697.245 1983.155 ;
        RECT 2697.935 1982.775 2698.195 1983.280 ;
        RECT 2697.260 1981.625 2697.505 1982.230 ;
        RECT 2696.985 1981.455 2698.215 1981.625 ;
        RECT 2696.985 1980.645 2697.325 1981.455 ;
        RECT 2697.495 1980.890 2698.245 1981.080 ;
        RECT 2696.985 1980.235 2697.500 1980.645 ;
        RECT 2698.075 1980.225 2698.245 1980.890 ;
        RECT 2698.415 1980.905 2698.605 1982.265 ;
        RECT 2698.775 1982.095 2699.050 1982.265 ;
        RECT 2698.775 1981.925 2699.055 1982.095 ;
        RECT 2698.775 1981.105 2699.050 1981.925 ;
        RECT 2699.240 1981.900 2699.770 1982.265 ;
        RECT 2699.595 1981.865 2699.770 1981.900 ;
        RECT 2699.255 1980.905 2699.425 1981.705 ;
        RECT 2698.415 1980.735 2699.425 1980.905 ;
        RECT 2699.595 1981.695 2700.525 1981.865 ;
        RECT 2700.695 1981.695 2700.950 1982.265 ;
        RECT 2699.595 1980.565 2699.765 1981.695 ;
        RECT 2700.355 1981.525 2700.525 1981.695 ;
        RECT 2698.640 1980.395 2699.765 1980.565 ;
        RECT 2699.935 1981.195 2700.130 1981.525 ;
        RECT 2700.355 1981.195 2700.610 1981.525 ;
        RECT 2699.935 1980.225 2700.105 1981.195 ;
        RECT 2700.780 1981.025 2700.950 1981.695 ;
        RECT 2701.630 1981.500 2701.815 1982.170 ;
        RECT 2702.300 1981.815 2702.630 1982.215 ;
        RECT 2703.345 1981.820 2703.675 1982.260 ;
        RECT 2703.345 1981.815 2704.575 1981.820 ;
        RECT 2702.300 1981.705 2704.575 1981.815 ;
        RECT 2702.420 1981.640 2704.575 1981.705 ;
        RECT 2701.180 1981.230 2701.815 1981.500 ;
        RECT 2701.995 1981.120 2702.280 1981.525 ;
        RECT 2702.450 1981.120 2702.780 1981.470 ;
        RECT 2698.075 1980.055 2700.105 1980.225 ;
        RECT 2700.615 1980.055 2700.950 1981.025 ;
        RECT 2701.215 1980.770 2702.325 1980.940 ;
        RECT 2701.215 1980.060 2701.410 1980.770 ;
        RECT 2702.095 1980.060 2702.325 1980.770 ;
        RECT 2702.505 1980.065 2702.780 1981.120 ;
        RECT 2702.950 1980.065 2703.285 1981.470 ;
        RECT 2703.485 1980.065 2703.935 1981.470 ;
        RECT 2704.190 1980.060 2704.575 1981.640 ;
        RECT 2696.985 1978.155 2697.325 1979.035 ;
        RECT 2697.495 1978.325 2697.665 1979.545 ;
        RECT 2698.690 1979.205 2699.165 1979.545 ;
        RECT 2697.905 1978.675 2698.155 1979.040 ;
        RECT 2698.875 1978.675 2699.590 1978.970 ;
        RECT 2699.760 1978.845 2700.035 1979.545 ;
        RECT 2697.905 1978.505 2699.695 1978.675 ;
        RECT 2697.495 1978.075 2698.290 1978.325 ;
        RECT 2697.495 1977.985 2697.745 1978.075 ;
        RECT 2697.415 1977.565 2697.745 1977.985 ;
        RECT 2698.460 1977.650 2698.715 1978.505 ;
        RECT 2697.925 1977.385 2698.715 1977.650 ;
        RECT 2698.885 1977.805 2699.295 1978.325 ;
        RECT 2699.465 1978.075 2699.695 1978.505 ;
        RECT 2699.865 1977.815 2700.035 1978.845 ;
        RECT 2698.885 1977.385 2699.085 1977.805 ;
        RECT 2699.775 1977.335 2700.035 1977.815 ;
        RECT 2522.640 1974.425 2523.160 1975.910 ;
        RECT 2523.330 1975.085 2523.850 1976.635 ;
        RECT 2697.075 1976.445 2697.245 1976.825 ;
        RECT 2697.075 1976.275 2697.740 1976.445 ;
        RECT 2697.935 1976.320 2698.195 1976.825 ;
        RECT 2697.005 1975.725 2697.335 1976.095 ;
        RECT 2697.570 1976.020 2697.740 1976.275 ;
        RECT 2697.570 1975.690 2697.855 1976.020 ;
        RECT 2697.570 1975.545 2697.740 1975.690 ;
        RECT 2697.075 1975.375 2697.740 1975.545 ;
        RECT 2698.025 1975.520 2698.195 1976.320 ;
        RECT 2697.075 1974.615 2697.245 1975.375 ;
        RECT 2697.925 1974.615 2698.195 1975.520 ;
        RECT 2698.455 1973.605 2698.625 1974.105 ;
        RECT 2699.415 1973.605 2699.585 1974.105 ;
        RECT 2700.255 1973.605 2700.425 1974.105 ;
        RECT 2698.455 1973.435 2700.425 1973.605 ;
        RECT 2700.595 1973.635 2700.925 1974.065 ;
        RECT 2701.535 1973.805 2701.875 1974.065 ;
        RECT 2700.595 1973.465 2701.445 1973.635 ;
        RECT 2698.390 1972.635 2698.645 1973.265 ;
        RECT 2698.875 1972.635 2699.255 1973.265 ;
        RECT 2700.125 1973.255 2700.425 1973.260 ;
        RECT 2700.125 1973.085 2700.435 1973.255 ;
        RECT 2700.125 1972.965 2700.425 1973.085 ;
        RECT 2698.875 1972.035 2699.080 1972.635 ;
        RECT 2699.515 1972.240 2699.735 1972.965 ;
        RECT 2700.045 1972.635 2700.425 1972.965 ;
        RECT 2700.625 1972.715 2700.955 1973.275 ;
        RECT 2701.275 1972.545 2701.445 1973.465 ;
        RECT 2700.625 1972.450 2701.445 1972.545 ;
        RECT 2700.430 1972.375 2701.445 1972.450 ;
        RECT 2699.310 1972.055 2700.260 1972.240 ;
        RECT 2700.430 1971.940 2700.845 1972.375 ;
        RECT 2701.615 1972.200 2701.875 1973.805 ;
        RECT 2701.535 1971.940 2701.875 1972.200 ;
        RECT 2698.335 1970.735 2698.665 1971.155 ;
        RECT 2698.845 1970.985 2699.105 1971.385 ;
        RECT 2699.775 1970.985 2699.945 1971.335 ;
        RECT 2698.845 1970.815 2700.510 1970.985 ;
        RECT 2700.680 1970.880 2700.955 1971.225 ;
        RECT 2522.640 1968.445 2523.160 1969.930 ;
        RECT 2523.330 1969.105 2523.850 1970.655 ;
        RECT 2698.415 1970.645 2698.665 1970.735 ;
        RECT 2700.340 1970.645 2700.510 1970.815 ;
        RECT 2697.910 1970.315 2698.245 1970.565 ;
        RECT 2698.415 1970.315 2699.130 1970.645 ;
        RECT 2699.345 1970.315 2700.170 1970.645 ;
        RECT 2700.340 1970.315 2700.615 1970.645 ;
        RECT 2698.415 1969.755 2698.585 1970.315 ;
        RECT 2698.845 1969.855 2699.175 1970.145 ;
        RECT 2699.345 1970.025 2699.590 1970.315 ;
        RECT 2700.340 1970.145 2700.510 1970.315 ;
        RECT 2700.785 1970.145 2700.955 1970.880 ;
        RECT 2699.850 1969.975 2700.510 1970.145 ;
        RECT 2699.850 1969.855 2700.020 1969.975 ;
        RECT 2698.845 1969.685 2700.020 1969.855 ;
        RECT 2698.405 1969.185 2700.020 1969.515 ;
        RECT 2700.680 1969.175 2700.955 1970.145 ;
        RECT 2701.125 1971.155 2701.715 1971.385 ;
        RECT 2701.125 1970.145 2701.415 1971.155 ;
        RECT 2703.290 1970.985 2703.715 1971.195 ;
        RECT 2701.585 1970.815 2703.715 1970.985 ;
        RECT 2701.585 1970.315 2701.755 1970.815 ;
        RECT 2702.045 1970.315 2702.375 1970.645 ;
        RECT 2702.565 1970.315 2702.835 1970.645 ;
        RECT 2703.025 1970.315 2703.375 1970.645 ;
        RECT 2701.125 1969.975 2702.670 1970.145 ;
        RECT 2703.545 1970.045 2703.715 1970.815 ;
        RECT 2701.125 1969.175 2701.715 1969.975 ;
        RECT 2702.340 1969.175 2702.670 1969.975 ;
        RECT 2703.290 1969.715 2703.715 1970.045 ;
        RECT 2697.075 1967.905 2697.245 1968.665 ;
        RECT 2697.075 1967.735 2697.740 1967.905 ;
        RECT 2697.925 1967.760 2698.195 1968.665 ;
        RECT 2697.570 1967.590 2697.740 1967.735 ;
        RECT 2697.005 1967.185 2697.335 1967.555 ;
        RECT 2697.570 1967.260 2697.855 1967.590 ;
        RECT 2697.570 1967.005 2697.740 1967.260 ;
        RECT 2697.075 1966.835 2697.740 1967.005 ;
        RECT 2698.025 1966.960 2698.195 1967.760 ;
        RECT 2699.255 1967.685 2699.585 1968.665 ;
        RECT 2698.845 1967.275 2699.180 1967.525 ;
        RECT 2699.350 1967.085 2699.520 1967.685 ;
        RECT 2699.690 1967.255 2700.025 1967.525 ;
        RECT 2697.075 1966.455 2697.245 1966.835 ;
        RECT 2697.935 1966.455 2698.195 1966.960 ;
        RECT 2698.825 1966.455 2699.520 1967.085 ;
        RECT 2697.260 1965.305 2697.505 1965.910 ;
        RECT 2696.985 1965.135 2698.215 1965.305 ;
        RECT 2522.640 1962.500 2523.160 1963.985 ;
        RECT 2523.330 1963.160 2523.850 1964.710 ;
        RECT 2696.985 1964.325 2697.325 1965.135 ;
        RECT 2697.495 1964.570 2698.245 1964.760 ;
        RECT 2696.985 1963.915 2697.500 1964.325 ;
        RECT 2698.075 1963.905 2698.245 1964.570 ;
        RECT 2698.415 1964.585 2698.605 1965.945 ;
        RECT 2698.775 1965.095 2699.050 1965.945 ;
        RECT 2699.240 1965.580 2699.770 1965.945 ;
        RECT 2699.595 1965.545 2699.770 1965.580 ;
        RECT 2698.775 1964.925 2699.055 1965.095 ;
        RECT 2698.775 1964.785 2699.050 1964.925 ;
        RECT 2699.255 1964.585 2699.425 1965.385 ;
        RECT 2698.415 1964.415 2699.425 1964.585 ;
        RECT 2699.595 1965.375 2700.525 1965.545 ;
        RECT 2700.695 1965.375 2700.950 1965.945 ;
        RECT 2699.595 1964.245 2699.765 1965.375 ;
        RECT 2700.355 1965.205 2700.525 1965.375 ;
        RECT 2698.640 1964.075 2699.765 1964.245 ;
        RECT 2699.935 1964.875 2700.130 1965.205 ;
        RECT 2700.355 1964.875 2700.610 1965.205 ;
        RECT 2699.935 1963.905 2700.105 1964.875 ;
        RECT 2700.780 1964.705 2700.950 1965.375 ;
        RECT 2698.075 1963.735 2700.105 1963.905 ;
        RECT 2700.615 1963.735 2700.950 1964.705 ;
        RECT 2697.075 1962.465 2697.245 1963.225 ;
        RECT 2697.075 1962.295 2697.740 1962.465 ;
        RECT 2697.925 1962.320 2698.195 1963.225 ;
        RECT 2697.570 1962.150 2697.740 1962.295 ;
        RECT 2697.005 1961.745 2697.335 1962.115 ;
        RECT 2697.570 1961.820 2697.855 1962.150 ;
        RECT 2697.570 1961.565 2697.740 1961.820 ;
        RECT 2697.075 1961.395 2697.740 1961.565 ;
        RECT 2698.025 1961.520 2698.195 1962.320 ;
        RECT 2697.075 1961.015 2697.245 1961.395 ;
        RECT 2697.935 1961.015 2698.195 1961.520 ;
        RECT 2522.640 1956.855 2523.160 1958.340 ;
        RECT 2523.330 1957.515 2523.850 1959.065 ;
        RECT 2697.075 1957.025 2697.245 1957.785 ;
        RECT 2697.075 1956.855 2697.740 1957.025 ;
        RECT 2697.925 1956.880 2698.195 1957.785 ;
        RECT 2697.570 1956.710 2697.740 1956.855 ;
        RECT 2697.005 1956.305 2697.335 1956.675 ;
        RECT 2697.570 1956.380 2697.855 1956.710 ;
        RECT 2697.570 1956.125 2697.740 1956.380 ;
        RECT 2697.075 1955.955 2697.740 1956.125 ;
        RECT 2698.025 1956.080 2698.195 1956.880 ;
        RECT 2697.075 1955.575 2697.245 1955.955 ;
        RECT 2697.935 1955.575 2698.195 1956.080 ;
        RECT 2358.650 1953.110 2358.825 1953.600 ;
        RECT 2359.175 1953.320 2359.345 1953.600 ;
        RECT 2359.175 1953.150 2359.405 1953.320 ;
        RECT 2358.650 1952.940 2358.820 1953.110 ;
        RECT 2358.650 1952.610 2359.060 1952.940 ;
        RECT 2358.650 1952.100 2358.820 1952.610 ;
        RECT 2358.650 1951.770 2359.060 1952.100 ;
        RECT 2358.650 1951.570 2358.820 1951.770 ;
        RECT 2358.650 1950.310 2358.825 1951.570 ;
        RECT 2359.235 1951.540 2359.405 1953.150 ;
        RECT 2359.605 1953.090 2359.780 1953.600 ;
        RECT 2369.465 1953.110 2369.640 1953.600 ;
        RECT 2369.465 1952.940 2369.635 1953.110 ;
        RECT 2370.420 1953.090 2370.595 1953.600 ;
        RECT 2370.850 1953.050 2371.025 1953.600 ;
        RECT 2375.080 1953.110 2375.255 1953.600 ;
        RECT 2375.605 1953.320 2375.775 1953.600 ;
        RECT 2375.605 1953.150 2375.835 1953.320 ;
        RECT 2369.465 1952.610 2369.875 1952.940 ;
        RECT 2359.175 1951.370 2359.405 1951.540 ;
        RECT 2359.605 1951.570 2359.775 1952.520 ;
        RECT 2369.465 1952.100 2369.635 1952.610 ;
        RECT 2369.465 1951.770 2369.875 1952.100 ;
        RECT 2369.465 1951.570 2369.635 1951.770 ;
        RECT 2370.420 1951.570 2370.590 1952.520 ;
        RECT 2359.175 1950.310 2359.345 1951.370 ;
        RECT 2359.605 1950.310 2359.780 1951.570 ;
        RECT 2369.465 1950.310 2369.640 1951.570 ;
        RECT 2370.420 1950.310 2370.595 1951.570 ;
        RECT 2370.850 1951.450 2371.020 1953.050 ;
        RECT 2375.080 1952.940 2375.250 1953.110 ;
        RECT 2375.080 1952.610 2375.490 1952.940 ;
        RECT 2375.080 1952.100 2375.250 1952.610 ;
        RECT 2375.080 1951.770 2375.490 1952.100 ;
        RECT 2375.080 1951.570 2375.250 1951.770 ;
        RECT 2370.850 1950.310 2371.025 1951.450 ;
        RECT 2375.080 1950.310 2375.255 1951.570 ;
        RECT 2375.665 1951.540 2375.835 1953.150 ;
        RECT 2376.035 1953.090 2376.210 1953.600 ;
        RECT 2376.465 1953.050 2376.640 1953.600 ;
        RECT 2377.830 1953.085 2378.000 1953.595 ;
        RECT 2378.820 1953.085 2378.990 1953.595 ;
        RECT 2388.025 1953.110 2388.200 1953.600 ;
        RECT 2375.605 1951.370 2375.835 1951.540 ;
        RECT 2376.035 1951.570 2376.205 1952.520 ;
        RECT 2375.605 1950.310 2375.775 1951.370 ;
        RECT 2376.035 1950.310 2376.210 1951.570 ;
        RECT 2376.465 1951.450 2376.635 1953.050 ;
        RECT 2388.025 1952.940 2388.195 1953.110 ;
        RECT 2388.980 1953.090 2389.155 1953.600 ;
        RECT 2389.410 1953.050 2389.585 1953.600 ;
        RECT 2393.640 1953.110 2393.815 1953.600 ;
        RECT 2394.165 1953.320 2394.335 1953.600 ;
        RECT 2394.165 1953.150 2394.395 1953.320 ;
        RECT 2377.395 1952.425 2377.625 1952.625 ;
        RECT 2388.025 1952.610 2388.435 1952.940 ;
        RECT 2377.395 1952.395 2377.925 1952.425 ;
        RECT 2377.455 1952.255 2377.925 1952.395 ;
        RECT 2378.445 1952.255 2378.915 1952.425 ;
        RECT 2377.455 1951.565 2377.625 1952.255 ;
        RECT 2377.825 1951.790 2377.995 1951.885 ;
        RECT 2378.445 1951.790 2378.615 1952.255 ;
        RECT 2388.025 1952.100 2388.195 1952.610 ;
        RECT 2377.825 1951.610 2378.615 1951.790 ;
        RECT 2376.465 1950.310 2376.640 1951.450 ;
        RECT 2377.825 1950.305 2378.000 1951.610 ;
        RECT 2378.445 1951.565 2378.615 1951.610 ;
        RECT 2378.815 1951.450 2378.985 1951.885 ;
        RECT 2388.025 1951.770 2388.435 1952.100 ;
        RECT 2388.025 1951.570 2388.195 1951.770 ;
        RECT 2388.980 1951.570 2389.150 1952.520 ;
        RECT 2378.815 1950.305 2378.990 1951.450 ;
        RECT 2388.025 1950.310 2388.200 1951.570 ;
        RECT 2388.980 1950.310 2389.155 1951.570 ;
        RECT 2389.410 1951.450 2389.580 1953.050 ;
        RECT 2393.640 1952.940 2393.810 1953.110 ;
        RECT 2393.640 1952.610 2394.050 1952.940 ;
        RECT 2393.640 1952.100 2393.810 1952.610 ;
        RECT 2393.640 1951.770 2394.050 1952.100 ;
        RECT 2393.640 1951.570 2393.810 1951.770 ;
        RECT 2389.410 1950.310 2389.585 1951.450 ;
        RECT 2393.640 1950.310 2393.815 1951.570 ;
        RECT 2394.225 1951.540 2394.395 1953.150 ;
        RECT 2394.595 1953.090 2394.770 1953.600 ;
        RECT 2395.025 1953.050 2395.200 1953.600 ;
        RECT 2396.390 1953.085 2396.560 1953.595 ;
        RECT 2397.380 1953.085 2397.550 1953.595 ;
        RECT 2406.585 1953.110 2406.760 1953.600 ;
        RECT 2394.165 1951.370 2394.395 1951.540 ;
        RECT 2394.595 1951.570 2394.765 1952.520 ;
        RECT 2394.165 1950.310 2394.335 1951.370 ;
        RECT 2394.595 1950.310 2394.770 1951.570 ;
        RECT 2395.025 1951.450 2395.195 1953.050 ;
        RECT 2406.585 1952.940 2406.755 1953.110 ;
        RECT 2407.540 1953.090 2407.715 1953.600 ;
        RECT 2407.970 1953.050 2408.145 1953.600 ;
        RECT 2412.200 1953.110 2412.375 1953.600 ;
        RECT 2412.725 1953.320 2412.895 1953.600 ;
        RECT 2412.725 1953.150 2412.955 1953.320 ;
        RECT 2395.955 1952.425 2396.185 1952.625 ;
        RECT 2406.585 1952.610 2406.995 1952.940 ;
        RECT 2395.955 1952.395 2396.485 1952.425 ;
        RECT 2396.015 1952.255 2396.485 1952.395 ;
        RECT 2397.005 1952.255 2397.475 1952.425 ;
        RECT 2396.015 1951.565 2396.185 1952.255 ;
        RECT 2396.385 1951.790 2396.555 1951.885 ;
        RECT 2397.005 1951.790 2397.175 1952.255 ;
        RECT 2406.585 1952.100 2406.755 1952.610 ;
        RECT 2396.385 1951.610 2397.175 1951.790 ;
        RECT 2395.025 1950.310 2395.200 1951.450 ;
        RECT 2396.385 1950.305 2396.560 1951.610 ;
        RECT 2397.005 1951.565 2397.175 1951.610 ;
        RECT 2397.375 1951.450 2397.545 1951.885 ;
        RECT 2406.585 1951.770 2406.995 1952.100 ;
        RECT 2406.585 1951.570 2406.755 1951.770 ;
        RECT 2407.540 1951.570 2407.710 1952.520 ;
        RECT 2397.375 1950.305 2397.550 1951.450 ;
        RECT 2406.585 1950.310 2406.760 1951.570 ;
        RECT 2407.540 1950.310 2407.715 1951.570 ;
        RECT 2407.970 1951.450 2408.140 1953.050 ;
        RECT 2412.200 1952.940 2412.370 1953.110 ;
        RECT 2412.200 1952.610 2412.610 1952.940 ;
        RECT 2412.200 1952.100 2412.370 1952.610 ;
        RECT 2412.200 1951.770 2412.610 1952.100 ;
        RECT 2412.200 1951.570 2412.370 1951.770 ;
        RECT 2407.970 1950.310 2408.145 1951.450 ;
        RECT 2412.200 1950.310 2412.375 1951.570 ;
        RECT 2412.785 1951.540 2412.955 1953.150 ;
        RECT 2413.155 1953.090 2413.330 1953.600 ;
        RECT 2413.585 1953.050 2413.760 1953.600 ;
        RECT 2414.950 1953.085 2415.120 1953.595 ;
        RECT 2415.940 1953.085 2416.110 1953.595 ;
        RECT 2425.145 1953.110 2425.320 1953.600 ;
        RECT 2412.725 1951.370 2412.955 1951.540 ;
        RECT 2413.155 1951.570 2413.325 1952.520 ;
        RECT 2412.725 1950.310 2412.895 1951.370 ;
        RECT 2413.155 1950.310 2413.330 1951.570 ;
        RECT 2413.585 1951.450 2413.755 1953.050 ;
        RECT 2425.145 1952.940 2425.315 1953.110 ;
        RECT 2426.100 1953.090 2426.275 1953.600 ;
        RECT 2426.530 1953.050 2426.705 1953.600 ;
        RECT 2430.760 1953.110 2430.935 1953.600 ;
        RECT 2431.285 1953.320 2431.455 1953.600 ;
        RECT 2431.285 1953.150 2431.515 1953.320 ;
        RECT 2414.515 1952.425 2414.745 1952.625 ;
        RECT 2425.145 1952.610 2425.555 1952.940 ;
        RECT 2414.515 1952.395 2415.045 1952.425 ;
        RECT 2414.575 1952.255 2415.045 1952.395 ;
        RECT 2415.565 1952.255 2416.035 1952.425 ;
        RECT 2414.575 1951.565 2414.745 1952.255 ;
        RECT 2414.945 1951.790 2415.115 1951.885 ;
        RECT 2415.565 1951.790 2415.735 1952.255 ;
        RECT 2425.145 1952.100 2425.315 1952.610 ;
        RECT 2414.945 1951.610 2415.735 1951.790 ;
        RECT 2413.585 1950.310 2413.760 1951.450 ;
        RECT 2414.945 1950.305 2415.120 1951.610 ;
        RECT 2415.565 1951.565 2415.735 1951.610 ;
        RECT 2415.935 1951.450 2416.105 1951.885 ;
        RECT 2425.145 1951.770 2425.555 1952.100 ;
        RECT 2425.145 1951.570 2425.315 1951.770 ;
        RECT 2426.100 1951.570 2426.270 1952.520 ;
        RECT 2415.935 1950.305 2416.110 1951.450 ;
        RECT 2425.145 1950.310 2425.320 1951.570 ;
        RECT 2426.100 1950.310 2426.275 1951.570 ;
        RECT 2426.530 1951.450 2426.700 1953.050 ;
        RECT 2430.760 1952.940 2430.930 1953.110 ;
        RECT 2430.760 1952.610 2431.170 1952.940 ;
        RECT 2430.760 1952.100 2430.930 1952.610 ;
        RECT 2430.760 1951.770 2431.170 1952.100 ;
        RECT 2430.760 1951.570 2430.930 1951.770 ;
        RECT 2426.530 1950.310 2426.705 1951.450 ;
        RECT 2430.760 1950.310 2430.935 1951.570 ;
        RECT 2431.345 1951.540 2431.515 1953.150 ;
        RECT 2431.715 1953.090 2431.890 1953.600 ;
        RECT 2432.145 1953.050 2432.320 1953.600 ;
        RECT 2433.510 1953.085 2433.680 1953.595 ;
        RECT 2434.500 1953.085 2434.670 1953.595 ;
        RECT 2443.705 1953.110 2443.880 1953.600 ;
        RECT 2431.285 1951.370 2431.515 1951.540 ;
        RECT 2431.715 1951.570 2431.885 1952.520 ;
        RECT 2431.285 1950.310 2431.455 1951.370 ;
        RECT 2431.715 1950.310 2431.890 1951.570 ;
        RECT 2432.145 1951.450 2432.315 1953.050 ;
        RECT 2443.705 1952.940 2443.875 1953.110 ;
        RECT 2444.660 1953.090 2444.835 1953.600 ;
        RECT 2445.090 1953.050 2445.265 1953.600 ;
        RECT 2449.320 1953.110 2449.495 1953.600 ;
        RECT 2449.845 1953.320 2450.015 1953.600 ;
        RECT 2449.845 1953.150 2450.075 1953.320 ;
        RECT 2433.075 1952.425 2433.305 1952.625 ;
        RECT 2443.705 1952.610 2444.115 1952.940 ;
        RECT 2433.075 1952.395 2433.605 1952.425 ;
        RECT 2433.135 1952.255 2433.605 1952.395 ;
        RECT 2434.125 1952.255 2434.595 1952.425 ;
        RECT 2433.135 1951.565 2433.305 1952.255 ;
        RECT 2433.505 1951.790 2433.675 1951.885 ;
        RECT 2434.125 1951.790 2434.295 1952.255 ;
        RECT 2443.705 1952.100 2443.875 1952.610 ;
        RECT 2433.505 1951.610 2434.295 1951.790 ;
        RECT 2432.145 1950.310 2432.320 1951.450 ;
        RECT 2433.505 1950.305 2433.680 1951.610 ;
        RECT 2434.125 1951.565 2434.295 1951.610 ;
        RECT 2434.495 1951.450 2434.665 1951.885 ;
        RECT 2443.705 1951.770 2444.115 1952.100 ;
        RECT 2443.705 1951.570 2443.875 1951.770 ;
        RECT 2444.660 1951.570 2444.830 1952.520 ;
        RECT 2434.495 1950.305 2434.670 1951.450 ;
        RECT 2443.705 1950.310 2443.880 1951.570 ;
        RECT 2444.660 1950.310 2444.835 1951.570 ;
        RECT 2445.090 1951.450 2445.260 1953.050 ;
        RECT 2449.320 1952.940 2449.490 1953.110 ;
        RECT 2449.320 1952.610 2449.730 1952.940 ;
        RECT 2449.320 1952.100 2449.490 1952.610 ;
        RECT 2449.320 1951.770 2449.730 1952.100 ;
        RECT 2449.320 1951.570 2449.490 1951.770 ;
        RECT 2445.090 1950.310 2445.265 1951.450 ;
        RECT 2449.320 1950.310 2449.495 1951.570 ;
        RECT 2449.905 1951.540 2450.075 1953.150 ;
        RECT 2450.275 1953.090 2450.450 1953.600 ;
        RECT 2450.705 1953.050 2450.880 1953.600 ;
        RECT 2452.070 1953.085 2452.240 1953.595 ;
        RECT 2453.060 1953.085 2453.230 1953.595 ;
        RECT 2449.845 1951.370 2450.075 1951.540 ;
        RECT 2450.275 1951.570 2450.445 1952.520 ;
        RECT 2449.845 1950.310 2450.015 1951.370 ;
        RECT 2450.275 1950.310 2450.450 1951.570 ;
        RECT 2450.705 1951.450 2450.875 1953.050 ;
        RECT 2451.635 1952.425 2451.865 1952.625 ;
        RECT 2451.635 1952.395 2452.165 1952.425 ;
        RECT 2451.695 1952.255 2452.165 1952.395 ;
        RECT 2452.685 1952.255 2453.155 1952.425 ;
        RECT 2451.695 1951.565 2451.865 1952.255 ;
        RECT 2452.065 1951.790 2452.235 1951.885 ;
        RECT 2452.685 1951.790 2452.855 1952.255 ;
        RECT 2452.065 1951.610 2452.855 1951.790 ;
        RECT 2450.705 1950.310 2450.880 1951.450 ;
        RECT 2452.065 1950.305 2452.240 1951.610 ;
        RECT 2452.685 1951.565 2452.855 1951.610 ;
        RECT 2453.055 1951.450 2453.225 1951.885 ;
        RECT 2453.055 1950.305 2453.230 1951.450 ;
        RECT 2522.640 1950.850 2523.160 1952.335 ;
        RECT 2523.330 1951.510 2523.850 1953.060 ;
        RECT 2697.075 1951.585 2697.245 1952.345 ;
        RECT 2697.075 1951.415 2697.740 1951.585 ;
        RECT 2697.925 1951.440 2698.195 1952.345 ;
        RECT 2697.570 1951.270 2697.740 1951.415 ;
        RECT 2697.005 1950.865 2697.335 1951.235 ;
        RECT 2697.570 1950.940 2697.855 1951.270 ;
        RECT 2697.570 1950.685 2697.740 1950.940 ;
        RECT 2697.075 1950.515 2697.740 1950.685 ;
        RECT 2698.025 1950.640 2698.195 1951.440 ;
        RECT 2698.455 1951.585 2698.625 1952.345 ;
        RECT 2698.455 1951.415 2699.120 1951.585 ;
        RECT 2699.305 1951.440 2699.575 1952.345 ;
        RECT 2698.950 1951.270 2699.120 1951.415 ;
        RECT 2698.385 1950.865 2698.715 1951.235 ;
        RECT 2698.950 1950.940 2699.235 1951.270 ;
        RECT 2698.950 1950.685 2699.120 1950.940 ;
        RECT 2697.075 1950.135 2697.245 1950.515 ;
        RECT 2697.935 1950.135 2698.195 1950.640 ;
        RECT 2698.455 1950.515 2699.120 1950.685 ;
        RECT 2699.405 1950.640 2699.575 1951.440 ;
        RECT 2698.455 1950.135 2698.625 1950.515 ;
        RECT 2699.315 1950.135 2699.575 1950.640 ;
        RECT 2361.875 1947.575 2362.045 1947.935 ;
        RECT 2362.835 1947.605 2363.005 1947.765 ;
        RECT 2364.795 1947.685 2364.965 1947.795 ;
        RECT 2362.215 1947.435 2363.005 1947.605 ;
        RECT 2363.755 1947.515 2365.045 1947.685 ;
        RECT 2362.215 1947.375 2362.385 1947.435 ;
        RECT 2362.115 1947.205 2362.385 1947.375 ;
        RECT 2362.835 1947.345 2363.005 1947.435 ;
        RECT 2365.275 1947.345 2365.445 1947.765 ;
        RECT 2365.755 1947.435 2365.925 1947.795 ;
        RECT 2366.675 1947.515 2367.165 1947.685 ;
        RECT 2362.115 1947.135 2362.285 1947.205 ;
        RECT 2361.875 1946.865 2362.285 1947.135 ;
        RECT 2362.115 1946.785 2362.285 1946.865 ;
        RECT 2362.595 1946.785 2362.765 1947.115 ;
        RECT 2363.745 1946.865 2364.325 1947.035 ;
        RECT 2363.745 1946.785 2363.915 1946.865 ;
        RECT 2364.555 1946.785 2364.725 1947.235 ;
        RECT 2366.275 1947.035 2366.445 1947.515 ;
        RECT 2366.995 1947.345 2368.005 1947.515 ;
        RECT 2368.195 1947.435 2368.365 1948.075 ;
        RECT 2368.715 1947.775 2368.885 1948.105 ;
        RECT 2369.675 1947.905 2370.325 1948.075 ;
        RECT 2370.035 1947.515 2370.325 1947.905 ;
        RECT 2371.035 1947.905 2371.325 1948.075 ;
        RECT 2367.835 1947.115 2368.005 1947.345 ;
        RECT 2368.715 1947.375 2368.885 1947.515 ;
        RECT 2370.155 1947.435 2370.325 1947.515 ;
        RECT 2368.715 1947.205 2369.605 1947.375 ;
        RECT 2370.675 1947.345 2370.845 1947.765 ;
        RECT 2371.035 1947.515 2371.205 1947.905 ;
        RECT 2371.875 1947.515 2372.845 1947.685 ;
        RECT 2371.035 1947.345 2371.325 1947.515 ;
        RECT 2371.875 1947.345 2372.045 1947.515 ;
        RECT 2365.435 1946.865 2365.925 1947.035 ;
        RECT 2366.275 1946.865 2366.765 1947.035 ;
        RECT 2365.755 1946.785 2365.925 1946.865 ;
        RECT 2366.995 1946.785 2367.165 1947.115 ;
        RECT 2367.475 1946.785 2367.645 1947.115 ;
        RECT 2367.835 1946.865 2368.125 1947.115 ;
        RECT 2367.955 1946.785 2368.125 1946.865 ;
        RECT 2368.715 1946.865 2369.205 1947.035 ;
        RECT 2368.715 1946.785 2368.885 1946.865 ;
        RECT 2369.435 1946.785 2369.605 1947.205 ;
        RECT 2370.155 1947.135 2370.325 1947.235 ;
        RECT 2369.915 1947.035 2370.325 1947.135 ;
        RECT 2371.035 1947.035 2371.205 1947.345 ;
        RECT 2369.835 1946.965 2370.325 1947.035 ;
        RECT 2369.835 1946.865 2370.165 1946.965 ;
        RECT 2370.835 1946.865 2371.205 1947.035 ;
        RECT 2371.395 1947.035 2371.565 1947.115 ;
        RECT 2371.395 1946.865 2372.125 1947.035 ;
        RECT 2371.395 1946.785 2371.565 1946.865 ;
        RECT 2372.355 1946.785 2372.525 1947.235 ;
        RECT 2375.080 1946.895 2375.255 1948.155 ;
        RECT 2375.605 1947.095 2375.775 1948.155 ;
        RECT 2375.605 1946.925 2375.835 1947.095 ;
        RECT 2375.080 1946.695 2375.250 1946.895 ;
        RECT 2361.875 1946.045 2362.045 1946.395 ;
        RECT 2362.835 1946.295 2363.005 1946.395 ;
        RECT 2365.275 1946.295 2365.445 1946.395 ;
        RECT 2366.755 1946.295 2366.925 1946.395 ;
        RECT 2362.835 1946.125 2363.565 1946.295 ;
        RECT 2364.715 1946.125 2365.445 1946.295 ;
        RECT 2366.195 1946.125 2366.925 1946.295 ;
        RECT 2367.715 1946.045 2367.885 1946.395 ;
        RECT 2368.715 1946.045 2368.885 1946.395 ;
        RECT 2369.675 1946.045 2369.845 1946.395 ;
        RECT 2371.155 1946.045 2371.325 1946.395 ;
        RECT 2372.115 1946.045 2372.285 1946.395 ;
        RECT 2375.080 1946.365 2375.490 1946.695 ;
        RECT 2375.080 1945.855 2375.250 1946.365 ;
        RECT 2375.080 1945.525 2375.490 1945.855 ;
        RECT 2375.080 1945.355 2375.250 1945.525 ;
        RECT 2375.080 1944.865 2375.255 1945.355 ;
        RECT 2375.665 1945.315 2375.835 1946.925 ;
        RECT 2376.035 1946.895 2376.210 1948.155 ;
        RECT 2376.465 1947.015 2376.640 1948.155 ;
        RECT 2376.035 1945.945 2376.205 1946.895 ;
        RECT 2376.465 1945.415 2376.635 1947.015 ;
        RECT 2377.455 1946.210 2377.625 1946.900 ;
        RECT 2377.825 1946.860 2378.000 1948.160 ;
        RECT 2378.810 1947.015 2378.985 1948.160 ;
        RECT 2380.435 1947.575 2380.605 1947.935 ;
        RECT 2381.395 1947.605 2381.565 1947.765 ;
        RECT 2383.355 1947.685 2383.525 1947.795 ;
        RECT 2380.775 1947.435 2381.565 1947.605 ;
        RECT 2382.315 1947.515 2383.605 1947.685 ;
        RECT 2380.775 1947.375 2380.945 1947.435 ;
        RECT 2380.675 1947.205 2380.945 1947.375 ;
        RECT 2381.395 1947.345 2381.565 1947.435 ;
        RECT 2383.835 1947.345 2384.005 1947.765 ;
        RECT 2384.315 1947.435 2384.485 1947.795 ;
        RECT 2385.235 1947.515 2385.725 1947.685 ;
        RECT 2380.675 1947.135 2380.845 1947.205 ;
        RECT 2378.440 1946.860 2378.610 1946.900 ;
        RECT 2377.825 1946.665 2378.610 1946.860 ;
        RECT 2377.825 1946.580 2377.995 1946.665 ;
        RECT 2378.440 1946.210 2378.610 1946.665 ;
        RECT 2378.810 1946.580 2378.980 1947.015 ;
        RECT 2380.435 1946.865 2380.845 1947.135 ;
        RECT 2380.675 1946.785 2380.845 1946.865 ;
        RECT 2381.155 1946.785 2381.325 1947.115 ;
        RECT 2382.305 1946.865 2382.885 1947.035 ;
        RECT 2382.305 1946.785 2382.475 1946.865 ;
        RECT 2383.115 1946.785 2383.285 1947.235 ;
        RECT 2384.835 1947.035 2385.005 1947.515 ;
        RECT 2385.555 1947.345 2386.565 1947.515 ;
        RECT 2386.755 1947.435 2386.925 1948.075 ;
        RECT 2387.275 1947.775 2387.445 1948.105 ;
        RECT 2388.235 1947.905 2388.885 1948.075 ;
        RECT 2388.595 1947.515 2388.885 1947.905 ;
        RECT 2389.595 1947.905 2389.885 1948.075 ;
        RECT 2386.395 1947.115 2386.565 1947.345 ;
        RECT 2387.275 1947.375 2387.445 1947.515 ;
        RECT 2388.715 1947.435 2388.885 1947.515 ;
        RECT 2387.275 1947.205 2388.165 1947.375 ;
        RECT 2389.235 1947.345 2389.405 1947.765 ;
        RECT 2389.595 1947.515 2389.765 1947.905 ;
        RECT 2390.435 1947.515 2391.405 1947.685 ;
        RECT 2389.595 1947.345 2389.885 1947.515 ;
        RECT 2390.435 1947.345 2390.605 1947.515 ;
        RECT 2383.995 1946.865 2384.485 1947.035 ;
        RECT 2384.835 1946.865 2385.325 1947.035 ;
        RECT 2384.315 1946.785 2384.485 1946.865 ;
        RECT 2385.555 1946.785 2385.725 1947.115 ;
        RECT 2386.035 1946.785 2386.205 1947.115 ;
        RECT 2386.395 1946.865 2386.685 1947.115 ;
        RECT 2386.515 1946.785 2386.685 1946.865 ;
        RECT 2387.275 1946.865 2387.765 1947.035 ;
        RECT 2387.275 1946.785 2387.445 1946.865 ;
        RECT 2387.995 1946.785 2388.165 1947.205 ;
        RECT 2388.715 1947.135 2388.885 1947.235 ;
        RECT 2388.475 1947.035 2388.885 1947.135 ;
        RECT 2389.595 1947.035 2389.765 1947.345 ;
        RECT 2388.395 1946.965 2388.885 1947.035 ;
        RECT 2388.395 1946.865 2388.725 1946.965 ;
        RECT 2389.395 1946.865 2389.765 1947.035 ;
        RECT 2389.955 1947.035 2390.125 1947.115 ;
        RECT 2389.955 1946.865 2390.685 1947.035 ;
        RECT 2389.955 1946.785 2390.125 1946.865 ;
        RECT 2390.915 1946.785 2391.085 1947.235 ;
        RECT 2393.640 1946.895 2393.815 1948.155 ;
        RECT 2394.165 1947.095 2394.335 1948.155 ;
        RECT 2394.165 1946.925 2394.395 1947.095 ;
        RECT 2393.640 1946.695 2393.810 1946.895 ;
        RECT 2377.455 1946.185 2377.925 1946.210 ;
        RECT 2377.400 1946.040 2377.925 1946.185 ;
        RECT 2378.440 1946.040 2378.910 1946.210 ;
        RECT 2380.435 1946.045 2380.605 1946.395 ;
        RECT 2381.395 1946.295 2381.565 1946.395 ;
        RECT 2383.835 1946.295 2384.005 1946.395 ;
        RECT 2385.315 1946.295 2385.485 1946.395 ;
        RECT 2381.395 1946.125 2382.125 1946.295 ;
        RECT 2383.275 1946.125 2384.005 1946.295 ;
        RECT 2384.755 1946.125 2385.485 1946.295 ;
        RECT 2386.275 1946.045 2386.445 1946.395 ;
        RECT 2387.275 1946.045 2387.445 1946.395 ;
        RECT 2388.235 1946.045 2388.405 1946.395 ;
        RECT 2389.715 1946.045 2389.885 1946.395 ;
        RECT 2390.675 1946.045 2390.845 1946.395 ;
        RECT 2393.640 1946.365 2394.050 1946.695 ;
        RECT 2377.400 1945.955 2377.630 1946.040 ;
        RECT 2393.640 1945.855 2393.810 1946.365 ;
        RECT 2393.640 1945.525 2394.050 1945.855 ;
        RECT 2375.605 1945.145 2375.835 1945.315 ;
        RECT 2375.605 1944.865 2375.775 1945.145 ;
        RECT 2376.035 1944.865 2376.210 1945.375 ;
        RECT 2376.465 1944.865 2376.640 1945.415 ;
        RECT 2377.830 1944.870 2378.000 1945.380 ;
        RECT 2378.815 1944.870 2378.985 1945.380 ;
        RECT 2393.640 1945.355 2393.810 1945.525 ;
        RECT 2393.640 1944.865 2393.815 1945.355 ;
        RECT 2394.225 1945.315 2394.395 1946.925 ;
        RECT 2394.595 1946.895 2394.770 1948.155 ;
        RECT 2395.025 1947.015 2395.200 1948.155 ;
        RECT 2394.595 1945.945 2394.765 1946.895 ;
        RECT 2395.025 1945.415 2395.195 1947.015 ;
        RECT 2396.015 1946.210 2396.185 1946.900 ;
        RECT 2396.385 1946.860 2396.560 1948.160 ;
        RECT 2397.370 1947.015 2397.545 1948.160 ;
        RECT 2398.995 1947.575 2399.165 1947.935 ;
        RECT 2399.955 1947.605 2400.125 1947.765 ;
        RECT 2401.915 1947.685 2402.085 1947.795 ;
        RECT 2399.335 1947.435 2400.125 1947.605 ;
        RECT 2400.875 1947.515 2402.165 1947.685 ;
        RECT 2399.335 1947.375 2399.505 1947.435 ;
        RECT 2399.235 1947.205 2399.505 1947.375 ;
        RECT 2399.955 1947.345 2400.125 1947.435 ;
        RECT 2402.395 1947.345 2402.565 1947.765 ;
        RECT 2402.875 1947.435 2403.045 1947.795 ;
        RECT 2403.795 1947.515 2404.285 1947.685 ;
        RECT 2399.235 1947.135 2399.405 1947.205 ;
        RECT 2397.000 1946.860 2397.170 1946.900 ;
        RECT 2396.385 1946.665 2397.170 1946.860 ;
        RECT 2396.385 1946.580 2396.555 1946.665 ;
        RECT 2397.000 1946.210 2397.170 1946.665 ;
        RECT 2397.370 1946.580 2397.540 1947.015 ;
        RECT 2398.995 1946.865 2399.405 1947.135 ;
        RECT 2399.235 1946.785 2399.405 1946.865 ;
        RECT 2399.715 1946.785 2399.885 1947.115 ;
        RECT 2400.865 1946.865 2401.445 1947.035 ;
        RECT 2400.865 1946.785 2401.035 1946.865 ;
        RECT 2401.675 1946.785 2401.845 1947.235 ;
        RECT 2403.395 1947.035 2403.565 1947.515 ;
        RECT 2404.115 1947.345 2405.125 1947.515 ;
        RECT 2405.315 1947.435 2405.485 1948.075 ;
        RECT 2405.835 1947.775 2406.005 1948.105 ;
        RECT 2406.795 1947.905 2407.445 1948.075 ;
        RECT 2407.155 1947.515 2407.445 1947.905 ;
        RECT 2408.155 1947.905 2408.445 1948.075 ;
        RECT 2404.955 1947.115 2405.125 1947.345 ;
        RECT 2405.835 1947.375 2406.005 1947.515 ;
        RECT 2407.275 1947.435 2407.445 1947.515 ;
        RECT 2405.835 1947.205 2406.725 1947.375 ;
        RECT 2407.795 1947.345 2407.965 1947.765 ;
        RECT 2408.155 1947.515 2408.325 1947.905 ;
        RECT 2408.995 1947.515 2409.965 1947.685 ;
        RECT 2408.155 1947.345 2408.445 1947.515 ;
        RECT 2408.995 1947.345 2409.165 1947.515 ;
        RECT 2402.555 1946.865 2403.045 1947.035 ;
        RECT 2403.395 1946.865 2403.885 1947.035 ;
        RECT 2402.875 1946.785 2403.045 1946.865 ;
        RECT 2404.115 1946.785 2404.285 1947.115 ;
        RECT 2404.595 1946.785 2404.765 1947.115 ;
        RECT 2404.955 1946.865 2405.245 1947.115 ;
        RECT 2405.075 1946.785 2405.245 1946.865 ;
        RECT 2405.835 1946.865 2406.325 1947.035 ;
        RECT 2405.835 1946.785 2406.005 1946.865 ;
        RECT 2406.555 1946.785 2406.725 1947.205 ;
        RECT 2407.275 1947.135 2407.445 1947.235 ;
        RECT 2407.035 1947.035 2407.445 1947.135 ;
        RECT 2408.155 1947.035 2408.325 1947.345 ;
        RECT 2406.955 1946.965 2407.445 1947.035 ;
        RECT 2406.955 1946.865 2407.285 1946.965 ;
        RECT 2407.955 1946.865 2408.325 1947.035 ;
        RECT 2408.515 1947.035 2408.685 1947.115 ;
        RECT 2408.515 1946.865 2409.245 1947.035 ;
        RECT 2408.515 1946.785 2408.685 1946.865 ;
        RECT 2409.475 1946.785 2409.645 1947.235 ;
        RECT 2412.200 1946.895 2412.375 1948.155 ;
        RECT 2412.725 1947.095 2412.895 1948.155 ;
        RECT 2412.725 1946.925 2412.955 1947.095 ;
        RECT 2412.200 1946.695 2412.370 1946.895 ;
        RECT 2396.015 1946.185 2396.485 1946.210 ;
        RECT 2395.960 1946.040 2396.485 1946.185 ;
        RECT 2397.000 1946.040 2397.470 1946.210 ;
        RECT 2398.995 1946.045 2399.165 1946.395 ;
        RECT 2399.955 1946.295 2400.125 1946.395 ;
        RECT 2402.395 1946.295 2402.565 1946.395 ;
        RECT 2403.875 1946.295 2404.045 1946.395 ;
        RECT 2399.955 1946.125 2400.685 1946.295 ;
        RECT 2401.835 1946.125 2402.565 1946.295 ;
        RECT 2403.315 1946.125 2404.045 1946.295 ;
        RECT 2404.835 1946.045 2405.005 1946.395 ;
        RECT 2405.835 1946.045 2406.005 1946.395 ;
        RECT 2406.795 1946.045 2406.965 1946.395 ;
        RECT 2408.275 1946.045 2408.445 1946.395 ;
        RECT 2409.235 1946.045 2409.405 1946.395 ;
        RECT 2412.200 1946.365 2412.610 1946.695 ;
        RECT 2395.960 1945.955 2396.190 1946.040 ;
        RECT 2412.200 1945.855 2412.370 1946.365 ;
        RECT 2412.200 1945.525 2412.610 1945.855 ;
        RECT 2394.165 1945.145 2394.395 1945.315 ;
        RECT 2394.165 1944.865 2394.335 1945.145 ;
        RECT 2394.595 1944.865 2394.770 1945.375 ;
        RECT 2395.025 1944.865 2395.200 1945.415 ;
        RECT 2396.390 1944.870 2396.560 1945.380 ;
        RECT 2397.375 1944.870 2397.545 1945.380 ;
        RECT 2412.200 1945.355 2412.370 1945.525 ;
        RECT 2412.200 1944.865 2412.375 1945.355 ;
        RECT 2412.785 1945.315 2412.955 1946.925 ;
        RECT 2413.155 1946.895 2413.330 1948.155 ;
        RECT 2413.585 1947.015 2413.760 1948.155 ;
        RECT 2413.155 1945.945 2413.325 1946.895 ;
        RECT 2413.585 1945.415 2413.755 1947.015 ;
        RECT 2414.575 1946.210 2414.745 1946.900 ;
        RECT 2414.945 1946.860 2415.120 1948.160 ;
        RECT 2415.930 1947.015 2416.105 1948.160 ;
        RECT 2417.555 1947.575 2417.725 1947.935 ;
        RECT 2418.515 1947.605 2418.685 1947.765 ;
        RECT 2420.475 1947.685 2420.645 1947.795 ;
        RECT 2417.895 1947.435 2418.685 1947.605 ;
        RECT 2419.435 1947.515 2420.725 1947.685 ;
        RECT 2417.895 1947.375 2418.065 1947.435 ;
        RECT 2417.795 1947.205 2418.065 1947.375 ;
        RECT 2418.515 1947.345 2418.685 1947.435 ;
        RECT 2420.955 1947.345 2421.125 1947.765 ;
        RECT 2421.435 1947.435 2421.605 1947.795 ;
        RECT 2422.355 1947.515 2422.845 1947.685 ;
        RECT 2417.795 1947.135 2417.965 1947.205 ;
        RECT 2415.560 1946.860 2415.730 1946.900 ;
        RECT 2414.945 1946.665 2415.730 1946.860 ;
        RECT 2414.945 1946.580 2415.115 1946.665 ;
        RECT 2415.560 1946.210 2415.730 1946.665 ;
        RECT 2415.930 1946.580 2416.100 1947.015 ;
        RECT 2417.555 1946.865 2417.965 1947.135 ;
        RECT 2417.795 1946.785 2417.965 1946.865 ;
        RECT 2418.275 1946.785 2418.445 1947.115 ;
        RECT 2419.425 1946.865 2420.005 1947.035 ;
        RECT 2419.425 1946.785 2419.595 1946.865 ;
        RECT 2420.235 1946.785 2420.405 1947.235 ;
        RECT 2421.955 1947.035 2422.125 1947.515 ;
        RECT 2422.675 1947.345 2423.685 1947.515 ;
        RECT 2423.875 1947.435 2424.045 1948.075 ;
        RECT 2424.395 1947.775 2424.565 1948.105 ;
        RECT 2425.355 1947.905 2426.005 1948.075 ;
        RECT 2425.715 1947.515 2426.005 1947.905 ;
        RECT 2426.715 1947.905 2427.005 1948.075 ;
        RECT 2423.515 1947.115 2423.685 1947.345 ;
        RECT 2424.395 1947.375 2424.565 1947.515 ;
        RECT 2425.835 1947.435 2426.005 1947.515 ;
        RECT 2424.395 1947.205 2425.285 1947.375 ;
        RECT 2426.355 1947.345 2426.525 1947.765 ;
        RECT 2426.715 1947.515 2426.885 1947.905 ;
        RECT 2427.555 1947.515 2428.525 1947.685 ;
        RECT 2426.715 1947.345 2427.005 1947.515 ;
        RECT 2427.555 1947.345 2427.725 1947.515 ;
        RECT 2421.115 1946.865 2421.605 1947.035 ;
        RECT 2421.955 1946.865 2422.445 1947.035 ;
        RECT 2421.435 1946.785 2421.605 1946.865 ;
        RECT 2422.675 1946.785 2422.845 1947.115 ;
        RECT 2423.155 1946.785 2423.325 1947.115 ;
        RECT 2423.515 1946.865 2423.805 1947.115 ;
        RECT 2423.635 1946.785 2423.805 1946.865 ;
        RECT 2424.395 1946.865 2424.885 1947.035 ;
        RECT 2424.395 1946.785 2424.565 1946.865 ;
        RECT 2425.115 1946.785 2425.285 1947.205 ;
        RECT 2425.835 1947.135 2426.005 1947.235 ;
        RECT 2425.595 1947.035 2426.005 1947.135 ;
        RECT 2426.715 1947.035 2426.885 1947.345 ;
        RECT 2425.515 1946.965 2426.005 1947.035 ;
        RECT 2425.515 1946.865 2425.845 1946.965 ;
        RECT 2426.515 1946.865 2426.885 1947.035 ;
        RECT 2427.075 1947.035 2427.245 1947.115 ;
        RECT 2427.075 1946.865 2427.805 1947.035 ;
        RECT 2427.075 1946.785 2427.245 1946.865 ;
        RECT 2428.035 1946.785 2428.205 1947.235 ;
        RECT 2430.760 1946.895 2430.935 1948.155 ;
        RECT 2431.285 1947.095 2431.455 1948.155 ;
        RECT 2431.285 1946.925 2431.515 1947.095 ;
        RECT 2430.760 1946.695 2430.930 1946.895 ;
        RECT 2414.575 1946.185 2415.045 1946.210 ;
        RECT 2414.520 1946.040 2415.045 1946.185 ;
        RECT 2415.560 1946.040 2416.030 1946.210 ;
        RECT 2417.555 1946.045 2417.725 1946.395 ;
        RECT 2418.515 1946.295 2418.685 1946.395 ;
        RECT 2420.955 1946.295 2421.125 1946.395 ;
        RECT 2422.435 1946.295 2422.605 1946.395 ;
        RECT 2418.515 1946.125 2419.245 1946.295 ;
        RECT 2420.395 1946.125 2421.125 1946.295 ;
        RECT 2421.875 1946.125 2422.605 1946.295 ;
        RECT 2423.395 1946.045 2423.565 1946.395 ;
        RECT 2424.395 1946.045 2424.565 1946.395 ;
        RECT 2425.355 1946.045 2425.525 1946.395 ;
        RECT 2426.835 1946.045 2427.005 1946.395 ;
        RECT 2427.795 1946.045 2427.965 1946.395 ;
        RECT 2430.760 1946.365 2431.170 1946.695 ;
        RECT 2414.520 1945.955 2414.750 1946.040 ;
        RECT 2430.760 1945.855 2430.930 1946.365 ;
        RECT 2430.760 1945.525 2431.170 1945.855 ;
        RECT 2412.725 1945.145 2412.955 1945.315 ;
        RECT 2412.725 1944.865 2412.895 1945.145 ;
        RECT 2413.155 1944.865 2413.330 1945.375 ;
        RECT 2413.585 1944.865 2413.760 1945.415 ;
        RECT 2414.950 1944.870 2415.120 1945.380 ;
        RECT 2415.935 1944.870 2416.105 1945.380 ;
        RECT 2430.760 1945.355 2430.930 1945.525 ;
        RECT 2430.760 1944.865 2430.935 1945.355 ;
        RECT 2431.345 1945.315 2431.515 1946.925 ;
        RECT 2431.715 1946.895 2431.890 1948.155 ;
        RECT 2432.145 1947.015 2432.320 1948.155 ;
        RECT 2431.715 1945.945 2431.885 1946.895 ;
        RECT 2432.145 1945.415 2432.315 1947.015 ;
        RECT 2433.135 1946.210 2433.305 1946.900 ;
        RECT 2433.505 1946.860 2433.680 1948.160 ;
        RECT 2434.490 1947.015 2434.665 1948.160 ;
        RECT 2436.115 1947.575 2436.285 1947.935 ;
        RECT 2437.075 1947.605 2437.245 1947.765 ;
        RECT 2439.035 1947.685 2439.205 1947.795 ;
        RECT 2436.455 1947.435 2437.245 1947.605 ;
        RECT 2437.995 1947.515 2439.285 1947.685 ;
        RECT 2436.455 1947.375 2436.625 1947.435 ;
        RECT 2436.355 1947.205 2436.625 1947.375 ;
        RECT 2437.075 1947.345 2437.245 1947.435 ;
        RECT 2439.515 1947.345 2439.685 1947.765 ;
        RECT 2439.995 1947.435 2440.165 1947.795 ;
        RECT 2440.915 1947.515 2441.405 1947.685 ;
        RECT 2436.355 1947.135 2436.525 1947.205 ;
        RECT 2434.120 1946.860 2434.290 1946.900 ;
        RECT 2433.505 1946.665 2434.290 1946.860 ;
        RECT 2433.505 1946.580 2433.675 1946.665 ;
        RECT 2434.120 1946.210 2434.290 1946.665 ;
        RECT 2434.490 1946.580 2434.660 1947.015 ;
        RECT 2436.115 1946.865 2436.525 1947.135 ;
        RECT 2436.355 1946.785 2436.525 1946.865 ;
        RECT 2436.835 1946.785 2437.005 1947.115 ;
        RECT 2437.985 1946.865 2438.565 1947.035 ;
        RECT 2437.985 1946.785 2438.155 1946.865 ;
        RECT 2438.795 1946.785 2438.965 1947.235 ;
        RECT 2440.515 1947.035 2440.685 1947.515 ;
        RECT 2441.235 1947.345 2442.245 1947.515 ;
        RECT 2442.435 1947.435 2442.605 1948.075 ;
        RECT 2442.955 1947.775 2443.125 1948.105 ;
        RECT 2443.915 1947.905 2444.565 1948.075 ;
        RECT 2444.275 1947.515 2444.565 1947.905 ;
        RECT 2445.275 1947.905 2445.565 1948.075 ;
        RECT 2442.075 1947.115 2442.245 1947.345 ;
        RECT 2442.955 1947.375 2443.125 1947.515 ;
        RECT 2444.395 1947.435 2444.565 1947.515 ;
        RECT 2442.955 1947.205 2443.845 1947.375 ;
        RECT 2444.915 1947.345 2445.085 1947.765 ;
        RECT 2445.275 1947.515 2445.445 1947.905 ;
        RECT 2446.115 1947.515 2447.085 1947.685 ;
        RECT 2445.275 1947.345 2445.565 1947.515 ;
        RECT 2446.115 1947.345 2446.285 1947.515 ;
        RECT 2439.675 1946.865 2440.165 1947.035 ;
        RECT 2440.515 1946.865 2441.005 1947.035 ;
        RECT 2439.995 1946.785 2440.165 1946.865 ;
        RECT 2441.235 1946.785 2441.405 1947.115 ;
        RECT 2441.715 1946.785 2441.885 1947.115 ;
        RECT 2442.075 1946.865 2442.365 1947.115 ;
        RECT 2442.195 1946.785 2442.365 1946.865 ;
        RECT 2442.955 1946.865 2443.445 1947.035 ;
        RECT 2442.955 1946.785 2443.125 1946.865 ;
        RECT 2443.675 1946.785 2443.845 1947.205 ;
        RECT 2444.395 1947.135 2444.565 1947.235 ;
        RECT 2444.155 1947.035 2444.565 1947.135 ;
        RECT 2445.275 1947.035 2445.445 1947.345 ;
        RECT 2444.075 1946.965 2444.565 1947.035 ;
        RECT 2444.075 1946.865 2444.405 1946.965 ;
        RECT 2445.075 1946.865 2445.445 1947.035 ;
        RECT 2445.635 1947.035 2445.805 1947.115 ;
        RECT 2445.635 1946.865 2446.365 1947.035 ;
        RECT 2445.635 1946.785 2445.805 1946.865 ;
        RECT 2446.595 1946.785 2446.765 1947.235 ;
        RECT 2449.320 1946.895 2449.495 1948.155 ;
        RECT 2449.845 1947.095 2450.015 1948.155 ;
        RECT 2449.845 1946.925 2450.075 1947.095 ;
        RECT 2449.320 1946.695 2449.490 1946.895 ;
        RECT 2433.135 1946.185 2433.605 1946.210 ;
        RECT 2433.080 1946.040 2433.605 1946.185 ;
        RECT 2434.120 1946.040 2434.590 1946.210 ;
        RECT 2436.115 1946.045 2436.285 1946.395 ;
        RECT 2437.075 1946.295 2437.245 1946.395 ;
        RECT 2439.515 1946.295 2439.685 1946.395 ;
        RECT 2440.995 1946.295 2441.165 1946.395 ;
        RECT 2437.075 1946.125 2437.805 1946.295 ;
        RECT 2438.955 1946.125 2439.685 1946.295 ;
        RECT 2440.435 1946.125 2441.165 1946.295 ;
        RECT 2441.955 1946.045 2442.125 1946.395 ;
        RECT 2442.955 1946.045 2443.125 1946.395 ;
        RECT 2443.915 1946.045 2444.085 1946.395 ;
        RECT 2445.395 1946.045 2445.565 1946.395 ;
        RECT 2446.355 1946.045 2446.525 1946.395 ;
        RECT 2449.320 1946.365 2449.730 1946.695 ;
        RECT 2433.080 1945.955 2433.310 1946.040 ;
        RECT 2449.320 1945.855 2449.490 1946.365 ;
        RECT 2449.320 1945.525 2449.730 1945.855 ;
        RECT 2431.285 1945.145 2431.515 1945.315 ;
        RECT 2431.285 1944.865 2431.455 1945.145 ;
        RECT 2431.715 1944.865 2431.890 1945.375 ;
        RECT 2432.145 1944.865 2432.320 1945.415 ;
        RECT 2433.510 1944.870 2433.680 1945.380 ;
        RECT 2434.495 1944.870 2434.665 1945.380 ;
        RECT 2449.320 1945.355 2449.490 1945.525 ;
        RECT 2449.320 1944.865 2449.495 1945.355 ;
        RECT 2449.905 1945.315 2450.075 1946.925 ;
        RECT 2450.275 1946.895 2450.450 1948.155 ;
        RECT 2450.705 1947.015 2450.880 1948.155 ;
        RECT 2450.275 1945.945 2450.445 1946.895 ;
        RECT 2450.705 1945.415 2450.875 1947.015 ;
        RECT 2451.695 1946.210 2451.865 1946.900 ;
        RECT 2452.065 1946.860 2452.240 1948.160 ;
        RECT 2453.050 1947.015 2453.225 1948.160 ;
        RECT 2452.680 1946.860 2452.850 1946.900 ;
        RECT 2452.065 1946.665 2452.850 1946.860 ;
        RECT 2452.065 1946.580 2452.235 1946.665 ;
        RECT 2452.680 1946.210 2452.850 1946.665 ;
        RECT 2453.050 1946.580 2453.220 1947.015 ;
        RECT 2451.695 1946.185 2452.165 1946.210 ;
        RECT 2451.640 1946.040 2452.165 1946.185 ;
        RECT 2452.680 1946.040 2453.150 1946.210 ;
        RECT 2451.640 1945.955 2451.870 1946.040 ;
        RECT 2449.845 1945.145 2450.075 1945.315 ;
        RECT 2449.845 1944.865 2450.015 1945.145 ;
        RECT 2450.275 1944.865 2450.450 1945.375 ;
        RECT 2450.705 1944.865 2450.880 1945.415 ;
        RECT 2452.070 1944.870 2452.240 1945.380 ;
        RECT 2453.055 1944.870 2453.225 1945.380 ;
        RECT 2882.085 1892.500 2882.605 1894.050 ;
        RECT 2696.985 1856.335 2697.245 1856.665 ;
        RECT 2696.985 1855.425 2697.155 1856.335 ;
        RECT 2697.940 1856.265 2698.145 1856.665 ;
        RECT 2697.940 1856.095 2698.625 1856.265 ;
        RECT 2697.865 1855.425 2698.115 1855.925 ;
        RECT 2696.985 1855.255 2698.115 1855.425 ;
        RECT 2696.985 1854.485 2697.255 1855.255 ;
        RECT 2698.285 1855.065 2698.625 1856.095 ;
        RECT 2697.960 1854.890 2698.625 1855.065 ;
        RECT 2698.825 1856.160 2699.085 1856.665 ;
        RECT 2699.775 1856.285 2699.945 1856.665 ;
        RECT 2698.825 1855.360 2698.995 1856.160 ;
        RECT 2699.280 1856.115 2699.945 1856.285 ;
        RECT 2700.205 1856.160 2700.465 1856.665 ;
        RECT 2701.155 1856.285 2701.325 1856.665 ;
        RECT 2699.280 1855.860 2699.450 1856.115 ;
        RECT 2699.165 1855.530 2699.450 1855.860 ;
        RECT 2699.685 1855.565 2700.015 1855.935 ;
        RECT 2699.280 1855.385 2699.450 1855.530 ;
        RECT 2697.960 1854.485 2698.145 1854.890 ;
        RECT 2698.825 1854.455 2699.095 1855.360 ;
        RECT 2699.280 1855.215 2699.945 1855.385 ;
        RECT 2699.775 1854.455 2699.945 1855.215 ;
        RECT 2700.205 1855.360 2700.375 1856.160 ;
        RECT 2700.660 1856.115 2701.325 1856.285 ;
        RECT 2709.035 1856.285 2709.205 1856.665 ;
        RECT 2709.035 1856.115 2709.750 1856.285 ;
        RECT 2700.660 1855.860 2700.830 1856.115 ;
        RECT 2700.545 1855.530 2700.830 1855.860 ;
        RECT 2701.065 1855.565 2701.395 1855.935 ;
        RECT 2709.580 1855.925 2709.750 1856.115 ;
        RECT 2709.920 1856.090 2710.175 1856.665 ;
        RECT 2722.335 1856.265 2722.540 1856.665 ;
        RECT 2723.235 1856.335 2723.495 1856.665 ;
        RECT 2709.580 1855.595 2709.835 1855.925 ;
        RECT 2700.660 1855.385 2700.830 1855.530 ;
        RECT 2709.580 1855.385 2709.750 1855.595 ;
        RECT 2700.205 1854.455 2700.475 1855.360 ;
        RECT 2700.660 1855.215 2701.325 1855.385 ;
        RECT 2701.155 1854.455 2701.325 1855.215 ;
        RECT 2709.035 1855.215 2709.750 1855.385 ;
        RECT 2710.005 1855.360 2710.175 1856.090 ;
        RECT 2709.035 1854.455 2709.205 1855.215 ;
        RECT 2709.920 1854.455 2710.175 1855.360 ;
        RECT 2721.855 1856.095 2722.540 1856.265 ;
        RECT 2721.855 1855.065 2722.195 1856.095 ;
        RECT 2722.365 1855.425 2722.615 1855.925 ;
        RECT 2723.325 1855.425 2723.495 1856.335 ;
        RECT 2722.365 1855.255 2723.495 1855.425 ;
        RECT 2721.855 1854.890 2722.520 1855.065 ;
        RECT 2722.335 1854.485 2722.520 1854.890 ;
        RECT 2723.225 1854.485 2723.495 1855.255 ;
        RECT 2731.485 1856.160 2731.745 1856.665 ;
        RECT 2732.435 1856.285 2732.605 1856.665 ;
        RECT 2731.485 1855.360 2731.665 1856.160 ;
        RECT 2731.940 1856.115 2732.605 1856.285 ;
        RECT 2731.940 1855.860 2732.110 1856.115 ;
        RECT 2731.835 1855.530 2732.110 1855.860 ;
        RECT 2731.940 1855.385 2732.110 1855.530 ;
        RECT 2731.485 1854.455 2731.755 1855.360 ;
        RECT 2731.940 1855.215 2732.615 1855.385 ;
        RECT 2732.435 1854.455 2732.615 1855.215 ;
        RECT 2697.075 1853.185 2697.245 1853.945 ;
        RECT 2697.075 1853.015 2697.740 1853.185 ;
        RECT 2697.925 1853.040 2698.195 1853.945 ;
        RECT 2697.570 1852.870 2697.740 1853.015 ;
        RECT 2697.005 1852.465 2697.335 1852.835 ;
        RECT 2697.570 1852.540 2697.855 1852.870 ;
        RECT 2697.570 1852.285 2697.740 1852.540 ;
        RECT 2697.075 1852.115 2697.740 1852.285 ;
        RECT 2698.025 1852.240 2698.195 1853.040 ;
        RECT 2697.075 1851.735 2697.245 1852.115 ;
        RECT 2697.935 1851.735 2698.195 1852.240 ;
        RECT 2697.075 1845.405 2697.245 1845.785 ;
        RECT 2697.075 1845.235 2697.740 1845.405 ;
        RECT 2697.935 1845.280 2698.195 1845.785 ;
        RECT 2697.005 1844.685 2697.335 1845.055 ;
        RECT 2697.570 1844.980 2697.740 1845.235 ;
        RECT 2697.570 1844.650 2697.855 1844.980 ;
        RECT 2697.570 1844.505 2697.740 1844.650 ;
        RECT 2697.075 1844.335 2697.740 1844.505 ;
        RECT 2698.025 1844.480 2698.195 1845.280 ;
        RECT 2697.075 1843.575 2697.245 1844.335 ;
        RECT 2697.925 1843.575 2698.195 1844.480 ;
        RECT 2697.075 1839.965 2697.245 1840.340 ;
        RECT 2697.915 1840.175 2698.990 1840.345 ;
        RECT 2697.915 1839.965 2698.085 1840.175 ;
        RECT 2697.075 1839.795 2698.085 1839.965 ;
        RECT 2698.310 1839.835 2698.650 1840.005 ;
        RECT 2698.820 1839.840 2698.990 1840.175 ;
        RECT 2700.280 1840.175 2701.880 1840.345 ;
        RECT 2698.310 1839.665 2698.600 1839.835 ;
        RECT 2697.050 1839.495 2697.395 1839.605 ;
        RECT 2697.045 1839.325 2697.395 1839.495 ;
        RECT 2697.050 1838.985 2697.395 1839.325 ;
        RECT 2697.705 1838.985 2698.140 1839.605 ;
        RECT 2698.310 1839.145 2698.480 1839.665 ;
        RECT 2699.160 1839.495 2699.520 1840.170 ;
        RECT 2700.280 1839.805 2700.450 1840.175 ;
        RECT 2701.525 1840.135 2701.880 1840.175 ;
        RECT 2700.620 1839.755 2700.950 1840.005 ;
        RECT 2700.635 1839.680 2700.950 1839.755 ;
        RECT 2701.120 1839.885 2701.290 1840.005 ;
        RECT 2702.395 1839.885 2702.640 1840.305 ;
        RECT 2703.410 1839.945 2703.585 1840.275 ;
        RECT 2703.930 1840.185 2704.100 1840.345 ;
        RECT 2703.930 1840.015 2704.460 1840.185 ;
        RECT 2704.630 1840.175 2705.625 1840.345 ;
        RECT 2704.630 1840.015 2704.800 1840.175 ;
        RECT 2701.120 1839.715 2702.640 1839.885 ;
        RECT 2698.980 1839.315 2699.520 1839.495 ;
        RECT 2699.160 1839.205 2699.520 1839.315 ;
        RECT 2698.310 1838.975 2698.945 1839.145 ;
        RECT 2699.160 1838.975 2699.965 1839.205 ;
        RECT 2697.075 1838.635 2698.605 1838.805 ;
        RECT 2697.075 1838.135 2697.245 1838.635 ;
        RECT 2698.435 1838.475 2698.605 1838.635 ;
        RECT 2698.775 1838.645 2698.945 1838.975 ;
        RECT 2698.775 1838.475 2699.105 1838.645 ;
        RECT 2697.915 1838.305 2698.085 1838.465 ;
        RECT 2699.275 1838.305 2699.445 1838.805 ;
        RECT 2697.915 1838.135 2699.445 1838.305 ;
        RECT 2699.615 1838.135 2699.965 1838.975 ;
        RECT 2700.165 1838.605 2700.465 1839.605 ;
        RECT 2700.635 1839.155 2700.805 1839.680 ;
        RECT 2701.120 1839.675 2701.290 1839.715 ;
        RECT 2700.975 1839.495 2701.305 1839.505 ;
        RECT 2700.975 1839.335 2701.360 1839.495 ;
        RECT 2701.190 1839.325 2701.360 1839.335 ;
        RECT 2701.700 1839.155 2701.945 1839.545 ;
        RECT 2700.635 1838.985 2701.395 1839.155 ;
        RECT 2701.645 1838.985 2701.945 1839.155 ;
        RECT 2700.725 1838.305 2700.895 1838.815 ;
        RECT 2701.065 1838.475 2701.395 1838.985 ;
        RECT 2701.700 1838.925 2701.945 1838.985 ;
        RECT 2702.150 1838.925 2702.480 1839.545 ;
        RECT 2702.955 1838.925 2703.245 1839.605 ;
        RECT 2703.415 1839.495 2703.585 1839.945 ;
        RECT 2703.880 1839.665 2704.120 1839.835 ;
        RECT 2703.415 1839.325 2703.705 1839.495 ;
        RECT 2701.565 1838.515 2702.630 1838.685 ;
        RECT 2701.565 1838.305 2701.735 1838.515 ;
        RECT 2700.725 1838.135 2701.735 1838.305 ;
        RECT 2702.460 1838.135 2702.630 1838.515 ;
        RECT 2703.415 1838.465 2703.585 1839.325 ;
        RECT 2703.400 1838.135 2703.585 1838.465 ;
        RECT 2703.880 1838.465 2704.050 1839.665 ;
        RECT 2704.290 1838.845 2704.460 1840.015 ;
        RECT 2705.110 1839.835 2705.285 1840.005 ;
        RECT 2704.870 1839.675 2705.285 1839.835 ;
        RECT 2705.455 1839.885 2705.625 1840.175 ;
        RECT 2705.455 1839.715 2706.025 1839.885 ;
        RECT 2704.870 1839.665 2705.280 1839.675 ;
        RECT 2705.090 1839.325 2705.545 1839.495 ;
        RECT 2705.855 1838.935 2706.025 1839.715 ;
        RECT 2704.290 1838.615 2705.075 1838.845 ;
        RECT 2704.745 1838.475 2705.075 1838.615 ;
        RECT 2705.375 1838.765 2706.025 1838.935 ;
        RECT 2703.880 1838.135 2704.090 1838.465 ;
        RECT 2704.260 1838.305 2704.590 1838.345 ;
        RECT 2705.375 1838.305 2705.545 1838.765 ;
        RECT 2704.260 1838.135 2705.545 1838.305 ;
        RECT 2706.215 1838.135 2706.475 1840.345 ;
        RECT 2697.075 1836.865 2697.245 1837.625 ;
        RECT 2697.075 1836.695 2697.740 1836.865 ;
        RECT 2697.925 1836.720 2698.195 1837.625 ;
        RECT 2697.570 1836.550 2697.740 1836.695 ;
        RECT 2697.005 1836.145 2697.335 1836.515 ;
        RECT 2697.570 1836.220 2697.855 1836.550 ;
        RECT 2697.570 1835.965 2697.740 1836.220 ;
        RECT 2697.075 1835.795 2697.740 1835.965 ;
        RECT 2698.025 1835.920 2698.195 1836.720 ;
        RECT 2697.075 1835.415 2697.245 1835.795 ;
        RECT 2697.935 1835.415 2698.195 1835.920 ;
        RECT 2697.075 1834.525 2697.245 1834.900 ;
        RECT 2697.915 1834.735 2698.990 1834.905 ;
        RECT 2697.915 1834.525 2698.085 1834.735 ;
        RECT 2697.075 1834.355 2698.085 1834.525 ;
        RECT 2698.310 1834.395 2698.650 1834.565 ;
        RECT 2698.820 1834.400 2698.990 1834.735 ;
        RECT 2700.280 1834.735 2701.880 1834.905 ;
        RECT 2698.310 1834.225 2698.600 1834.395 ;
        RECT 2697.050 1834.055 2697.395 1834.165 ;
        RECT 2697.045 1833.885 2697.395 1834.055 ;
        RECT 2697.050 1833.545 2697.395 1833.885 ;
        RECT 2697.705 1833.545 2698.140 1834.165 ;
        RECT 2698.310 1833.705 2698.480 1834.225 ;
        RECT 2699.160 1834.055 2699.520 1834.730 ;
        RECT 2700.280 1834.365 2700.450 1834.735 ;
        RECT 2701.525 1834.695 2701.880 1834.735 ;
        RECT 2700.620 1834.315 2700.950 1834.565 ;
        RECT 2700.635 1834.240 2700.950 1834.315 ;
        RECT 2701.120 1834.445 2701.290 1834.565 ;
        RECT 2702.395 1834.445 2702.640 1834.865 ;
        RECT 2703.410 1834.505 2703.585 1834.835 ;
        RECT 2703.930 1834.745 2704.100 1834.905 ;
        RECT 2703.930 1834.575 2704.460 1834.745 ;
        RECT 2704.630 1834.735 2705.625 1834.905 ;
        RECT 2704.630 1834.575 2704.800 1834.735 ;
        RECT 2701.120 1834.275 2702.640 1834.445 ;
        RECT 2698.980 1833.875 2699.520 1834.055 ;
        RECT 2699.160 1833.765 2699.520 1833.875 ;
        RECT 2698.310 1833.535 2698.945 1833.705 ;
        RECT 2699.160 1833.535 2699.965 1833.765 ;
        RECT 2697.075 1833.195 2698.605 1833.365 ;
        RECT 2697.075 1832.695 2697.245 1833.195 ;
        RECT 2698.435 1833.035 2698.605 1833.195 ;
        RECT 2698.775 1833.205 2698.945 1833.535 ;
        RECT 2698.775 1833.035 2699.105 1833.205 ;
        RECT 2697.915 1832.865 2698.085 1833.025 ;
        RECT 2699.275 1832.865 2699.445 1833.365 ;
        RECT 2697.915 1832.695 2699.445 1832.865 ;
        RECT 2699.615 1832.695 2699.965 1833.535 ;
        RECT 2700.165 1833.165 2700.465 1834.165 ;
        RECT 2700.635 1833.715 2700.805 1834.240 ;
        RECT 2701.120 1834.235 2701.290 1834.275 ;
        RECT 2700.975 1834.055 2701.305 1834.065 ;
        RECT 2700.975 1833.895 2701.360 1834.055 ;
        RECT 2701.190 1833.885 2701.360 1833.895 ;
        RECT 2701.700 1833.715 2701.945 1834.105 ;
        RECT 2700.635 1833.545 2701.395 1833.715 ;
        RECT 2701.645 1833.545 2701.945 1833.715 ;
        RECT 2700.725 1832.865 2700.895 1833.375 ;
        RECT 2701.065 1833.035 2701.395 1833.545 ;
        RECT 2701.700 1833.485 2701.945 1833.545 ;
        RECT 2702.150 1833.485 2702.480 1834.105 ;
        RECT 2702.955 1833.485 2703.245 1834.165 ;
        RECT 2703.415 1834.055 2703.585 1834.505 ;
        RECT 2703.880 1834.225 2704.120 1834.395 ;
        RECT 2703.415 1833.885 2703.705 1834.055 ;
        RECT 2701.565 1833.075 2702.630 1833.245 ;
        RECT 2701.565 1832.865 2701.735 1833.075 ;
        RECT 2700.725 1832.695 2701.735 1832.865 ;
        RECT 2702.460 1832.695 2702.630 1833.075 ;
        RECT 2703.415 1833.025 2703.585 1833.885 ;
        RECT 2703.400 1832.695 2703.585 1833.025 ;
        RECT 2703.880 1833.025 2704.050 1834.225 ;
        RECT 2704.290 1833.405 2704.460 1834.575 ;
        RECT 2705.110 1834.395 2705.285 1834.565 ;
        RECT 2704.870 1834.235 2705.285 1834.395 ;
        RECT 2705.455 1834.445 2705.625 1834.735 ;
        RECT 2705.455 1834.275 2706.025 1834.445 ;
        RECT 2704.870 1834.225 2705.280 1834.235 ;
        RECT 2705.090 1833.885 2705.545 1834.055 ;
        RECT 2705.855 1833.495 2706.025 1834.275 ;
        RECT 2704.290 1833.175 2705.075 1833.405 ;
        RECT 2704.745 1833.035 2705.075 1833.175 ;
        RECT 2705.375 1833.325 2706.025 1833.495 ;
        RECT 2703.880 1832.695 2704.090 1833.025 ;
        RECT 2704.260 1832.865 2704.590 1832.905 ;
        RECT 2705.375 1832.865 2705.545 1833.325 ;
        RECT 2704.260 1832.695 2705.545 1832.865 ;
        RECT 2706.215 1832.695 2706.475 1834.905 ;
        RECT 2697.075 1831.425 2697.245 1832.185 ;
        RECT 2697.075 1831.255 2697.740 1831.425 ;
        RECT 2697.925 1831.280 2698.195 1832.185 ;
        RECT 2697.570 1831.110 2697.740 1831.255 ;
        RECT 2697.005 1830.705 2697.335 1831.075 ;
        RECT 2697.570 1830.780 2697.855 1831.110 ;
        RECT 2697.570 1830.525 2697.740 1830.780 ;
        RECT 2697.075 1830.355 2697.740 1830.525 ;
        RECT 2698.025 1830.480 2698.195 1831.280 ;
        RECT 2697.075 1829.975 2697.245 1830.355 ;
        RECT 2697.935 1829.975 2698.195 1830.480 ;
        RECT 2701.590 1831.215 2701.925 1832.185 ;
        RECT 2702.435 1832.015 2704.465 1832.185 ;
        RECT 2701.590 1830.545 2701.760 1831.215 ;
        RECT 2702.435 1831.045 2702.605 1832.015 ;
        RECT 2701.930 1830.715 2702.185 1831.045 ;
        RECT 2702.410 1830.715 2702.605 1831.045 ;
        RECT 2702.775 1831.675 2703.900 1831.845 ;
        RECT 2702.015 1830.545 2702.185 1830.715 ;
        RECT 2702.775 1830.545 2702.945 1831.675 ;
        RECT 2701.590 1829.975 2701.845 1830.545 ;
        RECT 2702.015 1830.375 2702.945 1830.545 ;
        RECT 2703.115 1831.335 2704.125 1831.505 ;
        RECT 2703.115 1830.535 2703.285 1831.335 ;
        RECT 2703.490 1830.655 2703.765 1831.135 ;
        RECT 2703.485 1830.485 2703.765 1830.655 ;
        RECT 2702.770 1830.340 2702.945 1830.375 ;
        RECT 2702.770 1829.975 2703.300 1830.340 ;
        RECT 2703.490 1829.975 2703.765 1830.485 ;
        RECT 2703.935 1829.975 2704.125 1831.335 ;
        RECT 2704.295 1831.350 2704.465 1832.015 ;
        RECT 2705.040 1831.595 2705.555 1832.005 ;
        RECT 2704.295 1831.160 2705.045 1831.350 ;
        RECT 2705.215 1830.785 2705.555 1831.595 ;
        RECT 2704.325 1830.615 2705.555 1830.785 ;
        RECT 2705.035 1830.010 2705.280 1830.615 ;
        RECT 2697.075 1825.985 2697.245 1826.745 ;
        RECT 2697.075 1825.815 2697.740 1825.985 ;
        RECT 2697.925 1825.840 2698.195 1826.745 ;
        RECT 2697.570 1825.670 2697.740 1825.815 ;
        RECT 2697.005 1825.265 2697.335 1825.635 ;
        RECT 2697.570 1825.340 2697.855 1825.670 ;
        RECT 2697.570 1825.085 2697.740 1825.340 ;
        RECT 2697.075 1824.915 2697.740 1825.085 ;
        RECT 2698.025 1825.040 2698.195 1825.840 ;
        RECT 2697.075 1824.535 2697.245 1824.915 ;
        RECT 2697.935 1824.535 2698.195 1825.040 ;
        RECT 2701.595 1820.505 2701.925 1821.290 ;
        RECT 2701.595 1820.335 2702.275 1820.505 ;
        RECT 2701.585 1819.915 2701.935 1820.165 ;
        RECT 2702.105 1819.735 2702.275 1820.335 ;
        RECT 2702.445 1819.915 2702.795 1820.165 ;
        RECT 2702.015 1819.095 2702.345 1819.735 ;
        RECT 2697.075 1818.205 2697.245 1818.585 ;
        RECT 2697.075 1818.035 2697.740 1818.205 ;
        RECT 2697.935 1818.080 2698.195 1818.585 ;
        RECT 2697.005 1817.485 2697.335 1817.855 ;
        RECT 2697.570 1817.780 2697.740 1818.035 ;
        RECT 2697.570 1817.450 2697.855 1817.780 ;
        RECT 2697.570 1817.305 2697.740 1817.450 ;
        RECT 2697.075 1817.135 2697.740 1817.305 ;
        RECT 2698.025 1817.280 2698.195 1818.080 ;
        RECT 2702.565 1818.225 2702.885 1818.585 ;
        RECT 2703.880 1818.225 2704.225 1818.585 ;
        RECT 2702.565 1818.055 2704.225 1818.225 ;
        RECT 2697.075 1816.375 2697.245 1817.135 ;
        RECT 2697.925 1816.375 2698.195 1817.280 ;
        RECT 2702.105 1817.215 2702.380 1817.845 ;
        RECT 2702.090 1816.555 2702.395 1817.045 ;
        RECT 2702.565 1816.725 2702.865 1818.055 ;
        RECT 2703.245 1817.595 2703.575 1817.765 ;
        RECT 2703.250 1817.345 2703.575 1817.595 ;
        RECT 2703.755 1817.515 2704.365 1817.845 ;
        RECT 2704.535 1817.345 2705.035 1817.805 ;
        RECT 2703.250 1817.165 2705.035 1817.345 ;
        RECT 2703.035 1816.815 2705.070 1816.985 ;
        RECT 2703.035 1816.555 2703.365 1816.815 ;
        RECT 2702.090 1816.375 2703.365 1816.555 ;
        RECT 2703.960 1816.735 2705.070 1816.815 ;
        RECT 2703.960 1816.375 2704.130 1816.735 ;
        RECT 2704.810 1816.375 2705.070 1816.735 ;
        RECT 2725.935 1815.015 2726.265 1815.865 ;
        RECT 2726.775 1815.015 2727.105 1815.865 ;
        RECT 2725.935 1814.845 2727.435 1815.015 ;
        RECT 2725.555 1814.475 2727.080 1814.675 ;
        RECT 2727.260 1814.645 2727.435 1814.845 ;
        RECT 2727.260 1814.475 2729.885 1814.645 ;
        RECT 2727.260 1814.305 2727.435 1814.475 ;
        RECT 2726.015 1814.135 2727.435 1814.305 ;
        RECT 2726.015 1813.655 2726.185 1814.135 ;
        RECT 2726.855 1813.660 2727.025 1814.135 ;
        RECT 2697.075 1812.765 2697.245 1813.145 ;
        RECT 2697.075 1812.595 2697.740 1812.765 ;
        RECT 2697.935 1812.640 2698.195 1813.145 ;
        RECT 2697.005 1812.045 2697.335 1812.415 ;
        RECT 2697.570 1812.340 2697.740 1812.595 ;
        RECT 2697.570 1812.010 2697.855 1812.340 ;
        RECT 2697.570 1811.865 2697.740 1812.010 ;
        RECT 2697.075 1811.695 2697.740 1811.865 ;
        RECT 2698.025 1811.840 2698.195 1812.640 ;
        RECT 2697.075 1810.935 2697.245 1811.695 ;
        RECT 2697.925 1810.935 2698.195 1811.840 ;
        RECT 2697.310 1807.305 2697.480 1807.555 ;
        RECT 2522.640 1804.985 2523.160 1806.470 ;
        RECT 2523.330 1805.645 2523.850 1807.195 ;
        RECT 2696.985 1807.135 2697.480 1807.305 ;
        RECT 2698.215 1807.305 2698.385 1807.650 ;
        RECT 2699.055 1807.305 2699.575 1807.705 ;
        RECT 2698.215 1807.135 2699.575 1807.305 ;
        RECT 2696.985 1806.175 2697.155 1807.135 ;
        RECT 2697.325 1806.345 2697.675 1806.965 ;
        RECT 2697.845 1806.345 2698.185 1806.965 ;
        RECT 2698.355 1806.345 2698.595 1806.965 ;
        RECT 2698.775 1806.715 2699.235 1806.885 ;
        RECT 2698.775 1806.175 2698.945 1806.715 ;
        RECT 2699.405 1806.515 2699.575 1807.135 ;
        RECT 2696.985 1806.005 2698.945 1806.175 ;
        RECT 2699.115 1805.505 2699.575 1806.515 ;
        RECT 2697.075 1804.225 2697.245 1804.985 ;
        RECT 2697.075 1804.055 2697.740 1804.225 ;
        RECT 2697.925 1804.080 2698.195 1804.985 ;
        RECT 2697.570 1803.910 2697.740 1804.055 ;
        RECT 2697.005 1803.505 2697.335 1803.875 ;
        RECT 2697.570 1803.580 2697.855 1803.910 ;
        RECT 2697.570 1803.325 2697.740 1803.580 ;
        RECT 2697.075 1803.155 2697.740 1803.325 ;
        RECT 2698.025 1803.280 2698.195 1804.080 ;
        RECT 2697.075 1802.775 2697.245 1803.155 ;
        RECT 2697.935 1802.775 2698.195 1803.280 ;
        RECT 2697.260 1801.625 2697.505 1802.230 ;
        RECT 2696.985 1801.455 2698.215 1801.625 ;
        RECT 2696.985 1800.645 2697.325 1801.455 ;
        RECT 2697.495 1800.890 2698.245 1801.080 ;
        RECT 2696.985 1800.235 2697.500 1800.645 ;
        RECT 2698.075 1800.225 2698.245 1800.890 ;
        RECT 2698.415 1800.905 2698.605 1802.265 ;
        RECT 2698.775 1802.095 2699.050 1802.265 ;
        RECT 2698.775 1801.925 2699.055 1802.095 ;
        RECT 2698.775 1801.105 2699.050 1801.925 ;
        RECT 2699.240 1801.900 2699.770 1802.265 ;
        RECT 2699.595 1801.865 2699.770 1801.900 ;
        RECT 2699.255 1800.905 2699.425 1801.705 ;
        RECT 2698.415 1800.735 2699.425 1800.905 ;
        RECT 2699.595 1801.695 2700.525 1801.865 ;
        RECT 2700.695 1801.695 2700.950 1802.265 ;
        RECT 2699.595 1800.565 2699.765 1801.695 ;
        RECT 2700.355 1801.525 2700.525 1801.695 ;
        RECT 2698.640 1800.395 2699.765 1800.565 ;
        RECT 2699.935 1801.195 2700.130 1801.525 ;
        RECT 2700.355 1801.195 2700.610 1801.525 ;
        RECT 2699.935 1800.225 2700.105 1801.195 ;
        RECT 2700.780 1801.025 2700.950 1801.695 ;
        RECT 2701.630 1801.500 2701.815 1802.170 ;
        RECT 2702.300 1801.815 2702.630 1802.215 ;
        RECT 2703.345 1801.820 2703.675 1802.260 ;
        RECT 2703.345 1801.815 2704.575 1801.820 ;
        RECT 2702.300 1801.705 2704.575 1801.815 ;
        RECT 2702.420 1801.640 2704.575 1801.705 ;
        RECT 2701.180 1801.230 2701.815 1801.500 ;
        RECT 2701.995 1801.120 2702.280 1801.525 ;
        RECT 2702.450 1801.120 2702.780 1801.470 ;
        RECT 2698.075 1800.055 2700.105 1800.225 ;
        RECT 2700.615 1800.055 2700.950 1801.025 ;
        RECT 2701.215 1800.770 2702.325 1800.940 ;
        RECT 2701.215 1800.060 2701.410 1800.770 ;
        RECT 2702.095 1800.060 2702.325 1800.770 ;
        RECT 2702.505 1800.065 2702.780 1801.120 ;
        RECT 2702.950 1800.065 2703.285 1801.470 ;
        RECT 2703.485 1800.065 2703.935 1801.470 ;
        RECT 2704.190 1800.060 2704.575 1801.640 ;
        RECT 2522.640 1797.455 2523.160 1798.940 ;
        RECT 2523.330 1798.115 2523.850 1799.665 ;
        RECT 2696.985 1798.155 2697.325 1799.035 ;
        RECT 2697.495 1798.325 2697.665 1799.545 ;
        RECT 2698.690 1799.205 2699.165 1799.545 ;
        RECT 2697.905 1798.675 2698.155 1799.040 ;
        RECT 2698.875 1798.675 2699.590 1798.970 ;
        RECT 2699.760 1798.845 2700.035 1799.545 ;
        RECT 2697.905 1798.505 2699.695 1798.675 ;
        RECT 2697.495 1798.075 2698.290 1798.325 ;
        RECT 2697.495 1797.985 2697.745 1798.075 ;
        RECT 2697.415 1797.565 2697.745 1797.985 ;
        RECT 2698.460 1797.650 2698.715 1798.505 ;
        RECT 2697.925 1797.385 2698.715 1797.650 ;
        RECT 2698.885 1797.805 2699.295 1798.325 ;
        RECT 2699.465 1798.075 2699.695 1798.505 ;
        RECT 2699.865 1797.815 2700.035 1798.845 ;
        RECT 2698.885 1797.385 2699.085 1797.805 ;
        RECT 2699.775 1797.335 2700.035 1797.815 ;
        RECT 2697.075 1796.445 2697.245 1796.825 ;
        RECT 2697.075 1796.275 2697.740 1796.445 ;
        RECT 2697.935 1796.320 2698.195 1796.825 ;
        RECT 2697.005 1795.725 2697.335 1796.095 ;
        RECT 2697.570 1796.020 2697.740 1796.275 ;
        RECT 2697.570 1795.690 2697.855 1796.020 ;
        RECT 2697.570 1795.545 2697.740 1795.690 ;
        RECT 2697.075 1795.375 2697.740 1795.545 ;
        RECT 2698.025 1795.520 2698.195 1796.320 ;
        RECT 2697.075 1794.615 2697.245 1795.375 ;
        RECT 2697.925 1794.615 2698.195 1795.520 ;
        RECT 2522.640 1791.475 2523.160 1792.960 ;
        RECT 2523.330 1792.135 2523.850 1793.685 ;
        RECT 2698.455 1793.605 2698.625 1794.105 ;
        RECT 2699.415 1793.605 2699.585 1794.105 ;
        RECT 2700.255 1793.605 2700.425 1794.105 ;
        RECT 2698.455 1793.435 2700.425 1793.605 ;
        RECT 2700.595 1793.635 2700.925 1794.065 ;
        RECT 2701.535 1793.805 2701.875 1794.065 ;
        RECT 2700.595 1793.465 2701.445 1793.635 ;
        RECT 2698.390 1792.635 2698.645 1793.265 ;
        RECT 2698.875 1792.635 2699.255 1793.265 ;
        RECT 2700.125 1793.255 2700.425 1793.260 ;
        RECT 2700.125 1793.085 2700.435 1793.255 ;
        RECT 2700.125 1792.965 2700.425 1793.085 ;
        RECT 2698.875 1792.035 2699.080 1792.635 ;
        RECT 2699.515 1792.240 2699.735 1792.965 ;
        RECT 2700.045 1792.635 2700.425 1792.965 ;
        RECT 2700.625 1792.715 2700.955 1793.275 ;
        RECT 2701.275 1792.545 2701.445 1793.465 ;
        RECT 2700.625 1792.450 2701.445 1792.545 ;
        RECT 2700.430 1792.375 2701.445 1792.450 ;
        RECT 2699.310 1792.055 2700.260 1792.240 ;
        RECT 2700.430 1791.940 2700.845 1792.375 ;
        RECT 2701.615 1792.200 2701.875 1793.805 ;
        RECT 2701.535 1791.940 2701.875 1792.200 ;
        RECT 2698.335 1790.735 2698.665 1791.155 ;
        RECT 2698.845 1790.985 2699.105 1791.385 ;
        RECT 2699.775 1790.985 2699.945 1791.335 ;
        RECT 2698.845 1790.815 2700.510 1790.985 ;
        RECT 2700.680 1790.880 2700.955 1791.225 ;
        RECT 2698.415 1790.645 2698.665 1790.735 ;
        RECT 2700.340 1790.645 2700.510 1790.815 ;
        RECT 2368.595 1790.110 2368.770 1790.600 ;
        RECT 2369.120 1790.320 2369.290 1790.600 ;
        RECT 2369.120 1790.150 2369.350 1790.320 ;
        RECT 2368.595 1789.940 2368.765 1790.110 ;
        RECT 2368.595 1789.610 2369.005 1789.940 ;
        RECT 2368.595 1789.100 2368.765 1789.610 ;
        RECT 2368.595 1788.770 2369.005 1789.100 ;
        RECT 2368.595 1788.570 2368.765 1788.770 ;
        RECT 2368.595 1787.310 2368.770 1788.570 ;
        RECT 2369.180 1788.540 2369.350 1790.150 ;
        RECT 2369.550 1790.090 2369.725 1790.600 ;
        RECT 2376.110 1790.110 2376.285 1790.600 ;
        RECT 2376.110 1789.940 2376.280 1790.110 ;
        RECT 2377.065 1790.090 2377.240 1790.600 ;
        RECT 2377.495 1790.050 2377.670 1790.600 ;
        RECT 2381.725 1790.110 2381.900 1790.600 ;
        RECT 2382.250 1790.320 2382.420 1790.600 ;
        RECT 2382.250 1790.150 2382.480 1790.320 ;
        RECT 2376.110 1789.610 2376.520 1789.940 ;
        RECT 2369.120 1788.370 2369.350 1788.540 ;
        RECT 2369.550 1788.570 2369.720 1789.520 ;
        RECT 2376.110 1789.100 2376.280 1789.610 ;
        RECT 2376.110 1788.770 2376.520 1789.100 ;
        RECT 2376.110 1788.570 2376.280 1788.770 ;
        RECT 2377.065 1788.570 2377.235 1789.520 ;
        RECT 2369.120 1787.310 2369.290 1788.370 ;
        RECT 2369.550 1787.310 2369.725 1788.570 ;
        RECT 2376.110 1787.310 2376.285 1788.570 ;
        RECT 2377.065 1787.310 2377.240 1788.570 ;
        RECT 2377.495 1788.450 2377.665 1790.050 ;
        RECT 2381.725 1789.940 2381.895 1790.110 ;
        RECT 2381.725 1789.610 2382.135 1789.940 ;
        RECT 2381.725 1789.100 2381.895 1789.610 ;
        RECT 2381.725 1788.770 2382.135 1789.100 ;
        RECT 2381.725 1788.570 2381.895 1788.770 ;
        RECT 2377.495 1787.310 2377.670 1788.450 ;
        RECT 2381.725 1787.310 2381.900 1788.570 ;
        RECT 2382.310 1788.540 2382.480 1790.150 ;
        RECT 2382.680 1790.090 2382.855 1790.600 ;
        RECT 2383.110 1790.050 2383.285 1790.600 ;
        RECT 2384.475 1790.090 2384.645 1790.600 ;
        RECT 2385.465 1790.090 2385.635 1790.600 ;
        RECT 2391.370 1790.110 2391.545 1790.600 ;
        RECT 2382.250 1788.370 2382.480 1788.540 ;
        RECT 2382.680 1788.570 2382.850 1789.520 ;
        RECT 2382.250 1787.310 2382.420 1788.370 ;
        RECT 2382.680 1787.310 2382.855 1788.570 ;
        RECT 2383.110 1788.450 2383.280 1790.050 ;
        RECT 2391.370 1789.940 2391.540 1790.110 ;
        RECT 2392.325 1790.090 2392.500 1790.600 ;
        RECT 2392.755 1790.050 2392.930 1790.600 ;
        RECT 2396.985 1790.110 2397.160 1790.600 ;
        RECT 2397.510 1790.320 2397.680 1790.600 ;
        RECT 2397.510 1790.150 2397.740 1790.320 ;
        RECT 2391.370 1789.610 2391.780 1789.940 ;
        RECT 2383.650 1789.430 2383.880 1789.580 ;
        RECT 2383.650 1789.260 2384.570 1789.430 ;
        RECT 2385.090 1789.260 2385.560 1789.430 ;
        RECT 2384.100 1788.570 2384.270 1789.260 ;
        RECT 2384.470 1788.780 2384.640 1788.890 ;
        RECT 2385.090 1788.780 2385.260 1789.260 ;
        RECT 2391.370 1789.100 2391.540 1789.610 ;
        RECT 2384.470 1788.610 2385.260 1788.780 ;
        RECT 2383.110 1787.310 2383.285 1788.450 ;
        RECT 2384.470 1787.310 2384.645 1788.610 ;
        RECT 2385.090 1788.570 2385.260 1788.610 ;
        RECT 2385.460 1788.455 2385.630 1788.890 ;
        RECT 2391.370 1788.770 2391.780 1789.100 ;
        RECT 2391.370 1788.570 2391.540 1788.770 ;
        RECT 2392.325 1788.570 2392.495 1789.520 ;
        RECT 2385.460 1787.310 2385.635 1788.455 ;
        RECT 2391.370 1787.310 2391.545 1788.570 ;
        RECT 2392.325 1787.310 2392.500 1788.570 ;
        RECT 2392.755 1788.450 2392.925 1790.050 ;
        RECT 2396.985 1789.940 2397.155 1790.110 ;
        RECT 2396.985 1789.610 2397.395 1789.940 ;
        RECT 2396.985 1789.100 2397.155 1789.610 ;
        RECT 2396.985 1788.770 2397.395 1789.100 ;
        RECT 2396.985 1788.570 2397.155 1788.770 ;
        RECT 2392.755 1787.310 2392.930 1788.450 ;
        RECT 2396.985 1787.310 2397.160 1788.570 ;
        RECT 2397.570 1788.540 2397.740 1790.150 ;
        RECT 2397.940 1790.090 2398.115 1790.600 ;
        RECT 2398.370 1790.050 2398.545 1790.600 ;
        RECT 2399.735 1790.090 2399.905 1790.600 ;
        RECT 2400.725 1790.090 2400.895 1790.600 ;
        RECT 2406.630 1790.110 2406.805 1790.600 ;
        RECT 2397.510 1788.370 2397.740 1788.540 ;
        RECT 2397.940 1788.570 2398.110 1789.520 ;
        RECT 2397.510 1787.310 2397.680 1788.370 ;
        RECT 2397.940 1787.310 2398.115 1788.570 ;
        RECT 2398.370 1788.450 2398.540 1790.050 ;
        RECT 2406.630 1789.940 2406.800 1790.110 ;
        RECT 2407.585 1790.090 2407.760 1790.600 ;
        RECT 2408.015 1790.050 2408.190 1790.600 ;
        RECT 2412.245 1790.110 2412.420 1790.600 ;
        RECT 2412.770 1790.320 2412.940 1790.600 ;
        RECT 2412.770 1790.150 2413.000 1790.320 ;
        RECT 2406.630 1789.610 2407.040 1789.940 ;
        RECT 2398.910 1789.430 2399.140 1789.580 ;
        RECT 2398.910 1789.260 2399.830 1789.430 ;
        RECT 2400.350 1789.260 2400.820 1789.430 ;
        RECT 2399.360 1788.570 2399.530 1789.260 ;
        RECT 2399.730 1788.780 2399.900 1788.890 ;
        RECT 2400.350 1788.780 2400.520 1789.260 ;
        RECT 2406.630 1789.100 2406.800 1789.610 ;
        RECT 2399.730 1788.610 2400.520 1788.780 ;
        RECT 2398.370 1787.310 2398.545 1788.450 ;
        RECT 2399.730 1787.310 2399.905 1788.610 ;
        RECT 2400.350 1788.570 2400.520 1788.610 ;
        RECT 2400.720 1788.455 2400.890 1788.890 ;
        RECT 2406.630 1788.770 2407.040 1789.100 ;
        RECT 2406.630 1788.570 2406.800 1788.770 ;
        RECT 2407.585 1788.570 2407.755 1789.520 ;
        RECT 2400.720 1787.310 2400.895 1788.455 ;
        RECT 2406.630 1787.310 2406.805 1788.570 ;
        RECT 2407.585 1787.310 2407.760 1788.570 ;
        RECT 2408.015 1788.450 2408.185 1790.050 ;
        RECT 2412.245 1789.940 2412.415 1790.110 ;
        RECT 2412.245 1789.610 2412.655 1789.940 ;
        RECT 2412.245 1789.100 2412.415 1789.610 ;
        RECT 2412.245 1788.770 2412.655 1789.100 ;
        RECT 2412.245 1788.570 2412.415 1788.770 ;
        RECT 2408.015 1787.310 2408.190 1788.450 ;
        RECT 2412.245 1787.310 2412.420 1788.570 ;
        RECT 2412.830 1788.540 2413.000 1790.150 ;
        RECT 2413.200 1790.090 2413.375 1790.600 ;
        RECT 2413.630 1790.050 2413.805 1790.600 ;
        RECT 2414.995 1790.090 2415.165 1790.600 ;
        RECT 2415.985 1790.090 2416.155 1790.600 ;
        RECT 2421.890 1790.110 2422.065 1790.600 ;
        RECT 2412.770 1788.370 2413.000 1788.540 ;
        RECT 2413.200 1788.570 2413.370 1789.520 ;
        RECT 2412.770 1787.310 2412.940 1788.370 ;
        RECT 2413.200 1787.310 2413.375 1788.570 ;
        RECT 2413.630 1788.450 2413.800 1790.050 ;
        RECT 2421.890 1789.940 2422.060 1790.110 ;
        RECT 2422.845 1790.090 2423.020 1790.600 ;
        RECT 2423.275 1790.050 2423.450 1790.600 ;
        RECT 2427.505 1790.110 2427.680 1790.600 ;
        RECT 2428.030 1790.320 2428.200 1790.600 ;
        RECT 2428.030 1790.150 2428.260 1790.320 ;
        RECT 2421.890 1789.610 2422.300 1789.940 ;
        RECT 2414.170 1789.430 2414.400 1789.580 ;
        RECT 2414.170 1789.260 2415.090 1789.430 ;
        RECT 2415.610 1789.260 2416.080 1789.430 ;
        RECT 2414.620 1788.570 2414.790 1789.260 ;
        RECT 2414.990 1788.780 2415.160 1788.890 ;
        RECT 2415.610 1788.780 2415.780 1789.260 ;
        RECT 2421.890 1789.100 2422.060 1789.610 ;
        RECT 2414.990 1788.610 2415.780 1788.780 ;
        RECT 2413.630 1787.310 2413.805 1788.450 ;
        RECT 2414.990 1787.310 2415.165 1788.610 ;
        RECT 2415.610 1788.570 2415.780 1788.610 ;
        RECT 2415.980 1788.455 2416.150 1788.890 ;
        RECT 2421.890 1788.770 2422.300 1789.100 ;
        RECT 2421.890 1788.570 2422.060 1788.770 ;
        RECT 2422.845 1788.570 2423.015 1789.520 ;
        RECT 2415.980 1787.310 2416.155 1788.455 ;
        RECT 2421.890 1787.310 2422.065 1788.570 ;
        RECT 2422.845 1787.310 2423.020 1788.570 ;
        RECT 2423.275 1788.450 2423.445 1790.050 ;
        RECT 2427.505 1789.940 2427.675 1790.110 ;
        RECT 2427.505 1789.610 2427.915 1789.940 ;
        RECT 2427.505 1789.100 2427.675 1789.610 ;
        RECT 2427.505 1788.770 2427.915 1789.100 ;
        RECT 2427.505 1788.570 2427.675 1788.770 ;
        RECT 2423.275 1787.310 2423.450 1788.450 ;
        RECT 2427.505 1787.310 2427.680 1788.570 ;
        RECT 2428.090 1788.540 2428.260 1790.150 ;
        RECT 2428.460 1790.090 2428.635 1790.600 ;
        RECT 2428.890 1790.050 2429.065 1790.600 ;
        RECT 2430.255 1790.090 2430.425 1790.600 ;
        RECT 2431.245 1790.090 2431.415 1790.600 ;
        RECT 2437.150 1790.110 2437.325 1790.600 ;
        RECT 2428.030 1788.370 2428.260 1788.540 ;
        RECT 2428.460 1788.570 2428.630 1789.520 ;
        RECT 2428.030 1787.310 2428.200 1788.370 ;
        RECT 2428.460 1787.310 2428.635 1788.570 ;
        RECT 2428.890 1788.450 2429.060 1790.050 ;
        RECT 2437.150 1789.940 2437.320 1790.110 ;
        RECT 2438.105 1790.090 2438.280 1790.600 ;
        RECT 2438.535 1790.050 2438.710 1790.600 ;
        RECT 2442.765 1790.110 2442.940 1790.600 ;
        RECT 2443.290 1790.320 2443.460 1790.600 ;
        RECT 2443.290 1790.150 2443.520 1790.320 ;
        RECT 2437.150 1789.610 2437.560 1789.940 ;
        RECT 2429.430 1789.430 2429.660 1789.580 ;
        RECT 2429.430 1789.260 2430.350 1789.430 ;
        RECT 2430.870 1789.260 2431.340 1789.430 ;
        RECT 2429.880 1788.570 2430.050 1789.260 ;
        RECT 2430.250 1788.780 2430.420 1788.890 ;
        RECT 2430.870 1788.780 2431.040 1789.260 ;
        RECT 2437.150 1789.100 2437.320 1789.610 ;
        RECT 2430.250 1788.610 2431.040 1788.780 ;
        RECT 2428.890 1787.310 2429.065 1788.450 ;
        RECT 2430.250 1787.310 2430.425 1788.610 ;
        RECT 2430.870 1788.570 2431.040 1788.610 ;
        RECT 2431.240 1788.455 2431.410 1788.890 ;
        RECT 2437.150 1788.770 2437.560 1789.100 ;
        RECT 2437.150 1788.570 2437.320 1788.770 ;
        RECT 2438.105 1788.570 2438.275 1789.520 ;
        RECT 2431.240 1787.310 2431.415 1788.455 ;
        RECT 2437.150 1787.310 2437.325 1788.570 ;
        RECT 2438.105 1787.310 2438.280 1788.570 ;
        RECT 2438.535 1788.450 2438.705 1790.050 ;
        RECT 2442.765 1789.940 2442.935 1790.110 ;
        RECT 2442.765 1789.610 2443.175 1789.940 ;
        RECT 2442.765 1789.100 2442.935 1789.610 ;
        RECT 2442.765 1788.770 2443.175 1789.100 ;
        RECT 2442.765 1788.570 2442.935 1788.770 ;
        RECT 2438.535 1787.310 2438.710 1788.450 ;
        RECT 2442.765 1787.310 2442.940 1788.570 ;
        RECT 2443.350 1788.540 2443.520 1790.150 ;
        RECT 2443.720 1790.090 2443.895 1790.600 ;
        RECT 2444.150 1790.050 2444.325 1790.600 ;
        RECT 2445.515 1790.090 2445.685 1790.600 ;
        RECT 2446.505 1790.090 2446.675 1790.600 ;
        RECT 2697.910 1790.315 2698.245 1790.565 ;
        RECT 2698.415 1790.315 2699.130 1790.645 ;
        RECT 2699.345 1790.315 2700.170 1790.645 ;
        RECT 2700.340 1790.315 2700.615 1790.645 ;
        RECT 2443.290 1788.370 2443.520 1788.540 ;
        RECT 2443.720 1788.570 2443.890 1789.520 ;
        RECT 2443.290 1787.310 2443.460 1788.370 ;
        RECT 2443.720 1787.310 2443.895 1788.570 ;
        RECT 2444.150 1788.450 2444.320 1790.050 ;
        RECT 2698.415 1789.755 2698.585 1790.315 ;
        RECT 2698.845 1789.855 2699.175 1790.145 ;
        RECT 2699.345 1790.025 2699.590 1790.315 ;
        RECT 2700.340 1790.145 2700.510 1790.315 ;
        RECT 2700.785 1790.145 2700.955 1790.880 ;
        RECT 2699.850 1789.975 2700.510 1790.145 ;
        RECT 2699.850 1789.855 2700.020 1789.975 ;
        RECT 2698.845 1789.685 2700.020 1789.855 ;
        RECT 2444.690 1789.430 2444.920 1789.580 ;
        RECT 2444.690 1789.260 2445.610 1789.430 ;
        RECT 2446.130 1789.260 2446.600 1789.430 ;
        RECT 2445.140 1788.570 2445.310 1789.260 ;
        RECT 2445.510 1788.780 2445.680 1788.890 ;
        RECT 2446.130 1788.780 2446.300 1789.260 ;
        RECT 2698.405 1789.185 2700.020 1789.515 ;
        RECT 2700.680 1789.175 2700.955 1790.145 ;
        RECT 2701.125 1791.155 2701.715 1791.385 ;
        RECT 2701.125 1790.145 2701.415 1791.155 ;
        RECT 2703.290 1790.985 2703.715 1791.195 ;
        RECT 2701.585 1790.815 2703.715 1790.985 ;
        RECT 2701.585 1790.315 2701.755 1790.815 ;
        RECT 2702.045 1790.315 2702.375 1790.645 ;
        RECT 2702.565 1790.315 2702.835 1790.645 ;
        RECT 2703.025 1790.315 2703.375 1790.645 ;
        RECT 2701.125 1789.975 2702.670 1790.145 ;
        RECT 2703.545 1790.045 2703.715 1790.815 ;
        RECT 2701.125 1789.175 2701.715 1789.975 ;
        RECT 2702.340 1789.175 2702.670 1789.975 ;
        RECT 2703.290 1789.715 2703.715 1790.045 ;
        RECT 2445.510 1788.610 2446.300 1788.780 ;
        RECT 2444.150 1787.310 2444.325 1788.450 ;
        RECT 2445.510 1787.310 2445.685 1788.610 ;
        RECT 2446.130 1788.570 2446.300 1788.610 ;
        RECT 2446.500 1788.455 2446.670 1788.890 ;
        RECT 2446.500 1787.310 2446.675 1788.455 ;
        RECT 2697.075 1787.905 2697.245 1788.665 ;
        RECT 2522.640 1785.530 2523.160 1787.015 ;
        RECT 2523.330 1786.190 2523.850 1787.740 ;
        RECT 2697.075 1787.735 2697.740 1787.905 ;
        RECT 2697.925 1787.760 2698.195 1788.665 ;
        RECT 2697.570 1787.590 2697.740 1787.735 ;
        RECT 2697.005 1787.185 2697.335 1787.555 ;
        RECT 2697.570 1787.260 2697.855 1787.590 ;
        RECT 2697.570 1787.005 2697.740 1787.260 ;
        RECT 2697.075 1786.835 2697.740 1787.005 ;
        RECT 2698.025 1786.960 2698.195 1787.760 ;
        RECT 2699.255 1787.685 2699.585 1788.665 ;
        RECT 2698.845 1787.275 2699.180 1787.525 ;
        RECT 2699.350 1787.085 2699.520 1787.685 ;
        RECT 2699.690 1787.255 2700.025 1787.525 ;
        RECT 2697.075 1786.455 2697.245 1786.835 ;
        RECT 2697.935 1786.455 2698.195 1786.960 ;
        RECT 2698.825 1786.455 2699.520 1787.085 ;
        RECT 2697.260 1785.305 2697.505 1785.910 ;
        RECT 2371.825 1784.435 2371.995 1784.795 ;
        RECT 2372.765 1784.435 2372.935 1784.795 ;
        RECT 2373.245 1784.345 2373.415 1784.765 ;
        RECT 2373.605 1784.515 2373.895 1785.075 ;
        RECT 2374.685 1784.775 2374.855 1785.105 ;
        RECT 2375.165 1784.685 2375.335 1785.075 ;
        RECT 2377.060 1784.775 2377.235 1785.105 ;
        RECT 2379.005 1784.905 2379.515 1785.075 ;
        RECT 2377.585 1784.685 2377.765 1784.795 ;
        RECT 2379.345 1784.765 2379.515 1784.905 ;
        RECT 2375.055 1784.515 2375.390 1784.685 ;
        RECT 2375.885 1784.515 2376.375 1784.685 ;
        RECT 2377.585 1784.515 2378.935 1784.685 ;
        RECT 2379.345 1784.515 2379.630 1784.765 ;
        RECT 2373.725 1784.435 2373.895 1784.515 ;
        RECT 2372.525 1783.785 2372.695 1784.235 ;
        RECT 2373.005 1783.785 2373.175 1784.115 ;
        RECT 2373.965 1783.785 2374.135 1784.115 ;
        RECT 2374.445 1783.785 2374.615 1784.515 ;
        RECT 2375.885 1784.345 2376.055 1784.515 ;
        RECT 2377.585 1784.435 2377.765 1784.515 ;
        RECT 2378.765 1784.345 2378.935 1784.515 ;
        RECT 2379.455 1784.435 2379.630 1784.515 ;
        RECT 2374.925 1783.785 2375.095 1784.235 ;
        RECT 2375.405 1783.785 2375.575 1784.115 ;
        RECT 2375.885 1783.785 2376.055 1784.115 ;
        RECT 2376.365 1783.785 2376.535 1784.235 ;
        RECT 2377.325 1784.135 2377.495 1784.235 ;
        RECT 2376.845 1784.035 2377.495 1784.135 ;
        RECT 2376.765 1783.865 2377.575 1784.035 ;
        RECT 2377.805 1783.785 2377.975 1784.115 ;
        RECT 2378.285 1783.785 2378.455 1784.235 ;
        RECT 2378.765 1783.785 2378.935 1784.115 ;
        RECT 2379.245 1784.035 2379.515 1784.235 ;
        RECT 2379.125 1783.825 2379.515 1784.035 ;
        RECT 2381.725 1783.895 2381.900 1785.155 ;
        RECT 2382.250 1784.095 2382.420 1785.155 ;
        RECT 2382.250 1783.925 2382.480 1784.095 ;
        RECT 2381.725 1783.695 2381.895 1783.895 ;
        RECT 2376.845 1783.615 2377.015 1783.655 ;
        RECT 2376.485 1783.445 2377.015 1783.615 ;
        RECT 2371.825 1783.045 2371.995 1783.395 ;
        RECT 2373.725 1783.045 2373.895 1783.395 ;
        RECT 2375.125 1783.375 2375.295 1783.395 ;
        RECT 2375.125 1783.345 2375.335 1783.375 ;
        RECT 2375.025 1783.125 2375.335 1783.345 ;
        RECT 2375.165 1783.045 2375.335 1783.125 ;
        RECT 2376.125 1783.275 2376.295 1783.395 ;
        RECT 2376.125 1783.105 2377.365 1783.275 ;
        RECT 2378.045 1783.045 2378.215 1783.395 ;
        RECT 2379.005 1783.045 2379.175 1783.395 ;
        RECT 2381.725 1783.365 2382.135 1783.695 ;
        RECT 2381.725 1782.855 2381.895 1783.365 ;
        RECT 2381.725 1782.525 2382.135 1782.855 ;
        RECT 2381.725 1782.355 2381.895 1782.525 ;
        RECT 2381.725 1781.865 2381.900 1782.355 ;
        RECT 2382.310 1782.315 2382.480 1783.925 ;
        RECT 2382.680 1783.895 2382.855 1785.155 ;
        RECT 2383.110 1784.015 2383.285 1785.155 ;
        RECT 2382.680 1782.945 2382.850 1783.895 ;
        RECT 2383.110 1782.415 2383.280 1784.015 ;
        RECT 2384.470 1784.010 2384.645 1785.155 ;
        RECT 2385.455 1784.010 2385.630 1785.155 ;
        RECT 2387.085 1784.435 2387.255 1784.795 ;
        RECT 2388.025 1784.435 2388.195 1784.795 ;
        RECT 2388.505 1784.345 2388.675 1784.765 ;
        RECT 2388.865 1784.515 2389.155 1785.075 ;
        RECT 2389.945 1784.775 2390.115 1785.105 ;
        RECT 2390.425 1784.685 2390.595 1785.075 ;
        RECT 2392.320 1784.775 2392.495 1785.105 ;
        RECT 2394.265 1784.905 2394.775 1785.075 ;
        RECT 2392.845 1784.685 2393.025 1784.795 ;
        RECT 2394.605 1784.765 2394.775 1784.905 ;
        RECT 2390.315 1784.515 2390.650 1784.685 ;
        RECT 2391.145 1784.515 2391.635 1784.685 ;
        RECT 2392.845 1784.515 2394.195 1784.685 ;
        RECT 2394.605 1784.515 2394.890 1784.765 ;
        RECT 2388.985 1784.435 2389.155 1784.515 ;
        RECT 2384.100 1783.205 2384.270 1783.895 ;
        RECT 2384.470 1783.795 2384.640 1784.010 ;
        RECT 2385.085 1783.795 2385.255 1783.895 ;
        RECT 2384.470 1783.625 2385.255 1783.795 ;
        RECT 2384.470 1783.575 2384.640 1783.625 ;
        RECT 2385.085 1783.205 2385.255 1783.625 ;
        RECT 2385.455 1783.575 2385.625 1784.010 ;
        RECT 2387.785 1783.785 2387.955 1784.235 ;
        RECT 2388.265 1783.785 2388.435 1784.115 ;
        RECT 2389.225 1783.785 2389.395 1784.115 ;
        RECT 2389.705 1783.785 2389.875 1784.515 ;
        RECT 2391.145 1784.345 2391.315 1784.515 ;
        RECT 2392.845 1784.435 2393.025 1784.515 ;
        RECT 2394.025 1784.345 2394.195 1784.515 ;
        RECT 2394.715 1784.435 2394.890 1784.515 ;
        RECT 2390.185 1783.785 2390.355 1784.235 ;
        RECT 2390.665 1783.785 2390.835 1784.115 ;
        RECT 2391.145 1783.785 2391.315 1784.115 ;
        RECT 2391.625 1783.785 2391.795 1784.235 ;
        RECT 2392.585 1784.135 2392.755 1784.235 ;
        RECT 2392.105 1784.035 2392.755 1784.135 ;
        RECT 2392.025 1783.865 2392.835 1784.035 ;
        RECT 2393.065 1783.785 2393.235 1784.115 ;
        RECT 2393.545 1783.785 2393.715 1784.235 ;
        RECT 2394.025 1783.785 2394.195 1784.115 ;
        RECT 2394.505 1784.035 2394.775 1784.235 ;
        RECT 2394.385 1783.825 2394.775 1784.035 ;
        RECT 2396.985 1783.895 2397.160 1785.155 ;
        RECT 2397.510 1784.095 2397.680 1785.155 ;
        RECT 2397.510 1783.925 2397.740 1784.095 ;
        RECT 2396.985 1783.695 2397.155 1783.895 ;
        RECT 2392.105 1783.615 2392.275 1783.655 ;
        RECT 2391.745 1783.445 2392.275 1783.615 ;
        RECT 2383.650 1783.035 2384.570 1783.205 ;
        RECT 2385.085 1783.035 2385.555 1783.205 ;
        RECT 2387.085 1783.045 2387.255 1783.395 ;
        RECT 2388.985 1783.045 2389.155 1783.395 ;
        RECT 2390.385 1783.375 2390.555 1783.395 ;
        RECT 2390.385 1783.345 2390.595 1783.375 ;
        RECT 2390.285 1783.125 2390.595 1783.345 ;
        RECT 2390.425 1783.045 2390.595 1783.125 ;
        RECT 2391.385 1783.275 2391.555 1783.395 ;
        RECT 2391.385 1783.105 2392.625 1783.275 ;
        RECT 2393.305 1783.045 2393.475 1783.395 ;
        RECT 2394.265 1783.045 2394.435 1783.395 ;
        RECT 2396.985 1783.365 2397.395 1783.695 ;
        RECT 2383.650 1782.885 2383.880 1783.035 ;
        RECT 2396.985 1782.855 2397.155 1783.365 ;
        RECT 2396.985 1782.525 2397.395 1782.855 ;
        RECT 2382.250 1782.145 2382.480 1782.315 ;
        RECT 2382.250 1781.865 2382.420 1782.145 ;
        RECT 2382.680 1781.865 2382.855 1782.375 ;
        RECT 2383.110 1781.865 2383.285 1782.415 ;
        RECT 2384.475 1781.865 2384.645 1782.375 ;
        RECT 2385.460 1781.865 2385.630 1782.375 ;
        RECT 2396.985 1782.355 2397.155 1782.525 ;
        RECT 2396.985 1781.865 2397.160 1782.355 ;
        RECT 2397.570 1782.315 2397.740 1783.925 ;
        RECT 2397.940 1783.895 2398.115 1785.155 ;
        RECT 2398.370 1784.015 2398.545 1785.155 ;
        RECT 2397.940 1782.945 2398.110 1783.895 ;
        RECT 2398.370 1782.415 2398.540 1784.015 ;
        RECT 2399.730 1784.010 2399.905 1785.155 ;
        RECT 2400.715 1784.010 2400.890 1785.155 ;
        RECT 2402.345 1784.435 2402.515 1784.795 ;
        RECT 2403.285 1784.435 2403.455 1784.795 ;
        RECT 2403.765 1784.345 2403.935 1784.765 ;
        RECT 2404.125 1784.515 2404.415 1785.075 ;
        RECT 2405.205 1784.775 2405.375 1785.105 ;
        RECT 2405.685 1784.685 2405.855 1785.075 ;
        RECT 2407.580 1784.775 2407.755 1785.105 ;
        RECT 2409.525 1784.905 2410.035 1785.075 ;
        RECT 2408.105 1784.685 2408.285 1784.795 ;
        RECT 2409.865 1784.765 2410.035 1784.905 ;
        RECT 2405.575 1784.515 2405.910 1784.685 ;
        RECT 2406.405 1784.515 2406.895 1784.685 ;
        RECT 2408.105 1784.515 2409.455 1784.685 ;
        RECT 2409.865 1784.515 2410.150 1784.765 ;
        RECT 2404.245 1784.435 2404.415 1784.515 ;
        RECT 2399.360 1783.205 2399.530 1783.895 ;
        RECT 2399.730 1783.795 2399.900 1784.010 ;
        RECT 2400.345 1783.795 2400.515 1783.895 ;
        RECT 2399.730 1783.625 2400.515 1783.795 ;
        RECT 2399.730 1783.575 2399.900 1783.625 ;
        RECT 2400.345 1783.205 2400.515 1783.625 ;
        RECT 2400.715 1783.575 2400.885 1784.010 ;
        RECT 2403.045 1783.785 2403.215 1784.235 ;
        RECT 2403.525 1783.785 2403.695 1784.115 ;
        RECT 2404.485 1783.785 2404.655 1784.115 ;
        RECT 2404.965 1783.785 2405.135 1784.515 ;
        RECT 2406.405 1784.345 2406.575 1784.515 ;
        RECT 2408.105 1784.435 2408.285 1784.515 ;
        RECT 2409.285 1784.345 2409.455 1784.515 ;
        RECT 2409.975 1784.435 2410.150 1784.515 ;
        RECT 2405.445 1783.785 2405.615 1784.235 ;
        RECT 2405.925 1783.785 2406.095 1784.115 ;
        RECT 2406.405 1783.785 2406.575 1784.115 ;
        RECT 2406.885 1783.785 2407.055 1784.235 ;
        RECT 2407.845 1784.135 2408.015 1784.235 ;
        RECT 2407.365 1784.035 2408.015 1784.135 ;
        RECT 2407.285 1783.865 2408.095 1784.035 ;
        RECT 2408.325 1783.785 2408.495 1784.115 ;
        RECT 2408.805 1783.785 2408.975 1784.235 ;
        RECT 2409.285 1783.785 2409.455 1784.115 ;
        RECT 2409.765 1784.035 2410.035 1784.235 ;
        RECT 2409.645 1783.825 2410.035 1784.035 ;
        RECT 2412.245 1783.895 2412.420 1785.155 ;
        RECT 2412.770 1784.095 2412.940 1785.155 ;
        RECT 2412.770 1783.925 2413.000 1784.095 ;
        RECT 2412.245 1783.695 2412.415 1783.895 ;
        RECT 2407.365 1783.615 2407.535 1783.655 ;
        RECT 2407.005 1783.445 2407.535 1783.615 ;
        RECT 2398.910 1783.035 2399.830 1783.205 ;
        RECT 2400.345 1783.035 2400.815 1783.205 ;
        RECT 2402.345 1783.045 2402.515 1783.395 ;
        RECT 2404.245 1783.045 2404.415 1783.395 ;
        RECT 2405.645 1783.375 2405.815 1783.395 ;
        RECT 2405.645 1783.345 2405.855 1783.375 ;
        RECT 2405.545 1783.125 2405.855 1783.345 ;
        RECT 2405.685 1783.045 2405.855 1783.125 ;
        RECT 2406.645 1783.275 2406.815 1783.395 ;
        RECT 2406.645 1783.105 2407.885 1783.275 ;
        RECT 2408.565 1783.045 2408.735 1783.395 ;
        RECT 2409.525 1783.045 2409.695 1783.395 ;
        RECT 2412.245 1783.365 2412.655 1783.695 ;
        RECT 2398.910 1782.885 2399.140 1783.035 ;
        RECT 2412.245 1782.855 2412.415 1783.365 ;
        RECT 2412.245 1782.525 2412.655 1782.855 ;
        RECT 2397.510 1782.145 2397.740 1782.315 ;
        RECT 2397.510 1781.865 2397.680 1782.145 ;
        RECT 2397.940 1781.865 2398.115 1782.375 ;
        RECT 2398.370 1781.865 2398.545 1782.415 ;
        RECT 2399.735 1781.865 2399.905 1782.375 ;
        RECT 2400.720 1781.865 2400.890 1782.375 ;
        RECT 2412.245 1782.355 2412.415 1782.525 ;
        RECT 2412.245 1781.865 2412.420 1782.355 ;
        RECT 2412.830 1782.315 2413.000 1783.925 ;
        RECT 2413.200 1783.895 2413.375 1785.155 ;
        RECT 2413.630 1784.015 2413.805 1785.155 ;
        RECT 2413.200 1782.945 2413.370 1783.895 ;
        RECT 2413.630 1782.415 2413.800 1784.015 ;
        RECT 2414.990 1784.010 2415.165 1785.155 ;
        RECT 2415.975 1784.010 2416.150 1785.155 ;
        RECT 2417.605 1784.435 2417.775 1784.795 ;
        RECT 2418.545 1784.435 2418.715 1784.795 ;
        RECT 2419.025 1784.345 2419.195 1784.765 ;
        RECT 2419.385 1784.515 2419.675 1785.075 ;
        RECT 2420.465 1784.775 2420.635 1785.105 ;
        RECT 2420.945 1784.685 2421.115 1785.075 ;
        RECT 2422.840 1784.775 2423.015 1785.105 ;
        RECT 2424.785 1784.905 2425.295 1785.075 ;
        RECT 2423.365 1784.685 2423.545 1784.795 ;
        RECT 2425.125 1784.765 2425.295 1784.905 ;
        RECT 2420.835 1784.515 2421.170 1784.685 ;
        RECT 2421.665 1784.515 2422.155 1784.685 ;
        RECT 2423.365 1784.515 2424.715 1784.685 ;
        RECT 2425.125 1784.515 2425.410 1784.765 ;
        RECT 2419.505 1784.435 2419.675 1784.515 ;
        RECT 2414.620 1783.205 2414.790 1783.895 ;
        RECT 2414.990 1783.795 2415.160 1784.010 ;
        RECT 2415.605 1783.795 2415.775 1783.895 ;
        RECT 2414.990 1783.625 2415.775 1783.795 ;
        RECT 2414.990 1783.575 2415.160 1783.625 ;
        RECT 2415.605 1783.205 2415.775 1783.625 ;
        RECT 2415.975 1783.575 2416.145 1784.010 ;
        RECT 2418.305 1783.785 2418.475 1784.235 ;
        RECT 2418.785 1783.785 2418.955 1784.115 ;
        RECT 2419.745 1783.785 2419.915 1784.115 ;
        RECT 2420.225 1783.785 2420.395 1784.515 ;
        RECT 2421.665 1784.345 2421.835 1784.515 ;
        RECT 2423.365 1784.435 2423.545 1784.515 ;
        RECT 2424.545 1784.345 2424.715 1784.515 ;
        RECT 2425.235 1784.435 2425.410 1784.515 ;
        RECT 2420.705 1783.785 2420.875 1784.235 ;
        RECT 2421.185 1783.785 2421.355 1784.115 ;
        RECT 2421.665 1783.785 2421.835 1784.115 ;
        RECT 2422.145 1783.785 2422.315 1784.235 ;
        RECT 2423.105 1784.135 2423.275 1784.235 ;
        RECT 2422.625 1784.035 2423.275 1784.135 ;
        RECT 2422.545 1783.865 2423.355 1784.035 ;
        RECT 2423.585 1783.785 2423.755 1784.115 ;
        RECT 2424.065 1783.785 2424.235 1784.235 ;
        RECT 2424.545 1783.785 2424.715 1784.115 ;
        RECT 2425.025 1784.035 2425.295 1784.235 ;
        RECT 2424.905 1783.825 2425.295 1784.035 ;
        RECT 2427.505 1783.895 2427.680 1785.155 ;
        RECT 2428.030 1784.095 2428.200 1785.155 ;
        RECT 2428.030 1783.925 2428.260 1784.095 ;
        RECT 2427.505 1783.695 2427.675 1783.895 ;
        RECT 2422.625 1783.615 2422.795 1783.655 ;
        RECT 2422.265 1783.445 2422.795 1783.615 ;
        RECT 2414.170 1783.035 2415.090 1783.205 ;
        RECT 2415.605 1783.035 2416.075 1783.205 ;
        RECT 2417.605 1783.045 2417.775 1783.395 ;
        RECT 2419.505 1783.045 2419.675 1783.395 ;
        RECT 2420.905 1783.375 2421.075 1783.395 ;
        RECT 2420.905 1783.345 2421.115 1783.375 ;
        RECT 2420.805 1783.125 2421.115 1783.345 ;
        RECT 2420.945 1783.045 2421.115 1783.125 ;
        RECT 2421.905 1783.275 2422.075 1783.395 ;
        RECT 2421.905 1783.105 2423.145 1783.275 ;
        RECT 2423.825 1783.045 2423.995 1783.395 ;
        RECT 2424.785 1783.045 2424.955 1783.395 ;
        RECT 2427.505 1783.365 2427.915 1783.695 ;
        RECT 2414.170 1782.885 2414.400 1783.035 ;
        RECT 2427.505 1782.855 2427.675 1783.365 ;
        RECT 2427.505 1782.525 2427.915 1782.855 ;
        RECT 2412.770 1782.145 2413.000 1782.315 ;
        RECT 2412.770 1781.865 2412.940 1782.145 ;
        RECT 2413.200 1781.865 2413.375 1782.375 ;
        RECT 2413.630 1781.865 2413.805 1782.415 ;
        RECT 2414.995 1781.865 2415.165 1782.375 ;
        RECT 2415.980 1781.865 2416.150 1782.375 ;
        RECT 2427.505 1782.355 2427.675 1782.525 ;
        RECT 2427.505 1781.865 2427.680 1782.355 ;
        RECT 2428.090 1782.315 2428.260 1783.925 ;
        RECT 2428.460 1783.895 2428.635 1785.155 ;
        RECT 2428.890 1784.015 2429.065 1785.155 ;
        RECT 2428.460 1782.945 2428.630 1783.895 ;
        RECT 2428.890 1782.415 2429.060 1784.015 ;
        RECT 2430.250 1784.010 2430.425 1785.155 ;
        RECT 2431.235 1784.010 2431.410 1785.155 ;
        RECT 2432.865 1784.435 2433.035 1784.795 ;
        RECT 2433.805 1784.435 2433.975 1784.795 ;
        RECT 2434.285 1784.345 2434.455 1784.765 ;
        RECT 2434.645 1784.515 2434.935 1785.075 ;
        RECT 2435.725 1784.775 2435.895 1785.105 ;
        RECT 2436.205 1784.685 2436.375 1785.075 ;
        RECT 2438.100 1784.775 2438.275 1785.105 ;
        RECT 2440.045 1784.905 2440.555 1785.075 ;
        RECT 2438.625 1784.685 2438.805 1784.795 ;
        RECT 2440.385 1784.765 2440.555 1784.905 ;
        RECT 2436.095 1784.515 2436.430 1784.685 ;
        RECT 2436.925 1784.515 2437.415 1784.685 ;
        RECT 2438.625 1784.515 2439.975 1784.685 ;
        RECT 2440.385 1784.515 2440.670 1784.765 ;
        RECT 2434.765 1784.435 2434.935 1784.515 ;
        RECT 2429.880 1783.205 2430.050 1783.895 ;
        RECT 2430.250 1783.795 2430.420 1784.010 ;
        RECT 2430.865 1783.795 2431.035 1783.895 ;
        RECT 2430.250 1783.625 2431.035 1783.795 ;
        RECT 2430.250 1783.575 2430.420 1783.625 ;
        RECT 2430.865 1783.205 2431.035 1783.625 ;
        RECT 2431.235 1783.575 2431.405 1784.010 ;
        RECT 2433.565 1783.785 2433.735 1784.235 ;
        RECT 2434.045 1783.785 2434.215 1784.115 ;
        RECT 2435.005 1783.785 2435.175 1784.115 ;
        RECT 2435.485 1783.785 2435.655 1784.515 ;
        RECT 2436.925 1784.345 2437.095 1784.515 ;
        RECT 2438.625 1784.435 2438.805 1784.515 ;
        RECT 2439.805 1784.345 2439.975 1784.515 ;
        RECT 2440.495 1784.435 2440.670 1784.515 ;
        RECT 2435.965 1783.785 2436.135 1784.235 ;
        RECT 2436.445 1783.785 2436.615 1784.115 ;
        RECT 2436.925 1783.785 2437.095 1784.115 ;
        RECT 2437.405 1783.785 2437.575 1784.235 ;
        RECT 2438.365 1784.135 2438.535 1784.235 ;
        RECT 2437.885 1784.035 2438.535 1784.135 ;
        RECT 2437.805 1783.865 2438.615 1784.035 ;
        RECT 2438.845 1783.785 2439.015 1784.115 ;
        RECT 2439.325 1783.785 2439.495 1784.235 ;
        RECT 2439.805 1783.785 2439.975 1784.115 ;
        RECT 2440.285 1784.035 2440.555 1784.235 ;
        RECT 2440.165 1783.825 2440.555 1784.035 ;
        RECT 2442.765 1783.895 2442.940 1785.155 ;
        RECT 2443.290 1784.095 2443.460 1785.155 ;
        RECT 2443.290 1783.925 2443.520 1784.095 ;
        RECT 2442.765 1783.695 2442.935 1783.895 ;
        RECT 2437.885 1783.615 2438.055 1783.655 ;
        RECT 2437.525 1783.445 2438.055 1783.615 ;
        RECT 2429.430 1783.035 2430.350 1783.205 ;
        RECT 2430.865 1783.035 2431.335 1783.205 ;
        RECT 2432.865 1783.045 2433.035 1783.395 ;
        RECT 2434.765 1783.045 2434.935 1783.395 ;
        RECT 2436.165 1783.375 2436.335 1783.395 ;
        RECT 2436.165 1783.345 2436.375 1783.375 ;
        RECT 2436.065 1783.125 2436.375 1783.345 ;
        RECT 2436.205 1783.045 2436.375 1783.125 ;
        RECT 2437.165 1783.275 2437.335 1783.395 ;
        RECT 2437.165 1783.105 2438.405 1783.275 ;
        RECT 2439.085 1783.045 2439.255 1783.395 ;
        RECT 2440.045 1783.045 2440.215 1783.395 ;
        RECT 2442.765 1783.365 2443.175 1783.695 ;
        RECT 2429.430 1782.885 2429.660 1783.035 ;
        RECT 2442.765 1782.855 2442.935 1783.365 ;
        RECT 2442.765 1782.525 2443.175 1782.855 ;
        RECT 2428.030 1782.145 2428.260 1782.315 ;
        RECT 2428.030 1781.865 2428.200 1782.145 ;
        RECT 2428.460 1781.865 2428.635 1782.375 ;
        RECT 2428.890 1781.865 2429.065 1782.415 ;
        RECT 2430.255 1781.865 2430.425 1782.375 ;
        RECT 2431.240 1781.865 2431.410 1782.375 ;
        RECT 2442.765 1782.355 2442.935 1782.525 ;
        RECT 2442.765 1781.865 2442.940 1782.355 ;
        RECT 2443.350 1782.315 2443.520 1783.925 ;
        RECT 2443.720 1783.895 2443.895 1785.155 ;
        RECT 2444.150 1784.015 2444.325 1785.155 ;
        RECT 2443.720 1782.945 2443.890 1783.895 ;
        RECT 2444.150 1782.415 2444.320 1784.015 ;
        RECT 2445.510 1784.010 2445.685 1785.155 ;
        RECT 2446.495 1784.010 2446.670 1785.155 ;
        RECT 2696.985 1785.135 2698.215 1785.305 ;
        RECT 2696.985 1784.325 2697.325 1785.135 ;
        RECT 2697.495 1784.570 2698.245 1784.760 ;
        RECT 2445.140 1783.205 2445.310 1783.895 ;
        RECT 2445.510 1783.795 2445.680 1784.010 ;
        RECT 2446.125 1783.795 2446.295 1783.895 ;
        RECT 2445.510 1783.625 2446.295 1783.795 ;
        RECT 2445.510 1783.575 2445.680 1783.625 ;
        RECT 2446.125 1783.205 2446.295 1783.625 ;
        RECT 2446.495 1783.575 2446.665 1784.010 ;
        RECT 2696.985 1783.915 2697.500 1784.325 ;
        RECT 2698.075 1783.905 2698.245 1784.570 ;
        RECT 2698.415 1784.585 2698.605 1785.945 ;
        RECT 2698.775 1785.095 2699.050 1785.945 ;
        RECT 2699.240 1785.580 2699.770 1785.945 ;
        RECT 2699.595 1785.545 2699.770 1785.580 ;
        RECT 2698.775 1784.925 2699.055 1785.095 ;
        RECT 2698.775 1784.785 2699.050 1784.925 ;
        RECT 2699.255 1784.585 2699.425 1785.385 ;
        RECT 2698.415 1784.415 2699.425 1784.585 ;
        RECT 2699.595 1785.375 2700.525 1785.545 ;
        RECT 2700.695 1785.375 2700.950 1785.945 ;
        RECT 2699.595 1784.245 2699.765 1785.375 ;
        RECT 2700.355 1785.205 2700.525 1785.375 ;
        RECT 2698.640 1784.075 2699.765 1784.245 ;
        RECT 2699.935 1784.875 2700.130 1785.205 ;
        RECT 2700.355 1784.875 2700.610 1785.205 ;
        RECT 2699.935 1783.905 2700.105 1784.875 ;
        RECT 2700.780 1784.705 2700.950 1785.375 ;
        RECT 2698.075 1783.735 2700.105 1783.905 ;
        RECT 2700.615 1783.735 2700.950 1784.705 ;
        RECT 2444.690 1783.035 2445.610 1783.205 ;
        RECT 2446.125 1783.035 2446.595 1783.205 ;
        RECT 2444.690 1782.885 2444.920 1783.035 ;
        RECT 2697.075 1782.465 2697.245 1783.225 ;
        RECT 2443.290 1782.145 2443.520 1782.315 ;
        RECT 2443.290 1781.865 2443.460 1782.145 ;
        RECT 2443.720 1781.865 2443.895 1782.375 ;
        RECT 2444.150 1781.865 2444.325 1782.415 ;
        RECT 2445.515 1781.865 2445.685 1782.375 ;
        RECT 2446.500 1781.865 2446.670 1782.375 ;
        RECT 2697.075 1782.295 2697.740 1782.465 ;
        RECT 2697.925 1782.320 2698.195 1783.225 ;
        RECT 2697.570 1782.150 2697.740 1782.295 ;
        RECT 2522.640 1779.885 2523.160 1781.370 ;
        RECT 2523.330 1780.545 2523.850 1782.095 ;
        RECT 2697.005 1781.745 2697.335 1782.115 ;
        RECT 2697.570 1781.820 2697.855 1782.150 ;
        RECT 2697.570 1781.565 2697.740 1781.820 ;
        RECT 2697.075 1781.395 2697.740 1781.565 ;
        RECT 2698.025 1781.520 2698.195 1782.320 ;
        RECT 2697.075 1781.015 2697.245 1781.395 ;
        RECT 2697.935 1781.015 2698.195 1781.520 ;
        RECT 2697.075 1777.025 2697.245 1777.785 ;
        RECT 2697.075 1776.855 2697.740 1777.025 ;
        RECT 2697.925 1776.880 2698.195 1777.785 ;
        RECT 2697.570 1776.710 2697.740 1776.855 ;
        RECT 2697.005 1776.305 2697.335 1776.675 ;
        RECT 2697.570 1776.380 2697.855 1776.710 ;
        RECT 2697.570 1776.125 2697.740 1776.380 ;
        RECT 2697.075 1775.955 2697.740 1776.125 ;
        RECT 2698.025 1776.080 2698.195 1776.880 ;
        RECT 2697.075 1775.575 2697.245 1775.955 ;
        RECT 2697.935 1775.575 2698.195 1776.080 ;
        RECT 2697.075 1771.585 2697.245 1772.345 ;
        RECT 2697.075 1771.415 2697.740 1771.585 ;
        RECT 2697.925 1771.440 2698.195 1772.345 ;
        RECT 2697.570 1771.270 2697.740 1771.415 ;
        RECT 2697.005 1770.865 2697.335 1771.235 ;
        RECT 2697.570 1770.940 2697.855 1771.270 ;
        RECT 2697.570 1770.685 2697.740 1770.940 ;
        RECT 2522.640 1768.415 2523.160 1769.900 ;
        RECT 2523.330 1769.075 2523.850 1770.625 ;
        RECT 2697.075 1770.515 2697.740 1770.685 ;
        RECT 2698.025 1770.640 2698.195 1771.440 ;
        RECT 2698.455 1771.585 2698.625 1772.345 ;
        RECT 2698.455 1771.415 2699.120 1771.585 ;
        RECT 2699.305 1771.440 2699.575 1772.345 ;
        RECT 2698.950 1771.270 2699.120 1771.415 ;
        RECT 2698.385 1770.865 2698.715 1771.235 ;
        RECT 2698.950 1770.940 2699.235 1771.270 ;
        RECT 2698.950 1770.685 2699.120 1770.940 ;
        RECT 2697.075 1770.135 2697.245 1770.515 ;
        RECT 2697.935 1770.135 2698.195 1770.640 ;
        RECT 2698.455 1770.515 2699.120 1770.685 ;
        RECT 2699.405 1770.640 2699.575 1771.440 ;
        RECT 2698.455 1770.135 2698.625 1770.515 ;
        RECT 2699.315 1770.135 2699.575 1770.640 ;
        RECT 2359.015 1710.095 2359.190 1710.585 ;
        RECT 2359.540 1710.305 2359.710 1710.585 ;
        RECT 2359.540 1710.135 2359.770 1710.305 ;
        RECT 2359.015 1709.925 2359.185 1710.095 ;
        RECT 2359.015 1709.595 2359.425 1709.925 ;
        RECT 2359.015 1709.085 2359.185 1709.595 ;
        RECT 2359.015 1708.755 2359.425 1709.085 ;
        RECT 2359.015 1708.555 2359.185 1708.755 ;
        RECT 2359.015 1707.295 2359.190 1708.555 ;
        RECT 2359.600 1708.525 2359.770 1710.135 ;
        RECT 2359.970 1710.075 2360.145 1710.585 ;
        RECT 2362.245 1710.095 2362.420 1710.585 ;
        RECT 2362.245 1709.925 2362.415 1710.095 ;
        RECT 2363.200 1710.075 2363.375 1710.585 ;
        RECT 2363.630 1710.035 2363.805 1710.585 ;
        RECT 2373.470 1710.100 2373.645 1710.590 ;
        RECT 2373.995 1710.310 2374.165 1710.590 ;
        RECT 2373.995 1710.140 2374.225 1710.310 ;
        RECT 2362.245 1709.595 2362.655 1709.925 ;
        RECT 2359.540 1708.355 2359.770 1708.525 ;
        RECT 2359.970 1708.555 2360.140 1709.505 ;
        RECT 2362.245 1709.085 2362.415 1709.595 ;
        RECT 2362.245 1708.755 2362.655 1709.085 ;
        RECT 2362.245 1708.555 2362.415 1708.755 ;
        RECT 2363.200 1708.555 2363.370 1709.505 ;
        RECT 2359.540 1707.295 2359.710 1708.355 ;
        RECT 2359.970 1707.295 2360.145 1708.555 ;
        RECT 2362.245 1707.295 2362.420 1708.555 ;
        RECT 2363.200 1707.295 2363.375 1708.555 ;
        RECT 2363.630 1708.435 2363.800 1710.035 ;
        RECT 2373.470 1709.930 2373.640 1710.100 ;
        RECT 2373.470 1709.600 2373.880 1709.930 ;
        RECT 2373.470 1709.090 2373.640 1709.600 ;
        RECT 2373.470 1708.760 2373.880 1709.090 ;
        RECT 2373.470 1708.560 2373.640 1708.760 ;
        RECT 2363.630 1707.295 2363.805 1708.435 ;
        RECT 2365.420 1707.895 2365.980 1708.185 ;
        RECT 2367.020 1708.055 2367.280 1708.085 ;
        RECT 2365.420 1706.525 2365.670 1707.895 ;
        RECT 2367.020 1707.725 2367.350 1708.055 ;
        RECT 2368.730 1707.935 2370.040 1708.185 ;
        RECT 2368.730 1707.785 2368.910 1707.935 ;
        RECT 2365.960 1707.535 2367.350 1707.725 ;
        RECT 2368.180 1707.615 2368.910 1707.785 ;
        RECT 2365.960 1707.445 2366.130 1707.535 ;
        RECT 2365.840 1707.115 2366.130 1707.445 ;
        RECT 2366.860 1707.115 2367.540 1707.365 ;
        RECT 2365.960 1706.865 2366.130 1707.115 ;
        RECT 2365.960 1706.695 2366.905 1706.865 ;
        RECT 2367.270 1706.755 2367.540 1707.115 ;
        RECT 2368.180 1706.945 2368.350 1707.615 ;
        RECT 2369.160 1707.365 2369.370 1707.765 ;
        RECT 2369.020 1707.165 2369.370 1707.365 ;
        RECT 2369.620 1707.365 2369.870 1707.765 ;
        RECT 2369.620 1707.165 2370.090 1707.365 ;
        RECT 2370.280 1707.165 2370.730 1707.675 ;
        RECT 2373.470 1707.300 2373.645 1708.560 ;
        RECT 2374.055 1708.530 2374.225 1710.140 ;
        RECT 2374.425 1710.080 2374.600 1710.590 ;
        RECT 2374.855 1710.040 2375.030 1710.590 ;
        RECT 2376.220 1710.080 2376.390 1710.590 ;
        RECT 2377.210 1710.080 2377.380 1710.590 ;
        RECT 2378.830 1710.095 2379.005 1710.585 ;
        RECT 2373.995 1708.360 2374.225 1708.530 ;
        RECT 2374.425 1708.560 2374.595 1709.510 ;
        RECT 2373.995 1707.300 2374.165 1708.360 ;
        RECT 2374.425 1707.300 2374.600 1708.560 ;
        RECT 2374.855 1708.440 2375.025 1710.040 ;
        RECT 2378.830 1709.925 2379.000 1710.095 ;
        RECT 2379.785 1710.075 2379.960 1710.585 ;
        RECT 2380.215 1710.035 2380.390 1710.585 ;
        RECT 2390.055 1710.100 2390.230 1710.590 ;
        RECT 2390.580 1710.310 2390.750 1710.590 ;
        RECT 2390.580 1710.140 2390.810 1710.310 ;
        RECT 2378.830 1709.595 2379.240 1709.925 ;
        RECT 2375.395 1709.420 2375.625 1709.570 ;
        RECT 2375.395 1709.250 2376.315 1709.420 ;
        RECT 2376.835 1709.250 2377.305 1709.420 ;
        RECT 2375.845 1708.560 2376.015 1709.250 ;
        RECT 2376.215 1708.770 2376.385 1708.880 ;
        RECT 2376.835 1708.770 2377.005 1709.250 ;
        RECT 2378.830 1709.085 2379.000 1709.595 ;
        RECT 2376.215 1708.600 2377.005 1708.770 ;
        RECT 2374.855 1707.300 2375.030 1708.440 ;
        RECT 2376.215 1707.300 2376.390 1708.600 ;
        RECT 2376.835 1708.560 2377.005 1708.600 ;
        RECT 2377.205 1708.445 2377.375 1708.880 ;
        RECT 2378.830 1708.755 2379.240 1709.085 ;
        RECT 2378.830 1708.555 2379.000 1708.755 ;
        RECT 2379.785 1708.555 2379.955 1709.505 ;
        RECT 2377.205 1707.300 2377.380 1708.445 ;
        RECT 2378.830 1707.295 2379.005 1708.555 ;
        RECT 2379.785 1707.295 2379.960 1708.555 ;
        RECT 2380.215 1708.435 2380.385 1710.035 ;
        RECT 2390.055 1709.930 2390.225 1710.100 ;
        RECT 2390.055 1709.600 2390.465 1709.930 ;
        RECT 2390.055 1709.090 2390.225 1709.600 ;
        RECT 2390.055 1708.760 2390.465 1709.090 ;
        RECT 2390.055 1708.560 2390.225 1708.760 ;
        RECT 2380.215 1707.295 2380.390 1708.435 ;
        RECT 2382.005 1707.895 2382.565 1708.185 ;
        RECT 2383.605 1708.055 2383.865 1708.085 ;
        RECT 2369.020 1706.945 2370.760 1706.995 ;
        RECT 2368.180 1706.815 2370.760 1706.945 ;
        RECT 2368.180 1706.775 2369.240 1706.815 ;
        RECT 2365.420 1705.975 2365.880 1706.525 ;
        RECT 2366.600 1705.975 2366.905 1706.695 ;
        RECT 2369.380 1706.605 2370.260 1706.645 ;
        RECT 2368.730 1706.405 2370.260 1706.605 ;
        RECT 2368.730 1706.275 2368.900 1706.405 ;
        RECT 2369.650 1706.355 2370.260 1706.405 ;
        RECT 2370.030 1706.315 2370.260 1706.355 ;
        RECT 2370.430 1706.315 2370.760 1706.815 ;
        RECT 2382.005 1706.525 2382.255 1707.895 ;
        RECT 2383.605 1707.725 2383.935 1708.055 ;
        RECT 2385.315 1707.935 2386.625 1708.185 ;
        RECT 2385.315 1707.785 2385.495 1707.935 ;
        RECT 2382.545 1707.535 2383.935 1707.725 ;
        RECT 2384.765 1707.615 2385.495 1707.785 ;
        RECT 2382.545 1707.445 2382.715 1707.535 ;
        RECT 2382.425 1707.115 2382.715 1707.445 ;
        RECT 2383.445 1707.115 2384.125 1707.365 ;
        RECT 2382.545 1706.865 2382.715 1707.115 ;
        RECT 2382.545 1706.695 2383.490 1706.865 ;
        RECT 2383.855 1706.755 2384.125 1707.115 ;
        RECT 2384.765 1706.945 2384.935 1707.615 ;
        RECT 2385.745 1707.365 2385.955 1707.765 ;
        RECT 2385.605 1707.165 2385.955 1707.365 ;
        RECT 2386.205 1707.365 2386.455 1707.765 ;
        RECT 2386.205 1707.165 2386.675 1707.365 ;
        RECT 2386.865 1707.165 2387.315 1707.675 ;
        RECT 2390.055 1707.300 2390.230 1708.560 ;
        RECT 2390.640 1708.530 2390.810 1710.140 ;
        RECT 2391.010 1710.080 2391.185 1710.590 ;
        RECT 2391.440 1710.040 2391.615 1710.590 ;
        RECT 2392.805 1710.080 2392.975 1710.590 ;
        RECT 2393.795 1710.080 2393.965 1710.590 ;
        RECT 2395.415 1710.100 2395.590 1710.590 ;
        RECT 2390.580 1708.360 2390.810 1708.530 ;
        RECT 2391.010 1708.560 2391.180 1709.510 ;
        RECT 2390.580 1707.300 2390.750 1708.360 ;
        RECT 2391.010 1707.300 2391.185 1708.560 ;
        RECT 2391.440 1708.440 2391.610 1710.040 ;
        RECT 2395.415 1709.930 2395.585 1710.100 ;
        RECT 2396.370 1710.080 2396.545 1710.590 ;
        RECT 2396.800 1710.040 2396.975 1710.590 ;
        RECT 2406.640 1710.105 2406.815 1710.595 ;
        RECT 2407.165 1710.315 2407.335 1710.595 ;
        RECT 2407.165 1710.145 2407.395 1710.315 ;
        RECT 2395.415 1709.600 2395.825 1709.930 ;
        RECT 2391.980 1709.420 2392.210 1709.570 ;
        RECT 2391.980 1709.250 2392.900 1709.420 ;
        RECT 2393.420 1709.250 2393.890 1709.420 ;
        RECT 2392.430 1708.560 2392.600 1709.250 ;
        RECT 2392.800 1708.770 2392.970 1708.880 ;
        RECT 2393.420 1708.770 2393.590 1709.250 ;
        RECT 2395.415 1709.090 2395.585 1709.600 ;
        RECT 2392.800 1708.600 2393.590 1708.770 ;
        RECT 2391.440 1707.300 2391.615 1708.440 ;
        RECT 2392.800 1707.300 2392.975 1708.600 ;
        RECT 2393.420 1708.560 2393.590 1708.600 ;
        RECT 2393.790 1708.445 2393.960 1708.880 ;
        RECT 2395.415 1708.760 2395.825 1709.090 ;
        RECT 2395.415 1708.560 2395.585 1708.760 ;
        RECT 2396.370 1708.560 2396.540 1709.510 ;
        RECT 2393.790 1707.300 2393.965 1708.445 ;
        RECT 2395.415 1707.300 2395.590 1708.560 ;
        RECT 2396.370 1707.300 2396.545 1708.560 ;
        RECT 2396.800 1708.440 2396.970 1710.040 ;
        RECT 2406.640 1709.935 2406.810 1710.105 ;
        RECT 2406.640 1709.605 2407.050 1709.935 ;
        RECT 2406.640 1709.095 2406.810 1709.605 ;
        RECT 2406.640 1708.765 2407.050 1709.095 ;
        RECT 2406.640 1708.565 2406.810 1708.765 ;
        RECT 2396.800 1707.300 2396.975 1708.440 ;
        RECT 2398.590 1707.900 2399.150 1708.190 ;
        RECT 2400.190 1708.060 2400.450 1708.090 ;
        RECT 2385.605 1706.945 2387.345 1706.995 ;
        RECT 2384.765 1706.815 2387.345 1706.945 ;
        RECT 2384.765 1706.775 2385.825 1706.815 ;
        RECT 2369.590 1706.145 2369.920 1706.185 ;
        RECT 2370.430 1706.145 2371.250 1706.315 ;
        RECT 2369.590 1705.975 2370.760 1706.145 ;
        RECT 2382.005 1705.975 2382.465 1706.525 ;
        RECT 2383.185 1705.975 2383.490 1706.695 ;
        RECT 2385.965 1706.605 2386.845 1706.645 ;
        RECT 2385.315 1706.405 2386.845 1706.605 ;
        RECT 2385.315 1706.275 2385.485 1706.405 ;
        RECT 2386.235 1706.355 2386.845 1706.405 ;
        RECT 2386.615 1706.315 2386.845 1706.355 ;
        RECT 2387.015 1706.315 2387.345 1706.815 ;
        RECT 2398.590 1706.530 2398.840 1707.900 ;
        RECT 2400.190 1707.730 2400.520 1708.060 ;
        RECT 2401.900 1707.940 2403.210 1708.190 ;
        RECT 2401.900 1707.790 2402.080 1707.940 ;
        RECT 2399.130 1707.540 2400.520 1707.730 ;
        RECT 2401.350 1707.620 2402.080 1707.790 ;
        RECT 2399.130 1707.450 2399.300 1707.540 ;
        RECT 2399.010 1707.120 2399.300 1707.450 ;
        RECT 2400.030 1707.120 2400.710 1707.370 ;
        RECT 2399.130 1706.870 2399.300 1707.120 ;
        RECT 2399.130 1706.700 2400.075 1706.870 ;
        RECT 2400.440 1706.760 2400.710 1707.120 ;
        RECT 2401.350 1706.950 2401.520 1707.620 ;
        RECT 2402.330 1707.370 2402.540 1707.770 ;
        RECT 2402.190 1707.170 2402.540 1707.370 ;
        RECT 2402.790 1707.370 2403.040 1707.770 ;
        RECT 2402.790 1707.170 2403.260 1707.370 ;
        RECT 2403.450 1707.170 2403.900 1707.680 ;
        RECT 2406.640 1707.305 2406.815 1708.565 ;
        RECT 2407.225 1708.535 2407.395 1710.145 ;
        RECT 2407.595 1710.085 2407.770 1710.595 ;
        RECT 2408.025 1710.045 2408.200 1710.595 ;
        RECT 2409.390 1710.085 2409.560 1710.595 ;
        RECT 2410.380 1710.085 2410.550 1710.595 ;
        RECT 2412.000 1710.105 2412.175 1710.595 ;
        RECT 2407.165 1708.365 2407.395 1708.535 ;
        RECT 2407.595 1708.565 2407.765 1709.515 ;
        RECT 2407.165 1707.305 2407.335 1708.365 ;
        RECT 2407.595 1707.305 2407.770 1708.565 ;
        RECT 2408.025 1708.445 2408.195 1710.045 ;
        RECT 2412.000 1709.935 2412.170 1710.105 ;
        RECT 2412.955 1710.085 2413.130 1710.595 ;
        RECT 2413.385 1710.045 2413.560 1710.595 ;
        RECT 2423.225 1710.110 2423.400 1710.600 ;
        RECT 2423.750 1710.320 2423.920 1710.600 ;
        RECT 2423.750 1710.150 2423.980 1710.320 ;
        RECT 2412.000 1709.605 2412.410 1709.935 ;
        RECT 2408.565 1709.425 2408.795 1709.575 ;
        RECT 2408.565 1709.255 2409.485 1709.425 ;
        RECT 2410.005 1709.255 2410.475 1709.425 ;
        RECT 2409.015 1708.565 2409.185 1709.255 ;
        RECT 2409.385 1708.775 2409.555 1708.885 ;
        RECT 2410.005 1708.775 2410.175 1709.255 ;
        RECT 2412.000 1709.095 2412.170 1709.605 ;
        RECT 2409.385 1708.605 2410.175 1708.775 ;
        RECT 2408.025 1707.305 2408.200 1708.445 ;
        RECT 2409.385 1707.305 2409.560 1708.605 ;
        RECT 2410.005 1708.565 2410.175 1708.605 ;
        RECT 2410.375 1708.450 2410.545 1708.885 ;
        RECT 2412.000 1708.765 2412.410 1709.095 ;
        RECT 2412.000 1708.565 2412.170 1708.765 ;
        RECT 2412.955 1708.565 2413.125 1709.515 ;
        RECT 2410.375 1707.305 2410.550 1708.450 ;
        RECT 2412.000 1707.305 2412.175 1708.565 ;
        RECT 2412.955 1707.305 2413.130 1708.565 ;
        RECT 2413.385 1708.445 2413.555 1710.045 ;
        RECT 2423.225 1709.940 2423.395 1710.110 ;
        RECT 2423.225 1709.610 2423.635 1709.940 ;
        RECT 2423.225 1709.100 2423.395 1709.610 ;
        RECT 2423.225 1708.770 2423.635 1709.100 ;
        RECT 2423.225 1708.570 2423.395 1708.770 ;
        RECT 2413.385 1707.305 2413.560 1708.445 ;
        RECT 2415.175 1707.905 2415.735 1708.195 ;
        RECT 2416.775 1708.065 2417.035 1708.095 ;
        RECT 2402.190 1706.950 2403.930 1707.000 ;
        RECT 2401.350 1706.820 2403.930 1706.950 ;
        RECT 2401.350 1706.780 2402.410 1706.820 ;
        RECT 2386.175 1706.145 2386.505 1706.185 ;
        RECT 2387.015 1706.145 2387.835 1706.315 ;
        RECT 2386.175 1705.975 2387.345 1706.145 ;
        RECT 2398.590 1705.980 2399.050 1706.530 ;
        RECT 2399.770 1705.980 2400.075 1706.700 ;
        RECT 2402.550 1706.610 2403.430 1706.650 ;
        RECT 2401.900 1706.410 2403.430 1706.610 ;
        RECT 2401.900 1706.280 2402.070 1706.410 ;
        RECT 2402.820 1706.360 2403.430 1706.410 ;
        RECT 2403.200 1706.320 2403.430 1706.360 ;
        RECT 2403.600 1706.320 2403.930 1706.820 ;
        RECT 2415.175 1706.535 2415.425 1707.905 ;
        RECT 2416.775 1707.735 2417.105 1708.065 ;
        RECT 2418.485 1707.945 2419.795 1708.195 ;
        RECT 2418.485 1707.795 2418.665 1707.945 ;
        RECT 2415.715 1707.545 2417.105 1707.735 ;
        RECT 2417.935 1707.625 2418.665 1707.795 ;
        RECT 2415.715 1707.455 2415.885 1707.545 ;
        RECT 2415.595 1707.125 2415.885 1707.455 ;
        RECT 2416.615 1707.125 2417.295 1707.375 ;
        RECT 2415.715 1706.875 2415.885 1707.125 ;
        RECT 2415.715 1706.705 2416.660 1706.875 ;
        RECT 2417.025 1706.765 2417.295 1707.125 ;
        RECT 2417.935 1706.955 2418.105 1707.625 ;
        RECT 2418.915 1707.375 2419.125 1707.775 ;
        RECT 2418.775 1707.175 2419.125 1707.375 ;
        RECT 2419.375 1707.375 2419.625 1707.775 ;
        RECT 2419.375 1707.175 2419.845 1707.375 ;
        RECT 2420.035 1707.175 2420.485 1707.685 ;
        RECT 2423.225 1707.310 2423.400 1708.570 ;
        RECT 2423.810 1708.540 2423.980 1710.150 ;
        RECT 2424.180 1710.090 2424.355 1710.600 ;
        RECT 2424.610 1710.050 2424.785 1710.600 ;
        RECT 2425.975 1710.090 2426.145 1710.600 ;
        RECT 2426.965 1710.090 2427.135 1710.600 ;
        RECT 2428.580 1710.105 2428.755 1710.595 ;
        RECT 2423.750 1708.370 2423.980 1708.540 ;
        RECT 2424.180 1708.570 2424.350 1709.520 ;
        RECT 2423.750 1707.310 2423.920 1708.370 ;
        RECT 2424.180 1707.310 2424.355 1708.570 ;
        RECT 2424.610 1708.450 2424.780 1710.050 ;
        RECT 2428.580 1709.935 2428.750 1710.105 ;
        RECT 2429.535 1710.085 2429.710 1710.595 ;
        RECT 2429.965 1710.045 2430.140 1710.595 ;
        RECT 2439.805 1710.110 2439.980 1710.600 ;
        RECT 2440.330 1710.320 2440.500 1710.600 ;
        RECT 2440.330 1710.150 2440.560 1710.320 ;
        RECT 2428.580 1709.605 2428.990 1709.935 ;
        RECT 2425.150 1709.430 2425.380 1709.580 ;
        RECT 2425.150 1709.260 2426.070 1709.430 ;
        RECT 2426.590 1709.260 2427.060 1709.430 ;
        RECT 2425.600 1708.570 2425.770 1709.260 ;
        RECT 2425.970 1708.780 2426.140 1708.890 ;
        RECT 2426.590 1708.780 2426.760 1709.260 ;
        RECT 2428.580 1709.095 2428.750 1709.605 ;
        RECT 2425.970 1708.610 2426.760 1708.780 ;
        RECT 2424.610 1707.310 2424.785 1708.450 ;
        RECT 2425.970 1707.310 2426.145 1708.610 ;
        RECT 2426.590 1708.570 2426.760 1708.610 ;
        RECT 2426.960 1708.455 2427.130 1708.890 ;
        RECT 2428.580 1708.765 2428.990 1709.095 ;
        RECT 2428.580 1708.565 2428.750 1708.765 ;
        RECT 2429.535 1708.565 2429.705 1709.515 ;
        RECT 2426.960 1707.310 2427.135 1708.455 ;
        RECT 2428.580 1707.305 2428.755 1708.565 ;
        RECT 2429.535 1707.305 2429.710 1708.565 ;
        RECT 2429.965 1708.445 2430.135 1710.045 ;
        RECT 2439.805 1709.940 2439.975 1710.110 ;
        RECT 2439.805 1709.610 2440.215 1709.940 ;
        RECT 2439.805 1709.100 2439.975 1709.610 ;
        RECT 2439.805 1708.770 2440.215 1709.100 ;
        RECT 2439.805 1708.570 2439.975 1708.770 ;
        RECT 2429.965 1707.305 2430.140 1708.445 ;
        RECT 2431.755 1707.905 2432.315 1708.195 ;
        RECT 2433.355 1708.065 2433.615 1708.095 ;
        RECT 2418.775 1706.955 2420.515 1707.005 ;
        RECT 2417.935 1706.825 2420.515 1706.955 ;
        RECT 2417.935 1706.785 2418.995 1706.825 ;
        RECT 2402.760 1706.150 2403.090 1706.190 ;
        RECT 2403.600 1706.150 2404.420 1706.320 ;
        RECT 2402.760 1705.980 2403.930 1706.150 ;
        RECT 2415.175 1705.985 2415.635 1706.535 ;
        RECT 2416.355 1705.985 2416.660 1706.705 ;
        RECT 2419.135 1706.615 2420.015 1706.655 ;
        RECT 2418.485 1706.415 2420.015 1706.615 ;
        RECT 2418.485 1706.285 2418.655 1706.415 ;
        RECT 2419.405 1706.365 2420.015 1706.415 ;
        RECT 2419.785 1706.325 2420.015 1706.365 ;
        RECT 2420.185 1706.325 2420.515 1706.825 ;
        RECT 2431.755 1706.535 2432.005 1707.905 ;
        RECT 2433.355 1707.735 2433.685 1708.065 ;
        RECT 2435.065 1707.945 2436.375 1708.195 ;
        RECT 2435.065 1707.795 2435.245 1707.945 ;
        RECT 2432.295 1707.545 2433.685 1707.735 ;
        RECT 2434.515 1707.625 2435.245 1707.795 ;
        RECT 2432.295 1707.455 2432.465 1707.545 ;
        RECT 2432.175 1707.125 2432.465 1707.455 ;
        RECT 2433.195 1707.125 2433.875 1707.375 ;
        RECT 2432.295 1706.875 2432.465 1707.125 ;
        RECT 2432.295 1706.705 2433.240 1706.875 ;
        RECT 2433.605 1706.765 2433.875 1707.125 ;
        RECT 2434.515 1706.955 2434.685 1707.625 ;
        RECT 2435.495 1707.375 2435.705 1707.775 ;
        RECT 2435.355 1707.175 2435.705 1707.375 ;
        RECT 2435.955 1707.375 2436.205 1707.775 ;
        RECT 2435.955 1707.175 2436.425 1707.375 ;
        RECT 2436.615 1707.175 2437.065 1707.685 ;
        RECT 2439.805 1707.310 2439.980 1708.570 ;
        RECT 2440.390 1708.540 2440.560 1710.150 ;
        RECT 2440.760 1710.090 2440.935 1710.600 ;
        RECT 2441.190 1710.050 2441.365 1710.600 ;
        RECT 2442.555 1710.090 2442.725 1710.600 ;
        RECT 2443.545 1710.090 2443.715 1710.600 ;
        RECT 2440.330 1708.370 2440.560 1708.540 ;
        RECT 2440.760 1708.570 2440.930 1709.520 ;
        RECT 2440.330 1707.310 2440.500 1708.370 ;
        RECT 2440.760 1707.310 2440.935 1708.570 ;
        RECT 2441.190 1708.450 2441.360 1710.050 ;
        RECT 2441.730 1709.430 2441.960 1709.580 ;
        RECT 2441.730 1709.260 2442.650 1709.430 ;
        RECT 2443.170 1709.260 2443.640 1709.430 ;
        RECT 2442.180 1708.570 2442.350 1709.260 ;
        RECT 2442.550 1708.780 2442.720 1708.890 ;
        RECT 2443.170 1708.780 2443.340 1709.260 ;
        RECT 2442.550 1708.610 2443.340 1708.780 ;
        RECT 2441.190 1707.310 2441.365 1708.450 ;
        RECT 2442.550 1707.310 2442.725 1708.610 ;
        RECT 2443.170 1708.570 2443.340 1708.610 ;
        RECT 2443.540 1708.455 2443.710 1708.890 ;
        RECT 2443.540 1707.310 2443.715 1708.455 ;
        RECT 2435.355 1706.955 2437.095 1707.005 ;
        RECT 2434.515 1706.825 2437.095 1706.955 ;
        RECT 2434.515 1706.785 2435.575 1706.825 ;
        RECT 2419.345 1706.155 2419.675 1706.195 ;
        RECT 2420.185 1706.155 2421.005 1706.325 ;
        RECT 2419.345 1705.985 2420.515 1706.155 ;
        RECT 2431.755 1705.985 2432.215 1706.535 ;
        RECT 2432.935 1705.985 2433.240 1706.705 ;
        RECT 2435.715 1706.615 2436.595 1706.655 ;
        RECT 2435.065 1706.415 2436.595 1706.615 ;
        RECT 2435.065 1706.285 2435.235 1706.415 ;
        RECT 2435.985 1706.365 2436.595 1706.415 ;
        RECT 2436.365 1706.325 2436.595 1706.365 ;
        RECT 2436.765 1706.325 2437.095 1706.825 ;
        RECT 2435.925 1706.155 2436.255 1706.195 ;
        RECT 2436.765 1706.155 2437.585 1706.325 ;
        RECT 2435.925 1705.985 2437.095 1706.155 ;
        RECT 2365.175 1705.125 2365.345 1705.465 ;
        RECT 2366.670 1705.125 2367.140 1705.465 ;
        RECT 2365.170 1705.065 2365.345 1705.125 ;
        RECT 2364.660 1704.075 2365.000 1704.955 ;
        RECT 2365.170 1704.245 2365.340 1705.065 ;
        RECT 2365.880 1704.595 2366.130 1704.965 ;
        RECT 2366.850 1704.595 2367.570 1704.895 ;
        RECT 2367.740 1704.765 2368.010 1705.465 ;
        RECT 2368.960 1705.125 2369.440 1705.465 ;
        RECT 2365.880 1704.425 2367.670 1704.595 ;
        RECT 2365.170 1703.995 2366.270 1704.245 ;
        RECT 2365.170 1703.905 2365.420 1703.995 ;
        RECT 2365.120 1703.485 2365.420 1703.905 ;
        RECT 2366.440 1703.575 2366.690 1704.425 ;
        RECT 2365.900 1703.305 2366.690 1703.575 ;
        RECT 2366.860 1703.725 2367.270 1704.245 ;
        RECT 2367.440 1703.995 2367.670 1704.425 ;
        RECT 2367.840 1703.735 2368.010 1704.765 ;
        RECT 2368.180 1704.365 2368.440 1704.815 ;
        RECT 2369.110 1704.635 2369.870 1704.885 ;
        RECT 2370.040 1704.765 2370.310 1705.465 ;
        RECT 2369.100 1704.605 2369.870 1704.635 ;
        RECT 2369.080 1704.595 2369.870 1704.605 ;
        RECT 2369.080 1704.575 2369.970 1704.595 ;
        RECT 2369.060 1704.565 2369.970 1704.575 ;
        RECT 2369.040 1704.555 2369.970 1704.565 ;
        RECT 2369.010 1704.545 2369.970 1704.555 ;
        RECT 2368.940 1704.515 2369.970 1704.545 ;
        RECT 2368.920 1704.485 2369.970 1704.515 ;
        RECT 2368.900 1704.455 2369.970 1704.485 ;
        RECT 2368.870 1704.425 2369.970 1704.455 ;
        RECT 2368.840 1704.395 2369.970 1704.425 ;
        RECT 2368.810 1704.385 2369.970 1704.395 ;
        RECT 2368.810 1704.375 2369.170 1704.385 ;
        RECT 2368.810 1704.365 2369.160 1704.375 ;
        RECT 2368.180 1704.355 2369.140 1704.365 ;
        RECT 2368.180 1704.345 2369.130 1704.355 ;
        RECT 2368.180 1704.325 2369.110 1704.345 ;
        RECT 2368.180 1704.315 2369.100 1704.325 ;
        RECT 2368.180 1704.195 2369.070 1704.315 ;
        RECT 2366.860 1703.305 2367.060 1703.725 ;
        RECT 2367.750 1703.265 2368.010 1703.735 ;
        RECT 2368.180 1703.635 2368.730 1704.025 ;
        RECT 2368.900 1703.465 2369.070 1704.195 ;
        RECT 2368.180 1703.295 2369.070 1703.465 ;
        RECT 2369.240 1703.795 2369.570 1704.215 ;
        RECT 2369.740 1703.995 2369.970 1704.385 ;
        RECT 2370.140 1704.275 2370.310 1704.765 ;
        RECT 2370.490 1704.665 2370.820 1705.455 ;
        RECT 2370.490 1704.495 2371.170 1704.665 ;
        RECT 2370.480 1704.275 2370.830 1704.325 ;
        RECT 2370.140 1704.105 2370.830 1704.275 ;
        RECT 2369.240 1703.305 2369.460 1703.795 ;
        RECT 2370.140 1703.735 2370.310 1704.105 ;
        RECT 2370.480 1704.075 2370.830 1704.105 ;
        RECT 2371.000 1703.895 2371.170 1704.495 ;
        RECT 2371.340 1704.075 2371.690 1704.325 ;
        RECT 2373.470 1703.900 2373.645 1705.160 ;
        RECT 2373.995 1704.100 2374.165 1705.160 ;
        RECT 2373.995 1703.930 2374.225 1704.100 ;
        RECT 2370.050 1703.265 2370.310 1703.735 ;
        RECT 2370.910 1703.265 2371.240 1703.895 ;
        RECT 2373.470 1703.700 2373.640 1703.900 ;
        RECT 2373.470 1703.370 2373.880 1703.700 ;
        RECT 2373.470 1702.860 2373.640 1703.370 ;
        RECT 2373.470 1702.530 2373.880 1702.860 ;
        RECT 2373.470 1702.360 2373.640 1702.530 ;
        RECT 2373.470 1701.870 2373.645 1702.360 ;
        RECT 2374.055 1702.320 2374.225 1703.930 ;
        RECT 2374.425 1703.900 2374.600 1705.160 ;
        RECT 2374.855 1704.020 2375.030 1705.160 ;
        RECT 2374.425 1702.950 2374.595 1703.900 ;
        RECT 2374.855 1702.420 2375.025 1704.020 ;
        RECT 2376.215 1704.015 2376.390 1705.160 ;
        RECT 2377.205 1704.015 2377.380 1705.160 ;
        RECT 2381.760 1705.125 2381.930 1705.465 ;
        RECT 2383.255 1705.125 2383.725 1705.465 ;
        RECT 2381.755 1705.065 2381.930 1705.125 ;
        RECT 2381.245 1704.075 2381.585 1704.955 ;
        RECT 2381.755 1704.245 2381.925 1705.065 ;
        RECT 2382.465 1704.595 2382.715 1704.965 ;
        RECT 2383.435 1704.595 2384.155 1704.895 ;
        RECT 2384.325 1704.765 2384.595 1705.465 ;
        RECT 2385.545 1705.125 2386.025 1705.465 ;
        RECT 2382.465 1704.425 2384.255 1704.595 ;
        RECT 2375.845 1703.210 2376.015 1703.900 ;
        RECT 2376.215 1703.800 2376.385 1704.015 ;
        RECT 2376.835 1703.800 2377.005 1703.900 ;
        RECT 2376.215 1703.630 2377.005 1703.800 ;
        RECT 2376.215 1703.580 2376.385 1703.630 ;
        RECT 2376.835 1703.210 2377.005 1703.630 ;
        RECT 2377.205 1703.580 2377.375 1704.015 ;
        RECT 2381.755 1703.995 2382.855 1704.245 ;
        RECT 2381.755 1703.905 2382.005 1703.995 ;
        RECT 2381.705 1703.485 2382.005 1703.905 ;
        RECT 2383.025 1703.575 2383.275 1704.425 ;
        RECT 2382.485 1703.305 2383.275 1703.575 ;
        RECT 2383.445 1703.725 2383.855 1704.245 ;
        RECT 2384.025 1703.995 2384.255 1704.425 ;
        RECT 2384.425 1703.735 2384.595 1704.765 ;
        RECT 2384.765 1704.365 2385.025 1704.815 ;
        RECT 2385.695 1704.635 2386.455 1704.885 ;
        RECT 2386.625 1704.765 2386.895 1705.465 ;
        RECT 2385.685 1704.605 2386.455 1704.635 ;
        RECT 2385.665 1704.595 2386.455 1704.605 ;
        RECT 2385.665 1704.575 2386.555 1704.595 ;
        RECT 2385.645 1704.565 2386.555 1704.575 ;
        RECT 2385.625 1704.555 2386.555 1704.565 ;
        RECT 2385.595 1704.545 2386.555 1704.555 ;
        RECT 2385.525 1704.515 2386.555 1704.545 ;
        RECT 2385.505 1704.485 2386.555 1704.515 ;
        RECT 2385.485 1704.455 2386.555 1704.485 ;
        RECT 2385.455 1704.425 2386.555 1704.455 ;
        RECT 2385.425 1704.395 2386.555 1704.425 ;
        RECT 2385.395 1704.385 2386.555 1704.395 ;
        RECT 2385.395 1704.375 2385.755 1704.385 ;
        RECT 2385.395 1704.365 2385.745 1704.375 ;
        RECT 2384.765 1704.355 2385.725 1704.365 ;
        RECT 2384.765 1704.345 2385.715 1704.355 ;
        RECT 2384.765 1704.325 2385.695 1704.345 ;
        RECT 2384.765 1704.315 2385.685 1704.325 ;
        RECT 2384.765 1704.195 2385.655 1704.315 ;
        RECT 2383.445 1703.305 2383.645 1703.725 ;
        RECT 2384.335 1703.265 2384.595 1703.735 ;
        RECT 2384.765 1703.635 2385.315 1704.025 ;
        RECT 2385.485 1703.465 2385.655 1704.195 ;
        RECT 2384.765 1703.295 2385.655 1703.465 ;
        RECT 2385.825 1703.795 2386.155 1704.215 ;
        RECT 2386.325 1703.995 2386.555 1704.385 ;
        RECT 2386.725 1704.275 2386.895 1704.765 ;
        RECT 2387.075 1704.665 2387.405 1705.455 ;
        RECT 2387.075 1704.495 2387.755 1704.665 ;
        RECT 2387.065 1704.275 2387.415 1704.325 ;
        RECT 2386.725 1704.105 2387.415 1704.275 ;
        RECT 2385.825 1703.305 2386.045 1703.795 ;
        RECT 2386.725 1703.735 2386.895 1704.105 ;
        RECT 2387.065 1704.075 2387.415 1704.105 ;
        RECT 2387.585 1703.895 2387.755 1704.495 ;
        RECT 2387.925 1704.075 2388.275 1704.325 ;
        RECT 2390.055 1703.900 2390.230 1705.160 ;
        RECT 2390.580 1704.100 2390.750 1705.160 ;
        RECT 2390.580 1703.930 2390.810 1704.100 ;
        RECT 2386.635 1703.265 2386.895 1703.735 ;
        RECT 2387.495 1703.265 2387.825 1703.895 ;
        RECT 2390.055 1703.700 2390.225 1703.900 ;
        RECT 2390.055 1703.370 2390.465 1703.700 ;
        RECT 2375.395 1703.040 2376.315 1703.210 ;
        RECT 2376.835 1703.040 2377.305 1703.210 ;
        RECT 2375.395 1702.890 2375.625 1703.040 ;
        RECT 2390.055 1702.860 2390.225 1703.370 ;
        RECT 2390.055 1702.530 2390.465 1702.860 ;
        RECT 2373.995 1702.150 2374.225 1702.320 ;
        RECT 2373.995 1701.870 2374.165 1702.150 ;
        RECT 2374.425 1701.870 2374.600 1702.380 ;
        RECT 2374.855 1701.870 2375.030 1702.420 ;
        RECT 2376.220 1701.870 2376.390 1702.380 ;
        RECT 2377.210 1701.785 2377.380 1702.380 ;
        RECT 2390.055 1702.360 2390.225 1702.530 ;
        RECT 2390.055 1701.870 2390.230 1702.360 ;
        RECT 2390.640 1702.320 2390.810 1703.930 ;
        RECT 2391.010 1703.900 2391.185 1705.160 ;
        RECT 2391.440 1704.020 2391.615 1705.160 ;
        RECT 2391.010 1702.950 2391.180 1703.900 ;
        RECT 2391.440 1702.420 2391.610 1704.020 ;
        RECT 2392.800 1704.015 2392.975 1705.160 ;
        RECT 2393.790 1704.015 2393.965 1705.160 ;
        RECT 2398.345 1705.130 2398.515 1705.470 ;
        RECT 2399.840 1705.130 2400.310 1705.470 ;
        RECT 2398.340 1705.070 2398.515 1705.130 ;
        RECT 2397.830 1704.080 2398.170 1704.960 ;
        RECT 2398.340 1704.250 2398.510 1705.070 ;
        RECT 2399.050 1704.600 2399.300 1704.970 ;
        RECT 2400.020 1704.600 2400.740 1704.900 ;
        RECT 2400.910 1704.770 2401.180 1705.470 ;
        RECT 2402.130 1705.130 2402.610 1705.470 ;
        RECT 2399.050 1704.430 2400.840 1704.600 ;
        RECT 2392.430 1703.210 2392.600 1703.900 ;
        RECT 2392.800 1703.800 2392.970 1704.015 ;
        RECT 2393.420 1703.800 2393.590 1703.900 ;
        RECT 2392.800 1703.630 2393.590 1703.800 ;
        RECT 2392.800 1703.580 2392.970 1703.630 ;
        RECT 2393.420 1703.210 2393.590 1703.630 ;
        RECT 2393.790 1703.580 2393.960 1704.015 ;
        RECT 2398.340 1704.000 2399.440 1704.250 ;
        RECT 2398.340 1703.910 2398.590 1704.000 ;
        RECT 2398.290 1703.490 2398.590 1703.910 ;
        RECT 2399.610 1703.580 2399.860 1704.430 ;
        RECT 2399.070 1703.310 2399.860 1703.580 ;
        RECT 2400.030 1703.730 2400.440 1704.250 ;
        RECT 2400.610 1704.000 2400.840 1704.430 ;
        RECT 2401.010 1703.740 2401.180 1704.770 ;
        RECT 2401.350 1704.370 2401.610 1704.820 ;
        RECT 2402.280 1704.640 2403.040 1704.890 ;
        RECT 2403.210 1704.770 2403.480 1705.470 ;
        RECT 2402.270 1704.610 2403.040 1704.640 ;
        RECT 2402.250 1704.600 2403.040 1704.610 ;
        RECT 2402.250 1704.580 2403.140 1704.600 ;
        RECT 2402.230 1704.570 2403.140 1704.580 ;
        RECT 2402.210 1704.560 2403.140 1704.570 ;
        RECT 2402.180 1704.550 2403.140 1704.560 ;
        RECT 2402.110 1704.520 2403.140 1704.550 ;
        RECT 2402.090 1704.490 2403.140 1704.520 ;
        RECT 2402.070 1704.460 2403.140 1704.490 ;
        RECT 2402.040 1704.430 2403.140 1704.460 ;
        RECT 2402.010 1704.400 2403.140 1704.430 ;
        RECT 2401.980 1704.390 2403.140 1704.400 ;
        RECT 2401.980 1704.380 2402.340 1704.390 ;
        RECT 2401.980 1704.370 2402.330 1704.380 ;
        RECT 2401.350 1704.360 2402.310 1704.370 ;
        RECT 2401.350 1704.350 2402.300 1704.360 ;
        RECT 2401.350 1704.330 2402.280 1704.350 ;
        RECT 2401.350 1704.320 2402.270 1704.330 ;
        RECT 2401.350 1704.200 2402.240 1704.320 ;
        RECT 2400.030 1703.310 2400.230 1703.730 ;
        RECT 2400.920 1703.270 2401.180 1703.740 ;
        RECT 2401.350 1703.640 2401.900 1704.030 ;
        RECT 2402.070 1703.470 2402.240 1704.200 ;
        RECT 2401.350 1703.300 2402.240 1703.470 ;
        RECT 2402.410 1703.800 2402.740 1704.220 ;
        RECT 2402.910 1704.000 2403.140 1704.390 ;
        RECT 2403.310 1704.280 2403.480 1704.770 ;
        RECT 2403.660 1704.670 2403.990 1705.460 ;
        RECT 2403.660 1704.500 2404.340 1704.670 ;
        RECT 2403.650 1704.280 2404.000 1704.330 ;
        RECT 2403.310 1704.110 2404.000 1704.280 ;
        RECT 2402.410 1703.310 2402.630 1703.800 ;
        RECT 2403.310 1703.740 2403.480 1704.110 ;
        RECT 2403.650 1704.080 2404.000 1704.110 ;
        RECT 2404.170 1703.900 2404.340 1704.500 ;
        RECT 2404.510 1704.080 2404.860 1704.330 ;
        RECT 2406.640 1703.905 2406.815 1705.165 ;
        RECT 2407.165 1704.105 2407.335 1705.165 ;
        RECT 2407.165 1703.935 2407.395 1704.105 ;
        RECT 2403.220 1703.270 2403.480 1703.740 ;
        RECT 2404.080 1703.270 2404.410 1703.900 ;
        RECT 2406.640 1703.705 2406.810 1703.905 ;
        RECT 2406.640 1703.375 2407.050 1703.705 ;
        RECT 2391.980 1703.040 2392.900 1703.210 ;
        RECT 2393.420 1703.040 2393.890 1703.210 ;
        RECT 2391.980 1702.890 2392.210 1703.040 ;
        RECT 2406.640 1702.865 2406.810 1703.375 ;
        RECT 2406.640 1702.535 2407.050 1702.865 ;
        RECT 2390.580 1702.150 2390.810 1702.320 ;
        RECT 2390.580 1701.870 2390.750 1702.150 ;
        RECT 2391.010 1701.870 2391.185 1702.380 ;
        RECT 2391.440 1701.870 2391.615 1702.420 ;
        RECT 2392.805 1701.870 2392.975 1702.380 ;
        RECT 2393.795 1701.785 2393.965 1702.380 ;
        RECT 2406.640 1702.365 2406.810 1702.535 ;
        RECT 2406.640 1701.875 2406.815 1702.365 ;
        RECT 2407.225 1702.325 2407.395 1703.935 ;
        RECT 2407.595 1703.905 2407.770 1705.165 ;
        RECT 2408.025 1704.025 2408.200 1705.165 ;
        RECT 2407.595 1702.955 2407.765 1703.905 ;
        RECT 2408.025 1702.425 2408.195 1704.025 ;
        RECT 2409.385 1704.020 2409.560 1705.165 ;
        RECT 2410.375 1704.020 2410.550 1705.165 ;
        RECT 2414.930 1705.135 2415.100 1705.475 ;
        RECT 2416.425 1705.135 2416.895 1705.475 ;
        RECT 2414.925 1705.075 2415.100 1705.135 ;
        RECT 2414.415 1704.085 2414.755 1704.965 ;
        RECT 2414.925 1704.255 2415.095 1705.075 ;
        RECT 2415.635 1704.605 2415.885 1704.975 ;
        RECT 2416.605 1704.605 2417.325 1704.905 ;
        RECT 2417.495 1704.775 2417.765 1705.475 ;
        RECT 2418.715 1705.135 2419.195 1705.475 ;
        RECT 2415.635 1704.435 2417.425 1704.605 ;
        RECT 2409.015 1703.215 2409.185 1703.905 ;
        RECT 2409.385 1703.805 2409.555 1704.020 ;
        RECT 2410.005 1703.805 2410.175 1703.905 ;
        RECT 2409.385 1703.635 2410.175 1703.805 ;
        RECT 2409.385 1703.585 2409.555 1703.635 ;
        RECT 2410.005 1703.215 2410.175 1703.635 ;
        RECT 2410.375 1703.585 2410.545 1704.020 ;
        RECT 2414.925 1704.005 2416.025 1704.255 ;
        RECT 2414.925 1703.915 2415.175 1704.005 ;
        RECT 2414.875 1703.495 2415.175 1703.915 ;
        RECT 2416.195 1703.585 2416.445 1704.435 ;
        RECT 2415.655 1703.315 2416.445 1703.585 ;
        RECT 2416.615 1703.735 2417.025 1704.255 ;
        RECT 2417.195 1704.005 2417.425 1704.435 ;
        RECT 2417.595 1703.745 2417.765 1704.775 ;
        RECT 2417.935 1704.375 2418.195 1704.825 ;
        RECT 2418.865 1704.645 2419.625 1704.895 ;
        RECT 2419.795 1704.775 2420.065 1705.475 ;
        RECT 2418.855 1704.615 2419.625 1704.645 ;
        RECT 2418.835 1704.605 2419.625 1704.615 ;
        RECT 2418.835 1704.585 2419.725 1704.605 ;
        RECT 2418.815 1704.575 2419.725 1704.585 ;
        RECT 2418.795 1704.565 2419.725 1704.575 ;
        RECT 2418.765 1704.555 2419.725 1704.565 ;
        RECT 2418.695 1704.525 2419.725 1704.555 ;
        RECT 2418.675 1704.495 2419.725 1704.525 ;
        RECT 2418.655 1704.465 2419.725 1704.495 ;
        RECT 2418.625 1704.435 2419.725 1704.465 ;
        RECT 2418.595 1704.405 2419.725 1704.435 ;
        RECT 2418.565 1704.395 2419.725 1704.405 ;
        RECT 2418.565 1704.385 2418.925 1704.395 ;
        RECT 2418.565 1704.375 2418.915 1704.385 ;
        RECT 2417.935 1704.365 2418.895 1704.375 ;
        RECT 2417.935 1704.355 2418.885 1704.365 ;
        RECT 2417.935 1704.335 2418.865 1704.355 ;
        RECT 2417.935 1704.325 2418.855 1704.335 ;
        RECT 2417.935 1704.205 2418.825 1704.325 ;
        RECT 2416.615 1703.315 2416.815 1703.735 ;
        RECT 2417.505 1703.275 2417.765 1703.745 ;
        RECT 2417.935 1703.645 2418.485 1704.035 ;
        RECT 2418.655 1703.475 2418.825 1704.205 ;
        RECT 2417.935 1703.305 2418.825 1703.475 ;
        RECT 2418.995 1703.805 2419.325 1704.225 ;
        RECT 2419.495 1704.005 2419.725 1704.395 ;
        RECT 2419.895 1704.285 2420.065 1704.775 ;
        RECT 2420.245 1704.675 2420.575 1705.465 ;
        RECT 2420.245 1704.505 2420.925 1704.675 ;
        RECT 2420.235 1704.285 2420.585 1704.335 ;
        RECT 2419.895 1704.115 2420.585 1704.285 ;
        RECT 2418.995 1703.315 2419.215 1703.805 ;
        RECT 2419.895 1703.745 2420.065 1704.115 ;
        RECT 2420.235 1704.085 2420.585 1704.115 ;
        RECT 2420.755 1703.905 2420.925 1704.505 ;
        RECT 2421.095 1704.085 2421.445 1704.335 ;
        RECT 2423.225 1703.910 2423.400 1705.170 ;
        RECT 2423.750 1704.110 2423.920 1705.170 ;
        RECT 2423.750 1703.940 2423.980 1704.110 ;
        RECT 2419.805 1703.275 2420.065 1703.745 ;
        RECT 2420.665 1703.275 2420.995 1703.905 ;
        RECT 2423.225 1703.710 2423.395 1703.910 ;
        RECT 2423.225 1703.380 2423.635 1703.710 ;
        RECT 2408.565 1703.045 2409.485 1703.215 ;
        RECT 2410.005 1703.045 2410.475 1703.215 ;
        RECT 2408.565 1702.895 2408.795 1703.045 ;
        RECT 2423.225 1702.870 2423.395 1703.380 ;
        RECT 2423.225 1702.540 2423.635 1702.870 ;
        RECT 2407.165 1702.155 2407.395 1702.325 ;
        RECT 2407.165 1701.875 2407.335 1702.155 ;
        RECT 2407.595 1701.875 2407.770 1702.385 ;
        RECT 2408.025 1701.875 2408.200 1702.425 ;
        RECT 2409.390 1701.875 2409.560 1702.385 ;
        RECT 2410.380 1701.875 2410.550 1702.385 ;
        RECT 2423.225 1702.370 2423.395 1702.540 ;
        RECT 2423.225 1701.880 2423.400 1702.370 ;
        RECT 2423.810 1702.330 2423.980 1703.940 ;
        RECT 2424.180 1703.910 2424.355 1705.170 ;
        RECT 2424.610 1704.030 2424.785 1705.170 ;
        RECT 2424.180 1702.960 2424.350 1703.910 ;
        RECT 2424.610 1702.430 2424.780 1704.030 ;
        RECT 2425.970 1704.025 2426.145 1705.170 ;
        RECT 2426.960 1704.025 2427.135 1705.170 ;
        RECT 2431.510 1705.135 2431.680 1705.475 ;
        RECT 2433.005 1705.135 2433.475 1705.475 ;
        RECT 2431.505 1705.075 2431.680 1705.135 ;
        RECT 2430.995 1704.085 2431.335 1704.965 ;
        RECT 2431.505 1704.255 2431.675 1705.075 ;
        RECT 2432.215 1704.605 2432.465 1704.975 ;
        RECT 2433.185 1704.605 2433.905 1704.905 ;
        RECT 2434.075 1704.775 2434.345 1705.475 ;
        RECT 2435.295 1705.135 2435.775 1705.475 ;
        RECT 2432.215 1704.435 2434.005 1704.605 ;
        RECT 2425.600 1703.220 2425.770 1703.910 ;
        RECT 2425.970 1703.810 2426.140 1704.025 ;
        RECT 2426.590 1703.810 2426.760 1703.910 ;
        RECT 2425.970 1703.640 2426.760 1703.810 ;
        RECT 2425.970 1703.590 2426.140 1703.640 ;
        RECT 2426.590 1703.220 2426.760 1703.640 ;
        RECT 2426.960 1703.590 2427.130 1704.025 ;
        RECT 2431.505 1704.005 2432.605 1704.255 ;
        RECT 2431.505 1703.915 2431.755 1704.005 ;
        RECT 2431.455 1703.495 2431.755 1703.915 ;
        RECT 2432.775 1703.585 2433.025 1704.435 ;
        RECT 2432.235 1703.315 2433.025 1703.585 ;
        RECT 2433.195 1703.735 2433.605 1704.255 ;
        RECT 2433.775 1704.005 2434.005 1704.435 ;
        RECT 2434.175 1703.745 2434.345 1704.775 ;
        RECT 2434.515 1704.375 2434.775 1704.825 ;
        RECT 2435.445 1704.645 2436.205 1704.895 ;
        RECT 2436.375 1704.775 2436.645 1705.475 ;
        RECT 2435.435 1704.615 2436.205 1704.645 ;
        RECT 2435.415 1704.605 2436.205 1704.615 ;
        RECT 2435.415 1704.585 2436.305 1704.605 ;
        RECT 2435.395 1704.575 2436.305 1704.585 ;
        RECT 2435.375 1704.565 2436.305 1704.575 ;
        RECT 2435.345 1704.555 2436.305 1704.565 ;
        RECT 2435.275 1704.525 2436.305 1704.555 ;
        RECT 2435.255 1704.495 2436.305 1704.525 ;
        RECT 2435.235 1704.465 2436.305 1704.495 ;
        RECT 2435.205 1704.435 2436.305 1704.465 ;
        RECT 2435.175 1704.405 2436.305 1704.435 ;
        RECT 2435.145 1704.395 2436.305 1704.405 ;
        RECT 2435.145 1704.385 2435.505 1704.395 ;
        RECT 2435.145 1704.375 2435.495 1704.385 ;
        RECT 2434.515 1704.365 2435.475 1704.375 ;
        RECT 2434.515 1704.355 2435.465 1704.365 ;
        RECT 2434.515 1704.335 2435.445 1704.355 ;
        RECT 2434.515 1704.325 2435.435 1704.335 ;
        RECT 2434.515 1704.205 2435.405 1704.325 ;
        RECT 2433.195 1703.315 2433.395 1703.735 ;
        RECT 2434.085 1703.275 2434.345 1703.745 ;
        RECT 2434.515 1703.645 2435.065 1704.035 ;
        RECT 2435.235 1703.475 2435.405 1704.205 ;
        RECT 2434.515 1703.305 2435.405 1703.475 ;
        RECT 2435.575 1703.805 2435.905 1704.225 ;
        RECT 2436.075 1704.005 2436.305 1704.395 ;
        RECT 2436.475 1704.285 2436.645 1704.775 ;
        RECT 2436.825 1704.675 2437.155 1705.465 ;
        RECT 2436.825 1704.505 2437.505 1704.675 ;
        RECT 2436.815 1704.285 2437.165 1704.335 ;
        RECT 2436.475 1704.115 2437.165 1704.285 ;
        RECT 2435.575 1703.315 2435.795 1703.805 ;
        RECT 2436.475 1703.745 2436.645 1704.115 ;
        RECT 2436.815 1704.085 2437.165 1704.115 ;
        RECT 2437.335 1703.905 2437.505 1704.505 ;
        RECT 2437.675 1704.085 2438.025 1704.335 ;
        RECT 2439.805 1703.910 2439.980 1705.170 ;
        RECT 2440.330 1704.110 2440.500 1705.170 ;
        RECT 2440.330 1703.940 2440.560 1704.110 ;
        RECT 2436.385 1703.275 2436.645 1703.745 ;
        RECT 2437.245 1703.275 2437.575 1703.905 ;
        RECT 2439.805 1703.710 2439.975 1703.910 ;
        RECT 2439.805 1703.380 2440.215 1703.710 ;
        RECT 2425.150 1703.050 2426.070 1703.220 ;
        RECT 2426.590 1703.050 2427.060 1703.220 ;
        RECT 2425.150 1702.900 2425.380 1703.050 ;
        RECT 2439.805 1702.870 2439.975 1703.380 ;
        RECT 2439.805 1702.540 2440.215 1702.870 ;
        RECT 2423.750 1702.160 2423.980 1702.330 ;
        RECT 2423.750 1701.880 2423.920 1702.160 ;
        RECT 2424.180 1701.880 2424.355 1702.390 ;
        RECT 2424.610 1701.880 2424.785 1702.430 ;
        RECT 2425.975 1701.880 2426.145 1702.390 ;
        RECT 2426.965 1701.880 2427.135 1702.390 ;
        RECT 2439.805 1702.370 2439.975 1702.540 ;
        RECT 2439.805 1701.880 2439.980 1702.370 ;
        RECT 2440.390 1702.330 2440.560 1703.940 ;
        RECT 2440.760 1703.910 2440.935 1705.170 ;
        RECT 2441.190 1704.030 2441.365 1705.170 ;
        RECT 2440.760 1702.960 2440.930 1703.910 ;
        RECT 2441.190 1702.430 2441.360 1704.030 ;
        RECT 2442.550 1704.025 2442.725 1705.170 ;
        RECT 2443.540 1704.025 2443.715 1705.170 ;
        RECT 2442.180 1703.220 2442.350 1703.910 ;
        RECT 2442.550 1703.810 2442.720 1704.025 ;
        RECT 2443.170 1703.810 2443.340 1703.910 ;
        RECT 2442.550 1703.640 2443.340 1703.810 ;
        RECT 2442.550 1703.590 2442.720 1703.640 ;
        RECT 2443.170 1703.220 2443.340 1703.640 ;
        RECT 2443.540 1703.590 2443.710 1704.025 ;
        RECT 2441.730 1703.050 2442.650 1703.220 ;
        RECT 2443.170 1703.050 2443.640 1703.220 ;
        RECT 2441.730 1702.900 2441.960 1703.050 ;
        RECT 2440.330 1702.160 2440.560 1702.330 ;
        RECT 2440.330 1701.880 2440.500 1702.160 ;
        RECT 2440.760 1701.880 2440.935 1702.390 ;
        RECT 2441.190 1701.880 2441.365 1702.430 ;
        RECT 2442.555 1701.880 2442.725 1702.390 ;
        RECT 2443.545 1701.880 2443.715 1702.390 ;
        RECT 2696.985 1676.335 2697.245 1676.665 ;
        RECT 2696.985 1675.425 2697.155 1676.335 ;
        RECT 2697.940 1676.265 2698.145 1676.665 ;
        RECT 2697.940 1676.095 2698.625 1676.265 ;
        RECT 2697.865 1675.425 2698.115 1675.925 ;
        RECT 2696.985 1675.255 2698.115 1675.425 ;
        RECT 2696.985 1674.485 2697.255 1675.255 ;
        RECT 2698.285 1675.065 2698.625 1676.095 ;
        RECT 2697.960 1674.890 2698.625 1675.065 ;
        RECT 2698.825 1676.160 2699.085 1676.665 ;
        RECT 2699.775 1676.285 2699.945 1676.665 ;
        RECT 2698.825 1675.360 2698.995 1676.160 ;
        RECT 2699.280 1676.115 2699.945 1676.285 ;
        RECT 2700.205 1676.160 2700.465 1676.665 ;
        RECT 2701.155 1676.285 2701.325 1676.665 ;
        RECT 2699.280 1675.860 2699.450 1676.115 ;
        RECT 2699.165 1675.530 2699.450 1675.860 ;
        RECT 2699.685 1675.565 2700.015 1675.935 ;
        RECT 2699.280 1675.385 2699.450 1675.530 ;
        RECT 2697.960 1674.485 2698.145 1674.890 ;
        RECT 2698.825 1674.455 2699.095 1675.360 ;
        RECT 2699.280 1675.215 2699.945 1675.385 ;
        RECT 2699.775 1674.455 2699.945 1675.215 ;
        RECT 2700.205 1675.360 2700.375 1676.160 ;
        RECT 2700.660 1676.115 2701.325 1676.285 ;
        RECT 2709.035 1676.285 2709.205 1676.665 ;
        RECT 2709.035 1676.115 2709.750 1676.285 ;
        RECT 2700.660 1675.860 2700.830 1676.115 ;
        RECT 2700.545 1675.530 2700.830 1675.860 ;
        RECT 2701.065 1675.565 2701.395 1675.935 ;
        RECT 2709.580 1675.925 2709.750 1676.115 ;
        RECT 2709.920 1676.090 2710.175 1676.665 ;
        RECT 2722.335 1676.265 2722.540 1676.665 ;
        RECT 2723.235 1676.335 2723.495 1676.665 ;
        RECT 2709.580 1675.595 2709.835 1675.925 ;
        RECT 2700.660 1675.385 2700.830 1675.530 ;
        RECT 2709.580 1675.385 2709.750 1675.595 ;
        RECT 2700.205 1674.455 2700.475 1675.360 ;
        RECT 2700.660 1675.215 2701.325 1675.385 ;
        RECT 2701.155 1674.455 2701.325 1675.215 ;
        RECT 2709.035 1675.215 2709.750 1675.385 ;
        RECT 2710.005 1675.360 2710.175 1676.090 ;
        RECT 2709.035 1674.455 2709.205 1675.215 ;
        RECT 2709.920 1674.455 2710.175 1675.360 ;
        RECT 2721.855 1676.095 2722.540 1676.265 ;
        RECT 2721.855 1675.065 2722.195 1676.095 ;
        RECT 2722.365 1675.425 2722.615 1675.925 ;
        RECT 2723.325 1675.425 2723.495 1676.335 ;
        RECT 2722.365 1675.255 2723.495 1675.425 ;
        RECT 2721.855 1674.890 2722.520 1675.065 ;
        RECT 2722.335 1674.485 2722.520 1674.890 ;
        RECT 2723.225 1674.485 2723.495 1675.255 ;
        RECT 2731.485 1676.160 2731.745 1676.665 ;
        RECT 2732.435 1676.285 2732.605 1676.665 ;
        RECT 2731.485 1675.360 2731.665 1676.160 ;
        RECT 2731.940 1676.115 2732.605 1676.285 ;
        RECT 2731.940 1675.860 2732.110 1676.115 ;
        RECT 2731.835 1675.530 2732.110 1675.860 ;
        RECT 2731.940 1675.385 2732.110 1675.530 ;
        RECT 2731.485 1674.455 2731.755 1675.360 ;
        RECT 2731.940 1675.215 2732.615 1675.385 ;
        RECT 2732.435 1674.455 2732.615 1675.215 ;
        RECT 2697.075 1673.185 2697.245 1673.945 ;
        RECT 2697.075 1673.015 2697.740 1673.185 ;
        RECT 2697.925 1673.040 2698.195 1673.945 ;
        RECT 2697.570 1672.870 2697.740 1673.015 ;
        RECT 2697.005 1672.465 2697.335 1672.835 ;
        RECT 2697.570 1672.540 2697.855 1672.870 ;
        RECT 2697.570 1672.285 2697.740 1672.540 ;
        RECT 2697.075 1672.115 2697.740 1672.285 ;
        RECT 2698.025 1672.240 2698.195 1673.040 ;
        RECT 2697.075 1671.735 2697.245 1672.115 ;
        RECT 2697.935 1671.735 2698.195 1672.240 ;
        RECT 2697.075 1665.405 2697.245 1665.785 ;
        RECT 2697.075 1665.235 2697.740 1665.405 ;
        RECT 2697.935 1665.280 2698.195 1665.785 ;
        RECT 2697.005 1664.685 2697.335 1665.055 ;
        RECT 2697.570 1664.980 2697.740 1665.235 ;
        RECT 2697.570 1664.650 2697.855 1664.980 ;
        RECT 2697.570 1664.505 2697.740 1664.650 ;
        RECT 2697.075 1664.335 2697.740 1664.505 ;
        RECT 2698.025 1664.480 2698.195 1665.280 ;
        RECT 2697.075 1663.575 2697.245 1664.335 ;
        RECT 2697.925 1663.575 2698.195 1664.480 ;
        RECT 2697.075 1659.965 2697.245 1660.340 ;
        RECT 2697.915 1660.175 2698.990 1660.345 ;
        RECT 2697.915 1659.965 2698.085 1660.175 ;
        RECT 2697.075 1659.795 2698.085 1659.965 ;
        RECT 2698.310 1659.835 2698.650 1660.005 ;
        RECT 2698.820 1659.840 2698.990 1660.175 ;
        RECT 2700.280 1660.175 2701.880 1660.345 ;
        RECT 2698.310 1659.665 2698.600 1659.835 ;
        RECT 2697.050 1659.495 2697.395 1659.605 ;
        RECT 2697.045 1659.325 2697.395 1659.495 ;
        RECT 2697.050 1658.985 2697.395 1659.325 ;
        RECT 2697.705 1658.985 2698.140 1659.605 ;
        RECT 2698.310 1659.145 2698.480 1659.665 ;
        RECT 2699.160 1659.495 2699.520 1660.170 ;
        RECT 2700.280 1659.805 2700.450 1660.175 ;
        RECT 2701.525 1660.135 2701.880 1660.175 ;
        RECT 2700.620 1659.755 2700.950 1660.005 ;
        RECT 2700.635 1659.680 2700.950 1659.755 ;
        RECT 2701.120 1659.885 2701.290 1660.005 ;
        RECT 2702.395 1659.885 2702.640 1660.305 ;
        RECT 2703.410 1659.945 2703.585 1660.275 ;
        RECT 2703.930 1660.185 2704.100 1660.345 ;
        RECT 2703.930 1660.015 2704.460 1660.185 ;
        RECT 2704.630 1660.175 2705.625 1660.345 ;
        RECT 2704.630 1660.015 2704.800 1660.175 ;
        RECT 2701.120 1659.715 2702.640 1659.885 ;
        RECT 2698.980 1659.315 2699.520 1659.495 ;
        RECT 2699.160 1659.205 2699.520 1659.315 ;
        RECT 2698.310 1658.975 2698.945 1659.145 ;
        RECT 2699.160 1658.975 2699.965 1659.205 ;
        RECT 2697.075 1658.635 2698.605 1658.805 ;
        RECT 2697.075 1658.135 2697.245 1658.635 ;
        RECT 2698.435 1658.475 2698.605 1658.635 ;
        RECT 2698.775 1658.645 2698.945 1658.975 ;
        RECT 2698.775 1658.475 2699.105 1658.645 ;
        RECT 2697.915 1658.305 2698.085 1658.465 ;
        RECT 2699.275 1658.305 2699.445 1658.805 ;
        RECT 2697.915 1658.135 2699.445 1658.305 ;
        RECT 2699.615 1658.135 2699.965 1658.975 ;
        RECT 2700.165 1658.605 2700.465 1659.605 ;
        RECT 2700.635 1659.155 2700.805 1659.680 ;
        RECT 2701.120 1659.675 2701.290 1659.715 ;
        RECT 2700.975 1659.495 2701.305 1659.505 ;
        RECT 2700.975 1659.335 2701.360 1659.495 ;
        RECT 2701.190 1659.325 2701.360 1659.335 ;
        RECT 2701.700 1659.155 2701.945 1659.545 ;
        RECT 2700.635 1658.985 2701.395 1659.155 ;
        RECT 2701.645 1658.985 2701.945 1659.155 ;
        RECT 2700.725 1658.305 2700.895 1658.815 ;
        RECT 2701.065 1658.475 2701.395 1658.985 ;
        RECT 2701.700 1658.925 2701.945 1658.985 ;
        RECT 2702.150 1658.925 2702.480 1659.545 ;
        RECT 2702.955 1658.925 2703.245 1659.605 ;
        RECT 2703.415 1659.495 2703.585 1659.945 ;
        RECT 2703.880 1659.665 2704.120 1659.835 ;
        RECT 2703.415 1659.325 2703.705 1659.495 ;
        RECT 2701.565 1658.515 2702.630 1658.685 ;
        RECT 2701.565 1658.305 2701.735 1658.515 ;
        RECT 2700.725 1658.135 2701.735 1658.305 ;
        RECT 2702.460 1658.135 2702.630 1658.515 ;
        RECT 2703.415 1658.465 2703.585 1659.325 ;
        RECT 2703.400 1658.135 2703.585 1658.465 ;
        RECT 2703.880 1658.465 2704.050 1659.665 ;
        RECT 2704.290 1658.845 2704.460 1660.015 ;
        RECT 2705.110 1659.835 2705.285 1660.005 ;
        RECT 2704.870 1659.675 2705.285 1659.835 ;
        RECT 2705.455 1659.885 2705.625 1660.175 ;
        RECT 2705.455 1659.715 2706.025 1659.885 ;
        RECT 2704.870 1659.665 2705.280 1659.675 ;
        RECT 2705.090 1659.325 2705.545 1659.495 ;
        RECT 2705.855 1658.935 2706.025 1659.715 ;
        RECT 2704.290 1658.615 2705.075 1658.845 ;
        RECT 2704.745 1658.475 2705.075 1658.615 ;
        RECT 2705.375 1658.765 2706.025 1658.935 ;
        RECT 2703.880 1658.135 2704.090 1658.465 ;
        RECT 2704.260 1658.305 2704.590 1658.345 ;
        RECT 2705.375 1658.305 2705.545 1658.765 ;
        RECT 2704.260 1658.135 2705.545 1658.305 ;
        RECT 2706.215 1658.135 2706.475 1660.345 ;
        RECT 2697.075 1656.865 2697.245 1657.625 ;
        RECT 2697.075 1656.695 2697.740 1656.865 ;
        RECT 2697.925 1656.720 2698.195 1657.625 ;
        RECT 2697.570 1656.550 2697.740 1656.695 ;
        RECT 2697.005 1656.145 2697.335 1656.515 ;
        RECT 2697.570 1656.220 2697.855 1656.550 ;
        RECT 2697.570 1655.965 2697.740 1656.220 ;
        RECT 2697.075 1655.795 2697.740 1655.965 ;
        RECT 2698.025 1655.920 2698.195 1656.720 ;
        RECT 2697.075 1655.415 2697.245 1655.795 ;
        RECT 2697.935 1655.415 2698.195 1655.920 ;
        RECT 2697.075 1654.525 2697.245 1654.900 ;
        RECT 2697.915 1654.735 2698.990 1654.905 ;
        RECT 2697.915 1654.525 2698.085 1654.735 ;
        RECT 2697.075 1654.355 2698.085 1654.525 ;
        RECT 2698.310 1654.395 2698.650 1654.565 ;
        RECT 2698.820 1654.400 2698.990 1654.735 ;
        RECT 2700.280 1654.735 2701.880 1654.905 ;
        RECT 2698.310 1654.225 2698.600 1654.395 ;
        RECT 2697.050 1654.055 2697.395 1654.165 ;
        RECT 2697.045 1653.885 2697.395 1654.055 ;
        RECT 2697.050 1653.545 2697.395 1653.885 ;
        RECT 2697.705 1653.545 2698.140 1654.165 ;
        RECT 2698.310 1653.705 2698.480 1654.225 ;
        RECT 2699.160 1654.055 2699.520 1654.730 ;
        RECT 2700.280 1654.365 2700.450 1654.735 ;
        RECT 2701.525 1654.695 2701.880 1654.735 ;
        RECT 2700.620 1654.315 2700.950 1654.565 ;
        RECT 2700.635 1654.240 2700.950 1654.315 ;
        RECT 2701.120 1654.445 2701.290 1654.565 ;
        RECT 2702.395 1654.445 2702.640 1654.865 ;
        RECT 2703.410 1654.505 2703.585 1654.835 ;
        RECT 2703.930 1654.745 2704.100 1654.905 ;
        RECT 2703.930 1654.575 2704.460 1654.745 ;
        RECT 2704.630 1654.735 2705.625 1654.905 ;
        RECT 2704.630 1654.575 2704.800 1654.735 ;
        RECT 2701.120 1654.275 2702.640 1654.445 ;
        RECT 2698.980 1653.875 2699.520 1654.055 ;
        RECT 2699.160 1653.765 2699.520 1653.875 ;
        RECT 2698.310 1653.535 2698.945 1653.705 ;
        RECT 2699.160 1653.535 2699.965 1653.765 ;
        RECT 2697.075 1653.195 2698.605 1653.365 ;
        RECT 2697.075 1652.695 2697.245 1653.195 ;
        RECT 2698.435 1653.035 2698.605 1653.195 ;
        RECT 2698.775 1653.205 2698.945 1653.535 ;
        RECT 2698.775 1653.035 2699.105 1653.205 ;
        RECT 2697.915 1652.865 2698.085 1653.025 ;
        RECT 2699.275 1652.865 2699.445 1653.365 ;
        RECT 2697.915 1652.695 2699.445 1652.865 ;
        RECT 2699.615 1652.695 2699.965 1653.535 ;
        RECT 2700.165 1653.165 2700.465 1654.165 ;
        RECT 2700.635 1653.715 2700.805 1654.240 ;
        RECT 2701.120 1654.235 2701.290 1654.275 ;
        RECT 2700.975 1654.055 2701.305 1654.065 ;
        RECT 2700.975 1653.895 2701.360 1654.055 ;
        RECT 2701.190 1653.885 2701.360 1653.895 ;
        RECT 2701.700 1653.715 2701.945 1654.105 ;
        RECT 2700.635 1653.545 2701.395 1653.715 ;
        RECT 2701.645 1653.545 2701.945 1653.715 ;
        RECT 2700.725 1652.865 2700.895 1653.375 ;
        RECT 2701.065 1653.035 2701.395 1653.545 ;
        RECT 2701.700 1653.485 2701.945 1653.545 ;
        RECT 2702.150 1653.485 2702.480 1654.105 ;
        RECT 2702.955 1653.485 2703.245 1654.165 ;
        RECT 2703.415 1654.055 2703.585 1654.505 ;
        RECT 2703.880 1654.225 2704.120 1654.395 ;
        RECT 2703.415 1653.885 2703.705 1654.055 ;
        RECT 2701.565 1653.075 2702.630 1653.245 ;
        RECT 2701.565 1652.865 2701.735 1653.075 ;
        RECT 2700.725 1652.695 2701.735 1652.865 ;
        RECT 2702.460 1652.695 2702.630 1653.075 ;
        RECT 2703.415 1653.025 2703.585 1653.885 ;
        RECT 2703.400 1652.695 2703.585 1653.025 ;
        RECT 2703.880 1653.025 2704.050 1654.225 ;
        RECT 2704.290 1653.405 2704.460 1654.575 ;
        RECT 2705.110 1654.395 2705.285 1654.565 ;
        RECT 2704.870 1654.235 2705.285 1654.395 ;
        RECT 2705.455 1654.445 2705.625 1654.735 ;
        RECT 2705.455 1654.275 2706.025 1654.445 ;
        RECT 2704.870 1654.225 2705.280 1654.235 ;
        RECT 2705.090 1653.885 2705.545 1654.055 ;
        RECT 2705.855 1653.495 2706.025 1654.275 ;
        RECT 2704.290 1653.175 2705.075 1653.405 ;
        RECT 2704.745 1653.035 2705.075 1653.175 ;
        RECT 2705.375 1653.325 2706.025 1653.495 ;
        RECT 2703.880 1652.695 2704.090 1653.025 ;
        RECT 2704.260 1652.865 2704.590 1652.905 ;
        RECT 2705.375 1652.865 2705.545 1653.325 ;
        RECT 2704.260 1652.695 2705.545 1652.865 ;
        RECT 2706.215 1652.695 2706.475 1654.905 ;
        RECT 2697.075 1651.425 2697.245 1652.185 ;
        RECT 2697.075 1651.255 2697.740 1651.425 ;
        RECT 2697.925 1651.280 2698.195 1652.185 ;
        RECT 2697.570 1651.110 2697.740 1651.255 ;
        RECT 2697.005 1650.705 2697.335 1651.075 ;
        RECT 2697.570 1650.780 2697.855 1651.110 ;
        RECT 2697.570 1650.525 2697.740 1650.780 ;
        RECT 2697.075 1650.355 2697.740 1650.525 ;
        RECT 2698.025 1650.480 2698.195 1651.280 ;
        RECT 2697.075 1649.975 2697.245 1650.355 ;
        RECT 2697.935 1649.975 2698.195 1650.480 ;
        RECT 2701.590 1651.215 2701.925 1652.185 ;
        RECT 2702.435 1652.015 2704.465 1652.185 ;
        RECT 2701.590 1650.545 2701.760 1651.215 ;
        RECT 2702.435 1651.045 2702.605 1652.015 ;
        RECT 2701.930 1650.715 2702.185 1651.045 ;
        RECT 2702.410 1650.715 2702.605 1651.045 ;
        RECT 2702.775 1651.675 2703.900 1651.845 ;
        RECT 2702.015 1650.545 2702.185 1650.715 ;
        RECT 2702.775 1650.545 2702.945 1651.675 ;
        RECT 2701.590 1649.975 2701.845 1650.545 ;
        RECT 2702.015 1650.375 2702.945 1650.545 ;
        RECT 2703.115 1651.335 2704.125 1651.505 ;
        RECT 2703.115 1650.535 2703.285 1651.335 ;
        RECT 2703.490 1650.655 2703.765 1651.135 ;
        RECT 2703.485 1650.485 2703.765 1650.655 ;
        RECT 2702.770 1650.340 2702.945 1650.375 ;
        RECT 2702.770 1649.975 2703.300 1650.340 ;
        RECT 2703.490 1649.975 2703.765 1650.485 ;
        RECT 2703.935 1649.975 2704.125 1651.335 ;
        RECT 2704.295 1651.350 2704.465 1652.015 ;
        RECT 2705.040 1651.595 2705.555 1652.005 ;
        RECT 2704.295 1651.160 2705.045 1651.350 ;
        RECT 2705.215 1650.785 2705.555 1651.595 ;
        RECT 2704.325 1650.615 2705.555 1650.785 ;
        RECT 2705.035 1650.010 2705.280 1650.615 ;
        RECT 2697.075 1645.985 2697.245 1646.745 ;
        RECT 2697.075 1645.815 2697.740 1645.985 ;
        RECT 2697.925 1645.840 2698.195 1646.745 ;
        RECT 2697.570 1645.670 2697.740 1645.815 ;
        RECT 2697.005 1645.265 2697.335 1645.635 ;
        RECT 2697.570 1645.340 2697.855 1645.670 ;
        RECT 2697.570 1645.085 2697.740 1645.340 ;
        RECT 2697.075 1644.915 2697.740 1645.085 ;
        RECT 2698.025 1645.040 2698.195 1645.840 ;
        RECT 2697.075 1644.535 2697.245 1644.915 ;
        RECT 2697.935 1644.535 2698.195 1645.040 ;
        RECT 2701.595 1640.505 2701.925 1641.290 ;
        RECT 2701.595 1640.335 2702.275 1640.505 ;
        RECT 2701.585 1639.915 2701.935 1640.165 ;
        RECT 2702.105 1639.735 2702.275 1640.335 ;
        RECT 2702.445 1639.915 2702.795 1640.165 ;
        RECT 2702.015 1639.095 2702.345 1639.735 ;
        RECT 2697.075 1638.205 2697.245 1638.585 ;
        RECT 2697.075 1638.035 2697.740 1638.205 ;
        RECT 2697.935 1638.080 2698.195 1638.585 ;
        RECT 2697.005 1637.485 2697.335 1637.855 ;
        RECT 2697.570 1637.780 2697.740 1638.035 ;
        RECT 2697.570 1637.450 2697.855 1637.780 ;
        RECT 2697.570 1637.305 2697.740 1637.450 ;
        RECT 2697.075 1637.135 2697.740 1637.305 ;
        RECT 2698.025 1637.280 2698.195 1638.080 ;
        RECT 2702.565 1638.225 2702.885 1638.585 ;
        RECT 2703.880 1638.225 2704.225 1638.585 ;
        RECT 2702.565 1638.055 2704.225 1638.225 ;
        RECT 2697.075 1636.375 2697.245 1637.135 ;
        RECT 2697.925 1636.375 2698.195 1637.280 ;
        RECT 2702.105 1637.215 2702.380 1637.845 ;
        RECT 2702.090 1636.555 2702.395 1637.045 ;
        RECT 2702.565 1636.725 2702.865 1638.055 ;
        RECT 2703.245 1637.595 2703.575 1637.765 ;
        RECT 2703.250 1637.345 2703.575 1637.595 ;
        RECT 2703.755 1637.515 2704.365 1637.845 ;
        RECT 2704.535 1637.345 2705.035 1637.805 ;
        RECT 2703.250 1637.165 2705.035 1637.345 ;
        RECT 2703.035 1636.815 2705.070 1636.985 ;
        RECT 2703.035 1636.555 2703.365 1636.815 ;
        RECT 2702.090 1636.375 2703.365 1636.555 ;
        RECT 2703.960 1636.735 2705.070 1636.815 ;
        RECT 2703.960 1636.375 2704.130 1636.735 ;
        RECT 2704.810 1636.375 2705.070 1636.735 ;
        RECT 2725.935 1635.015 2726.265 1635.865 ;
        RECT 2726.775 1635.015 2727.105 1635.865 ;
        RECT 2725.935 1634.845 2727.435 1635.015 ;
        RECT 2725.555 1634.475 2727.080 1634.675 ;
        RECT 2727.260 1634.645 2727.435 1634.845 ;
        RECT 2727.260 1634.475 2729.885 1634.645 ;
        RECT 2727.260 1634.305 2727.435 1634.475 ;
        RECT 2726.015 1634.135 2727.435 1634.305 ;
        RECT 2726.015 1633.655 2726.185 1634.135 ;
        RECT 2726.855 1633.660 2727.025 1634.135 ;
        RECT 2697.075 1632.765 2697.245 1633.145 ;
        RECT 2697.075 1632.595 2697.740 1632.765 ;
        RECT 2697.935 1632.640 2698.195 1633.145 ;
        RECT 2697.005 1632.045 2697.335 1632.415 ;
        RECT 2697.570 1632.340 2697.740 1632.595 ;
        RECT 2697.570 1632.010 2697.855 1632.340 ;
        RECT 2697.570 1631.865 2697.740 1632.010 ;
        RECT 2697.075 1631.695 2697.740 1631.865 ;
        RECT 2698.025 1631.840 2698.195 1632.640 ;
        RECT 2697.075 1630.935 2697.245 1631.695 ;
        RECT 2697.925 1630.935 2698.195 1631.840 ;
        RECT 2697.310 1627.305 2697.480 1627.555 ;
        RECT 2696.985 1627.135 2697.480 1627.305 ;
        RECT 2698.215 1627.305 2698.385 1627.650 ;
        RECT 2699.055 1627.305 2699.575 1627.705 ;
        RECT 2698.215 1627.135 2699.575 1627.305 ;
        RECT 2696.985 1626.175 2697.155 1627.135 ;
        RECT 2697.325 1626.345 2697.675 1626.965 ;
        RECT 2697.845 1626.345 2698.185 1626.965 ;
        RECT 2698.355 1626.345 2698.595 1626.965 ;
        RECT 2698.775 1626.715 2699.235 1626.885 ;
        RECT 2698.775 1626.175 2698.945 1626.715 ;
        RECT 2699.405 1626.515 2699.575 1627.135 ;
        RECT 2882.085 1626.620 2882.605 1628.170 ;
        RECT 2522.640 1623.850 2523.160 1625.335 ;
        RECT 2523.330 1624.510 2523.850 1626.060 ;
        RECT 2696.985 1626.005 2698.945 1626.175 ;
        RECT 2699.115 1625.505 2699.575 1626.515 ;
        RECT 2697.075 1624.225 2697.245 1624.985 ;
        RECT 2697.075 1624.055 2697.740 1624.225 ;
        RECT 2697.925 1624.080 2698.195 1624.985 ;
        RECT 2697.570 1623.910 2697.740 1624.055 ;
        RECT 2697.005 1623.505 2697.335 1623.875 ;
        RECT 2697.570 1623.580 2697.855 1623.910 ;
        RECT 2697.570 1623.325 2697.740 1623.580 ;
        RECT 2697.075 1623.155 2697.740 1623.325 ;
        RECT 2698.025 1623.280 2698.195 1624.080 ;
        RECT 2697.075 1622.775 2697.245 1623.155 ;
        RECT 2697.935 1622.775 2698.195 1623.280 ;
        RECT 2697.260 1621.625 2697.505 1622.230 ;
        RECT 2696.985 1621.455 2698.215 1621.625 ;
        RECT 2696.985 1620.645 2697.325 1621.455 ;
        RECT 2697.495 1620.890 2698.245 1621.080 ;
        RECT 2696.985 1620.235 2697.500 1620.645 ;
        RECT 2698.075 1620.225 2698.245 1620.890 ;
        RECT 2698.415 1620.905 2698.605 1622.265 ;
        RECT 2698.775 1622.095 2699.050 1622.265 ;
        RECT 2698.775 1621.925 2699.055 1622.095 ;
        RECT 2698.775 1621.105 2699.050 1621.925 ;
        RECT 2699.240 1621.900 2699.770 1622.265 ;
        RECT 2699.595 1621.865 2699.770 1621.900 ;
        RECT 2699.255 1620.905 2699.425 1621.705 ;
        RECT 2698.415 1620.735 2699.425 1620.905 ;
        RECT 2699.595 1621.695 2700.525 1621.865 ;
        RECT 2700.695 1621.695 2700.950 1622.265 ;
        RECT 2699.595 1620.565 2699.765 1621.695 ;
        RECT 2700.355 1621.525 2700.525 1621.695 ;
        RECT 2698.640 1620.395 2699.765 1620.565 ;
        RECT 2699.935 1621.195 2700.130 1621.525 ;
        RECT 2700.355 1621.195 2700.610 1621.525 ;
        RECT 2699.935 1620.225 2700.105 1621.195 ;
        RECT 2700.780 1621.025 2700.950 1621.695 ;
        RECT 2701.630 1621.500 2701.815 1622.170 ;
        RECT 2702.300 1621.815 2702.630 1622.215 ;
        RECT 2703.345 1621.820 2703.675 1622.260 ;
        RECT 2703.345 1621.815 2704.575 1621.820 ;
        RECT 2702.300 1621.705 2704.575 1621.815 ;
        RECT 2702.420 1621.640 2704.575 1621.705 ;
        RECT 2701.180 1621.230 2701.815 1621.500 ;
        RECT 2701.995 1621.120 2702.280 1621.525 ;
        RECT 2702.450 1621.120 2702.780 1621.470 ;
        RECT 2698.075 1620.055 2700.105 1620.225 ;
        RECT 2700.615 1620.055 2700.950 1621.025 ;
        RECT 2701.215 1620.770 2702.325 1620.940 ;
        RECT 2701.215 1620.060 2701.410 1620.770 ;
        RECT 2702.095 1620.060 2702.325 1620.770 ;
        RECT 2702.505 1620.065 2702.780 1621.120 ;
        RECT 2702.950 1620.065 2703.285 1621.470 ;
        RECT 2703.485 1620.065 2703.935 1621.470 ;
        RECT 2704.190 1620.060 2704.575 1621.640 ;
        RECT 2522.640 1617.435 2523.160 1618.920 ;
        RECT 2523.330 1618.095 2523.850 1619.645 ;
        RECT 2696.985 1618.155 2697.325 1619.035 ;
        RECT 2697.495 1618.325 2697.665 1619.545 ;
        RECT 2698.690 1619.205 2699.165 1619.545 ;
        RECT 2697.905 1618.675 2698.155 1619.040 ;
        RECT 2698.875 1618.675 2699.590 1618.970 ;
        RECT 2699.760 1618.845 2700.035 1619.545 ;
        RECT 2697.905 1618.505 2699.695 1618.675 ;
        RECT 2697.495 1618.075 2698.290 1618.325 ;
        RECT 2697.495 1617.985 2697.745 1618.075 ;
        RECT 2697.415 1617.565 2697.745 1617.985 ;
        RECT 2698.460 1617.650 2698.715 1618.505 ;
        RECT 2697.925 1617.385 2698.715 1617.650 ;
        RECT 2698.885 1617.805 2699.295 1618.325 ;
        RECT 2699.465 1618.075 2699.695 1618.505 ;
        RECT 2699.865 1617.815 2700.035 1618.845 ;
        RECT 2698.885 1617.385 2699.085 1617.805 ;
        RECT 2699.775 1617.335 2700.035 1617.815 ;
        RECT 2697.075 1616.445 2697.245 1616.825 ;
        RECT 2697.075 1616.275 2697.740 1616.445 ;
        RECT 2697.935 1616.320 2698.195 1616.825 ;
        RECT 2697.005 1615.725 2697.335 1616.095 ;
        RECT 2697.570 1616.020 2697.740 1616.275 ;
        RECT 2697.570 1615.690 2697.855 1616.020 ;
        RECT 2697.570 1615.545 2697.740 1615.690 ;
        RECT 2697.075 1615.375 2697.740 1615.545 ;
        RECT 2698.025 1615.520 2698.195 1616.320 ;
        RECT 2697.075 1614.615 2697.245 1615.375 ;
        RECT 2697.925 1614.615 2698.195 1615.520 ;
        RECT 2698.455 1613.605 2698.625 1614.105 ;
        RECT 2699.415 1613.605 2699.585 1614.105 ;
        RECT 2700.255 1613.605 2700.425 1614.105 ;
        RECT 2698.455 1613.435 2700.425 1613.605 ;
        RECT 2700.595 1613.635 2700.925 1614.065 ;
        RECT 2701.535 1613.805 2701.875 1614.065 ;
        RECT 2700.595 1613.465 2701.445 1613.635 ;
        RECT 2698.390 1612.635 2698.645 1613.265 ;
        RECT 2698.875 1612.635 2699.255 1613.265 ;
        RECT 2700.125 1613.255 2700.425 1613.260 ;
        RECT 2700.125 1613.085 2700.435 1613.255 ;
        RECT 2700.125 1612.965 2700.425 1613.085 ;
        RECT 2698.875 1612.035 2699.080 1612.635 ;
        RECT 2699.515 1612.240 2699.735 1612.965 ;
        RECT 2700.045 1612.635 2700.425 1612.965 ;
        RECT 2700.625 1612.715 2700.955 1613.275 ;
        RECT 2701.275 1612.545 2701.445 1613.465 ;
        RECT 2700.625 1612.450 2701.445 1612.545 ;
        RECT 2700.430 1612.375 2701.445 1612.450 ;
        RECT 2699.310 1612.055 2700.260 1612.240 ;
        RECT 2700.430 1611.940 2700.845 1612.375 ;
        RECT 2701.615 1612.200 2701.875 1613.805 ;
        RECT 2701.535 1611.940 2701.875 1612.200 ;
        RECT 2698.335 1610.735 2698.665 1611.155 ;
        RECT 2698.845 1610.985 2699.105 1611.385 ;
        RECT 2699.775 1610.985 2699.945 1611.335 ;
        RECT 2698.845 1610.815 2700.510 1610.985 ;
        RECT 2700.680 1610.880 2700.955 1611.225 ;
        RECT 2698.415 1610.645 2698.665 1610.735 ;
        RECT 2700.340 1610.645 2700.510 1610.815 ;
        RECT 2358.645 1610.105 2358.820 1610.595 ;
        RECT 2359.170 1610.315 2359.340 1610.595 ;
        RECT 2359.170 1610.145 2359.400 1610.315 ;
        RECT 2358.645 1609.935 2358.815 1610.105 ;
        RECT 2358.645 1609.605 2359.055 1609.935 ;
        RECT 2358.645 1609.095 2358.815 1609.605 ;
        RECT 2358.645 1608.765 2359.055 1609.095 ;
        RECT 2358.645 1608.565 2358.815 1608.765 ;
        RECT 2358.645 1607.305 2358.820 1608.565 ;
        RECT 2359.230 1608.535 2359.400 1610.145 ;
        RECT 2359.600 1610.085 2359.775 1610.595 ;
        RECT 2362.055 1610.105 2362.230 1610.595 ;
        RECT 2362.055 1609.935 2362.225 1610.105 ;
        RECT 2363.010 1610.085 2363.185 1610.595 ;
        RECT 2363.440 1610.045 2363.615 1610.595 ;
        RECT 2373.740 1610.105 2373.915 1610.595 ;
        RECT 2374.265 1610.315 2374.435 1610.595 ;
        RECT 2374.265 1610.145 2374.495 1610.315 ;
        RECT 2362.055 1609.605 2362.465 1609.935 ;
        RECT 2359.170 1608.365 2359.400 1608.535 ;
        RECT 2359.600 1608.565 2359.770 1609.515 ;
        RECT 2362.055 1609.095 2362.225 1609.605 ;
        RECT 2362.055 1608.765 2362.465 1609.095 ;
        RECT 2362.055 1608.565 2362.225 1608.765 ;
        RECT 2363.010 1608.565 2363.180 1609.515 ;
        RECT 2359.170 1607.305 2359.340 1608.365 ;
        RECT 2359.600 1607.305 2359.775 1608.565 ;
        RECT 2362.055 1607.305 2362.230 1608.565 ;
        RECT 2363.010 1607.305 2363.185 1608.565 ;
        RECT 2363.440 1608.445 2363.610 1610.045 ;
        RECT 2373.740 1609.935 2373.910 1610.105 ;
        RECT 2373.740 1609.605 2374.150 1609.935 ;
        RECT 2373.740 1609.095 2373.910 1609.605 ;
        RECT 2373.740 1608.765 2374.150 1609.095 ;
        RECT 2373.740 1608.565 2373.910 1608.765 ;
        RECT 2363.440 1607.305 2363.615 1608.445 ;
        RECT 2365.645 1607.560 2366.340 1608.190 ;
        RECT 2365.645 1606.960 2365.815 1607.560 ;
        RECT 2365.985 1607.340 2366.320 1607.370 ;
        RECT 2366.710 1607.340 2366.880 1608.020 ;
        RECT 2365.985 1607.170 2366.880 1607.340 ;
        RECT 2367.945 1607.560 2368.640 1608.190 ;
        RECT 2368.810 1607.560 2369.505 1608.190 ;
        RECT 2370.190 1607.560 2370.885 1608.190 ;
        RECT 2365.985 1607.120 2366.320 1607.170 ;
        RECT 2367.945 1606.960 2368.115 1607.560 ;
        RECT 2368.285 1607.340 2368.620 1607.370 ;
        RECT 2368.830 1607.340 2369.165 1607.370 ;
        RECT 2368.285 1607.170 2369.165 1607.340 ;
        RECT 2368.285 1607.120 2368.620 1607.170 ;
        RECT 2368.830 1607.120 2369.165 1607.170 ;
        RECT 2369.335 1606.960 2369.505 1607.560 ;
        RECT 2369.675 1607.120 2370.010 1607.390 ;
        RECT 2370.210 1607.120 2370.545 1607.370 ;
        RECT 2370.715 1606.960 2370.885 1607.560 ;
        RECT 2371.055 1607.120 2371.390 1607.390 ;
        RECT 2373.740 1607.305 2373.915 1608.565 ;
        RECT 2374.325 1608.535 2374.495 1610.145 ;
        RECT 2374.695 1610.085 2374.870 1610.595 ;
        RECT 2375.125 1610.045 2375.300 1610.595 ;
        RECT 2376.490 1610.085 2376.660 1610.595 ;
        RECT 2377.480 1610.085 2377.650 1610.595 ;
        RECT 2379.275 1610.105 2379.450 1610.595 ;
        RECT 2374.265 1608.365 2374.495 1608.535 ;
        RECT 2374.695 1608.565 2374.865 1609.515 ;
        RECT 2374.265 1607.305 2374.435 1608.365 ;
        RECT 2374.695 1607.305 2374.870 1608.565 ;
        RECT 2375.125 1608.445 2375.295 1610.045 ;
        RECT 2379.275 1609.935 2379.445 1610.105 ;
        RECT 2380.230 1610.085 2380.405 1610.595 ;
        RECT 2380.660 1610.045 2380.835 1610.595 ;
        RECT 2390.960 1610.105 2391.135 1610.595 ;
        RECT 2391.485 1610.315 2391.655 1610.595 ;
        RECT 2391.485 1610.145 2391.715 1610.315 ;
        RECT 2376.055 1609.425 2376.285 1609.615 ;
        RECT 2379.275 1609.605 2379.685 1609.935 ;
        RECT 2376.055 1609.385 2376.585 1609.425 ;
        RECT 2376.115 1609.255 2376.585 1609.385 ;
        RECT 2377.105 1609.255 2377.575 1609.425 ;
        RECT 2376.115 1608.565 2376.285 1609.255 ;
        RECT 2376.485 1608.780 2376.655 1608.885 ;
        RECT 2377.105 1608.780 2377.275 1609.255 ;
        RECT 2379.275 1609.095 2379.445 1609.605 ;
        RECT 2376.485 1608.605 2377.275 1608.780 ;
        RECT 2375.125 1607.305 2375.300 1608.445 ;
        RECT 2376.485 1607.305 2376.660 1608.605 ;
        RECT 2377.105 1608.565 2377.275 1608.605 ;
        RECT 2377.475 1608.450 2377.645 1608.885 ;
        RECT 2379.275 1608.765 2379.685 1609.095 ;
        RECT 2379.275 1608.565 2379.445 1608.765 ;
        RECT 2380.230 1608.565 2380.400 1609.515 ;
        RECT 2377.475 1607.305 2377.650 1608.450 ;
        RECT 2379.275 1607.305 2379.450 1608.565 ;
        RECT 2380.230 1607.305 2380.405 1608.565 ;
        RECT 2380.660 1608.445 2380.830 1610.045 ;
        RECT 2390.960 1609.935 2391.130 1610.105 ;
        RECT 2390.960 1609.605 2391.370 1609.935 ;
        RECT 2390.960 1609.095 2391.130 1609.605 ;
        RECT 2390.960 1608.765 2391.370 1609.095 ;
        RECT 2390.960 1608.565 2391.130 1608.765 ;
        RECT 2380.660 1607.305 2380.835 1608.445 ;
        RECT 2382.865 1607.560 2383.560 1608.190 ;
        RECT 2382.865 1606.960 2383.035 1607.560 ;
        RECT 2383.205 1607.340 2383.540 1607.370 ;
        RECT 2383.930 1607.340 2384.100 1608.020 ;
        RECT 2383.205 1607.170 2384.100 1607.340 ;
        RECT 2385.165 1607.560 2385.860 1608.190 ;
        RECT 2386.030 1607.560 2386.725 1608.190 ;
        RECT 2387.410 1607.560 2388.105 1608.190 ;
        RECT 2383.205 1607.120 2383.540 1607.170 ;
        RECT 2385.165 1606.960 2385.335 1607.560 ;
        RECT 2385.505 1607.340 2385.840 1607.370 ;
        RECT 2386.050 1607.340 2386.385 1607.370 ;
        RECT 2385.505 1607.170 2386.385 1607.340 ;
        RECT 2385.505 1607.120 2385.840 1607.170 ;
        RECT 2386.050 1607.120 2386.385 1607.170 ;
        RECT 2386.555 1606.960 2386.725 1607.560 ;
        RECT 2386.895 1607.120 2387.230 1607.390 ;
        RECT 2387.430 1607.120 2387.765 1607.370 ;
        RECT 2387.935 1606.960 2388.105 1607.560 ;
        RECT 2388.275 1607.120 2388.610 1607.390 ;
        RECT 2390.960 1607.305 2391.135 1608.565 ;
        RECT 2391.545 1608.535 2391.715 1610.145 ;
        RECT 2391.915 1610.085 2392.090 1610.595 ;
        RECT 2392.345 1610.045 2392.520 1610.595 ;
        RECT 2393.710 1610.085 2393.880 1610.595 ;
        RECT 2394.700 1610.085 2394.870 1610.595 ;
        RECT 2396.495 1610.110 2396.670 1610.600 ;
        RECT 2391.485 1608.365 2391.715 1608.535 ;
        RECT 2391.915 1608.565 2392.085 1609.515 ;
        RECT 2391.485 1607.305 2391.655 1608.365 ;
        RECT 2391.915 1607.305 2392.090 1608.565 ;
        RECT 2392.345 1608.445 2392.515 1610.045 ;
        RECT 2396.495 1609.940 2396.665 1610.110 ;
        RECT 2397.450 1610.090 2397.625 1610.600 ;
        RECT 2397.880 1610.050 2398.055 1610.600 ;
        RECT 2408.180 1610.110 2408.355 1610.600 ;
        RECT 2408.705 1610.320 2408.875 1610.600 ;
        RECT 2408.705 1610.150 2408.935 1610.320 ;
        RECT 2393.275 1609.425 2393.505 1609.615 ;
        RECT 2396.495 1609.610 2396.905 1609.940 ;
        RECT 2393.275 1609.385 2393.805 1609.425 ;
        RECT 2393.335 1609.255 2393.805 1609.385 ;
        RECT 2394.325 1609.255 2394.795 1609.425 ;
        RECT 2393.335 1608.565 2393.505 1609.255 ;
        RECT 2393.705 1608.780 2393.875 1608.885 ;
        RECT 2394.325 1608.780 2394.495 1609.255 ;
        RECT 2396.495 1609.100 2396.665 1609.610 ;
        RECT 2393.705 1608.605 2394.495 1608.780 ;
        RECT 2392.345 1607.305 2392.520 1608.445 ;
        RECT 2393.705 1607.305 2393.880 1608.605 ;
        RECT 2394.325 1608.565 2394.495 1608.605 ;
        RECT 2394.695 1608.450 2394.865 1608.885 ;
        RECT 2396.495 1608.770 2396.905 1609.100 ;
        RECT 2396.495 1608.570 2396.665 1608.770 ;
        RECT 2397.450 1608.570 2397.620 1609.520 ;
        RECT 2394.695 1607.305 2394.870 1608.450 ;
        RECT 2396.495 1607.310 2396.670 1608.570 ;
        RECT 2397.450 1607.310 2397.625 1608.570 ;
        RECT 2397.880 1608.450 2398.050 1610.050 ;
        RECT 2408.180 1609.940 2408.350 1610.110 ;
        RECT 2408.180 1609.610 2408.590 1609.940 ;
        RECT 2408.180 1609.100 2408.350 1609.610 ;
        RECT 2408.180 1608.770 2408.590 1609.100 ;
        RECT 2408.180 1608.570 2408.350 1608.770 ;
        RECT 2397.880 1607.310 2398.055 1608.450 ;
        RECT 2400.085 1607.565 2400.780 1608.195 ;
        RECT 2400.085 1606.965 2400.255 1607.565 ;
        RECT 2400.425 1607.345 2400.760 1607.375 ;
        RECT 2401.150 1607.345 2401.320 1608.025 ;
        RECT 2400.425 1607.175 2401.320 1607.345 ;
        RECT 2402.385 1607.565 2403.080 1608.195 ;
        RECT 2403.250 1607.565 2403.945 1608.195 ;
        RECT 2404.630 1607.565 2405.325 1608.195 ;
        RECT 2400.425 1607.125 2400.760 1607.175 ;
        RECT 2402.385 1606.965 2402.555 1607.565 ;
        RECT 2402.725 1607.345 2403.060 1607.375 ;
        RECT 2403.270 1607.345 2403.605 1607.375 ;
        RECT 2402.725 1607.175 2403.605 1607.345 ;
        RECT 2402.725 1607.125 2403.060 1607.175 ;
        RECT 2403.270 1607.125 2403.605 1607.175 ;
        RECT 2403.775 1606.965 2403.945 1607.565 ;
        RECT 2404.115 1607.125 2404.450 1607.395 ;
        RECT 2404.650 1607.125 2404.985 1607.375 ;
        RECT 2405.155 1606.965 2405.325 1607.565 ;
        RECT 2405.495 1607.125 2405.830 1607.395 ;
        RECT 2408.180 1607.310 2408.355 1608.570 ;
        RECT 2408.765 1608.540 2408.935 1610.150 ;
        RECT 2409.135 1610.090 2409.310 1610.600 ;
        RECT 2409.565 1610.050 2409.740 1610.600 ;
        RECT 2410.930 1610.090 2411.100 1610.600 ;
        RECT 2411.920 1610.090 2412.090 1610.600 ;
        RECT 2413.715 1610.105 2413.890 1610.595 ;
        RECT 2408.705 1608.370 2408.935 1608.540 ;
        RECT 2409.135 1608.570 2409.305 1609.520 ;
        RECT 2408.705 1607.310 2408.875 1608.370 ;
        RECT 2409.135 1607.310 2409.310 1608.570 ;
        RECT 2409.565 1608.450 2409.735 1610.050 ;
        RECT 2413.715 1609.935 2413.885 1610.105 ;
        RECT 2414.670 1610.085 2414.845 1610.595 ;
        RECT 2415.100 1610.045 2415.275 1610.595 ;
        RECT 2425.400 1610.105 2425.575 1610.595 ;
        RECT 2425.925 1610.315 2426.095 1610.595 ;
        RECT 2425.925 1610.145 2426.155 1610.315 ;
        RECT 2410.495 1609.430 2410.725 1609.620 ;
        RECT 2413.715 1609.605 2414.125 1609.935 ;
        RECT 2410.495 1609.390 2411.025 1609.430 ;
        RECT 2410.555 1609.260 2411.025 1609.390 ;
        RECT 2411.545 1609.260 2412.015 1609.430 ;
        RECT 2410.555 1608.570 2410.725 1609.260 ;
        RECT 2410.925 1608.785 2411.095 1608.890 ;
        RECT 2411.545 1608.785 2411.715 1609.260 ;
        RECT 2413.715 1609.095 2413.885 1609.605 ;
        RECT 2410.925 1608.610 2411.715 1608.785 ;
        RECT 2409.565 1607.310 2409.740 1608.450 ;
        RECT 2410.925 1607.310 2411.100 1608.610 ;
        RECT 2411.545 1608.570 2411.715 1608.610 ;
        RECT 2411.915 1608.455 2412.085 1608.890 ;
        RECT 2413.715 1608.765 2414.125 1609.095 ;
        RECT 2413.715 1608.565 2413.885 1608.765 ;
        RECT 2414.670 1608.565 2414.840 1609.515 ;
        RECT 2411.915 1607.310 2412.090 1608.455 ;
        RECT 2413.715 1607.305 2413.890 1608.565 ;
        RECT 2414.670 1607.305 2414.845 1608.565 ;
        RECT 2415.100 1608.445 2415.270 1610.045 ;
        RECT 2425.400 1609.935 2425.570 1610.105 ;
        RECT 2425.400 1609.605 2425.810 1609.935 ;
        RECT 2425.400 1609.095 2425.570 1609.605 ;
        RECT 2425.400 1608.765 2425.810 1609.095 ;
        RECT 2425.400 1608.565 2425.570 1608.765 ;
        RECT 2415.100 1607.305 2415.275 1608.445 ;
        RECT 2417.305 1607.560 2418.000 1608.190 ;
        RECT 2365.580 1605.980 2365.910 1606.960 ;
        RECT 2367.880 1605.980 2368.210 1606.960 ;
        RECT 2369.240 1605.980 2369.570 1606.960 ;
        RECT 2370.620 1605.980 2370.950 1606.960 ;
        RECT 2382.800 1605.980 2383.130 1606.960 ;
        RECT 2385.100 1605.980 2385.430 1606.960 ;
        RECT 2386.460 1605.980 2386.790 1606.960 ;
        RECT 2387.840 1605.980 2388.170 1606.960 ;
        RECT 2400.020 1605.985 2400.350 1606.965 ;
        RECT 2402.320 1605.985 2402.650 1606.965 ;
        RECT 2403.680 1605.985 2404.010 1606.965 ;
        RECT 2405.060 1605.985 2405.390 1606.965 ;
        RECT 2417.305 1606.960 2417.475 1607.560 ;
        RECT 2417.645 1607.340 2417.980 1607.370 ;
        RECT 2418.370 1607.340 2418.540 1608.020 ;
        RECT 2417.645 1607.170 2418.540 1607.340 ;
        RECT 2419.605 1607.560 2420.300 1608.190 ;
        RECT 2420.470 1607.560 2421.165 1608.190 ;
        RECT 2421.850 1607.560 2422.545 1608.190 ;
        RECT 2417.645 1607.120 2417.980 1607.170 ;
        RECT 2419.605 1606.960 2419.775 1607.560 ;
        RECT 2419.945 1607.340 2420.280 1607.370 ;
        RECT 2420.490 1607.340 2420.825 1607.370 ;
        RECT 2419.945 1607.170 2420.825 1607.340 ;
        RECT 2419.945 1607.120 2420.280 1607.170 ;
        RECT 2420.490 1607.120 2420.825 1607.170 ;
        RECT 2420.995 1606.960 2421.165 1607.560 ;
        RECT 2421.335 1607.120 2421.670 1607.390 ;
        RECT 2421.870 1607.120 2422.205 1607.370 ;
        RECT 2422.375 1606.960 2422.545 1607.560 ;
        RECT 2422.715 1607.120 2423.050 1607.390 ;
        RECT 2425.400 1607.305 2425.575 1608.565 ;
        RECT 2425.985 1608.535 2426.155 1610.145 ;
        RECT 2426.355 1610.085 2426.530 1610.595 ;
        RECT 2426.785 1610.045 2426.960 1610.595 ;
        RECT 2428.150 1610.085 2428.320 1610.595 ;
        RECT 2429.140 1610.085 2429.310 1610.595 ;
        RECT 2430.935 1610.105 2431.110 1610.595 ;
        RECT 2425.925 1608.365 2426.155 1608.535 ;
        RECT 2426.355 1608.565 2426.525 1609.515 ;
        RECT 2425.925 1607.305 2426.095 1608.365 ;
        RECT 2426.355 1607.305 2426.530 1608.565 ;
        RECT 2426.785 1608.445 2426.955 1610.045 ;
        RECT 2430.935 1609.935 2431.105 1610.105 ;
        RECT 2431.890 1610.085 2432.065 1610.595 ;
        RECT 2432.320 1610.045 2432.495 1610.595 ;
        RECT 2442.620 1610.105 2442.795 1610.595 ;
        RECT 2443.145 1610.315 2443.315 1610.595 ;
        RECT 2443.145 1610.145 2443.375 1610.315 ;
        RECT 2427.715 1609.425 2427.945 1609.615 ;
        RECT 2430.935 1609.605 2431.345 1609.935 ;
        RECT 2427.715 1609.385 2428.245 1609.425 ;
        RECT 2427.775 1609.255 2428.245 1609.385 ;
        RECT 2428.765 1609.255 2429.235 1609.425 ;
        RECT 2427.775 1608.565 2427.945 1609.255 ;
        RECT 2428.145 1608.780 2428.315 1608.885 ;
        RECT 2428.765 1608.780 2428.935 1609.255 ;
        RECT 2430.935 1609.095 2431.105 1609.605 ;
        RECT 2428.145 1608.605 2428.935 1608.780 ;
        RECT 2426.785 1607.305 2426.960 1608.445 ;
        RECT 2428.145 1607.305 2428.320 1608.605 ;
        RECT 2428.765 1608.565 2428.935 1608.605 ;
        RECT 2429.135 1608.450 2429.305 1608.885 ;
        RECT 2430.935 1608.765 2431.345 1609.095 ;
        RECT 2430.935 1608.565 2431.105 1608.765 ;
        RECT 2431.890 1608.565 2432.060 1609.515 ;
        RECT 2429.135 1607.305 2429.310 1608.450 ;
        RECT 2430.935 1607.305 2431.110 1608.565 ;
        RECT 2431.890 1607.305 2432.065 1608.565 ;
        RECT 2432.320 1608.445 2432.490 1610.045 ;
        RECT 2442.620 1609.935 2442.790 1610.105 ;
        RECT 2442.620 1609.605 2443.030 1609.935 ;
        RECT 2442.620 1609.095 2442.790 1609.605 ;
        RECT 2442.620 1608.765 2443.030 1609.095 ;
        RECT 2442.620 1608.565 2442.790 1608.765 ;
        RECT 2432.320 1607.305 2432.495 1608.445 ;
        RECT 2434.525 1607.560 2435.220 1608.190 ;
        RECT 2434.525 1606.960 2434.695 1607.560 ;
        RECT 2434.865 1607.340 2435.200 1607.370 ;
        RECT 2435.590 1607.340 2435.760 1608.020 ;
        RECT 2434.865 1607.170 2435.760 1607.340 ;
        RECT 2436.825 1607.560 2437.520 1608.190 ;
        RECT 2437.690 1607.560 2438.385 1608.190 ;
        RECT 2439.070 1607.560 2439.765 1608.190 ;
        RECT 2434.865 1607.120 2435.200 1607.170 ;
        RECT 2436.825 1606.960 2436.995 1607.560 ;
        RECT 2437.165 1607.340 2437.500 1607.370 ;
        RECT 2437.710 1607.340 2438.045 1607.370 ;
        RECT 2437.165 1607.170 2438.045 1607.340 ;
        RECT 2437.165 1607.120 2437.500 1607.170 ;
        RECT 2437.710 1607.120 2438.045 1607.170 ;
        RECT 2438.215 1606.960 2438.385 1607.560 ;
        RECT 2438.555 1607.120 2438.890 1607.390 ;
        RECT 2439.090 1607.120 2439.425 1607.370 ;
        RECT 2439.595 1606.960 2439.765 1607.560 ;
        RECT 2439.935 1607.120 2440.270 1607.390 ;
        RECT 2442.620 1607.305 2442.795 1608.565 ;
        RECT 2443.205 1608.535 2443.375 1610.145 ;
        RECT 2443.575 1610.085 2443.750 1610.595 ;
        RECT 2444.005 1610.045 2444.180 1610.595 ;
        RECT 2445.370 1610.085 2445.540 1610.595 ;
        RECT 2446.360 1610.085 2446.530 1610.595 ;
        RECT 2697.910 1610.315 2698.245 1610.565 ;
        RECT 2698.415 1610.315 2699.130 1610.645 ;
        RECT 2699.345 1610.315 2700.170 1610.645 ;
        RECT 2700.340 1610.315 2700.615 1610.645 ;
        RECT 2443.145 1608.365 2443.375 1608.535 ;
        RECT 2443.575 1608.565 2443.745 1609.515 ;
        RECT 2443.145 1607.305 2443.315 1608.365 ;
        RECT 2443.575 1607.305 2443.750 1608.565 ;
        RECT 2444.005 1608.445 2444.175 1610.045 ;
        RECT 2698.415 1609.755 2698.585 1610.315 ;
        RECT 2698.845 1609.855 2699.175 1610.145 ;
        RECT 2699.345 1610.025 2699.590 1610.315 ;
        RECT 2700.340 1610.145 2700.510 1610.315 ;
        RECT 2700.785 1610.145 2700.955 1610.880 ;
        RECT 2699.850 1609.975 2700.510 1610.145 ;
        RECT 2699.850 1609.855 2700.020 1609.975 ;
        RECT 2698.845 1609.685 2700.020 1609.855 ;
        RECT 2444.935 1609.425 2445.165 1609.615 ;
        RECT 2444.935 1609.385 2445.465 1609.425 ;
        RECT 2444.995 1609.255 2445.465 1609.385 ;
        RECT 2445.985 1609.255 2446.455 1609.425 ;
        RECT 2444.995 1608.565 2445.165 1609.255 ;
        RECT 2445.365 1608.780 2445.535 1608.885 ;
        RECT 2445.985 1608.780 2446.155 1609.255 ;
        RECT 2698.405 1609.185 2700.020 1609.515 ;
        RECT 2700.680 1609.175 2700.955 1610.145 ;
        RECT 2701.125 1611.155 2701.715 1611.385 ;
        RECT 2701.125 1610.145 2701.415 1611.155 ;
        RECT 2703.290 1610.985 2703.715 1611.195 ;
        RECT 2701.585 1610.815 2703.715 1610.985 ;
        RECT 2701.585 1610.315 2701.755 1610.815 ;
        RECT 2702.045 1610.315 2702.375 1610.645 ;
        RECT 2702.565 1610.315 2702.835 1610.645 ;
        RECT 2703.025 1610.315 2703.375 1610.645 ;
        RECT 2701.125 1609.975 2702.670 1610.145 ;
        RECT 2703.545 1610.045 2703.715 1610.815 ;
        RECT 2701.125 1609.175 2701.715 1609.975 ;
        RECT 2702.340 1609.175 2702.670 1609.975 ;
        RECT 2703.290 1609.715 2703.715 1610.045 ;
        RECT 2445.365 1608.605 2446.155 1608.780 ;
        RECT 2444.005 1607.305 2444.180 1608.445 ;
        RECT 2445.365 1607.305 2445.540 1608.605 ;
        RECT 2445.985 1608.565 2446.155 1608.605 ;
        RECT 2446.355 1608.450 2446.525 1608.885 ;
        RECT 2446.355 1607.305 2446.530 1608.450 ;
        RECT 2697.075 1607.905 2697.245 1608.665 ;
        RECT 2697.075 1607.735 2697.740 1607.905 ;
        RECT 2697.925 1607.760 2698.195 1608.665 ;
        RECT 2697.570 1607.590 2697.740 1607.735 ;
        RECT 2697.005 1607.185 2697.335 1607.555 ;
        RECT 2697.570 1607.260 2697.855 1607.590 ;
        RECT 2697.570 1607.005 2697.740 1607.260 ;
        RECT 2417.240 1605.980 2417.570 1606.960 ;
        RECT 2419.540 1605.980 2419.870 1606.960 ;
        RECT 2420.900 1605.980 2421.230 1606.960 ;
        RECT 2422.280 1605.980 2422.610 1606.960 ;
        RECT 2434.460 1605.980 2434.790 1606.960 ;
        RECT 2436.760 1605.980 2437.090 1606.960 ;
        RECT 2438.120 1605.980 2438.450 1606.960 ;
        RECT 2439.500 1605.980 2439.830 1606.960 ;
        RECT 2697.075 1606.835 2697.740 1607.005 ;
        RECT 2698.025 1606.960 2698.195 1607.760 ;
        RECT 2699.255 1607.685 2699.585 1608.665 ;
        RECT 2698.845 1607.275 2699.180 1607.525 ;
        RECT 2699.350 1607.085 2699.520 1607.685 ;
        RECT 2699.690 1607.255 2700.025 1607.525 ;
        RECT 2697.075 1606.455 2697.245 1606.835 ;
        RECT 2697.935 1606.455 2698.195 1606.960 ;
        RECT 2698.825 1606.455 2699.520 1607.085 ;
        RECT 2365.110 1604.490 2365.440 1605.470 ;
        RECT 2366.920 1604.670 2367.250 1605.455 ;
        RECT 2366.570 1604.500 2367.250 1604.670 ;
        RECT 2367.440 1604.670 2367.770 1605.455 ;
        RECT 2367.440 1604.500 2368.120 1604.670 ;
        RECT 2365.110 1603.890 2365.360 1604.490 ;
        RECT 2365.530 1604.280 2365.860 1604.330 ;
        RECT 2366.050 1604.280 2366.400 1604.330 ;
        RECT 2365.530 1604.110 2366.400 1604.280 ;
        RECT 2365.530 1604.080 2365.860 1604.110 ;
        RECT 2366.050 1604.080 2366.400 1604.110 ;
        RECT 2366.570 1603.900 2366.740 1604.500 ;
        RECT 2366.910 1604.080 2367.260 1604.330 ;
        RECT 2367.430 1604.080 2367.780 1604.330 ;
        RECT 2367.950 1603.900 2368.120 1604.500 ;
        RECT 2368.810 1604.620 2369.130 1605.470 ;
        RECT 2369.310 1604.960 2369.710 1605.470 ;
        RECT 2370.220 1604.960 2370.550 1605.470 ;
        RECT 2369.310 1604.790 2370.550 1604.960 ;
        RECT 2371.130 1604.620 2371.300 1605.300 ;
        RECT 2371.480 1604.790 2371.860 1605.470 ;
        RECT 2368.810 1604.540 2369.260 1604.620 ;
        RECT 2368.810 1604.370 2369.440 1604.540 ;
        RECT 2368.290 1604.080 2368.640 1604.330 ;
        RECT 2365.110 1603.260 2365.440 1603.890 ;
        RECT 2366.500 1603.260 2366.830 1603.900 ;
        RECT 2367.860 1603.260 2368.190 1603.900 ;
        RECT 2369.270 1603.490 2369.440 1604.370 ;
        RECT 2370.215 1604.450 2371.520 1604.620 ;
        RECT 2369.610 1603.830 2369.840 1604.330 ;
        RECT 2370.215 1604.250 2370.385 1604.450 ;
        RECT 2370.010 1604.080 2370.385 1604.250 ;
        RECT 2370.555 1604.080 2371.105 1604.280 ;
        RECT 2371.275 1604.000 2371.520 1604.450 ;
        RECT 2371.690 1603.830 2371.860 1604.790 ;
        RECT 2369.610 1603.660 2371.860 1603.830 ;
        RECT 2373.740 1603.895 2373.915 1605.155 ;
        RECT 2374.265 1604.095 2374.435 1605.155 ;
        RECT 2374.265 1603.925 2374.495 1604.095 ;
        RECT 2373.740 1603.695 2373.910 1603.895 ;
        RECT 2369.270 1603.320 2370.225 1603.490 ;
        RECT 2371.140 1603.340 2371.310 1603.660 ;
        RECT 2373.740 1603.365 2374.150 1603.695 ;
        RECT 2373.740 1602.855 2373.910 1603.365 ;
        RECT 2373.740 1602.525 2374.150 1602.855 ;
        RECT 2373.740 1602.355 2373.910 1602.525 ;
        RECT 2373.740 1601.865 2373.915 1602.355 ;
        RECT 2374.325 1602.315 2374.495 1603.925 ;
        RECT 2374.695 1603.895 2374.870 1605.155 ;
        RECT 2375.125 1604.015 2375.300 1605.155 ;
        RECT 2374.695 1602.945 2374.865 1603.895 ;
        RECT 2375.125 1602.415 2375.295 1604.015 ;
        RECT 2376.485 1604.010 2376.660 1605.155 ;
        RECT 2377.470 1604.010 2377.645 1605.155 ;
        RECT 2382.330 1604.490 2382.660 1605.470 ;
        RECT 2384.140 1604.670 2384.470 1605.455 ;
        RECT 2383.790 1604.500 2384.470 1604.670 ;
        RECT 2384.660 1604.670 2384.990 1605.455 ;
        RECT 2384.660 1604.500 2385.340 1604.670 ;
        RECT 2376.115 1603.205 2376.285 1603.895 ;
        RECT 2376.485 1603.805 2376.655 1604.010 ;
        RECT 2377.100 1603.805 2377.270 1603.895 ;
        RECT 2376.485 1603.625 2377.270 1603.805 ;
        RECT 2376.485 1603.575 2376.655 1603.625 ;
        RECT 2377.100 1603.205 2377.270 1603.625 ;
        RECT 2377.470 1603.575 2377.640 1604.010 ;
        RECT 2382.330 1603.890 2382.580 1604.490 ;
        RECT 2382.750 1604.280 2383.080 1604.330 ;
        RECT 2383.270 1604.280 2383.620 1604.330 ;
        RECT 2382.750 1604.110 2383.620 1604.280 ;
        RECT 2382.750 1604.080 2383.080 1604.110 ;
        RECT 2383.270 1604.080 2383.620 1604.110 ;
        RECT 2383.790 1603.900 2383.960 1604.500 ;
        RECT 2384.130 1604.080 2384.480 1604.330 ;
        RECT 2384.650 1604.080 2385.000 1604.330 ;
        RECT 2385.170 1603.900 2385.340 1604.500 ;
        RECT 2386.030 1604.620 2386.350 1605.470 ;
        RECT 2386.530 1604.960 2386.930 1605.470 ;
        RECT 2387.440 1604.960 2387.770 1605.470 ;
        RECT 2386.530 1604.790 2387.770 1604.960 ;
        RECT 2388.350 1604.620 2388.520 1605.300 ;
        RECT 2388.700 1604.790 2389.080 1605.470 ;
        RECT 2386.030 1604.540 2386.480 1604.620 ;
        RECT 2386.030 1604.370 2386.660 1604.540 ;
        RECT 2385.510 1604.080 2385.860 1604.330 ;
        RECT 2382.330 1603.260 2382.660 1603.890 ;
        RECT 2383.720 1603.260 2384.050 1603.900 ;
        RECT 2385.080 1603.260 2385.410 1603.900 ;
        RECT 2386.490 1603.490 2386.660 1604.370 ;
        RECT 2387.435 1604.450 2388.740 1604.620 ;
        RECT 2386.830 1603.830 2387.060 1604.330 ;
        RECT 2387.435 1604.250 2387.605 1604.450 ;
        RECT 2387.230 1604.080 2387.605 1604.250 ;
        RECT 2387.775 1604.080 2388.325 1604.280 ;
        RECT 2388.495 1604.000 2388.740 1604.450 ;
        RECT 2388.910 1603.830 2389.080 1604.790 ;
        RECT 2386.830 1603.660 2389.080 1603.830 ;
        RECT 2390.960 1603.895 2391.135 1605.155 ;
        RECT 2391.485 1604.095 2391.655 1605.155 ;
        RECT 2391.485 1603.925 2391.715 1604.095 ;
        RECT 2390.960 1603.695 2391.130 1603.895 ;
        RECT 2386.490 1603.320 2387.445 1603.490 ;
        RECT 2388.360 1603.340 2388.530 1603.660 ;
        RECT 2390.960 1603.365 2391.370 1603.695 ;
        RECT 2376.115 1603.175 2376.585 1603.205 ;
        RECT 2376.030 1603.035 2376.585 1603.175 ;
        RECT 2377.100 1603.035 2377.570 1603.205 ;
        RECT 2376.030 1602.945 2376.260 1603.035 ;
        RECT 2390.960 1602.855 2391.130 1603.365 ;
        RECT 2390.960 1602.525 2391.370 1602.855 ;
        RECT 2374.265 1602.145 2374.495 1602.315 ;
        RECT 2374.265 1601.865 2374.435 1602.145 ;
        RECT 2374.695 1601.865 2374.870 1602.375 ;
        RECT 2375.125 1601.865 2375.300 1602.415 ;
        RECT 2376.490 1601.865 2376.660 1602.375 ;
        RECT 2377.475 1601.865 2377.645 1602.375 ;
        RECT 2390.960 1602.355 2391.130 1602.525 ;
        RECT 2390.960 1601.865 2391.135 1602.355 ;
        RECT 2391.545 1602.315 2391.715 1603.925 ;
        RECT 2391.915 1603.895 2392.090 1605.155 ;
        RECT 2392.345 1604.015 2392.520 1605.155 ;
        RECT 2391.915 1602.945 2392.085 1603.895 ;
        RECT 2392.345 1602.415 2392.515 1604.015 ;
        RECT 2393.705 1604.010 2393.880 1605.155 ;
        RECT 2394.690 1604.010 2394.865 1605.155 ;
        RECT 2399.550 1604.495 2399.880 1605.475 ;
        RECT 2401.360 1604.675 2401.690 1605.460 ;
        RECT 2401.010 1604.505 2401.690 1604.675 ;
        RECT 2401.880 1604.675 2402.210 1605.460 ;
        RECT 2401.880 1604.505 2402.560 1604.675 ;
        RECT 2393.335 1603.205 2393.505 1603.895 ;
        RECT 2393.705 1603.805 2393.875 1604.010 ;
        RECT 2394.320 1603.805 2394.490 1603.895 ;
        RECT 2393.705 1603.625 2394.490 1603.805 ;
        RECT 2393.705 1603.575 2393.875 1603.625 ;
        RECT 2394.320 1603.205 2394.490 1603.625 ;
        RECT 2394.690 1603.575 2394.860 1604.010 ;
        RECT 2399.550 1603.895 2399.800 1604.495 ;
        RECT 2399.970 1604.285 2400.300 1604.335 ;
        RECT 2400.490 1604.285 2400.840 1604.335 ;
        RECT 2399.970 1604.115 2400.840 1604.285 ;
        RECT 2399.970 1604.085 2400.300 1604.115 ;
        RECT 2400.490 1604.085 2400.840 1604.115 ;
        RECT 2401.010 1603.905 2401.180 1604.505 ;
        RECT 2401.350 1604.085 2401.700 1604.335 ;
        RECT 2401.870 1604.085 2402.220 1604.335 ;
        RECT 2402.390 1603.905 2402.560 1604.505 ;
        RECT 2403.250 1604.625 2403.570 1605.475 ;
        RECT 2403.750 1604.965 2404.150 1605.475 ;
        RECT 2404.660 1604.965 2404.990 1605.475 ;
        RECT 2403.750 1604.795 2404.990 1604.965 ;
        RECT 2405.570 1604.625 2405.740 1605.305 ;
        RECT 2405.920 1604.795 2406.300 1605.475 ;
        RECT 2403.250 1604.545 2403.700 1604.625 ;
        RECT 2403.250 1604.375 2403.880 1604.545 ;
        RECT 2402.730 1604.085 2403.080 1604.335 ;
        RECT 2399.550 1603.265 2399.880 1603.895 ;
        RECT 2400.940 1603.265 2401.270 1603.905 ;
        RECT 2402.300 1603.265 2402.630 1603.905 ;
        RECT 2403.710 1603.495 2403.880 1604.375 ;
        RECT 2404.655 1604.455 2405.960 1604.625 ;
        RECT 2404.050 1603.835 2404.280 1604.335 ;
        RECT 2404.655 1604.255 2404.825 1604.455 ;
        RECT 2404.450 1604.085 2404.825 1604.255 ;
        RECT 2404.995 1604.085 2405.545 1604.285 ;
        RECT 2405.715 1604.005 2405.960 1604.455 ;
        RECT 2406.130 1603.835 2406.300 1604.795 ;
        RECT 2404.050 1603.665 2406.300 1603.835 ;
        RECT 2408.180 1603.900 2408.355 1605.160 ;
        RECT 2408.705 1604.100 2408.875 1605.160 ;
        RECT 2408.705 1603.930 2408.935 1604.100 ;
        RECT 2408.180 1603.700 2408.350 1603.900 ;
        RECT 2403.710 1603.325 2404.665 1603.495 ;
        RECT 2405.580 1603.345 2405.750 1603.665 ;
        RECT 2408.180 1603.370 2408.590 1603.700 ;
        RECT 2393.335 1603.175 2393.805 1603.205 ;
        RECT 2393.250 1603.035 2393.805 1603.175 ;
        RECT 2394.320 1603.035 2394.790 1603.205 ;
        RECT 2393.250 1602.945 2393.480 1603.035 ;
        RECT 2408.180 1602.860 2408.350 1603.370 ;
        RECT 2408.180 1602.530 2408.590 1602.860 ;
        RECT 2391.485 1602.145 2391.715 1602.315 ;
        RECT 2391.485 1601.865 2391.655 1602.145 ;
        RECT 2391.915 1601.865 2392.090 1602.375 ;
        RECT 2392.345 1601.865 2392.520 1602.415 ;
        RECT 2393.710 1601.865 2393.880 1602.375 ;
        RECT 2394.695 1601.825 2394.865 1602.375 ;
        RECT 2408.180 1602.360 2408.350 1602.530 ;
        RECT 2408.180 1601.870 2408.355 1602.360 ;
        RECT 2408.765 1602.320 2408.935 1603.930 ;
        RECT 2409.135 1603.900 2409.310 1605.160 ;
        RECT 2409.565 1604.020 2409.740 1605.160 ;
        RECT 2409.135 1602.950 2409.305 1603.900 ;
        RECT 2409.565 1602.420 2409.735 1604.020 ;
        RECT 2410.925 1604.015 2411.100 1605.160 ;
        RECT 2411.910 1604.015 2412.085 1605.160 ;
        RECT 2416.770 1604.490 2417.100 1605.470 ;
        RECT 2418.580 1604.670 2418.910 1605.455 ;
        RECT 2418.230 1604.500 2418.910 1604.670 ;
        RECT 2419.100 1604.670 2419.430 1605.455 ;
        RECT 2419.100 1604.500 2419.780 1604.670 ;
        RECT 2410.555 1603.210 2410.725 1603.900 ;
        RECT 2410.925 1603.810 2411.095 1604.015 ;
        RECT 2411.540 1603.810 2411.710 1603.900 ;
        RECT 2410.925 1603.630 2411.710 1603.810 ;
        RECT 2410.925 1603.580 2411.095 1603.630 ;
        RECT 2411.540 1603.210 2411.710 1603.630 ;
        RECT 2411.910 1603.580 2412.080 1604.015 ;
        RECT 2416.770 1603.890 2417.020 1604.490 ;
        RECT 2417.190 1604.280 2417.520 1604.330 ;
        RECT 2417.710 1604.280 2418.060 1604.330 ;
        RECT 2417.190 1604.110 2418.060 1604.280 ;
        RECT 2417.190 1604.080 2417.520 1604.110 ;
        RECT 2417.710 1604.080 2418.060 1604.110 ;
        RECT 2418.230 1603.900 2418.400 1604.500 ;
        RECT 2418.570 1604.080 2418.920 1604.330 ;
        RECT 2419.090 1604.080 2419.440 1604.330 ;
        RECT 2419.610 1603.900 2419.780 1604.500 ;
        RECT 2420.470 1604.620 2420.790 1605.470 ;
        RECT 2420.970 1604.960 2421.370 1605.470 ;
        RECT 2421.880 1604.960 2422.210 1605.470 ;
        RECT 2420.970 1604.790 2422.210 1604.960 ;
        RECT 2422.790 1604.620 2422.960 1605.300 ;
        RECT 2423.140 1604.790 2423.520 1605.470 ;
        RECT 2420.470 1604.540 2420.920 1604.620 ;
        RECT 2420.470 1604.370 2421.100 1604.540 ;
        RECT 2419.950 1604.080 2420.300 1604.330 ;
        RECT 2416.770 1603.260 2417.100 1603.890 ;
        RECT 2418.160 1603.260 2418.490 1603.900 ;
        RECT 2419.520 1603.260 2419.850 1603.900 ;
        RECT 2420.930 1603.490 2421.100 1604.370 ;
        RECT 2421.875 1604.450 2423.180 1604.620 ;
        RECT 2421.270 1603.830 2421.500 1604.330 ;
        RECT 2421.875 1604.250 2422.045 1604.450 ;
        RECT 2421.670 1604.080 2422.045 1604.250 ;
        RECT 2422.215 1604.080 2422.765 1604.280 ;
        RECT 2422.935 1604.000 2423.180 1604.450 ;
        RECT 2423.350 1603.830 2423.520 1604.790 ;
        RECT 2421.270 1603.660 2423.520 1603.830 ;
        RECT 2425.400 1603.895 2425.575 1605.155 ;
        RECT 2425.925 1604.095 2426.095 1605.155 ;
        RECT 2425.925 1603.925 2426.155 1604.095 ;
        RECT 2425.400 1603.695 2425.570 1603.895 ;
        RECT 2420.930 1603.320 2421.885 1603.490 ;
        RECT 2422.800 1603.340 2422.970 1603.660 ;
        RECT 2425.400 1603.365 2425.810 1603.695 ;
        RECT 2410.555 1603.180 2411.025 1603.210 ;
        RECT 2410.470 1603.040 2411.025 1603.180 ;
        RECT 2411.540 1603.040 2412.010 1603.210 ;
        RECT 2410.470 1602.950 2410.700 1603.040 ;
        RECT 2425.400 1602.855 2425.570 1603.365 ;
        RECT 2425.400 1602.525 2425.810 1602.855 ;
        RECT 2408.705 1602.150 2408.935 1602.320 ;
        RECT 2408.705 1601.870 2408.875 1602.150 ;
        RECT 2409.135 1601.870 2409.310 1602.380 ;
        RECT 2409.565 1601.870 2409.740 1602.420 ;
        RECT 2410.930 1601.870 2411.100 1602.380 ;
        RECT 2411.915 1601.870 2412.085 1602.380 ;
        RECT 2425.400 1602.355 2425.570 1602.525 ;
        RECT 2425.400 1601.865 2425.575 1602.355 ;
        RECT 2425.985 1602.315 2426.155 1603.925 ;
        RECT 2426.355 1603.895 2426.530 1605.155 ;
        RECT 2426.785 1604.015 2426.960 1605.155 ;
        RECT 2426.355 1602.945 2426.525 1603.895 ;
        RECT 2426.785 1602.415 2426.955 1604.015 ;
        RECT 2428.145 1604.010 2428.320 1605.155 ;
        RECT 2429.130 1604.010 2429.305 1605.155 ;
        RECT 2433.990 1604.490 2434.320 1605.470 ;
        RECT 2435.800 1604.670 2436.130 1605.455 ;
        RECT 2435.450 1604.500 2436.130 1604.670 ;
        RECT 2436.320 1604.670 2436.650 1605.455 ;
        RECT 2436.320 1604.500 2437.000 1604.670 ;
        RECT 2427.775 1603.205 2427.945 1603.895 ;
        RECT 2428.145 1603.805 2428.315 1604.010 ;
        RECT 2428.760 1603.805 2428.930 1603.895 ;
        RECT 2428.145 1603.625 2428.930 1603.805 ;
        RECT 2428.145 1603.575 2428.315 1603.625 ;
        RECT 2428.760 1603.205 2428.930 1603.625 ;
        RECT 2429.130 1603.575 2429.300 1604.010 ;
        RECT 2433.990 1603.890 2434.240 1604.490 ;
        RECT 2434.410 1604.280 2434.740 1604.330 ;
        RECT 2434.930 1604.280 2435.280 1604.330 ;
        RECT 2434.410 1604.110 2435.280 1604.280 ;
        RECT 2434.410 1604.080 2434.740 1604.110 ;
        RECT 2434.930 1604.080 2435.280 1604.110 ;
        RECT 2435.450 1603.900 2435.620 1604.500 ;
        RECT 2435.790 1604.080 2436.140 1604.330 ;
        RECT 2436.310 1604.080 2436.660 1604.330 ;
        RECT 2436.830 1603.900 2437.000 1604.500 ;
        RECT 2437.690 1604.620 2438.010 1605.470 ;
        RECT 2438.190 1604.960 2438.590 1605.470 ;
        RECT 2439.100 1604.960 2439.430 1605.470 ;
        RECT 2438.190 1604.790 2439.430 1604.960 ;
        RECT 2440.010 1604.620 2440.180 1605.300 ;
        RECT 2440.360 1604.790 2440.740 1605.470 ;
        RECT 2697.260 1605.305 2697.505 1605.910 ;
        RECT 2437.690 1604.540 2438.140 1604.620 ;
        RECT 2437.690 1604.370 2438.320 1604.540 ;
        RECT 2437.170 1604.080 2437.520 1604.330 ;
        RECT 2433.990 1603.260 2434.320 1603.890 ;
        RECT 2435.380 1603.260 2435.710 1603.900 ;
        RECT 2436.740 1603.260 2437.070 1603.900 ;
        RECT 2438.150 1603.490 2438.320 1604.370 ;
        RECT 2439.095 1604.450 2440.400 1604.620 ;
        RECT 2438.490 1603.830 2438.720 1604.330 ;
        RECT 2439.095 1604.250 2439.265 1604.450 ;
        RECT 2438.890 1604.080 2439.265 1604.250 ;
        RECT 2439.435 1604.080 2439.985 1604.280 ;
        RECT 2440.155 1604.000 2440.400 1604.450 ;
        RECT 2440.570 1603.830 2440.740 1604.790 ;
        RECT 2438.490 1603.660 2440.740 1603.830 ;
        RECT 2442.620 1603.895 2442.795 1605.155 ;
        RECT 2443.145 1604.095 2443.315 1605.155 ;
        RECT 2443.145 1603.925 2443.375 1604.095 ;
        RECT 2442.620 1603.695 2442.790 1603.895 ;
        RECT 2438.150 1603.320 2439.105 1603.490 ;
        RECT 2440.020 1603.340 2440.190 1603.660 ;
        RECT 2442.620 1603.365 2443.030 1603.695 ;
        RECT 2427.775 1603.175 2428.245 1603.205 ;
        RECT 2427.690 1603.035 2428.245 1603.175 ;
        RECT 2428.760 1603.035 2429.230 1603.205 ;
        RECT 2427.690 1602.945 2427.920 1603.035 ;
        RECT 2442.620 1602.855 2442.790 1603.365 ;
        RECT 2442.620 1602.525 2443.030 1602.855 ;
        RECT 2425.925 1602.145 2426.155 1602.315 ;
        RECT 2425.925 1601.865 2426.095 1602.145 ;
        RECT 2426.355 1601.865 2426.530 1602.375 ;
        RECT 2426.785 1601.865 2426.960 1602.415 ;
        RECT 2428.150 1601.865 2428.320 1602.375 ;
        RECT 2429.135 1601.825 2429.305 1602.375 ;
        RECT 2442.620 1602.355 2442.790 1602.525 ;
        RECT 2442.620 1601.865 2442.795 1602.355 ;
        RECT 2443.205 1602.315 2443.375 1603.925 ;
        RECT 2443.575 1603.895 2443.750 1605.155 ;
        RECT 2444.005 1604.015 2444.180 1605.155 ;
        RECT 2443.575 1602.945 2443.745 1603.895 ;
        RECT 2444.005 1602.415 2444.175 1604.015 ;
        RECT 2445.365 1604.010 2445.540 1605.155 ;
        RECT 2446.350 1604.010 2446.525 1605.155 ;
        RECT 2696.985 1605.135 2698.215 1605.305 ;
        RECT 2696.985 1604.325 2697.325 1605.135 ;
        RECT 2697.495 1604.570 2698.245 1604.760 ;
        RECT 2444.995 1603.205 2445.165 1603.895 ;
        RECT 2445.365 1603.805 2445.535 1604.010 ;
        RECT 2445.980 1603.805 2446.150 1603.895 ;
        RECT 2445.365 1603.625 2446.150 1603.805 ;
        RECT 2445.365 1603.575 2445.535 1603.625 ;
        RECT 2445.980 1603.205 2446.150 1603.625 ;
        RECT 2446.350 1603.575 2446.520 1604.010 ;
        RECT 2696.985 1603.915 2697.500 1604.325 ;
        RECT 2698.075 1603.905 2698.245 1604.570 ;
        RECT 2698.415 1604.585 2698.605 1605.945 ;
        RECT 2698.775 1605.095 2699.050 1605.945 ;
        RECT 2699.240 1605.580 2699.770 1605.945 ;
        RECT 2699.595 1605.545 2699.770 1605.580 ;
        RECT 2698.775 1604.925 2699.055 1605.095 ;
        RECT 2698.775 1604.785 2699.050 1604.925 ;
        RECT 2699.255 1604.585 2699.425 1605.385 ;
        RECT 2698.415 1604.415 2699.425 1604.585 ;
        RECT 2699.595 1605.375 2700.525 1605.545 ;
        RECT 2700.695 1605.375 2700.950 1605.945 ;
        RECT 2699.595 1604.245 2699.765 1605.375 ;
        RECT 2700.355 1605.205 2700.525 1605.375 ;
        RECT 2698.640 1604.075 2699.765 1604.245 ;
        RECT 2699.935 1604.875 2700.130 1605.205 ;
        RECT 2700.355 1604.875 2700.610 1605.205 ;
        RECT 2699.935 1603.905 2700.105 1604.875 ;
        RECT 2700.780 1604.705 2700.950 1605.375 ;
        RECT 2698.075 1603.735 2700.105 1603.905 ;
        RECT 2700.615 1603.735 2700.950 1604.705 ;
        RECT 2444.995 1603.175 2445.465 1603.205 ;
        RECT 2444.910 1603.035 2445.465 1603.175 ;
        RECT 2445.980 1603.035 2446.450 1603.205 ;
        RECT 2444.910 1602.945 2445.140 1603.035 ;
        RECT 2697.075 1602.465 2697.245 1603.225 ;
        RECT 2443.145 1602.145 2443.375 1602.315 ;
        RECT 2443.145 1601.865 2443.315 1602.145 ;
        RECT 2443.575 1601.865 2443.750 1602.375 ;
        RECT 2444.005 1601.865 2444.180 1602.415 ;
        RECT 2445.370 1601.865 2445.540 1602.375 ;
        RECT 2446.355 1601.865 2446.525 1602.375 ;
        RECT 2697.075 1602.295 2697.740 1602.465 ;
        RECT 2697.925 1602.320 2698.195 1603.225 ;
        RECT 2697.570 1602.150 2697.740 1602.295 ;
        RECT 2697.005 1601.745 2697.335 1602.115 ;
        RECT 2697.570 1601.820 2697.855 1602.150 ;
        RECT 2697.570 1601.565 2697.740 1601.820 ;
        RECT 2697.075 1601.395 2697.740 1601.565 ;
        RECT 2698.025 1601.520 2698.195 1602.320 ;
        RECT 2697.075 1601.015 2697.245 1601.395 ;
        RECT 2697.935 1601.015 2698.195 1601.520 ;
        RECT 2697.075 1597.025 2697.245 1597.785 ;
        RECT 2697.075 1596.855 2697.740 1597.025 ;
        RECT 2697.925 1596.880 2698.195 1597.785 ;
        RECT 2697.570 1596.710 2697.740 1596.855 ;
        RECT 2697.005 1596.305 2697.335 1596.675 ;
        RECT 2697.570 1596.380 2697.855 1596.710 ;
        RECT 2697.570 1596.125 2697.740 1596.380 ;
        RECT 2697.075 1595.955 2697.740 1596.125 ;
        RECT 2698.025 1596.080 2698.195 1596.880 ;
        RECT 2697.075 1595.575 2697.245 1595.955 ;
        RECT 2697.935 1595.575 2698.195 1596.080 ;
        RECT 2697.075 1591.585 2697.245 1592.345 ;
        RECT 2697.075 1591.415 2697.740 1591.585 ;
        RECT 2697.925 1591.440 2698.195 1592.345 ;
        RECT 2697.570 1591.270 2697.740 1591.415 ;
        RECT 2697.005 1590.865 2697.335 1591.235 ;
        RECT 2697.570 1590.940 2697.855 1591.270 ;
        RECT 2697.570 1590.685 2697.740 1590.940 ;
        RECT 2697.075 1590.515 2697.740 1590.685 ;
        RECT 2698.025 1590.640 2698.195 1591.440 ;
        RECT 2698.455 1591.585 2698.625 1592.345 ;
        RECT 2698.455 1591.415 2699.120 1591.585 ;
        RECT 2699.305 1591.440 2699.575 1592.345 ;
        RECT 2698.950 1591.270 2699.120 1591.415 ;
        RECT 2698.385 1590.865 2698.715 1591.235 ;
        RECT 2698.950 1590.940 2699.235 1591.270 ;
        RECT 2698.950 1590.685 2699.120 1590.940 ;
        RECT 2522.640 1588.190 2523.160 1589.675 ;
        RECT 2523.330 1588.850 2523.850 1590.400 ;
        RECT 2697.075 1590.135 2697.245 1590.515 ;
        RECT 2697.935 1590.135 2698.195 1590.640 ;
        RECT 2698.455 1590.515 2699.120 1590.685 ;
        RECT 2699.405 1590.640 2699.575 1591.440 ;
        RECT 2698.455 1590.135 2698.625 1590.515 ;
        RECT 2699.315 1590.135 2699.575 1590.640 ;
        RECT 2522.640 1580.660 2523.160 1582.145 ;
        RECT 2523.330 1581.320 2523.850 1582.870 ;
        RECT 2522.640 1574.680 2523.160 1576.165 ;
        RECT 2523.330 1575.340 2523.850 1576.890 ;
        RECT 2522.640 1566.265 2523.160 1567.750 ;
        RECT 2523.330 1566.925 2523.850 1568.475 ;
        RECT 2358.645 1533.105 2358.820 1533.595 ;
        RECT 2359.170 1533.315 2359.340 1533.595 ;
        RECT 2359.170 1533.145 2359.400 1533.315 ;
        RECT 2358.645 1532.935 2358.815 1533.105 ;
        RECT 2358.645 1532.605 2359.055 1532.935 ;
        RECT 2358.645 1532.095 2358.815 1532.605 ;
        RECT 2358.645 1531.765 2359.055 1532.095 ;
        RECT 2358.645 1531.565 2358.815 1531.765 ;
        RECT 2358.645 1530.305 2358.820 1531.565 ;
        RECT 2359.230 1531.535 2359.400 1533.145 ;
        RECT 2359.600 1533.085 2359.775 1533.595 ;
        RECT 2367.225 1533.105 2367.400 1533.595 ;
        RECT 2367.225 1532.935 2367.395 1533.105 ;
        RECT 2368.180 1533.085 2368.355 1533.595 ;
        RECT 2368.610 1533.045 2368.785 1533.595 ;
        RECT 2372.840 1533.105 2373.015 1533.595 ;
        RECT 2373.365 1533.315 2373.535 1533.595 ;
        RECT 2373.365 1533.145 2373.595 1533.315 ;
        RECT 2367.225 1532.605 2367.635 1532.935 ;
        RECT 2359.170 1531.365 2359.400 1531.535 ;
        RECT 2359.600 1531.565 2359.770 1532.515 ;
        RECT 2367.225 1532.095 2367.395 1532.605 ;
        RECT 2367.225 1531.765 2367.635 1532.095 ;
        RECT 2367.225 1531.565 2367.395 1531.765 ;
        RECT 2368.180 1531.565 2368.350 1532.515 ;
        RECT 2359.170 1530.305 2359.340 1531.365 ;
        RECT 2359.600 1530.305 2359.775 1531.565 ;
        RECT 2367.225 1530.305 2367.400 1531.565 ;
        RECT 2368.180 1530.305 2368.355 1531.565 ;
        RECT 2368.610 1531.445 2368.780 1533.045 ;
        RECT 2372.840 1532.935 2373.010 1533.105 ;
        RECT 2372.840 1532.605 2373.250 1532.935 ;
        RECT 2372.840 1532.095 2373.010 1532.605 ;
        RECT 2372.840 1531.765 2373.250 1532.095 ;
        RECT 2372.840 1531.565 2373.010 1531.765 ;
        RECT 2368.610 1530.305 2368.785 1531.445 ;
        RECT 2372.840 1530.305 2373.015 1531.565 ;
        RECT 2373.425 1531.535 2373.595 1533.145 ;
        RECT 2373.795 1533.085 2373.970 1533.595 ;
        RECT 2374.225 1533.045 2374.400 1533.595 ;
        RECT 2375.590 1533.085 2375.760 1533.595 ;
        RECT 2376.585 1533.080 2376.755 1533.590 ;
        RECT 2383.550 1533.105 2383.725 1533.595 ;
        RECT 2373.365 1531.365 2373.595 1531.535 ;
        RECT 2373.795 1531.565 2373.965 1532.515 ;
        RECT 2373.365 1530.305 2373.535 1531.365 ;
        RECT 2373.795 1530.305 2373.970 1531.565 ;
        RECT 2374.225 1531.445 2374.395 1533.045 ;
        RECT 2383.550 1532.935 2383.720 1533.105 ;
        RECT 2384.505 1533.085 2384.680 1533.595 ;
        RECT 2384.935 1533.045 2385.110 1533.595 ;
        RECT 2389.165 1533.105 2389.340 1533.595 ;
        RECT 2389.690 1533.315 2389.860 1533.595 ;
        RECT 2389.690 1533.145 2389.920 1533.315 ;
        RECT 2383.550 1532.605 2383.960 1532.935 ;
        RECT 2374.765 1532.425 2374.995 1532.575 ;
        RECT 2374.765 1532.255 2375.685 1532.425 ;
        RECT 2375.215 1531.565 2375.385 1532.255 ;
        RECT 2376.210 1532.250 2376.680 1532.420 ;
        RECT 2375.585 1531.775 2375.755 1531.885 ;
        RECT 2376.210 1531.775 2376.380 1532.250 ;
        RECT 2383.550 1532.095 2383.720 1532.605 ;
        RECT 2375.585 1531.605 2376.380 1531.775 ;
        RECT 2374.225 1530.305 2374.400 1531.445 ;
        RECT 2375.585 1530.305 2375.760 1531.605 ;
        RECT 2376.210 1531.560 2376.380 1531.605 ;
        RECT 2376.580 1531.445 2376.750 1531.880 ;
        RECT 2383.550 1531.765 2383.960 1532.095 ;
        RECT 2383.550 1531.565 2383.720 1531.765 ;
        RECT 2384.505 1531.565 2384.675 1532.515 ;
        RECT 2376.580 1530.300 2376.755 1531.445 ;
        RECT 2383.550 1530.305 2383.725 1531.565 ;
        RECT 2384.505 1530.305 2384.680 1531.565 ;
        RECT 2384.935 1531.445 2385.105 1533.045 ;
        RECT 2389.165 1532.935 2389.335 1533.105 ;
        RECT 2389.165 1532.605 2389.575 1532.935 ;
        RECT 2389.165 1532.095 2389.335 1532.605 ;
        RECT 2389.165 1531.765 2389.575 1532.095 ;
        RECT 2389.165 1531.565 2389.335 1531.765 ;
        RECT 2384.935 1530.305 2385.110 1531.445 ;
        RECT 2389.165 1530.305 2389.340 1531.565 ;
        RECT 2389.750 1531.535 2389.920 1533.145 ;
        RECT 2390.120 1533.085 2390.295 1533.595 ;
        RECT 2390.550 1533.045 2390.725 1533.595 ;
        RECT 2391.915 1533.085 2392.085 1533.595 ;
        RECT 2392.910 1533.080 2393.080 1533.590 ;
        RECT 2399.875 1533.105 2400.050 1533.595 ;
        RECT 2389.690 1531.365 2389.920 1531.535 ;
        RECT 2390.120 1531.565 2390.290 1532.515 ;
        RECT 2389.690 1530.305 2389.860 1531.365 ;
        RECT 2390.120 1530.305 2390.295 1531.565 ;
        RECT 2390.550 1531.445 2390.720 1533.045 ;
        RECT 2399.875 1532.935 2400.045 1533.105 ;
        RECT 2400.830 1533.085 2401.005 1533.595 ;
        RECT 2401.260 1533.045 2401.435 1533.595 ;
        RECT 2405.490 1533.105 2405.665 1533.595 ;
        RECT 2406.015 1533.315 2406.185 1533.595 ;
        RECT 2406.015 1533.145 2406.245 1533.315 ;
        RECT 2399.875 1532.605 2400.285 1532.935 ;
        RECT 2391.090 1532.425 2391.320 1532.575 ;
        RECT 2391.090 1532.255 2392.010 1532.425 ;
        RECT 2391.540 1531.565 2391.710 1532.255 ;
        RECT 2392.535 1532.250 2393.005 1532.420 ;
        RECT 2391.910 1531.775 2392.080 1531.885 ;
        RECT 2392.535 1531.775 2392.705 1532.250 ;
        RECT 2399.875 1532.095 2400.045 1532.605 ;
        RECT 2391.910 1531.605 2392.705 1531.775 ;
        RECT 2390.550 1530.305 2390.725 1531.445 ;
        RECT 2391.910 1530.305 2392.085 1531.605 ;
        RECT 2392.535 1531.560 2392.705 1531.605 ;
        RECT 2392.905 1531.445 2393.075 1531.880 ;
        RECT 2399.875 1531.765 2400.285 1532.095 ;
        RECT 2399.875 1531.565 2400.045 1531.765 ;
        RECT 2400.830 1531.565 2401.000 1532.515 ;
        RECT 2392.905 1530.300 2393.080 1531.445 ;
        RECT 2399.875 1530.305 2400.050 1531.565 ;
        RECT 2400.830 1530.305 2401.005 1531.565 ;
        RECT 2401.260 1531.445 2401.430 1533.045 ;
        RECT 2405.490 1532.935 2405.660 1533.105 ;
        RECT 2405.490 1532.605 2405.900 1532.935 ;
        RECT 2405.490 1532.095 2405.660 1532.605 ;
        RECT 2405.490 1531.765 2405.900 1532.095 ;
        RECT 2405.490 1531.565 2405.660 1531.765 ;
        RECT 2401.260 1530.305 2401.435 1531.445 ;
        RECT 2405.490 1530.305 2405.665 1531.565 ;
        RECT 2406.075 1531.535 2406.245 1533.145 ;
        RECT 2406.445 1533.085 2406.620 1533.595 ;
        RECT 2406.875 1533.045 2407.050 1533.595 ;
        RECT 2408.240 1533.085 2408.410 1533.595 ;
        RECT 2409.235 1533.080 2409.405 1533.590 ;
        RECT 2416.200 1533.105 2416.375 1533.595 ;
        RECT 2406.015 1531.365 2406.245 1531.535 ;
        RECT 2406.445 1531.565 2406.615 1532.515 ;
        RECT 2406.015 1530.305 2406.185 1531.365 ;
        RECT 2406.445 1530.305 2406.620 1531.565 ;
        RECT 2406.875 1531.445 2407.045 1533.045 ;
        RECT 2416.200 1532.935 2416.370 1533.105 ;
        RECT 2417.155 1533.085 2417.330 1533.595 ;
        RECT 2417.585 1533.045 2417.760 1533.595 ;
        RECT 2421.815 1533.105 2421.990 1533.595 ;
        RECT 2422.340 1533.315 2422.510 1533.595 ;
        RECT 2422.340 1533.145 2422.570 1533.315 ;
        RECT 2416.200 1532.605 2416.610 1532.935 ;
        RECT 2407.415 1532.425 2407.645 1532.575 ;
        RECT 2407.415 1532.255 2408.335 1532.425 ;
        RECT 2407.865 1531.565 2408.035 1532.255 ;
        RECT 2408.860 1532.250 2409.330 1532.420 ;
        RECT 2408.235 1531.775 2408.405 1531.885 ;
        RECT 2408.860 1531.775 2409.030 1532.250 ;
        RECT 2416.200 1532.095 2416.370 1532.605 ;
        RECT 2408.235 1531.605 2409.030 1531.775 ;
        RECT 2406.875 1530.305 2407.050 1531.445 ;
        RECT 2408.235 1530.305 2408.410 1531.605 ;
        RECT 2408.860 1531.560 2409.030 1531.605 ;
        RECT 2409.230 1531.445 2409.400 1531.880 ;
        RECT 2416.200 1531.765 2416.610 1532.095 ;
        RECT 2416.200 1531.565 2416.370 1531.765 ;
        RECT 2417.155 1531.565 2417.325 1532.515 ;
        RECT 2409.230 1530.300 2409.405 1531.445 ;
        RECT 2416.200 1530.305 2416.375 1531.565 ;
        RECT 2417.155 1530.305 2417.330 1531.565 ;
        RECT 2417.585 1531.445 2417.755 1533.045 ;
        RECT 2421.815 1532.935 2421.985 1533.105 ;
        RECT 2421.815 1532.605 2422.225 1532.935 ;
        RECT 2421.815 1532.095 2421.985 1532.605 ;
        RECT 2421.815 1531.765 2422.225 1532.095 ;
        RECT 2421.815 1531.565 2421.985 1531.765 ;
        RECT 2417.585 1530.305 2417.760 1531.445 ;
        RECT 2421.815 1530.305 2421.990 1531.565 ;
        RECT 2422.400 1531.535 2422.570 1533.145 ;
        RECT 2422.770 1533.085 2422.945 1533.595 ;
        RECT 2423.200 1533.045 2423.375 1533.595 ;
        RECT 2424.565 1533.085 2424.735 1533.595 ;
        RECT 2425.560 1533.080 2425.730 1533.590 ;
        RECT 2432.525 1533.105 2432.700 1533.595 ;
        RECT 2422.340 1531.365 2422.570 1531.535 ;
        RECT 2422.770 1531.565 2422.940 1532.515 ;
        RECT 2422.340 1530.305 2422.510 1531.365 ;
        RECT 2422.770 1530.305 2422.945 1531.565 ;
        RECT 2423.200 1531.445 2423.370 1533.045 ;
        RECT 2432.525 1532.935 2432.695 1533.105 ;
        RECT 2433.480 1533.085 2433.655 1533.595 ;
        RECT 2433.910 1533.045 2434.085 1533.595 ;
        RECT 2438.140 1533.105 2438.315 1533.595 ;
        RECT 2438.665 1533.315 2438.835 1533.595 ;
        RECT 2438.665 1533.145 2438.895 1533.315 ;
        RECT 2432.525 1532.605 2432.935 1532.935 ;
        RECT 2423.740 1532.425 2423.970 1532.575 ;
        RECT 2423.740 1532.255 2424.660 1532.425 ;
        RECT 2424.190 1531.565 2424.360 1532.255 ;
        RECT 2425.185 1532.250 2425.655 1532.420 ;
        RECT 2424.560 1531.775 2424.730 1531.885 ;
        RECT 2425.185 1531.775 2425.355 1532.250 ;
        RECT 2432.525 1532.095 2432.695 1532.605 ;
        RECT 2424.560 1531.605 2425.355 1531.775 ;
        RECT 2423.200 1530.305 2423.375 1531.445 ;
        RECT 2424.560 1530.305 2424.735 1531.605 ;
        RECT 2425.185 1531.560 2425.355 1531.605 ;
        RECT 2425.555 1531.445 2425.725 1531.880 ;
        RECT 2432.525 1531.765 2432.935 1532.095 ;
        RECT 2432.525 1531.565 2432.695 1531.765 ;
        RECT 2433.480 1531.565 2433.650 1532.515 ;
        RECT 2425.555 1530.300 2425.730 1531.445 ;
        RECT 2432.525 1530.305 2432.700 1531.565 ;
        RECT 2433.480 1530.305 2433.655 1531.565 ;
        RECT 2433.910 1531.445 2434.080 1533.045 ;
        RECT 2438.140 1532.935 2438.310 1533.105 ;
        RECT 2438.140 1532.605 2438.550 1532.935 ;
        RECT 2438.140 1532.095 2438.310 1532.605 ;
        RECT 2438.140 1531.765 2438.550 1532.095 ;
        RECT 2438.140 1531.565 2438.310 1531.765 ;
        RECT 2433.910 1530.305 2434.085 1531.445 ;
        RECT 2438.140 1530.305 2438.315 1531.565 ;
        RECT 2438.725 1531.535 2438.895 1533.145 ;
        RECT 2439.095 1533.085 2439.270 1533.595 ;
        RECT 2439.525 1533.045 2439.700 1533.595 ;
        RECT 2440.890 1533.085 2441.060 1533.595 ;
        RECT 2441.885 1533.080 2442.055 1533.590 ;
        RECT 2438.665 1531.365 2438.895 1531.535 ;
        RECT 2439.095 1531.565 2439.265 1532.515 ;
        RECT 2438.665 1530.305 2438.835 1531.365 ;
        RECT 2439.095 1530.305 2439.270 1531.565 ;
        RECT 2439.525 1531.445 2439.695 1533.045 ;
        RECT 2440.065 1532.425 2440.295 1532.575 ;
        RECT 2440.065 1532.255 2440.985 1532.425 ;
        RECT 2440.515 1531.565 2440.685 1532.255 ;
        RECT 2441.510 1532.250 2441.980 1532.420 ;
        RECT 2440.885 1531.775 2441.055 1531.885 ;
        RECT 2441.510 1531.775 2441.680 1532.250 ;
        RECT 2440.885 1531.605 2441.680 1531.775 ;
        RECT 2439.525 1530.305 2439.700 1531.445 ;
        RECT 2440.885 1530.305 2441.060 1531.605 ;
        RECT 2441.510 1531.560 2441.680 1531.605 ;
        RECT 2441.880 1531.445 2442.050 1531.880 ;
        RECT 2441.880 1530.300 2442.055 1531.445 ;
        RECT 2362.225 1527.795 2362.515 1527.965 ;
        RECT 2361.865 1527.235 2362.035 1527.655 ;
        RECT 2362.225 1526.925 2362.395 1527.795 ;
        RECT 2363.545 1527.515 2363.955 1527.685 ;
        RECT 2362.025 1526.755 2362.395 1526.925 ;
        RECT 2362.585 1527.235 2363.235 1527.405 ;
        RECT 2363.785 1527.325 2363.955 1527.515 ;
        RECT 2364.305 1527.235 2364.475 1527.655 ;
        RECT 2364.665 1527.515 2364.955 1527.685 ;
        RECT 2362.585 1526.675 2362.755 1527.235 ;
        RECT 2363.065 1526.675 2363.235 1527.005 ;
        RECT 2364.665 1526.925 2364.835 1527.515 ;
        RECT 2365.745 1527.325 2365.915 1527.685 ;
        RECT 2368.185 1527.665 2368.355 1527.995 ;
        RECT 2369.185 1527.665 2369.355 1527.995 ;
        RECT 2366.665 1527.495 2367.955 1527.575 ;
        RECT 2368.585 1527.495 2368.915 1527.575 ;
        RECT 2366.665 1527.405 2368.915 1527.495 ;
        RECT 2370.065 1527.405 2370.395 1527.575 ;
        RECT 2367.705 1527.325 2368.835 1527.405 ;
        RECT 2369.305 1527.235 2370.315 1527.405 ;
        RECT 2363.465 1526.755 2363.955 1526.925 ;
        RECT 2364.465 1526.755 2364.835 1526.925 ;
        RECT 2363.785 1526.675 2363.955 1526.755 ;
        RECT 2365.025 1526.675 2365.195 1527.005 ;
        RECT 2365.505 1526.675 2365.675 1527.125 ;
        RECT 2365.905 1526.755 2367.235 1526.925 ;
        RECT 2366.985 1526.675 2367.155 1526.755 ;
        RECT 2367.465 1526.675 2367.635 1527.005 ;
        RECT 2367.945 1526.675 2368.115 1527.125 ;
        RECT 2369.305 1527.005 2369.475 1527.235 ;
        RECT 2369.305 1526.755 2369.595 1527.005 ;
        RECT 2369.425 1526.675 2369.595 1526.755 ;
        RECT 2369.905 1526.675 2370.075 1527.005 ;
        RECT 2372.840 1526.895 2373.015 1528.155 ;
        RECT 2373.365 1527.095 2373.535 1528.155 ;
        RECT 2373.365 1526.925 2373.595 1527.095 ;
        RECT 2372.840 1526.695 2373.010 1526.895 ;
        RECT 2365.985 1526.525 2366.155 1526.565 ;
        RECT 2365.985 1526.355 2366.475 1526.525 ;
        RECT 2368.425 1526.395 2368.835 1526.565 ;
        RECT 2362.345 1525.935 2362.515 1526.285 ;
        RECT 2363.305 1525.935 2363.475 1526.285 ;
        RECT 2364.785 1525.935 2364.955 1526.285 ;
        RECT 2366.745 1525.935 2366.915 1526.285 ;
        RECT 2368.665 1525.935 2368.835 1526.395 ;
        RECT 2372.840 1526.365 2373.250 1526.695 ;
        RECT 2369.185 1525.935 2369.355 1526.285 ;
        RECT 2370.145 1526.185 2370.315 1526.285 ;
        RECT 2370.145 1526.015 2370.875 1526.185 ;
        RECT 2372.840 1525.855 2373.010 1526.365 ;
        RECT 2372.840 1525.525 2373.250 1525.855 ;
        RECT 2372.840 1525.355 2373.010 1525.525 ;
        RECT 2372.840 1524.865 2373.015 1525.355 ;
        RECT 2373.425 1525.315 2373.595 1526.925 ;
        RECT 2373.795 1526.895 2373.970 1528.155 ;
        RECT 2374.225 1527.015 2374.400 1528.155 ;
        RECT 2373.795 1525.945 2373.965 1526.895 ;
        RECT 2374.225 1525.415 2374.395 1527.015 ;
        RECT 2375.585 1527.010 2375.760 1528.155 ;
        RECT 2376.575 1528.100 2376.750 1528.160 ;
        RECT 2376.570 1527.755 2376.750 1528.100 ;
        RECT 2376.575 1527.015 2376.750 1527.755 ;
        RECT 2378.550 1527.795 2378.840 1527.965 ;
        RECT 2378.190 1527.235 2378.360 1527.655 ;
        RECT 2375.215 1526.205 2375.385 1526.895 ;
        RECT 2375.585 1526.795 2375.755 1527.010 ;
        RECT 2376.205 1526.795 2376.375 1526.900 ;
        RECT 2375.585 1526.625 2376.375 1526.795 ;
        RECT 2375.585 1526.575 2375.755 1526.625 ;
        RECT 2376.205 1526.210 2376.375 1526.625 ;
        RECT 2376.575 1526.580 2376.745 1527.015 ;
        RECT 2378.550 1526.925 2378.720 1527.795 ;
        RECT 2379.870 1527.515 2380.280 1527.685 ;
        RECT 2378.350 1526.755 2378.720 1526.925 ;
        RECT 2378.910 1527.235 2379.560 1527.405 ;
        RECT 2380.110 1527.325 2380.280 1527.515 ;
        RECT 2380.630 1527.235 2380.800 1527.655 ;
        RECT 2380.990 1527.515 2381.280 1527.685 ;
        RECT 2378.910 1526.675 2379.080 1527.235 ;
        RECT 2379.390 1526.675 2379.560 1527.005 ;
        RECT 2380.990 1526.925 2381.160 1527.515 ;
        RECT 2382.070 1527.325 2382.240 1527.685 ;
        RECT 2384.510 1527.665 2384.680 1527.995 ;
        RECT 2385.510 1527.665 2385.680 1527.995 ;
        RECT 2382.990 1527.495 2384.280 1527.575 ;
        RECT 2384.910 1527.495 2385.240 1527.575 ;
        RECT 2382.990 1527.405 2385.240 1527.495 ;
        RECT 2386.390 1527.405 2386.720 1527.575 ;
        RECT 2384.030 1527.325 2385.160 1527.405 ;
        RECT 2385.630 1527.235 2386.640 1527.405 ;
        RECT 2379.790 1526.755 2380.280 1526.925 ;
        RECT 2380.790 1526.755 2381.160 1526.925 ;
        RECT 2380.110 1526.675 2380.280 1526.755 ;
        RECT 2381.350 1526.675 2381.520 1527.005 ;
        RECT 2381.830 1526.675 2382.000 1527.125 ;
        RECT 2382.230 1526.755 2383.560 1526.925 ;
        RECT 2383.310 1526.675 2383.480 1526.755 ;
        RECT 2383.790 1526.675 2383.960 1527.005 ;
        RECT 2384.270 1526.675 2384.440 1527.125 ;
        RECT 2385.630 1527.005 2385.800 1527.235 ;
        RECT 2385.630 1526.755 2385.920 1527.005 ;
        RECT 2385.750 1526.675 2385.920 1526.755 ;
        RECT 2386.230 1526.675 2386.400 1527.005 ;
        RECT 2389.165 1526.895 2389.340 1528.155 ;
        RECT 2389.690 1527.095 2389.860 1528.155 ;
        RECT 2389.690 1526.925 2389.920 1527.095 ;
        RECT 2389.165 1526.695 2389.335 1526.895 ;
        RECT 2382.310 1526.525 2382.480 1526.565 ;
        RECT 2382.310 1526.355 2382.800 1526.525 ;
        RECT 2384.750 1526.395 2385.160 1526.565 ;
        RECT 2374.765 1526.035 2375.685 1526.205 ;
        RECT 2376.205 1526.040 2376.675 1526.210 ;
        RECT 2374.765 1525.885 2374.995 1526.035 ;
        RECT 2378.670 1525.935 2378.840 1526.285 ;
        RECT 2379.630 1525.935 2379.800 1526.285 ;
        RECT 2381.110 1525.935 2381.280 1526.285 ;
        RECT 2383.070 1525.935 2383.240 1526.285 ;
        RECT 2384.990 1525.935 2385.160 1526.395 ;
        RECT 2389.165 1526.365 2389.575 1526.695 ;
        RECT 2385.510 1525.935 2385.680 1526.285 ;
        RECT 2386.470 1526.185 2386.640 1526.285 ;
        RECT 2386.470 1526.015 2387.200 1526.185 ;
        RECT 2389.165 1525.855 2389.335 1526.365 ;
        RECT 2389.165 1525.525 2389.575 1525.855 ;
        RECT 2373.365 1525.145 2373.595 1525.315 ;
        RECT 2373.365 1524.865 2373.535 1525.145 ;
        RECT 2373.795 1524.865 2373.970 1525.375 ;
        RECT 2374.225 1524.865 2374.400 1525.415 ;
        RECT 2375.590 1524.865 2375.760 1525.375 ;
        RECT 2376.580 1524.870 2376.750 1525.380 ;
        RECT 2389.165 1525.355 2389.335 1525.525 ;
        RECT 2389.165 1524.865 2389.340 1525.355 ;
        RECT 2389.750 1525.315 2389.920 1526.925 ;
        RECT 2390.120 1526.895 2390.295 1528.155 ;
        RECT 2390.550 1527.015 2390.725 1528.155 ;
        RECT 2390.120 1525.945 2390.290 1526.895 ;
        RECT 2390.550 1525.415 2390.720 1527.015 ;
        RECT 2391.910 1527.010 2392.085 1528.155 ;
        RECT 2392.900 1528.100 2393.075 1528.160 ;
        RECT 2392.895 1527.755 2393.075 1528.100 ;
        RECT 2392.900 1527.015 2393.075 1527.755 ;
        RECT 2394.875 1527.795 2395.165 1527.965 ;
        RECT 2394.515 1527.235 2394.685 1527.655 ;
        RECT 2391.540 1526.205 2391.710 1526.895 ;
        RECT 2391.910 1526.795 2392.080 1527.010 ;
        RECT 2392.530 1526.795 2392.700 1526.900 ;
        RECT 2391.910 1526.625 2392.700 1526.795 ;
        RECT 2391.910 1526.575 2392.080 1526.625 ;
        RECT 2392.530 1526.210 2392.700 1526.625 ;
        RECT 2392.900 1526.580 2393.070 1527.015 ;
        RECT 2394.875 1526.925 2395.045 1527.795 ;
        RECT 2396.195 1527.515 2396.605 1527.685 ;
        RECT 2394.675 1526.755 2395.045 1526.925 ;
        RECT 2395.235 1527.235 2395.885 1527.405 ;
        RECT 2396.435 1527.325 2396.605 1527.515 ;
        RECT 2396.955 1527.235 2397.125 1527.655 ;
        RECT 2397.315 1527.515 2397.605 1527.685 ;
        RECT 2395.235 1526.675 2395.405 1527.235 ;
        RECT 2395.715 1526.675 2395.885 1527.005 ;
        RECT 2397.315 1526.925 2397.485 1527.515 ;
        RECT 2398.395 1527.325 2398.565 1527.685 ;
        RECT 2400.835 1527.665 2401.005 1527.995 ;
        RECT 2401.835 1527.665 2402.005 1527.995 ;
        RECT 2399.315 1527.495 2400.605 1527.575 ;
        RECT 2401.235 1527.495 2401.565 1527.575 ;
        RECT 2399.315 1527.405 2401.565 1527.495 ;
        RECT 2402.715 1527.405 2403.045 1527.575 ;
        RECT 2400.355 1527.325 2401.485 1527.405 ;
        RECT 2401.955 1527.235 2402.965 1527.405 ;
        RECT 2396.115 1526.755 2396.605 1526.925 ;
        RECT 2397.115 1526.755 2397.485 1526.925 ;
        RECT 2396.435 1526.675 2396.605 1526.755 ;
        RECT 2397.675 1526.675 2397.845 1527.005 ;
        RECT 2398.155 1526.675 2398.325 1527.125 ;
        RECT 2398.555 1526.755 2399.885 1526.925 ;
        RECT 2399.635 1526.675 2399.805 1526.755 ;
        RECT 2400.115 1526.675 2400.285 1527.005 ;
        RECT 2400.595 1526.675 2400.765 1527.125 ;
        RECT 2401.955 1527.005 2402.125 1527.235 ;
        RECT 2401.955 1526.755 2402.245 1527.005 ;
        RECT 2402.075 1526.675 2402.245 1526.755 ;
        RECT 2402.555 1526.675 2402.725 1527.005 ;
        RECT 2405.490 1526.895 2405.665 1528.155 ;
        RECT 2406.015 1527.095 2406.185 1528.155 ;
        RECT 2406.015 1526.925 2406.245 1527.095 ;
        RECT 2405.490 1526.695 2405.660 1526.895 ;
        RECT 2398.635 1526.525 2398.805 1526.565 ;
        RECT 2398.635 1526.355 2399.125 1526.525 ;
        RECT 2401.075 1526.395 2401.485 1526.565 ;
        RECT 2391.090 1526.035 2392.010 1526.205 ;
        RECT 2392.530 1526.040 2393.000 1526.210 ;
        RECT 2391.090 1525.885 2391.320 1526.035 ;
        RECT 2394.995 1525.935 2395.165 1526.285 ;
        RECT 2395.955 1525.935 2396.125 1526.285 ;
        RECT 2397.435 1525.935 2397.605 1526.285 ;
        RECT 2399.395 1525.935 2399.565 1526.285 ;
        RECT 2401.315 1525.935 2401.485 1526.395 ;
        RECT 2405.490 1526.365 2405.900 1526.695 ;
        RECT 2401.835 1525.935 2402.005 1526.285 ;
        RECT 2402.795 1526.185 2402.965 1526.285 ;
        RECT 2402.795 1526.015 2403.525 1526.185 ;
        RECT 2405.490 1525.855 2405.660 1526.365 ;
        RECT 2405.490 1525.525 2405.900 1525.855 ;
        RECT 2389.690 1525.145 2389.920 1525.315 ;
        RECT 2389.690 1524.865 2389.860 1525.145 ;
        RECT 2390.120 1524.865 2390.295 1525.375 ;
        RECT 2390.550 1524.865 2390.725 1525.415 ;
        RECT 2391.915 1524.865 2392.085 1525.375 ;
        RECT 2392.905 1524.870 2393.075 1525.380 ;
        RECT 2405.490 1525.355 2405.660 1525.525 ;
        RECT 2405.490 1524.865 2405.665 1525.355 ;
        RECT 2406.075 1525.315 2406.245 1526.925 ;
        RECT 2406.445 1526.895 2406.620 1528.155 ;
        RECT 2406.875 1527.015 2407.050 1528.155 ;
        RECT 2406.445 1525.945 2406.615 1526.895 ;
        RECT 2406.875 1525.415 2407.045 1527.015 ;
        RECT 2408.235 1527.010 2408.410 1528.155 ;
        RECT 2409.225 1528.100 2409.400 1528.160 ;
        RECT 2409.220 1527.755 2409.400 1528.100 ;
        RECT 2409.225 1527.015 2409.400 1527.755 ;
        RECT 2411.200 1527.795 2411.490 1527.965 ;
        RECT 2410.840 1527.235 2411.010 1527.655 ;
        RECT 2407.865 1526.205 2408.035 1526.895 ;
        RECT 2408.235 1526.795 2408.405 1527.010 ;
        RECT 2408.855 1526.795 2409.025 1526.900 ;
        RECT 2408.235 1526.625 2409.025 1526.795 ;
        RECT 2408.235 1526.575 2408.405 1526.625 ;
        RECT 2408.855 1526.210 2409.025 1526.625 ;
        RECT 2409.225 1526.580 2409.395 1527.015 ;
        RECT 2411.200 1526.925 2411.370 1527.795 ;
        RECT 2412.520 1527.515 2412.930 1527.685 ;
        RECT 2411.000 1526.755 2411.370 1526.925 ;
        RECT 2411.560 1527.235 2412.210 1527.405 ;
        RECT 2412.760 1527.325 2412.930 1527.515 ;
        RECT 2413.280 1527.235 2413.450 1527.655 ;
        RECT 2413.640 1527.515 2413.930 1527.685 ;
        RECT 2411.560 1526.675 2411.730 1527.235 ;
        RECT 2412.040 1526.675 2412.210 1527.005 ;
        RECT 2413.640 1526.925 2413.810 1527.515 ;
        RECT 2414.720 1527.325 2414.890 1527.685 ;
        RECT 2417.160 1527.665 2417.330 1527.995 ;
        RECT 2418.160 1527.665 2418.330 1527.995 ;
        RECT 2415.640 1527.495 2416.930 1527.575 ;
        RECT 2417.560 1527.495 2417.890 1527.575 ;
        RECT 2415.640 1527.405 2417.890 1527.495 ;
        RECT 2419.040 1527.405 2419.370 1527.575 ;
        RECT 2416.680 1527.325 2417.810 1527.405 ;
        RECT 2418.280 1527.235 2419.290 1527.405 ;
        RECT 2412.440 1526.755 2412.930 1526.925 ;
        RECT 2413.440 1526.755 2413.810 1526.925 ;
        RECT 2412.760 1526.675 2412.930 1526.755 ;
        RECT 2414.000 1526.675 2414.170 1527.005 ;
        RECT 2414.480 1526.675 2414.650 1527.125 ;
        RECT 2414.880 1526.755 2416.210 1526.925 ;
        RECT 2415.960 1526.675 2416.130 1526.755 ;
        RECT 2416.440 1526.675 2416.610 1527.005 ;
        RECT 2416.920 1526.675 2417.090 1527.125 ;
        RECT 2418.280 1527.005 2418.450 1527.235 ;
        RECT 2418.280 1526.755 2418.570 1527.005 ;
        RECT 2418.400 1526.675 2418.570 1526.755 ;
        RECT 2418.880 1526.675 2419.050 1527.005 ;
        RECT 2421.815 1526.895 2421.990 1528.155 ;
        RECT 2422.340 1527.095 2422.510 1528.155 ;
        RECT 2422.340 1526.925 2422.570 1527.095 ;
        RECT 2421.815 1526.695 2421.985 1526.895 ;
        RECT 2414.960 1526.525 2415.130 1526.565 ;
        RECT 2414.960 1526.355 2415.450 1526.525 ;
        RECT 2417.400 1526.395 2417.810 1526.565 ;
        RECT 2407.415 1526.035 2408.335 1526.205 ;
        RECT 2408.855 1526.040 2409.325 1526.210 ;
        RECT 2407.415 1525.885 2407.645 1526.035 ;
        RECT 2411.320 1525.935 2411.490 1526.285 ;
        RECT 2412.280 1525.935 2412.450 1526.285 ;
        RECT 2413.760 1525.935 2413.930 1526.285 ;
        RECT 2415.720 1525.935 2415.890 1526.285 ;
        RECT 2417.640 1525.935 2417.810 1526.395 ;
        RECT 2421.815 1526.365 2422.225 1526.695 ;
        RECT 2418.160 1525.935 2418.330 1526.285 ;
        RECT 2419.120 1526.185 2419.290 1526.285 ;
        RECT 2419.120 1526.015 2419.850 1526.185 ;
        RECT 2421.815 1525.855 2421.985 1526.365 ;
        RECT 2421.815 1525.525 2422.225 1525.855 ;
        RECT 2406.015 1525.145 2406.245 1525.315 ;
        RECT 2406.015 1524.865 2406.185 1525.145 ;
        RECT 2406.445 1524.865 2406.620 1525.375 ;
        RECT 2406.875 1524.865 2407.050 1525.415 ;
        RECT 2408.240 1524.865 2408.410 1525.375 ;
        RECT 2409.230 1524.870 2409.400 1525.380 ;
        RECT 2421.815 1525.355 2421.985 1525.525 ;
        RECT 2421.815 1524.865 2421.990 1525.355 ;
        RECT 2422.400 1525.315 2422.570 1526.925 ;
        RECT 2422.770 1526.895 2422.945 1528.155 ;
        RECT 2423.200 1527.015 2423.375 1528.155 ;
        RECT 2422.770 1525.945 2422.940 1526.895 ;
        RECT 2423.200 1525.415 2423.370 1527.015 ;
        RECT 2424.560 1527.010 2424.735 1528.155 ;
        RECT 2425.550 1528.100 2425.725 1528.160 ;
        RECT 2425.545 1527.755 2425.725 1528.100 ;
        RECT 2425.550 1527.015 2425.725 1527.755 ;
        RECT 2427.525 1527.795 2427.815 1527.965 ;
        RECT 2427.165 1527.235 2427.335 1527.655 ;
        RECT 2424.190 1526.205 2424.360 1526.895 ;
        RECT 2424.560 1526.795 2424.730 1527.010 ;
        RECT 2425.180 1526.795 2425.350 1526.900 ;
        RECT 2424.560 1526.625 2425.350 1526.795 ;
        RECT 2424.560 1526.575 2424.730 1526.625 ;
        RECT 2425.180 1526.210 2425.350 1526.625 ;
        RECT 2425.550 1526.580 2425.720 1527.015 ;
        RECT 2427.525 1526.925 2427.695 1527.795 ;
        RECT 2428.845 1527.515 2429.255 1527.685 ;
        RECT 2427.325 1526.755 2427.695 1526.925 ;
        RECT 2427.885 1527.235 2428.535 1527.405 ;
        RECT 2429.085 1527.325 2429.255 1527.515 ;
        RECT 2429.605 1527.235 2429.775 1527.655 ;
        RECT 2429.965 1527.515 2430.255 1527.685 ;
        RECT 2427.885 1526.675 2428.055 1527.235 ;
        RECT 2428.365 1526.675 2428.535 1527.005 ;
        RECT 2429.965 1526.925 2430.135 1527.515 ;
        RECT 2431.045 1527.325 2431.215 1527.685 ;
        RECT 2433.485 1527.665 2433.655 1527.995 ;
        RECT 2434.485 1527.665 2434.655 1527.995 ;
        RECT 2431.965 1527.495 2433.255 1527.575 ;
        RECT 2433.885 1527.495 2434.215 1527.575 ;
        RECT 2431.965 1527.405 2434.215 1527.495 ;
        RECT 2435.365 1527.405 2435.695 1527.575 ;
        RECT 2433.005 1527.325 2434.135 1527.405 ;
        RECT 2434.605 1527.235 2435.615 1527.405 ;
        RECT 2428.765 1526.755 2429.255 1526.925 ;
        RECT 2429.765 1526.755 2430.135 1526.925 ;
        RECT 2429.085 1526.675 2429.255 1526.755 ;
        RECT 2430.325 1526.675 2430.495 1527.005 ;
        RECT 2430.805 1526.675 2430.975 1527.125 ;
        RECT 2431.205 1526.755 2432.535 1526.925 ;
        RECT 2432.285 1526.675 2432.455 1526.755 ;
        RECT 2432.765 1526.675 2432.935 1527.005 ;
        RECT 2433.245 1526.675 2433.415 1527.125 ;
        RECT 2434.605 1527.005 2434.775 1527.235 ;
        RECT 2434.605 1526.755 2434.895 1527.005 ;
        RECT 2434.725 1526.675 2434.895 1526.755 ;
        RECT 2435.205 1526.675 2435.375 1527.005 ;
        RECT 2438.140 1526.895 2438.315 1528.155 ;
        RECT 2438.665 1527.095 2438.835 1528.155 ;
        RECT 2438.665 1526.925 2438.895 1527.095 ;
        RECT 2438.140 1526.695 2438.310 1526.895 ;
        RECT 2431.285 1526.525 2431.455 1526.565 ;
        RECT 2431.285 1526.355 2431.775 1526.525 ;
        RECT 2433.725 1526.395 2434.135 1526.565 ;
        RECT 2423.740 1526.035 2424.660 1526.205 ;
        RECT 2425.180 1526.040 2425.650 1526.210 ;
        RECT 2423.740 1525.885 2423.970 1526.035 ;
        RECT 2427.645 1525.935 2427.815 1526.285 ;
        RECT 2428.605 1525.935 2428.775 1526.285 ;
        RECT 2430.085 1525.935 2430.255 1526.285 ;
        RECT 2432.045 1525.935 2432.215 1526.285 ;
        RECT 2433.965 1525.935 2434.135 1526.395 ;
        RECT 2438.140 1526.365 2438.550 1526.695 ;
        RECT 2434.485 1525.935 2434.655 1526.285 ;
        RECT 2435.445 1526.185 2435.615 1526.285 ;
        RECT 2435.445 1526.015 2436.175 1526.185 ;
        RECT 2438.140 1525.855 2438.310 1526.365 ;
        RECT 2438.140 1525.525 2438.550 1525.855 ;
        RECT 2422.340 1525.145 2422.570 1525.315 ;
        RECT 2422.340 1524.865 2422.510 1525.145 ;
        RECT 2422.770 1524.865 2422.945 1525.375 ;
        RECT 2423.200 1524.865 2423.375 1525.415 ;
        RECT 2424.565 1524.865 2424.735 1525.375 ;
        RECT 2425.555 1524.870 2425.725 1525.380 ;
        RECT 2438.140 1525.355 2438.310 1525.525 ;
        RECT 2438.140 1524.865 2438.315 1525.355 ;
        RECT 2438.725 1525.315 2438.895 1526.925 ;
        RECT 2439.095 1526.895 2439.270 1528.155 ;
        RECT 2439.525 1527.015 2439.700 1528.155 ;
        RECT 2439.095 1525.945 2439.265 1526.895 ;
        RECT 2439.525 1525.415 2439.695 1527.015 ;
        RECT 2440.885 1527.010 2441.060 1528.155 ;
        RECT 2441.875 1528.100 2442.050 1528.160 ;
        RECT 2441.870 1527.755 2442.050 1528.100 ;
        RECT 2441.875 1527.015 2442.050 1527.755 ;
        RECT 2440.515 1526.205 2440.685 1526.895 ;
        RECT 2440.885 1526.795 2441.055 1527.010 ;
        RECT 2441.505 1526.795 2441.675 1526.900 ;
        RECT 2440.885 1526.625 2441.675 1526.795 ;
        RECT 2440.885 1526.575 2441.055 1526.625 ;
        RECT 2441.505 1526.210 2441.675 1526.625 ;
        RECT 2441.875 1526.580 2442.045 1527.015 ;
        RECT 2440.065 1526.035 2440.985 1526.205 ;
        RECT 2441.505 1526.040 2441.975 1526.210 ;
        RECT 2440.065 1525.885 2440.295 1526.035 ;
        RECT 2438.665 1525.145 2438.895 1525.315 ;
        RECT 2438.665 1524.865 2438.835 1525.145 ;
        RECT 2439.095 1524.865 2439.270 1525.375 ;
        RECT 2439.525 1524.865 2439.700 1525.415 ;
        RECT 2440.890 1524.865 2441.060 1525.375 ;
        RECT 2441.880 1524.870 2442.050 1525.380 ;
        RECT 2696.985 1496.335 2697.245 1496.665 ;
        RECT 2696.985 1495.425 2697.155 1496.335 ;
        RECT 2697.940 1496.265 2698.145 1496.665 ;
        RECT 2697.940 1496.095 2698.625 1496.265 ;
        RECT 2697.865 1495.425 2698.115 1495.925 ;
        RECT 2696.985 1495.255 2698.115 1495.425 ;
        RECT 2696.985 1494.485 2697.255 1495.255 ;
        RECT 2698.285 1495.065 2698.625 1496.095 ;
        RECT 2697.960 1494.890 2698.625 1495.065 ;
        RECT 2698.825 1496.160 2699.085 1496.665 ;
        RECT 2699.775 1496.285 2699.945 1496.665 ;
        RECT 2698.825 1495.360 2698.995 1496.160 ;
        RECT 2699.280 1496.115 2699.945 1496.285 ;
        RECT 2700.205 1496.160 2700.465 1496.665 ;
        RECT 2701.155 1496.285 2701.325 1496.665 ;
        RECT 2699.280 1495.860 2699.450 1496.115 ;
        RECT 2699.165 1495.530 2699.450 1495.860 ;
        RECT 2699.685 1495.565 2700.015 1495.935 ;
        RECT 2699.280 1495.385 2699.450 1495.530 ;
        RECT 2697.960 1494.485 2698.145 1494.890 ;
        RECT 2698.825 1494.455 2699.095 1495.360 ;
        RECT 2699.280 1495.215 2699.945 1495.385 ;
        RECT 2699.775 1494.455 2699.945 1495.215 ;
        RECT 2700.205 1495.360 2700.375 1496.160 ;
        RECT 2700.660 1496.115 2701.325 1496.285 ;
        RECT 2709.035 1496.285 2709.205 1496.665 ;
        RECT 2709.035 1496.115 2709.750 1496.285 ;
        RECT 2700.660 1495.860 2700.830 1496.115 ;
        RECT 2700.545 1495.530 2700.830 1495.860 ;
        RECT 2701.065 1495.565 2701.395 1495.935 ;
        RECT 2709.580 1495.925 2709.750 1496.115 ;
        RECT 2709.920 1496.090 2710.175 1496.665 ;
        RECT 2722.335 1496.265 2722.540 1496.665 ;
        RECT 2723.235 1496.335 2723.495 1496.665 ;
        RECT 2709.580 1495.595 2709.835 1495.925 ;
        RECT 2700.660 1495.385 2700.830 1495.530 ;
        RECT 2709.580 1495.385 2709.750 1495.595 ;
        RECT 2700.205 1494.455 2700.475 1495.360 ;
        RECT 2700.660 1495.215 2701.325 1495.385 ;
        RECT 2701.155 1494.455 2701.325 1495.215 ;
        RECT 2709.035 1495.215 2709.750 1495.385 ;
        RECT 2710.005 1495.360 2710.175 1496.090 ;
        RECT 2709.035 1494.455 2709.205 1495.215 ;
        RECT 2709.920 1494.455 2710.175 1495.360 ;
        RECT 2721.855 1496.095 2722.540 1496.265 ;
        RECT 2721.855 1495.065 2722.195 1496.095 ;
        RECT 2722.365 1495.425 2722.615 1495.925 ;
        RECT 2723.325 1495.425 2723.495 1496.335 ;
        RECT 2722.365 1495.255 2723.495 1495.425 ;
        RECT 2721.855 1494.890 2722.520 1495.065 ;
        RECT 2722.335 1494.485 2722.520 1494.890 ;
        RECT 2723.225 1494.485 2723.495 1495.255 ;
        RECT 2731.485 1496.160 2731.745 1496.665 ;
        RECT 2732.435 1496.285 2732.605 1496.665 ;
        RECT 2731.485 1495.360 2731.665 1496.160 ;
        RECT 2731.940 1496.115 2732.605 1496.285 ;
        RECT 2731.940 1495.860 2732.110 1496.115 ;
        RECT 2731.835 1495.530 2732.110 1495.860 ;
        RECT 2731.940 1495.385 2732.110 1495.530 ;
        RECT 2731.485 1494.455 2731.755 1495.360 ;
        RECT 2731.940 1495.215 2732.615 1495.385 ;
        RECT 2732.435 1494.455 2732.615 1495.215 ;
        RECT 2697.075 1493.185 2697.245 1493.945 ;
        RECT 2697.075 1493.015 2697.740 1493.185 ;
        RECT 2697.925 1493.040 2698.195 1493.945 ;
        RECT 2697.570 1492.870 2697.740 1493.015 ;
        RECT 2697.005 1492.465 2697.335 1492.835 ;
        RECT 2697.570 1492.540 2697.855 1492.870 ;
        RECT 2697.570 1492.285 2697.740 1492.540 ;
        RECT 2697.075 1492.115 2697.740 1492.285 ;
        RECT 2698.025 1492.240 2698.195 1493.040 ;
        RECT 2697.075 1491.735 2697.245 1492.115 ;
        RECT 2697.935 1491.735 2698.195 1492.240 ;
        RECT 2697.075 1485.405 2697.245 1485.785 ;
        RECT 2697.075 1485.235 2697.740 1485.405 ;
        RECT 2697.935 1485.280 2698.195 1485.785 ;
        RECT 2697.005 1484.685 2697.335 1485.055 ;
        RECT 2697.570 1484.980 2697.740 1485.235 ;
        RECT 2697.570 1484.650 2697.855 1484.980 ;
        RECT 2697.570 1484.505 2697.740 1484.650 ;
        RECT 2697.075 1484.335 2697.740 1484.505 ;
        RECT 2698.025 1484.480 2698.195 1485.280 ;
        RECT 2697.075 1483.575 2697.245 1484.335 ;
        RECT 2697.925 1483.575 2698.195 1484.480 ;
        RECT 2697.075 1479.965 2697.245 1480.340 ;
        RECT 2697.915 1480.175 2698.990 1480.345 ;
        RECT 2697.915 1479.965 2698.085 1480.175 ;
        RECT 2697.075 1479.795 2698.085 1479.965 ;
        RECT 2698.310 1479.835 2698.650 1480.005 ;
        RECT 2698.820 1479.840 2698.990 1480.175 ;
        RECT 2700.280 1480.175 2701.880 1480.345 ;
        RECT 2698.310 1479.665 2698.600 1479.835 ;
        RECT 2697.050 1479.495 2697.395 1479.605 ;
        RECT 2697.045 1479.325 2697.395 1479.495 ;
        RECT 2697.050 1478.985 2697.395 1479.325 ;
        RECT 2697.705 1478.985 2698.140 1479.605 ;
        RECT 2698.310 1479.145 2698.480 1479.665 ;
        RECT 2699.160 1479.495 2699.520 1480.170 ;
        RECT 2700.280 1479.805 2700.450 1480.175 ;
        RECT 2701.525 1480.135 2701.880 1480.175 ;
        RECT 2700.620 1479.755 2700.950 1480.005 ;
        RECT 2700.635 1479.680 2700.950 1479.755 ;
        RECT 2701.120 1479.885 2701.290 1480.005 ;
        RECT 2702.395 1479.885 2702.640 1480.305 ;
        RECT 2703.410 1479.945 2703.585 1480.275 ;
        RECT 2703.930 1480.185 2704.100 1480.345 ;
        RECT 2703.930 1480.015 2704.460 1480.185 ;
        RECT 2704.630 1480.175 2705.625 1480.345 ;
        RECT 2704.630 1480.015 2704.800 1480.175 ;
        RECT 2701.120 1479.715 2702.640 1479.885 ;
        RECT 2698.980 1479.315 2699.520 1479.495 ;
        RECT 2699.160 1479.205 2699.520 1479.315 ;
        RECT 2698.310 1478.975 2698.945 1479.145 ;
        RECT 2699.160 1478.975 2699.965 1479.205 ;
        RECT 2697.075 1478.635 2698.605 1478.805 ;
        RECT 2697.075 1478.135 2697.245 1478.635 ;
        RECT 2698.435 1478.475 2698.605 1478.635 ;
        RECT 2698.775 1478.645 2698.945 1478.975 ;
        RECT 2698.775 1478.475 2699.105 1478.645 ;
        RECT 2697.915 1478.305 2698.085 1478.465 ;
        RECT 2699.275 1478.305 2699.445 1478.805 ;
        RECT 2697.915 1478.135 2699.445 1478.305 ;
        RECT 2699.615 1478.135 2699.965 1478.975 ;
        RECT 2700.165 1478.605 2700.465 1479.605 ;
        RECT 2700.635 1479.155 2700.805 1479.680 ;
        RECT 2701.120 1479.675 2701.290 1479.715 ;
        RECT 2700.975 1479.495 2701.305 1479.505 ;
        RECT 2700.975 1479.335 2701.360 1479.495 ;
        RECT 2701.190 1479.325 2701.360 1479.335 ;
        RECT 2701.700 1479.155 2701.945 1479.545 ;
        RECT 2700.635 1478.985 2701.395 1479.155 ;
        RECT 2701.645 1478.985 2701.945 1479.155 ;
        RECT 2700.725 1478.305 2700.895 1478.815 ;
        RECT 2701.065 1478.475 2701.395 1478.985 ;
        RECT 2701.700 1478.925 2701.945 1478.985 ;
        RECT 2702.150 1478.925 2702.480 1479.545 ;
        RECT 2702.955 1478.925 2703.245 1479.605 ;
        RECT 2703.415 1479.495 2703.585 1479.945 ;
        RECT 2703.880 1479.665 2704.120 1479.835 ;
        RECT 2703.415 1479.325 2703.705 1479.495 ;
        RECT 2701.565 1478.515 2702.630 1478.685 ;
        RECT 2701.565 1478.305 2701.735 1478.515 ;
        RECT 2700.725 1478.135 2701.735 1478.305 ;
        RECT 2702.460 1478.135 2702.630 1478.515 ;
        RECT 2703.415 1478.465 2703.585 1479.325 ;
        RECT 2703.400 1478.135 2703.585 1478.465 ;
        RECT 2703.880 1478.465 2704.050 1479.665 ;
        RECT 2704.290 1478.845 2704.460 1480.015 ;
        RECT 2705.110 1479.835 2705.285 1480.005 ;
        RECT 2704.870 1479.675 2705.285 1479.835 ;
        RECT 2705.455 1479.885 2705.625 1480.175 ;
        RECT 2705.455 1479.715 2706.025 1479.885 ;
        RECT 2704.870 1479.665 2705.280 1479.675 ;
        RECT 2705.090 1479.325 2705.545 1479.495 ;
        RECT 2705.855 1478.935 2706.025 1479.715 ;
        RECT 2704.290 1478.615 2705.075 1478.845 ;
        RECT 2704.745 1478.475 2705.075 1478.615 ;
        RECT 2705.375 1478.765 2706.025 1478.935 ;
        RECT 2703.880 1478.135 2704.090 1478.465 ;
        RECT 2704.260 1478.305 2704.590 1478.345 ;
        RECT 2705.375 1478.305 2705.545 1478.765 ;
        RECT 2704.260 1478.135 2705.545 1478.305 ;
        RECT 2706.215 1478.135 2706.475 1480.345 ;
        RECT 2697.075 1476.865 2697.245 1477.625 ;
        RECT 2697.075 1476.695 2697.740 1476.865 ;
        RECT 2697.925 1476.720 2698.195 1477.625 ;
        RECT 2697.570 1476.550 2697.740 1476.695 ;
        RECT 2697.005 1476.145 2697.335 1476.515 ;
        RECT 2697.570 1476.220 2697.855 1476.550 ;
        RECT 2697.570 1475.965 2697.740 1476.220 ;
        RECT 2697.075 1475.795 2697.740 1475.965 ;
        RECT 2698.025 1475.920 2698.195 1476.720 ;
        RECT 2697.075 1475.415 2697.245 1475.795 ;
        RECT 2697.935 1475.415 2698.195 1475.920 ;
        RECT 2697.075 1474.525 2697.245 1474.900 ;
        RECT 2697.915 1474.735 2698.990 1474.905 ;
        RECT 2697.915 1474.525 2698.085 1474.735 ;
        RECT 2697.075 1474.355 2698.085 1474.525 ;
        RECT 2698.310 1474.395 2698.650 1474.565 ;
        RECT 2698.820 1474.400 2698.990 1474.735 ;
        RECT 2700.280 1474.735 2701.880 1474.905 ;
        RECT 2698.310 1474.225 2698.600 1474.395 ;
        RECT 2697.050 1474.055 2697.395 1474.165 ;
        RECT 2697.045 1473.885 2697.395 1474.055 ;
        RECT 2697.050 1473.545 2697.395 1473.885 ;
        RECT 2697.705 1473.545 2698.140 1474.165 ;
        RECT 2698.310 1473.705 2698.480 1474.225 ;
        RECT 2699.160 1474.055 2699.520 1474.730 ;
        RECT 2700.280 1474.365 2700.450 1474.735 ;
        RECT 2701.525 1474.695 2701.880 1474.735 ;
        RECT 2700.620 1474.315 2700.950 1474.565 ;
        RECT 2700.635 1474.240 2700.950 1474.315 ;
        RECT 2701.120 1474.445 2701.290 1474.565 ;
        RECT 2702.395 1474.445 2702.640 1474.865 ;
        RECT 2703.410 1474.505 2703.585 1474.835 ;
        RECT 2703.930 1474.745 2704.100 1474.905 ;
        RECT 2703.930 1474.575 2704.460 1474.745 ;
        RECT 2704.630 1474.735 2705.625 1474.905 ;
        RECT 2704.630 1474.575 2704.800 1474.735 ;
        RECT 2701.120 1474.275 2702.640 1474.445 ;
        RECT 2698.980 1473.875 2699.520 1474.055 ;
        RECT 2699.160 1473.765 2699.520 1473.875 ;
        RECT 2698.310 1473.535 2698.945 1473.705 ;
        RECT 2699.160 1473.535 2699.965 1473.765 ;
        RECT 2697.075 1473.195 2698.605 1473.365 ;
        RECT 2697.075 1472.695 2697.245 1473.195 ;
        RECT 2698.435 1473.035 2698.605 1473.195 ;
        RECT 2698.775 1473.205 2698.945 1473.535 ;
        RECT 2698.775 1473.035 2699.105 1473.205 ;
        RECT 2697.915 1472.865 2698.085 1473.025 ;
        RECT 2699.275 1472.865 2699.445 1473.365 ;
        RECT 2697.915 1472.695 2699.445 1472.865 ;
        RECT 2699.615 1472.695 2699.965 1473.535 ;
        RECT 2700.165 1473.165 2700.465 1474.165 ;
        RECT 2700.635 1473.715 2700.805 1474.240 ;
        RECT 2701.120 1474.235 2701.290 1474.275 ;
        RECT 2700.975 1474.055 2701.305 1474.065 ;
        RECT 2700.975 1473.895 2701.360 1474.055 ;
        RECT 2701.190 1473.885 2701.360 1473.895 ;
        RECT 2701.700 1473.715 2701.945 1474.105 ;
        RECT 2700.635 1473.545 2701.395 1473.715 ;
        RECT 2701.645 1473.545 2701.945 1473.715 ;
        RECT 2700.725 1472.865 2700.895 1473.375 ;
        RECT 2701.065 1473.035 2701.395 1473.545 ;
        RECT 2701.700 1473.485 2701.945 1473.545 ;
        RECT 2702.150 1473.485 2702.480 1474.105 ;
        RECT 2702.955 1473.485 2703.245 1474.165 ;
        RECT 2703.415 1474.055 2703.585 1474.505 ;
        RECT 2703.880 1474.225 2704.120 1474.395 ;
        RECT 2703.415 1473.885 2703.705 1474.055 ;
        RECT 2701.565 1473.075 2702.630 1473.245 ;
        RECT 2701.565 1472.865 2701.735 1473.075 ;
        RECT 2700.725 1472.695 2701.735 1472.865 ;
        RECT 2702.460 1472.695 2702.630 1473.075 ;
        RECT 2703.415 1473.025 2703.585 1473.885 ;
        RECT 2703.400 1472.695 2703.585 1473.025 ;
        RECT 2703.880 1473.025 2704.050 1474.225 ;
        RECT 2704.290 1473.405 2704.460 1474.575 ;
        RECT 2705.110 1474.395 2705.285 1474.565 ;
        RECT 2704.870 1474.235 2705.285 1474.395 ;
        RECT 2705.455 1474.445 2705.625 1474.735 ;
        RECT 2705.455 1474.275 2706.025 1474.445 ;
        RECT 2704.870 1474.225 2705.280 1474.235 ;
        RECT 2705.090 1473.885 2705.545 1474.055 ;
        RECT 2705.855 1473.495 2706.025 1474.275 ;
        RECT 2704.290 1473.175 2705.075 1473.405 ;
        RECT 2704.745 1473.035 2705.075 1473.175 ;
        RECT 2705.375 1473.325 2706.025 1473.495 ;
        RECT 2703.880 1472.695 2704.090 1473.025 ;
        RECT 2704.260 1472.865 2704.590 1472.905 ;
        RECT 2705.375 1472.865 2705.545 1473.325 ;
        RECT 2704.260 1472.695 2705.545 1472.865 ;
        RECT 2706.215 1472.695 2706.475 1474.905 ;
        RECT 2697.075 1471.425 2697.245 1472.185 ;
        RECT 2697.075 1471.255 2697.740 1471.425 ;
        RECT 2697.925 1471.280 2698.195 1472.185 ;
        RECT 2697.570 1471.110 2697.740 1471.255 ;
        RECT 2697.005 1470.705 2697.335 1471.075 ;
        RECT 2697.570 1470.780 2697.855 1471.110 ;
        RECT 2697.570 1470.525 2697.740 1470.780 ;
        RECT 2697.075 1470.355 2697.740 1470.525 ;
        RECT 2698.025 1470.480 2698.195 1471.280 ;
        RECT 2697.075 1469.975 2697.245 1470.355 ;
        RECT 2697.935 1469.975 2698.195 1470.480 ;
        RECT 2701.590 1471.215 2701.925 1472.185 ;
        RECT 2702.435 1472.015 2704.465 1472.185 ;
        RECT 2701.590 1470.545 2701.760 1471.215 ;
        RECT 2702.435 1471.045 2702.605 1472.015 ;
        RECT 2701.930 1470.715 2702.185 1471.045 ;
        RECT 2702.410 1470.715 2702.605 1471.045 ;
        RECT 2702.775 1471.675 2703.900 1471.845 ;
        RECT 2702.015 1470.545 2702.185 1470.715 ;
        RECT 2702.775 1470.545 2702.945 1471.675 ;
        RECT 2701.590 1469.975 2701.845 1470.545 ;
        RECT 2702.015 1470.375 2702.945 1470.545 ;
        RECT 2703.115 1471.335 2704.125 1471.505 ;
        RECT 2703.115 1470.535 2703.285 1471.335 ;
        RECT 2703.490 1470.655 2703.765 1471.135 ;
        RECT 2703.485 1470.485 2703.765 1470.655 ;
        RECT 2702.770 1470.340 2702.945 1470.375 ;
        RECT 2702.770 1469.975 2703.300 1470.340 ;
        RECT 2703.490 1469.975 2703.765 1470.485 ;
        RECT 2703.935 1469.975 2704.125 1471.335 ;
        RECT 2704.295 1471.350 2704.465 1472.015 ;
        RECT 2705.040 1471.595 2705.555 1472.005 ;
        RECT 2704.295 1471.160 2705.045 1471.350 ;
        RECT 2705.215 1470.785 2705.555 1471.595 ;
        RECT 2704.325 1470.615 2705.555 1470.785 ;
        RECT 2705.035 1470.010 2705.280 1470.615 ;
        RECT 2697.075 1465.985 2697.245 1466.745 ;
        RECT 2697.075 1465.815 2697.740 1465.985 ;
        RECT 2697.925 1465.840 2698.195 1466.745 ;
        RECT 2697.570 1465.670 2697.740 1465.815 ;
        RECT 2697.005 1465.265 2697.335 1465.635 ;
        RECT 2697.570 1465.340 2697.855 1465.670 ;
        RECT 2697.570 1465.085 2697.740 1465.340 ;
        RECT 2697.075 1464.915 2697.740 1465.085 ;
        RECT 2698.025 1465.040 2698.195 1465.840 ;
        RECT 2697.075 1464.535 2697.245 1464.915 ;
        RECT 2697.935 1464.535 2698.195 1465.040 ;
        RECT 2701.595 1460.505 2701.925 1461.290 ;
        RECT 2701.595 1460.335 2702.275 1460.505 ;
        RECT 2701.585 1459.915 2701.935 1460.165 ;
        RECT 2702.105 1459.735 2702.275 1460.335 ;
        RECT 2702.445 1459.915 2702.795 1460.165 ;
        RECT 2702.015 1459.095 2702.345 1459.735 ;
        RECT 2697.075 1458.205 2697.245 1458.585 ;
        RECT 2697.075 1458.035 2697.740 1458.205 ;
        RECT 2697.935 1458.080 2698.195 1458.585 ;
        RECT 2697.005 1457.485 2697.335 1457.855 ;
        RECT 2697.570 1457.780 2697.740 1458.035 ;
        RECT 2697.570 1457.450 2697.855 1457.780 ;
        RECT 2697.570 1457.305 2697.740 1457.450 ;
        RECT 2697.075 1457.135 2697.740 1457.305 ;
        RECT 2698.025 1457.280 2698.195 1458.080 ;
        RECT 2702.565 1458.225 2702.885 1458.585 ;
        RECT 2703.880 1458.225 2704.225 1458.585 ;
        RECT 2702.565 1458.055 2704.225 1458.225 ;
        RECT 2697.075 1456.375 2697.245 1457.135 ;
        RECT 2697.925 1456.375 2698.195 1457.280 ;
        RECT 2702.105 1457.215 2702.380 1457.845 ;
        RECT 2702.090 1456.555 2702.395 1457.045 ;
        RECT 2702.565 1456.725 2702.865 1458.055 ;
        RECT 2703.245 1457.595 2703.575 1457.765 ;
        RECT 2703.250 1457.345 2703.575 1457.595 ;
        RECT 2703.755 1457.515 2704.365 1457.845 ;
        RECT 2704.535 1457.345 2705.035 1457.805 ;
        RECT 2703.250 1457.165 2705.035 1457.345 ;
        RECT 2703.035 1456.815 2705.070 1456.985 ;
        RECT 2703.035 1456.555 2703.365 1456.815 ;
        RECT 2702.090 1456.375 2703.365 1456.555 ;
        RECT 2703.960 1456.735 2705.070 1456.815 ;
        RECT 2703.960 1456.375 2704.130 1456.735 ;
        RECT 2704.810 1456.375 2705.070 1456.735 ;
        RECT 2725.935 1455.015 2726.265 1455.865 ;
        RECT 2726.775 1455.015 2727.105 1455.865 ;
        RECT 2725.935 1454.845 2727.435 1455.015 ;
        RECT 2725.555 1454.475 2727.080 1454.675 ;
        RECT 2727.260 1454.645 2727.435 1454.845 ;
        RECT 2727.260 1454.475 2729.885 1454.645 ;
        RECT 2727.260 1454.305 2727.435 1454.475 ;
        RECT 2726.015 1454.135 2727.435 1454.305 ;
        RECT 2726.015 1453.655 2726.185 1454.135 ;
        RECT 2726.855 1453.660 2727.025 1454.135 ;
        RECT 2697.075 1452.765 2697.245 1453.145 ;
        RECT 2697.075 1452.595 2697.740 1452.765 ;
        RECT 2697.935 1452.640 2698.195 1453.145 ;
        RECT 2697.005 1452.045 2697.335 1452.415 ;
        RECT 2697.570 1452.340 2697.740 1452.595 ;
        RECT 2697.570 1452.010 2697.855 1452.340 ;
        RECT 2697.570 1451.865 2697.740 1452.010 ;
        RECT 2697.075 1451.695 2697.740 1451.865 ;
        RECT 2698.025 1451.840 2698.195 1452.640 ;
        RECT 2697.075 1450.935 2697.245 1451.695 ;
        RECT 2697.925 1450.935 2698.195 1451.840 ;
        RECT 2697.310 1447.305 2697.480 1447.555 ;
        RECT 2696.985 1447.135 2697.480 1447.305 ;
        RECT 2698.215 1447.305 2698.385 1447.650 ;
        RECT 2699.055 1447.305 2699.575 1447.705 ;
        RECT 2698.215 1447.135 2699.575 1447.305 ;
        RECT 2696.985 1446.175 2697.155 1447.135 ;
        RECT 2697.325 1446.345 2697.675 1446.965 ;
        RECT 2697.845 1446.345 2698.185 1446.965 ;
        RECT 2698.355 1446.345 2698.595 1446.965 ;
        RECT 2698.775 1446.715 2699.235 1446.885 ;
        RECT 2698.775 1446.175 2698.945 1446.715 ;
        RECT 2699.405 1446.515 2699.575 1447.135 ;
        RECT 2696.985 1446.005 2698.945 1446.175 ;
        RECT 2699.115 1445.505 2699.575 1446.515 ;
        RECT 2697.075 1444.225 2697.245 1444.985 ;
        RECT 2697.075 1444.055 2697.740 1444.225 ;
        RECT 2697.925 1444.080 2698.195 1444.985 ;
        RECT 2697.570 1443.910 2697.740 1444.055 ;
        RECT 2697.005 1443.505 2697.335 1443.875 ;
        RECT 2697.570 1443.580 2697.855 1443.910 ;
        RECT 2697.570 1443.325 2697.740 1443.580 ;
        RECT 2697.075 1443.155 2697.740 1443.325 ;
        RECT 2698.025 1443.280 2698.195 1444.080 ;
        RECT 2697.075 1442.775 2697.245 1443.155 ;
        RECT 2697.935 1442.775 2698.195 1443.280 ;
        RECT 2697.260 1441.625 2697.505 1442.230 ;
        RECT 2696.985 1441.455 2698.215 1441.625 ;
        RECT 2696.985 1440.645 2697.325 1441.455 ;
        RECT 2697.495 1440.890 2698.245 1441.080 ;
        RECT 2696.985 1440.235 2697.500 1440.645 ;
        RECT 2698.075 1440.225 2698.245 1440.890 ;
        RECT 2698.415 1440.905 2698.605 1442.265 ;
        RECT 2698.775 1442.095 2699.050 1442.265 ;
        RECT 2698.775 1441.925 2699.055 1442.095 ;
        RECT 2698.775 1441.105 2699.050 1441.925 ;
        RECT 2699.240 1441.900 2699.770 1442.265 ;
        RECT 2699.595 1441.865 2699.770 1441.900 ;
        RECT 2699.255 1440.905 2699.425 1441.705 ;
        RECT 2698.415 1440.735 2699.425 1440.905 ;
        RECT 2699.595 1441.695 2700.525 1441.865 ;
        RECT 2700.695 1441.695 2700.950 1442.265 ;
        RECT 2699.595 1440.565 2699.765 1441.695 ;
        RECT 2700.355 1441.525 2700.525 1441.695 ;
        RECT 2698.640 1440.395 2699.765 1440.565 ;
        RECT 2699.935 1441.195 2700.130 1441.525 ;
        RECT 2700.355 1441.195 2700.610 1441.525 ;
        RECT 2699.935 1440.225 2700.105 1441.195 ;
        RECT 2700.780 1441.025 2700.950 1441.695 ;
        RECT 2701.630 1441.500 2701.815 1442.170 ;
        RECT 2702.300 1441.815 2702.630 1442.215 ;
        RECT 2703.345 1441.820 2703.675 1442.260 ;
        RECT 2703.345 1441.815 2704.575 1441.820 ;
        RECT 2702.300 1441.705 2704.575 1441.815 ;
        RECT 2702.420 1441.640 2704.575 1441.705 ;
        RECT 2701.180 1441.230 2701.815 1441.500 ;
        RECT 2701.995 1441.120 2702.280 1441.525 ;
        RECT 2702.450 1441.120 2702.780 1441.470 ;
        RECT 2698.075 1440.055 2700.105 1440.225 ;
        RECT 2700.615 1440.055 2700.950 1441.025 ;
        RECT 2701.215 1440.770 2702.325 1440.940 ;
        RECT 2701.215 1440.060 2701.410 1440.770 ;
        RECT 2702.095 1440.060 2702.325 1440.770 ;
        RECT 2702.505 1440.065 2702.780 1441.120 ;
        RECT 2702.950 1440.065 2703.285 1441.470 ;
        RECT 2703.485 1440.065 2703.935 1441.470 ;
        RECT 2704.190 1440.060 2704.575 1441.640 ;
        RECT 2522.640 1436.565 2523.160 1438.050 ;
        RECT 2523.330 1437.225 2523.850 1438.775 ;
        RECT 2696.985 1438.155 2697.325 1439.035 ;
        RECT 2697.495 1438.325 2697.665 1439.545 ;
        RECT 2698.690 1439.205 2699.165 1439.545 ;
        RECT 2697.905 1438.675 2698.155 1439.040 ;
        RECT 2698.875 1438.675 2699.590 1438.970 ;
        RECT 2699.760 1438.845 2700.035 1439.545 ;
        RECT 2697.905 1438.505 2699.695 1438.675 ;
        RECT 2697.495 1438.075 2698.290 1438.325 ;
        RECT 2697.495 1437.985 2697.745 1438.075 ;
        RECT 2697.415 1437.565 2697.745 1437.985 ;
        RECT 2698.460 1437.650 2698.715 1438.505 ;
        RECT 2697.925 1437.385 2698.715 1437.650 ;
        RECT 2698.885 1437.805 2699.295 1438.325 ;
        RECT 2699.465 1438.075 2699.695 1438.505 ;
        RECT 2699.865 1437.815 2700.035 1438.845 ;
        RECT 2698.885 1437.385 2699.085 1437.805 ;
        RECT 2699.775 1437.335 2700.035 1437.815 ;
        RECT 2697.075 1436.445 2697.245 1436.825 ;
        RECT 2697.075 1436.275 2697.740 1436.445 ;
        RECT 2697.935 1436.320 2698.195 1436.825 ;
        RECT 2697.005 1435.725 2697.335 1436.095 ;
        RECT 2697.570 1436.020 2697.740 1436.275 ;
        RECT 2697.570 1435.690 2697.855 1436.020 ;
        RECT 2358.645 1435.110 2358.820 1435.600 ;
        RECT 2359.170 1435.320 2359.340 1435.600 ;
        RECT 2359.170 1435.150 2359.400 1435.320 ;
        RECT 2358.645 1434.940 2358.815 1435.110 ;
        RECT 2358.645 1434.610 2359.055 1434.940 ;
        RECT 2358.645 1434.100 2358.815 1434.610 ;
        RECT 2358.645 1433.770 2359.055 1434.100 ;
        RECT 2358.645 1433.570 2358.815 1433.770 ;
        RECT 2358.645 1432.310 2358.820 1433.570 ;
        RECT 2359.230 1433.540 2359.400 1435.150 ;
        RECT 2359.600 1435.090 2359.775 1435.600 ;
        RECT 2369.460 1435.110 2369.635 1435.600 ;
        RECT 2369.460 1434.940 2369.630 1435.110 ;
        RECT 2370.415 1435.090 2370.590 1435.600 ;
        RECT 2370.845 1435.050 2371.020 1435.600 ;
        RECT 2375.075 1435.110 2375.250 1435.600 ;
        RECT 2375.600 1435.320 2375.770 1435.600 ;
        RECT 2375.600 1435.150 2375.830 1435.320 ;
        RECT 2369.460 1434.610 2369.870 1434.940 ;
        RECT 2359.170 1433.370 2359.400 1433.540 ;
        RECT 2359.600 1433.570 2359.770 1434.520 ;
        RECT 2369.460 1434.100 2369.630 1434.610 ;
        RECT 2369.460 1433.770 2369.870 1434.100 ;
        RECT 2369.460 1433.570 2369.630 1433.770 ;
        RECT 2370.415 1433.570 2370.585 1434.520 ;
        RECT 2359.170 1432.310 2359.340 1433.370 ;
        RECT 2359.600 1432.310 2359.775 1433.570 ;
        RECT 2369.460 1432.310 2369.635 1433.570 ;
        RECT 2370.415 1432.310 2370.590 1433.570 ;
        RECT 2370.845 1433.450 2371.015 1435.050 ;
        RECT 2375.075 1434.940 2375.245 1435.110 ;
        RECT 2375.075 1434.610 2375.485 1434.940 ;
        RECT 2375.075 1434.100 2375.245 1434.610 ;
        RECT 2375.075 1433.770 2375.485 1434.100 ;
        RECT 2375.075 1433.570 2375.245 1433.770 ;
        RECT 2370.845 1432.310 2371.020 1433.450 ;
        RECT 2375.075 1432.310 2375.250 1433.570 ;
        RECT 2375.660 1433.540 2375.830 1435.150 ;
        RECT 2376.030 1435.090 2376.205 1435.600 ;
        RECT 2376.460 1435.050 2376.635 1435.600 ;
        RECT 2377.825 1435.090 2377.995 1435.600 ;
        RECT 2378.820 1435.085 2378.990 1435.595 ;
        RECT 2388.020 1435.110 2388.195 1435.600 ;
        RECT 2375.600 1433.370 2375.830 1433.540 ;
        RECT 2376.030 1433.570 2376.200 1434.520 ;
        RECT 2375.600 1432.310 2375.770 1433.370 ;
        RECT 2376.030 1432.310 2376.205 1433.570 ;
        RECT 2376.460 1433.450 2376.630 1435.050 ;
        RECT 2388.020 1434.940 2388.190 1435.110 ;
        RECT 2388.975 1435.090 2389.150 1435.600 ;
        RECT 2389.405 1435.050 2389.580 1435.600 ;
        RECT 2393.635 1435.110 2393.810 1435.600 ;
        RECT 2394.160 1435.320 2394.330 1435.600 ;
        RECT 2394.160 1435.150 2394.390 1435.320 ;
        RECT 2388.020 1434.610 2388.430 1434.940 ;
        RECT 2377.390 1434.430 2377.620 1434.600 ;
        RECT 2377.390 1434.370 2377.920 1434.430 ;
        RECT 2377.450 1434.260 2377.920 1434.370 ;
        RECT 2377.450 1433.570 2377.620 1434.260 ;
        RECT 2378.445 1434.255 2378.915 1434.425 ;
        RECT 2377.820 1433.810 2377.990 1433.890 ;
        RECT 2378.445 1433.810 2378.615 1434.255 ;
        RECT 2388.020 1434.100 2388.190 1434.610 ;
        RECT 2377.820 1433.610 2378.615 1433.810 ;
        RECT 2376.460 1432.310 2376.635 1433.450 ;
        RECT 2377.820 1432.310 2377.995 1433.610 ;
        RECT 2378.445 1433.565 2378.615 1433.610 ;
        RECT 2378.815 1433.450 2378.985 1433.885 ;
        RECT 2388.020 1433.770 2388.430 1434.100 ;
        RECT 2388.020 1433.570 2388.190 1433.770 ;
        RECT 2388.975 1433.570 2389.145 1434.520 ;
        RECT 2378.815 1432.305 2378.990 1433.450 ;
        RECT 2388.020 1432.310 2388.195 1433.570 ;
        RECT 2388.975 1432.310 2389.150 1433.570 ;
        RECT 2389.405 1433.450 2389.575 1435.050 ;
        RECT 2393.635 1434.940 2393.805 1435.110 ;
        RECT 2393.635 1434.610 2394.045 1434.940 ;
        RECT 2393.635 1434.100 2393.805 1434.610 ;
        RECT 2393.635 1433.770 2394.045 1434.100 ;
        RECT 2393.635 1433.570 2393.805 1433.770 ;
        RECT 2389.405 1432.310 2389.580 1433.450 ;
        RECT 2393.635 1432.310 2393.810 1433.570 ;
        RECT 2394.220 1433.540 2394.390 1435.150 ;
        RECT 2394.590 1435.090 2394.765 1435.600 ;
        RECT 2395.020 1435.050 2395.195 1435.600 ;
        RECT 2396.385 1435.090 2396.555 1435.600 ;
        RECT 2397.380 1435.085 2397.550 1435.595 ;
        RECT 2406.580 1435.110 2406.755 1435.600 ;
        RECT 2394.160 1433.370 2394.390 1433.540 ;
        RECT 2394.590 1433.570 2394.760 1434.520 ;
        RECT 2394.160 1432.310 2394.330 1433.370 ;
        RECT 2394.590 1432.310 2394.765 1433.570 ;
        RECT 2395.020 1433.450 2395.190 1435.050 ;
        RECT 2406.580 1434.940 2406.750 1435.110 ;
        RECT 2407.535 1435.090 2407.710 1435.600 ;
        RECT 2407.965 1435.050 2408.140 1435.600 ;
        RECT 2412.195 1435.110 2412.370 1435.600 ;
        RECT 2412.720 1435.320 2412.890 1435.600 ;
        RECT 2412.720 1435.150 2412.950 1435.320 ;
        RECT 2406.580 1434.610 2406.990 1434.940 ;
        RECT 2395.950 1434.430 2396.180 1434.600 ;
        RECT 2395.950 1434.370 2396.480 1434.430 ;
        RECT 2396.010 1434.260 2396.480 1434.370 ;
        RECT 2396.010 1433.570 2396.180 1434.260 ;
        RECT 2397.005 1434.255 2397.475 1434.425 ;
        RECT 2396.380 1433.810 2396.550 1433.890 ;
        RECT 2397.005 1433.810 2397.175 1434.255 ;
        RECT 2406.580 1434.100 2406.750 1434.610 ;
        RECT 2396.380 1433.610 2397.175 1433.810 ;
        RECT 2395.020 1432.310 2395.195 1433.450 ;
        RECT 2396.380 1432.310 2396.555 1433.610 ;
        RECT 2397.005 1433.565 2397.175 1433.610 ;
        RECT 2397.375 1433.450 2397.545 1433.885 ;
        RECT 2406.580 1433.770 2406.990 1434.100 ;
        RECT 2406.580 1433.570 2406.750 1433.770 ;
        RECT 2407.535 1433.570 2407.705 1434.520 ;
        RECT 2397.375 1432.305 2397.550 1433.450 ;
        RECT 2406.580 1432.310 2406.755 1433.570 ;
        RECT 2407.535 1432.310 2407.710 1433.570 ;
        RECT 2407.965 1433.450 2408.135 1435.050 ;
        RECT 2412.195 1434.940 2412.365 1435.110 ;
        RECT 2412.195 1434.610 2412.605 1434.940 ;
        RECT 2412.195 1434.100 2412.365 1434.610 ;
        RECT 2412.195 1433.770 2412.605 1434.100 ;
        RECT 2412.195 1433.570 2412.365 1433.770 ;
        RECT 2407.965 1432.310 2408.140 1433.450 ;
        RECT 2412.195 1432.310 2412.370 1433.570 ;
        RECT 2412.780 1433.540 2412.950 1435.150 ;
        RECT 2413.150 1435.090 2413.325 1435.600 ;
        RECT 2413.580 1435.050 2413.755 1435.600 ;
        RECT 2414.945 1435.090 2415.115 1435.600 ;
        RECT 2415.940 1435.085 2416.110 1435.595 ;
        RECT 2425.140 1435.110 2425.315 1435.600 ;
        RECT 2412.720 1433.370 2412.950 1433.540 ;
        RECT 2413.150 1433.570 2413.320 1434.520 ;
        RECT 2412.720 1432.310 2412.890 1433.370 ;
        RECT 2413.150 1432.310 2413.325 1433.570 ;
        RECT 2413.580 1433.450 2413.750 1435.050 ;
        RECT 2425.140 1434.940 2425.310 1435.110 ;
        RECT 2426.095 1435.090 2426.270 1435.600 ;
        RECT 2426.525 1435.050 2426.700 1435.600 ;
        RECT 2430.755 1435.110 2430.930 1435.600 ;
        RECT 2431.280 1435.320 2431.450 1435.600 ;
        RECT 2431.280 1435.150 2431.510 1435.320 ;
        RECT 2425.140 1434.610 2425.550 1434.940 ;
        RECT 2414.510 1434.430 2414.740 1434.600 ;
        RECT 2414.510 1434.370 2415.040 1434.430 ;
        RECT 2414.570 1434.260 2415.040 1434.370 ;
        RECT 2414.570 1433.570 2414.740 1434.260 ;
        RECT 2415.565 1434.255 2416.035 1434.425 ;
        RECT 2414.940 1433.810 2415.110 1433.890 ;
        RECT 2415.565 1433.810 2415.735 1434.255 ;
        RECT 2425.140 1434.100 2425.310 1434.610 ;
        RECT 2414.940 1433.610 2415.735 1433.810 ;
        RECT 2413.580 1432.310 2413.755 1433.450 ;
        RECT 2414.940 1432.310 2415.115 1433.610 ;
        RECT 2415.565 1433.565 2415.735 1433.610 ;
        RECT 2415.935 1433.450 2416.105 1433.885 ;
        RECT 2425.140 1433.770 2425.550 1434.100 ;
        RECT 2425.140 1433.570 2425.310 1433.770 ;
        RECT 2426.095 1433.570 2426.265 1434.520 ;
        RECT 2415.935 1432.305 2416.110 1433.450 ;
        RECT 2425.140 1432.310 2425.315 1433.570 ;
        RECT 2426.095 1432.310 2426.270 1433.570 ;
        RECT 2426.525 1433.450 2426.695 1435.050 ;
        RECT 2430.755 1434.940 2430.925 1435.110 ;
        RECT 2430.755 1434.610 2431.165 1434.940 ;
        RECT 2430.755 1434.100 2430.925 1434.610 ;
        RECT 2430.755 1433.770 2431.165 1434.100 ;
        RECT 2430.755 1433.570 2430.925 1433.770 ;
        RECT 2426.525 1432.310 2426.700 1433.450 ;
        RECT 2430.755 1432.310 2430.930 1433.570 ;
        RECT 2431.340 1433.540 2431.510 1435.150 ;
        RECT 2431.710 1435.090 2431.885 1435.600 ;
        RECT 2432.140 1435.050 2432.315 1435.600 ;
        RECT 2433.505 1435.090 2433.675 1435.600 ;
        RECT 2434.500 1435.085 2434.670 1435.595 ;
        RECT 2443.700 1435.110 2443.875 1435.600 ;
        RECT 2431.280 1433.370 2431.510 1433.540 ;
        RECT 2431.710 1433.570 2431.880 1434.520 ;
        RECT 2431.280 1432.310 2431.450 1433.370 ;
        RECT 2431.710 1432.310 2431.885 1433.570 ;
        RECT 2432.140 1433.450 2432.310 1435.050 ;
        RECT 2443.700 1434.940 2443.870 1435.110 ;
        RECT 2444.655 1435.090 2444.830 1435.600 ;
        RECT 2445.085 1435.050 2445.260 1435.600 ;
        RECT 2449.315 1435.110 2449.490 1435.600 ;
        RECT 2449.840 1435.320 2450.010 1435.600 ;
        RECT 2449.840 1435.150 2450.070 1435.320 ;
        RECT 2443.700 1434.610 2444.110 1434.940 ;
        RECT 2433.070 1434.430 2433.300 1434.600 ;
        RECT 2433.070 1434.370 2433.600 1434.430 ;
        RECT 2433.130 1434.260 2433.600 1434.370 ;
        RECT 2433.130 1433.570 2433.300 1434.260 ;
        RECT 2434.125 1434.255 2434.595 1434.425 ;
        RECT 2433.500 1433.810 2433.670 1433.890 ;
        RECT 2434.125 1433.810 2434.295 1434.255 ;
        RECT 2443.700 1434.100 2443.870 1434.610 ;
        RECT 2433.500 1433.610 2434.295 1433.810 ;
        RECT 2432.140 1432.310 2432.315 1433.450 ;
        RECT 2433.500 1432.310 2433.675 1433.610 ;
        RECT 2434.125 1433.565 2434.295 1433.610 ;
        RECT 2434.495 1433.450 2434.665 1433.885 ;
        RECT 2443.700 1433.770 2444.110 1434.100 ;
        RECT 2443.700 1433.570 2443.870 1433.770 ;
        RECT 2444.655 1433.570 2444.825 1434.520 ;
        RECT 2434.495 1432.305 2434.670 1433.450 ;
        RECT 2443.700 1432.310 2443.875 1433.570 ;
        RECT 2444.655 1432.310 2444.830 1433.570 ;
        RECT 2445.085 1433.450 2445.255 1435.050 ;
        RECT 2449.315 1434.940 2449.485 1435.110 ;
        RECT 2449.315 1434.610 2449.725 1434.940 ;
        RECT 2449.315 1434.100 2449.485 1434.610 ;
        RECT 2449.315 1433.770 2449.725 1434.100 ;
        RECT 2449.315 1433.570 2449.485 1433.770 ;
        RECT 2445.085 1432.310 2445.260 1433.450 ;
        RECT 2449.315 1432.310 2449.490 1433.570 ;
        RECT 2449.900 1433.540 2450.070 1435.150 ;
        RECT 2450.270 1435.090 2450.445 1435.600 ;
        RECT 2450.700 1435.050 2450.875 1435.600 ;
        RECT 2452.065 1435.090 2452.235 1435.600 ;
        RECT 2453.060 1435.085 2453.230 1435.595 ;
        RECT 2697.570 1435.545 2697.740 1435.690 ;
        RECT 2697.075 1435.375 2697.740 1435.545 ;
        RECT 2698.025 1435.520 2698.195 1436.320 ;
        RECT 2449.840 1433.370 2450.070 1433.540 ;
        RECT 2450.270 1433.570 2450.440 1434.520 ;
        RECT 2449.840 1432.310 2450.010 1433.370 ;
        RECT 2450.270 1432.310 2450.445 1433.570 ;
        RECT 2450.700 1433.450 2450.870 1435.050 ;
        RECT 2697.075 1434.615 2697.245 1435.375 ;
        RECT 2697.925 1434.615 2698.195 1435.520 ;
        RECT 2451.630 1434.430 2451.860 1434.600 ;
        RECT 2451.630 1434.370 2452.160 1434.430 ;
        RECT 2451.690 1434.260 2452.160 1434.370 ;
        RECT 2451.690 1433.570 2451.860 1434.260 ;
        RECT 2452.685 1434.255 2453.155 1434.425 ;
        RECT 2452.060 1433.810 2452.230 1433.890 ;
        RECT 2452.685 1433.810 2452.855 1434.255 ;
        RECT 2452.060 1433.610 2452.855 1433.810 ;
        RECT 2450.700 1432.310 2450.875 1433.450 ;
        RECT 2452.060 1432.310 2452.235 1433.610 ;
        RECT 2452.685 1433.565 2452.855 1433.610 ;
        RECT 2453.055 1433.450 2453.225 1433.885 ;
        RECT 2698.455 1433.605 2698.625 1434.105 ;
        RECT 2699.415 1433.605 2699.585 1434.105 ;
        RECT 2700.255 1433.605 2700.425 1434.105 ;
        RECT 2453.055 1432.305 2453.230 1433.450 ;
        RECT 2698.455 1433.435 2700.425 1433.605 ;
        RECT 2700.595 1433.635 2700.925 1434.065 ;
        RECT 2701.535 1433.805 2701.875 1434.065 ;
        RECT 2700.595 1433.465 2701.445 1433.635 ;
        RECT 2698.390 1432.635 2698.645 1433.265 ;
        RECT 2698.875 1432.635 2699.255 1433.265 ;
        RECT 2700.125 1433.255 2700.425 1433.260 ;
        RECT 2700.125 1433.085 2700.435 1433.255 ;
        RECT 2700.125 1432.965 2700.425 1433.085 ;
        RECT 2361.870 1429.575 2362.040 1429.935 ;
        RECT 2362.830 1429.605 2363.000 1429.765 ;
        RECT 2364.790 1429.685 2364.960 1429.795 ;
        RECT 2362.210 1429.435 2363.000 1429.605 ;
        RECT 2363.750 1429.515 2365.040 1429.685 ;
        RECT 2362.210 1429.375 2362.380 1429.435 ;
        RECT 2362.110 1429.205 2362.380 1429.375 ;
        RECT 2362.830 1429.345 2363.000 1429.435 ;
        RECT 2365.270 1429.345 2365.440 1429.765 ;
        RECT 2365.750 1429.435 2365.920 1429.795 ;
        RECT 2366.670 1429.515 2367.160 1429.685 ;
        RECT 2362.110 1429.135 2362.280 1429.205 ;
        RECT 2361.870 1428.865 2362.280 1429.135 ;
        RECT 2362.110 1428.785 2362.280 1428.865 ;
        RECT 2362.590 1428.785 2362.760 1429.115 ;
        RECT 2363.740 1428.865 2364.320 1429.035 ;
        RECT 2363.740 1428.785 2363.910 1428.865 ;
        RECT 2364.550 1428.785 2364.720 1429.235 ;
        RECT 2366.270 1429.035 2366.440 1429.515 ;
        RECT 2366.990 1429.345 2368.000 1429.515 ;
        RECT 2368.190 1429.435 2368.360 1430.075 ;
        RECT 2368.710 1429.775 2368.880 1430.105 ;
        RECT 2369.670 1429.905 2370.320 1430.075 ;
        RECT 2370.030 1429.515 2370.320 1429.905 ;
        RECT 2371.030 1429.905 2371.320 1430.075 ;
        RECT 2367.830 1429.115 2368.000 1429.345 ;
        RECT 2368.710 1429.375 2368.880 1429.515 ;
        RECT 2370.150 1429.435 2370.320 1429.515 ;
        RECT 2368.710 1429.205 2369.600 1429.375 ;
        RECT 2370.670 1429.345 2370.840 1429.765 ;
        RECT 2371.030 1429.515 2371.200 1429.905 ;
        RECT 2371.870 1429.515 2372.840 1429.685 ;
        RECT 2371.030 1429.345 2371.320 1429.515 ;
        RECT 2371.870 1429.345 2372.040 1429.515 ;
        RECT 2365.430 1428.865 2365.920 1429.035 ;
        RECT 2366.270 1428.865 2366.760 1429.035 ;
        RECT 2365.750 1428.785 2365.920 1428.865 ;
        RECT 2366.990 1428.785 2367.160 1429.115 ;
        RECT 2367.470 1428.785 2367.640 1429.115 ;
        RECT 2367.830 1428.865 2368.120 1429.115 ;
        RECT 2367.950 1428.785 2368.120 1428.865 ;
        RECT 2368.710 1428.865 2369.200 1429.035 ;
        RECT 2368.710 1428.785 2368.880 1428.865 ;
        RECT 2369.430 1428.785 2369.600 1429.205 ;
        RECT 2370.150 1429.135 2370.320 1429.235 ;
        RECT 2369.910 1429.035 2370.320 1429.135 ;
        RECT 2371.030 1429.035 2371.200 1429.345 ;
        RECT 2369.830 1428.965 2370.320 1429.035 ;
        RECT 2369.830 1428.865 2370.160 1428.965 ;
        RECT 2370.830 1428.865 2371.200 1429.035 ;
        RECT 2371.390 1429.035 2371.560 1429.115 ;
        RECT 2371.390 1428.865 2372.120 1429.035 ;
        RECT 2371.390 1428.785 2371.560 1428.865 ;
        RECT 2372.350 1428.785 2372.520 1429.235 ;
        RECT 2375.075 1428.895 2375.250 1430.155 ;
        RECT 2375.600 1429.095 2375.770 1430.155 ;
        RECT 2375.600 1428.925 2375.830 1429.095 ;
        RECT 2375.075 1428.695 2375.245 1428.895 ;
        RECT 2361.870 1428.045 2362.040 1428.395 ;
        RECT 2362.830 1428.295 2363.000 1428.395 ;
        RECT 2365.270 1428.295 2365.440 1428.395 ;
        RECT 2366.750 1428.295 2366.920 1428.395 ;
        RECT 2362.830 1428.125 2363.560 1428.295 ;
        RECT 2364.710 1428.125 2365.440 1428.295 ;
        RECT 2366.190 1428.125 2366.920 1428.295 ;
        RECT 2367.710 1428.045 2367.880 1428.395 ;
        RECT 2368.710 1428.045 2368.880 1428.395 ;
        RECT 2369.670 1428.045 2369.840 1428.395 ;
        RECT 2371.150 1428.045 2371.320 1428.395 ;
        RECT 2372.110 1428.045 2372.280 1428.395 ;
        RECT 2375.075 1428.365 2375.485 1428.695 ;
        RECT 2375.075 1427.855 2375.245 1428.365 ;
        RECT 2375.075 1427.525 2375.485 1427.855 ;
        RECT 2375.075 1427.355 2375.245 1427.525 ;
        RECT 2375.075 1426.865 2375.250 1427.355 ;
        RECT 2375.660 1427.315 2375.830 1428.925 ;
        RECT 2376.030 1428.895 2376.205 1430.155 ;
        RECT 2376.460 1429.015 2376.635 1430.155 ;
        RECT 2376.030 1427.945 2376.200 1428.895 ;
        RECT 2376.460 1427.415 2376.630 1429.015 ;
        RECT 2377.820 1429.010 2377.995 1430.155 ;
        RECT 2378.810 1429.015 2378.985 1430.160 ;
        RECT 2380.430 1429.575 2380.600 1429.935 ;
        RECT 2381.390 1429.605 2381.560 1429.765 ;
        RECT 2383.350 1429.685 2383.520 1429.795 ;
        RECT 2380.770 1429.435 2381.560 1429.605 ;
        RECT 2382.310 1429.515 2383.600 1429.685 ;
        RECT 2380.770 1429.375 2380.940 1429.435 ;
        RECT 2380.670 1429.205 2380.940 1429.375 ;
        RECT 2381.390 1429.345 2381.560 1429.435 ;
        RECT 2383.830 1429.345 2384.000 1429.765 ;
        RECT 2384.310 1429.435 2384.480 1429.795 ;
        RECT 2385.230 1429.515 2385.720 1429.685 ;
        RECT 2380.670 1429.135 2380.840 1429.205 ;
        RECT 2377.450 1428.205 2377.620 1428.895 ;
        RECT 2377.820 1428.805 2377.990 1429.010 ;
        RECT 2378.440 1428.805 2378.610 1428.900 ;
        RECT 2377.820 1428.625 2378.610 1428.805 ;
        RECT 2377.820 1428.575 2377.990 1428.625 ;
        RECT 2378.440 1428.210 2378.610 1428.625 ;
        RECT 2378.810 1428.580 2378.980 1429.015 ;
        RECT 2380.430 1428.865 2380.840 1429.135 ;
        RECT 2380.670 1428.785 2380.840 1428.865 ;
        RECT 2381.150 1428.785 2381.320 1429.115 ;
        RECT 2382.300 1428.865 2382.880 1429.035 ;
        RECT 2382.300 1428.785 2382.470 1428.865 ;
        RECT 2383.110 1428.785 2383.280 1429.235 ;
        RECT 2384.830 1429.035 2385.000 1429.515 ;
        RECT 2385.550 1429.345 2386.560 1429.515 ;
        RECT 2386.750 1429.435 2386.920 1430.075 ;
        RECT 2387.270 1429.775 2387.440 1430.105 ;
        RECT 2388.230 1429.905 2388.880 1430.075 ;
        RECT 2388.590 1429.515 2388.880 1429.905 ;
        RECT 2389.590 1429.905 2389.880 1430.075 ;
        RECT 2386.390 1429.115 2386.560 1429.345 ;
        RECT 2387.270 1429.375 2387.440 1429.515 ;
        RECT 2388.710 1429.435 2388.880 1429.515 ;
        RECT 2387.270 1429.205 2388.160 1429.375 ;
        RECT 2389.230 1429.345 2389.400 1429.765 ;
        RECT 2389.590 1429.515 2389.760 1429.905 ;
        RECT 2390.430 1429.515 2391.400 1429.685 ;
        RECT 2389.590 1429.345 2389.880 1429.515 ;
        RECT 2390.430 1429.345 2390.600 1429.515 ;
        RECT 2383.990 1428.865 2384.480 1429.035 ;
        RECT 2384.830 1428.865 2385.320 1429.035 ;
        RECT 2384.310 1428.785 2384.480 1428.865 ;
        RECT 2385.550 1428.785 2385.720 1429.115 ;
        RECT 2386.030 1428.785 2386.200 1429.115 ;
        RECT 2386.390 1428.865 2386.680 1429.115 ;
        RECT 2386.510 1428.785 2386.680 1428.865 ;
        RECT 2387.270 1428.865 2387.760 1429.035 ;
        RECT 2387.270 1428.785 2387.440 1428.865 ;
        RECT 2387.990 1428.785 2388.160 1429.205 ;
        RECT 2388.710 1429.135 2388.880 1429.235 ;
        RECT 2388.470 1429.035 2388.880 1429.135 ;
        RECT 2389.590 1429.035 2389.760 1429.345 ;
        RECT 2388.390 1428.965 2388.880 1429.035 ;
        RECT 2388.390 1428.865 2388.720 1428.965 ;
        RECT 2389.390 1428.865 2389.760 1429.035 ;
        RECT 2389.950 1429.035 2390.120 1429.115 ;
        RECT 2389.950 1428.865 2390.680 1429.035 ;
        RECT 2389.950 1428.785 2390.120 1428.865 ;
        RECT 2390.910 1428.785 2391.080 1429.235 ;
        RECT 2393.635 1428.895 2393.810 1430.155 ;
        RECT 2394.160 1429.095 2394.330 1430.155 ;
        RECT 2394.160 1428.925 2394.390 1429.095 ;
        RECT 2393.635 1428.695 2393.805 1428.895 ;
        RECT 2377.450 1428.175 2377.920 1428.205 ;
        RECT 2377.390 1428.035 2377.920 1428.175 ;
        RECT 2378.440 1428.040 2378.910 1428.210 ;
        RECT 2380.430 1428.045 2380.600 1428.395 ;
        RECT 2381.390 1428.295 2381.560 1428.395 ;
        RECT 2383.830 1428.295 2384.000 1428.395 ;
        RECT 2385.310 1428.295 2385.480 1428.395 ;
        RECT 2381.390 1428.125 2382.120 1428.295 ;
        RECT 2383.270 1428.125 2384.000 1428.295 ;
        RECT 2384.750 1428.125 2385.480 1428.295 ;
        RECT 2386.270 1428.045 2386.440 1428.395 ;
        RECT 2387.270 1428.045 2387.440 1428.395 ;
        RECT 2388.230 1428.045 2388.400 1428.395 ;
        RECT 2389.710 1428.045 2389.880 1428.395 ;
        RECT 2390.670 1428.045 2390.840 1428.395 ;
        RECT 2393.635 1428.365 2394.045 1428.695 ;
        RECT 2377.390 1427.945 2377.620 1428.035 ;
        RECT 2393.635 1427.855 2393.805 1428.365 ;
        RECT 2393.635 1427.525 2394.045 1427.855 ;
        RECT 2375.600 1427.145 2375.830 1427.315 ;
        RECT 2375.600 1426.865 2375.770 1427.145 ;
        RECT 2376.030 1426.865 2376.205 1427.375 ;
        RECT 2376.460 1426.865 2376.635 1427.415 ;
        RECT 2377.825 1426.865 2377.995 1427.375 ;
        RECT 2378.815 1426.870 2378.985 1427.380 ;
        RECT 2393.635 1427.355 2393.805 1427.525 ;
        RECT 2393.635 1426.865 2393.810 1427.355 ;
        RECT 2394.220 1427.315 2394.390 1428.925 ;
        RECT 2394.590 1428.895 2394.765 1430.155 ;
        RECT 2395.020 1429.015 2395.195 1430.155 ;
        RECT 2394.590 1427.945 2394.760 1428.895 ;
        RECT 2395.020 1427.415 2395.190 1429.015 ;
        RECT 2396.380 1429.010 2396.555 1430.155 ;
        RECT 2397.370 1429.015 2397.545 1430.160 ;
        RECT 2398.990 1429.575 2399.160 1429.935 ;
        RECT 2399.950 1429.605 2400.120 1429.765 ;
        RECT 2401.910 1429.685 2402.080 1429.795 ;
        RECT 2399.330 1429.435 2400.120 1429.605 ;
        RECT 2400.870 1429.515 2402.160 1429.685 ;
        RECT 2399.330 1429.375 2399.500 1429.435 ;
        RECT 2399.230 1429.205 2399.500 1429.375 ;
        RECT 2399.950 1429.345 2400.120 1429.435 ;
        RECT 2402.390 1429.345 2402.560 1429.765 ;
        RECT 2402.870 1429.435 2403.040 1429.795 ;
        RECT 2403.790 1429.515 2404.280 1429.685 ;
        RECT 2399.230 1429.135 2399.400 1429.205 ;
        RECT 2396.010 1428.205 2396.180 1428.895 ;
        RECT 2396.380 1428.805 2396.550 1429.010 ;
        RECT 2397.000 1428.805 2397.170 1428.900 ;
        RECT 2396.380 1428.625 2397.170 1428.805 ;
        RECT 2396.380 1428.575 2396.550 1428.625 ;
        RECT 2397.000 1428.210 2397.170 1428.625 ;
        RECT 2397.370 1428.580 2397.540 1429.015 ;
        RECT 2398.990 1428.865 2399.400 1429.135 ;
        RECT 2399.230 1428.785 2399.400 1428.865 ;
        RECT 2399.710 1428.785 2399.880 1429.115 ;
        RECT 2400.860 1428.865 2401.440 1429.035 ;
        RECT 2400.860 1428.785 2401.030 1428.865 ;
        RECT 2401.670 1428.785 2401.840 1429.235 ;
        RECT 2403.390 1429.035 2403.560 1429.515 ;
        RECT 2404.110 1429.345 2405.120 1429.515 ;
        RECT 2405.310 1429.435 2405.480 1430.075 ;
        RECT 2405.830 1429.775 2406.000 1430.105 ;
        RECT 2406.790 1429.905 2407.440 1430.075 ;
        RECT 2407.150 1429.515 2407.440 1429.905 ;
        RECT 2408.150 1429.905 2408.440 1430.075 ;
        RECT 2404.950 1429.115 2405.120 1429.345 ;
        RECT 2405.830 1429.375 2406.000 1429.515 ;
        RECT 2407.270 1429.435 2407.440 1429.515 ;
        RECT 2405.830 1429.205 2406.720 1429.375 ;
        RECT 2407.790 1429.345 2407.960 1429.765 ;
        RECT 2408.150 1429.515 2408.320 1429.905 ;
        RECT 2408.990 1429.515 2409.960 1429.685 ;
        RECT 2408.150 1429.345 2408.440 1429.515 ;
        RECT 2408.990 1429.345 2409.160 1429.515 ;
        RECT 2402.550 1428.865 2403.040 1429.035 ;
        RECT 2403.390 1428.865 2403.880 1429.035 ;
        RECT 2402.870 1428.785 2403.040 1428.865 ;
        RECT 2404.110 1428.785 2404.280 1429.115 ;
        RECT 2404.590 1428.785 2404.760 1429.115 ;
        RECT 2404.950 1428.865 2405.240 1429.115 ;
        RECT 2405.070 1428.785 2405.240 1428.865 ;
        RECT 2405.830 1428.865 2406.320 1429.035 ;
        RECT 2405.830 1428.785 2406.000 1428.865 ;
        RECT 2406.550 1428.785 2406.720 1429.205 ;
        RECT 2407.270 1429.135 2407.440 1429.235 ;
        RECT 2407.030 1429.035 2407.440 1429.135 ;
        RECT 2408.150 1429.035 2408.320 1429.345 ;
        RECT 2406.950 1428.965 2407.440 1429.035 ;
        RECT 2406.950 1428.865 2407.280 1428.965 ;
        RECT 2407.950 1428.865 2408.320 1429.035 ;
        RECT 2408.510 1429.035 2408.680 1429.115 ;
        RECT 2408.510 1428.865 2409.240 1429.035 ;
        RECT 2408.510 1428.785 2408.680 1428.865 ;
        RECT 2409.470 1428.785 2409.640 1429.235 ;
        RECT 2412.195 1428.895 2412.370 1430.155 ;
        RECT 2412.720 1429.095 2412.890 1430.155 ;
        RECT 2412.720 1428.925 2412.950 1429.095 ;
        RECT 2412.195 1428.695 2412.365 1428.895 ;
        RECT 2396.010 1428.175 2396.480 1428.205 ;
        RECT 2395.950 1428.035 2396.480 1428.175 ;
        RECT 2397.000 1428.040 2397.470 1428.210 ;
        RECT 2398.990 1428.045 2399.160 1428.395 ;
        RECT 2399.950 1428.295 2400.120 1428.395 ;
        RECT 2402.390 1428.295 2402.560 1428.395 ;
        RECT 2403.870 1428.295 2404.040 1428.395 ;
        RECT 2399.950 1428.125 2400.680 1428.295 ;
        RECT 2401.830 1428.125 2402.560 1428.295 ;
        RECT 2403.310 1428.125 2404.040 1428.295 ;
        RECT 2404.830 1428.045 2405.000 1428.395 ;
        RECT 2405.830 1428.045 2406.000 1428.395 ;
        RECT 2406.790 1428.045 2406.960 1428.395 ;
        RECT 2408.270 1428.045 2408.440 1428.395 ;
        RECT 2409.230 1428.045 2409.400 1428.395 ;
        RECT 2412.195 1428.365 2412.605 1428.695 ;
        RECT 2395.950 1427.945 2396.180 1428.035 ;
        RECT 2412.195 1427.855 2412.365 1428.365 ;
        RECT 2412.195 1427.525 2412.605 1427.855 ;
        RECT 2394.160 1427.145 2394.390 1427.315 ;
        RECT 2394.160 1426.865 2394.330 1427.145 ;
        RECT 2394.590 1426.865 2394.765 1427.375 ;
        RECT 2395.020 1426.865 2395.195 1427.415 ;
        RECT 2396.385 1426.865 2396.555 1427.375 ;
        RECT 2397.375 1426.870 2397.545 1427.380 ;
        RECT 2412.195 1427.355 2412.365 1427.525 ;
        RECT 2412.195 1426.865 2412.370 1427.355 ;
        RECT 2412.780 1427.315 2412.950 1428.925 ;
        RECT 2413.150 1428.895 2413.325 1430.155 ;
        RECT 2413.580 1429.015 2413.755 1430.155 ;
        RECT 2413.150 1427.945 2413.320 1428.895 ;
        RECT 2413.580 1427.415 2413.750 1429.015 ;
        RECT 2414.940 1429.010 2415.115 1430.155 ;
        RECT 2415.930 1429.015 2416.105 1430.160 ;
        RECT 2417.550 1429.575 2417.720 1429.935 ;
        RECT 2418.510 1429.605 2418.680 1429.765 ;
        RECT 2420.470 1429.685 2420.640 1429.795 ;
        RECT 2417.890 1429.435 2418.680 1429.605 ;
        RECT 2419.430 1429.515 2420.720 1429.685 ;
        RECT 2417.890 1429.375 2418.060 1429.435 ;
        RECT 2417.790 1429.205 2418.060 1429.375 ;
        RECT 2418.510 1429.345 2418.680 1429.435 ;
        RECT 2420.950 1429.345 2421.120 1429.765 ;
        RECT 2421.430 1429.435 2421.600 1429.795 ;
        RECT 2422.350 1429.515 2422.840 1429.685 ;
        RECT 2417.790 1429.135 2417.960 1429.205 ;
        RECT 2414.570 1428.205 2414.740 1428.895 ;
        RECT 2414.940 1428.805 2415.110 1429.010 ;
        RECT 2415.560 1428.805 2415.730 1428.900 ;
        RECT 2414.940 1428.625 2415.730 1428.805 ;
        RECT 2414.940 1428.575 2415.110 1428.625 ;
        RECT 2415.560 1428.210 2415.730 1428.625 ;
        RECT 2415.930 1428.580 2416.100 1429.015 ;
        RECT 2417.550 1428.865 2417.960 1429.135 ;
        RECT 2417.790 1428.785 2417.960 1428.865 ;
        RECT 2418.270 1428.785 2418.440 1429.115 ;
        RECT 2419.420 1428.865 2420.000 1429.035 ;
        RECT 2419.420 1428.785 2419.590 1428.865 ;
        RECT 2420.230 1428.785 2420.400 1429.235 ;
        RECT 2421.950 1429.035 2422.120 1429.515 ;
        RECT 2422.670 1429.345 2423.680 1429.515 ;
        RECT 2423.870 1429.435 2424.040 1430.075 ;
        RECT 2424.390 1429.775 2424.560 1430.105 ;
        RECT 2425.350 1429.905 2426.000 1430.075 ;
        RECT 2425.710 1429.515 2426.000 1429.905 ;
        RECT 2426.710 1429.905 2427.000 1430.075 ;
        RECT 2423.510 1429.115 2423.680 1429.345 ;
        RECT 2424.390 1429.375 2424.560 1429.515 ;
        RECT 2425.830 1429.435 2426.000 1429.515 ;
        RECT 2424.390 1429.205 2425.280 1429.375 ;
        RECT 2426.350 1429.345 2426.520 1429.765 ;
        RECT 2426.710 1429.515 2426.880 1429.905 ;
        RECT 2427.550 1429.515 2428.520 1429.685 ;
        RECT 2426.710 1429.345 2427.000 1429.515 ;
        RECT 2427.550 1429.345 2427.720 1429.515 ;
        RECT 2421.110 1428.865 2421.600 1429.035 ;
        RECT 2421.950 1428.865 2422.440 1429.035 ;
        RECT 2421.430 1428.785 2421.600 1428.865 ;
        RECT 2422.670 1428.785 2422.840 1429.115 ;
        RECT 2423.150 1428.785 2423.320 1429.115 ;
        RECT 2423.510 1428.865 2423.800 1429.115 ;
        RECT 2423.630 1428.785 2423.800 1428.865 ;
        RECT 2424.390 1428.865 2424.880 1429.035 ;
        RECT 2424.390 1428.785 2424.560 1428.865 ;
        RECT 2425.110 1428.785 2425.280 1429.205 ;
        RECT 2425.830 1429.135 2426.000 1429.235 ;
        RECT 2425.590 1429.035 2426.000 1429.135 ;
        RECT 2426.710 1429.035 2426.880 1429.345 ;
        RECT 2425.510 1428.965 2426.000 1429.035 ;
        RECT 2425.510 1428.865 2425.840 1428.965 ;
        RECT 2426.510 1428.865 2426.880 1429.035 ;
        RECT 2427.070 1429.035 2427.240 1429.115 ;
        RECT 2427.070 1428.865 2427.800 1429.035 ;
        RECT 2427.070 1428.785 2427.240 1428.865 ;
        RECT 2428.030 1428.785 2428.200 1429.235 ;
        RECT 2430.755 1428.895 2430.930 1430.155 ;
        RECT 2431.280 1429.095 2431.450 1430.155 ;
        RECT 2431.280 1428.925 2431.510 1429.095 ;
        RECT 2430.755 1428.695 2430.925 1428.895 ;
        RECT 2414.570 1428.175 2415.040 1428.205 ;
        RECT 2414.510 1428.035 2415.040 1428.175 ;
        RECT 2415.560 1428.040 2416.030 1428.210 ;
        RECT 2417.550 1428.045 2417.720 1428.395 ;
        RECT 2418.510 1428.295 2418.680 1428.395 ;
        RECT 2420.950 1428.295 2421.120 1428.395 ;
        RECT 2422.430 1428.295 2422.600 1428.395 ;
        RECT 2418.510 1428.125 2419.240 1428.295 ;
        RECT 2420.390 1428.125 2421.120 1428.295 ;
        RECT 2421.870 1428.125 2422.600 1428.295 ;
        RECT 2423.390 1428.045 2423.560 1428.395 ;
        RECT 2424.390 1428.045 2424.560 1428.395 ;
        RECT 2425.350 1428.045 2425.520 1428.395 ;
        RECT 2426.830 1428.045 2427.000 1428.395 ;
        RECT 2427.790 1428.045 2427.960 1428.395 ;
        RECT 2430.755 1428.365 2431.165 1428.695 ;
        RECT 2414.510 1427.945 2414.740 1428.035 ;
        RECT 2430.755 1427.855 2430.925 1428.365 ;
        RECT 2430.755 1427.525 2431.165 1427.855 ;
        RECT 2412.720 1427.145 2412.950 1427.315 ;
        RECT 2412.720 1426.865 2412.890 1427.145 ;
        RECT 2413.150 1426.865 2413.325 1427.375 ;
        RECT 2413.580 1426.865 2413.755 1427.415 ;
        RECT 2414.945 1426.865 2415.115 1427.375 ;
        RECT 2415.935 1426.870 2416.105 1427.380 ;
        RECT 2430.755 1427.355 2430.925 1427.525 ;
        RECT 2430.755 1426.865 2430.930 1427.355 ;
        RECT 2431.340 1427.315 2431.510 1428.925 ;
        RECT 2431.710 1428.895 2431.885 1430.155 ;
        RECT 2432.140 1429.015 2432.315 1430.155 ;
        RECT 2431.710 1427.945 2431.880 1428.895 ;
        RECT 2432.140 1427.415 2432.310 1429.015 ;
        RECT 2433.500 1429.010 2433.675 1430.155 ;
        RECT 2434.490 1429.015 2434.665 1430.160 ;
        RECT 2436.110 1429.575 2436.280 1429.935 ;
        RECT 2437.070 1429.605 2437.240 1429.765 ;
        RECT 2439.030 1429.685 2439.200 1429.795 ;
        RECT 2436.450 1429.435 2437.240 1429.605 ;
        RECT 2437.990 1429.515 2439.280 1429.685 ;
        RECT 2436.450 1429.375 2436.620 1429.435 ;
        RECT 2436.350 1429.205 2436.620 1429.375 ;
        RECT 2437.070 1429.345 2437.240 1429.435 ;
        RECT 2439.510 1429.345 2439.680 1429.765 ;
        RECT 2439.990 1429.435 2440.160 1429.795 ;
        RECT 2440.910 1429.515 2441.400 1429.685 ;
        RECT 2436.350 1429.135 2436.520 1429.205 ;
        RECT 2433.130 1428.205 2433.300 1428.895 ;
        RECT 2433.500 1428.805 2433.670 1429.010 ;
        RECT 2434.120 1428.805 2434.290 1428.900 ;
        RECT 2433.500 1428.625 2434.290 1428.805 ;
        RECT 2433.500 1428.575 2433.670 1428.625 ;
        RECT 2434.120 1428.210 2434.290 1428.625 ;
        RECT 2434.490 1428.580 2434.660 1429.015 ;
        RECT 2436.110 1428.865 2436.520 1429.135 ;
        RECT 2436.350 1428.785 2436.520 1428.865 ;
        RECT 2436.830 1428.785 2437.000 1429.115 ;
        RECT 2437.980 1428.865 2438.560 1429.035 ;
        RECT 2437.980 1428.785 2438.150 1428.865 ;
        RECT 2438.790 1428.785 2438.960 1429.235 ;
        RECT 2440.510 1429.035 2440.680 1429.515 ;
        RECT 2441.230 1429.345 2442.240 1429.515 ;
        RECT 2442.430 1429.435 2442.600 1430.075 ;
        RECT 2442.950 1429.775 2443.120 1430.105 ;
        RECT 2443.910 1429.905 2444.560 1430.075 ;
        RECT 2444.270 1429.515 2444.560 1429.905 ;
        RECT 2445.270 1429.905 2445.560 1430.075 ;
        RECT 2442.070 1429.115 2442.240 1429.345 ;
        RECT 2442.950 1429.375 2443.120 1429.515 ;
        RECT 2444.390 1429.435 2444.560 1429.515 ;
        RECT 2442.950 1429.205 2443.840 1429.375 ;
        RECT 2444.910 1429.345 2445.080 1429.765 ;
        RECT 2445.270 1429.515 2445.440 1429.905 ;
        RECT 2446.110 1429.515 2447.080 1429.685 ;
        RECT 2445.270 1429.345 2445.560 1429.515 ;
        RECT 2446.110 1429.345 2446.280 1429.515 ;
        RECT 2439.670 1428.865 2440.160 1429.035 ;
        RECT 2440.510 1428.865 2441.000 1429.035 ;
        RECT 2439.990 1428.785 2440.160 1428.865 ;
        RECT 2441.230 1428.785 2441.400 1429.115 ;
        RECT 2441.710 1428.785 2441.880 1429.115 ;
        RECT 2442.070 1428.865 2442.360 1429.115 ;
        RECT 2442.190 1428.785 2442.360 1428.865 ;
        RECT 2442.950 1428.865 2443.440 1429.035 ;
        RECT 2442.950 1428.785 2443.120 1428.865 ;
        RECT 2443.670 1428.785 2443.840 1429.205 ;
        RECT 2444.390 1429.135 2444.560 1429.235 ;
        RECT 2444.150 1429.035 2444.560 1429.135 ;
        RECT 2445.270 1429.035 2445.440 1429.345 ;
        RECT 2444.070 1428.965 2444.560 1429.035 ;
        RECT 2444.070 1428.865 2444.400 1428.965 ;
        RECT 2445.070 1428.865 2445.440 1429.035 ;
        RECT 2445.630 1429.035 2445.800 1429.115 ;
        RECT 2445.630 1428.865 2446.360 1429.035 ;
        RECT 2445.630 1428.785 2445.800 1428.865 ;
        RECT 2446.590 1428.785 2446.760 1429.235 ;
        RECT 2449.315 1428.895 2449.490 1430.155 ;
        RECT 2449.840 1429.095 2450.010 1430.155 ;
        RECT 2449.840 1428.925 2450.070 1429.095 ;
        RECT 2449.315 1428.695 2449.485 1428.895 ;
        RECT 2433.130 1428.175 2433.600 1428.205 ;
        RECT 2433.070 1428.035 2433.600 1428.175 ;
        RECT 2434.120 1428.040 2434.590 1428.210 ;
        RECT 2436.110 1428.045 2436.280 1428.395 ;
        RECT 2437.070 1428.295 2437.240 1428.395 ;
        RECT 2439.510 1428.295 2439.680 1428.395 ;
        RECT 2440.990 1428.295 2441.160 1428.395 ;
        RECT 2437.070 1428.125 2437.800 1428.295 ;
        RECT 2438.950 1428.125 2439.680 1428.295 ;
        RECT 2440.430 1428.125 2441.160 1428.295 ;
        RECT 2441.950 1428.045 2442.120 1428.395 ;
        RECT 2442.950 1428.045 2443.120 1428.395 ;
        RECT 2443.910 1428.045 2444.080 1428.395 ;
        RECT 2445.390 1428.045 2445.560 1428.395 ;
        RECT 2446.350 1428.045 2446.520 1428.395 ;
        RECT 2449.315 1428.365 2449.725 1428.695 ;
        RECT 2433.070 1427.945 2433.300 1428.035 ;
        RECT 2449.315 1427.855 2449.485 1428.365 ;
        RECT 2449.315 1427.525 2449.725 1427.855 ;
        RECT 2431.280 1427.145 2431.510 1427.315 ;
        RECT 2431.280 1426.865 2431.450 1427.145 ;
        RECT 2431.710 1426.865 2431.885 1427.375 ;
        RECT 2432.140 1426.865 2432.315 1427.415 ;
        RECT 2433.505 1426.865 2433.675 1427.375 ;
        RECT 2434.495 1426.870 2434.665 1427.380 ;
        RECT 2449.315 1427.355 2449.485 1427.525 ;
        RECT 2449.315 1426.865 2449.490 1427.355 ;
        RECT 2449.900 1427.315 2450.070 1428.925 ;
        RECT 2450.270 1428.895 2450.445 1430.155 ;
        RECT 2450.700 1429.015 2450.875 1430.155 ;
        RECT 2450.270 1427.945 2450.440 1428.895 ;
        RECT 2450.700 1427.415 2450.870 1429.015 ;
        RECT 2452.060 1429.010 2452.235 1430.155 ;
        RECT 2453.050 1429.015 2453.225 1430.160 ;
        RECT 2522.640 1430.150 2523.160 1431.635 ;
        RECT 2523.330 1430.810 2523.850 1432.360 ;
        RECT 2698.875 1432.035 2699.080 1432.635 ;
        RECT 2699.515 1432.240 2699.735 1432.965 ;
        RECT 2700.045 1432.635 2700.425 1432.965 ;
        RECT 2700.625 1432.715 2700.955 1433.275 ;
        RECT 2701.275 1432.545 2701.445 1433.465 ;
        RECT 2700.625 1432.450 2701.445 1432.545 ;
        RECT 2700.430 1432.375 2701.445 1432.450 ;
        RECT 2699.310 1432.055 2700.260 1432.240 ;
        RECT 2700.430 1431.940 2700.845 1432.375 ;
        RECT 2701.615 1432.200 2701.875 1433.805 ;
        RECT 2701.535 1431.940 2701.875 1432.200 ;
        RECT 2698.335 1430.735 2698.665 1431.155 ;
        RECT 2698.845 1430.985 2699.105 1431.385 ;
        RECT 2699.775 1430.985 2699.945 1431.335 ;
        RECT 2698.845 1430.815 2700.510 1430.985 ;
        RECT 2700.680 1430.880 2700.955 1431.225 ;
        RECT 2698.415 1430.645 2698.665 1430.735 ;
        RECT 2700.340 1430.645 2700.510 1430.815 ;
        RECT 2697.910 1430.315 2698.245 1430.565 ;
        RECT 2698.415 1430.315 2699.130 1430.645 ;
        RECT 2699.345 1430.315 2700.170 1430.645 ;
        RECT 2700.340 1430.315 2700.615 1430.645 ;
        RECT 2698.415 1429.755 2698.585 1430.315 ;
        RECT 2698.845 1429.855 2699.175 1430.145 ;
        RECT 2699.345 1430.025 2699.590 1430.315 ;
        RECT 2700.340 1430.145 2700.510 1430.315 ;
        RECT 2700.785 1430.145 2700.955 1430.880 ;
        RECT 2699.850 1429.975 2700.510 1430.145 ;
        RECT 2699.850 1429.855 2700.020 1429.975 ;
        RECT 2698.845 1429.685 2700.020 1429.855 ;
        RECT 2698.405 1429.185 2700.020 1429.515 ;
        RECT 2700.680 1429.175 2700.955 1430.145 ;
        RECT 2701.125 1431.155 2701.715 1431.385 ;
        RECT 2701.125 1430.145 2701.415 1431.155 ;
        RECT 2703.290 1430.985 2703.715 1431.195 ;
        RECT 2701.585 1430.815 2703.715 1430.985 ;
        RECT 2701.585 1430.315 2701.755 1430.815 ;
        RECT 2702.045 1430.315 2702.375 1430.645 ;
        RECT 2702.565 1430.315 2702.835 1430.645 ;
        RECT 2703.025 1430.315 2703.375 1430.645 ;
        RECT 2701.125 1429.975 2702.670 1430.145 ;
        RECT 2703.545 1430.045 2703.715 1430.815 ;
        RECT 2701.125 1429.175 2701.715 1429.975 ;
        RECT 2702.340 1429.175 2702.670 1429.975 ;
        RECT 2703.290 1429.715 2703.715 1430.045 ;
        RECT 2451.690 1428.205 2451.860 1428.895 ;
        RECT 2452.060 1428.805 2452.230 1429.010 ;
        RECT 2452.680 1428.805 2452.850 1428.900 ;
        RECT 2452.060 1428.625 2452.850 1428.805 ;
        RECT 2452.060 1428.575 2452.230 1428.625 ;
        RECT 2452.680 1428.210 2452.850 1428.625 ;
        RECT 2453.050 1428.580 2453.220 1429.015 ;
        RECT 2451.690 1428.175 2452.160 1428.205 ;
        RECT 2451.630 1428.035 2452.160 1428.175 ;
        RECT 2452.680 1428.040 2453.150 1428.210 ;
        RECT 2451.630 1427.945 2451.860 1428.035 ;
        RECT 2697.075 1427.905 2697.245 1428.665 ;
        RECT 2697.075 1427.735 2697.740 1427.905 ;
        RECT 2697.925 1427.760 2698.195 1428.665 ;
        RECT 2697.570 1427.590 2697.740 1427.735 ;
        RECT 2449.840 1427.145 2450.070 1427.315 ;
        RECT 2449.840 1426.865 2450.010 1427.145 ;
        RECT 2450.270 1426.865 2450.445 1427.375 ;
        RECT 2450.700 1426.865 2450.875 1427.415 ;
        RECT 2452.065 1426.865 2452.235 1427.375 ;
        RECT 2453.055 1426.870 2453.225 1427.380 ;
        RECT 2697.005 1427.185 2697.335 1427.555 ;
        RECT 2697.570 1427.260 2697.855 1427.590 ;
        RECT 2697.570 1427.005 2697.740 1427.260 ;
        RECT 2697.075 1426.835 2697.740 1427.005 ;
        RECT 2698.025 1426.960 2698.195 1427.760 ;
        RECT 2699.255 1427.685 2699.585 1428.665 ;
        RECT 2698.845 1427.275 2699.180 1427.525 ;
        RECT 2699.350 1427.085 2699.520 1427.685 ;
        RECT 2699.690 1427.255 2700.025 1427.525 ;
        RECT 2697.075 1426.455 2697.245 1426.835 ;
        RECT 2697.935 1426.455 2698.195 1426.960 ;
        RECT 2698.825 1426.455 2699.520 1427.085 ;
        RECT 2697.260 1425.305 2697.505 1425.910 ;
        RECT 2696.985 1425.135 2698.215 1425.305 ;
        RECT 2696.985 1424.325 2697.325 1425.135 ;
        RECT 2697.495 1424.570 2698.245 1424.760 ;
        RECT 2696.985 1423.915 2697.500 1424.325 ;
        RECT 2698.075 1423.905 2698.245 1424.570 ;
        RECT 2698.415 1424.585 2698.605 1425.945 ;
        RECT 2698.775 1425.095 2699.050 1425.945 ;
        RECT 2699.240 1425.580 2699.770 1425.945 ;
        RECT 2699.595 1425.545 2699.770 1425.580 ;
        RECT 2698.775 1424.925 2699.055 1425.095 ;
        RECT 2698.775 1424.785 2699.050 1424.925 ;
        RECT 2699.255 1424.585 2699.425 1425.385 ;
        RECT 2698.415 1424.415 2699.425 1424.585 ;
        RECT 2699.595 1425.375 2700.525 1425.545 ;
        RECT 2700.695 1425.375 2700.950 1425.945 ;
        RECT 2699.595 1424.245 2699.765 1425.375 ;
        RECT 2700.355 1425.205 2700.525 1425.375 ;
        RECT 2698.640 1424.075 2699.765 1424.245 ;
        RECT 2699.935 1424.875 2700.130 1425.205 ;
        RECT 2700.355 1424.875 2700.610 1425.205 ;
        RECT 2699.935 1423.905 2700.105 1424.875 ;
        RECT 2700.780 1424.705 2700.950 1425.375 ;
        RECT 2698.075 1423.735 2700.105 1423.905 ;
        RECT 2700.615 1423.735 2700.950 1424.705 ;
        RECT 2697.075 1422.465 2697.245 1423.225 ;
        RECT 2697.075 1422.295 2697.740 1422.465 ;
        RECT 2697.925 1422.320 2698.195 1423.225 ;
        RECT 2697.570 1422.150 2697.740 1422.295 ;
        RECT 2697.005 1421.745 2697.335 1422.115 ;
        RECT 2697.570 1421.820 2697.855 1422.150 ;
        RECT 2697.570 1421.565 2697.740 1421.820 ;
        RECT 2697.075 1421.395 2697.740 1421.565 ;
        RECT 2698.025 1421.520 2698.195 1422.320 ;
        RECT 2697.075 1421.015 2697.245 1421.395 ;
        RECT 2697.935 1421.015 2698.195 1421.520 ;
        RECT 2522.640 1415.960 2523.160 1417.445 ;
        RECT 2523.330 1416.620 2523.850 1418.170 ;
        RECT 2697.075 1417.025 2697.245 1417.785 ;
        RECT 2697.075 1416.855 2697.740 1417.025 ;
        RECT 2697.925 1416.880 2698.195 1417.785 ;
        RECT 2697.570 1416.710 2697.740 1416.855 ;
        RECT 2697.005 1416.305 2697.335 1416.675 ;
        RECT 2697.570 1416.380 2697.855 1416.710 ;
        RECT 2697.570 1416.125 2697.740 1416.380 ;
        RECT 2697.075 1415.955 2697.740 1416.125 ;
        RECT 2698.025 1416.080 2698.195 1416.880 ;
        RECT 2697.075 1415.575 2697.245 1415.955 ;
        RECT 2697.935 1415.575 2698.195 1416.080 ;
        RECT 2697.075 1411.585 2697.245 1412.345 ;
        RECT 2697.075 1411.415 2697.740 1411.585 ;
        RECT 2697.925 1411.440 2698.195 1412.345 ;
        RECT 2697.570 1411.270 2697.740 1411.415 ;
        RECT 2697.005 1410.865 2697.335 1411.235 ;
        RECT 2697.570 1410.940 2697.855 1411.270 ;
        RECT 2697.570 1410.685 2697.740 1410.940 ;
        RECT 2522.640 1408.430 2523.160 1409.915 ;
        RECT 2523.330 1409.090 2523.850 1410.640 ;
        RECT 2697.075 1410.515 2697.740 1410.685 ;
        RECT 2698.025 1410.640 2698.195 1411.440 ;
        RECT 2698.455 1411.585 2698.625 1412.345 ;
        RECT 2698.455 1411.415 2699.120 1411.585 ;
        RECT 2699.305 1411.440 2699.575 1412.345 ;
        RECT 2698.950 1411.270 2699.120 1411.415 ;
        RECT 2698.385 1410.865 2698.715 1411.235 ;
        RECT 2698.950 1410.940 2699.235 1411.270 ;
        RECT 2698.950 1410.685 2699.120 1410.940 ;
        RECT 2697.075 1410.135 2697.245 1410.515 ;
        RECT 2697.935 1410.135 2698.195 1410.640 ;
        RECT 2698.455 1410.515 2699.120 1410.685 ;
        RECT 2699.405 1410.640 2699.575 1411.440 ;
        RECT 2698.455 1410.135 2698.625 1410.515 ;
        RECT 2699.315 1410.135 2699.575 1410.640 ;
        RECT 2522.640 1402.450 2523.160 1403.935 ;
        RECT 2523.330 1403.110 2523.850 1404.660 ;
        RECT 2522.640 1394.035 2523.160 1395.520 ;
        RECT 2523.330 1394.695 2523.850 1396.245 ;
        RECT 2882.085 1361.420 2882.605 1362.970 ;
        RECT 2368.645 1335.110 2368.820 1335.600 ;
        RECT 2369.170 1335.320 2369.340 1335.600 ;
        RECT 2369.170 1335.150 2369.400 1335.320 ;
        RECT 2368.645 1334.940 2368.815 1335.110 ;
        RECT 2368.645 1334.610 2369.055 1334.940 ;
        RECT 2368.645 1334.100 2368.815 1334.610 ;
        RECT 2368.645 1333.770 2369.055 1334.100 ;
        RECT 2368.645 1333.570 2368.815 1333.770 ;
        RECT 2368.645 1332.310 2368.820 1333.570 ;
        RECT 2369.230 1333.540 2369.400 1335.150 ;
        RECT 2369.600 1335.090 2369.775 1335.600 ;
        RECT 2376.160 1335.110 2376.335 1335.600 ;
        RECT 2376.160 1334.940 2376.330 1335.110 ;
        RECT 2377.115 1335.090 2377.290 1335.600 ;
        RECT 2377.545 1335.050 2377.720 1335.600 ;
        RECT 2381.775 1335.110 2381.950 1335.600 ;
        RECT 2382.300 1335.320 2382.470 1335.600 ;
        RECT 2382.300 1335.150 2382.530 1335.320 ;
        RECT 2376.160 1334.610 2376.570 1334.940 ;
        RECT 2369.170 1333.370 2369.400 1333.540 ;
        RECT 2369.600 1333.570 2369.770 1334.520 ;
        RECT 2376.160 1334.100 2376.330 1334.610 ;
        RECT 2376.160 1333.770 2376.570 1334.100 ;
        RECT 2376.160 1333.570 2376.330 1333.770 ;
        RECT 2377.115 1333.570 2377.285 1334.520 ;
        RECT 2369.170 1332.310 2369.340 1333.370 ;
        RECT 2369.600 1332.310 2369.775 1333.570 ;
        RECT 2376.160 1332.310 2376.335 1333.570 ;
        RECT 2377.115 1332.310 2377.290 1333.570 ;
        RECT 2377.545 1333.450 2377.715 1335.050 ;
        RECT 2381.775 1334.940 2381.945 1335.110 ;
        RECT 2381.775 1334.610 2382.185 1334.940 ;
        RECT 2381.775 1334.100 2381.945 1334.610 ;
        RECT 2381.775 1333.770 2382.185 1334.100 ;
        RECT 2381.775 1333.570 2381.945 1333.770 ;
        RECT 2377.545 1332.310 2377.720 1333.450 ;
        RECT 2381.775 1332.310 2381.950 1333.570 ;
        RECT 2382.360 1333.540 2382.530 1335.150 ;
        RECT 2382.730 1335.090 2382.905 1335.600 ;
        RECT 2383.160 1335.050 2383.335 1335.600 ;
        RECT 2384.525 1335.090 2384.695 1335.600 ;
        RECT 2385.515 1335.090 2385.685 1335.600 ;
        RECT 2391.420 1335.110 2391.595 1335.600 ;
        RECT 2382.300 1333.370 2382.530 1333.540 ;
        RECT 2382.730 1333.570 2382.900 1334.520 ;
        RECT 2382.300 1332.310 2382.470 1333.370 ;
        RECT 2382.730 1332.310 2382.905 1333.570 ;
        RECT 2383.160 1333.450 2383.330 1335.050 ;
        RECT 2391.420 1334.940 2391.590 1335.110 ;
        RECT 2392.375 1335.090 2392.550 1335.600 ;
        RECT 2392.805 1335.050 2392.980 1335.600 ;
        RECT 2397.035 1335.110 2397.210 1335.600 ;
        RECT 2397.560 1335.320 2397.730 1335.600 ;
        RECT 2397.560 1335.150 2397.790 1335.320 ;
        RECT 2391.420 1334.610 2391.830 1334.940 ;
        RECT 2384.090 1334.430 2384.320 1334.585 ;
        RECT 2384.090 1334.355 2384.620 1334.430 ;
        RECT 2384.150 1334.260 2384.620 1334.355 ;
        RECT 2385.140 1334.260 2385.610 1334.430 ;
        RECT 2384.150 1333.570 2384.320 1334.260 ;
        RECT 2384.520 1333.810 2384.690 1333.890 ;
        RECT 2385.140 1333.810 2385.310 1334.260 ;
        RECT 2391.420 1334.100 2391.590 1334.610 ;
        RECT 2384.520 1333.610 2385.310 1333.810 ;
        RECT 2383.160 1332.310 2383.335 1333.450 ;
        RECT 2384.520 1332.310 2384.695 1333.610 ;
        RECT 2385.140 1333.570 2385.310 1333.610 ;
        RECT 2385.510 1333.455 2385.680 1333.890 ;
        RECT 2391.420 1333.770 2391.830 1334.100 ;
        RECT 2391.420 1333.570 2391.590 1333.770 ;
        RECT 2392.375 1333.570 2392.545 1334.520 ;
        RECT 2385.510 1332.310 2385.685 1333.455 ;
        RECT 2391.420 1332.310 2391.595 1333.570 ;
        RECT 2392.375 1332.310 2392.550 1333.570 ;
        RECT 2392.805 1333.450 2392.975 1335.050 ;
        RECT 2397.035 1334.940 2397.205 1335.110 ;
        RECT 2397.035 1334.610 2397.445 1334.940 ;
        RECT 2397.035 1334.100 2397.205 1334.610 ;
        RECT 2397.035 1333.770 2397.445 1334.100 ;
        RECT 2397.035 1333.570 2397.205 1333.770 ;
        RECT 2392.805 1332.310 2392.980 1333.450 ;
        RECT 2397.035 1332.310 2397.210 1333.570 ;
        RECT 2397.620 1333.540 2397.790 1335.150 ;
        RECT 2397.990 1335.090 2398.165 1335.600 ;
        RECT 2398.420 1335.050 2398.595 1335.600 ;
        RECT 2399.785 1335.090 2399.955 1335.600 ;
        RECT 2400.775 1335.090 2400.945 1335.600 ;
        RECT 2406.680 1335.110 2406.855 1335.600 ;
        RECT 2397.560 1333.370 2397.790 1333.540 ;
        RECT 2397.990 1333.570 2398.160 1334.520 ;
        RECT 2397.560 1332.310 2397.730 1333.370 ;
        RECT 2397.990 1332.310 2398.165 1333.570 ;
        RECT 2398.420 1333.450 2398.590 1335.050 ;
        RECT 2406.680 1334.940 2406.850 1335.110 ;
        RECT 2407.635 1335.090 2407.810 1335.600 ;
        RECT 2408.065 1335.050 2408.240 1335.600 ;
        RECT 2412.295 1335.110 2412.470 1335.600 ;
        RECT 2412.820 1335.320 2412.990 1335.600 ;
        RECT 2412.820 1335.150 2413.050 1335.320 ;
        RECT 2406.680 1334.610 2407.090 1334.940 ;
        RECT 2399.350 1334.430 2399.580 1334.585 ;
        RECT 2399.350 1334.355 2399.880 1334.430 ;
        RECT 2399.410 1334.260 2399.880 1334.355 ;
        RECT 2400.400 1334.260 2400.870 1334.430 ;
        RECT 2399.410 1333.570 2399.580 1334.260 ;
        RECT 2399.780 1333.810 2399.950 1333.890 ;
        RECT 2400.400 1333.810 2400.570 1334.260 ;
        RECT 2406.680 1334.100 2406.850 1334.610 ;
        RECT 2399.780 1333.610 2400.570 1333.810 ;
        RECT 2398.420 1332.310 2398.595 1333.450 ;
        RECT 2399.780 1332.310 2399.955 1333.610 ;
        RECT 2400.400 1333.570 2400.570 1333.610 ;
        RECT 2400.770 1333.455 2400.940 1333.890 ;
        RECT 2406.680 1333.770 2407.090 1334.100 ;
        RECT 2406.680 1333.570 2406.850 1333.770 ;
        RECT 2407.635 1333.570 2407.805 1334.520 ;
        RECT 2400.770 1332.310 2400.945 1333.455 ;
        RECT 2406.680 1332.310 2406.855 1333.570 ;
        RECT 2407.635 1332.310 2407.810 1333.570 ;
        RECT 2408.065 1333.450 2408.235 1335.050 ;
        RECT 2412.295 1334.940 2412.465 1335.110 ;
        RECT 2412.295 1334.610 2412.705 1334.940 ;
        RECT 2412.295 1334.100 2412.465 1334.610 ;
        RECT 2412.295 1333.770 2412.705 1334.100 ;
        RECT 2412.295 1333.570 2412.465 1333.770 ;
        RECT 2408.065 1332.310 2408.240 1333.450 ;
        RECT 2412.295 1332.310 2412.470 1333.570 ;
        RECT 2412.880 1333.540 2413.050 1335.150 ;
        RECT 2413.250 1335.090 2413.425 1335.600 ;
        RECT 2413.680 1335.050 2413.855 1335.600 ;
        RECT 2415.045 1335.090 2415.215 1335.600 ;
        RECT 2416.035 1335.090 2416.205 1335.600 ;
        RECT 2421.940 1335.110 2422.115 1335.600 ;
        RECT 2412.820 1333.370 2413.050 1333.540 ;
        RECT 2413.250 1333.570 2413.420 1334.520 ;
        RECT 2412.820 1332.310 2412.990 1333.370 ;
        RECT 2413.250 1332.310 2413.425 1333.570 ;
        RECT 2413.680 1333.450 2413.850 1335.050 ;
        RECT 2421.940 1334.940 2422.110 1335.110 ;
        RECT 2422.895 1335.090 2423.070 1335.600 ;
        RECT 2423.325 1335.050 2423.500 1335.600 ;
        RECT 2427.555 1335.110 2427.730 1335.600 ;
        RECT 2428.080 1335.320 2428.250 1335.600 ;
        RECT 2428.080 1335.150 2428.310 1335.320 ;
        RECT 2421.940 1334.610 2422.350 1334.940 ;
        RECT 2414.610 1334.430 2414.840 1334.585 ;
        RECT 2414.610 1334.355 2415.140 1334.430 ;
        RECT 2414.670 1334.260 2415.140 1334.355 ;
        RECT 2415.660 1334.260 2416.130 1334.430 ;
        RECT 2414.670 1333.570 2414.840 1334.260 ;
        RECT 2415.040 1333.810 2415.210 1333.890 ;
        RECT 2415.660 1333.810 2415.830 1334.260 ;
        RECT 2421.940 1334.100 2422.110 1334.610 ;
        RECT 2415.040 1333.610 2415.830 1333.810 ;
        RECT 2413.680 1332.310 2413.855 1333.450 ;
        RECT 2415.040 1332.310 2415.215 1333.610 ;
        RECT 2415.660 1333.570 2415.830 1333.610 ;
        RECT 2416.030 1333.455 2416.200 1333.890 ;
        RECT 2421.940 1333.770 2422.350 1334.100 ;
        RECT 2421.940 1333.570 2422.110 1333.770 ;
        RECT 2422.895 1333.570 2423.065 1334.520 ;
        RECT 2416.030 1332.310 2416.205 1333.455 ;
        RECT 2421.940 1332.310 2422.115 1333.570 ;
        RECT 2422.895 1332.310 2423.070 1333.570 ;
        RECT 2423.325 1333.450 2423.495 1335.050 ;
        RECT 2427.555 1334.940 2427.725 1335.110 ;
        RECT 2427.555 1334.610 2427.965 1334.940 ;
        RECT 2427.555 1334.100 2427.725 1334.610 ;
        RECT 2427.555 1333.770 2427.965 1334.100 ;
        RECT 2427.555 1333.570 2427.725 1333.770 ;
        RECT 2423.325 1332.310 2423.500 1333.450 ;
        RECT 2427.555 1332.310 2427.730 1333.570 ;
        RECT 2428.140 1333.540 2428.310 1335.150 ;
        RECT 2428.510 1335.090 2428.685 1335.600 ;
        RECT 2428.940 1335.050 2429.115 1335.600 ;
        RECT 2430.305 1335.090 2430.475 1335.600 ;
        RECT 2431.295 1335.090 2431.465 1335.600 ;
        RECT 2437.200 1335.110 2437.375 1335.600 ;
        RECT 2428.080 1333.370 2428.310 1333.540 ;
        RECT 2428.510 1333.570 2428.680 1334.520 ;
        RECT 2428.080 1332.310 2428.250 1333.370 ;
        RECT 2428.510 1332.310 2428.685 1333.570 ;
        RECT 2428.940 1333.450 2429.110 1335.050 ;
        RECT 2437.200 1334.940 2437.370 1335.110 ;
        RECT 2438.155 1335.090 2438.330 1335.600 ;
        RECT 2438.585 1335.050 2438.760 1335.600 ;
        RECT 2442.815 1335.110 2442.990 1335.600 ;
        RECT 2443.340 1335.320 2443.510 1335.600 ;
        RECT 2443.340 1335.150 2443.570 1335.320 ;
        RECT 2437.200 1334.610 2437.610 1334.940 ;
        RECT 2429.870 1334.430 2430.100 1334.585 ;
        RECT 2429.870 1334.355 2430.400 1334.430 ;
        RECT 2429.930 1334.260 2430.400 1334.355 ;
        RECT 2430.920 1334.260 2431.390 1334.430 ;
        RECT 2429.930 1333.570 2430.100 1334.260 ;
        RECT 2430.300 1333.810 2430.470 1333.890 ;
        RECT 2430.920 1333.810 2431.090 1334.260 ;
        RECT 2437.200 1334.100 2437.370 1334.610 ;
        RECT 2430.300 1333.610 2431.090 1333.810 ;
        RECT 2428.940 1332.310 2429.115 1333.450 ;
        RECT 2430.300 1332.310 2430.475 1333.610 ;
        RECT 2430.920 1333.570 2431.090 1333.610 ;
        RECT 2431.290 1333.455 2431.460 1333.890 ;
        RECT 2437.200 1333.770 2437.610 1334.100 ;
        RECT 2437.200 1333.570 2437.370 1333.770 ;
        RECT 2438.155 1333.570 2438.325 1334.520 ;
        RECT 2431.290 1332.310 2431.465 1333.455 ;
        RECT 2437.200 1332.310 2437.375 1333.570 ;
        RECT 2438.155 1332.310 2438.330 1333.570 ;
        RECT 2438.585 1333.450 2438.755 1335.050 ;
        RECT 2442.815 1334.940 2442.985 1335.110 ;
        RECT 2442.815 1334.610 2443.225 1334.940 ;
        RECT 2442.815 1334.100 2442.985 1334.610 ;
        RECT 2442.815 1333.770 2443.225 1334.100 ;
        RECT 2442.815 1333.570 2442.985 1333.770 ;
        RECT 2438.585 1332.310 2438.760 1333.450 ;
        RECT 2442.815 1332.310 2442.990 1333.570 ;
        RECT 2443.400 1333.540 2443.570 1335.150 ;
        RECT 2443.770 1335.090 2443.945 1335.600 ;
        RECT 2444.200 1335.050 2444.375 1335.600 ;
        RECT 2445.565 1335.090 2445.735 1335.600 ;
        RECT 2446.555 1335.090 2446.725 1335.600 ;
        RECT 2443.340 1333.370 2443.570 1333.540 ;
        RECT 2443.770 1333.570 2443.940 1334.520 ;
        RECT 2443.340 1332.310 2443.510 1333.370 ;
        RECT 2443.770 1332.310 2443.945 1333.570 ;
        RECT 2444.200 1333.450 2444.370 1335.050 ;
        RECT 2445.130 1334.430 2445.360 1334.585 ;
        RECT 2445.130 1334.355 2445.660 1334.430 ;
        RECT 2445.190 1334.260 2445.660 1334.355 ;
        RECT 2446.180 1334.260 2446.650 1334.430 ;
        RECT 2445.190 1333.570 2445.360 1334.260 ;
        RECT 2445.560 1333.810 2445.730 1333.890 ;
        RECT 2446.180 1333.810 2446.350 1334.260 ;
        RECT 2445.560 1333.610 2446.350 1333.810 ;
        RECT 2444.200 1332.310 2444.375 1333.450 ;
        RECT 2445.560 1332.310 2445.735 1333.610 ;
        RECT 2446.180 1333.570 2446.350 1333.610 ;
        RECT 2446.550 1333.455 2446.720 1333.890 ;
        RECT 2446.550 1332.310 2446.725 1333.455 ;
        RECT 2371.875 1329.435 2372.045 1329.795 ;
        RECT 2372.815 1329.435 2372.985 1329.795 ;
        RECT 2373.295 1329.345 2373.465 1329.765 ;
        RECT 2373.655 1329.515 2373.945 1330.075 ;
        RECT 2374.735 1329.775 2374.905 1330.105 ;
        RECT 2375.215 1329.685 2375.385 1330.075 ;
        RECT 2377.110 1329.775 2377.285 1330.105 ;
        RECT 2379.055 1329.905 2379.565 1330.075 ;
        RECT 2377.635 1329.685 2377.815 1329.795 ;
        RECT 2379.395 1329.765 2379.565 1329.905 ;
        RECT 2375.105 1329.515 2375.440 1329.685 ;
        RECT 2375.935 1329.515 2376.425 1329.685 ;
        RECT 2377.635 1329.515 2378.985 1329.685 ;
        RECT 2379.395 1329.515 2379.680 1329.765 ;
        RECT 2373.775 1329.435 2373.945 1329.515 ;
        RECT 2372.575 1328.785 2372.745 1329.235 ;
        RECT 2373.055 1328.785 2373.225 1329.115 ;
        RECT 2374.015 1328.785 2374.185 1329.115 ;
        RECT 2374.495 1328.785 2374.665 1329.515 ;
        RECT 2375.935 1329.345 2376.105 1329.515 ;
        RECT 2377.635 1329.435 2377.815 1329.515 ;
        RECT 2378.815 1329.345 2378.985 1329.515 ;
        RECT 2379.505 1329.435 2379.680 1329.515 ;
        RECT 2374.975 1328.785 2375.145 1329.235 ;
        RECT 2375.455 1328.785 2375.625 1329.115 ;
        RECT 2375.935 1328.785 2376.105 1329.115 ;
        RECT 2376.415 1328.785 2376.585 1329.235 ;
        RECT 2377.375 1329.135 2377.545 1329.235 ;
        RECT 2376.895 1329.035 2377.545 1329.135 ;
        RECT 2376.815 1328.865 2377.625 1329.035 ;
        RECT 2377.855 1328.785 2378.025 1329.115 ;
        RECT 2378.335 1328.785 2378.505 1329.235 ;
        RECT 2378.815 1328.785 2378.985 1329.115 ;
        RECT 2379.295 1329.035 2379.565 1329.235 ;
        RECT 2379.175 1328.825 2379.565 1329.035 ;
        RECT 2381.775 1328.895 2381.950 1330.155 ;
        RECT 2382.300 1329.095 2382.470 1330.155 ;
        RECT 2382.300 1328.925 2382.530 1329.095 ;
        RECT 2381.775 1328.695 2381.945 1328.895 ;
        RECT 2376.895 1328.615 2377.065 1328.655 ;
        RECT 2376.535 1328.445 2377.065 1328.615 ;
        RECT 2371.875 1328.045 2372.045 1328.395 ;
        RECT 2373.775 1328.045 2373.945 1328.395 ;
        RECT 2375.175 1328.375 2375.345 1328.395 ;
        RECT 2375.175 1328.345 2375.385 1328.375 ;
        RECT 2375.075 1328.125 2375.385 1328.345 ;
        RECT 2375.215 1328.045 2375.385 1328.125 ;
        RECT 2376.175 1328.275 2376.345 1328.395 ;
        RECT 2376.175 1328.105 2377.415 1328.275 ;
        RECT 2378.095 1328.045 2378.265 1328.395 ;
        RECT 2379.055 1328.045 2379.225 1328.395 ;
        RECT 2381.775 1328.365 2382.185 1328.695 ;
        RECT 2381.775 1327.855 2381.945 1328.365 ;
        RECT 2381.775 1327.525 2382.185 1327.855 ;
        RECT 2381.775 1327.355 2381.945 1327.525 ;
        RECT 2381.775 1326.865 2381.950 1327.355 ;
        RECT 2382.360 1327.315 2382.530 1328.925 ;
        RECT 2382.730 1328.895 2382.905 1330.155 ;
        RECT 2383.160 1329.015 2383.335 1330.155 ;
        RECT 2382.730 1327.945 2382.900 1328.895 ;
        RECT 2383.160 1327.415 2383.330 1329.015 ;
        RECT 2384.520 1329.010 2384.695 1330.155 ;
        RECT 2385.505 1329.010 2385.680 1330.155 ;
        RECT 2387.135 1329.435 2387.305 1329.795 ;
        RECT 2388.075 1329.435 2388.245 1329.795 ;
        RECT 2388.555 1329.345 2388.725 1329.765 ;
        RECT 2388.915 1329.515 2389.205 1330.075 ;
        RECT 2389.995 1329.775 2390.165 1330.105 ;
        RECT 2390.475 1329.685 2390.645 1330.075 ;
        RECT 2392.370 1329.775 2392.545 1330.105 ;
        RECT 2394.315 1329.905 2394.825 1330.075 ;
        RECT 2392.895 1329.685 2393.075 1329.795 ;
        RECT 2394.655 1329.765 2394.825 1329.905 ;
        RECT 2390.365 1329.515 2390.700 1329.685 ;
        RECT 2391.195 1329.515 2391.685 1329.685 ;
        RECT 2392.895 1329.515 2394.245 1329.685 ;
        RECT 2394.655 1329.515 2394.940 1329.765 ;
        RECT 2389.035 1329.435 2389.205 1329.515 ;
        RECT 2384.150 1328.205 2384.320 1328.895 ;
        RECT 2384.520 1328.820 2384.690 1329.010 ;
        RECT 2385.135 1328.820 2385.305 1328.895 ;
        RECT 2384.520 1328.625 2385.305 1328.820 ;
        RECT 2384.520 1328.575 2384.690 1328.625 ;
        RECT 2385.135 1328.205 2385.305 1328.625 ;
        RECT 2385.505 1328.575 2385.675 1329.010 ;
        RECT 2387.835 1328.785 2388.005 1329.235 ;
        RECT 2388.315 1328.785 2388.485 1329.115 ;
        RECT 2389.275 1328.785 2389.445 1329.115 ;
        RECT 2389.755 1328.785 2389.925 1329.515 ;
        RECT 2391.195 1329.345 2391.365 1329.515 ;
        RECT 2392.895 1329.435 2393.075 1329.515 ;
        RECT 2394.075 1329.345 2394.245 1329.515 ;
        RECT 2394.765 1329.435 2394.940 1329.515 ;
        RECT 2390.235 1328.785 2390.405 1329.235 ;
        RECT 2390.715 1328.785 2390.885 1329.115 ;
        RECT 2391.195 1328.785 2391.365 1329.115 ;
        RECT 2391.675 1328.785 2391.845 1329.235 ;
        RECT 2392.635 1329.135 2392.805 1329.235 ;
        RECT 2392.155 1329.035 2392.805 1329.135 ;
        RECT 2392.075 1328.865 2392.885 1329.035 ;
        RECT 2393.115 1328.785 2393.285 1329.115 ;
        RECT 2393.595 1328.785 2393.765 1329.235 ;
        RECT 2394.075 1328.785 2394.245 1329.115 ;
        RECT 2394.555 1329.035 2394.825 1329.235 ;
        RECT 2394.435 1328.825 2394.825 1329.035 ;
        RECT 2397.035 1328.895 2397.210 1330.155 ;
        RECT 2397.560 1329.095 2397.730 1330.155 ;
        RECT 2397.560 1328.925 2397.790 1329.095 ;
        RECT 2397.035 1328.695 2397.205 1328.895 ;
        RECT 2392.155 1328.615 2392.325 1328.655 ;
        RECT 2391.795 1328.445 2392.325 1328.615 ;
        RECT 2384.150 1328.170 2384.620 1328.205 ;
        RECT 2384.090 1328.035 2384.620 1328.170 ;
        RECT 2385.135 1328.035 2385.605 1328.205 ;
        RECT 2387.135 1328.045 2387.305 1328.395 ;
        RECT 2389.035 1328.045 2389.205 1328.395 ;
        RECT 2390.435 1328.375 2390.605 1328.395 ;
        RECT 2390.435 1328.345 2390.645 1328.375 ;
        RECT 2390.335 1328.125 2390.645 1328.345 ;
        RECT 2390.475 1328.045 2390.645 1328.125 ;
        RECT 2391.435 1328.275 2391.605 1328.395 ;
        RECT 2391.435 1328.105 2392.675 1328.275 ;
        RECT 2393.355 1328.045 2393.525 1328.395 ;
        RECT 2394.315 1328.045 2394.485 1328.395 ;
        RECT 2397.035 1328.365 2397.445 1328.695 ;
        RECT 2384.090 1327.940 2384.320 1328.035 ;
        RECT 2397.035 1327.855 2397.205 1328.365 ;
        RECT 2397.035 1327.525 2397.445 1327.855 ;
        RECT 2382.300 1327.145 2382.530 1327.315 ;
        RECT 2382.300 1326.865 2382.470 1327.145 ;
        RECT 2382.730 1326.865 2382.905 1327.375 ;
        RECT 2383.160 1326.865 2383.335 1327.415 ;
        RECT 2384.525 1326.865 2384.695 1327.375 ;
        RECT 2385.510 1326.865 2385.680 1327.375 ;
        RECT 2397.035 1327.355 2397.205 1327.525 ;
        RECT 2397.035 1326.865 2397.210 1327.355 ;
        RECT 2397.620 1327.315 2397.790 1328.925 ;
        RECT 2397.990 1328.895 2398.165 1330.155 ;
        RECT 2398.420 1329.015 2398.595 1330.155 ;
        RECT 2397.990 1327.945 2398.160 1328.895 ;
        RECT 2398.420 1327.415 2398.590 1329.015 ;
        RECT 2399.780 1329.010 2399.955 1330.155 ;
        RECT 2400.765 1329.010 2400.940 1330.155 ;
        RECT 2402.395 1329.435 2402.565 1329.795 ;
        RECT 2403.335 1329.435 2403.505 1329.795 ;
        RECT 2403.815 1329.345 2403.985 1329.765 ;
        RECT 2404.175 1329.515 2404.465 1330.075 ;
        RECT 2405.255 1329.775 2405.425 1330.105 ;
        RECT 2405.735 1329.685 2405.905 1330.075 ;
        RECT 2407.630 1329.775 2407.805 1330.105 ;
        RECT 2409.575 1329.905 2410.085 1330.075 ;
        RECT 2408.155 1329.685 2408.335 1329.795 ;
        RECT 2409.915 1329.765 2410.085 1329.905 ;
        RECT 2405.625 1329.515 2405.960 1329.685 ;
        RECT 2406.455 1329.515 2406.945 1329.685 ;
        RECT 2408.155 1329.515 2409.505 1329.685 ;
        RECT 2409.915 1329.515 2410.200 1329.765 ;
        RECT 2404.295 1329.435 2404.465 1329.515 ;
        RECT 2399.410 1328.205 2399.580 1328.895 ;
        RECT 2399.780 1328.820 2399.950 1329.010 ;
        RECT 2400.395 1328.820 2400.565 1328.895 ;
        RECT 2399.780 1328.625 2400.565 1328.820 ;
        RECT 2399.780 1328.575 2399.950 1328.625 ;
        RECT 2400.395 1328.205 2400.565 1328.625 ;
        RECT 2400.765 1328.575 2400.935 1329.010 ;
        RECT 2403.095 1328.785 2403.265 1329.235 ;
        RECT 2403.575 1328.785 2403.745 1329.115 ;
        RECT 2404.535 1328.785 2404.705 1329.115 ;
        RECT 2405.015 1328.785 2405.185 1329.515 ;
        RECT 2406.455 1329.345 2406.625 1329.515 ;
        RECT 2408.155 1329.435 2408.335 1329.515 ;
        RECT 2409.335 1329.345 2409.505 1329.515 ;
        RECT 2410.025 1329.435 2410.200 1329.515 ;
        RECT 2405.495 1328.785 2405.665 1329.235 ;
        RECT 2405.975 1328.785 2406.145 1329.115 ;
        RECT 2406.455 1328.785 2406.625 1329.115 ;
        RECT 2406.935 1328.785 2407.105 1329.235 ;
        RECT 2407.895 1329.135 2408.065 1329.235 ;
        RECT 2407.415 1329.035 2408.065 1329.135 ;
        RECT 2407.335 1328.865 2408.145 1329.035 ;
        RECT 2408.375 1328.785 2408.545 1329.115 ;
        RECT 2408.855 1328.785 2409.025 1329.235 ;
        RECT 2409.335 1328.785 2409.505 1329.115 ;
        RECT 2409.815 1329.035 2410.085 1329.235 ;
        RECT 2409.695 1328.825 2410.085 1329.035 ;
        RECT 2412.295 1328.895 2412.470 1330.155 ;
        RECT 2412.820 1329.095 2412.990 1330.155 ;
        RECT 2412.820 1328.925 2413.050 1329.095 ;
        RECT 2412.295 1328.695 2412.465 1328.895 ;
        RECT 2407.415 1328.615 2407.585 1328.655 ;
        RECT 2407.055 1328.445 2407.585 1328.615 ;
        RECT 2399.410 1328.170 2399.880 1328.205 ;
        RECT 2399.350 1328.035 2399.880 1328.170 ;
        RECT 2400.395 1328.035 2400.865 1328.205 ;
        RECT 2402.395 1328.045 2402.565 1328.395 ;
        RECT 2404.295 1328.045 2404.465 1328.395 ;
        RECT 2405.695 1328.375 2405.865 1328.395 ;
        RECT 2405.695 1328.345 2405.905 1328.375 ;
        RECT 2405.595 1328.125 2405.905 1328.345 ;
        RECT 2405.735 1328.045 2405.905 1328.125 ;
        RECT 2406.695 1328.275 2406.865 1328.395 ;
        RECT 2406.695 1328.105 2407.935 1328.275 ;
        RECT 2408.615 1328.045 2408.785 1328.395 ;
        RECT 2409.575 1328.045 2409.745 1328.395 ;
        RECT 2412.295 1328.365 2412.705 1328.695 ;
        RECT 2399.350 1327.940 2399.580 1328.035 ;
        RECT 2412.295 1327.855 2412.465 1328.365 ;
        RECT 2412.295 1327.525 2412.705 1327.855 ;
        RECT 2397.560 1327.145 2397.790 1327.315 ;
        RECT 2397.560 1326.865 2397.730 1327.145 ;
        RECT 2397.990 1326.865 2398.165 1327.375 ;
        RECT 2398.420 1326.865 2398.595 1327.415 ;
        RECT 2399.785 1326.865 2399.955 1327.375 ;
        RECT 2400.770 1326.865 2400.940 1327.375 ;
        RECT 2412.295 1327.355 2412.465 1327.525 ;
        RECT 2412.295 1326.865 2412.470 1327.355 ;
        RECT 2412.880 1327.315 2413.050 1328.925 ;
        RECT 2413.250 1328.895 2413.425 1330.155 ;
        RECT 2413.680 1329.015 2413.855 1330.155 ;
        RECT 2413.250 1327.945 2413.420 1328.895 ;
        RECT 2413.680 1327.415 2413.850 1329.015 ;
        RECT 2415.040 1329.010 2415.215 1330.155 ;
        RECT 2416.025 1329.010 2416.200 1330.155 ;
        RECT 2417.655 1329.435 2417.825 1329.795 ;
        RECT 2418.595 1329.435 2418.765 1329.795 ;
        RECT 2419.075 1329.345 2419.245 1329.765 ;
        RECT 2419.435 1329.515 2419.725 1330.075 ;
        RECT 2420.515 1329.775 2420.685 1330.105 ;
        RECT 2420.995 1329.685 2421.165 1330.075 ;
        RECT 2422.890 1329.775 2423.065 1330.105 ;
        RECT 2424.835 1329.905 2425.345 1330.075 ;
        RECT 2423.415 1329.685 2423.595 1329.795 ;
        RECT 2425.175 1329.765 2425.345 1329.905 ;
        RECT 2420.885 1329.515 2421.220 1329.685 ;
        RECT 2421.715 1329.515 2422.205 1329.685 ;
        RECT 2423.415 1329.515 2424.765 1329.685 ;
        RECT 2425.175 1329.515 2425.460 1329.765 ;
        RECT 2419.555 1329.435 2419.725 1329.515 ;
        RECT 2414.670 1328.205 2414.840 1328.895 ;
        RECT 2415.040 1328.820 2415.210 1329.010 ;
        RECT 2415.655 1328.820 2415.825 1328.895 ;
        RECT 2415.040 1328.625 2415.825 1328.820 ;
        RECT 2415.040 1328.575 2415.210 1328.625 ;
        RECT 2415.655 1328.205 2415.825 1328.625 ;
        RECT 2416.025 1328.575 2416.195 1329.010 ;
        RECT 2418.355 1328.785 2418.525 1329.235 ;
        RECT 2418.835 1328.785 2419.005 1329.115 ;
        RECT 2419.795 1328.785 2419.965 1329.115 ;
        RECT 2420.275 1328.785 2420.445 1329.515 ;
        RECT 2421.715 1329.345 2421.885 1329.515 ;
        RECT 2423.415 1329.435 2423.595 1329.515 ;
        RECT 2424.595 1329.345 2424.765 1329.515 ;
        RECT 2425.285 1329.435 2425.460 1329.515 ;
        RECT 2420.755 1328.785 2420.925 1329.235 ;
        RECT 2421.235 1328.785 2421.405 1329.115 ;
        RECT 2421.715 1328.785 2421.885 1329.115 ;
        RECT 2422.195 1328.785 2422.365 1329.235 ;
        RECT 2423.155 1329.135 2423.325 1329.235 ;
        RECT 2422.675 1329.035 2423.325 1329.135 ;
        RECT 2422.595 1328.865 2423.405 1329.035 ;
        RECT 2423.635 1328.785 2423.805 1329.115 ;
        RECT 2424.115 1328.785 2424.285 1329.235 ;
        RECT 2424.595 1328.785 2424.765 1329.115 ;
        RECT 2425.075 1329.035 2425.345 1329.235 ;
        RECT 2424.955 1328.825 2425.345 1329.035 ;
        RECT 2427.555 1328.895 2427.730 1330.155 ;
        RECT 2428.080 1329.095 2428.250 1330.155 ;
        RECT 2428.080 1328.925 2428.310 1329.095 ;
        RECT 2427.555 1328.695 2427.725 1328.895 ;
        RECT 2422.675 1328.615 2422.845 1328.655 ;
        RECT 2422.315 1328.445 2422.845 1328.615 ;
        RECT 2414.670 1328.170 2415.140 1328.205 ;
        RECT 2414.610 1328.035 2415.140 1328.170 ;
        RECT 2415.655 1328.035 2416.125 1328.205 ;
        RECT 2417.655 1328.045 2417.825 1328.395 ;
        RECT 2419.555 1328.045 2419.725 1328.395 ;
        RECT 2420.955 1328.375 2421.125 1328.395 ;
        RECT 2420.955 1328.345 2421.165 1328.375 ;
        RECT 2420.855 1328.125 2421.165 1328.345 ;
        RECT 2420.995 1328.045 2421.165 1328.125 ;
        RECT 2421.955 1328.275 2422.125 1328.395 ;
        RECT 2421.955 1328.105 2423.195 1328.275 ;
        RECT 2423.875 1328.045 2424.045 1328.395 ;
        RECT 2424.835 1328.045 2425.005 1328.395 ;
        RECT 2427.555 1328.365 2427.965 1328.695 ;
        RECT 2414.610 1327.940 2414.840 1328.035 ;
        RECT 2427.555 1327.855 2427.725 1328.365 ;
        RECT 2427.555 1327.525 2427.965 1327.855 ;
        RECT 2412.820 1327.145 2413.050 1327.315 ;
        RECT 2412.820 1326.865 2412.990 1327.145 ;
        RECT 2413.250 1326.865 2413.425 1327.375 ;
        RECT 2413.680 1326.865 2413.855 1327.415 ;
        RECT 2415.045 1326.865 2415.215 1327.375 ;
        RECT 2416.030 1326.865 2416.200 1327.375 ;
        RECT 2427.555 1327.355 2427.725 1327.525 ;
        RECT 2427.555 1326.865 2427.730 1327.355 ;
        RECT 2428.140 1327.315 2428.310 1328.925 ;
        RECT 2428.510 1328.895 2428.685 1330.155 ;
        RECT 2428.940 1329.015 2429.115 1330.155 ;
        RECT 2428.510 1327.945 2428.680 1328.895 ;
        RECT 2428.940 1327.415 2429.110 1329.015 ;
        RECT 2430.300 1329.010 2430.475 1330.155 ;
        RECT 2431.285 1329.010 2431.460 1330.155 ;
        RECT 2432.915 1329.435 2433.085 1329.795 ;
        RECT 2433.855 1329.435 2434.025 1329.795 ;
        RECT 2434.335 1329.345 2434.505 1329.765 ;
        RECT 2434.695 1329.515 2434.985 1330.075 ;
        RECT 2435.775 1329.775 2435.945 1330.105 ;
        RECT 2436.255 1329.685 2436.425 1330.075 ;
        RECT 2438.150 1329.775 2438.325 1330.105 ;
        RECT 2440.095 1329.905 2440.605 1330.075 ;
        RECT 2438.675 1329.685 2438.855 1329.795 ;
        RECT 2440.435 1329.765 2440.605 1329.905 ;
        RECT 2436.145 1329.515 2436.480 1329.685 ;
        RECT 2436.975 1329.515 2437.465 1329.685 ;
        RECT 2438.675 1329.515 2440.025 1329.685 ;
        RECT 2440.435 1329.515 2440.720 1329.765 ;
        RECT 2434.815 1329.435 2434.985 1329.515 ;
        RECT 2429.930 1328.205 2430.100 1328.895 ;
        RECT 2430.300 1328.820 2430.470 1329.010 ;
        RECT 2430.915 1328.820 2431.085 1328.895 ;
        RECT 2430.300 1328.625 2431.085 1328.820 ;
        RECT 2430.300 1328.575 2430.470 1328.625 ;
        RECT 2430.915 1328.205 2431.085 1328.625 ;
        RECT 2431.285 1328.575 2431.455 1329.010 ;
        RECT 2433.615 1328.785 2433.785 1329.235 ;
        RECT 2434.095 1328.785 2434.265 1329.115 ;
        RECT 2435.055 1328.785 2435.225 1329.115 ;
        RECT 2435.535 1328.785 2435.705 1329.515 ;
        RECT 2436.975 1329.345 2437.145 1329.515 ;
        RECT 2438.675 1329.435 2438.855 1329.515 ;
        RECT 2439.855 1329.345 2440.025 1329.515 ;
        RECT 2440.545 1329.435 2440.720 1329.515 ;
        RECT 2436.015 1328.785 2436.185 1329.235 ;
        RECT 2436.495 1328.785 2436.665 1329.115 ;
        RECT 2436.975 1328.785 2437.145 1329.115 ;
        RECT 2437.455 1328.785 2437.625 1329.235 ;
        RECT 2438.415 1329.135 2438.585 1329.235 ;
        RECT 2437.935 1329.035 2438.585 1329.135 ;
        RECT 2437.855 1328.865 2438.665 1329.035 ;
        RECT 2438.895 1328.785 2439.065 1329.115 ;
        RECT 2439.375 1328.785 2439.545 1329.235 ;
        RECT 2439.855 1328.785 2440.025 1329.115 ;
        RECT 2440.335 1329.035 2440.605 1329.235 ;
        RECT 2440.215 1328.825 2440.605 1329.035 ;
        RECT 2442.815 1328.895 2442.990 1330.155 ;
        RECT 2443.340 1329.095 2443.510 1330.155 ;
        RECT 2443.340 1328.925 2443.570 1329.095 ;
        RECT 2442.815 1328.695 2442.985 1328.895 ;
        RECT 2437.935 1328.615 2438.105 1328.655 ;
        RECT 2437.575 1328.445 2438.105 1328.615 ;
        RECT 2429.930 1328.170 2430.400 1328.205 ;
        RECT 2429.870 1328.035 2430.400 1328.170 ;
        RECT 2430.915 1328.035 2431.385 1328.205 ;
        RECT 2432.915 1328.045 2433.085 1328.395 ;
        RECT 2434.815 1328.045 2434.985 1328.395 ;
        RECT 2436.215 1328.375 2436.385 1328.395 ;
        RECT 2436.215 1328.345 2436.425 1328.375 ;
        RECT 2436.115 1328.125 2436.425 1328.345 ;
        RECT 2436.255 1328.045 2436.425 1328.125 ;
        RECT 2437.215 1328.275 2437.385 1328.395 ;
        RECT 2437.215 1328.105 2438.455 1328.275 ;
        RECT 2439.135 1328.045 2439.305 1328.395 ;
        RECT 2440.095 1328.045 2440.265 1328.395 ;
        RECT 2442.815 1328.365 2443.225 1328.695 ;
        RECT 2429.870 1327.940 2430.100 1328.035 ;
        RECT 2442.815 1327.855 2442.985 1328.365 ;
        RECT 2442.815 1327.525 2443.225 1327.855 ;
        RECT 2428.080 1327.145 2428.310 1327.315 ;
        RECT 2428.080 1326.865 2428.250 1327.145 ;
        RECT 2428.510 1326.865 2428.685 1327.375 ;
        RECT 2428.940 1326.865 2429.115 1327.415 ;
        RECT 2430.305 1326.865 2430.475 1327.375 ;
        RECT 2431.290 1326.865 2431.460 1327.375 ;
        RECT 2442.815 1327.355 2442.985 1327.525 ;
        RECT 2442.815 1326.865 2442.990 1327.355 ;
        RECT 2443.400 1327.315 2443.570 1328.925 ;
        RECT 2443.770 1328.895 2443.945 1330.155 ;
        RECT 2444.200 1329.015 2444.375 1330.155 ;
        RECT 2443.770 1327.945 2443.940 1328.895 ;
        RECT 2444.200 1327.415 2444.370 1329.015 ;
        RECT 2445.560 1329.010 2445.735 1330.155 ;
        RECT 2446.545 1329.010 2446.720 1330.155 ;
        RECT 2445.190 1328.205 2445.360 1328.895 ;
        RECT 2445.560 1328.820 2445.730 1329.010 ;
        RECT 2446.175 1328.820 2446.345 1328.895 ;
        RECT 2445.560 1328.625 2446.345 1328.820 ;
        RECT 2445.560 1328.575 2445.730 1328.625 ;
        RECT 2446.175 1328.205 2446.345 1328.625 ;
        RECT 2446.545 1328.575 2446.715 1329.010 ;
        RECT 2445.190 1328.170 2445.660 1328.205 ;
        RECT 2445.130 1328.035 2445.660 1328.170 ;
        RECT 2446.175 1328.035 2446.645 1328.205 ;
        RECT 2445.130 1327.940 2445.360 1328.035 ;
        RECT 2443.340 1327.145 2443.570 1327.315 ;
        RECT 2443.340 1326.865 2443.510 1327.145 ;
        RECT 2443.770 1326.865 2443.945 1327.375 ;
        RECT 2444.200 1326.865 2444.375 1327.415 ;
        RECT 2445.565 1326.865 2445.735 1327.375 ;
        RECT 2446.550 1326.865 2446.720 1327.375 ;
        RECT 2882.085 1162.180 2882.605 1163.730 ;
      LAYER met1 ;
        RECT 2359.550 2255.045 2359.840 2255.275 ;
        RECT 2362.780 2255.045 2363.070 2255.275 ;
        RECT 2374.005 2255.050 2374.295 2255.280 ;
        RECT 2359.610 2254.585 2359.780 2255.045 ;
        RECT 2362.840 2254.675 2363.010 2255.045 ;
        RECT 2359.520 2254.305 2359.860 2254.585 ;
        RECT 2362.740 2254.305 2363.110 2254.675 ;
        RECT 2374.065 2254.575 2374.235 2255.050 ;
        RECT 2375.795 2255.020 2376.090 2255.280 ;
        RECT 2376.785 2255.020 2377.080 2255.280 ;
        RECT 2379.365 2255.045 2379.655 2255.275 ;
        RECT 2390.590 2255.050 2390.880 2255.280 ;
        RECT 2374.975 2254.575 2375.325 2254.600 ;
        RECT 2374.065 2254.540 2375.325 2254.575 ;
        RECT 2374.005 2254.405 2375.325 2254.540 ;
        RECT 2374.005 2254.310 2374.295 2254.405 ;
        RECT 2374.975 2254.310 2375.325 2254.405 ;
        RECT 2363.240 2254.165 2363.580 2254.195 ;
        RECT 2374.460 2254.170 2374.785 2254.265 ;
        RECT 2363.210 2254.135 2363.580 2254.165 ;
        RECT 2374.435 2254.140 2374.785 2254.170 ;
        RECT 2363.040 2253.965 2363.580 2254.135 ;
        RECT 2374.265 2253.970 2374.785 2254.140 ;
        RECT 2363.210 2253.935 2363.580 2253.965 ;
        RECT 2374.435 2253.940 2374.785 2253.970 ;
        RECT 2363.240 2253.915 2363.580 2253.935 ;
        RECT 2375.855 2253.920 2376.025 2255.020 ;
        RECT 2376.845 2254.270 2377.015 2255.020 ;
        RECT 2379.425 2254.675 2379.595 2255.045 ;
        RECT 2379.325 2254.305 2379.695 2254.675 ;
        RECT 2390.650 2254.575 2390.820 2255.050 ;
        RECT 2392.380 2255.020 2392.675 2255.280 ;
        RECT 2393.370 2255.020 2393.665 2255.280 ;
        RECT 2395.950 2255.045 2396.240 2255.275 ;
        RECT 2407.175 2255.050 2407.465 2255.280 ;
        RECT 2391.560 2254.575 2391.910 2254.600 ;
        RECT 2390.650 2254.540 2391.910 2254.575 ;
        RECT 2390.590 2254.405 2391.910 2254.540 ;
        RECT 2390.590 2254.310 2390.880 2254.405 ;
        RECT 2391.560 2254.310 2391.910 2254.405 ;
        RECT 2376.845 2253.945 2377.175 2254.270 ;
        RECT 2379.825 2254.165 2380.165 2254.195 ;
        RECT 2391.045 2254.170 2391.370 2254.265 ;
        RECT 2379.795 2254.135 2380.165 2254.165 ;
        RECT 2391.020 2254.140 2391.370 2254.170 ;
        RECT 2379.625 2253.965 2380.165 2254.135 ;
        RECT 2390.850 2253.970 2391.370 2254.140 ;
        RECT 2376.845 2253.920 2377.135 2253.945 ;
        RECT 2379.795 2253.935 2380.165 2253.965 ;
        RECT 2391.020 2253.940 2391.370 2253.970 ;
        RECT 2375.795 2253.915 2376.025 2253.920 ;
        RECT 2359.145 2253.775 2359.485 2253.845 ;
        RECT 2373.660 2253.810 2373.980 2253.890 ;
        RECT 2373.635 2253.780 2373.980 2253.810 ;
        RECT 2359.005 2253.605 2359.485 2253.775 ;
        RECT 2373.460 2253.610 2373.980 2253.780 ;
        RECT 2375.795 2253.680 2376.085 2253.915 ;
        RECT 2376.785 2253.795 2377.135 2253.920 ;
        RECT 2379.825 2253.915 2380.165 2253.935 ;
        RECT 2392.440 2253.920 2392.610 2255.020 ;
        RECT 2393.430 2254.270 2393.600 2255.020 ;
        RECT 2396.010 2254.675 2396.180 2255.045 ;
        RECT 2395.910 2254.305 2396.280 2254.675 ;
        RECT 2407.235 2254.575 2407.405 2255.050 ;
        RECT 2408.965 2255.020 2409.260 2255.280 ;
        RECT 2409.955 2255.020 2410.250 2255.280 ;
        RECT 2412.535 2255.045 2412.825 2255.275 ;
        RECT 2423.760 2255.050 2424.050 2255.280 ;
        RECT 2408.145 2254.575 2408.495 2254.600 ;
        RECT 2407.235 2254.540 2408.495 2254.575 ;
        RECT 2407.175 2254.405 2408.495 2254.540 ;
        RECT 2407.175 2254.310 2407.465 2254.405 ;
        RECT 2408.145 2254.310 2408.495 2254.405 ;
        RECT 2393.430 2253.945 2393.760 2254.270 ;
        RECT 2396.410 2254.165 2396.750 2254.195 ;
        RECT 2407.630 2254.170 2407.955 2254.265 ;
        RECT 2396.380 2254.135 2396.750 2254.165 ;
        RECT 2407.605 2254.140 2407.955 2254.170 ;
        RECT 2396.210 2253.965 2396.750 2254.135 ;
        RECT 2407.435 2253.970 2407.955 2254.140 ;
        RECT 2393.430 2253.920 2393.720 2253.945 ;
        RECT 2396.380 2253.935 2396.750 2253.965 ;
        RECT 2407.605 2253.940 2407.955 2253.970 ;
        RECT 2392.380 2253.915 2392.610 2253.920 ;
        RECT 2390.245 2253.810 2390.565 2253.890 ;
        RECT 2376.785 2253.680 2377.075 2253.795 ;
        RECT 2390.220 2253.780 2390.565 2253.810 ;
        RECT 2390.045 2253.610 2390.565 2253.780 ;
        RECT 2392.380 2253.680 2392.670 2253.915 ;
        RECT 2393.370 2253.805 2393.720 2253.920 ;
        RECT 2396.410 2253.915 2396.750 2253.935 ;
        RECT 2409.025 2253.920 2409.195 2255.020 ;
        RECT 2410.015 2254.270 2410.185 2255.020 ;
        RECT 2412.595 2254.675 2412.765 2255.045 ;
        RECT 2412.495 2254.305 2412.865 2254.675 ;
        RECT 2423.820 2254.575 2423.990 2255.050 ;
        RECT 2425.550 2255.020 2425.845 2255.280 ;
        RECT 2426.540 2255.020 2426.835 2255.280 ;
        RECT 2429.115 2255.045 2429.405 2255.275 ;
        RECT 2440.340 2255.050 2440.630 2255.280 ;
        RECT 2424.730 2254.575 2425.080 2254.600 ;
        RECT 2423.820 2254.540 2425.080 2254.575 ;
        RECT 2423.760 2254.405 2425.080 2254.540 ;
        RECT 2423.760 2254.310 2424.050 2254.405 ;
        RECT 2424.730 2254.310 2425.080 2254.405 ;
        RECT 2410.015 2253.945 2410.345 2254.270 ;
        RECT 2412.995 2254.165 2413.335 2254.195 ;
        RECT 2424.215 2254.170 2424.540 2254.265 ;
        RECT 2412.965 2254.135 2413.335 2254.165 ;
        RECT 2424.190 2254.140 2424.540 2254.170 ;
        RECT 2412.795 2253.965 2413.335 2254.135 ;
        RECT 2424.020 2253.970 2424.540 2254.140 ;
        RECT 2410.015 2253.920 2410.305 2253.945 ;
        RECT 2412.965 2253.935 2413.335 2253.965 ;
        RECT 2424.190 2253.940 2424.540 2253.970 ;
        RECT 2408.965 2253.915 2409.195 2253.920 ;
        RECT 2406.830 2253.810 2407.150 2253.890 ;
        RECT 2393.370 2253.680 2393.660 2253.805 ;
        RECT 2406.805 2253.780 2407.150 2253.810 ;
        RECT 2406.630 2253.610 2407.150 2253.780 ;
        RECT 2408.965 2253.680 2409.255 2253.915 ;
        RECT 2409.955 2253.805 2410.305 2253.920 ;
        RECT 2412.995 2253.915 2413.335 2253.935 ;
        RECT 2425.610 2253.920 2425.780 2255.020 ;
        RECT 2426.600 2254.270 2426.770 2255.020 ;
        RECT 2429.175 2254.675 2429.345 2255.045 ;
        RECT 2429.075 2254.305 2429.445 2254.675 ;
        RECT 2440.400 2254.575 2440.570 2255.050 ;
        RECT 2442.130 2255.020 2442.425 2255.280 ;
        RECT 2443.120 2255.020 2443.415 2255.280 ;
        RECT 2441.310 2254.575 2441.660 2254.600 ;
        RECT 2440.400 2254.540 2441.660 2254.575 ;
        RECT 2440.340 2254.405 2441.660 2254.540 ;
        RECT 2440.340 2254.310 2440.630 2254.405 ;
        RECT 2441.310 2254.310 2441.660 2254.405 ;
        RECT 2426.600 2253.945 2426.930 2254.270 ;
        RECT 2429.575 2254.165 2429.915 2254.195 ;
        RECT 2440.795 2254.170 2441.120 2254.265 ;
        RECT 2429.545 2254.135 2429.915 2254.165 ;
        RECT 2440.770 2254.140 2441.120 2254.170 ;
        RECT 2429.375 2253.965 2429.915 2254.135 ;
        RECT 2440.600 2253.970 2441.120 2254.140 ;
        RECT 2426.600 2253.920 2426.890 2253.945 ;
        RECT 2429.545 2253.935 2429.915 2253.965 ;
        RECT 2440.770 2253.940 2441.120 2253.970 ;
        RECT 2425.550 2253.915 2425.780 2253.920 ;
        RECT 2423.415 2253.810 2423.735 2253.890 ;
        RECT 2409.955 2253.680 2410.245 2253.805 ;
        RECT 2423.390 2253.780 2423.735 2253.810 ;
        RECT 2423.215 2253.610 2423.735 2253.780 ;
        RECT 2425.550 2253.680 2425.840 2253.915 ;
        RECT 2426.540 2253.805 2426.890 2253.920 ;
        RECT 2429.575 2253.915 2429.915 2253.935 ;
        RECT 2442.190 2253.920 2442.360 2255.020 ;
        RECT 2443.150 2254.985 2443.415 2255.020 ;
        RECT 2443.150 2254.585 2443.475 2254.985 ;
        RECT 2443.180 2253.920 2443.350 2254.585 ;
        RECT 2442.130 2253.915 2442.360 2253.920 ;
        RECT 2443.120 2253.915 2443.350 2253.920 ;
        RECT 2439.995 2253.810 2440.315 2253.890 ;
        RECT 2426.540 2253.680 2426.830 2253.805 ;
        RECT 2439.970 2253.780 2440.315 2253.810 ;
        RECT 2439.795 2253.610 2440.315 2253.780 ;
        RECT 2442.130 2253.680 2442.420 2253.915 ;
        RECT 2443.120 2253.680 2443.410 2253.915 ;
        RECT 2359.145 2253.565 2359.485 2253.605 ;
        RECT 2373.635 2253.580 2373.980 2253.610 ;
        RECT 2390.220 2253.580 2390.565 2253.610 ;
        RECT 2406.805 2253.580 2407.150 2253.610 ;
        RECT 2423.390 2253.580 2423.735 2253.610 ;
        RECT 2439.970 2253.580 2440.315 2253.610 ;
        RECT 2373.660 2253.565 2373.980 2253.580 ;
        RECT 2390.245 2253.565 2390.565 2253.580 ;
        RECT 2406.830 2253.565 2407.150 2253.580 ;
        RECT 2423.415 2253.565 2423.735 2253.580 ;
        RECT 2439.995 2253.565 2440.315 2253.580 ;
        RECT 2366.920 2252.325 2367.210 2252.365 ;
        RECT 2367.590 2252.325 2367.910 2252.385 ;
        RECT 2366.920 2252.185 2367.910 2252.325 ;
        RECT 2366.920 2252.135 2367.210 2252.185 ;
        RECT 2367.590 2252.125 2367.910 2252.185 ;
        RECT 2368.610 2252.125 2368.930 2252.385 ;
        RECT 2369.300 2252.135 2369.590 2252.365 ;
        RECT 2369.970 2252.325 2370.290 2252.385 ;
        RECT 2383.505 2252.325 2383.795 2252.365 ;
        RECT 2384.175 2252.325 2384.495 2252.385 ;
        RECT 2369.970 2252.185 2370.560 2252.325 ;
        RECT 2383.505 2252.185 2384.495 2252.325 ;
        RECT 2367.680 2251.985 2367.820 2252.125 ;
        RECT 2369.380 2251.985 2369.520 2252.135 ;
        RECT 2369.970 2252.125 2370.290 2252.185 ;
        RECT 2383.505 2252.135 2383.795 2252.185 ;
        RECT 2384.175 2252.125 2384.495 2252.185 ;
        RECT 2385.195 2252.125 2385.515 2252.385 ;
        RECT 2385.885 2252.135 2386.175 2252.365 ;
        RECT 2386.555 2252.325 2386.875 2252.385 ;
        RECT 2400.090 2252.325 2400.380 2252.365 ;
        RECT 2400.760 2252.325 2401.080 2252.385 ;
        RECT 2386.555 2252.185 2387.145 2252.325 ;
        RECT 2400.090 2252.185 2401.080 2252.325 ;
        RECT 2367.680 2251.845 2369.520 2251.985 ;
        RECT 2384.265 2251.985 2384.405 2252.125 ;
        RECT 2385.965 2251.985 2386.105 2252.135 ;
        RECT 2386.555 2252.125 2386.875 2252.185 ;
        RECT 2400.090 2252.135 2400.380 2252.185 ;
        RECT 2400.760 2252.125 2401.080 2252.185 ;
        RECT 2401.780 2252.125 2402.100 2252.385 ;
        RECT 2402.470 2252.135 2402.760 2252.365 ;
        RECT 2403.140 2252.325 2403.460 2252.385 ;
        RECT 2416.675 2252.325 2416.965 2252.365 ;
        RECT 2417.345 2252.325 2417.665 2252.385 ;
        RECT 2403.140 2252.185 2403.730 2252.325 ;
        RECT 2416.675 2252.185 2417.665 2252.325 ;
        RECT 2384.265 2251.845 2386.105 2251.985 ;
        RECT 2400.850 2251.985 2400.990 2252.125 ;
        RECT 2402.550 2251.985 2402.690 2252.135 ;
        RECT 2403.140 2252.125 2403.460 2252.185 ;
        RECT 2416.675 2252.135 2416.965 2252.185 ;
        RECT 2417.345 2252.125 2417.665 2252.185 ;
        RECT 2418.365 2252.125 2418.685 2252.385 ;
        RECT 2419.055 2252.135 2419.345 2252.365 ;
        RECT 2419.725 2252.325 2420.045 2252.385 ;
        RECT 2433.255 2252.325 2433.545 2252.365 ;
        RECT 2433.925 2252.325 2434.245 2252.385 ;
        RECT 2419.725 2252.185 2420.315 2252.325 ;
        RECT 2433.255 2252.185 2434.245 2252.325 ;
        RECT 2400.850 2251.845 2402.690 2251.985 ;
        RECT 2417.435 2251.985 2417.575 2252.125 ;
        RECT 2419.135 2251.985 2419.275 2252.135 ;
        RECT 2419.725 2252.125 2420.045 2252.185 ;
        RECT 2433.255 2252.135 2433.545 2252.185 ;
        RECT 2433.925 2252.125 2434.245 2252.185 ;
        RECT 2434.945 2252.125 2435.265 2252.385 ;
        RECT 2435.635 2252.135 2435.925 2252.365 ;
        RECT 2436.305 2252.325 2436.625 2252.385 ;
        RECT 2436.305 2252.185 2436.895 2252.325 ;
        RECT 2417.435 2251.845 2419.275 2251.985 ;
        RECT 2434.015 2251.985 2434.155 2252.125 ;
        RECT 2435.715 2251.985 2435.855 2252.135 ;
        RECT 2436.305 2252.125 2436.625 2252.185 ;
        RECT 2434.015 2251.845 2435.855 2251.985 ;
        RECT 2365.220 2251.305 2365.510 2251.345 ;
        RECT 2367.930 2251.305 2368.250 2251.365 ;
        RECT 2365.220 2251.165 2368.250 2251.305 ;
        RECT 2365.220 2251.115 2365.510 2251.165 ;
        RECT 2367.930 2251.105 2368.250 2251.165 ;
        RECT 2370.660 2251.105 2371.310 2251.365 ;
        RECT 2381.805 2251.305 2382.095 2251.345 ;
        RECT 2384.515 2251.305 2384.835 2251.365 ;
        RECT 2381.805 2251.165 2384.835 2251.305 ;
        RECT 2381.805 2251.115 2382.095 2251.165 ;
        RECT 2384.515 2251.105 2384.835 2251.165 ;
        RECT 2387.245 2251.105 2387.895 2251.365 ;
        RECT 2398.390 2251.305 2398.680 2251.345 ;
        RECT 2401.100 2251.305 2401.420 2251.365 ;
        RECT 2398.390 2251.165 2401.420 2251.305 ;
        RECT 2398.390 2251.115 2398.680 2251.165 ;
        RECT 2401.100 2251.105 2401.420 2251.165 ;
        RECT 2403.830 2251.105 2404.480 2251.365 ;
        RECT 2414.975 2251.305 2415.265 2251.345 ;
        RECT 2417.685 2251.305 2418.005 2251.365 ;
        RECT 2414.975 2251.165 2418.005 2251.305 ;
        RECT 2414.975 2251.115 2415.265 2251.165 ;
        RECT 2417.685 2251.105 2418.005 2251.165 ;
        RECT 2420.415 2251.105 2421.065 2251.365 ;
        RECT 2431.555 2251.305 2431.845 2251.345 ;
        RECT 2434.265 2251.305 2434.585 2251.365 ;
        RECT 2431.555 2251.165 2434.585 2251.305 ;
        RECT 2431.555 2251.115 2431.845 2251.165 ;
        RECT 2434.265 2251.105 2434.585 2251.165 ;
        RECT 2436.995 2251.105 2437.645 2251.365 ;
        RECT 2366.410 2250.285 2366.700 2250.325 ;
        RECT 2368.620 2250.285 2368.910 2250.325 ;
        RECT 2369.290 2250.285 2369.610 2250.345 ;
        RECT 2366.410 2250.145 2369.610 2250.285 ;
        RECT 2366.410 2250.095 2366.700 2250.145 ;
        RECT 2368.620 2250.095 2368.910 2250.145 ;
        RECT 2369.290 2250.085 2369.610 2250.145 ;
        RECT 2382.995 2250.285 2383.285 2250.325 ;
        RECT 2385.205 2250.285 2385.495 2250.325 ;
        RECT 2385.875 2250.285 2386.195 2250.345 ;
        RECT 2382.995 2250.145 2386.195 2250.285 ;
        RECT 2382.995 2250.095 2383.285 2250.145 ;
        RECT 2385.205 2250.095 2385.495 2250.145 ;
        RECT 2385.875 2250.085 2386.195 2250.145 ;
        RECT 2399.580 2250.285 2399.870 2250.325 ;
        RECT 2401.790 2250.285 2402.080 2250.325 ;
        RECT 2402.460 2250.285 2402.780 2250.345 ;
        RECT 2399.580 2250.145 2402.780 2250.285 ;
        RECT 2399.580 2250.095 2399.870 2250.145 ;
        RECT 2401.790 2250.095 2402.080 2250.145 ;
        RECT 2402.460 2250.085 2402.780 2250.145 ;
        RECT 2416.165 2250.285 2416.455 2250.325 ;
        RECT 2418.375 2250.285 2418.665 2250.325 ;
        RECT 2419.045 2250.285 2419.365 2250.345 ;
        RECT 2416.165 2250.145 2419.365 2250.285 ;
        RECT 2416.165 2250.095 2416.455 2250.145 ;
        RECT 2418.375 2250.095 2418.665 2250.145 ;
        RECT 2419.045 2250.085 2419.365 2250.145 ;
        RECT 2432.745 2250.285 2433.035 2250.325 ;
        RECT 2434.955 2250.285 2435.245 2250.325 ;
        RECT 2435.625 2250.285 2435.945 2250.345 ;
        RECT 2432.745 2250.145 2435.945 2250.285 ;
        RECT 2432.745 2250.095 2433.035 2250.145 ;
        RECT 2434.955 2250.095 2435.245 2250.145 ;
        RECT 2435.625 2250.085 2435.945 2250.145 ;
        RECT 2368.610 2249.605 2368.930 2249.665 ;
        RECT 2370.580 2249.605 2370.870 2249.645 ;
        RECT 2371.405 2249.620 2371.730 2249.805 ;
        RECT 2371.305 2249.605 2371.730 2249.620 ;
        RECT 2368.610 2249.480 2371.730 2249.605 ;
        RECT 2385.195 2249.605 2385.515 2249.665 ;
        RECT 2387.165 2249.605 2387.455 2249.645 ;
        RECT 2387.990 2249.620 2388.315 2249.805 ;
        RECT 2387.890 2249.605 2388.315 2249.620 ;
        RECT 2385.195 2249.480 2388.315 2249.605 ;
        RECT 2401.780 2249.605 2402.100 2249.665 ;
        RECT 2403.750 2249.605 2404.040 2249.645 ;
        RECT 2404.575 2249.620 2404.900 2249.805 ;
        RECT 2404.475 2249.605 2404.900 2249.620 ;
        RECT 2401.780 2249.480 2404.900 2249.605 ;
        RECT 2418.365 2249.605 2418.685 2249.665 ;
        RECT 2420.335 2249.605 2420.625 2249.645 ;
        RECT 2421.160 2249.620 2421.485 2249.805 ;
        RECT 2421.060 2249.605 2421.485 2249.620 ;
        RECT 2418.365 2249.480 2421.485 2249.605 ;
        RECT 2434.945 2249.605 2435.265 2249.665 ;
        RECT 2436.915 2249.605 2437.205 2249.645 ;
        RECT 2437.740 2249.620 2438.065 2249.805 ;
        RECT 2437.640 2249.605 2438.065 2249.620 ;
        RECT 2434.945 2249.480 2438.065 2249.605 ;
        RECT 2368.610 2249.465 2371.445 2249.480 ;
        RECT 2385.195 2249.465 2388.030 2249.480 ;
        RECT 2401.780 2249.465 2404.615 2249.480 ;
        RECT 2418.365 2249.465 2421.200 2249.480 ;
        RECT 2434.945 2249.465 2437.780 2249.480 ;
        RECT 2368.610 2249.405 2368.930 2249.465 ;
        RECT 2370.580 2249.415 2370.870 2249.465 ;
        RECT 2385.195 2249.405 2385.515 2249.465 ;
        RECT 2387.165 2249.415 2387.455 2249.465 ;
        RECT 2401.780 2249.405 2402.100 2249.465 ;
        RECT 2403.750 2249.415 2404.040 2249.465 ;
        RECT 2418.365 2249.405 2418.685 2249.465 ;
        RECT 2420.335 2249.415 2420.625 2249.465 ;
        RECT 2434.945 2249.405 2435.265 2249.465 ;
        RECT 2436.915 2249.415 2437.205 2249.465 ;
        RECT 2364.250 2249.265 2364.540 2249.305 ;
        RECT 2366.985 2249.265 2367.855 2249.295 ;
        RECT 2369.290 2249.265 2369.610 2249.325 ;
        RECT 2370.990 2249.265 2371.310 2249.325 ;
        RECT 2364.250 2249.155 2369.610 2249.265 ;
        RECT 2364.250 2249.125 2367.125 2249.155 ;
        RECT 2367.715 2249.125 2369.610 2249.155 ;
        RECT 2370.710 2249.125 2371.310 2249.265 ;
        RECT 2364.250 2249.075 2364.540 2249.125 ;
        RECT 2369.290 2249.065 2369.610 2249.125 ;
        RECT 2370.990 2249.065 2371.310 2249.125 ;
        RECT 2380.835 2249.265 2381.125 2249.305 ;
        RECT 2383.570 2249.265 2384.440 2249.295 ;
        RECT 2385.875 2249.265 2386.195 2249.325 ;
        RECT 2387.575 2249.265 2387.895 2249.325 ;
        RECT 2380.835 2249.155 2386.195 2249.265 ;
        RECT 2380.835 2249.125 2383.710 2249.155 ;
        RECT 2384.300 2249.125 2386.195 2249.155 ;
        RECT 2387.295 2249.125 2387.895 2249.265 ;
        RECT 2380.835 2249.075 2381.125 2249.125 ;
        RECT 2385.875 2249.065 2386.195 2249.125 ;
        RECT 2387.575 2249.065 2387.895 2249.125 ;
        RECT 2397.420 2249.265 2397.710 2249.305 ;
        RECT 2400.155 2249.265 2401.025 2249.295 ;
        RECT 2402.460 2249.265 2402.780 2249.325 ;
        RECT 2404.160 2249.265 2404.480 2249.325 ;
        RECT 2397.420 2249.155 2402.780 2249.265 ;
        RECT 2397.420 2249.125 2400.295 2249.155 ;
        RECT 2400.885 2249.125 2402.780 2249.155 ;
        RECT 2403.880 2249.125 2404.480 2249.265 ;
        RECT 2397.420 2249.075 2397.710 2249.125 ;
        RECT 2402.460 2249.065 2402.780 2249.125 ;
        RECT 2404.160 2249.065 2404.480 2249.125 ;
        RECT 2414.005 2249.265 2414.295 2249.305 ;
        RECT 2416.740 2249.265 2417.610 2249.295 ;
        RECT 2419.045 2249.265 2419.365 2249.325 ;
        RECT 2420.745 2249.265 2421.065 2249.325 ;
        RECT 2414.005 2249.155 2419.365 2249.265 ;
        RECT 2414.005 2249.125 2416.880 2249.155 ;
        RECT 2417.470 2249.125 2419.365 2249.155 ;
        RECT 2420.465 2249.125 2421.065 2249.265 ;
        RECT 2414.005 2249.075 2414.295 2249.125 ;
        RECT 2419.045 2249.065 2419.365 2249.125 ;
        RECT 2420.745 2249.065 2421.065 2249.125 ;
        RECT 2430.585 2249.265 2430.875 2249.305 ;
        RECT 2433.320 2249.265 2434.190 2249.295 ;
        RECT 2435.625 2249.265 2435.945 2249.325 ;
        RECT 2437.325 2249.265 2437.645 2249.325 ;
        RECT 2430.585 2249.155 2435.945 2249.265 ;
        RECT 2430.585 2249.125 2433.460 2249.155 ;
        RECT 2434.050 2249.125 2435.945 2249.155 ;
        RECT 2437.045 2249.125 2437.645 2249.265 ;
        RECT 2430.585 2249.075 2430.875 2249.125 ;
        RECT 2435.625 2249.065 2435.945 2249.125 ;
        RECT 2437.325 2249.065 2437.645 2249.125 ;
        RECT 2367.250 2248.965 2367.570 2248.975 ;
        RECT 2366.580 2248.735 2366.870 2248.965 ;
        RECT 2367.250 2248.925 2367.710 2248.965 ;
        RECT 2367.930 2248.925 2368.250 2248.985 ;
        RECT 2369.380 2248.925 2369.520 2249.065 ;
        RECT 2367.250 2248.785 2367.730 2248.925 ;
        RECT 2367.930 2248.785 2368.520 2248.925 ;
        RECT 2369.380 2248.785 2369.860 2248.925 ;
        RECT 2373.660 2248.880 2373.980 2248.980 ;
        RECT 2383.835 2248.965 2384.155 2248.975 ;
        RECT 2373.635 2248.860 2373.980 2248.880 ;
        RECT 2367.250 2248.735 2367.710 2248.785 ;
        RECT 2366.660 2248.535 2366.800 2248.735 ;
        RECT 2367.250 2248.715 2367.570 2248.735 ;
        RECT 2367.930 2248.725 2368.250 2248.785 ;
        RECT 2368.980 2248.665 2369.240 2248.695 ;
        RECT 2368.950 2248.645 2369.270 2248.665 ;
        RECT 2369.720 2248.645 2369.860 2248.785 ;
        RECT 2373.345 2248.690 2373.980 2248.860 ;
        RECT 2373.460 2248.680 2373.980 2248.690 ;
        RECT 2373.635 2248.660 2373.980 2248.680 ;
        RECT 2373.635 2248.650 2373.925 2248.660 ;
        RECT 2368.850 2248.535 2369.270 2248.645 ;
        RECT 2366.660 2248.405 2369.270 2248.535 ;
        RECT 2369.640 2248.415 2369.930 2248.645 ;
        RECT 2371.990 2248.490 2372.315 2248.615 ;
        RECT 2374.435 2248.490 2374.785 2248.610 ;
        RECT 2375.795 2248.545 2376.085 2248.780 ;
        RECT 2376.785 2248.545 2377.075 2248.780 ;
        RECT 2383.165 2248.735 2383.455 2248.965 ;
        RECT 2383.835 2248.925 2384.295 2248.965 ;
        RECT 2384.515 2248.925 2384.835 2248.985 ;
        RECT 2385.965 2248.925 2386.105 2249.065 ;
        RECT 2383.835 2248.785 2384.315 2248.925 ;
        RECT 2384.515 2248.785 2385.105 2248.925 ;
        RECT 2385.965 2248.785 2386.445 2248.925 ;
        RECT 2390.245 2248.880 2390.565 2248.980 ;
        RECT 2400.420 2248.965 2400.740 2248.975 ;
        RECT 2390.220 2248.860 2390.565 2248.880 ;
        RECT 2383.835 2248.735 2384.295 2248.785 ;
        RECT 2375.795 2248.540 2376.025 2248.545 ;
        RECT 2376.785 2248.540 2377.015 2248.545 ;
        RECT 2366.660 2248.395 2368.910 2248.405 ;
        RECT 2371.990 2248.320 2374.785 2248.490 ;
        RECT 2371.990 2248.290 2372.315 2248.320 ;
        RECT 2374.435 2248.260 2374.785 2248.320 ;
        RECT 2374.005 2248.120 2374.295 2248.150 ;
        RECT 2374.975 2248.120 2375.325 2248.150 ;
        RECT 2374.005 2247.950 2375.325 2248.120 ;
        RECT 2374.005 2247.920 2374.295 2247.950 ;
        RECT 2374.065 2247.410 2374.235 2247.920 ;
        RECT 2374.975 2247.860 2375.325 2247.950 ;
        RECT 2375.855 2247.440 2376.025 2248.540 ;
        RECT 2376.845 2247.440 2377.015 2248.540 ;
        RECT 2383.245 2248.535 2383.385 2248.735 ;
        RECT 2383.835 2248.715 2384.155 2248.735 ;
        RECT 2384.515 2248.725 2384.835 2248.785 ;
        RECT 2385.565 2248.665 2385.825 2248.695 ;
        RECT 2385.535 2248.645 2385.855 2248.665 ;
        RECT 2386.305 2248.645 2386.445 2248.785 ;
        RECT 2389.930 2248.690 2390.565 2248.860 ;
        RECT 2390.045 2248.680 2390.565 2248.690 ;
        RECT 2390.220 2248.660 2390.565 2248.680 ;
        RECT 2390.220 2248.650 2390.510 2248.660 ;
        RECT 2385.435 2248.535 2385.855 2248.645 ;
        RECT 2383.245 2248.405 2385.855 2248.535 ;
        RECT 2386.225 2248.415 2386.515 2248.645 ;
        RECT 2388.575 2248.490 2388.900 2248.615 ;
        RECT 2391.020 2248.490 2391.370 2248.610 ;
        RECT 2392.380 2248.545 2392.670 2248.780 ;
        RECT 2393.370 2248.545 2393.660 2248.780 ;
        RECT 2399.750 2248.735 2400.040 2248.965 ;
        RECT 2400.420 2248.925 2400.880 2248.965 ;
        RECT 2401.100 2248.925 2401.420 2248.985 ;
        RECT 2402.550 2248.925 2402.690 2249.065 ;
        RECT 2400.420 2248.785 2400.900 2248.925 ;
        RECT 2401.100 2248.785 2401.690 2248.925 ;
        RECT 2402.550 2248.785 2403.030 2248.925 ;
        RECT 2406.830 2248.880 2407.150 2248.980 ;
        RECT 2417.005 2248.965 2417.325 2248.975 ;
        RECT 2406.805 2248.860 2407.150 2248.880 ;
        RECT 2400.420 2248.735 2400.880 2248.785 ;
        RECT 2392.380 2248.540 2392.610 2248.545 ;
        RECT 2393.370 2248.540 2393.600 2248.545 ;
        RECT 2383.245 2248.395 2385.495 2248.405 ;
        RECT 2388.575 2248.320 2391.370 2248.490 ;
        RECT 2388.575 2248.290 2388.900 2248.320 ;
        RECT 2391.020 2248.260 2391.370 2248.320 ;
        RECT 2390.590 2248.120 2390.880 2248.150 ;
        RECT 2391.560 2248.120 2391.910 2248.150 ;
        RECT 2390.590 2247.950 2391.910 2248.120 ;
        RECT 2390.590 2247.920 2390.880 2247.950 ;
        RECT 2374.005 2247.180 2374.295 2247.410 ;
        RECT 2375.795 2247.180 2376.090 2247.440 ;
        RECT 2376.785 2247.180 2377.210 2247.440 ;
        RECT 2390.650 2247.410 2390.820 2247.920 ;
        RECT 2391.560 2247.860 2391.910 2247.950 ;
        RECT 2392.440 2247.440 2392.610 2248.540 ;
        RECT 2393.430 2247.440 2393.600 2248.540 ;
        RECT 2399.830 2248.535 2399.970 2248.735 ;
        RECT 2400.420 2248.715 2400.740 2248.735 ;
        RECT 2401.100 2248.725 2401.420 2248.785 ;
        RECT 2402.150 2248.665 2402.410 2248.695 ;
        RECT 2402.120 2248.645 2402.440 2248.665 ;
        RECT 2402.890 2248.645 2403.030 2248.785 ;
        RECT 2406.515 2248.690 2407.150 2248.860 ;
        RECT 2406.630 2248.680 2407.150 2248.690 ;
        RECT 2406.805 2248.660 2407.150 2248.680 ;
        RECT 2406.805 2248.650 2407.095 2248.660 ;
        RECT 2402.020 2248.535 2402.440 2248.645 ;
        RECT 2399.830 2248.405 2402.440 2248.535 ;
        RECT 2402.810 2248.415 2403.100 2248.645 ;
        RECT 2405.160 2248.490 2405.485 2248.615 ;
        RECT 2407.605 2248.490 2407.955 2248.610 ;
        RECT 2408.965 2248.545 2409.255 2248.780 ;
        RECT 2409.955 2248.545 2410.245 2248.780 ;
        RECT 2416.335 2248.735 2416.625 2248.965 ;
        RECT 2417.005 2248.925 2417.465 2248.965 ;
        RECT 2417.685 2248.925 2418.005 2248.985 ;
        RECT 2419.135 2248.925 2419.275 2249.065 ;
        RECT 2417.005 2248.785 2417.485 2248.925 ;
        RECT 2417.685 2248.785 2418.275 2248.925 ;
        RECT 2419.135 2248.785 2419.615 2248.925 ;
        RECT 2423.415 2248.880 2423.735 2248.980 ;
        RECT 2433.585 2248.965 2433.905 2248.975 ;
        RECT 2423.390 2248.860 2423.735 2248.880 ;
        RECT 2417.005 2248.735 2417.465 2248.785 ;
        RECT 2408.965 2248.540 2409.195 2248.545 ;
        RECT 2409.955 2248.540 2410.185 2248.545 ;
        RECT 2399.830 2248.395 2402.080 2248.405 ;
        RECT 2405.160 2248.320 2407.955 2248.490 ;
        RECT 2405.160 2248.290 2405.485 2248.320 ;
        RECT 2407.605 2248.260 2407.955 2248.320 ;
        RECT 2407.175 2248.120 2407.465 2248.150 ;
        RECT 2408.145 2248.120 2408.495 2248.150 ;
        RECT 2407.175 2247.950 2408.495 2248.120 ;
        RECT 2407.175 2247.920 2407.465 2247.950 ;
        RECT 2390.590 2247.180 2390.880 2247.410 ;
        RECT 2392.380 2247.180 2392.675 2247.440 ;
        RECT 2393.370 2247.180 2393.770 2247.440 ;
        RECT 2407.235 2247.410 2407.405 2247.920 ;
        RECT 2408.145 2247.860 2408.495 2247.950 ;
        RECT 2409.025 2247.440 2409.195 2248.540 ;
        RECT 2410.015 2247.440 2410.185 2248.540 ;
        RECT 2416.415 2248.535 2416.555 2248.735 ;
        RECT 2417.005 2248.715 2417.325 2248.735 ;
        RECT 2417.685 2248.725 2418.005 2248.785 ;
        RECT 2418.735 2248.665 2418.995 2248.695 ;
        RECT 2418.705 2248.645 2419.025 2248.665 ;
        RECT 2419.475 2248.645 2419.615 2248.785 ;
        RECT 2423.100 2248.690 2423.735 2248.860 ;
        RECT 2423.215 2248.680 2423.735 2248.690 ;
        RECT 2423.390 2248.660 2423.735 2248.680 ;
        RECT 2423.390 2248.650 2423.680 2248.660 ;
        RECT 2418.605 2248.535 2419.025 2248.645 ;
        RECT 2416.415 2248.405 2419.025 2248.535 ;
        RECT 2419.395 2248.415 2419.685 2248.645 ;
        RECT 2421.745 2248.490 2422.070 2248.615 ;
        RECT 2424.190 2248.490 2424.540 2248.610 ;
        RECT 2425.550 2248.545 2425.840 2248.780 ;
        RECT 2426.540 2248.545 2426.830 2248.780 ;
        RECT 2432.915 2248.735 2433.205 2248.965 ;
        RECT 2433.585 2248.925 2434.045 2248.965 ;
        RECT 2434.265 2248.925 2434.585 2248.985 ;
        RECT 2435.715 2248.925 2435.855 2249.065 ;
        RECT 2433.585 2248.785 2434.065 2248.925 ;
        RECT 2434.265 2248.785 2434.855 2248.925 ;
        RECT 2435.715 2248.785 2436.195 2248.925 ;
        RECT 2439.995 2248.880 2440.315 2248.980 ;
        RECT 2439.970 2248.860 2440.315 2248.880 ;
        RECT 2433.585 2248.735 2434.045 2248.785 ;
        RECT 2425.550 2248.540 2425.780 2248.545 ;
        RECT 2426.540 2248.540 2426.770 2248.545 ;
        RECT 2416.415 2248.395 2418.665 2248.405 ;
        RECT 2421.745 2248.320 2424.540 2248.490 ;
        RECT 2421.745 2248.290 2422.070 2248.320 ;
        RECT 2424.190 2248.260 2424.540 2248.320 ;
        RECT 2423.760 2248.120 2424.050 2248.150 ;
        RECT 2424.730 2248.120 2425.080 2248.150 ;
        RECT 2423.760 2247.950 2425.080 2248.120 ;
        RECT 2423.760 2247.920 2424.050 2247.950 ;
        RECT 2407.175 2247.180 2407.465 2247.410 ;
        RECT 2408.965 2247.180 2409.260 2247.440 ;
        RECT 2409.955 2247.180 2410.330 2247.440 ;
        RECT 2423.820 2247.410 2423.990 2247.920 ;
        RECT 2424.730 2247.860 2425.080 2247.950 ;
        RECT 2425.610 2247.440 2425.780 2248.540 ;
        RECT 2426.600 2247.440 2426.770 2248.540 ;
        RECT 2432.995 2248.535 2433.135 2248.735 ;
        RECT 2433.585 2248.715 2433.905 2248.735 ;
        RECT 2434.265 2248.725 2434.585 2248.785 ;
        RECT 2435.315 2248.665 2435.575 2248.695 ;
        RECT 2435.285 2248.645 2435.605 2248.665 ;
        RECT 2436.055 2248.645 2436.195 2248.785 ;
        RECT 2439.680 2248.690 2440.315 2248.860 ;
        RECT 2439.795 2248.680 2440.315 2248.690 ;
        RECT 2439.970 2248.660 2440.315 2248.680 ;
        RECT 2439.970 2248.650 2440.260 2248.660 ;
        RECT 2435.185 2248.535 2435.605 2248.645 ;
        RECT 2432.995 2248.405 2435.605 2248.535 ;
        RECT 2435.975 2248.415 2436.265 2248.645 ;
        RECT 2438.325 2248.490 2438.650 2248.615 ;
        RECT 2440.770 2248.490 2441.120 2248.610 ;
        RECT 2442.130 2248.545 2442.420 2248.780 ;
        RECT 2443.120 2248.545 2443.410 2248.780 ;
        RECT 2442.130 2248.540 2442.360 2248.545 ;
        RECT 2443.120 2248.540 2443.350 2248.545 ;
        RECT 2432.995 2248.395 2435.245 2248.405 ;
        RECT 2438.325 2248.320 2441.120 2248.490 ;
        RECT 2438.325 2248.290 2438.650 2248.320 ;
        RECT 2440.770 2248.260 2441.120 2248.320 ;
        RECT 2440.340 2248.120 2440.630 2248.150 ;
        RECT 2441.310 2248.120 2441.660 2248.150 ;
        RECT 2440.340 2247.950 2441.660 2248.120 ;
        RECT 2440.340 2247.920 2440.630 2247.950 ;
        RECT 2423.760 2247.180 2424.050 2247.410 ;
        RECT 2425.550 2247.180 2425.845 2247.440 ;
        RECT 2426.540 2247.180 2426.890 2247.440 ;
        RECT 2440.400 2247.410 2440.570 2247.920 ;
        RECT 2441.310 2247.860 2441.660 2247.950 ;
        RECT 2442.190 2247.440 2442.360 2248.540 ;
        RECT 2443.180 2247.440 2443.350 2248.540 ;
        RECT 2440.340 2247.180 2440.630 2247.410 ;
        RECT 2442.130 2247.180 2442.425 2247.440 ;
        RECT 2443.120 2247.180 2443.415 2247.440 ;
        RECT 2443.220 2246.960 2443.360 2247.180 ;
        RECT 2459.690 2246.960 2460.010 2247.020 ;
        RECT 2443.220 2246.820 2460.010 2246.960 ;
        RECT 2459.690 2246.760 2460.010 2246.820 ;
        RECT 2393.450 2231.320 2393.770 2231.380 ;
        RECT 2393.450 2231.180 2401.270 2231.320 ;
        RECT 2393.450 2231.120 2393.770 2231.180 ;
        RECT 2401.130 2229.620 2401.270 2231.180 ;
        RECT 2576.990 2229.620 2577.310 2229.680 ;
        RECT 2401.130 2229.480 2577.310 2229.620 ;
        RECT 2576.990 2229.420 2577.310 2229.480 ;
        RECT 2410.010 2229.080 2410.330 2229.340 ;
        RECT 2426.570 2229.280 2426.890 2229.340 ;
        RECT 2618.390 2229.280 2618.710 2229.340 ;
        RECT 2426.570 2229.140 2618.710 2229.280 ;
        RECT 2426.570 2229.080 2426.890 2229.140 ;
        RECT 2618.390 2229.080 2618.710 2229.140 ;
        RECT 2410.100 2228.940 2410.240 2229.080 ;
        RECT 2604.590 2228.940 2604.910 2229.000 ;
        RECT 2410.100 2228.800 2604.910 2228.940 ;
        RECT 2604.590 2228.740 2604.910 2228.800 ;
        RECT 2376.890 2228.600 2377.210 2228.660 ;
        RECT 2677.270 2228.600 2677.590 2228.660 ;
        RECT 2376.890 2228.460 2677.590 2228.600 ;
        RECT 2376.890 2228.400 2377.210 2228.460 ;
        RECT 2677.270 2228.400 2677.590 2228.460 ;
        RECT 2695.590 2216.480 2695.910 2216.540 ;
        RECT 2698.810 2216.480 2699.130 2216.540 ;
        RECT 2700.205 2216.480 2700.495 2216.525 ;
        RECT 2695.590 2216.340 2698.120 2216.480 ;
        RECT 2695.590 2216.280 2695.910 2216.340 ;
        RECT 2697.980 2216.140 2698.120 2216.340 ;
        RECT 2698.810 2216.340 2700.495 2216.480 ;
        RECT 2698.810 2216.280 2699.130 2216.340 ;
        RECT 2700.205 2216.295 2700.495 2216.340 ;
        RECT 2702.490 2216.480 2702.810 2216.540 ;
        RECT 2709.865 2216.480 2710.155 2216.525 ;
        RECT 2702.490 2216.340 2710.155 2216.480 ;
        RECT 2702.490 2216.280 2702.810 2216.340 ;
        RECT 2709.865 2216.295 2710.155 2216.340 ;
        RECT 2697.980 2216.000 2701.340 2216.140 ;
        RECT 2695.130 2215.800 2695.450 2215.860 ;
        RECT 2701.200 2215.845 2701.340 2216.000 ;
        RECT 2699.745 2215.800 2700.035 2215.845 ;
        RECT 2695.130 2215.660 2700.035 2215.800 ;
        RECT 2695.130 2215.600 2695.450 2215.660 ;
        RECT 2699.745 2215.615 2700.035 2215.660 ;
        RECT 2701.125 2215.615 2701.415 2215.845 ;
        RECT 2698.365 2215.460 2698.655 2215.505 ;
        RECT 2701.570 2215.460 2701.890 2215.520 ;
        RECT 2698.365 2215.320 2701.890 2215.460 ;
        RECT 2698.365 2215.275 2698.655 2215.320 ;
        RECT 2701.570 2215.260 2701.890 2215.320 ;
        RECT 2452.790 2215.000 2453.110 2215.060 ;
        RECT 2677.270 2215.000 2677.590 2215.060 ;
        RECT 2452.790 2214.860 2677.590 2215.000 ;
        RECT 2721.810 2214.920 2722.130 2215.180 ;
        RECT 2452.790 2214.800 2453.110 2214.860 ;
        RECT 2677.270 2214.800 2677.590 2214.860 ;
        RECT 2698.350 2214.780 2698.670 2214.840 ;
        RECT 2698.825 2214.780 2699.115 2214.825 ;
        RECT 2698.350 2214.640 2699.115 2214.780 ;
        RECT 2698.350 2214.580 2698.670 2214.640 ;
        RECT 2698.825 2214.595 2699.115 2214.640 ;
        RECT 2731.470 2214.580 2731.790 2214.840 ;
        RECT 2694.670 2212.740 2694.990 2212.800 ;
        RECT 2696.985 2212.740 2697.275 2212.785 ;
        RECT 2694.670 2212.600 2697.275 2212.740 ;
        RECT 2694.670 2212.540 2694.990 2212.600 ;
        RECT 2696.985 2212.555 2697.275 2212.600 ;
        RECT 2697.890 2211.860 2698.210 2212.120 ;
        RECT 2466.590 2208.200 2466.910 2208.260 ;
        RECT 2677.270 2208.200 2677.590 2208.260 ;
        RECT 2466.590 2208.060 2677.590 2208.200 ;
        RECT 2466.590 2208.000 2466.910 2208.060 ;
        RECT 2677.270 2208.000 2677.590 2208.060 ;
        RECT 2694.670 2204.920 2694.990 2204.980 ;
        RECT 2696.985 2204.920 2697.275 2204.965 ;
        RECT 2694.670 2204.780 2697.275 2204.920 ;
        RECT 2694.670 2204.720 2694.990 2204.780 ;
        RECT 2696.985 2204.735 2697.275 2204.780 ;
        RECT 2696.970 2203.900 2697.290 2203.960 ;
        RECT 2697.905 2203.900 2698.195 2203.945 ;
        RECT 2696.970 2203.760 2698.195 2203.900 ;
        RECT 2696.970 2203.700 2697.290 2203.760 ;
        RECT 2697.905 2203.715 2698.195 2203.760 ;
        RECT 2697.430 2202.200 2697.750 2202.260 ;
        RECT 2698.350 2202.200 2698.670 2202.260 ;
        RECT 2697.430 2202.060 2698.670 2202.200 ;
        RECT 2697.430 2202.000 2697.750 2202.060 ;
        RECT 2698.350 2202.000 2698.670 2202.060 ;
        RECT 2473.490 2201.400 2473.810 2201.460 ;
        RECT 2677.270 2201.400 2677.590 2201.460 ;
        RECT 2473.490 2201.260 2677.590 2201.400 ;
        RECT 2473.490 2201.200 2473.810 2201.260 ;
        RECT 2677.270 2201.200 2677.590 2201.260 ;
        RECT 2698.370 2199.820 2698.660 2199.865 ;
        RECT 2703.890 2199.820 2704.180 2199.865 ;
        RECT 2704.810 2199.820 2705.100 2199.865 ;
        RECT 2698.370 2199.680 2705.100 2199.820 ;
        RECT 2698.370 2199.635 2698.660 2199.680 ;
        RECT 2703.890 2199.635 2704.180 2199.680 ;
        RECT 2704.810 2199.635 2705.100 2199.680 ;
        RECT 2696.985 2199.480 2697.275 2199.525 ;
        RECT 2697.430 2199.480 2697.750 2199.540 ;
        RECT 2696.985 2199.340 2697.750 2199.480 ;
        RECT 2696.985 2199.295 2697.275 2199.340 ;
        RECT 2697.430 2199.280 2697.750 2199.340 ;
        RECT 2697.890 2199.280 2698.210 2199.540 ;
        RECT 2699.290 2199.480 2699.580 2199.525 ;
        RECT 2701.130 2199.480 2701.420 2199.525 ;
        RECT 2699.290 2199.340 2701.420 2199.480 ;
        RECT 2699.290 2199.295 2699.580 2199.340 ;
        RECT 2701.130 2199.295 2701.420 2199.340 ;
        RECT 2703.475 2199.480 2703.765 2199.525 ;
        RECT 2705.315 2199.480 2705.605 2199.525 ;
        RECT 2703.475 2199.340 2705.605 2199.480 ;
        RECT 2703.475 2199.295 2703.765 2199.340 ;
        RECT 2705.315 2199.295 2705.605 2199.340 ;
        RECT 2721.810 2199.280 2722.130 2199.540 ;
        RECT 2702.030 2199.185 2702.350 2199.200 ;
        RECT 2701.585 2199.140 2701.875 2199.185 ;
        RECT 2697.520 2199.000 2701.875 2199.140 ;
        RECT 2697.520 2198.860 2697.660 2199.000 ;
        RECT 2701.585 2198.955 2701.875 2199.000 ;
        RECT 2702.030 2198.955 2702.460 2199.185 ;
        RECT 2702.950 2199.140 2703.270 2199.200 ;
        RECT 2721.900 2199.140 2722.040 2199.280 ;
        RECT 2702.950 2199.000 2722.040 2199.140 ;
        RECT 2702.030 2198.940 2702.350 2198.955 ;
        RECT 2702.950 2198.940 2703.270 2199.000 ;
        RECT 2697.430 2198.600 2697.750 2198.860 ;
        RECT 2700.205 2198.615 2700.495 2198.845 ;
        RECT 2701.165 2198.800 2701.455 2198.845 ;
        RECT 2704.395 2198.800 2704.685 2198.845 ;
        RECT 2701.165 2198.660 2704.685 2198.800 ;
        RECT 2701.165 2198.615 2701.455 2198.660 ;
        RECT 2704.395 2198.615 2704.685 2198.660 ;
        RECT 2700.280 2198.460 2700.420 2198.615 ;
        RECT 2702.490 2198.460 2702.810 2198.520 ;
        RECT 2700.280 2198.320 2702.810 2198.460 ;
        RECT 2702.490 2198.260 2702.810 2198.320 ;
        RECT 2703.870 2198.460 2704.190 2198.520 ;
        RECT 2706.185 2198.460 2706.475 2198.505 ;
        RECT 2703.870 2198.320 2706.475 2198.460 ;
        RECT 2703.870 2198.260 2704.190 2198.320 ;
        RECT 2706.185 2198.275 2706.475 2198.320 ;
        RECT 2697.905 2197.440 2698.195 2197.485 ;
        RECT 2702.030 2197.440 2702.350 2197.500 ;
        RECT 2697.905 2197.300 2702.350 2197.440 ;
        RECT 2697.905 2197.255 2698.195 2197.300 ;
        RECT 2702.030 2197.240 2702.350 2197.300 ;
        RECT 2694.670 2196.420 2694.990 2196.480 ;
        RECT 2696.985 2196.420 2697.275 2196.465 ;
        RECT 2694.670 2196.280 2697.275 2196.420 ;
        RECT 2694.670 2196.220 2694.990 2196.280 ;
        RECT 2696.985 2196.235 2697.275 2196.280 ;
        RECT 2480.390 2194.600 2480.710 2194.660 ;
        RECT 2677.270 2194.600 2677.590 2194.660 ;
        RECT 2480.390 2194.460 2677.590 2194.600 ;
        RECT 2480.390 2194.400 2480.710 2194.460 ;
        RECT 2677.270 2194.400 2677.590 2194.460 ;
        RECT 2698.370 2194.380 2698.660 2194.425 ;
        RECT 2703.890 2194.380 2704.180 2194.425 ;
        RECT 2704.810 2194.380 2705.100 2194.425 ;
        RECT 2698.370 2194.240 2705.100 2194.380 ;
        RECT 2698.370 2194.195 2698.660 2194.240 ;
        RECT 2703.890 2194.195 2704.180 2194.240 ;
        RECT 2704.810 2194.195 2705.100 2194.240 ;
        RECT 2696.970 2193.840 2697.290 2194.100 ;
        RECT 2697.890 2193.840 2698.210 2194.100 ;
        RECT 2699.290 2194.040 2699.580 2194.085 ;
        RECT 2701.130 2194.040 2701.420 2194.085 ;
        RECT 2699.290 2193.900 2701.420 2194.040 ;
        RECT 2699.290 2193.855 2699.580 2193.900 ;
        RECT 2701.130 2193.855 2701.420 2193.900 ;
        RECT 2702.950 2193.840 2703.270 2194.100 ;
        RECT 2703.475 2194.040 2703.765 2194.085 ;
        RECT 2705.315 2194.040 2705.605 2194.085 ;
        RECT 2703.475 2193.900 2705.605 2194.040 ;
        RECT 2703.475 2193.855 2703.765 2193.900 ;
        RECT 2705.315 2193.855 2705.605 2193.900 ;
        RECT 2698.810 2193.700 2699.130 2193.760 ;
        RECT 2702.030 2193.745 2702.350 2193.760 ;
        RECT 2701.585 2193.700 2701.875 2193.745 ;
        RECT 2698.810 2193.560 2701.875 2193.700 ;
        RECT 2698.810 2193.500 2699.130 2193.560 ;
        RECT 2701.585 2193.515 2701.875 2193.560 ;
        RECT 2702.030 2193.515 2702.460 2193.745 ;
        RECT 2702.030 2193.500 2702.350 2193.515 ;
        RECT 2700.205 2193.175 2700.495 2193.405 ;
        RECT 2701.165 2193.360 2701.455 2193.405 ;
        RECT 2704.395 2193.360 2704.685 2193.405 ;
        RECT 2701.165 2193.220 2704.685 2193.360 ;
        RECT 2701.165 2193.175 2701.455 2193.220 ;
        RECT 2704.395 2193.175 2704.685 2193.220 ;
        RECT 2698.350 2193.020 2698.670 2193.080 ;
        RECT 2700.280 2193.020 2700.420 2193.175 ;
        RECT 2702.490 2193.020 2702.810 2193.080 ;
        RECT 2698.350 2192.880 2702.810 2193.020 ;
        RECT 2698.350 2192.820 2698.670 2192.880 ;
        RECT 2702.490 2192.820 2702.810 2192.880 ;
        RECT 2706.170 2192.820 2706.490 2193.080 ;
        RECT 2697.905 2192.000 2698.195 2192.045 ;
        RECT 2702.030 2192.000 2702.350 2192.060 ;
        RECT 2706.170 2192.000 2706.490 2192.060 ;
        RECT 2697.905 2191.860 2702.350 2192.000 ;
        RECT 2697.905 2191.815 2698.195 2191.860 ;
        RECT 2702.030 2191.800 2702.350 2191.860 ;
        RECT 2703.960 2191.860 2706.490 2192.000 ;
        RECT 2697.890 2191.320 2698.210 2191.380 ;
        RECT 2701.570 2191.320 2701.890 2191.380 ;
        RECT 2703.960 2191.365 2704.100 2191.860 ;
        RECT 2706.170 2191.800 2706.490 2191.860 ;
        RECT 2697.890 2191.180 2703.640 2191.320 ;
        RECT 2697.890 2191.120 2698.210 2191.180 ;
        RECT 2701.570 2191.120 2701.890 2191.180 ;
        RECT 2694.670 2190.980 2694.990 2191.040 ;
        RECT 2696.985 2190.980 2697.275 2191.025 ;
        RECT 2694.670 2190.840 2697.275 2190.980 ;
        RECT 2703.500 2190.980 2703.640 2191.180 ;
        RECT 2703.885 2191.135 2704.175 2191.365 ;
        RECT 2704.345 2191.135 2704.635 2191.365 ;
        RECT 2704.420 2190.980 2704.560 2191.135 ;
        RECT 2703.500 2190.840 2704.560 2190.980 ;
        RECT 2694.670 2190.780 2694.990 2190.840 ;
        RECT 2696.985 2190.795 2697.275 2190.840 ;
        RECT 2703.425 2190.640 2703.715 2190.685 ;
        RECT 2703.870 2190.640 2704.190 2190.700 ;
        RECT 2703.425 2190.500 2704.190 2190.640 ;
        RECT 2703.425 2190.455 2703.715 2190.500 ;
        RECT 2703.870 2190.440 2704.190 2190.500 ;
        RECT 2701.570 2190.100 2701.890 2190.360 ;
        RECT 2487.290 2187.460 2487.610 2187.520 ;
        RECT 2677.270 2187.460 2677.590 2187.520 ;
        RECT 2487.290 2187.320 2677.590 2187.460 ;
        RECT 2487.290 2187.260 2487.610 2187.320 ;
        RECT 2677.270 2187.260 2677.590 2187.320 ;
        RECT 2697.430 2186.560 2697.750 2186.620 ;
        RECT 2697.905 2186.560 2698.195 2186.605 ;
        RECT 2697.430 2186.420 2698.195 2186.560 ;
        RECT 2697.430 2186.360 2697.750 2186.420 ;
        RECT 2697.905 2186.375 2698.195 2186.420 ;
        RECT 2694.670 2185.540 2694.990 2185.600 ;
        RECT 2696.985 2185.540 2697.275 2185.585 ;
        RECT 2694.670 2185.400 2697.275 2185.540 ;
        RECT 2694.670 2185.340 2694.990 2185.400 ;
        RECT 2696.985 2185.355 2697.275 2185.400 ;
        RECT 2494.190 2180.660 2494.510 2180.720 ;
        RECT 2677.270 2180.660 2677.590 2180.720 ;
        RECT 2494.190 2180.520 2677.590 2180.660 ;
        RECT 2494.190 2180.460 2494.510 2180.520 ;
        RECT 2677.270 2180.460 2677.590 2180.520 ;
        RECT 2701.570 2179.900 2701.890 2180.160 ;
        RECT 2702.505 2180.100 2702.795 2180.145 ;
        RECT 2703.870 2180.100 2704.190 2180.160 ;
        RECT 2731.470 2180.100 2731.790 2180.160 ;
        RECT 2702.505 2179.960 2731.790 2180.100 ;
        RECT 2702.505 2179.915 2702.795 2179.960 ;
        RECT 2703.870 2179.900 2704.190 2179.960 ;
        RECT 2731.470 2179.900 2731.790 2179.960 ;
        RECT 2702.030 2179.220 2702.350 2179.480 ;
        RECT 2697.905 2178.400 2698.195 2178.445 ;
        RECT 2698.810 2178.400 2699.130 2178.460 ;
        RECT 2697.905 2178.260 2699.130 2178.400 ;
        RECT 2697.905 2178.215 2698.195 2178.260 ;
        RECT 2698.810 2178.200 2699.130 2178.260 ;
        RECT 2702.030 2178.200 2702.350 2178.460 ;
        RECT 2703.870 2178.200 2704.190 2178.460 ;
        RECT 2694.670 2177.720 2694.990 2177.780 ;
        RECT 2702.120 2177.765 2702.260 2178.200 ;
        RECT 2703.960 2177.765 2704.100 2178.200 ;
        RECT 2696.985 2177.720 2697.275 2177.765 ;
        RECT 2694.670 2177.580 2697.275 2177.720 ;
        RECT 2694.670 2177.520 2694.990 2177.580 ;
        RECT 2696.985 2177.535 2697.275 2177.580 ;
        RECT 2702.045 2177.535 2702.335 2177.765 ;
        RECT 2703.885 2177.535 2704.175 2177.765 ;
        RECT 2704.790 2177.180 2705.110 2177.440 ;
        RECT 2702.490 2176.840 2702.810 2177.100 ;
        RECT 2702.490 2175.680 2702.810 2175.740 ;
        RECT 2702.490 2175.540 2724.570 2175.680 ;
        RECT 2702.490 2175.480 2702.810 2175.540 ;
        RECT 2724.430 2174.660 2724.570 2175.540 ;
        RECT 2725.505 2174.660 2725.795 2174.705 ;
        RECT 2724.430 2174.520 2725.795 2174.660 ;
        RECT 2725.505 2174.475 2725.795 2174.520 ;
        RECT 2501.090 2173.860 2501.410 2173.920 ;
        RECT 2677.270 2173.860 2677.590 2173.920 ;
        RECT 2501.090 2173.720 2677.590 2173.860 ;
        RECT 2501.090 2173.660 2501.410 2173.720 ;
        RECT 2677.270 2173.660 2677.590 2173.720 ;
        RECT 2694.670 2172.280 2694.990 2172.340 ;
        RECT 2696.985 2172.280 2697.275 2172.325 ;
        RECT 2694.670 2172.140 2697.275 2172.280 ;
        RECT 2694.670 2172.080 2694.990 2172.140 ;
        RECT 2696.985 2172.095 2697.275 2172.140 ;
        RECT 2697.430 2171.260 2697.750 2171.320 ;
        RECT 2697.905 2171.260 2698.195 2171.305 ;
        RECT 2697.430 2171.120 2698.195 2171.260 ;
        RECT 2697.430 2171.060 2697.750 2171.120 ;
        RECT 2697.905 2171.075 2698.195 2171.120 ;
        RECT 2507.990 2166.720 2508.310 2166.780 ;
        RECT 2677.270 2166.720 2677.590 2166.780 ;
        RECT 2507.990 2166.580 2677.590 2166.720 ;
        RECT 2697.890 2166.640 2698.210 2166.900 ;
        RECT 2698.350 2166.640 2698.670 2166.900 ;
        RECT 2507.990 2166.520 2508.310 2166.580 ;
        RECT 2677.270 2166.520 2677.590 2166.580 ;
        RECT 2697.430 2166.300 2697.750 2166.560 ;
        RECT 2697.980 2166.500 2698.120 2166.640 ;
        RECT 2702.030 2166.500 2702.350 2166.560 ;
        RECT 2697.980 2166.360 2702.350 2166.500 ;
        RECT 2702.030 2166.300 2702.350 2166.360 ;
        RECT 2699.285 2165.820 2699.575 2165.865 ;
        RECT 2702.950 2165.820 2703.270 2165.880 ;
        RECT 2699.285 2165.680 2703.270 2165.820 ;
        RECT 2699.285 2165.635 2699.575 2165.680 ;
        RECT 2702.950 2165.620 2703.270 2165.680 ;
        RECT 2694.670 2163.780 2694.990 2163.840 ;
        RECT 2696.985 2163.780 2697.275 2163.825 ;
        RECT 2694.670 2163.640 2697.275 2163.780 ;
        RECT 2694.670 2163.580 2694.990 2163.640 ;
        RECT 2696.985 2163.595 2697.275 2163.640 ;
        RECT 2359.565 2163.055 2359.855 2163.285 ;
        RECT 2359.625 2162.590 2359.795 2163.055 ;
        RECT 2362.975 2163.045 2363.265 2163.275 ;
        RECT 2374.660 2163.055 2374.950 2163.285 ;
        RECT 2363.035 2162.680 2363.205 2163.045 ;
        RECT 2359.535 2162.310 2359.875 2162.590 ;
        RECT 2362.940 2162.310 2363.310 2162.680 ;
        RECT 2374.720 2162.575 2374.890 2163.055 ;
        RECT 2376.450 2163.025 2376.745 2163.285 ;
        RECT 2377.440 2163.025 2377.735 2163.285 ;
        RECT 2380.195 2163.045 2380.485 2163.275 ;
        RECT 2391.880 2163.055 2392.170 2163.285 ;
        RECT 2376.080 2162.650 2376.310 2162.670 ;
        RECT 2376.050 2162.575 2376.340 2162.650 ;
        RECT 2374.720 2162.545 2376.340 2162.575 ;
        RECT 2374.660 2162.405 2376.340 2162.545 ;
        RECT 2374.660 2162.315 2374.950 2162.405 ;
        RECT 2376.050 2162.340 2376.340 2162.405 ;
        RECT 2376.080 2162.315 2376.310 2162.340 ;
        RECT 2362.975 2162.305 2363.265 2162.310 ;
        RECT 2375.115 2162.175 2375.440 2162.265 ;
        RECT 2363.405 2162.140 2363.695 2162.165 ;
        RECT 2375.090 2162.145 2375.440 2162.175 ;
        RECT 2363.385 2162.135 2363.725 2162.140 ;
        RECT 2363.235 2161.965 2363.725 2162.135 ;
        RECT 2374.920 2161.975 2375.440 2162.145 ;
        RECT 2363.385 2161.860 2363.725 2161.965 ;
        RECT 2375.090 2161.945 2375.440 2161.975 ;
        RECT 2375.115 2161.940 2375.440 2161.945 ;
        RECT 2376.510 2161.925 2376.680 2163.025 ;
        RECT 2377.500 2162.270 2377.670 2163.025 ;
        RECT 2380.255 2162.680 2380.425 2163.045 ;
        RECT 2380.160 2162.310 2380.530 2162.680 ;
        RECT 2391.940 2162.575 2392.110 2163.055 ;
        RECT 2393.670 2163.025 2393.965 2163.285 ;
        RECT 2394.660 2163.025 2394.955 2163.285 ;
        RECT 2397.415 2163.045 2397.705 2163.275 ;
        RECT 2409.100 2163.055 2409.390 2163.285 ;
        RECT 2393.300 2162.650 2393.530 2162.670 ;
        RECT 2393.270 2162.575 2393.560 2162.650 ;
        RECT 2391.940 2162.545 2393.560 2162.575 ;
        RECT 2391.880 2162.405 2393.560 2162.545 ;
        RECT 2391.880 2162.315 2392.170 2162.405 ;
        RECT 2393.270 2162.340 2393.560 2162.405 ;
        RECT 2393.300 2162.315 2393.530 2162.340 ;
        RECT 2380.195 2162.305 2380.485 2162.310 ;
        RECT 2377.500 2161.945 2377.830 2162.270 ;
        RECT 2392.335 2162.175 2392.660 2162.265 ;
        RECT 2380.625 2162.140 2380.915 2162.165 ;
        RECT 2392.310 2162.145 2392.660 2162.175 ;
        RECT 2380.605 2162.135 2380.945 2162.140 ;
        RECT 2380.455 2161.965 2380.945 2162.135 ;
        RECT 2392.140 2161.975 2392.660 2162.145 ;
        RECT 2377.500 2161.925 2377.790 2161.945 ;
        RECT 2376.450 2161.920 2376.680 2161.925 ;
        RECT 2359.160 2161.785 2359.500 2161.850 ;
        RECT 2374.315 2161.815 2374.635 2161.890 ;
        RECT 2374.290 2161.785 2374.635 2161.815 ;
        RECT 2359.020 2161.615 2359.500 2161.785 ;
        RECT 2374.115 2161.615 2374.635 2161.785 ;
        RECT 2376.450 2161.685 2376.740 2161.920 ;
        RECT 2377.440 2161.835 2377.790 2161.925 ;
        RECT 2380.605 2161.860 2380.945 2161.965 ;
        RECT 2392.310 2161.945 2392.660 2161.975 ;
        RECT 2392.335 2161.940 2392.660 2161.945 ;
        RECT 2393.730 2161.925 2393.900 2163.025 ;
        RECT 2394.720 2162.270 2394.890 2163.025 ;
        RECT 2397.475 2162.680 2397.645 2163.045 ;
        RECT 2397.380 2162.310 2397.750 2162.680 ;
        RECT 2409.160 2162.575 2409.330 2163.055 ;
        RECT 2410.890 2163.025 2411.185 2163.285 ;
        RECT 2411.880 2163.025 2412.175 2163.285 ;
        RECT 2414.635 2163.045 2414.925 2163.275 ;
        RECT 2426.320 2163.055 2426.610 2163.285 ;
        RECT 2410.520 2162.650 2410.750 2162.670 ;
        RECT 2410.490 2162.575 2410.780 2162.650 ;
        RECT 2409.160 2162.545 2410.780 2162.575 ;
        RECT 2409.100 2162.405 2410.780 2162.545 ;
        RECT 2409.100 2162.315 2409.390 2162.405 ;
        RECT 2410.490 2162.340 2410.780 2162.405 ;
        RECT 2410.520 2162.315 2410.750 2162.340 ;
        RECT 2397.415 2162.305 2397.705 2162.310 ;
        RECT 2394.720 2161.945 2395.050 2162.270 ;
        RECT 2409.555 2162.175 2409.880 2162.265 ;
        RECT 2397.845 2162.140 2398.135 2162.165 ;
        RECT 2409.530 2162.145 2409.880 2162.175 ;
        RECT 2397.825 2162.135 2398.165 2162.140 ;
        RECT 2397.675 2161.965 2398.165 2162.135 ;
        RECT 2409.360 2161.975 2409.880 2162.145 ;
        RECT 2394.720 2161.925 2395.010 2161.945 ;
        RECT 2393.670 2161.920 2393.900 2161.925 ;
        RECT 2377.440 2161.685 2377.730 2161.835 ;
        RECT 2391.535 2161.815 2391.855 2161.890 ;
        RECT 2391.510 2161.785 2391.855 2161.815 ;
        RECT 2391.335 2161.615 2391.855 2161.785 ;
        RECT 2393.670 2161.685 2393.960 2161.920 ;
        RECT 2394.660 2161.845 2395.010 2161.925 ;
        RECT 2397.825 2161.860 2398.165 2161.965 ;
        RECT 2409.530 2161.945 2409.880 2161.975 ;
        RECT 2409.555 2161.940 2409.880 2161.945 ;
        RECT 2410.950 2161.925 2411.120 2163.025 ;
        RECT 2411.940 2162.270 2412.110 2163.025 ;
        RECT 2414.695 2162.680 2414.865 2163.045 ;
        RECT 2414.600 2162.310 2414.970 2162.680 ;
        RECT 2426.380 2162.575 2426.550 2163.055 ;
        RECT 2428.110 2163.025 2428.405 2163.285 ;
        RECT 2429.100 2163.025 2429.395 2163.285 ;
        RECT 2431.855 2163.045 2432.145 2163.275 ;
        RECT 2443.540 2163.055 2443.830 2163.285 ;
        RECT 2427.740 2162.650 2427.970 2162.670 ;
        RECT 2427.710 2162.575 2428.000 2162.650 ;
        RECT 2426.380 2162.545 2428.000 2162.575 ;
        RECT 2426.320 2162.405 2428.000 2162.545 ;
        RECT 2426.320 2162.315 2426.610 2162.405 ;
        RECT 2427.710 2162.340 2428.000 2162.405 ;
        RECT 2427.740 2162.315 2427.970 2162.340 ;
        RECT 2414.635 2162.305 2414.925 2162.310 ;
        RECT 2411.940 2161.945 2412.270 2162.270 ;
        RECT 2426.775 2162.175 2427.100 2162.265 ;
        RECT 2415.065 2162.140 2415.355 2162.165 ;
        RECT 2426.750 2162.145 2427.100 2162.175 ;
        RECT 2415.045 2162.135 2415.385 2162.140 ;
        RECT 2414.895 2161.965 2415.385 2162.135 ;
        RECT 2426.580 2161.975 2427.100 2162.145 ;
        RECT 2411.940 2161.925 2412.230 2161.945 ;
        RECT 2410.890 2161.920 2411.120 2161.925 ;
        RECT 2394.660 2161.685 2394.950 2161.845 ;
        RECT 2408.755 2161.815 2409.075 2161.890 ;
        RECT 2408.730 2161.785 2409.075 2161.815 ;
        RECT 2408.555 2161.615 2409.075 2161.785 ;
        RECT 2410.890 2161.685 2411.180 2161.920 ;
        RECT 2411.880 2161.825 2412.230 2161.925 ;
        RECT 2415.045 2161.860 2415.385 2161.965 ;
        RECT 2426.750 2161.945 2427.100 2161.975 ;
        RECT 2426.775 2161.940 2427.100 2161.945 ;
        RECT 2428.170 2161.925 2428.340 2163.025 ;
        RECT 2429.160 2162.270 2429.330 2163.025 ;
        RECT 2431.915 2162.680 2432.085 2163.045 ;
        RECT 2431.820 2162.310 2432.190 2162.680 ;
        RECT 2443.600 2162.575 2443.770 2163.055 ;
        RECT 2445.330 2163.025 2445.625 2163.285 ;
        RECT 2446.320 2163.025 2446.615 2163.285 ;
        RECT 2444.960 2162.650 2445.190 2162.670 ;
        RECT 2444.930 2162.575 2445.220 2162.650 ;
        RECT 2443.600 2162.545 2445.220 2162.575 ;
        RECT 2443.540 2162.405 2445.220 2162.545 ;
        RECT 2443.540 2162.315 2443.830 2162.405 ;
        RECT 2444.930 2162.340 2445.220 2162.405 ;
        RECT 2444.960 2162.315 2445.190 2162.340 ;
        RECT 2431.855 2162.305 2432.145 2162.310 ;
        RECT 2429.160 2161.945 2429.490 2162.270 ;
        RECT 2443.995 2162.175 2444.320 2162.265 ;
        RECT 2432.285 2162.140 2432.575 2162.165 ;
        RECT 2443.970 2162.145 2444.320 2162.175 ;
        RECT 2432.265 2162.135 2432.605 2162.140 ;
        RECT 2432.115 2161.965 2432.605 2162.135 ;
        RECT 2443.800 2161.975 2444.320 2162.145 ;
        RECT 2429.160 2161.925 2429.450 2161.945 ;
        RECT 2428.110 2161.920 2428.340 2161.925 ;
        RECT 2411.880 2161.685 2412.170 2161.825 ;
        RECT 2425.975 2161.815 2426.295 2161.890 ;
        RECT 2425.950 2161.785 2426.295 2161.815 ;
        RECT 2425.775 2161.615 2426.295 2161.785 ;
        RECT 2428.110 2161.685 2428.400 2161.920 ;
        RECT 2429.100 2161.805 2429.450 2161.925 ;
        RECT 2432.265 2161.860 2432.605 2161.965 ;
        RECT 2443.970 2161.945 2444.320 2161.975 ;
        RECT 2443.995 2161.940 2444.320 2161.945 ;
        RECT 2445.390 2161.925 2445.560 2163.025 ;
        RECT 2446.350 2163.010 2446.615 2163.025 ;
        RECT 2446.350 2162.585 2446.675 2163.010 ;
        RECT 2697.890 2162.900 2698.210 2163.160 ;
        RECT 2446.380 2161.925 2446.550 2162.585 ;
        RECT 2445.330 2161.920 2445.560 2161.925 ;
        RECT 2446.320 2161.920 2446.550 2161.925 ;
        RECT 2697.890 2162.080 2698.210 2162.140 ;
        RECT 2698.825 2162.080 2699.115 2162.125 ;
        RECT 2697.890 2161.940 2699.115 2162.080 ;
        RECT 2443.195 2161.815 2443.515 2161.890 ;
        RECT 2429.100 2161.685 2429.390 2161.805 ;
        RECT 2443.170 2161.785 2443.515 2161.815 ;
        RECT 2442.995 2161.615 2443.515 2161.785 ;
        RECT 2445.330 2161.685 2445.620 2161.920 ;
        RECT 2446.320 2161.685 2446.610 2161.920 ;
        RECT 2697.890 2161.880 2698.210 2161.940 ;
        RECT 2698.825 2161.895 2699.115 2161.940 ;
        RECT 2700.665 2162.080 2700.955 2162.125 ;
        RECT 2701.585 2162.080 2701.875 2162.125 ;
        RECT 2700.665 2161.940 2701.875 2162.080 ;
        RECT 2700.665 2161.895 2700.955 2161.940 ;
        RECT 2701.585 2161.895 2701.875 2161.940 ;
        RECT 2702.030 2161.880 2702.350 2162.140 ;
        RECT 2702.950 2161.880 2703.270 2162.140 ;
        RECT 2703.410 2161.880 2703.730 2162.140 ;
        RECT 2698.350 2161.740 2698.670 2161.800 ;
        RECT 2359.160 2161.570 2359.500 2161.615 ;
        RECT 2374.290 2161.585 2374.635 2161.615 ;
        RECT 2391.510 2161.585 2391.855 2161.615 ;
        RECT 2408.730 2161.585 2409.075 2161.615 ;
        RECT 2425.950 2161.585 2426.295 2161.615 ;
        RECT 2443.170 2161.585 2443.515 2161.615 ;
        RECT 2374.315 2161.565 2374.635 2161.585 ;
        RECT 2391.535 2161.565 2391.855 2161.585 ;
        RECT 2408.755 2161.565 2409.075 2161.585 ;
        RECT 2425.975 2161.565 2426.295 2161.585 ;
        RECT 2443.195 2161.565 2443.515 2161.585 ;
        RECT 2697.980 2161.600 2698.670 2161.740 ;
        RECT 2697.980 2161.105 2698.120 2161.600 ;
        RECT 2698.350 2161.540 2698.670 2161.600 ;
        RECT 2702.120 2161.445 2702.260 2161.880 ;
        RECT 2702.045 2161.215 2702.335 2161.445 ;
        RECT 2702.490 2161.200 2702.810 2161.460 ;
        RECT 2703.040 2161.445 2703.180 2161.880 ;
        RECT 2702.965 2161.215 2703.255 2161.445 ;
        RECT 2366.675 2161.005 2366.965 2161.050 ;
        RECT 2367.680 2161.005 2368.000 2161.035 ;
        RECT 2369.040 2161.005 2369.360 2161.050 ;
        RECT 2366.675 2160.865 2368.590 2161.005 ;
        RECT 2366.675 2160.820 2366.965 2160.865 ;
        RECT 2367.675 2160.835 2368.005 2160.865 ;
        RECT 2367.680 2160.775 2368.000 2160.835 ;
        RECT 2368.450 2160.650 2368.590 2160.865 ;
        RECT 2369.040 2160.865 2369.635 2161.005 ;
        RECT 2369.040 2160.790 2369.360 2160.865 ;
        RECT 2370.415 2160.805 2371.060 2161.050 ;
        RECT 2383.895 2161.005 2384.185 2161.050 ;
        RECT 2384.900 2161.005 2385.220 2161.035 ;
        RECT 2386.260 2161.005 2386.580 2161.050 ;
        RECT 2383.895 2160.865 2385.810 2161.005 ;
        RECT 2383.895 2160.820 2384.185 2160.865 ;
        RECT 2384.895 2160.835 2385.225 2160.865 ;
        RECT 2370.740 2160.775 2371.060 2160.805 ;
        RECT 2384.900 2160.775 2385.220 2160.835 ;
        RECT 2385.670 2160.650 2385.810 2160.865 ;
        RECT 2386.260 2160.865 2386.855 2161.005 ;
        RECT 2386.260 2160.790 2386.580 2160.865 ;
        RECT 2387.635 2160.805 2388.280 2161.050 ;
        RECT 2401.115 2161.005 2401.405 2161.050 ;
        RECT 2402.120 2161.005 2402.440 2161.035 ;
        RECT 2403.480 2161.005 2403.800 2161.050 ;
        RECT 2401.115 2160.865 2403.030 2161.005 ;
        RECT 2401.115 2160.820 2401.405 2160.865 ;
        RECT 2402.115 2160.835 2402.445 2160.865 ;
        RECT 2387.960 2160.775 2388.280 2160.805 ;
        RECT 2402.120 2160.775 2402.440 2160.835 ;
        RECT 2402.890 2160.650 2403.030 2160.865 ;
        RECT 2403.480 2160.865 2404.075 2161.005 ;
        RECT 2403.480 2160.790 2403.800 2160.865 ;
        RECT 2404.855 2160.805 2405.500 2161.050 ;
        RECT 2418.335 2161.005 2418.625 2161.050 ;
        RECT 2419.340 2161.005 2419.660 2161.035 ;
        RECT 2420.700 2161.005 2421.020 2161.050 ;
        RECT 2418.335 2160.865 2420.250 2161.005 ;
        RECT 2418.335 2160.820 2418.625 2160.865 ;
        RECT 2419.335 2160.835 2419.665 2160.865 ;
        RECT 2405.180 2160.775 2405.500 2160.805 ;
        RECT 2419.340 2160.775 2419.660 2160.835 ;
        RECT 2420.110 2160.650 2420.250 2160.865 ;
        RECT 2420.700 2160.865 2421.295 2161.005 ;
        RECT 2420.700 2160.790 2421.020 2160.865 ;
        RECT 2422.075 2160.805 2422.720 2161.050 ;
        RECT 2435.555 2161.005 2435.845 2161.050 ;
        RECT 2436.560 2161.005 2436.880 2161.035 ;
        RECT 2437.920 2161.005 2438.240 2161.050 ;
        RECT 2435.555 2160.865 2437.470 2161.005 ;
        RECT 2435.555 2160.820 2435.845 2160.865 ;
        RECT 2436.555 2160.835 2436.885 2160.865 ;
        RECT 2422.400 2160.775 2422.720 2160.805 ;
        RECT 2436.560 2160.775 2436.880 2160.835 ;
        RECT 2437.330 2160.650 2437.470 2160.865 ;
        RECT 2437.920 2160.865 2438.515 2161.005 ;
        RECT 2437.920 2160.790 2438.240 2160.865 ;
        RECT 2439.295 2160.805 2439.940 2161.050 ;
        RECT 2697.905 2160.875 2698.195 2161.105 ;
        RECT 2698.350 2160.860 2698.670 2161.120 ;
        RECT 2702.580 2161.060 2702.720 2161.200 ;
        RECT 2703.425 2161.060 2703.715 2161.105 ;
        RECT 2702.580 2160.920 2703.715 2161.060 ;
        RECT 2703.425 2160.875 2703.715 2160.920 ;
        RECT 2439.620 2160.775 2439.940 2160.805 ;
        RECT 2368.450 2160.510 2370.460 2160.650 ;
        RECT 2385.670 2160.510 2387.680 2160.650 ;
        RECT 2402.890 2160.510 2404.900 2160.650 ;
        RECT 2420.110 2160.510 2422.120 2160.650 ;
        RECT 2437.330 2160.510 2439.340 2160.650 ;
        RECT 2370.320 2160.370 2370.460 2160.510 ;
        RECT 2387.540 2160.370 2387.680 2160.510 ;
        RECT 2404.760 2160.370 2404.900 2160.510 ;
        RECT 2421.980 2160.370 2422.120 2160.510 ;
        RECT 2439.200 2160.370 2439.340 2160.510 ;
        RECT 2368.365 2160.125 2369.010 2160.370 ;
        RECT 2368.690 2160.110 2369.010 2160.125 ;
        RECT 2369.720 2160.110 2370.040 2160.370 ;
        RECT 2370.245 2160.140 2370.535 2160.370 ;
        RECT 2371.095 2160.140 2371.385 2160.370 ;
        RECT 2369.810 2159.970 2369.950 2160.110 ;
        RECT 2371.170 2159.970 2371.310 2160.140 ;
        RECT 2385.585 2160.125 2386.230 2160.370 ;
        RECT 2385.910 2160.110 2386.230 2160.125 ;
        RECT 2386.940 2160.110 2387.260 2160.370 ;
        RECT 2387.465 2160.140 2387.755 2160.370 ;
        RECT 2388.315 2160.140 2388.605 2160.370 ;
        RECT 2369.810 2159.830 2371.310 2159.970 ;
        RECT 2387.030 2159.970 2387.170 2160.110 ;
        RECT 2388.390 2159.970 2388.530 2160.140 ;
        RECT 2402.805 2160.125 2403.450 2160.370 ;
        RECT 2403.130 2160.110 2403.450 2160.125 ;
        RECT 2404.160 2160.110 2404.480 2160.370 ;
        RECT 2404.685 2160.140 2404.975 2160.370 ;
        RECT 2405.535 2160.140 2405.825 2160.370 ;
        RECT 2387.030 2159.830 2388.530 2159.970 ;
        RECT 2404.250 2159.970 2404.390 2160.110 ;
        RECT 2405.610 2159.970 2405.750 2160.140 ;
        RECT 2420.025 2160.125 2420.670 2160.370 ;
        RECT 2420.350 2160.110 2420.670 2160.125 ;
        RECT 2421.380 2160.110 2421.700 2160.370 ;
        RECT 2421.905 2160.140 2422.195 2160.370 ;
        RECT 2422.755 2160.140 2423.045 2160.370 ;
        RECT 2404.250 2159.830 2405.750 2159.970 ;
        RECT 2421.470 2159.970 2421.610 2160.110 ;
        RECT 2422.830 2159.970 2422.970 2160.140 ;
        RECT 2437.245 2160.125 2437.890 2160.370 ;
        RECT 2437.570 2160.110 2437.890 2160.125 ;
        RECT 2438.600 2160.110 2438.920 2160.370 ;
        RECT 2439.125 2160.140 2439.415 2160.370 ;
        RECT 2439.975 2160.140 2440.265 2160.370 ;
        RECT 2702.490 2160.180 2702.810 2160.440 ;
        RECT 2421.470 2159.830 2422.970 2159.970 ;
        RECT 2438.690 2159.970 2438.830 2160.110 ;
        RECT 2440.050 2159.970 2440.190 2160.140 ;
        RECT 2438.690 2159.830 2440.190 2159.970 ;
        RECT 2514.890 2159.920 2515.210 2159.980 ;
        RECT 2677.270 2159.920 2677.590 2159.980 ;
        RECT 2514.890 2159.780 2677.590 2159.920 ;
        RECT 2514.890 2159.720 2515.210 2159.780 ;
        RECT 2677.270 2159.720 2677.590 2159.780 ;
        RECT 2365.640 2159.305 2365.960 2159.365 ;
        RECT 2365.365 2159.165 2365.960 2159.305 ;
        RECT 2365.640 2159.105 2365.960 2159.165 ;
        RECT 2367.915 2159.305 2368.205 2159.350 ;
        RECT 2370.060 2159.305 2370.380 2159.365 ;
        RECT 2382.860 2159.305 2383.180 2159.365 ;
        RECT 2367.915 2159.165 2370.380 2159.305 ;
        RECT 2382.585 2159.165 2383.180 2159.305 ;
        RECT 2367.915 2159.120 2368.205 2159.165 ;
        RECT 2370.060 2159.105 2370.380 2159.165 ;
        RECT 2382.860 2159.105 2383.180 2159.165 ;
        RECT 2385.135 2159.305 2385.425 2159.350 ;
        RECT 2387.280 2159.305 2387.600 2159.365 ;
        RECT 2400.080 2159.305 2400.400 2159.365 ;
        RECT 2385.135 2159.165 2387.600 2159.305 ;
        RECT 2399.805 2159.165 2400.400 2159.305 ;
        RECT 2385.135 2159.120 2385.425 2159.165 ;
        RECT 2387.280 2159.105 2387.600 2159.165 ;
        RECT 2400.080 2159.105 2400.400 2159.165 ;
        RECT 2402.355 2159.305 2402.645 2159.350 ;
        RECT 2404.500 2159.305 2404.820 2159.365 ;
        RECT 2417.300 2159.305 2417.620 2159.365 ;
        RECT 2402.355 2159.165 2404.820 2159.305 ;
        RECT 2417.025 2159.165 2417.620 2159.305 ;
        RECT 2402.355 2159.120 2402.645 2159.165 ;
        RECT 2404.500 2159.105 2404.820 2159.165 ;
        RECT 2417.300 2159.105 2417.620 2159.165 ;
        RECT 2419.575 2159.305 2419.865 2159.350 ;
        RECT 2421.720 2159.305 2422.040 2159.365 ;
        RECT 2434.520 2159.305 2434.840 2159.365 ;
        RECT 2419.575 2159.165 2422.040 2159.305 ;
        RECT 2434.245 2159.165 2434.840 2159.305 ;
        RECT 2419.575 2159.120 2419.865 2159.165 ;
        RECT 2421.720 2159.105 2422.040 2159.165 ;
        RECT 2434.520 2159.105 2434.840 2159.165 ;
        RECT 2436.795 2159.305 2437.085 2159.350 ;
        RECT 2438.940 2159.305 2439.260 2159.365 ;
        RECT 2436.795 2159.165 2439.260 2159.305 ;
        RECT 2436.795 2159.120 2437.085 2159.165 ;
        RECT 2438.940 2159.105 2439.260 2159.165 ;
        RECT 2698.810 2159.160 2699.130 2159.420 ;
        RECT 2699.745 2159.360 2700.035 2159.405 ;
        RECT 2702.490 2159.360 2702.810 2159.420 ;
        RECT 2699.745 2159.220 2702.810 2159.360 ;
        RECT 2699.745 2159.175 2700.035 2159.220 ;
        RECT 2702.490 2159.160 2702.810 2159.220 ;
        RECT 2696.985 2159.020 2697.275 2159.065 ;
        RECT 2697.430 2159.020 2697.750 2159.080 ;
        RECT 2696.985 2158.880 2697.750 2159.020 ;
        RECT 2698.900 2159.020 2699.040 2159.160 ;
        RECT 2702.030 2159.020 2702.350 2159.080 ;
        RECT 2698.900 2158.880 2702.350 2159.020 ;
        RECT 2696.985 2158.835 2697.275 2158.880 ;
        RECT 2697.430 2158.820 2697.750 2158.880 ;
        RECT 2702.030 2158.820 2702.350 2158.880 ;
        RECT 2367.015 2158.285 2367.305 2158.330 ;
        RECT 2369.380 2158.285 2369.700 2158.345 ;
        RECT 2367.015 2158.145 2369.700 2158.285 ;
        RECT 2367.015 2158.100 2367.305 2158.145 ;
        RECT 2369.380 2158.085 2369.700 2158.145 ;
        RECT 2370.060 2158.285 2370.380 2158.345 ;
        RECT 2371.095 2158.285 2371.385 2158.330 ;
        RECT 2370.060 2158.145 2371.385 2158.285 ;
        RECT 2370.060 2158.085 2370.380 2158.145 ;
        RECT 2371.095 2158.100 2371.385 2158.145 ;
        RECT 2384.235 2158.285 2384.525 2158.330 ;
        RECT 2386.600 2158.285 2386.920 2158.345 ;
        RECT 2384.235 2158.145 2386.920 2158.285 ;
        RECT 2384.235 2158.100 2384.525 2158.145 ;
        RECT 2386.600 2158.085 2386.920 2158.145 ;
        RECT 2387.280 2158.285 2387.600 2158.345 ;
        RECT 2388.315 2158.285 2388.605 2158.330 ;
        RECT 2387.280 2158.145 2388.605 2158.285 ;
        RECT 2387.280 2158.085 2387.600 2158.145 ;
        RECT 2388.315 2158.100 2388.605 2158.145 ;
        RECT 2401.455 2158.285 2401.745 2158.330 ;
        RECT 2403.820 2158.285 2404.140 2158.345 ;
        RECT 2401.455 2158.145 2404.140 2158.285 ;
        RECT 2401.455 2158.100 2401.745 2158.145 ;
        RECT 2403.820 2158.085 2404.140 2158.145 ;
        RECT 2404.500 2158.285 2404.820 2158.345 ;
        RECT 2405.535 2158.285 2405.825 2158.330 ;
        RECT 2404.500 2158.145 2405.825 2158.285 ;
        RECT 2404.500 2158.085 2404.820 2158.145 ;
        RECT 2405.535 2158.100 2405.825 2158.145 ;
        RECT 2418.675 2158.285 2418.965 2158.330 ;
        RECT 2421.040 2158.285 2421.360 2158.345 ;
        RECT 2418.675 2158.145 2421.360 2158.285 ;
        RECT 2418.675 2158.100 2418.965 2158.145 ;
        RECT 2421.040 2158.085 2421.360 2158.145 ;
        RECT 2421.720 2158.285 2422.040 2158.345 ;
        RECT 2422.755 2158.285 2423.045 2158.330 ;
        RECT 2421.720 2158.145 2423.045 2158.285 ;
        RECT 2421.720 2158.085 2422.040 2158.145 ;
        RECT 2422.755 2158.100 2423.045 2158.145 ;
        RECT 2435.895 2158.285 2436.185 2158.330 ;
        RECT 2438.260 2158.285 2438.580 2158.345 ;
        RECT 2435.895 2158.145 2438.580 2158.285 ;
        RECT 2435.895 2158.100 2436.185 2158.145 ;
        RECT 2438.260 2158.085 2438.580 2158.145 ;
        RECT 2438.940 2158.285 2439.260 2158.345 ;
        RECT 2439.975 2158.285 2440.265 2158.330 ;
        RECT 2438.940 2158.145 2440.265 2158.285 ;
        RECT 2438.940 2158.085 2439.260 2158.145 ;
        RECT 2439.975 2158.100 2440.265 2158.145 ;
        RECT 2365.145 2157.945 2365.435 2157.990 ;
        RECT 2368.020 2157.945 2368.340 2158.005 ;
        RECT 2365.145 2157.805 2368.340 2157.945 ;
        RECT 2365.145 2157.760 2365.435 2157.805 ;
        RECT 2365.640 2157.265 2365.960 2157.325 ;
        RECT 2367.600 2157.315 2367.740 2157.805 ;
        RECT 2368.020 2157.745 2368.340 2157.805 ;
        RECT 2382.365 2157.945 2382.655 2157.990 ;
        RECT 2385.240 2157.945 2385.560 2158.005 ;
        RECT 2382.365 2157.805 2385.560 2157.945 ;
        RECT 2382.365 2157.760 2382.655 2157.805 ;
        RECT 2369.040 2157.605 2369.360 2157.665 ;
        RECT 2368.765 2157.465 2369.360 2157.605 ;
        RECT 2369.040 2157.405 2369.360 2157.465 ;
        RECT 2367.015 2157.270 2367.305 2157.315 ;
        RECT 2365.365 2157.125 2365.960 2157.265 ;
        RECT 2365.640 2157.065 2365.960 2157.125 ;
        RECT 2366.410 2157.130 2367.305 2157.270 ;
        RECT 2366.410 2156.985 2366.550 2157.130 ;
        RECT 2367.015 2157.085 2367.305 2157.130 ;
        RECT 2367.525 2157.085 2367.815 2157.315 ;
        RECT 2368.360 2157.265 2368.680 2157.325 ;
        RECT 2370.740 2157.265 2371.060 2157.325 ;
        RECT 2382.860 2157.265 2383.180 2157.325 ;
        RECT 2384.820 2157.315 2384.960 2157.805 ;
        RECT 2385.240 2157.745 2385.560 2157.805 ;
        RECT 2399.585 2157.945 2399.875 2157.990 ;
        RECT 2402.460 2157.945 2402.780 2158.005 ;
        RECT 2399.585 2157.805 2402.780 2157.945 ;
        RECT 2399.585 2157.760 2399.875 2157.805 ;
        RECT 2386.260 2157.605 2386.580 2157.665 ;
        RECT 2385.985 2157.465 2386.580 2157.605 ;
        RECT 2386.260 2157.405 2386.580 2157.465 ;
        RECT 2384.235 2157.270 2384.525 2157.315 ;
        RECT 2368.085 2157.125 2368.680 2157.265 ;
        RECT 2370.465 2157.125 2371.060 2157.265 ;
        RECT 2382.585 2157.125 2383.180 2157.265 ;
        RECT 2368.360 2157.065 2368.680 2157.125 ;
        RECT 2370.740 2157.065 2371.060 2157.125 ;
        RECT 2382.860 2157.065 2383.180 2157.125 ;
        RECT 2383.630 2157.130 2384.525 2157.270 ;
        RECT 2383.630 2156.985 2383.770 2157.130 ;
        RECT 2384.235 2157.085 2384.525 2157.130 ;
        RECT 2384.745 2157.085 2385.035 2157.315 ;
        RECT 2385.580 2157.265 2385.900 2157.325 ;
        RECT 2387.960 2157.265 2388.280 2157.325 ;
        RECT 2400.080 2157.265 2400.400 2157.325 ;
        RECT 2402.040 2157.315 2402.180 2157.805 ;
        RECT 2402.460 2157.745 2402.780 2157.805 ;
        RECT 2416.805 2157.945 2417.095 2157.990 ;
        RECT 2419.680 2157.945 2420.000 2158.005 ;
        RECT 2416.805 2157.805 2420.000 2157.945 ;
        RECT 2416.805 2157.760 2417.095 2157.805 ;
        RECT 2403.480 2157.605 2403.800 2157.665 ;
        RECT 2403.205 2157.465 2403.800 2157.605 ;
        RECT 2403.480 2157.405 2403.800 2157.465 ;
        RECT 2401.455 2157.270 2401.745 2157.315 ;
        RECT 2385.305 2157.125 2385.900 2157.265 ;
        RECT 2387.685 2157.125 2388.280 2157.265 ;
        RECT 2394.830 2157.245 2395.150 2157.260 ;
        RECT 2385.580 2157.065 2385.900 2157.125 ;
        RECT 2387.960 2157.065 2388.280 2157.125 ;
        RECT 2394.655 2157.015 2395.150 2157.245 ;
        RECT 2399.805 2157.125 2400.400 2157.265 ;
        RECT 2400.080 2157.065 2400.400 2157.125 ;
        RECT 2400.850 2157.130 2401.745 2157.270 ;
        RECT 2394.830 2157.000 2395.150 2157.015 ;
        RECT 2400.850 2156.985 2400.990 2157.130 ;
        RECT 2401.455 2157.085 2401.745 2157.130 ;
        RECT 2401.965 2157.085 2402.255 2157.315 ;
        RECT 2402.800 2157.265 2403.120 2157.325 ;
        RECT 2405.180 2157.265 2405.500 2157.325 ;
        RECT 2417.300 2157.265 2417.620 2157.325 ;
        RECT 2419.260 2157.315 2419.400 2157.805 ;
        RECT 2419.680 2157.745 2420.000 2157.805 ;
        RECT 2434.025 2157.945 2434.315 2157.990 ;
        RECT 2436.900 2157.945 2437.220 2158.005 ;
        RECT 2434.025 2157.805 2437.220 2157.945 ;
        RECT 2434.025 2157.760 2434.315 2157.805 ;
        RECT 2420.700 2157.605 2421.020 2157.665 ;
        RECT 2420.425 2157.465 2421.020 2157.605 ;
        RECT 2420.700 2157.405 2421.020 2157.465 ;
        RECT 2418.675 2157.270 2418.965 2157.315 ;
        RECT 2402.525 2157.125 2403.120 2157.265 ;
        RECT 2404.905 2157.125 2405.500 2157.265 ;
        RECT 2417.025 2157.125 2417.620 2157.265 ;
        RECT 2402.800 2157.065 2403.120 2157.125 ;
        RECT 2405.180 2157.065 2405.500 2157.125 ;
        RECT 2417.300 2157.065 2417.620 2157.125 ;
        RECT 2418.070 2157.130 2418.965 2157.270 ;
        RECT 2418.070 2156.985 2418.210 2157.130 ;
        RECT 2418.675 2157.085 2418.965 2157.130 ;
        RECT 2419.185 2157.085 2419.475 2157.315 ;
        RECT 2420.020 2157.265 2420.340 2157.325 ;
        RECT 2422.400 2157.265 2422.720 2157.325 ;
        RECT 2434.520 2157.265 2434.840 2157.325 ;
        RECT 2436.480 2157.315 2436.620 2157.805 ;
        RECT 2436.900 2157.745 2437.220 2157.805 ;
        RECT 2437.920 2157.605 2438.240 2157.665 ;
        RECT 2437.645 2157.465 2438.240 2157.605 ;
        RECT 2437.920 2157.405 2438.240 2157.465 ;
        RECT 2698.810 2157.460 2699.130 2157.720 ;
        RECT 2435.895 2157.270 2436.185 2157.315 ;
        RECT 2419.745 2157.125 2420.340 2157.265 ;
        RECT 2422.125 2157.125 2422.720 2157.265 ;
        RECT 2420.020 2157.065 2420.340 2157.125 ;
        RECT 2422.400 2157.065 2422.720 2157.125 ;
        RECT 2428.870 2157.245 2429.190 2157.260 ;
        RECT 2428.870 2157.015 2429.385 2157.245 ;
        RECT 2434.245 2157.125 2434.840 2157.265 ;
        RECT 2434.520 2157.065 2434.840 2157.125 ;
        RECT 2435.290 2157.130 2436.185 2157.270 ;
        RECT 2428.870 2157.000 2429.190 2157.015 ;
        RECT 2435.290 2156.985 2435.430 2157.130 ;
        RECT 2435.895 2157.085 2436.185 2157.130 ;
        RECT 2436.405 2157.085 2436.695 2157.315 ;
        RECT 2437.240 2157.265 2437.560 2157.325 ;
        RECT 2439.620 2157.265 2439.940 2157.325 ;
        RECT 2436.965 2157.125 2437.560 2157.265 ;
        RECT 2439.345 2157.125 2439.940 2157.265 ;
        RECT 2437.240 2157.065 2437.560 2157.125 ;
        RECT 2439.620 2157.065 2439.940 2157.125 ;
        RECT 2366.320 2156.725 2366.640 2156.985 ;
        RECT 2374.315 2156.875 2374.635 2156.980 ;
        RECT 2374.290 2156.860 2374.635 2156.875 ;
        RECT 2367.680 2156.800 2368.000 2156.815 ;
        RECT 2367.680 2156.755 2368.185 2156.800 ;
        RECT 2367.590 2156.615 2368.185 2156.755 ;
        RECT 2374.000 2156.690 2374.635 2156.860 ;
        RECT 2374.115 2156.675 2374.635 2156.690 ;
        RECT 2374.290 2156.660 2374.635 2156.675 ;
        RECT 2374.290 2156.645 2374.580 2156.660 ;
        RECT 2367.680 2156.570 2368.185 2156.615 ;
        RECT 2367.680 2156.555 2368.000 2156.570 ;
        RECT 2372.645 2156.290 2372.970 2156.615 ;
        RECT 2375.090 2156.485 2375.440 2156.610 ;
        RECT 2376.450 2156.540 2376.740 2156.775 ;
        RECT 2377.435 2156.540 2377.725 2156.775 ;
        RECT 2383.540 2156.725 2383.860 2156.985 ;
        RECT 2391.535 2156.875 2391.855 2156.980 ;
        RECT 2391.510 2156.860 2391.855 2156.875 ;
        RECT 2384.900 2156.800 2385.220 2156.815 ;
        RECT 2384.900 2156.755 2385.405 2156.800 ;
        RECT 2384.810 2156.615 2385.405 2156.755 ;
        RECT 2391.220 2156.690 2391.855 2156.860 ;
        RECT 2391.335 2156.675 2391.855 2156.690 ;
        RECT 2391.510 2156.660 2391.855 2156.675 ;
        RECT 2391.510 2156.645 2391.800 2156.660 ;
        RECT 2384.900 2156.570 2385.405 2156.615 ;
        RECT 2384.900 2156.555 2385.220 2156.570 ;
        RECT 2376.450 2156.535 2376.680 2156.540 ;
        RECT 2377.435 2156.535 2377.665 2156.540 ;
        RECT 2374.920 2156.315 2375.440 2156.485 ;
        RECT 2375.090 2156.260 2375.440 2156.315 ;
        RECT 2376.090 2156.225 2376.325 2156.235 ;
        RECT 2374.660 2156.120 2374.950 2156.145 ;
        RECT 2376.030 2156.120 2376.370 2156.225 ;
        RECT 2374.660 2155.950 2376.370 2156.120 ;
        RECT 2374.660 2155.915 2374.950 2155.950 ;
        RECT 2374.720 2155.405 2374.890 2155.915 ;
        RECT 2376.030 2155.910 2376.370 2155.950 ;
        RECT 2376.090 2155.885 2376.325 2155.910 ;
        RECT 2376.510 2155.435 2376.680 2156.535 ;
        RECT 2377.495 2155.435 2377.665 2156.535 ;
        RECT 2389.865 2156.290 2390.190 2156.615 ;
        RECT 2392.310 2156.485 2392.660 2156.610 ;
        RECT 2393.670 2156.540 2393.960 2156.775 ;
        RECT 2394.655 2156.540 2394.945 2156.775 ;
        RECT 2400.760 2156.725 2401.080 2156.985 ;
        RECT 2408.755 2156.875 2409.075 2156.980 ;
        RECT 2408.730 2156.860 2409.075 2156.875 ;
        RECT 2402.120 2156.800 2402.440 2156.815 ;
        RECT 2402.120 2156.755 2402.625 2156.800 ;
        RECT 2402.030 2156.615 2402.625 2156.755 ;
        RECT 2408.440 2156.690 2409.075 2156.860 ;
        RECT 2408.555 2156.675 2409.075 2156.690 ;
        RECT 2408.730 2156.660 2409.075 2156.675 ;
        RECT 2408.730 2156.645 2409.020 2156.660 ;
        RECT 2402.120 2156.570 2402.625 2156.615 ;
        RECT 2402.120 2156.555 2402.440 2156.570 ;
        RECT 2393.670 2156.535 2393.900 2156.540 ;
        RECT 2394.655 2156.535 2394.885 2156.540 ;
        RECT 2392.140 2156.315 2392.660 2156.485 ;
        RECT 2392.310 2156.260 2392.660 2156.315 ;
        RECT 2393.310 2156.225 2393.545 2156.235 ;
        RECT 2391.880 2156.120 2392.170 2156.145 ;
        RECT 2393.250 2156.120 2393.590 2156.225 ;
        RECT 2391.880 2155.950 2393.590 2156.120 ;
        RECT 2391.880 2155.915 2392.170 2155.950 ;
        RECT 2374.660 2155.175 2374.950 2155.405 ;
        RECT 2376.450 2155.175 2376.745 2155.435 ;
        RECT 2377.350 2155.175 2377.730 2155.435 ;
        RECT 2391.940 2155.405 2392.110 2155.915 ;
        RECT 2393.250 2155.910 2393.590 2155.950 ;
        RECT 2393.310 2155.885 2393.545 2155.910 ;
        RECT 2393.730 2155.435 2393.900 2156.535 ;
        RECT 2394.715 2155.435 2394.885 2156.535 ;
        RECT 2407.085 2156.290 2407.410 2156.615 ;
        RECT 2409.530 2156.485 2409.880 2156.610 ;
        RECT 2410.890 2156.540 2411.180 2156.775 ;
        RECT 2411.875 2156.540 2412.165 2156.775 ;
        RECT 2417.980 2156.725 2418.300 2156.985 ;
        RECT 2425.975 2156.875 2426.295 2156.980 ;
        RECT 2425.950 2156.860 2426.295 2156.875 ;
        RECT 2419.340 2156.800 2419.660 2156.815 ;
        RECT 2419.340 2156.755 2419.845 2156.800 ;
        RECT 2419.250 2156.615 2419.845 2156.755 ;
        RECT 2425.660 2156.690 2426.295 2156.860 ;
        RECT 2425.775 2156.675 2426.295 2156.690 ;
        RECT 2425.950 2156.660 2426.295 2156.675 ;
        RECT 2425.950 2156.645 2426.240 2156.660 ;
        RECT 2419.340 2156.570 2419.845 2156.615 ;
        RECT 2419.340 2156.555 2419.660 2156.570 ;
        RECT 2410.890 2156.535 2411.120 2156.540 ;
        RECT 2411.875 2156.535 2412.105 2156.540 ;
        RECT 2409.360 2156.315 2409.880 2156.485 ;
        RECT 2409.530 2156.260 2409.880 2156.315 ;
        RECT 2410.530 2156.225 2410.765 2156.235 ;
        RECT 2409.100 2156.120 2409.390 2156.145 ;
        RECT 2410.470 2156.120 2410.810 2156.225 ;
        RECT 2409.100 2155.950 2410.810 2156.120 ;
        RECT 2409.100 2155.915 2409.390 2155.950 ;
        RECT 2391.880 2155.175 2392.170 2155.405 ;
        RECT 2393.670 2155.175 2393.965 2155.435 ;
        RECT 2394.655 2155.175 2394.950 2155.435 ;
        RECT 2409.160 2155.405 2409.330 2155.915 ;
        RECT 2410.470 2155.910 2410.810 2155.950 ;
        RECT 2410.530 2155.885 2410.765 2155.910 ;
        RECT 2410.950 2155.435 2411.120 2156.535 ;
        RECT 2411.935 2155.435 2412.105 2156.535 ;
        RECT 2424.305 2156.290 2424.630 2156.615 ;
        RECT 2426.750 2156.485 2427.100 2156.610 ;
        RECT 2428.110 2156.540 2428.400 2156.775 ;
        RECT 2429.095 2156.540 2429.385 2156.775 ;
        RECT 2435.200 2156.725 2435.520 2156.985 ;
        RECT 2443.195 2156.875 2443.515 2156.980 ;
        RECT 2443.170 2156.860 2443.515 2156.875 ;
        RECT 2436.560 2156.800 2436.880 2156.815 ;
        RECT 2436.560 2156.755 2437.065 2156.800 ;
        RECT 2436.470 2156.615 2437.065 2156.755 ;
        RECT 2442.880 2156.690 2443.515 2156.860 ;
        RECT 2442.995 2156.675 2443.515 2156.690 ;
        RECT 2443.170 2156.660 2443.515 2156.675 ;
        RECT 2443.170 2156.645 2443.460 2156.660 ;
        RECT 2436.560 2156.570 2437.065 2156.615 ;
        RECT 2436.560 2156.555 2436.880 2156.570 ;
        RECT 2428.110 2156.535 2428.340 2156.540 ;
        RECT 2429.095 2156.535 2429.325 2156.540 ;
        RECT 2426.580 2156.315 2427.100 2156.485 ;
        RECT 2426.750 2156.260 2427.100 2156.315 ;
        RECT 2427.750 2156.225 2427.985 2156.235 ;
        RECT 2426.320 2156.120 2426.610 2156.145 ;
        RECT 2427.690 2156.120 2428.030 2156.225 ;
        RECT 2426.320 2155.950 2428.030 2156.120 ;
        RECT 2426.320 2155.915 2426.610 2155.950 ;
        RECT 2409.100 2155.175 2409.390 2155.405 ;
        RECT 2410.890 2155.175 2411.185 2155.435 ;
        RECT 2411.850 2155.175 2412.170 2155.435 ;
        RECT 2426.380 2155.405 2426.550 2155.915 ;
        RECT 2427.690 2155.910 2428.030 2155.950 ;
        RECT 2427.750 2155.885 2427.985 2155.910 ;
        RECT 2428.170 2155.435 2428.340 2156.535 ;
        RECT 2429.155 2155.435 2429.325 2156.535 ;
        RECT 2441.525 2156.290 2441.850 2156.615 ;
        RECT 2443.970 2156.485 2444.320 2156.610 ;
        RECT 2445.330 2156.540 2445.620 2156.775 ;
        RECT 2446.315 2156.540 2446.605 2156.775 ;
        RECT 2697.905 2156.640 2698.195 2156.685 ;
        RECT 2698.810 2156.640 2699.130 2156.700 ;
        RECT 2445.330 2156.535 2445.560 2156.540 ;
        RECT 2446.315 2156.535 2446.545 2156.540 ;
        RECT 2443.800 2156.315 2444.320 2156.485 ;
        RECT 2443.970 2156.260 2444.320 2156.315 ;
        RECT 2444.970 2156.225 2445.205 2156.235 ;
        RECT 2443.540 2156.120 2443.830 2156.145 ;
        RECT 2444.910 2156.120 2445.250 2156.225 ;
        RECT 2443.540 2155.950 2445.250 2156.120 ;
        RECT 2443.540 2155.915 2443.830 2155.950 ;
        RECT 2426.320 2155.175 2426.610 2155.405 ;
        RECT 2428.110 2155.175 2428.405 2155.435 ;
        RECT 2429.095 2155.175 2429.390 2155.435 ;
        RECT 2443.600 2155.405 2443.770 2155.915 ;
        RECT 2444.910 2155.910 2445.250 2155.950 ;
        RECT 2444.970 2155.885 2445.205 2155.910 ;
        RECT 2445.390 2155.435 2445.560 2156.535 ;
        RECT 2446.375 2155.435 2446.545 2156.535 ;
        RECT 2697.905 2156.500 2699.130 2156.640 ;
        RECT 2697.905 2156.455 2698.195 2156.500 ;
        RECT 2698.810 2156.440 2699.130 2156.500 ;
        RECT 2694.670 2155.960 2694.990 2156.020 ;
        RECT 2696.985 2155.960 2697.275 2156.005 ;
        RECT 2694.670 2155.820 2697.275 2155.960 ;
        RECT 2694.670 2155.760 2694.990 2155.820 ;
        RECT 2696.985 2155.775 2697.275 2155.820 ;
        RECT 2443.540 2155.175 2443.830 2155.405 ;
        RECT 2445.330 2155.175 2445.625 2155.435 ;
        RECT 2446.315 2155.375 2446.610 2155.435 ;
        RECT 2446.315 2155.235 2447.960 2155.375 ;
        RECT 2446.315 2155.175 2446.610 2155.235 ;
        RECT 2447.820 2155.160 2447.960 2155.235 ;
        RECT 2460.150 2155.160 2460.470 2155.220 ;
        RECT 2447.820 2155.020 2460.470 2155.160 ;
        RECT 2460.150 2154.960 2460.470 2155.020 ;
        RECT 2700.205 2153.240 2700.495 2153.285 ;
        RECT 2701.570 2153.240 2701.890 2153.300 ;
        RECT 2700.205 2153.100 2701.890 2153.240 ;
        RECT 2700.205 2153.055 2700.495 2153.100 ;
        RECT 2701.570 2153.040 2701.890 2153.100 ;
        RECT 2698.365 2152.900 2698.655 2152.945 ;
        RECT 2699.730 2152.900 2700.050 2152.960 ;
        RECT 2698.365 2152.760 2700.050 2152.900 ;
        RECT 2698.365 2152.715 2698.655 2152.760 ;
        RECT 2699.730 2152.700 2700.050 2152.760 ;
        RECT 2700.665 2152.900 2700.955 2152.945 ;
        RECT 2703.410 2152.900 2703.730 2152.960 ;
        RECT 2700.665 2152.760 2703.730 2152.900 ;
        RECT 2700.665 2152.715 2700.955 2152.760 ;
        RECT 2703.410 2152.700 2703.730 2152.760 ;
        RECT 2696.970 2152.560 2697.290 2152.620 ;
        RECT 2702.030 2152.560 2702.350 2152.620 ;
        RECT 2696.970 2152.420 2702.350 2152.560 ;
        RECT 2696.970 2152.360 2697.290 2152.420 ;
        RECT 2702.030 2152.360 2702.350 2152.420 ;
        RECT 2698.810 2152.020 2699.130 2152.280 ;
        RECT 2699.270 2152.020 2699.590 2152.280 ;
        RECT 2701.585 2152.220 2701.875 2152.265 ;
        RECT 2703.870 2152.220 2704.190 2152.280 ;
        RECT 2701.585 2152.080 2704.190 2152.220 ;
        RECT 2701.585 2152.035 2701.875 2152.080 ;
        RECT 2703.870 2152.020 2704.190 2152.080 ;
        RECT 2698.810 2151.200 2699.130 2151.260 ;
        RECT 2701.125 2151.200 2701.415 2151.245 ;
        RECT 2698.810 2151.060 2701.415 2151.200 ;
        RECT 2698.810 2151.000 2699.130 2151.060 ;
        RECT 2701.125 2151.015 2701.415 2151.060 ;
        RECT 2699.730 2150.860 2700.050 2150.920 ;
        RECT 2697.520 2150.720 2699.500 2150.860 ;
        RECT 2697.520 2150.580 2697.660 2150.720 ;
        RECT 2697.430 2150.320 2697.750 2150.580 ;
        RECT 2697.890 2150.320 2698.210 2150.580 ;
        RECT 2699.360 2150.225 2699.500 2150.720 ;
        RECT 2699.730 2150.720 2700.880 2150.860 ;
        RECT 2699.730 2150.660 2700.050 2150.720 ;
        RECT 2699.285 2149.995 2699.575 2150.225 ;
        RECT 2696.970 2149.500 2697.290 2149.560 ;
        RECT 2698.365 2149.500 2698.655 2149.545 ;
        RECT 2696.970 2149.360 2698.655 2149.500 ;
        RECT 2699.360 2149.500 2699.500 2149.995 ;
        RECT 2700.740 2149.885 2700.880 2150.720 ;
        RECT 2702.030 2150.320 2702.350 2150.580 ;
        RECT 2702.490 2150.320 2702.810 2150.580 ;
        RECT 2702.965 2150.335 2703.255 2150.565 ;
        RECT 2703.040 2150.180 2703.180 2150.335 ;
        RECT 2702.580 2150.040 2703.180 2150.180 ;
        RECT 2700.665 2149.655 2700.955 2149.885 ;
        RECT 2702.580 2149.500 2702.720 2150.040 ;
        RECT 2699.360 2149.360 2702.720 2149.500 ;
        RECT 2696.970 2149.300 2697.290 2149.360 ;
        RECT 2698.365 2149.315 2698.655 2149.360 ;
        RECT 2697.905 2148.480 2698.195 2148.525 ;
        RECT 2698.350 2148.480 2698.670 2148.540 ;
        RECT 2697.905 2148.340 2698.670 2148.480 ;
        RECT 2697.905 2148.295 2698.195 2148.340 ;
        RECT 2698.350 2148.280 2698.670 2148.340 ;
        RECT 2698.810 2148.480 2699.130 2148.540 ;
        RECT 2699.285 2148.480 2699.575 2148.525 ;
        RECT 2698.810 2148.340 2699.575 2148.480 ;
        RECT 2698.810 2148.280 2699.130 2148.340 ;
        RECT 2699.285 2148.295 2699.575 2148.340 ;
        RECT 2694.670 2147.460 2694.990 2147.520 ;
        RECT 2696.985 2147.460 2697.275 2147.505 ;
        RECT 2694.670 2147.320 2697.275 2147.460 ;
        RECT 2694.670 2147.260 2694.990 2147.320 ;
        RECT 2696.985 2147.275 2697.275 2147.320 ;
        RECT 2697.430 2147.460 2697.750 2147.520 ;
        RECT 2698.825 2147.460 2699.115 2147.505 ;
        RECT 2697.430 2147.320 2699.115 2147.460 ;
        RECT 2697.430 2147.260 2697.750 2147.320 ;
        RECT 2698.825 2147.275 2699.115 2147.320 ;
        RECT 2699.730 2147.260 2700.050 2147.520 ;
        RECT 2699.730 2145.760 2700.050 2145.820 ;
        RECT 2700.665 2145.760 2700.955 2145.805 ;
        RECT 2377.350 2145.640 2377.670 2145.700 ;
        RECT 2452.790 2145.640 2453.110 2145.700 ;
        RECT 2377.350 2145.500 2453.110 2145.640 ;
        RECT 2699.730 2145.620 2700.955 2145.760 ;
        RECT 2699.730 2145.560 2700.050 2145.620 ;
        RECT 2700.665 2145.575 2700.955 2145.620 ;
        RECT 2377.350 2145.440 2377.670 2145.500 ;
        RECT 2452.790 2145.440 2453.110 2145.500 ;
        RECT 2698.810 2144.880 2699.130 2145.140 ;
        RECT 2696.970 2144.740 2697.290 2144.800 ;
        RECT 2697.445 2144.740 2697.735 2144.785 ;
        RECT 2696.970 2144.600 2697.735 2144.740 ;
        RECT 2696.970 2144.540 2697.290 2144.600 ;
        RECT 2697.445 2144.555 2697.735 2144.600 ;
        RECT 2698.350 2144.540 2698.670 2144.800 ;
        RECT 2697.890 2142.840 2698.210 2143.100 ;
        RECT 2694.670 2142.020 2694.990 2142.080 ;
        RECT 2696.985 2142.020 2697.275 2142.065 ;
        RECT 2694.670 2141.880 2697.275 2142.020 ;
        RECT 2694.670 2141.820 2694.990 2141.880 ;
        RECT 2696.985 2141.835 2697.275 2141.880 ;
        RECT 2411.850 2139.180 2412.170 2139.240 ;
        RECT 2611.490 2139.180 2611.810 2139.240 ;
        RECT 2411.850 2139.040 2611.810 2139.180 ;
        RECT 2411.850 2138.980 2412.170 2139.040 ;
        RECT 2611.490 2138.980 2611.810 2139.040 ;
        RECT 2697.905 2137.600 2698.195 2137.645 ;
        RECT 2698.810 2137.600 2699.130 2137.660 ;
        RECT 2697.905 2137.460 2699.130 2137.600 ;
        RECT 2697.905 2137.415 2698.195 2137.460 ;
        RECT 2698.810 2137.400 2699.130 2137.460 ;
        RECT 2694.670 2136.580 2694.990 2136.640 ;
        RECT 2696.985 2136.580 2697.275 2136.625 ;
        RECT 2694.670 2136.440 2697.275 2136.580 ;
        RECT 2694.670 2136.380 2694.990 2136.440 ;
        RECT 2696.985 2136.395 2697.275 2136.440 ;
        RECT 2523.545 2135.005 2523.865 2135.265 ;
        RECT 2698.350 2132.160 2698.670 2132.220 ;
        RECT 2699.285 2132.160 2699.575 2132.205 ;
        RECT 2698.350 2132.020 2699.575 2132.160 ;
        RECT 2698.350 2131.960 2698.670 2132.020 ;
        RECT 2699.285 2131.975 2699.575 2132.020 ;
        RECT 2702.490 2131.960 2702.810 2132.220 ;
        RECT 2697.905 2131.820 2698.195 2131.865 ;
        RECT 2702.580 2131.820 2702.720 2131.960 ;
        RECT 2697.905 2131.680 2702.720 2131.820 ;
        RECT 2697.905 2131.635 2698.195 2131.680 ;
        RECT 2694.670 2131.140 2694.990 2131.200 ;
        RECT 2696.985 2131.140 2697.275 2131.185 ;
        RECT 2694.670 2131.000 2697.275 2131.140 ;
        RECT 2694.670 2130.940 2694.990 2131.000 ;
        RECT 2696.985 2130.955 2697.275 2131.000 ;
        RECT 2698.350 2130.940 2698.670 2131.200 ;
        RECT 2523.545 2127.475 2523.865 2127.735 ;
        RECT 2523.545 2121.495 2523.865 2121.755 ;
        RECT 2523.545 2115.550 2523.865 2115.810 ;
        RECT 2523.545 2109.905 2523.865 2110.165 ;
        RECT 2523.545 2103.900 2523.865 2104.160 ;
        RECT 2359.545 2058.055 2359.835 2058.285 ;
        RECT 2368.125 2058.055 2368.415 2058.285 ;
        RECT 2373.740 2058.055 2374.030 2058.285 ;
        RECT 2359.605 2057.605 2359.775 2058.055 ;
        RECT 2368.185 2057.710 2368.355 2058.055 ;
        RECT 2359.515 2057.315 2359.865 2057.605 ;
        RECT 2368.105 2057.360 2368.475 2057.710 ;
        RECT 2373.800 2057.575 2373.970 2058.055 ;
        RECT 2375.530 2058.025 2375.825 2058.285 ;
        RECT 2374.710 2057.575 2375.060 2057.605 ;
        RECT 2373.800 2057.545 2375.060 2057.575 ;
        RECT 2373.740 2057.405 2375.060 2057.545 ;
        RECT 2368.105 2057.340 2368.415 2057.360 ;
        RECT 2368.125 2057.315 2368.415 2057.340 ;
        RECT 2373.740 2057.315 2374.030 2057.405 ;
        RECT 2374.710 2057.315 2375.060 2057.405 ;
        RECT 2368.555 2057.145 2368.845 2057.175 ;
        RECT 2368.385 2057.140 2368.845 2057.145 ;
        RECT 2369.590 2057.140 2369.940 2057.240 ;
        RECT 2374.195 2057.175 2374.520 2057.265 ;
        RECT 2374.170 2057.145 2374.520 2057.175 ;
        RECT 2374.000 2057.140 2374.520 2057.145 ;
        RECT 2368.385 2056.975 2374.520 2057.140 ;
        RECT 2368.555 2056.970 2374.520 2056.975 ;
        RECT 2368.555 2056.945 2368.845 2056.970 ;
        RECT 2369.590 2056.890 2369.940 2056.970 ;
        RECT 2374.170 2056.945 2374.520 2056.970 ;
        RECT 2374.195 2056.940 2374.520 2056.945 ;
        RECT 2375.590 2056.925 2375.760 2058.025 ;
        RECT 2376.525 2058.020 2376.820 2058.280 ;
        RECT 2384.450 2058.055 2384.740 2058.285 ;
        RECT 2390.065 2058.055 2390.355 2058.285 ;
        RECT 2376.585 2057.290 2376.755 2058.020 ;
        RECT 2384.510 2057.710 2384.680 2058.055 ;
        RECT 2384.430 2057.360 2384.800 2057.710 ;
        RECT 2390.125 2057.575 2390.295 2058.055 ;
        RECT 2391.855 2058.025 2392.150 2058.285 ;
        RECT 2391.035 2057.575 2391.385 2057.605 ;
        RECT 2390.125 2057.545 2391.385 2057.575 ;
        RECT 2390.065 2057.405 2391.385 2057.545 ;
        RECT 2384.430 2057.340 2384.740 2057.360 ;
        RECT 2384.450 2057.315 2384.740 2057.340 ;
        RECT 2390.065 2057.315 2390.355 2057.405 ;
        RECT 2391.035 2057.315 2391.385 2057.405 ;
        RECT 2375.530 2056.920 2375.760 2056.925 ;
        RECT 2376.575 2056.940 2376.925 2057.290 ;
        RECT 2385.080 2057.175 2385.430 2057.245 ;
        RECT 2390.520 2057.175 2390.845 2057.265 ;
        RECT 2384.880 2057.145 2385.430 2057.175 ;
        RECT 2390.495 2057.145 2390.845 2057.175 ;
        RECT 2384.710 2057.140 2385.430 2057.145 ;
        RECT 2390.325 2057.140 2390.845 2057.145 ;
        RECT 2384.710 2056.975 2390.845 2057.140 ;
        RECT 2384.880 2056.970 2390.845 2056.975 ;
        RECT 2384.880 2056.945 2385.430 2056.970 ;
        RECT 2390.495 2056.945 2390.845 2056.970 ;
        RECT 2376.575 2056.920 2376.875 2056.940 ;
        RECT 2359.140 2056.785 2359.490 2056.860 ;
        RECT 2373.395 2056.815 2373.715 2056.830 ;
        RECT 2373.370 2056.785 2373.715 2056.815 ;
        RECT 2359.000 2056.615 2359.490 2056.785 ;
        RECT 2373.195 2056.615 2373.715 2056.785 ;
        RECT 2375.530 2056.685 2375.820 2056.920 ;
        RECT 2376.525 2056.835 2376.875 2056.920 ;
        RECT 2385.080 2056.895 2385.430 2056.945 ;
        RECT 2390.520 2056.940 2390.845 2056.945 ;
        RECT 2391.915 2056.925 2392.085 2058.025 ;
        RECT 2392.850 2058.020 2393.145 2058.280 ;
        RECT 2400.775 2058.055 2401.065 2058.285 ;
        RECT 2406.390 2058.055 2406.680 2058.285 ;
        RECT 2392.910 2057.300 2393.080 2058.020 ;
        RECT 2400.835 2057.710 2401.005 2058.055 ;
        RECT 2400.755 2057.360 2401.125 2057.710 ;
        RECT 2406.450 2057.575 2406.620 2058.055 ;
        RECT 2408.180 2058.025 2408.475 2058.285 ;
        RECT 2407.360 2057.575 2407.710 2057.605 ;
        RECT 2406.450 2057.545 2407.710 2057.575 ;
        RECT 2406.390 2057.405 2407.710 2057.545 ;
        RECT 2400.755 2057.340 2401.065 2057.360 ;
        RECT 2400.775 2057.315 2401.065 2057.340 ;
        RECT 2406.390 2057.315 2406.680 2057.405 ;
        RECT 2407.360 2057.315 2407.710 2057.405 ;
        RECT 2391.855 2056.920 2392.085 2056.925 ;
        RECT 2392.895 2056.945 2393.250 2057.300 ;
        RECT 2401.405 2057.175 2401.755 2057.250 ;
        RECT 2406.845 2057.175 2407.170 2057.265 ;
        RECT 2401.205 2057.145 2401.755 2057.175 ;
        RECT 2406.820 2057.145 2407.170 2057.175 ;
        RECT 2401.035 2057.140 2401.755 2057.145 ;
        RECT 2406.650 2057.140 2407.170 2057.145 ;
        RECT 2401.035 2056.975 2407.170 2057.140 ;
        RECT 2401.205 2056.970 2407.170 2056.975 ;
        RECT 2401.205 2056.945 2401.755 2056.970 ;
        RECT 2406.820 2056.945 2407.170 2056.970 ;
        RECT 2392.895 2056.920 2393.200 2056.945 ;
        RECT 2376.525 2056.680 2376.815 2056.835 ;
        RECT 2389.720 2056.815 2390.040 2056.830 ;
        RECT 2389.695 2056.785 2390.040 2056.815 ;
        RECT 2389.520 2056.615 2390.040 2056.785 ;
        RECT 2391.855 2056.685 2392.145 2056.920 ;
        RECT 2392.850 2056.840 2393.200 2056.920 ;
        RECT 2401.405 2056.900 2401.755 2056.945 ;
        RECT 2406.845 2056.940 2407.170 2056.945 ;
        RECT 2408.240 2056.925 2408.410 2058.025 ;
        RECT 2409.175 2058.020 2409.470 2058.280 ;
        RECT 2417.100 2058.055 2417.390 2058.285 ;
        RECT 2422.715 2058.055 2423.005 2058.285 ;
        RECT 2409.235 2057.290 2409.405 2058.020 ;
        RECT 2417.160 2057.710 2417.330 2058.055 ;
        RECT 2417.080 2057.360 2417.450 2057.710 ;
        RECT 2422.775 2057.575 2422.945 2058.055 ;
        RECT 2424.505 2058.025 2424.800 2058.285 ;
        RECT 2423.685 2057.575 2424.035 2057.605 ;
        RECT 2422.775 2057.545 2424.035 2057.575 ;
        RECT 2422.715 2057.405 2424.035 2057.545 ;
        RECT 2417.080 2057.340 2417.390 2057.360 ;
        RECT 2417.100 2057.315 2417.390 2057.340 ;
        RECT 2422.715 2057.315 2423.005 2057.405 ;
        RECT 2423.685 2057.315 2424.035 2057.405 ;
        RECT 2408.180 2056.920 2408.410 2056.925 ;
        RECT 2409.180 2056.940 2409.530 2057.290 ;
        RECT 2417.730 2057.175 2418.080 2057.245 ;
        RECT 2423.170 2057.175 2423.495 2057.265 ;
        RECT 2417.530 2057.145 2418.080 2057.175 ;
        RECT 2423.145 2057.145 2423.495 2057.175 ;
        RECT 2417.360 2057.140 2418.080 2057.145 ;
        RECT 2422.975 2057.140 2423.495 2057.145 ;
        RECT 2417.360 2056.975 2423.495 2057.140 ;
        RECT 2417.530 2056.970 2423.495 2056.975 ;
        RECT 2417.530 2056.945 2418.080 2056.970 ;
        RECT 2423.145 2056.945 2423.495 2056.970 ;
        RECT 2409.180 2056.920 2409.525 2056.940 ;
        RECT 2392.850 2056.680 2393.140 2056.840 ;
        RECT 2406.045 2056.815 2406.365 2056.830 ;
        RECT 2406.020 2056.785 2406.365 2056.815 ;
        RECT 2405.845 2056.615 2406.365 2056.785 ;
        RECT 2408.180 2056.685 2408.470 2056.920 ;
        RECT 2409.175 2056.840 2409.525 2056.920 ;
        RECT 2417.730 2056.895 2418.080 2056.945 ;
        RECT 2423.170 2056.940 2423.495 2056.945 ;
        RECT 2424.565 2056.925 2424.735 2058.025 ;
        RECT 2425.500 2058.020 2425.795 2058.280 ;
        RECT 2433.425 2058.055 2433.715 2058.285 ;
        RECT 2439.040 2058.055 2439.330 2058.285 ;
        RECT 2425.560 2057.290 2425.730 2058.020 ;
        RECT 2433.485 2057.710 2433.655 2058.055 ;
        RECT 2433.405 2057.360 2433.775 2057.710 ;
        RECT 2439.100 2057.575 2439.270 2058.055 ;
        RECT 2440.830 2058.025 2441.125 2058.285 ;
        RECT 2440.010 2057.575 2440.360 2057.605 ;
        RECT 2439.100 2057.545 2440.360 2057.575 ;
        RECT 2439.040 2057.405 2440.360 2057.545 ;
        RECT 2433.405 2057.340 2433.715 2057.360 ;
        RECT 2433.425 2057.315 2433.715 2057.340 ;
        RECT 2439.040 2057.315 2439.330 2057.405 ;
        RECT 2440.010 2057.315 2440.360 2057.405 ;
        RECT 2424.505 2056.920 2424.735 2056.925 ;
        RECT 2425.505 2056.940 2425.855 2057.290 ;
        RECT 2434.060 2057.175 2434.410 2057.245 ;
        RECT 2439.495 2057.175 2439.820 2057.265 ;
        RECT 2433.855 2057.145 2434.410 2057.175 ;
        RECT 2439.470 2057.145 2439.820 2057.175 ;
        RECT 2433.685 2057.140 2434.410 2057.145 ;
        RECT 2439.300 2057.140 2439.820 2057.145 ;
        RECT 2433.685 2056.975 2439.820 2057.140 ;
        RECT 2433.855 2056.970 2439.820 2056.975 ;
        RECT 2433.855 2056.945 2434.410 2056.970 ;
        RECT 2439.470 2056.945 2439.820 2056.970 ;
        RECT 2425.505 2056.920 2425.850 2056.940 ;
        RECT 2409.175 2056.680 2409.465 2056.840 ;
        RECT 2422.370 2056.815 2422.690 2056.830 ;
        RECT 2422.345 2056.785 2422.690 2056.815 ;
        RECT 2422.170 2056.615 2422.690 2056.785 ;
        RECT 2424.505 2056.685 2424.795 2056.920 ;
        RECT 2425.500 2056.845 2425.850 2056.920 ;
        RECT 2434.060 2056.895 2434.410 2056.945 ;
        RECT 2439.495 2056.940 2439.820 2056.945 ;
        RECT 2440.890 2056.925 2441.060 2058.025 ;
        RECT 2441.825 2058.020 2442.120 2058.280 ;
        RECT 2441.855 2058.005 2442.120 2058.020 ;
        RECT 2441.855 2057.910 2442.180 2058.005 ;
        RECT 2441.855 2057.560 2442.205 2057.910 ;
        RECT 2440.830 2056.920 2441.060 2056.925 ;
        RECT 2441.885 2056.920 2442.055 2057.560 ;
        RECT 2425.500 2056.680 2425.790 2056.845 ;
        RECT 2438.695 2056.815 2439.015 2056.830 ;
        RECT 2438.670 2056.785 2439.015 2056.815 ;
        RECT 2438.495 2056.615 2439.015 2056.785 ;
        RECT 2440.830 2056.685 2441.120 2056.920 ;
        RECT 2441.825 2056.915 2442.055 2056.920 ;
        RECT 2441.825 2056.680 2442.115 2056.915 ;
        RECT 2359.140 2056.570 2359.490 2056.615 ;
        RECT 2373.370 2056.585 2373.715 2056.615 ;
        RECT 2389.695 2056.585 2390.040 2056.615 ;
        RECT 2406.020 2056.585 2406.365 2056.615 ;
        RECT 2422.345 2056.585 2422.690 2056.615 ;
        RECT 2438.670 2056.585 2439.015 2056.615 ;
        RECT 2373.395 2056.540 2373.715 2056.585 ;
        RECT 2389.720 2056.540 2390.040 2056.585 ;
        RECT 2406.045 2056.540 2406.365 2056.585 ;
        RECT 2422.370 2056.540 2422.690 2056.585 ;
        RECT 2438.695 2056.540 2439.015 2056.585 ;
        RECT 2362.290 2053.065 2362.580 2053.105 ;
        RECT 2362.990 2053.065 2363.310 2053.125 ;
        RECT 2362.290 2052.925 2363.310 2053.065 ;
        RECT 2362.290 2052.875 2362.620 2052.925 ;
        RECT 2362.990 2052.865 2363.310 2052.925 ;
        RECT 2368.130 2053.065 2368.420 2053.105 ;
        RECT 2368.130 2052.875 2368.460 2053.065 ;
        RECT 2363.490 2052.785 2363.780 2052.825 ;
        RECT 2364.710 2052.785 2365.030 2052.845 ;
        RECT 2365.550 2052.825 2365.870 2052.845 ;
        RECT 2365.550 2052.785 2365.980 2052.825 ;
        RECT 2363.490 2052.595 2363.940 2052.785 ;
        RECT 2361.790 2052.305 2362.110 2052.565 ;
        RECT 2362.750 2052.545 2363.070 2052.565 ;
        RECT 2362.750 2052.315 2363.300 2052.545 ;
        RECT 2363.800 2052.365 2363.940 2052.595 ;
        RECT 2364.710 2052.645 2365.980 2052.785 ;
        RECT 2364.710 2052.585 2365.030 2052.645 ;
        RECT 2365.550 2052.595 2365.980 2052.645 ;
        RECT 2365.550 2052.585 2365.870 2052.595 ;
        RECT 2362.750 2052.305 2363.070 2052.315 ;
        RECT 2361.880 2051.385 2362.020 2052.305 ;
        RECT 2363.440 2052.225 2363.940 2052.365 ;
        RECT 2364.250 2052.315 2364.540 2052.545 ;
        RECT 2362.750 2051.985 2363.070 2052.005 ;
        RECT 2362.750 2051.755 2363.300 2051.985 ;
        RECT 2362.750 2051.745 2363.070 2051.755 ;
        RECT 2363.440 2051.445 2363.580 2052.225 ;
        RECT 2364.320 2052.005 2364.460 2052.315 ;
        RECT 2365.520 2052.265 2368.100 2052.365 ;
        RECT 2365.450 2052.225 2368.180 2052.265 ;
        RECT 2365.450 2052.035 2366.110 2052.225 ;
        RECT 2367.890 2052.035 2368.180 2052.225 ;
        RECT 2365.790 2052.025 2366.110 2052.035 ;
        RECT 2363.970 2051.985 2364.460 2052.005 ;
        RECT 2363.730 2051.755 2364.460 2051.985 ;
        RECT 2363.970 2051.745 2364.460 2051.755 ;
        RECT 2364.950 2051.745 2365.270 2052.005 ;
        RECT 2366.790 2051.985 2367.110 2052.005 ;
        RECT 2366.790 2051.755 2367.220 2051.985 ;
        RECT 2366.790 2051.745 2367.110 2051.755 ;
        RECT 2367.390 2051.745 2367.710 2052.005 ;
        RECT 2362.290 2051.385 2362.580 2051.425 ;
        RECT 2361.880 2051.245 2362.580 2051.385 ;
        RECT 2362.290 2051.195 2362.580 2051.245 ;
        RECT 2363.230 2051.245 2363.580 2051.445 ;
        RECT 2364.320 2051.385 2364.460 2051.745 ;
        RECT 2365.430 2051.665 2365.750 2051.725 ;
        RECT 2368.320 2051.705 2368.460 2052.875 ;
        RECT 2369.130 2052.845 2369.420 2053.105 ;
        RECT 2378.615 2053.065 2378.905 2053.105 ;
        RECT 2379.315 2053.065 2379.635 2053.125 ;
        RECT 2378.615 2052.925 2379.635 2053.065 ;
        RECT 2378.615 2052.875 2378.945 2052.925 ;
        RECT 2379.315 2052.865 2379.635 2052.925 ;
        RECT 2384.455 2053.065 2384.745 2053.105 ;
        RECT 2384.455 2052.875 2384.785 2053.065 ;
        RECT 2369.110 2052.585 2369.430 2052.845 ;
        RECT 2379.815 2052.785 2380.105 2052.825 ;
        RECT 2381.035 2052.785 2381.355 2052.845 ;
        RECT 2381.875 2052.825 2382.195 2052.845 ;
        RECT 2381.875 2052.785 2382.305 2052.825 ;
        RECT 2379.815 2052.595 2380.265 2052.785 ;
        RECT 2378.115 2052.305 2378.435 2052.565 ;
        RECT 2379.075 2052.545 2379.395 2052.565 ;
        RECT 2379.075 2052.315 2379.625 2052.545 ;
        RECT 2380.125 2052.365 2380.265 2052.595 ;
        RECT 2381.035 2052.645 2382.305 2052.785 ;
        RECT 2381.035 2052.585 2381.355 2052.645 ;
        RECT 2381.875 2052.595 2382.305 2052.645 ;
        RECT 2381.875 2052.585 2382.195 2052.595 ;
        RECT 2379.075 2052.305 2379.395 2052.315 ;
        RECT 2369.230 2051.985 2369.550 2052.005 ;
        RECT 2369.230 2051.745 2369.700 2051.985 ;
        RECT 2369.850 2051.945 2370.140 2051.985 ;
        RECT 2369.850 2051.805 2370.300 2051.945 ;
        RECT 2373.395 2051.875 2373.715 2051.945 ;
        RECT 2373.370 2051.845 2373.715 2051.875 ;
        RECT 2369.850 2051.755 2370.780 2051.805 ;
        RECT 2365.930 2051.665 2366.220 2051.705 ;
        RECT 2368.320 2051.665 2368.660 2051.705 ;
        RECT 2365.430 2051.525 2366.220 2051.665 ;
        RECT 2365.430 2051.465 2365.750 2051.525 ;
        RECT 2365.930 2051.475 2366.220 2051.525 ;
        RECT 2367.960 2051.525 2368.660 2051.665 ;
        RECT 2367.960 2051.505 2368.100 2051.525 ;
        RECT 2366.500 2051.445 2368.100 2051.505 ;
        RECT 2368.370 2051.475 2368.660 2051.525 ;
        RECT 2369.560 2051.505 2369.700 2051.745 ;
        RECT 2370.160 2051.725 2370.780 2051.755 ;
        RECT 2370.160 2051.665 2370.870 2051.725 ;
        RECT 2373.195 2051.675 2373.715 2051.845 ;
        RECT 2364.730 2051.385 2365.020 2051.425 ;
        RECT 2364.320 2051.245 2365.020 2051.385 ;
        RECT 2363.230 2051.185 2363.550 2051.245 ;
        RECT 2364.730 2051.195 2365.020 2051.245 ;
        RECT 2366.410 2051.365 2368.100 2051.445 ;
        RECT 2368.850 2051.425 2369.170 2051.445 ;
        RECT 2366.410 2051.195 2366.980 2051.365 ;
        RECT 2368.850 2051.195 2369.420 2051.425 ;
        RECT 2369.560 2051.385 2369.820 2051.505 ;
        RECT 2370.550 2051.465 2370.870 2051.665 ;
        RECT 2373.370 2051.645 2373.715 2051.675 ;
        RECT 2374.170 2051.490 2374.520 2051.610 ;
        RECT 2375.530 2051.540 2375.820 2051.775 ;
        RECT 2376.520 2051.545 2376.810 2051.780 ;
        RECT 2376.520 2051.540 2376.750 2051.545 ;
        RECT 2375.530 2051.535 2375.760 2051.540 ;
        RECT 2370.090 2051.385 2370.380 2051.425 ;
        RECT 2369.560 2051.365 2370.380 2051.385 ;
        RECT 2369.680 2051.245 2370.380 2051.365 ;
        RECT 2370.090 2051.195 2370.380 2051.245 ;
        RECT 2371.865 2051.320 2374.520 2051.490 ;
        RECT 2366.410 2051.185 2366.730 2051.195 ;
        RECT 2368.850 2051.185 2369.170 2051.195 ;
        RECT 2371.865 2051.105 2372.035 2051.320 ;
        RECT 2374.000 2051.315 2374.520 2051.320 ;
        RECT 2374.170 2051.260 2374.520 2051.315 ;
        RECT 2373.740 2051.120 2374.030 2051.145 ;
        RECT 2374.710 2051.120 2375.060 2051.145 ;
        RECT 2371.775 2050.755 2372.115 2051.105 ;
        RECT 2373.740 2050.950 2375.060 2051.120 ;
        RECT 2373.740 2050.915 2374.030 2050.950 ;
        RECT 2373.800 2050.405 2373.970 2050.915 ;
        RECT 2374.710 2050.855 2375.060 2050.950 ;
        RECT 2375.590 2050.435 2375.760 2051.535 ;
        RECT 2376.580 2050.440 2376.750 2051.540 ;
        RECT 2378.205 2051.385 2378.345 2052.305 ;
        RECT 2379.765 2052.225 2380.265 2052.365 ;
        RECT 2380.575 2052.315 2380.865 2052.545 ;
        RECT 2379.075 2051.985 2379.395 2052.005 ;
        RECT 2379.075 2051.755 2379.625 2051.985 ;
        RECT 2379.075 2051.745 2379.395 2051.755 ;
        RECT 2379.765 2051.445 2379.905 2052.225 ;
        RECT 2380.645 2052.005 2380.785 2052.315 ;
        RECT 2381.845 2052.265 2384.425 2052.365 ;
        RECT 2381.775 2052.225 2384.505 2052.265 ;
        RECT 2381.775 2052.035 2382.435 2052.225 ;
        RECT 2384.215 2052.035 2384.505 2052.225 ;
        RECT 2382.115 2052.025 2382.435 2052.035 ;
        RECT 2380.295 2051.985 2380.785 2052.005 ;
        RECT 2380.055 2051.755 2380.785 2051.985 ;
        RECT 2380.295 2051.745 2380.785 2051.755 ;
        RECT 2381.275 2051.745 2381.595 2052.005 ;
        RECT 2383.115 2051.985 2383.435 2052.005 ;
        RECT 2383.115 2051.755 2383.545 2051.985 ;
        RECT 2383.115 2051.745 2383.435 2051.755 ;
        RECT 2383.715 2051.745 2384.035 2052.005 ;
        RECT 2378.615 2051.385 2378.905 2051.425 ;
        RECT 2378.205 2051.245 2378.905 2051.385 ;
        RECT 2378.615 2051.195 2378.905 2051.245 ;
        RECT 2379.555 2051.245 2379.905 2051.445 ;
        RECT 2380.645 2051.385 2380.785 2051.745 ;
        RECT 2381.755 2051.665 2382.075 2051.725 ;
        RECT 2384.645 2051.705 2384.785 2052.875 ;
        RECT 2385.455 2052.845 2385.745 2053.105 ;
        RECT 2394.940 2053.065 2395.230 2053.105 ;
        RECT 2395.640 2053.065 2395.960 2053.125 ;
        RECT 2394.940 2052.925 2395.960 2053.065 ;
        RECT 2394.940 2052.875 2395.270 2052.925 ;
        RECT 2395.640 2052.865 2395.960 2052.925 ;
        RECT 2400.780 2053.065 2401.070 2053.105 ;
        RECT 2400.780 2052.875 2401.110 2053.065 ;
        RECT 2385.435 2052.585 2385.755 2052.845 ;
        RECT 2396.140 2052.785 2396.430 2052.825 ;
        RECT 2397.360 2052.785 2397.680 2052.845 ;
        RECT 2398.200 2052.825 2398.520 2052.845 ;
        RECT 2398.200 2052.785 2398.630 2052.825 ;
        RECT 2396.140 2052.595 2396.590 2052.785 ;
        RECT 2394.440 2052.305 2394.760 2052.565 ;
        RECT 2395.400 2052.545 2395.720 2052.565 ;
        RECT 2395.400 2052.315 2395.950 2052.545 ;
        RECT 2396.450 2052.365 2396.590 2052.595 ;
        RECT 2397.360 2052.645 2398.630 2052.785 ;
        RECT 2397.360 2052.585 2397.680 2052.645 ;
        RECT 2398.200 2052.595 2398.630 2052.645 ;
        RECT 2398.200 2052.585 2398.520 2052.595 ;
        RECT 2395.400 2052.305 2395.720 2052.315 ;
        RECT 2392.990 2052.185 2393.310 2052.200 ;
        RECT 2385.555 2051.985 2385.875 2052.005 ;
        RECT 2385.555 2051.745 2386.025 2051.985 ;
        RECT 2386.175 2051.945 2386.465 2051.985 ;
        RECT 2392.845 2051.955 2393.310 2052.185 ;
        RECT 2386.175 2051.805 2386.625 2051.945 ;
        RECT 2389.720 2051.875 2390.040 2051.945 ;
        RECT 2392.990 2051.940 2393.310 2051.955 ;
        RECT 2389.695 2051.845 2390.040 2051.875 ;
        RECT 2386.175 2051.755 2387.105 2051.805 ;
        RECT 2382.255 2051.665 2382.545 2051.705 ;
        RECT 2384.645 2051.665 2384.985 2051.705 ;
        RECT 2381.755 2051.525 2382.545 2051.665 ;
        RECT 2381.755 2051.465 2382.075 2051.525 ;
        RECT 2382.255 2051.475 2382.545 2051.525 ;
        RECT 2384.285 2051.525 2384.985 2051.665 ;
        RECT 2384.285 2051.505 2384.425 2051.525 ;
        RECT 2382.825 2051.445 2384.425 2051.505 ;
        RECT 2384.695 2051.475 2384.985 2051.525 ;
        RECT 2385.885 2051.505 2386.025 2051.745 ;
        RECT 2386.485 2051.725 2387.105 2051.755 ;
        RECT 2386.485 2051.665 2387.195 2051.725 ;
        RECT 2389.520 2051.675 2390.040 2051.845 ;
        RECT 2381.055 2051.385 2381.345 2051.425 ;
        RECT 2380.645 2051.245 2381.345 2051.385 ;
        RECT 2379.555 2051.185 2379.875 2051.245 ;
        RECT 2381.055 2051.195 2381.345 2051.245 ;
        RECT 2382.735 2051.365 2384.425 2051.445 ;
        RECT 2385.175 2051.425 2385.495 2051.445 ;
        RECT 2382.735 2051.195 2383.305 2051.365 ;
        RECT 2385.175 2051.195 2385.745 2051.425 ;
        RECT 2385.885 2051.385 2386.145 2051.505 ;
        RECT 2386.875 2051.465 2387.195 2051.665 ;
        RECT 2389.695 2051.645 2390.040 2051.675 ;
        RECT 2390.495 2051.490 2390.845 2051.610 ;
        RECT 2391.855 2051.540 2392.145 2051.775 ;
        RECT 2392.845 2051.545 2393.135 2051.780 ;
        RECT 2392.845 2051.540 2393.075 2051.545 ;
        RECT 2391.855 2051.535 2392.085 2051.540 ;
        RECT 2386.415 2051.385 2386.705 2051.425 ;
        RECT 2385.885 2051.365 2386.705 2051.385 ;
        RECT 2386.005 2051.245 2386.705 2051.365 ;
        RECT 2386.415 2051.195 2386.705 2051.245 ;
        RECT 2388.190 2051.320 2390.845 2051.490 ;
        RECT 2382.735 2051.185 2383.055 2051.195 ;
        RECT 2385.175 2051.185 2385.495 2051.195 ;
        RECT 2388.190 2051.105 2388.360 2051.320 ;
        RECT 2390.325 2051.315 2390.845 2051.320 ;
        RECT 2390.495 2051.260 2390.845 2051.315 ;
        RECT 2390.065 2051.120 2390.355 2051.145 ;
        RECT 2391.035 2051.120 2391.385 2051.145 ;
        RECT 2388.100 2050.755 2388.440 2051.105 ;
        RECT 2390.065 2050.950 2391.385 2051.120 ;
        RECT 2390.065 2050.915 2390.355 2050.950 ;
        RECT 2373.740 2050.175 2374.030 2050.405 ;
        RECT 2375.530 2050.175 2375.825 2050.435 ;
        RECT 2376.430 2050.180 2376.815 2050.440 ;
        RECT 2390.125 2050.405 2390.295 2050.915 ;
        RECT 2391.035 2050.855 2391.385 2050.950 ;
        RECT 2391.915 2050.435 2392.085 2051.535 ;
        RECT 2392.905 2050.440 2393.075 2051.540 ;
        RECT 2394.530 2051.385 2394.670 2052.305 ;
        RECT 2396.090 2052.225 2396.590 2052.365 ;
        RECT 2396.900 2052.315 2397.190 2052.545 ;
        RECT 2395.400 2051.985 2395.720 2052.005 ;
        RECT 2395.400 2051.755 2395.950 2051.985 ;
        RECT 2395.400 2051.745 2395.720 2051.755 ;
        RECT 2396.090 2051.445 2396.230 2052.225 ;
        RECT 2396.970 2052.005 2397.110 2052.315 ;
        RECT 2398.170 2052.265 2400.750 2052.365 ;
        RECT 2398.100 2052.225 2400.830 2052.265 ;
        RECT 2398.100 2052.035 2398.760 2052.225 ;
        RECT 2400.540 2052.035 2400.830 2052.225 ;
        RECT 2398.440 2052.025 2398.760 2052.035 ;
        RECT 2396.620 2051.985 2397.110 2052.005 ;
        RECT 2396.380 2051.755 2397.110 2051.985 ;
        RECT 2396.620 2051.745 2397.110 2051.755 ;
        RECT 2397.600 2051.745 2397.920 2052.005 ;
        RECT 2399.440 2051.985 2399.760 2052.005 ;
        RECT 2399.440 2051.755 2399.870 2051.985 ;
        RECT 2399.440 2051.745 2399.760 2051.755 ;
        RECT 2400.040 2051.745 2400.360 2052.005 ;
        RECT 2394.940 2051.385 2395.230 2051.425 ;
        RECT 2394.530 2051.245 2395.230 2051.385 ;
        RECT 2394.940 2051.195 2395.230 2051.245 ;
        RECT 2395.880 2051.245 2396.230 2051.445 ;
        RECT 2396.970 2051.385 2397.110 2051.745 ;
        RECT 2398.080 2051.665 2398.400 2051.725 ;
        RECT 2400.970 2051.705 2401.110 2052.875 ;
        RECT 2401.780 2052.845 2402.070 2053.105 ;
        RECT 2411.265 2053.065 2411.555 2053.105 ;
        RECT 2411.965 2053.065 2412.285 2053.125 ;
        RECT 2411.265 2052.925 2412.285 2053.065 ;
        RECT 2411.265 2052.875 2411.595 2052.925 ;
        RECT 2411.965 2052.865 2412.285 2052.925 ;
        RECT 2417.105 2053.065 2417.395 2053.105 ;
        RECT 2417.105 2052.875 2417.435 2053.065 ;
        RECT 2401.760 2052.585 2402.080 2052.845 ;
        RECT 2412.465 2052.785 2412.755 2052.825 ;
        RECT 2413.685 2052.785 2414.005 2052.845 ;
        RECT 2414.525 2052.825 2414.845 2052.845 ;
        RECT 2414.525 2052.785 2414.955 2052.825 ;
        RECT 2412.465 2052.595 2412.915 2052.785 ;
        RECT 2410.765 2052.305 2411.085 2052.565 ;
        RECT 2411.725 2052.545 2412.045 2052.565 ;
        RECT 2411.725 2052.315 2412.275 2052.545 ;
        RECT 2412.775 2052.365 2412.915 2052.595 ;
        RECT 2413.685 2052.645 2414.955 2052.785 ;
        RECT 2413.685 2052.585 2414.005 2052.645 ;
        RECT 2414.525 2052.595 2414.955 2052.645 ;
        RECT 2414.525 2052.585 2414.845 2052.595 ;
        RECT 2411.725 2052.305 2412.045 2052.315 ;
        RECT 2401.880 2051.985 2402.200 2052.005 ;
        RECT 2401.880 2051.745 2402.350 2051.985 ;
        RECT 2402.500 2051.945 2402.790 2051.985 ;
        RECT 2402.500 2051.805 2402.950 2051.945 ;
        RECT 2406.045 2051.875 2406.365 2051.945 ;
        RECT 2406.020 2051.845 2406.365 2051.875 ;
        RECT 2402.500 2051.755 2403.430 2051.805 ;
        RECT 2398.580 2051.665 2398.870 2051.705 ;
        RECT 2400.970 2051.665 2401.310 2051.705 ;
        RECT 2398.080 2051.525 2398.870 2051.665 ;
        RECT 2398.080 2051.465 2398.400 2051.525 ;
        RECT 2398.580 2051.475 2398.870 2051.525 ;
        RECT 2400.610 2051.525 2401.310 2051.665 ;
        RECT 2400.610 2051.505 2400.750 2051.525 ;
        RECT 2399.150 2051.445 2400.750 2051.505 ;
        RECT 2401.020 2051.475 2401.310 2051.525 ;
        RECT 2402.210 2051.505 2402.350 2051.745 ;
        RECT 2402.810 2051.725 2403.430 2051.755 ;
        RECT 2402.810 2051.665 2403.520 2051.725 ;
        RECT 2405.845 2051.675 2406.365 2051.845 ;
        RECT 2397.380 2051.385 2397.670 2051.425 ;
        RECT 2396.970 2051.245 2397.670 2051.385 ;
        RECT 2395.880 2051.185 2396.200 2051.245 ;
        RECT 2397.380 2051.195 2397.670 2051.245 ;
        RECT 2399.060 2051.365 2400.750 2051.445 ;
        RECT 2401.500 2051.425 2401.820 2051.445 ;
        RECT 2399.060 2051.195 2399.630 2051.365 ;
        RECT 2401.500 2051.195 2402.070 2051.425 ;
        RECT 2402.210 2051.385 2402.470 2051.505 ;
        RECT 2403.200 2051.465 2403.520 2051.665 ;
        RECT 2406.020 2051.645 2406.365 2051.675 ;
        RECT 2406.820 2051.490 2407.170 2051.610 ;
        RECT 2408.180 2051.540 2408.470 2051.775 ;
        RECT 2409.170 2051.545 2409.460 2051.780 ;
        RECT 2409.170 2051.540 2409.400 2051.545 ;
        RECT 2408.180 2051.535 2408.410 2051.540 ;
        RECT 2402.740 2051.385 2403.030 2051.425 ;
        RECT 2402.210 2051.365 2403.030 2051.385 ;
        RECT 2402.330 2051.245 2403.030 2051.365 ;
        RECT 2402.740 2051.195 2403.030 2051.245 ;
        RECT 2404.515 2051.320 2407.170 2051.490 ;
        RECT 2399.060 2051.185 2399.380 2051.195 ;
        RECT 2401.500 2051.185 2401.820 2051.195 ;
        RECT 2404.515 2051.105 2404.685 2051.320 ;
        RECT 2406.650 2051.315 2407.170 2051.320 ;
        RECT 2406.820 2051.260 2407.170 2051.315 ;
        RECT 2406.390 2051.120 2406.680 2051.145 ;
        RECT 2407.360 2051.120 2407.710 2051.145 ;
        RECT 2404.425 2050.755 2404.765 2051.105 ;
        RECT 2406.390 2050.950 2407.710 2051.120 ;
        RECT 2406.390 2050.915 2406.680 2050.950 ;
        RECT 2390.065 2050.175 2390.355 2050.405 ;
        RECT 2391.855 2050.175 2392.150 2050.435 ;
        RECT 2392.845 2050.180 2393.140 2050.440 ;
        RECT 2406.450 2050.405 2406.620 2050.915 ;
        RECT 2407.360 2050.855 2407.710 2050.950 ;
        RECT 2408.240 2050.435 2408.410 2051.535 ;
        RECT 2409.230 2050.440 2409.400 2051.540 ;
        RECT 2410.855 2051.385 2410.995 2052.305 ;
        RECT 2412.415 2052.225 2412.915 2052.365 ;
        RECT 2413.225 2052.315 2413.515 2052.545 ;
        RECT 2411.725 2051.985 2412.045 2052.005 ;
        RECT 2411.725 2051.755 2412.275 2051.985 ;
        RECT 2411.725 2051.745 2412.045 2051.755 ;
        RECT 2412.415 2051.445 2412.555 2052.225 ;
        RECT 2413.295 2052.005 2413.435 2052.315 ;
        RECT 2414.495 2052.265 2417.075 2052.365 ;
        RECT 2414.425 2052.225 2417.155 2052.265 ;
        RECT 2414.425 2052.035 2415.085 2052.225 ;
        RECT 2416.865 2052.035 2417.155 2052.225 ;
        RECT 2414.765 2052.025 2415.085 2052.035 ;
        RECT 2412.945 2051.985 2413.435 2052.005 ;
        RECT 2412.705 2051.755 2413.435 2051.985 ;
        RECT 2412.945 2051.745 2413.435 2051.755 ;
        RECT 2413.925 2051.745 2414.245 2052.005 ;
        RECT 2415.765 2051.985 2416.085 2052.005 ;
        RECT 2415.765 2051.755 2416.195 2051.985 ;
        RECT 2415.765 2051.745 2416.085 2051.755 ;
        RECT 2416.365 2051.745 2416.685 2052.005 ;
        RECT 2411.265 2051.385 2411.555 2051.425 ;
        RECT 2410.855 2051.245 2411.555 2051.385 ;
        RECT 2411.265 2051.195 2411.555 2051.245 ;
        RECT 2412.205 2051.245 2412.555 2051.445 ;
        RECT 2413.295 2051.385 2413.435 2051.745 ;
        RECT 2414.405 2051.665 2414.725 2051.725 ;
        RECT 2417.295 2051.705 2417.435 2052.875 ;
        RECT 2418.105 2052.845 2418.395 2053.105 ;
        RECT 2427.590 2053.065 2427.880 2053.105 ;
        RECT 2428.290 2053.065 2428.610 2053.125 ;
        RECT 2427.590 2052.925 2428.610 2053.065 ;
        RECT 2427.590 2052.875 2427.920 2052.925 ;
        RECT 2428.290 2052.865 2428.610 2052.925 ;
        RECT 2433.430 2053.065 2433.720 2053.105 ;
        RECT 2433.430 2052.875 2433.760 2053.065 ;
        RECT 2418.085 2052.585 2418.405 2052.845 ;
        RECT 2428.790 2052.785 2429.080 2052.825 ;
        RECT 2430.010 2052.785 2430.330 2052.845 ;
        RECT 2430.850 2052.825 2431.170 2052.845 ;
        RECT 2430.850 2052.785 2431.280 2052.825 ;
        RECT 2428.790 2052.595 2429.240 2052.785 ;
        RECT 2427.090 2052.305 2427.410 2052.565 ;
        RECT 2428.050 2052.545 2428.370 2052.565 ;
        RECT 2428.050 2052.315 2428.600 2052.545 ;
        RECT 2429.100 2052.365 2429.240 2052.595 ;
        RECT 2430.010 2052.645 2431.280 2052.785 ;
        RECT 2430.010 2052.585 2430.330 2052.645 ;
        RECT 2430.850 2052.595 2431.280 2052.645 ;
        RECT 2430.850 2052.585 2431.170 2052.595 ;
        RECT 2428.050 2052.305 2428.370 2052.315 ;
        RECT 2425.650 2052.185 2425.970 2052.200 ;
        RECT 2418.205 2051.985 2418.525 2052.005 ;
        RECT 2418.205 2051.745 2418.675 2051.985 ;
        RECT 2418.825 2051.945 2419.115 2051.985 ;
        RECT 2425.495 2051.955 2425.970 2052.185 ;
        RECT 2418.825 2051.805 2419.275 2051.945 ;
        RECT 2422.370 2051.875 2422.690 2051.945 ;
        RECT 2425.650 2051.940 2425.970 2051.955 ;
        RECT 2422.345 2051.845 2422.690 2051.875 ;
        RECT 2418.825 2051.755 2419.755 2051.805 ;
        RECT 2414.905 2051.665 2415.195 2051.705 ;
        RECT 2417.295 2051.665 2417.635 2051.705 ;
        RECT 2414.405 2051.525 2415.195 2051.665 ;
        RECT 2414.405 2051.465 2414.725 2051.525 ;
        RECT 2414.905 2051.475 2415.195 2051.525 ;
        RECT 2416.935 2051.525 2417.635 2051.665 ;
        RECT 2416.935 2051.505 2417.075 2051.525 ;
        RECT 2415.475 2051.445 2417.075 2051.505 ;
        RECT 2417.345 2051.475 2417.635 2051.525 ;
        RECT 2418.535 2051.505 2418.675 2051.745 ;
        RECT 2419.135 2051.725 2419.755 2051.755 ;
        RECT 2419.135 2051.665 2419.845 2051.725 ;
        RECT 2422.170 2051.675 2422.690 2051.845 ;
        RECT 2413.705 2051.385 2413.995 2051.425 ;
        RECT 2413.295 2051.245 2413.995 2051.385 ;
        RECT 2412.205 2051.185 2412.525 2051.245 ;
        RECT 2413.705 2051.195 2413.995 2051.245 ;
        RECT 2415.385 2051.365 2417.075 2051.445 ;
        RECT 2417.825 2051.425 2418.145 2051.445 ;
        RECT 2415.385 2051.195 2415.955 2051.365 ;
        RECT 2417.825 2051.195 2418.395 2051.425 ;
        RECT 2418.535 2051.385 2418.795 2051.505 ;
        RECT 2419.525 2051.465 2419.845 2051.665 ;
        RECT 2422.345 2051.645 2422.690 2051.675 ;
        RECT 2423.145 2051.490 2423.495 2051.610 ;
        RECT 2424.505 2051.540 2424.795 2051.775 ;
        RECT 2425.495 2051.545 2425.785 2051.780 ;
        RECT 2425.495 2051.540 2425.725 2051.545 ;
        RECT 2424.505 2051.535 2424.735 2051.540 ;
        RECT 2419.065 2051.385 2419.355 2051.425 ;
        RECT 2418.535 2051.365 2419.355 2051.385 ;
        RECT 2418.655 2051.245 2419.355 2051.365 ;
        RECT 2419.065 2051.195 2419.355 2051.245 ;
        RECT 2420.840 2051.320 2423.495 2051.490 ;
        RECT 2415.385 2051.185 2415.705 2051.195 ;
        RECT 2417.825 2051.185 2418.145 2051.195 ;
        RECT 2420.840 2051.105 2421.010 2051.320 ;
        RECT 2422.975 2051.315 2423.495 2051.320 ;
        RECT 2423.145 2051.260 2423.495 2051.315 ;
        RECT 2422.715 2051.120 2423.005 2051.145 ;
        RECT 2423.685 2051.120 2424.035 2051.145 ;
        RECT 2420.750 2050.755 2421.090 2051.105 ;
        RECT 2422.715 2050.950 2424.035 2051.120 ;
        RECT 2422.715 2050.915 2423.005 2050.950 ;
        RECT 2406.390 2050.175 2406.680 2050.405 ;
        RECT 2408.180 2050.175 2408.475 2050.435 ;
        RECT 2409.090 2050.180 2409.465 2050.440 ;
        RECT 2422.775 2050.405 2422.945 2050.915 ;
        RECT 2423.685 2050.855 2424.035 2050.950 ;
        RECT 2424.565 2050.435 2424.735 2051.535 ;
        RECT 2425.555 2050.440 2425.725 2051.540 ;
        RECT 2427.180 2051.385 2427.320 2052.305 ;
        RECT 2428.740 2052.225 2429.240 2052.365 ;
        RECT 2429.550 2052.315 2429.840 2052.545 ;
        RECT 2428.050 2051.985 2428.370 2052.005 ;
        RECT 2428.050 2051.755 2428.600 2051.985 ;
        RECT 2428.050 2051.745 2428.370 2051.755 ;
        RECT 2428.740 2051.445 2428.880 2052.225 ;
        RECT 2429.620 2052.005 2429.760 2052.315 ;
        RECT 2430.820 2052.265 2433.400 2052.365 ;
        RECT 2430.750 2052.225 2433.480 2052.265 ;
        RECT 2430.750 2052.035 2431.410 2052.225 ;
        RECT 2433.190 2052.035 2433.480 2052.225 ;
        RECT 2431.090 2052.025 2431.410 2052.035 ;
        RECT 2429.270 2051.985 2429.760 2052.005 ;
        RECT 2429.030 2051.755 2429.760 2051.985 ;
        RECT 2429.270 2051.745 2429.760 2051.755 ;
        RECT 2430.250 2051.745 2430.570 2052.005 ;
        RECT 2432.090 2051.985 2432.410 2052.005 ;
        RECT 2432.090 2051.755 2432.520 2051.985 ;
        RECT 2432.090 2051.745 2432.410 2051.755 ;
        RECT 2432.690 2051.745 2433.010 2052.005 ;
        RECT 2427.590 2051.385 2427.880 2051.425 ;
        RECT 2427.180 2051.245 2427.880 2051.385 ;
        RECT 2427.590 2051.195 2427.880 2051.245 ;
        RECT 2428.530 2051.245 2428.880 2051.445 ;
        RECT 2429.620 2051.385 2429.760 2051.745 ;
        RECT 2430.730 2051.665 2431.050 2051.725 ;
        RECT 2433.620 2051.705 2433.760 2052.875 ;
        RECT 2434.430 2052.845 2434.720 2053.105 ;
        RECT 2434.410 2052.585 2434.730 2052.845 ;
        RECT 2434.530 2051.985 2434.850 2052.005 ;
        RECT 2434.530 2051.745 2435.000 2051.985 ;
        RECT 2435.150 2051.945 2435.440 2051.985 ;
        RECT 2435.150 2051.805 2435.600 2051.945 ;
        RECT 2438.695 2051.875 2439.015 2051.945 ;
        RECT 2438.670 2051.845 2439.015 2051.875 ;
        RECT 2435.150 2051.755 2436.080 2051.805 ;
        RECT 2431.230 2051.665 2431.520 2051.705 ;
        RECT 2433.620 2051.665 2433.960 2051.705 ;
        RECT 2430.730 2051.525 2431.520 2051.665 ;
        RECT 2430.730 2051.465 2431.050 2051.525 ;
        RECT 2431.230 2051.475 2431.520 2051.525 ;
        RECT 2433.260 2051.525 2433.960 2051.665 ;
        RECT 2433.260 2051.505 2433.400 2051.525 ;
        RECT 2431.800 2051.445 2433.400 2051.505 ;
        RECT 2433.670 2051.475 2433.960 2051.525 ;
        RECT 2434.860 2051.505 2435.000 2051.745 ;
        RECT 2435.460 2051.725 2436.080 2051.755 ;
        RECT 2435.460 2051.665 2436.170 2051.725 ;
        RECT 2438.495 2051.675 2439.015 2051.845 ;
        RECT 2430.030 2051.385 2430.320 2051.425 ;
        RECT 2429.620 2051.245 2430.320 2051.385 ;
        RECT 2428.530 2051.185 2428.850 2051.245 ;
        RECT 2430.030 2051.195 2430.320 2051.245 ;
        RECT 2431.710 2051.365 2433.400 2051.445 ;
        RECT 2434.150 2051.425 2434.470 2051.445 ;
        RECT 2431.710 2051.195 2432.280 2051.365 ;
        RECT 2434.150 2051.195 2434.720 2051.425 ;
        RECT 2434.860 2051.385 2435.120 2051.505 ;
        RECT 2435.850 2051.465 2436.170 2051.665 ;
        RECT 2438.670 2051.645 2439.015 2051.675 ;
        RECT 2439.470 2051.490 2439.820 2051.610 ;
        RECT 2440.830 2051.540 2441.120 2051.775 ;
        RECT 2441.820 2051.545 2442.110 2051.780 ;
        RECT 2441.820 2051.540 2442.050 2051.545 ;
        RECT 2440.830 2051.535 2441.060 2051.540 ;
        RECT 2435.390 2051.385 2435.680 2051.425 ;
        RECT 2434.860 2051.365 2435.680 2051.385 ;
        RECT 2434.980 2051.245 2435.680 2051.365 ;
        RECT 2435.390 2051.195 2435.680 2051.245 ;
        RECT 2437.165 2051.320 2439.820 2051.490 ;
        RECT 2431.710 2051.185 2432.030 2051.195 ;
        RECT 2434.150 2051.185 2434.470 2051.195 ;
        RECT 2437.165 2051.105 2437.335 2051.320 ;
        RECT 2439.300 2051.315 2439.820 2051.320 ;
        RECT 2439.470 2051.260 2439.820 2051.315 ;
        RECT 2439.040 2051.120 2439.330 2051.145 ;
        RECT 2440.010 2051.120 2440.360 2051.145 ;
        RECT 2437.075 2050.755 2437.415 2051.105 ;
        RECT 2439.040 2050.950 2440.360 2051.120 ;
        RECT 2439.040 2050.915 2439.330 2050.950 ;
        RECT 2422.715 2050.175 2423.005 2050.405 ;
        RECT 2424.505 2050.175 2424.800 2050.435 ;
        RECT 2425.495 2050.180 2425.790 2050.440 ;
        RECT 2439.100 2050.405 2439.270 2050.915 ;
        RECT 2440.010 2050.855 2440.360 2050.950 ;
        RECT 2440.890 2050.435 2441.060 2051.535 ;
        RECT 2441.880 2050.440 2442.050 2051.540 ;
        RECT 2439.040 2050.175 2439.330 2050.405 ;
        RECT 2440.830 2050.175 2441.125 2050.435 ;
        RECT 2441.820 2050.380 2442.115 2050.440 ;
        RECT 2441.820 2050.240 2443.360 2050.380 ;
        RECT 2441.820 2050.180 2442.115 2050.240 ;
        RECT 2443.220 2050.100 2443.360 2050.240 ;
        RECT 2453.710 2050.100 2454.030 2050.160 ;
        RECT 2443.220 2049.960 2454.030 2050.100 ;
        RECT 2453.710 2049.900 2454.030 2049.960 ;
        RECT 2576.990 2049.080 2577.310 2049.140 ;
        RECT 2677.270 2049.080 2677.590 2049.140 ;
        RECT 2576.990 2048.940 2677.590 2049.080 ;
        RECT 2576.990 2048.880 2577.310 2048.940 ;
        RECT 2677.270 2048.880 2677.590 2048.940 ;
        RECT 2376.430 2042.280 2376.750 2042.340 ;
        RECT 2466.590 2042.280 2466.910 2042.340 ;
        RECT 2376.430 2042.140 2466.910 2042.280 ;
        RECT 2376.430 2042.080 2376.750 2042.140 ;
        RECT 2466.590 2042.080 2466.910 2042.140 ;
        RECT 2695.590 2036.480 2695.910 2036.540 ;
        RECT 2698.810 2036.480 2699.130 2036.540 ;
        RECT 2700.205 2036.480 2700.495 2036.525 ;
        RECT 2695.590 2036.340 2698.120 2036.480 ;
        RECT 2695.590 2036.280 2695.910 2036.340 ;
        RECT 2697.980 2036.140 2698.120 2036.340 ;
        RECT 2698.810 2036.340 2700.495 2036.480 ;
        RECT 2698.810 2036.280 2699.130 2036.340 ;
        RECT 2700.205 2036.295 2700.495 2036.340 ;
        RECT 2702.490 2036.480 2702.810 2036.540 ;
        RECT 2709.865 2036.480 2710.155 2036.525 ;
        RECT 2702.490 2036.340 2710.155 2036.480 ;
        RECT 2702.490 2036.280 2702.810 2036.340 ;
        RECT 2709.865 2036.295 2710.155 2036.340 ;
        RECT 2697.980 2036.000 2701.340 2036.140 ;
        RECT 2695.130 2035.800 2695.450 2035.860 ;
        RECT 2701.200 2035.845 2701.340 2036.000 ;
        RECT 2699.745 2035.800 2700.035 2035.845 ;
        RECT 2695.130 2035.660 2700.035 2035.800 ;
        RECT 2695.130 2035.600 2695.450 2035.660 ;
        RECT 2699.745 2035.615 2700.035 2035.660 ;
        RECT 2701.125 2035.615 2701.415 2035.845 ;
        RECT 2392.990 2035.480 2393.310 2035.540 ;
        RECT 2677.270 2035.480 2677.590 2035.540 ;
        RECT 2392.990 2035.340 2677.590 2035.480 ;
        RECT 2392.990 2035.280 2393.310 2035.340 ;
        RECT 2677.270 2035.280 2677.590 2035.340 ;
        RECT 2698.365 2035.460 2698.655 2035.505 ;
        RECT 2701.570 2035.460 2701.890 2035.520 ;
        RECT 2698.365 2035.320 2701.890 2035.460 ;
        RECT 2698.365 2035.275 2698.655 2035.320 ;
        RECT 2701.570 2035.260 2701.890 2035.320 ;
        RECT 2721.810 2034.920 2722.130 2035.180 ;
        RECT 2698.350 2034.780 2698.670 2034.840 ;
        RECT 2698.825 2034.780 2699.115 2034.825 ;
        RECT 2698.350 2034.640 2699.115 2034.780 ;
        RECT 2698.350 2034.580 2698.670 2034.640 ;
        RECT 2698.825 2034.595 2699.115 2034.640 ;
        RECT 2731.470 2034.580 2731.790 2034.840 ;
        RECT 2694.670 2032.740 2694.990 2032.800 ;
        RECT 2696.985 2032.740 2697.275 2032.785 ;
        RECT 2694.670 2032.600 2697.275 2032.740 ;
        RECT 2694.670 2032.540 2694.990 2032.600 ;
        RECT 2696.985 2032.555 2697.275 2032.600 ;
        RECT 2697.890 2031.860 2698.210 2032.120 ;
        RECT 2694.670 2024.920 2694.990 2024.980 ;
        RECT 2696.985 2024.920 2697.275 2024.965 ;
        RECT 2694.670 2024.780 2697.275 2024.920 ;
        RECT 2694.670 2024.720 2694.990 2024.780 ;
        RECT 2696.985 2024.735 2697.275 2024.780 ;
        RECT 2696.970 2023.900 2697.290 2023.960 ;
        RECT 2697.905 2023.900 2698.195 2023.945 ;
        RECT 2696.970 2023.760 2698.195 2023.900 ;
        RECT 2696.970 2023.700 2697.290 2023.760 ;
        RECT 2697.905 2023.715 2698.195 2023.760 ;
        RECT 2697.430 2022.200 2697.750 2022.260 ;
        RECT 2698.350 2022.200 2698.670 2022.260 ;
        RECT 2697.430 2022.060 2698.670 2022.200 ;
        RECT 2697.430 2022.000 2697.750 2022.060 ;
        RECT 2698.350 2022.000 2698.670 2022.060 ;
        RECT 2576.990 2021.880 2577.310 2021.940 ;
        RECT 2677.270 2021.880 2677.590 2021.940 ;
        RECT 2576.990 2021.740 2677.590 2021.880 ;
        RECT 2576.990 2021.680 2577.310 2021.740 ;
        RECT 2677.270 2021.680 2677.590 2021.740 ;
        RECT 2698.370 2019.820 2698.660 2019.865 ;
        RECT 2703.890 2019.820 2704.180 2019.865 ;
        RECT 2704.810 2019.820 2705.100 2019.865 ;
        RECT 2698.370 2019.680 2705.100 2019.820 ;
        RECT 2698.370 2019.635 2698.660 2019.680 ;
        RECT 2703.890 2019.635 2704.180 2019.680 ;
        RECT 2704.810 2019.635 2705.100 2019.680 ;
        RECT 2696.985 2019.480 2697.275 2019.525 ;
        RECT 2697.430 2019.480 2697.750 2019.540 ;
        RECT 2696.985 2019.340 2697.750 2019.480 ;
        RECT 2696.985 2019.295 2697.275 2019.340 ;
        RECT 2697.430 2019.280 2697.750 2019.340 ;
        RECT 2697.890 2019.280 2698.210 2019.540 ;
        RECT 2699.290 2019.480 2699.580 2019.525 ;
        RECT 2701.130 2019.480 2701.420 2019.525 ;
        RECT 2699.290 2019.340 2701.420 2019.480 ;
        RECT 2699.290 2019.295 2699.580 2019.340 ;
        RECT 2701.130 2019.295 2701.420 2019.340 ;
        RECT 2703.475 2019.480 2703.765 2019.525 ;
        RECT 2705.315 2019.480 2705.605 2019.525 ;
        RECT 2703.475 2019.340 2705.605 2019.480 ;
        RECT 2703.475 2019.295 2703.765 2019.340 ;
        RECT 2705.315 2019.295 2705.605 2019.340 ;
        RECT 2721.810 2019.280 2722.130 2019.540 ;
        RECT 2702.030 2019.185 2702.350 2019.200 ;
        RECT 2701.585 2019.140 2701.875 2019.185 ;
        RECT 2697.520 2019.000 2701.875 2019.140 ;
        RECT 2697.520 2018.860 2697.660 2019.000 ;
        RECT 2701.585 2018.955 2701.875 2019.000 ;
        RECT 2702.030 2018.955 2702.460 2019.185 ;
        RECT 2702.950 2019.140 2703.270 2019.200 ;
        RECT 2721.900 2019.140 2722.040 2019.280 ;
        RECT 2702.950 2019.000 2722.040 2019.140 ;
        RECT 2702.030 2018.940 2702.350 2018.955 ;
        RECT 2702.950 2018.940 2703.270 2019.000 ;
        RECT 2697.430 2018.600 2697.750 2018.860 ;
        RECT 2700.205 2018.615 2700.495 2018.845 ;
        RECT 2701.165 2018.800 2701.455 2018.845 ;
        RECT 2704.395 2018.800 2704.685 2018.845 ;
        RECT 2701.165 2018.660 2704.685 2018.800 ;
        RECT 2701.165 2018.615 2701.455 2018.660 ;
        RECT 2704.395 2018.615 2704.685 2018.660 ;
        RECT 2700.280 2018.460 2700.420 2018.615 ;
        RECT 2702.490 2018.460 2702.810 2018.520 ;
        RECT 2700.280 2018.320 2702.810 2018.460 ;
        RECT 2702.490 2018.260 2702.810 2018.320 ;
        RECT 2703.870 2018.460 2704.190 2018.520 ;
        RECT 2706.185 2018.460 2706.475 2018.505 ;
        RECT 2703.870 2018.320 2706.475 2018.460 ;
        RECT 2703.870 2018.260 2704.190 2018.320 ;
        RECT 2706.185 2018.275 2706.475 2018.320 ;
        RECT 2697.905 2017.440 2698.195 2017.485 ;
        RECT 2702.030 2017.440 2702.350 2017.500 ;
        RECT 2697.905 2017.300 2702.350 2017.440 ;
        RECT 2697.905 2017.255 2698.195 2017.300 ;
        RECT 2702.030 2017.240 2702.350 2017.300 ;
        RECT 2694.670 2016.420 2694.990 2016.480 ;
        RECT 2696.985 2016.420 2697.275 2016.465 ;
        RECT 2694.670 2016.280 2697.275 2016.420 ;
        RECT 2694.670 2016.220 2694.990 2016.280 ;
        RECT 2696.985 2016.235 2697.275 2016.280 ;
        RECT 2583.890 2015.080 2584.210 2015.140 ;
        RECT 2677.270 2015.080 2677.590 2015.140 ;
        RECT 2583.890 2014.940 2677.590 2015.080 ;
        RECT 2583.890 2014.880 2584.210 2014.940 ;
        RECT 2677.270 2014.880 2677.590 2014.940 ;
        RECT 2698.370 2014.380 2698.660 2014.425 ;
        RECT 2703.890 2014.380 2704.180 2014.425 ;
        RECT 2704.810 2014.380 2705.100 2014.425 ;
        RECT 2698.370 2014.240 2705.100 2014.380 ;
        RECT 2698.370 2014.195 2698.660 2014.240 ;
        RECT 2703.890 2014.195 2704.180 2014.240 ;
        RECT 2704.810 2014.195 2705.100 2014.240 ;
        RECT 2696.970 2013.840 2697.290 2014.100 ;
        RECT 2697.890 2013.840 2698.210 2014.100 ;
        RECT 2699.290 2014.040 2699.580 2014.085 ;
        RECT 2701.130 2014.040 2701.420 2014.085 ;
        RECT 2699.290 2013.900 2701.420 2014.040 ;
        RECT 2699.290 2013.855 2699.580 2013.900 ;
        RECT 2701.130 2013.855 2701.420 2013.900 ;
        RECT 2702.950 2013.840 2703.270 2014.100 ;
        RECT 2703.475 2014.040 2703.765 2014.085 ;
        RECT 2705.315 2014.040 2705.605 2014.085 ;
        RECT 2703.475 2013.900 2705.605 2014.040 ;
        RECT 2703.475 2013.855 2703.765 2013.900 ;
        RECT 2705.315 2013.855 2705.605 2013.900 ;
        RECT 2698.810 2013.700 2699.130 2013.760 ;
        RECT 2702.030 2013.745 2702.350 2013.760 ;
        RECT 2701.585 2013.700 2701.875 2013.745 ;
        RECT 2698.810 2013.560 2701.875 2013.700 ;
        RECT 2698.810 2013.500 2699.130 2013.560 ;
        RECT 2701.585 2013.515 2701.875 2013.560 ;
        RECT 2702.030 2013.515 2702.460 2013.745 ;
        RECT 2702.030 2013.500 2702.350 2013.515 ;
        RECT 2700.205 2013.175 2700.495 2013.405 ;
        RECT 2701.165 2013.360 2701.455 2013.405 ;
        RECT 2704.395 2013.360 2704.685 2013.405 ;
        RECT 2701.165 2013.220 2704.685 2013.360 ;
        RECT 2701.165 2013.175 2701.455 2013.220 ;
        RECT 2704.395 2013.175 2704.685 2013.220 ;
        RECT 2698.350 2013.020 2698.670 2013.080 ;
        RECT 2700.280 2013.020 2700.420 2013.175 ;
        RECT 2702.490 2013.020 2702.810 2013.080 ;
        RECT 2698.350 2012.880 2702.810 2013.020 ;
        RECT 2698.350 2012.820 2698.670 2012.880 ;
        RECT 2702.490 2012.820 2702.810 2012.880 ;
        RECT 2706.170 2012.820 2706.490 2013.080 ;
        RECT 2697.905 2012.000 2698.195 2012.045 ;
        RECT 2702.030 2012.000 2702.350 2012.060 ;
        RECT 2706.170 2012.000 2706.490 2012.060 ;
        RECT 2697.905 2011.860 2702.350 2012.000 ;
        RECT 2697.905 2011.815 2698.195 2011.860 ;
        RECT 2702.030 2011.800 2702.350 2011.860 ;
        RECT 2703.960 2011.860 2706.490 2012.000 ;
        RECT 2697.890 2011.320 2698.210 2011.380 ;
        RECT 2701.570 2011.320 2701.890 2011.380 ;
        RECT 2703.960 2011.365 2704.100 2011.860 ;
        RECT 2706.170 2011.800 2706.490 2011.860 ;
        RECT 2697.890 2011.180 2703.640 2011.320 ;
        RECT 2697.890 2011.120 2698.210 2011.180 ;
        RECT 2701.570 2011.120 2701.890 2011.180 ;
        RECT 2694.670 2010.980 2694.990 2011.040 ;
        RECT 2696.985 2010.980 2697.275 2011.025 ;
        RECT 2694.670 2010.840 2697.275 2010.980 ;
        RECT 2703.500 2010.980 2703.640 2011.180 ;
        RECT 2703.885 2011.135 2704.175 2011.365 ;
        RECT 2704.345 2011.135 2704.635 2011.365 ;
        RECT 2704.420 2010.980 2704.560 2011.135 ;
        RECT 2703.500 2010.840 2704.560 2010.980 ;
        RECT 2694.670 2010.780 2694.990 2010.840 ;
        RECT 2696.985 2010.795 2697.275 2010.840 ;
        RECT 2703.425 2010.640 2703.715 2010.685 ;
        RECT 2703.870 2010.640 2704.190 2010.700 ;
        RECT 2703.425 2010.500 2704.190 2010.640 ;
        RECT 2703.425 2010.455 2703.715 2010.500 ;
        RECT 2703.870 2010.440 2704.190 2010.500 ;
        RECT 2701.570 2010.100 2701.890 2010.360 ;
        RECT 2697.430 2006.560 2697.750 2006.620 ;
        RECT 2697.905 2006.560 2698.195 2006.605 ;
        RECT 2697.430 2006.420 2698.195 2006.560 ;
        RECT 2697.430 2006.360 2697.750 2006.420 ;
        RECT 2697.905 2006.375 2698.195 2006.420 ;
        RECT 2694.670 2005.540 2694.990 2005.600 ;
        RECT 2696.985 2005.540 2697.275 2005.585 ;
        RECT 2694.670 2005.400 2697.275 2005.540 ;
        RECT 2694.670 2005.340 2694.990 2005.400 ;
        RECT 2696.985 2005.355 2697.275 2005.400 ;
        RECT 2701.570 1999.900 2701.890 2000.160 ;
        RECT 2702.505 2000.100 2702.795 2000.145 ;
        RECT 2703.870 2000.100 2704.190 2000.160 ;
        RECT 2731.470 2000.100 2731.790 2000.160 ;
        RECT 2702.505 1999.960 2731.790 2000.100 ;
        RECT 2702.505 1999.915 2702.795 1999.960 ;
        RECT 2703.870 1999.900 2704.190 1999.960 ;
        RECT 2731.470 1999.900 2731.790 1999.960 ;
        RECT 2702.030 1999.220 2702.350 1999.480 ;
        RECT 2697.905 1998.400 2698.195 1998.445 ;
        RECT 2698.810 1998.400 2699.130 1998.460 ;
        RECT 2697.905 1998.260 2699.130 1998.400 ;
        RECT 2697.905 1998.215 2698.195 1998.260 ;
        RECT 2698.810 1998.200 2699.130 1998.260 ;
        RECT 2702.030 1998.200 2702.350 1998.460 ;
        RECT 2703.870 1998.200 2704.190 1998.460 ;
        RECT 2694.670 1997.720 2694.990 1997.780 ;
        RECT 2702.120 1997.765 2702.260 1998.200 ;
        RECT 2703.960 1997.765 2704.100 1998.200 ;
        RECT 2696.985 1997.720 2697.275 1997.765 ;
        RECT 2694.670 1997.580 2697.275 1997.720 ;
        RECT 2694.670 1997.520 2694.990 1997.580 ;
        RECT 2696.985 1997.535 2697.275 1997.580 ;
        RECT 2702.045 1997.535 2702.335 1997.765 ;
        RECT 2703.885 1997.535 2704.175 1997.765 ;
        RECT 2704.790 1997.180 2705.110 1997.440 ;
        RECT 2702.490 1996.840 2702.810 1997.100 ;
        RECT 2702.490 1995.680 2702.810 1995.740 ;
        RECT 2702.490 1995.540 2724.570 1995.680 ;
        RECT 2702.490 1995.480 2702.810 1995.540 ;
        RECT 2724.430 1994.660 2724.570 1995.540 ;
        RECT 2725.505 1994.660 2725.795 1994.705 ;
        RECT 2724.430 1994.520 2725.795 1994.660 ;
        RECT 2725.505 1994.475 2725.795 1994.520 ;
        RECT 2590.790 1994.340 2591.110 1994.400 ;
        RECT 2677.270 1994.340 2677.590 1994.400 ;
        RECT 2590.790 1994.200 2677.590 1994.340 ;
        RECT 2590.790 1994.140 2591.110 1994.200 ;
        RECT 2677.270 1994.140 2677.590 1994.200 ;
        RECT 2694.670 1992.280 2694.990 1992.340 ;
        RECT 2696.985 1992.280 2697.275 1992.325 ;
        RECT 2694.670 1992.140 2697.275 1992.280 ;
        RECT 2694.670 1992.080 2694.990 1992.140 ;
        RECT 2696.985 1992.095 2697.275 1992.140 ;
        RECT 2697.430 1991.260 2697.750 1991.320 ;
        RECT 2697.905 1991.260 2698.195 1991.305 ;
        RECT 2697.430 1991.120 2698.195 1991.260 ;
        RECT 2697.430 1991.060 2697.750 1991.120 ;
        RECT 2697.905 1991.075 2698.195 1991.120 ;
        RECT 2697.890 1986.640 2698.210 1986.900 ;
        RECT 2698.350 1986.640 2698.670 1986.900 ;
        RECT 2697.430 1986.300 2697.750 1986.560 ;
        RECT 2697.980 1986.500 2698.120 1986.640 ;
        RECT 2702.030 1986.500 2702.350 1986.560 ;
        RECT 2697.980 1986.360 2702.350 1986.500 ;
        RECT 2702.030 1986.300 2702.350 1986.360 ;
        RECT 2699.285 1985.820 2699.575 1985.865 ;
        RECT 2702.950 1985.820 2703.270 1985.880 ;
        RECT 2699.285 1985.680 2703.270 1985.820 ;
        RECT 2699.285 1985.635 2699.575 1985.680 ;
        RECT 2702.950 1985.620 2703.270 1985.680 ;
        RECT 2694.670 1983.780 2694.990 1983.840 ;
        RECT 2696.985 1983.780 2697.275 1983.825 ;
        RECT 2694.670 1983.640 2697.275 1983.780 ;
        RECT 2694.670 1983.580 2694.990 1983.640 ;
        RECT 2696.985 1983.595 2697.275 1983.640 ;
        RECT 2523.545 1982.750 2523.865 1983.010 ;
        RECT 2697.890 1982.900 2698.210 1983.160 ;
        RECT 2697.890 1982.080 2698.210 1982.140 ;
        RECT 2698.825 1982.080 2699.115 1982.125 ;
        RECT 2697.890 1981.940 2699.115 1982.080 ;
        RECT 2697.890 1981.880 2698.210 1981.940 ;
        RECT 2698.825 1981.895 2699.115 1981.940 ;
        RECT 2700.665 1982.080 2700.955 1982.125 ;
        RECT 2701.585 1982.080 2701.875 1982.125 ;
        RECT 2700.665 1981.940 2701.875 1982.080 ;
        RECT 2700.665 1981.895 2700.955 1981.940 ;
        RECT 2701.585 1981.895 2701.875 1981.940 ;
        RECT 2702.030 1981.880 2702.350 1982.140 ;
        RECT 2702.950 1981.880 2703.270 1982.140 ;
        RECT 2703.410 1981.880 2703.730 1982.140 ;
        RECT 2698.350 1981.740 2698.670 1981.800 ;
        RECT 2697.980 1981.600 2698.670 1981.740 ;
        RECT 2697.980 1981.105 2698.120 1981.600 ;
        RECT 2698.350 1981.540 2698.670 1981.600 ;
        RECT 2702.120 1981.445 2702.260 1981.880 ;
        RECT 2702.045 1981.215 2702.335 1981.445 ;
        RECT 2702.490 1981.200 2702.810 1981.460 ;
        RECT 2703.040 1981.445 2703.180 1981.880 ;
        RECT 2702.965 1981.215 2703.255 1981.445 ;
        RECT 2697.905 1980.875 2698.195 1981.105 ;
        RECT 2698.350 1980.860 2698.670 1981.120 ;
        RECT 2702.580 1981.060 2702.720 1981.200 ;
        RECT 2703.425 1981.060 2703.715 1981.105 ;
        RECT 2702.580 1980.920 2703.715 1981.060 ;
        RECT 2703.425 1980.875 2703.715 1980.920 ;
        RECT 2597.690 1980.400 2598.010 1980.460 ;
        RECT 2677.270 1980.400 2677.590 1980.460 ;
        RECT 2597.690 1980.260 2677.590 1980.400 ;
        RECT 2597.690 1980.200 2598.010 1980.260 ;
        RECT 2677.270 1980.200 2677.590 1980.260 ;
        RECT 2702.490 1980.180 2702.810 1980.440 ;
        RECT 2698.810 1979.160 2699.130 1979.420 ;
        RECT 2699.745 1979.360 2700.035 1979.405 ;
        RECT 2702.490 1979.360 2702.810 1979.420 ;
        RECT 2699.745 1979.220 2702.810 1979.360 ;
        RECT 2699.745 1979.175 2700.035 1979.220 ;
        RECT 2702.490 1979.160 2702.810 1979.220 ;
        RECT 2696.985 1979.020 2697.275 1979.065 ;
        RECT 2697.430 1979.020 2697.750 1979.080 ;
        RECT 2696.985 1978.880 2697.750 1979.020 ;
        RECT 2698.900 1979.020 2699.040 1979.160 ;
        RECT 2702.030 1979.020 2702.350 1979.080 ;
        RECT 2698.900 1978.880 2702.350 1979.020 ;
        RECT 2696.985 1978.835 2697.275 1978.880 ;
        RECT 2697.430 1978.820 2697.750 1978.880 ;
        RECT 2702.030 1978.820 2702.350 1978.880 ;
        RECT 2698.810 1977.460 2699.130 1977.720 ;
        RECT 2697.905 1976.640 2698.195 1976.685 ;
        RECT 2698.810 1976.640 2699.130 1976.700 ;
        RECT 2697.905 1976.500 2699.130 1976.640 ;
        RECT 2697.905 1976.455 2698.195 1976.500 ;
        RECT 2698.810 1976.440 2699.130 1976.500 ;
        RECT 2694.670 1975.960 2694.990 1976.020 ;
        RECT 2696.985 1975.960 2697.275 1976.005 ;
        RECT 2694.670 1975.820 2697.275 1975.960 ;
        RECT 2694.670 1975.760 2694.990 1975.820 ;
        RECT 2696.985 1975.775 2697.275 1975.820 ;
        RECT 2523.545 1975.220 2523.865 1975.480 ;
        RECT 2700.205 1973.240 2700.495 1973.285 ;
        RECT 2701.570 1973.240 2701.890 1973.300 ;
        RECT 2700.205 1973.100 2701.890 1973.240 ;
        RECT 2700.205 1973.055 2700.495 1973.100 ;
        RECT 2701.570 1973.040 2701.890 1973.100 ;
        RECT 2698.365 1972.900 2698.655 1972.945 ;
        RECT 2699.730 1972.900 2700.050 1972.960 ;
        RECT 2698.365 1972.760 2700.050 1972.900 ;
        RECT 2698.365 1972.715 2698.655 1972.760 ;
        RECT 2699.730 1972.700 2700.050 1972.760 ;
        RECT 2700.665 1972.900 2700.955 1972.945 ;
        RECT 2703.410 1972.900 2703.730 1972.960 ;
        RECT 2700.665 1972.760 2703.730 1972.900 ;
        RECT 2700.665 1972.715 2700.955 1972.760 ;
        RECT 2703.410 1972.700 2703.730 1972.760 ;
        RECT 2696.970 1972.560 2697.290 1972.620 ;
        RECT 2702.030 1972.560 2702.350 1972.620 ;
        RECT 2696.970 1972.420 2702.350 1972.560 ;
        RECT 2696.970 1972.360 2697.290 1972.420 ;
        RECT 2702.030 1972.360 2702.350 1972.420 ;
        RECT 2698.810 1972.020 2699.130 1972.280 ;
        RECT 2699.270 1972.020 2699.590 1972.280 ;
        RECT 2701.585 1972.220 2701.875 1972.265 ;
        RECT 2703.870 1972.220 2704.190 1972.280 ;
        RECT 2701.585 1972.080 2704.190 1972.220 ;
        RECT 2701.585 1972.035 2701.875 1972.080 ;
        RECT 2703.870 1972.020 2704.190 1972.080 ;
        RECT 2698.810 1971.200 2699.130 1971.260 ;
        RECT 2701.125 1971.200 2701.415 1971.245 ;
        RECT 2698.810 1971.060 2701.415 1971.200 ;
        RECT 2698.810 1971.000 2699.130 1971.060 ;
        RECT 2701.125 1971.015 2701.415 1971.060 ;
        RECT 2699.730 1970.860 2700.050 1970.920 ;
        RECT 2697.520 1970.720 2699.500 1970.860 ;
        RECT 2697.520 1970.580 2697.660 1970.720 ;
        RECT 2697.430 1970.320 2697.750 1970.580 ;
        RECT 2697.890 1970.320 2698.210 1970.580 ;
        RECT 2699.360 1970.225 2699.500 1970.720 ;
        RECT 2699.730 1970.720 2700.880 1970.860 ;
        RECT 2699.730 1970.660 2700.050 1970.720 ;
        RECT 2699.285 1969.995 2699.575 1970.225 ;
        RECT 2696.970 1969.500 2697.290 1969.560 ;
        RECT 2698.365 1969.500 2698.655 1969.545 ;
        RECT 2523.545 1969.240 2523.865 1969.500 ;
        RECT 2696.970 1969.360 2698.655 1969.500 ;
        RECT 2699.360 1969.500 2699.500 1969.995 ;
        RECT 2700.740 1969.885 2700.880 1970.720 ;
        RECT 2702.030 1970.320 2702.350 1970.580 ;
        RECT 2702.490 1970.320 2702.810 1970.580 ;
        RECT 2702.965 1970.335 2703.255 1970.565 ;
        RECT 2703.040 1970.180 2703.180 1970.335 ;
        RECT 2702.580 1970.040 2703.180 1970.180 ;
        RECT 2700.665 1969.655 2700.955 1969.885 ;
        RECT 2702.580 1969.500 2702.720 1970.040 ;
        RECT 2699.360 1969.360 2702.720 1969.500 ;
        RECT 2696.970 1969.300 2697.290 1969.360 ;
        RECT 2698.365 1969.315 2698.655 1969.360 ;
        RECT 2697.905 1968.480 2698.195 1968.525 ;
        RECT 2698.350 1968.480 2698.670 1968.540 ;
        RECT 2697.905 1968.340 2698.670 1968.480 ;
        RECT 2697.905 1968.295 2698.195 1968.340 ;
        RECT 2698.350 1968.280 2698.670 1968.340 ;
        RECT 2698.810 1968.480 2699.130 1968.540 ;
        RECT 2699.285 1968.480 2699.575 1968.525 ;
        RECT 2698.810 1968.340 2699.575 1968.480 ;
        RECT 2698.810 1968.280 2699.130 1968.340 ;
        RECT 2699.285 1968.295 2699.575 1968.340 ;
        RECT 2694.670 1967.460 2694.990 1967.520 ;
        RECT 2696.985 1967.460 2697.275 1967.505 ;
        RECT 2694.670 1967.320 2697.275 1967.460 ;
        RECT 2694.670 1967.260 2694.990 1967.320 ;
        RECT 2696.985 1967.275 2697.275 1967.320 ;
        RECT 2697.430 1967.460 2697.750 1967.520 ;
        RECT 2698.825 1967.460 2699.115 1967.505 ;
        RECT 2697.430 1967.320 2699.115 1967.460 ;
        RECT 2697.430 1967.260 2697.750 1967.320 ;
        RECT 2698.825 1967.275 2699.115 1967.320 ;
        RECT 2699.730 1967.260 2700.050 1967.520 ;
        RECT 2699.730 1965.760 2700.050 1965.820 ;
        RECT 2700.665 1965.760 2700.955 1965.805 ;
        RECT 2699.730 1965.620 2700.955 1965.760 ;
        RECT 2699.730 1965.560 2700.050 1965.620 ;
        RECT 2700.665 1965.575 2700.955 1965.620 ;
        RECT 2698.810 1964.880 2699.130 1965.140 ;
        RECT 2696.970 1964.740 2697.290 1964.800 ;
        RECT 2697.445 1964.740 2697.735 1964.785 ;
        RECT 2696.970 1964.600 2697.735 1964.740 ;
        RECT 2696.970 1964.540 2697.290 1964.600 ;
        RECT 2697.445 1964.555 2697.735 1964.600 ;
        RECT 2698.350 1964.540 2698.670 1964.800 ;
        RECT 2523.545 1963.295 2523.865 1963.555 ;
        RECT 2697.890 1962.840 2698.210 1963.100 ;
        RECT 2694.670 1962.020 2694.990 1962.080 ;
        RECT 2696.985 1962.020 2697.275 1962.065 ;
        RECT 2694.670 1961.880 2697.275 1962.020 ;
        RECT 2694.670 1961.820 2694.990 1961.880 ;
        RECT 2696.985 1961.835 2697.275 1961.880 ;
        RECT 2523.545 1957.650 2523.865 1957.910 ;
        RECT 2697.905 1957.600 2698.195 1957.645 ;
        RECT 2698.810 1957.600 2699.130 1957.660 ;
        RECT 2697.905 1957.460 2699.130 1957.600 ;
        RECT 2697.905 1957.415 2698.195 1957.460 ;
        RECT 2698.810 1957.400 2699.130 1957.460 ;
        RECT 2694.670 1956.580 2694.990 1956.640 ;
        RECT 2696.985 1956.580 2697.275 1956.625 ;
        RECT 2694.670 1956.440 2697.275 1956.580 ;
        RECT 2694.670 1956.380 2694.990 1956.440 ;
        RECT 2696.985 1956.395 2697.275 1956.440 ;
        RECT 2359.545 1953.060 2359.835 1953.290 ;
        RECT 2370.360 1953.060 2370.650 1953.290 ;
        RECT 2375.975 1953.060 2376.265 1953.290 ;
        RECT 2359.605 1952.610 2359.775 1953.060 ;
        RECT 2370.420 1952.715 2370.590 1953.060 ;
        RECT 2359.515 1952.320 2359.865 1952.610 ;
        RECT 2370.320 1952.345 2370.700 1952.715 ;
        RECT 2376.035 1952.580 2376.205 1953.060 ;
        RECT 2377.765 1953.025 2378.060 1953.285 ;
        RECT 2378.755 1953.025 2379.050 1953.285 ;
        RECT 2388.920 1953.060 2389.210 1953.290 ;
        RECT 2394.535 1953.060 2394.825 1953.290 ;
        RECT 2377.395 1952.655 2377.625 1952.685 ;
        RECT 2377.365 1952.580 2377.655 1952.655 ;
        RECT 2376.035 1952.550 2377.655 1952.580 ;
        RECT 2375.975 1952.410 2377.655 1952.550 ;
        RECT 2370.360 1952.320 2370.650 1952.345 ;
        RECT 2375.975 1952.320 2376.265 1952.410 ;
        RECT 2377.365 1952.350 2377.655 1952.410 ;
        RECT 2377.395 1952.335 2377.625 1952.350 ;
        RECT 2370.995 1952.180 2371.345 1952.245 ;
        RECT 2376.430 1952.180 2376.755 1952.270 ;
        RECT 2370.790 1952.150 2371.345 1952.180 ;
        RECT 2376.405 1952.150 2376.755 1952.180 ;
        RECT 2370.620 1952.145 2371.345 1952.150 ;
        RECT 2376.235 1952.145 2376.755 1952.150 ;
        RECT 2370.620 1951.975 2376.755 1952.145 ;
        RECT 2370.790 1951.950 2371.345 1951.975 ;
        RECT 2376.405 1951.950 2376.755 1951.975 ;
        RECT 2370.995 1951.895 2371.345 1951.950 ;
        RECT 2376.430 1951.945 2376.755 1951.950 ;
        RECT 2377.825 1951.925 2377.995 1953.025 ;
        RECT 2378.815 1952.295 2378.985 1953.025 ;
        RECT 2388.980 1952.715 2389.150 1953.060 ;
        RECT 2388.880 1952.345 2389.260 1952.715 ;
        RECT 2394.595 1952.580 2394.765 1953.060 ;
        RECT 2396.325 1953.025 2396.620 1953.285 ;
        RECT 2397.315 1953.025 2397.610 1953.285 ;
        RECT 2407.480 1953.060 2407.770 1953.290 ;
        RECT 2413.095 1953.060 2413.385 1953.290 ;
        RECT 2395.955 1952.655 2396.185 1952.685 ;
        RECT 2395.925 1952.580 2396.215 1952.655 ;
        RECT 2394.595 1952.550 2396.215 1952.580 ;
        RECT 2394.535 1952.410 2396.215 1952.550 ;
        RECT 2388.920 1952.320 2389.210 1952.345 ;
        RECT 2394.535 1952.320 2394.825 1952.410 ;
        RECT 2395.925 1952.350 2396.215 1952.410 ;
        RECT 2395.955 1952.335 2396.185 1952.350 ;
        RECT 2378.810 1951.945 2379.160 1952.295 ;
        RECT 2389.555 1952.180 2389.905 1952.250 ;
        RECT 2394.990 1952.180 2395.315 1952.270 ;
        RECT 2389.350 1952.150 2389.905 1952.180 ;
        RECT 2394.965 1952.150 2395.315 1952.180 ;
        RECT 2389.180 1952.145 2389.905 1952.150 ;
        RECT 2394.795 1952.145 2395.315 1952.150 ;
        RECT 2389.180 1951.975 2395.315 1952.145 ;
        RECT 2389.350 1951.950 2389.905 1951.975 ;
        RECT 2394.965 1951.950 2395.315 1951.975 ;
        RECT 2378.810 1951.925 2379.105 1951.945 ;
        RECT 2377.765 1951.920 2377.995 1951.925 ;
        RECT 2359.140 1951.790 2359.490 1951.865 ;
        RECT 2375.630 1951.820 2375.950 1951.835 ;
        RECT 2375.605 1951.790 2375.950 1951.820 ;
        RECT 2359.000 1951.620 2359.490 1951.790 ;
        RECT 2375.430 1951.620 2375.950 1951.790 ;
        RECT 2377.765 1951.685 2378.055 1951.920 ;
        RECT 2378.755 1951.855 2379.105 1951.925 ;
        RECT 2389.555 1951.900 2389.905 1951.950 ;
        RECT 2394.990 1951.945 2395.315 1951.950 ;
        RECT 2396.385 1951.925 2396.555 1953.025 ;
        RECT 2397.375 1952.305 2397.545 1953.025 ;
        RECT 2407.540 1952.715 2407.710 1953.060 ;
        RECT 2407.440 1952.345 2407.820 1952.715 ;
        RECT 2413.155 1952.580 2413.325 1953.060 ;
        RECT 2414.885 1953.025 2415.180 1953.285 ;
        RECT 2415.875 1953.025 2416.170 1953.285 ;
        RECT 2426.040 1953.060 2426.330 1953.290 ;
        RECT 2431.655 1953.060 2431.945 1953.290 ;
        RECT 2414.515 1952.655 2414.745 1952.685 ;
        RECT 2414.485 1952.580 2414.775 1952.655 ;
        RECT 2413.155 1952.550 2414.775 1952.580 ;
        RECT 2413.095 1952.410 2414.775 1952.550 ;
        RECT 2407.480 1952.320 2407.770 1952.345 ;
        RECT 2413.095 1952.320 2413.385 1952.410 ;
        RECT 2414.485 1952.350 2414.775 1952.410 ;
        RECT 2414.515 1952.335 2414.745 1952.350 ;
        RECT 2397.365 1951.950 2397.720 1952.305 ;
        RECT 2408.110 1952.180 2408.460 1952.255 ;
        RECT 2413.550 1952.180 2413.875 1952.270 ;
        RECT 2407.910 1952.150 2408.460 1952.180 ;
        RECT 2413.525 1952.150 2413.875 1952.180 ;
        RECT 2407.740 1952.145 2408.460 1952.150 ;
        RECT 2413.355 1952.145 2413.875 1952.150 ;
        RECT 2407.740 1951.975 2413.875 1952.145 ;
        RECT 2407.910 1951.950 2408.460 1951.975 ;
        RECT 2413.525 1951.950 2413.875 1951.975 ;
        RECT 2397.365 1951.925 2397.665 1951.950 ;
        RECT 2396.325 1951.920 2396.555 1951.925 ;
        RECT 2378.755 1951.685 2379.045 1951.855 ;
        RECT 2394.190 1951.820 2394.510 1951.835 ;
        RECT 2394.165 1951.790 2394.510 1951.820 ;
        RECT 2393.990 1951.620 2394.510 1951.790 ;
        RECT 2396.325 1951.685 2396.615 1951.920 ;
        RECT 2397.315 1951.855 2397.665 1951.925 ;
        RECT 2408.110 1951.905 2408.460 1951.950 ;
        RECT 2413.550 1951.945 2413.875 1951.950 ;
        RECT 2414.945 1951.925 2415.115 1953.025 ;
        RECT 2415.935 1952.295 2416.105 1953.025 ;
        RECT 2426.100 1952.715 2426.270 1953.060 ;
        RECT 2426.000 1952.345 2426.380 1952.715 ;
        RECT 2431.715 1952.580 2431.885 1953.060 ;
        RECT 2433.445 1953.025 2433.740 1953.285 ;
        RECT 2434.435 1953.025 2434.730 1953.285 ;
        RECT 2444.600 1953.060 2444.890 1953.290 ;
        RECT 2450.215 1953.060 2450.505 1953.290 ;
        RECT 2433.075 1952.655 2433.305 1952.685 ;
        RECT 2433.045 1952.580 2433.335 1952.655 ;
        RECT 2431.715 1952.550 2433.335 1952.580 ;
        RECT 2431.655 1952.410 2433.335 1952.550 ;
        RECT 2426.040 1952.320 2426.330 1952.345 ;
        RECT 2431.655 1952.320 2431.945 1952.410 ;
        RECT 2433.045 1952.350 2433.335 1952.410 ;
        RECT 2433.075 1952.335 2433.305 1952.350 ;
        RECT 2415.885 1951.945 2416.235 1952.295 ;
        RECT 2426.670 1952.180 2427.020 1952.250 ;
        RECT 2432.110 1952.180 2432.435 1952.270 ;
        RECT 2426.470 1952.150 2427.020 1952.180 ;
        RECT 2432.085 1952.150 2432.435 1952.180 ;
        RECT 2426.300 1952.145 2427.020 1952.150 ;
        RECT 2431.915 1952.145 2432.435 1952.150 ;
        RECT 2426.300 1951.975 2432.435 1952.145 ;
        RECT 2426.470 1951.950 2427.020 1951.975 ;
        RECT 2432.085 1951.950 2432.435 1951.975 ;
        RECT 2415.885 1951.925 2416.225 1951.945 ;
        RECT 2414.885 1951.920 2415.115 1951.925 ;
        RECT 2397.315 1951.685 2397.605 1951.855 ;
        RECT 2412.750 1951.820 2413.070 1951.835 ;
        RECT 2412.725 1951.790 2413.070 1951.820 ;
        RECT 2412.550 1951.620 2413.070 1951.790 ;
        RECT 2414.885 1951.685 2415.175 1951.920 ;
        RECT 2415.875 1951.855 2416.225 1951.925 ;
        RECT 2426.670 1951.900 2427.020 1951.950 ;
        RECT 2432.110 1951.945 2432.435 1951.950 ;
        RECT 2433.505 1951.925 2433.675 1953.025 ;
        RECT 2434.495 1952.295 2434.665 1953.025 ;
        RECT 2444.660 1952.715 2444.830 1953.060 ;
        RECT 2444.560 1952.345 2444.940 1952.715 ;
        RECT 2450.275 1952.580 2450.445 1953.060 ;
        RECT 2452.005 1953.025 2452.300 1953.285 ;
        RECT 2452.995 1953.025 2453.290 1953.285 ;
        RECT 2451.635 1952.655 2451.865 1952.685 ;
        RECT 2451.605 1952.580 2451.895 1952.655 ;
        RECT 2450.275 1952.550 2451.895 1952.580 ;
        RECT 2450.215 1952.410 2451.895 1952.550 ;
        RECT 2444.600 1952.320 2444.890 1952.345 ;
        RECT 2450.215 1952.320 2450.505 1952.410 ;
        RECT 2451.605 1952.350 2451.895 1952.410 ;
        RECT 2451.635 1952.335 2451.865 1952.350 ;
        RECT 2434.445 1951.945 2434.795 1952.295 ;
        RECT 2445.230 1952.180 2445.580 1952.250 ;
        RECT 2450.670 1952.180 2450.995 1952.270 ;
        RECT 2445.030 1952.150 2445.580 1952.180 ;
        RECT 2450.645 1952.150 2450.995 1952.180 ;
        RECT 2444.860 1952.145 2445.580 1952.150 ;
        RECT 2450.475 1952.145 2450.995 1952.150 ;
        RECT 2444.860 1951.975 2450.995 1952.145 ;
        RECT 2445.030 1951.950 2445.580 1951.975 ;
        RECT 2450.645 1951.950 2450.995 1951.975 ;
        RECT 2434.445 1951.925 2434.785 1951.945 ;
        RECT 2433.445 1951.920 2433.675 1951.925 ;
        RECT 2415.875 1951.685 2416.165 1951.855 ;
        RECT 2431.310 1951.820 2431.630 1951.835 ;
        RECT 2431.285 1951.790 2431.630 1951.820 ;
        RECT 2431.110 1951.620 2431.630 1951.790 ;
        RECT 2433.445 1951.685 2433.735 1951.920 ;
        RECT 2434.435 1951.855 2434.785 1951.925 ;
        RECT 2445.230 1951.900 2445.580 1951.950 ;
        RECT 2450.670 1951.945 2450.995 1951.950 ;
        RECT 2452.065 1951.925 2452.235 1953.025 ;
        RECT 2453.030 1953.000 2453.290 1953.025 ;
        RECT 2453.030 1952.915 2453.350 1953.000 ;
        RECT 2453.030 1952.565 2453.380 1952.915 ;
        RECT 2453.055 1951.925 2453.225 1952.565 ;
        RECT 2698.350 1952.160 2698.670 1952.220 ;
        RECT 2699.285 1952.160 2699.575 1952.205 ;
        RECT 2698.350 1952.020 2699.575 1952.160 ;
        RECT 2698.350 1951.960 2698.670 1952.020 ;
        RECT 2699.285 1951.975 2699.575 1952.020 ;
        RECT 2702.490 1951.960 2702.810 1952.220 ;
        RECT 2452.005 1951.920 2452.235 1951.925 ;
        RECT 2452.995 1951.920 2453.225 1951.925 ;
        RECT 2434.435 1951.685 2434.725 1951.855 ;
        RECT 2449.870 1951.820 2450.190 1951.835 ;
        RECT 2449.845 1951.790 2450.190 1951.820 ;
        RECT 2449.670 1951.620 2450.190 1951.790 ;
        RECT 2452.005 1951.685 2452.295 1951.920 ;
        RECT 2452.995 1951.685 2453.285 1951.920 ;
        RECT 2523.545 1951.645 2523.865 1951.905 ;
        RECT 2697.905 1951.820 2698.195 1951.865 ;
        RECT 2702.580 1951.820 2702.720 1951.960 ;
        RECT 2697.905 1951.680 2702.720 1951.820 ;
        RECT 2697.905 1951.635 2698.195 1951.680 ;
        RECT 2359.140 1951.575 2359.490 1951.620 ;
        RECT 2375.605 1951.590 2375.950 1951.620 ;
        RECT 2394.165 1951.590 2394.510 1951.620 ;
        RECT 2412.725 1951.590 2413.070 1951.620 ;
        RECT 2431.285 1951.590 2431.630 1951.620 ;
        RECT 2449.845 1951.590 2450.190 1951.620 ;
        RECT 2375.630 1951.545 2375.950 1951.590 ;
        RECT 2394.190 1951.545 2394.510 1951.590 ;
        RECT 2412.750 1951.545 2413.070 1951.590 ;
        RECT 2431.310 1951.545 2431.630 1951.590 ;
        RECT 2449.870 1951.545 2450.190 1951.590 ;
        RECT 2694.670 1951.140 2694.990 1951.200 ;
        RECT 2696.985 1951.140 2697.275 1951.185 ;
        RECT 2694.670 1951.000 2697.275 1951.140 ;
        RECT 2694.670 1950.940 2694.990 1951.000 ;
        RECT 2696.985 1950.955 2697.275 1951.000 ;
        RECT 2698.350 1950.940 2698.670 1951.200 ;
        RECT 2366.555 1948.065 2366.875 1948.125 ;
        RECT 2361.795 1947.555 2362.115 1947.965 ;
        RECT 2366.555 1947.925 2367.625 1948.065 ;
        RECT 2364.805 1947.825 2365.905 1947.895 ;
        RECT 2366.555 1947.865 2366.875 1947.925 ;
        RECT 2364.735 1947.755 2365.985 1947.825 ;
        RECT 2364.735 1947.595 2365.025 1947.755 ;
        RECT 2365.695 1947.595 2365.985 1947.755 ;
        RECT 2361.875 1946.425 2362.035 1947.555 ;
        RECT 2362.755 1947.305 2363.075 1947.565 ;
        RECT 2363.875 1947.445 2364.195 1947.565 ;
        RECT 2365.215 1947.505 2365.505 1947.545 ;
        RECT 2363.875 1947.305 2364.705 1947.445 ;
        RECT 2365.215 1947.315 2365.545 1947.505 ;
        RECT 2364.495 1947.265 2364.705 1947.305 ;
        RECT 2364.495 1947.035 2364.785 1947.265 ;
        RECT 2362.275 1946.985 2362.595 1947.005 ;
        RECT 2362.275 1946.845 2363.225 1946.985 ;
        RECT 2363.685 1946.945 2363.975 1946.985 ;
        RECT 2362.275 1946.755 2362.825 1946.845 ;
        RECT 2363.085 1946.805 2363.225 1946.845 ;
        RECT 2363.585 1946.805 2363.975 1946.945 ;
        RECT 2363.085 1946.755 2363.975 1946.805 ;
        RECT 2362.275 1946.745 2362.595 1946.755 ;
        RECT 2363.085 1946.665 2363.725 1946.755 ;
        RECT 2361.815 1946.195 2362.105 1946.425 ;
        RECT 2362.755 1946.385 2363.075 1946.445 ;
        RECT 2364.715 1946.385 2365.035 1946.445 ;
        RECT 2365.405 1946.425 2365.545 1947.315 ;
        RECT 2366.195 1947.305 2366.515 1947.565 ;
        RECT 2366.915 1947.305 2367.235 1947.565 ;
        RECT 2367.485 1947.505 2367.625 1947.925 ;
        RECT 2368.115 1947.865 2368.435 1948.125 ;
        RECT 2368.655 1948.065 2368.945 1948.105 ;
        RECT 2369.115 1948.065 2369.435 1948.125 ;
        RECT 2368.655 1947.925 2369.435 1948.065 ;
        RECT 2368.655 1947.875 2368.945 1947.925 ;
        RECT 2369.115 1947.865 2369.435 1947.925 ;
        RECT 2369.595 1947.865 2369.915 1948.125 ;
        RECT 2370.075 1947.865 2370.395 1948.125 ;
        RECT 2371.075 1947.895 2371.395 1948.125 ;
        RECT 2385.115 1948.065 2385.435 1948.125 ;
        RECT 2371.075 1947.865 2372.505 1947.895 ;
        RECT 2371.165 1947.755 2372.505 1947.865 ;
        RECT 2368.655 1947.505 2368.945 1947.545 ;
        RECT 2367.485 1947.365 2368.945 1947.505 ;
        RECT 2368.655 1947.315 2368.945 1947.365 ;
        RECT 2370.595 1947.305 2370.915 1947.565 ;
        RECT 2371.165 1947.545 2371.305 1947.755 ;
        RECT 2371.095 1947.315 2371.385 1947.545 ;
        RECT 2371.815 1947.505 2372.105 1947.545 ;
        RECT 2371.815 1947.315 2372.145 1947.505 ;
        RECT 2370.095 1947.225 2370.385 1947.265 ;
        RECT 2370.595 1947.225 2370.825 1947.305 ;
        RECT 2370.095 1947.085 2370.825 1947.225 ;
        RECT 2370.095 1947.035 2370.385 1947.085 ;
        RECT 2365.935 1946.985 2366.255 1947.005 ;
        RECT 2365.695 1946.945 2366.255 1946.985 ;
        RECT 2366.935 1946.945 2367.225 1946.985 ;
        RECT 2365.695 1946.805 2367.225 1946.945 ;
        RECT 2365.695 1946.755 2366.255 1946.805 ;
        RECT 2366.935 1946.755 2367.225 1946.805 ;
        RECT 2367.415 1946.945 2367.705 1946.985 ;
        RECT 2367.415 1946.805 2368.345 1946.945 ;
        RECT 2367.415 1946.755 2367.705 1946.805 ;
        RECT 2365.935 1946.745 2366.255 1946.755 ;
        RECT 2362.755 1946.245 2365.035 1946.385 ;
        RECT 2362.755 1946.185 2363.075 1946.245 ;
        RECT 2364.715 1946.185 2365.035 1946.245 ;
        RECT 2365.215 1946.385 2365.545 1946.425 ;
        RECT 2366.195 1946.385 2366.515 1946.445 ;
        RECT 2366.915 1946.425 2367.235 1946.445 ;
        RECT 2365.215 1946.245 2366.515 1946.385 ;
        RECT 2365.215 1946.195 2365.505 1946.245 ;
        RECT 2366.195 1946.185 2366.515 1946.245 ;
        RECT 2366.695 1946.195 2367.235 1946.425 ;
        RECT 2366.915 1946.185 2367.235 1946.195 ;
        RECT 2367.635 1946.185 2367.955 1946.445 ;
        RECT 2368.205 1946.385 2368.345 1946.805 ;
        RECT 2368.635 1946.805 2368.955 1947.005 ;
        RECT 2371.335 1946.805 2371.625 1946.985 ;
        RECT 2368.635 1946.755 2371.625 1946.805 ;
        RECT 2368.635 1946.745 2371.545 1946.755 ;
        RECT 2368.725 1946.665 2371.545 1946.745 ;
        RECT 2372.005 1946.445 2372.145 1947.315 ;
        RECT 2372.365 1947.265 2372.505 1947.755 ;
        RECT 2374.025 1947.445 2374.365 1947.795 ;
        RECT 2380.355 1947.555 2380.675 1947.965 ;
        RECT 2385.115 1947.925 2386.185 1948.065 ;
        RECT 2383.365 1947.825 2384.465 1947.895 ;
        RECT 2385.115 1947.865 2385.435 1947.925 ;
        RECT 2383.295 1947.755 2384.545 1947.825 ;
        RECT 2383.295 1947.595 2383.585 1947.755 ;
        RECT 2384.255 1947.595 2384.545 1947.755 ;
        RECT 2372.295 1947.035 2372.585 1947.265 ;
        RECT 2374.115 1946.490 2374.285 1947.445 ;
        RECT 2375.630 1946.875 2375.950 1946.980 ;
        RECT 2375.605 1946.860 2375.950 1946.875 ;
        RECT 2375.600 1946.845 2375.950 1946.860 ;
        RECT 2375.430 1946.675 2375.950 1946.845 ;
        RECT 2375.605 1946.660 2375.950 1946.675 ;
        RECT 2375.605 1946.645 2375.895 1946.660 ;
        RECT 2376.405 1946.490 2376.755 1946.610 ;
        RECT 2377.765 1946.545 2378.055 1946.780 ;
        RECT 2378.750 1946.545 2379.040 1946.780 ;
        RECT 2377.765 1946.540 2377.995 1946.545 ;
        RECT 2378.750 1946.540 2378.980 1946.545 ;
        RECT 2368.875 1946.425 2369.195 1946.445 ;
        RECT 2368.655 1946.385 2369.195 1946.425 ;
        RECT 2368.205 1946.245 2369.195 1946.385 ;
        RECT 2368.655 1946.195 2369.195 1946.245 ;
        RECT 2368.875 1946.185 2369.195 1946.195 ;
        RECT 2369.475 1946.185 2370.155 1946.445 ;
        RECT 2370.595 1946.385 2370.915 1946.445 ;
        RECT 2371.095 1946.385 2371.385 1946.425 ;
        RECT 2370.595 1946.245 2371.385 1946.385 ;
        RECT 2372.005 1946.245 2372.355 1946.445 ;
        RECT 2374.115 1946.320 2376.755 1946.490 ;
        RECT 2376.235 1946.315 2376.755 1946.320 ;
        RECT 2376.405 1946.260 2376.755 1946.315 ;
        RECT 2370.595 1946.185 2370.915 1946.245 ;
        RECT 2371.095 1946.195 2371.385 1946.245 ;
        RECT 2372.035 1946.185 2372.355 1946.245 ;
        RECT 2377.400 1946.225 2377.630 1946.245 ;
        RECT 2375.975 1946.120 2376.265 1946.145 ;
        RECT 2377.370 1946.120 2377.660 1946.225 ;
        RECT 2375.975 1945.950 2377.660 1946.120 ;
        RECT 2375.975 1945.915 2376.265 1945.950 ;
        RECT 2377.370 1945.915 2377.660 1945.950 ;
        RECT 2376.035 1945.405 2376.205 1945.915 ;
        RECT 2377.400 1945.895 2377.630 1945.915 ;
        RECT 2377.825 1945.440 2377.995 1946.540 ;
        RECT 2378.810 1945.440 2378.980 1946.540 ;
        RECT 2380.435 1946.425 2380.595 1947.555 ;
        RECT 2381.315 1947.305 2381.635 1947.565 ;
        RECT 2382.435 1947.445 2382.755 1947.565 ;
        RECT 2383.775 1947.505 2384.065 1947.545 ;
        RECT 2382.435 1947.305 2383.265 1947.445 ;
        RECT 2383.775 1947.315 2384.105 1947.505 ;
        RECT 2383.055 1947.265 2383.265 1947.305 ;
        RECT 2383.055 1947.035 2383.345 1947.265 ;
        RECT 2380.835 1946.985 2381.155 1947.005 ;
        RECT 2380.835 1946.845 2381.785 1946.985 ;
        RECT 2382.245 1946.945 2382.535 1946.985 ;
        RECT 2380.835 1946.755 2381.385 1946.845 ;
        RECT 2381.645 1946.805 2381.785 1946.845 ;
        RECT 2382.145 1946.805 2382.535 1946.945 ;
        RECT 2381.645 1946.755 2382.535 1946.805 ;
        RECT 2380.835 1946.745 2381.155 1946.755 ;
        RECT 2381.645 1946.665 2382.285 1946.755 ;
        RECT 2380.375 1946.195 2380.665 1946.425 ;
        RECT 2381.315 1946.385 2381.635 1946.445 ;
        RECT 2383.275 1946.385 2383.595 1946.445 ;
        RECT 2383.965 1946.425 2384.105 1947.315 ;
        RECT 2384.755 1947.305 2385.075 1947.565 ;
        RECT 2385.475 1947.305 2385.795 1947.565 ;
        RECT 2386.045 1947.505 2386.185 1947.925 ;
        RECT 2386.675 1947.865 2386.995 1948.125 ;
        RECT 2387.215 1948.065 2387.505 1948.105 ;
        RECT 2387.675 1948.065 2387.995 1948.125 ;
        RECT 2387.215 1947.925 2387.995 1948.065 ;
        RECT 2387.215 1947.875 2387.505 1947.925 ;
        RECT 2387.675 1947.865 2387.995 1947.925 ;
        RECT 2388.155 1947.865 2388.475 1948.125 ;
        RECT 2388.635 1947.865 2388.955 1948.125 ;
        RECT 2389.635 1947.895 2389.955 1948.125 ;
        RECT 2403.675 1948.065 2403.995 1948.125 ;
        RECT 2389.635 1947.865 2391.065 1947.895 ;
        RECT 2389.725 1947.755 2391.065 1947.865 ;
        RECT 2387.215 1947.505 2387.505 1947.545 ;
        RECT 2386.045 1947.365 2387.505 1947.505 ;
        RECT 2387.215 1947.315 2387.505 1947.365 ;
        RECT 2389.155 1947.305 2389.475 1947.565 ;
        RECT 2389.725 1947.545 2389.865 1947.755 ;
        RECT 2389.655 1947.315 2389.945 1947.545 ;
        RECT 2390.375 1947.505 2390.665 1947.545 ;
        RECT 2390.375 1947.315 2390.705 1947.505 ;
        RECT 2388.655 1947.225 2388.945 1947.265 ;
        RECT 2389.155 1947.225 2389.385 1947.305 ;
        RECT 2388.655 1947.085 2389.385 1947.225 ;
        RECT 2388.655 1947.035 2388.945 1947.085 ;
        RECT 2384.495 1946.985 2384.815 1947.005 ;
        RECT 2384.255 1946.945 2384.815 1946.985 ;
        RECT 2385.495 1946.945 2385.785 1946.985 ;
        RECT 2384.255 1946.805 2385.785 1946.945 ;
        RECT 2384.255 1946.755 2384.815 1946.805 ;
        RECT 2385.495 1946.755 2385.785 1946.805 ;
        RECT 2385.975 1946.945 2386.265 1946.985 ;
        RECT 2385.975 1946.805 2386.905 1946.945 ;
        RECT 2385.975 1946.755 2386.265 1946.805 ;
        RECT 2384.495 1946.745 2384.815 1946.755 ;
        RECT 2381.315 1946.245 2383.595 1946.385 ;
        RECT 2381.315 1946.185 2381.635 1946.245 ;
        RECT 2383.275 1946.185 2383.595 1946.245 ;
        RECT 2383.775 1946.385 2384.105 1946.425 ;
        RECT 2384.755 1946.385 2385.075 1946.445 ;
        RECT 2385.475 1946.425 2385.795 1946.445 ;
        RECT 2383.775 1946.245 2385.075 1946.385 ;
        RECT 2383.775 1946.195 2384.065 1946.245 ;
        RECT 2384.755 1946.185 2385.075 1946.245 ;
        RECT 2385.255 1946.195 2385.795 1946.425 ;
        RECT 2385.475 1946.185 2385.795 1946.195 ;
        RECT 2386.195 1946.185 2386.515 1946.445 ;
        RECT 2386.765 1946.385 2386.905 1946.805 ;
        RECT 2387.195 1946.805 2387.515 1947.005 ;
        RECT 2389.895 1946.805 2390.185 1946.985 ;
        RECT 2387.195 1946.755 2390.185 1946.805 ;
        RECT 2387.195 1946.745 2390.105 1946.755 ;
        RECT 2387.285 1946.665 2390.105 1946.745 ;
        RECT 2390.565 1946.445 2390.705 1947.315 ;
        RECT 2390.925 1947.265 2391.065 1947.755 ;
        RECT 2392.585 1947.445 2392.925 1947.795 ;
        RECT 2398.915 1947.555 2399.235 1947.965 ;
        RECT 2403.675 1947.925 2404.745 1948.065 ;
        RECT 2401.925 1947.825 2403.025 1947.895 ;
        RECT 2403.675 1947.865 2403.995 1947.925 ;
        RECT 2401.855 1947.755 2403.105 1947.825 ;
        RECT 2401.855 1947.595 2402.145 1947.755 ;
        RECT 2402.815 1947.595 2403.105 1947.755 ;
        RECT 2397.130 1947.465 2397.450 1947.480 ;
        RECT 2390.855 1947.035 2391.145 1947.265 ;
        RECT 2392.675 1946.490 2392.845 1947.445 ;
        RECT 2397.130 1947.235 2397.600 1947.465 ;
        RECT 2397.130 1947.220 2397.450 1947.235 ;
        RECT 2394.190 1946.875 2394.510 1946.980 ;
        RECT 2394.165 1946.860 2394.510 1946.875 ;
        RECT 2394.160 1946.845 2394.510 1946.860 ;
        RECT 2393.990 1946.675 2394.510 1946.845 ;
        RECT 2394.165 1946.660 2394.510 1946.675 ;
        RECT 2394.165 1946.645 2394.455 1946.660 ;
        RECT 2394.965 1946.490 2395.315 1946.610 ;
        RECT 2396.325 1946.545 2396.615 1946.780 ;
        RECT 2397.310 1946.545 2397.600 1946.780 ;
        RECT 2396.325 1946.540 2396.555 1946.545 ;
        RECT 2397.310 1946.540 2397.540 1946.545 ;
        RECT 2387.435 1946.425 2387.755 1946.445 ;
        RECT 2387.215 1946.385 2387.755 1946.425 ;
        RECT 2386.765 1946.245 2387.755 1946.385 ;
        RECT 2387.215 1946.195 2387.755 1946.245 ;
        RECT 2387.435 1946.185 2387.755 1946.195 ;
        RECT 2388.035 1946.185 2388.715 1946.445 ;
        RECT 2389.155 1946.385 2389.475 1946.445 ;
        RECT 2389.655 1946.385 2389.945 1946.425 ;
        RECT 2389.155 1946.245 2389.945 1946.385 ;
        RECT 2390.565 1946.245 2390.915 1946.445 ;
        RECT 2392.675 1946.320 2395.315 1946.490 ;
        RECT 2394.795 1946.315 2395.315 1946.320 ;
        RECT 2394.965 1946.260 2395.315 1946.315 ;
        RECT 2389.155 1946.185 2389.475 1946.245 ;
        RECT 2389.655 1946.195 2389.945 1946.245 ;
        RECT 2390.595 1946.185 2390.915 1946.245 ;
        RECT 2395.960 1946.225 2396.190 1946.245 ;
        RECT 2394.535 1946.120 2394.825 1946.145 ;
        RECT 2395.930 1946.120 2396.220 1946.225 ;
        RECT 2394.535 1945.950 2396.220 1946.120 ;
        RECT 2394.535 1945.915 2394.825 1945.950 ;
        RECT 2395.930 1945.915 2396.220 1945.950 ;
        RECT 2375.975 1945.175 2376.265 1945.405 ;
        RECT 2377.765 1945.180 2378.060 1945.440 ;
        RECT 2378.730 1945.180 2379.050 1945.440 ;
        RECT 2394.595 1945.405 2394.765 1945.915 ;
        RECT 2395.960 1945.895 2396.190 1945.915 ;
        RECT 2396.385 1945.440 2396.555 1946.540 ;
        RECT 2397.370 1945.440 2397.540 1946.540 ;
        RECT 2398.995 1946.425 2399.155 1947.555 ;
        RECT 2399.875 1947.305 2400.195 1947.565 ;
        RECT 2400.995 1947.445 2401.315 1947.565 ;
        RECT 2402.335 1947.505 2402.625 1947.545 ;
        RECT 2400.995 1947.305 2401.825 1947.445 ;
        RECT 2402.335 1947.315 2402.665 1947.505 ;
        RECT 2401.615 1947.265 2401.825 1947.305 ;
        RECT 2401.615 1947.035 2401.905 1947.265 ;
        RECT 2399.395 1946.985 2399.715 1947.005 ;
        RECT 2399.395 1946.845 2400.345 1946.985 ;
        RECT 2400.805 1946.945 2401.095 1946.985 ;
        RECT 2399.395 1946.755 2399.945 1946.845 ;
        RECT 2400.205 1946.805 2400.345 1946.845 ;
        RECT 2400.705 1946.805 2401.095 1946.945 ;
        RECT 2400.205 1946.755 2401.095 1946.805 ;
        RECT 2399.395 1946.745 2399.715 1946.755 ;
        RECT 2400.205 1946.665 2400.845 1946.755 ;
        RECT 2398.935 1946.195 2399.225 1946.425 ;
        RECT 2399.875 1946.385 2400.195 1946.445 ;
        RECT 2401.835 1946.385 2402.155 1946.445 ;
        RECT 2402.525 1946.425 2402.665 1947.315 ;
        RECT 2403.315 1947.305 2403.635 1947.565 ;
        RECT 2404.035 1947.305 2404.355 1947.565 ;
        RECT 2404.605 1947.505 2404.745 1947.925 ;
        RECT 2405.235 1947.865 2405.555 1948.125 ;
        RECT 2405.775 1948.065 2406.065 1948.105 ;
        RECT 2406.235 1948.065 2406.555 1948.125 ;
        RECT 2405.775 1947.925 2406.555 1948.065 ;
        RECT 2405.775 1947.875 2406.065 1947.925 ;
        RECT 2406.235 1947.865 2406.555 1947.925 ;
        RECT 2406.715 1947.865 2407.035 1948.125 ;
        RECT 2407.195 1947.865 2407.515 1948.125 ;
        RECT 2408.195 1947.895 2408.515 1948.125 ;
        RECT 2422.235 1948.065 2422.555 1948.125 ;
        RECT 2408.195 1947.865 2409.625 1947.895 ;
        RECT 2408.285 1947.755 2409.625 1947.865 ;
        RECT 2405.775 1947.505 2406.065 1947.545 ;
        RECT 2404.605 1947.365 2406.065 1947.505 ;
        RECT 2405.775 1947.315 2406.065 1947.365 ;
        RECT 2407.715 1947.305 2408.035 1947.565 ;
        RECT 2408.285 1947.545 2408.425 1947.755 ;
        RECT 2408.215 1947.315 2408.505 1947.545 ;
        RECT 2408.935 1947.505 2409.225 1947.545 ;
        RECT 2408.935 1947.315 2409.265 1947.505 ;
        RECT 2407.215 1947.225 2407.505 1947.265 ;
        RECT 2407.715 1947.225 2407.945 1947.305 ;
        RECT 2407.215 1947.085 2407.945 1947.225 ;
        RECT 2407.215 1947.035 2407.505 1947.085 ;
        RECT 2403.055 1946.985 2403.375 1947.005 ;
        RECT 2402.815 1946.945 2403.375 1946.985 ;
        RECT 2404.055 1946.945 2404.345 1946.985 ;
        RECT 2402.815 1946.805 2404.345 1946.945 ;
        RECT 2402.815 1946.755 2403.375 1946.805 ;
        RECT 2404.055 1946.755 2404.345 1946.805 ;
        RECT 2404.535 1946.945 2404.825 1946.985 ;
        RECT 2404.535 1946.805 2405.465 1946.945 ;
        RECT 2404.535 1946.755 2404.825 1946.805 ;
        RECT 2403.055 1946.745 2403.375 1946.755 ;
        RECT 2399.875 1946.245 2402.155 1946.385 ;
        RECT 2399.875 1946.185 2400.195 1946.245 ;
        RECT 2401.835 1946.185 2402.155 1946.245 ;
        RECT 2402.335 1946.385 2402.665 1946.425 ;
        RECT 2403.315 1946.385 2403.635 1946.445 ;
        RECT 2404.035 1946.425 2404.355 1946.445 ;
        RECT 2402.335 1946.245 2403.635 1946.385 ;
        RECT 2402.335 1946.195 2402.625 1946.245 ;
        RECT 2403.315 1946.185 2403.635 1946.245 ;
        RECT 2403.815 1946.195 2404.355 1946.425 ;
        RECT 2404.035 1946.185 2404.355 1946.195 ;
        RECT 2404.755 1946.185 2405.075 1946.445 ;
        RECT 2405.325 1946.385 2405.465 1946.805 ;
        RECT 2405.755 1946.805 2406.075 1947.005 ;
        RECT 2408.455 1946.805 2408.745 1946.985 ;
        RECT 2405.755 1946.755 2408.745 1946.805 ;
        RECT 2405.755 1946.745 2408.665 1946.755 ;
        RECT 2405.845 1946.665 2408.665 1946.745 ;
        RECT 2409.125 1946.445 2409.265 1947.315 ;
        RECT 2409.485 1947.265 2409.625 1947.755 ;
        RECT 2411.145 1947.445 2411.485 1947.795 ;
        RECT 2417.475 1947.555 2417.795 1947.965 ;
        RECT 2422.235 1947.925 2423.305 1948.065 ;
        RECT 2420.485 1947.825 2421.585 1947.895 ;
        RECT 2422.235 1947.865 2422.555 1947.925 ;
        RECT 2420.415 1947.755 2421.665 1947.825 ;
        RECT 2420.415 1947.595 2420.705 1947.755 ;
        RECT 2421.375 1947.595 2421.665 1947.755 ;
        RECT 2409.415 1947.035 2409.705 1947.265 ;
        RECT 2411.235 1946.490 2411.405 1947.445 ;
        RECT 2412.750 1946.875 2413.070 1946.980 ;
        RECT 2412.725 1946.860 2413.070 1946.875 ;
        RECT 2412.720 1946.845 2413.070 1946.860 ;
        RECT 2412.550 1946.675 2413.070 1946.845 ;
        RECT 2412.725 1946.660 2413.070 1946.675 ;
        RECT 2412.725 1946.645 2413.015 1946.660 ;
        RECT 2413.525 1946.490 2413.875 1946.610 ;
        RECT 2414.885 1946.545 2415.175 1946.780 ;
        RECT 2415.870 1946.545 2416.160 1946.780 ;
        RECT 2414.885 1946.540 2415.115 1946.545 ;
        RECT 2415.870 1946.540 2416.100 1946.545 ;
        RECT 2405.995 1946.425 2406.315 1946.445 ;
        RECT 2405.775 1946.385 2406.315 1946.425 ;
        RECT 2405.325 1946.245 2406.315 1946.385 ;
        RECT 2405.775 1946.195 2406.315 1946.245 ;
        RECT 2405.995 1946.185 2406.315 1946.195 ;
        RECT 2406.595 1946.185 2407.275 1946.445 ;
        RECT 2407.715 1946.385 2408.035 1946.445 ;
        RECT 2408.215 1946.385 2408.505 1946.425 ;
        RECT 2407.715 1946.245 2408.505 1946.385 ;
        RECT 2409.125 1946.245 2409.475 1946.445 ;
        RECT 2411.235 1946.320 2413.875 1946.490 ;
        RECT 2413.355 1946.315 2413.875 1946.320 ;
        RECT 2413.525 1946.260 2413.875 1946.315 ;
        RECT 2407.715 1946.185 2408.035 1946.245 ;
        RECT 2408.215 1946.195 2408.505 1946.245 ;
        RECT 2409.155 1946.185 2409.475 1946.245 ;
        RECT 2414.520 1946.225 2414.750 1946.245 ;
        RECT 2413.095 1946.120 2413.385 1946.145 ;
        RECT 2414.490 1946.120 2414.780 1946.225 ;
        RECT 2413.095 1945.950 2414.780 1946.120 ;
        RECT 2413.095 1945.915 2413.385 1945.950 ;
        RECT 2414.490 1945.915 2414.780 1945.950 ;
        RECT 2394.535 1945.175 2394.825 1945.405 ;
        RECT 2396.325 1945.180 2396.620 1945.440 ;
        RECT 2397.310 1945.180 2397.605 1945.440 ;
        RECT 2413.155 1945.405 2413.325 1945.915 ;
        RECT 2414.520 1945.895 2414.750 1945.915 ;
        RECT 2414.945 1945.440 2415.115 1946.540 ;
        RECT 2415.930 1945.440 2416.100 1946.540 ;
        RECT 2417.555 1946.425 2417.715 1947.555 ;
        RECT 2418.435 1947.305 2418.755 1947.565 ;
        RECT 2419.555 1947.445 2419.875 1947.565 ;
        RECT 2420.895 1947.505 2421.185 1947.545 ;
        RECT 2419.555 1947.305 2420.385 1947.445 ;
        RECT 2420.895 1947.315 2421.225 1947.505 ;
        RECT 2420.175 1947.265 2420.385 1947.305 ;
        RECT 2420.175 1947.035 2420.465 1947.265 ;
        RECT 2417.955 1946.985 2418.275 1947.005 ;
        RECT 2417.955 1946.845 2418.905 1946.985 ;
        RECT 2419.365 1946.945 2419.655 1946.985 ;
        RECT 2417.955 1946.755 2418.505 1946.845 ;
        RECT 2418.765 1946.805 2418.905 1946.845 ;
        RECT 2419.265 1946.805 2419.655 1946.945 ;
        RECT 2418.765 1946.755 2419.655 1946.805 ;
        RECT 2417.955 1946.745 2418.275 1946.755 ;
        RECT 2418.765 1946.665 2419.405 1946.755 ;
        RECT 2417.495 1946.195 2417.785 1946.425 ;
        RECT 2418.435 1946.385 2418.755 1946.445 ;
        RECT 2420.395 1946.385 2420.715 1946.445 ;
        RECT 2421.085 1946.425 2421.225 1947.315 ;
        RECT 2421.875 1947.305 2422.195 1947.565 ;
        RECT 2422.595 1947.305 2422.915 1947.565 ;
        RECT 2423.165 1947.505 2423.305 1947.925 ;
        RECT 2423.795 1947.865 2424.115 1948.125 ;
        RECT 2424.335 1948.065 2424.625 1948.105 ;
        RECT 2424.795 1948.065 2425.115 1948.125 ;
        RECT 2424.335 1947.925 2425.115 1948.065 ;
        RECT 2424.335 1947.875 2424.625 1947.925 ;
        RECT 2424.795 1947.865 2425.115 1947.925 ;
        RECT 2425.275 1947.865 2425.595 1948.125 ;
        RECT 2425.755 1947.865 2426.075 1948.125 ;
        RECT 2426.755 1947.895 2427.075 1948.125 ;
        RECT 2440.795 1948.065 2441.115 1948.125 ;
        RECT 2426.755 1947.865 2428.185 1947.895 ;
        RECT 2426.845 1947.755 2428.185 1947.865 ;
        RECT 2424.335 1947.505 2424.625 1947.545 ;
        RECT 2423.165 1947.365 2424.625 1947.505 ;
        RECT 2424.335 1947.315 2424.625 1947.365 ;
        RECT 2426.275 1947.305 2426.595 1947.565 ;
        RECT 2426.845 1947.545 2426.985 1947.755 ;
        RECT 2426.775 1947.315 2427.065 1947.545 ;
        RECT 2427.495 1947.505 2427.785 1947.545 ;
        RECT 2427.495 1947.315 2427.825 1947.505 ;
        RECT 2425.775 1947.225 2426.065 1947.265 ;
        RECT 2426.275 1947.225 2426.505 1947.305 ;
        RECT 2425.775 1947.085 2426.505 1947.225 ;
        RECT 2425.775 1947.035 2426.065 1947.085 ;
        RECT 2421.615 1946.985 2421.935 1947.005 ;
        RECT 2421.375 1946.945 2421.935 1946.985 ;
        RECT 2422.615 1946.945 2422.905 1946.985 ;
        RECT 2421.375 1946.805 2422.905 1946.945 ;
        RECT 2421.375 1946.755 2421.935 1946.805 ;
        RECT 2422.615 1946.755 2422.905 1946.805 ;
        RECT 2423.095 1946.945 2423.385 1946.985 ;
        RECT 2423.095 1946.805 2424.025 1946.945 ;
        RECT 2423.095 1946.755 2423.385 1946.805 ;
        RECT 2421.615 1946.745 2421.935 1946.755 ;
        RECT 2418.435 1946.245 2420.715 1946.385 ;
        RECT 2418.435 1946.185 2418.755 1946.245 ;
        RECT 2420.395 1946.185 2420.715 1946.245 ;
        RECT 2420.895 1946.385 2421.225 1946.425 ;
        RECT 2421.875 1946.385 2422.195 1946.445 ;
        RECT 2422.595 1946.425 2422.915 1946.445 ;
        RECT 2420.895 1946.245 2422.195 1946.385 ;
        RECT 2420.895 1946.195 2421.185 1946.245 ;
        RECT 2421.875 1946.185 2422.195 1946.245 ;
        RECT 2422.375 1946.195 2422.915 1946.425 ;
        RECT 2422.595 1946.185 2422.915 1946.195 ;
        RECT 2423.315 1946.185 2423.635 1946.445 ;
        RECT 2423.885 1946.385 2424.025 1946.805 ;
        RECT 2424.315 1946.805 2424.635 1947.005 ;
        RECT 2427.015 1946.805 2427.305 1946.985 ;
        RECT 2424.315 1946.755 2427.305 1946.805 ;
        RECT 2424.315 1946.745 2427.225 1946.755 ;
        RECT 2424.405 1946.665 2427.225 1946.745 ;
        RECT 2427.685 1946.445 2427.825 1947.315 ;
        RECT 2428.045 1947.265 2428.185 1947.755 ;
        RECT 2429.705 1947.445 2430.045 1947.795 ;
        RECT 2436.035 1947.555 2436.355 1947.965 ;
        RECT 2440.795 1947.925 2441.865 1948.065 ;
        RECT 2439.045 1947.825 2440.145 1947.895 ;
        RECT 2440.795 1947.865 2441.115 1947.925 ;
        RECT 2438.975 1947.755 2440.225 1947.825 ;
        RECT 2438.975 1947.595 2439.265 1947.755 ;
        RECT 2439.935 1947.595 2440.225 1947.755 ;
        RECT 2427.975 1947.035 2428.265 1947.265 ;
        RECT 2429.795 1946.490 2429.965 1947.445 ;
        RECT 2431.310 1946.875 2431.630 1946.980 ;
        RECT 2431.285 1946.860 2431.630 1946.875 ;
        RECT 2431.280 1946.845 2431.630 1946.860 ;
        RECT 2431.110 1946.675 2431.630 1946.845 ;
        RECT 2431.285 1946.660 2431.630 1946.675 ;
        RECT 2431.285 1946.645 2431.575 1946.660 ;
        RECT 2432.085 1946.490 2432.435 1946.610 ;
        RECT 2433.445 1946.545 2433.735 1946.780 ;
        RECT 2434.430 1946.545 2434.720 1946.780 ;
        RECT 2433.445 1946.540 2433.675 1946.545 ;
        RECT 2434.430 1946.540 2434.660 1946.545 ;
        RECT 2424.555 1946.425 2424.875 1946.445 ;
        RECT 2424.335 1946.385 2424.875 1946.425 ;
        RECT 2423.885 1946.245 2424.875 1946.385 ;
        RECT 2424.335 1946.195 2424.875 1946.245 ;
        RECT 2424.555 1946.185 2424.875 1946.195 ;
        RECT 2425.155 1946.185 2425.835 1946.445 ;
        RECT 2426.275 1946.385 2426.595 1946.445 ;
        RECT 2426.775 1946.385 2427.065 1946.425 ;
        RECT 2426.275 1946.245 2427.065 1946.385 ;
        RECT 2427.685 1946.245 2428.035 1946.445 ;
        RECT 2429.795 1946.320 2432.435 1946.490 ;
        RECT 2431.915 1946.315 2432.435 1946.320 ;
        RECT 2432.085 1946.260 2432.435 1946.315 ;
        RECT 2426.275 1946.185 2426.595 1946.245 ;
        RECT 2426.775 1946.195 2427.065 1946.245 ;
        RECT 2427.715 1946.185 2428.035 1946.245 ;
        RECT 2433.080 1946.225 2433.310 1946.245 ;
        RECT 2431.655 1946.120 2431.945 1946.145 ;
        RECT 2433.050 1946.120 2433.340 1946.225 ;
        RECT 2431.655 1945.950 2433.340 1946.120 ;
        RECT 2431.655 1945.915 2431.945 1945.950 ;
        RECT 2433.050 1945.915 2433.340 1945.950 ;
        RECT 2413.095 1945.175 2413.385 1945.405 ;
        RECT 2414.885 1945.180 2415.180 1945.440 ;
        RECT 2415.870 1945.180 2416.310 1945.440 ;
        RECT 2431.715 1945.405 2431.885 1945.915 ;
        RECT 2433.080 1945.895 2433.310 1945.915 ;
        RECT 2433.505 1945.440 2433.675 1946.540 ;
        RECT 2434.490 1945.440 2434.660 1946.540 ;
        RECT 2436.115 1946.425 2436.275 1947.555 ;
        RECT 2436.995 1947.305 2437.315 1947.565 ;
        RECT 2438.115 1947.445 2438.435 1947.565 ;
        RECT 2439.455 1947.505 2439.745 1947.545 ;
        RECT 2438.115 1947.305 2438.945 1947.445 ;
        RECT 2439.455 1947.315 2439.785 1947.505 ;
        RECT 2438.735 1947.265 2438.945 1947.305 ;
        RECT 2438.735 1947.035 2439.025 1947.265 ;
        RECT 2436.515 1946.985 2436.835 1947.005 ;
        RECT 2436.515 1946.845 2437.465 1946.985 ;
        RECT 2437.925 1946.945 2438.215 1946.985 ;
        RECT 2436.515 1946.755 2437.065 1946.845 ;
        RECT 2437.325 1946.805 2437.465 1946.845 ;
        RECT 2437.825 1946.805 2438.215 1946.945 ;
        RECT 2437.325 1946.755 2438.215 1946.805 ;
        RECT 2436.515 1946.745 2436.835 1946.755 ;
        RECT 2437.325 1946.665 2437.965 1946.755 ;
        RECT 2436.055 1946.195 2436.345 1946.425 ;
        RECT 2436.995 1946.385 2437.315 1946.445 ;
        RECT 2438.955 1946.385 2439.275 1946.445 ;
        RECT 2439.645 1946.425 2439.785 1947.315 ;
        RECT 2440.435 1947.305 2440.755 1947.565 ;
        RECT 2441.155 1947.305 2441.475 1947.565 ;
        RECT 2441.725 1947.505 2441.865 1947.925 ;
        RECT 2442.355 1947.865 2442.675 1948.125 ;
        RECT 2442.895 1948.065 2443.185 1948.105 ;
        RECT 2443.355 1948.065 2443.675 1948.125 ;
        RECT 2442.895 1947.925 2443.675 1948.065 ;
        RECT 2442.895 1947.875 2443.185 1947.925 ;
        RECT 2443.355 1947.865 2443.675 1947.925 ;
        RECT 2443.835 1947.865 2444.155 1948.125 ;
        RECT 2444.315 1947.865 2444.635 1948.125 ;
        RECT 2445.315 1947.895 2445.635 1948.125 ;
        RECT 2445.315 1947.865 2446.745 1947.895 ;
        RECT 2445.405 1947.755 2446.745 1947.865 ;
        RECT 2442.895 1947.505 2443.185 1947.545 ;
        RECT 2441.725 1947.365 2443.185 1947.505 ;
        RECT 2442.895 1947.315 2443.185 1947.365 ;
        RECT 2444.835 1947.305 2445.155 1947.565 ;
        RECT 2445.405 1947.545 2445.545 1947.755 ;
        RECT 2445.335 1947.315 2445.625 1947.545 ;
        RECT 2446.055 1947.505 2446.345 1947.545 ;
        RECT 2446.055 1947.315 2446.385 1947.505 ;
        RECT 2444.335 1947.225 2444.625 1947.265 ;
        RECT 2444.835 1947.225 2445.065 1947.305 ;
        RECT 2444.335 1947.085 2445.065 1947.225 ;
        RECT 2444.335 1947.035 2444.625 1947.085 ;
        RECT 2440.175 1946.985 2440.495 1947.005 ;
        RECT 2439.935 1946.945 2440.495 1946.985 ;
        RECT 2441.175 1946.945 2441.465 1946.985 ;
        RECT 2439.935 1946.805 2441.465 1946.945 ;
        RECT 2439.935 1946.755 2440.495 1946.805 ;
        RECT 2441.175 1946.755 2441.465 1946.805 ;
        RECT 2441.655 1946.945 2441.945 1946.985 ;
        RECT 2441.655 1946.805 2442.585 1946.945 ;
        RECT 2441.655 1946.755 2441.945 1946.805 ;
        RECT 2440.175 1946.745 2440.495 1946.755 ;
        RECT 2436.995 1946.245 2439.275 1946.385 ;
        RECT 2436.995 1946.185 2437.315 1946.245 ;
        RECT 2438.955 1946.185 2439.275 1946.245 ;
        RECT 2439.455 1946.385 2439.785 1946.425 ;
        RECT 2440.435 1946.385 2440.755 1946.445 ;
        RECT 2441.155 1946.425 2441.475 1946.445 ;
        RECT 2439.455 1946.245 2440.755 1946.385 ;
        RECT 2439.455 1946.195 2439.745 1946.245 ;
        RECT 2440.435 1946.185 2440.755 1946.245 ;
        RECT 2440.935 1946.195 2441.475 1946.425 ;
        RECT 2441.155 1946.185 2441.475 1946.195 ;
        RECT 2441.875 1946.185 2442.195 1946.445 ;
        RECT 2442.445 1946.385 2442.585 1946.805 ;
        RECT 2442.875 1946.805 2443.195 1947.005 ;
        RECT 2445.575 1946.805 2445.865 1946.985 ;
        RECT 2442.875 1946.755 2445.865 1946.805 ;
        RECT 2442.875 1946.745 2445.785 1946.755 ;
        RECT 2442.965 1946.665 2445.785 1946.745 ;
        RECT 2446.245 1946.445 2446.385 1947.315 ;
        RECT 2446.605 1947.265 2446.745 1947.755 ;
        RECT 2448.265 1947.445 2448.605 1947.795 ;
        RECT 2446.535 1947.035 2446.825 1947.265 ;
        RECT 2448.355 1946.490 2448.525 1947.445 ;
        RECT 2452.990 1947.420 2453.280 1947.465 ;
        RECT 2466.590 1947.420 2466.910 1947.480 ;
        RECT 2452.990 1947.280 2466.910 1947.420 ;
        RECT 2452.990 1947.235 2453.280 1947.280 ;
        RECT 2466.590 1947.220 2466.910 1947.280 ;
        RECT 2449.870 1946.875 2450.190 1946.980 ;
        RECT 2449.845 1946.860 2450.190 1946.875 ;
        RECT 2449.840 1946.845 2450.190 1946.860 ;
        RECT 2449.670 1946.675 2450.190 1946.845 ;
        RECT 2449.845 1946.660 2450.190 1946.675 ;
        RECT 2449.845 1946.645 2450.135 1946.660 ;
        RECT 2450.645 1946.490 2450.995 1946.610 ;
        RECT 2452.005 1946.545 2452.295 1946.780 ;
        RECT 2452.990 1946.545 2453.280 1946.780 ;
        RECT 2452.005 1946.540 2452.235 1946.545 ;
        RECT 2452.990 1946.540 2453.220 1946.545 ;
        RECT 2443.115 1946.425 2443.435 1946.445 ;
        RECT 2442.895 1946.385 2443.435 1946.425 ;
        RECT 2442.445 1946.245 2443.435 1946.385 ;
        RECT 2442.895 1946.195 2443.435 1946.245 ;
        RECT 2443.115 1946.185 2443.435 1946.195 ;
        RECT 2443.715 1946.185 2444.395 1946.445 ;
        RECT 2444.835 1946.385 2445.155 1946.445 ;
        RECT 2445.335 1946.385 2445.625 1946.425 ;
        RECT 2444.835 1946.245 2445.625 1946.385 ;
        RECT 2446.245 1946.245 2446.595 1946.445 ;
        RECT 2448.355 1946.320 2450.995 1946.490 ;
        RECT 2450.475 1946.315 2450.995 1946.320 ;
        RECT 2450.645 1946.260 2450.995 1946.315 ;
        RECT 2444.835 1946.185 2445.155 1946.245 ;
        RECT 2445.335 1946.195 2445.625 1946.245 ;
        RECT 2446.275 1946.185 2446.595 1946.245 ;
        RECT 2451.640 1946.225 2451.870 1946.245 ;
        RECT 2450.215 1946.120 2450.505 1946.145 ;
        RECT 2451.610 1946.120 2451.900 1946.225 ;
        RECT 2450.215 1945.950 2451.900 1946.120 ;
        RECT 2450.215 1945.915 2450.505 1945.950 ;
        RECT 2451.610 1945.915 2451.900 1945.950 ;
        RECT 2431.655 1945.175 2431.945 1945.405 ;
        RECT 2433.445 1945.180 2433.740 1945.440 ;
        RECT 2434.390 1945.180 2434.725 1945.440 ;
        RECT 2450.275 1945.405 2450.445 1945.915 ;
        RECT 2451.640 1945.895 2451.870 1945.915 ;
        RECT 2452.065 1945.440 2452.235 1946.540 ;
        RECT 2453.050 1945.440 2453.220 1946.540 ;
        RECT 2450.215 1945.175 2450.505 1945.405 ;
        RECT 2452.005 1945.180 2452.300 1945.440 ;
        RECT 2452.990 1945.180 2453.285 1945.440 ;
        RECT 2378.730 1938.720 2379.050 1938.980 ;
        RECT 2397.130 1938.920 2397.450 1938.980 ;
        RECT 2576.990 1938.920 2577.310 1938.980 ;
        RECT 2397.130 1938.780 2577.310 1938.920 ;
        RECT 2397.130 1938.720 2397.450 1938.780 ;
        RECT 2576.990 1938.720 2577.310 1938.780 ;
        RECT 2378.820 1938.580 2378.960 1938.720 ;
        RECT 2473.490 1938.580 2473.810 1938.640 ;
        RECT 2378.820 1938.440 2473.810 1938.580 ;
        RECT 2473.490 1938.380 2473.810 1938.440 ;
        RECT 2415.990 1932.120 2416.310 1932.180 ;
        RECT 2421.510 1932.120 2421.830 1932.180 ;
        RECT 2415.990 1931.980 2421.830 1932.120 ;
        RECT 2415.990 1931.920 2416.310 1931.980 ;
        RECT 2421.510 1931.920 2421.830 1931.980 ;
        RECT 2604.590 1869.900 2604.910 1869.960 ;
        RECT 2677.270 1869.900 2677.590 1869.960 ;
        RECT 2604.590 1869.760 2677.590 1869.900 ;
        RECT 2604.590 1869.700 2604.910 1869.760 ;
        RECT 2677.270 1869.700 2677.590 1869.760 ;
        RECT 2611.490 1862.760 2611.810 1862.820 ;
        RECT 2677.270 1862.760 2677.590 1862.820 ;
        RECT 2611.490 1862.620 2677.590 1862.760 ;
        RECT 2611.490 1862.560 2611.810 1862.620 ;
        RECT 2677.270 1862.560 2677.590 1862.620 ;
        RECT 2695.590 1856.480 2695.910 1856.540 ;
        RECT 2698.810 1856.480 2699.130 1856.540 ;
        RECT 2700.205 1856.480 2700.495 1856.525 ;
        RECT 2695.590 1856.340 2698.120 1856.480 ;
        RECT 2695.590 1856.280 2695.910 1856.340 ;
        RECT 2697.980 1856.140 2698.120 1856.340 ;
        RECT 2698.810 1856.340 2700.495 1856.480 ;
        RECT 2698.810 1856.280 2699.130 1856.340 ;
        RECT 2700.205 1856.295 2700.495 1856.340 ;
        RECT 2702.490 1856.480 2702.810 1856.540 ;
        RECT 2709.865 1856.480 2710.155 1856.525 ;
        RECT 2702.490 1856.340 2710.155 1856.480 ;
        RECT 2702.490 1856.280 2702.810 1856.340 ;
        RECT 2709.865 1856.295 2710.155 1856.340 ;
        RECT 2697.980 1856.000 2701.340 1856.140 ;
        RECT 2695.130 1855.800 2695.450 1855.860 ;
        RECT 2701.200 1855.845 2701.340 1856.000 ;
        RECT 2699.745 1855.800 2700.035 1855.845 ;
        RECT 2695.130 1855.660 2700.035 1855.800 ;
        RECT 2695.130 1855.600 2695.450 1855.660 ;
        RECT 2699.745 1855.615 2700.035 1855.660 ;
        RECT 2701.125 1855.615 2701.415 1855.845 ;
        RECT 2698.365 1855.460 2698.655 1855.505 ;
        RECT 2701.570 1855.460 2701.890 1855.520 ;
        RECT 2698.365 1855.320 2701.890 1855.460 ;
        RECT 2698.365 1855.275 2698.655 1855.320 ;
        RECT 2701.570 1855.260 2701.890 1855.320 ;
        RECT 2721.810 1854.920 2722.130 1855.180 ;
        RECT 2698.350 1854.780 2698.670 1854.840 ;
        RECT 2698.825 1854.780 2699.115 1854.825 ;
        RECT 2698.350 1854.640 2699.115 1854.780 ;
        RECT 2698.350 1854.580 2698.670 1854.640 ;
        RECT 2698.825 1854.595 2699.115 1854.640 ;
        RECT 2731.470 1854.580 2731.790 1854.840 ;
        RECT 2694.670 1852.740 2694.990 1852.800 ;
        RECT 2696.985 1852.740 2697.275 1852.785 ;
        RECT 2694.670 1852.600 2697.275 1852.740 ;
        RECT 2694.670 1852.540 2694.990 1852.600 ;
        RECT 2696.985 1852.555 2697.275 1852.600 ;
        RECT 2697.890 1851.860 2698.210 1852.120 ;
        RECT 2421.510 1849.160 2421.830 1849.220 ;
        RECT 2677.270 1849.160 2677.590 1849.220 ;
        RECT 2421.510 1849.020 2677.590 1849.160 ;
        RECT 2421.510 1848.960 2421.830 1849.020 ;
        RECT 2677.270 1848.960 2677.590 1849.020 ;
        RECT 2694.670 1844.920 2694.990 1844.980 ;
        RECT 2696.985 1844.920 2697.275 1844.965 ;
        RECT 2694.670 1844.780 2697.275 1844.920 ;
        RECT 2694.670 1844.720 2694.990 1844.780 ;
        RECT 2696.985 1844.735 2697.275 1844.780 ;
        RECT 2696.970 1843.900 2697.290 1843.960 ;
        RECT 2697.905 1843.900 2698.195 1843.945 ;
        RECT 2696.970 1843.760 2698.195 1843.900 ;
        RECT 2696.970 1843.700 2697.290 1843.760 ;
        RECT 2697.905 1843.715 2698.195 1843.760 ;
        RECT 2697.430 1842.200 2697.750 1842.260 ;
        RECT 2698.350 1842.200 2698.670 1842.260 ;
        RECT 2697.430 1842.060 2698.670 1842.200 ;
        RECT 2697.430 1842.000 2697.750 1842.060 ;
        RECT 2698.350 1842.000 2698.670 1842.060 ;
        RECT 2698.370 1839.820 2698.660 1839.865 ;
        RECT 2703.890 1839.820 2704.180 1839.865 ;
        RECT 2704.810 1839.820 2705.100 1839.865 ;
        RECT 2698.370 1839.680 2705.100 1839.820 ;
        RECT 2698.370 1839.635 2698.660 1839.680 ;
        RECT 2703.890 1839.635 2704.180 1839.680 ;
        RECT 2704.810 1839.635 2705.100 1839.680 ;
        RECT 2696.985 1839.480 2697.275 1839.525 ;
        RECT 2697.430 1839.480 2697.750 1839.540 ;
        RECT 2696.985 1839.340 2697.750 1839.480 ;
        RECT 2696.985 1839.295 2697.275 1839.340 ;
        RECT 2697.430 1839.280 2697.750 1839.340 ;
        RECT 2697.890 1839.280 2698.210 1839.540 ;
        RECT 2699.290 1839.480 2699.580 1839.525 ;
        RECT 2701.130 1839.480 2701.420 1839.525 ;
        RECT 2699.290 1839.340 2701.420 1839.480 ;
        RECT 2699.290 1839.295 2699.580 1839.340 ;
        RECT 2701.130 1839.295 2701.420 1839.340 ;
        RECT 2703.475 1839.480 2703.765 1839.525 ;
        RECT 2705.315 1839.480 2705.605 1839.525 ;
        RECT 2703.475 1839.340 2705.605 1839.480 ;
        RECT 2703.475 1839.295 2703.765 1839.340 ;
        RECT 2705.315 1839.295 2705.605 1839.340 ;
        RECT 2721.810 1839.280 2722.130 1839.540 ;
        RECT 2702.030 1839.185 2702.350 1839.200 ;
        RECT 2701.585 1839.140 2701.875 1839.185 ;
        RECT 2697.520 1839.000 2701.875 1839.140 ;
        RECT 2697.520 1838.860 2697.660 1839.000 ;
        RECT 2701.585 1838.955 2701.875 1839.000 ;
        RECT 2702.030 1838.955 2702.460 1839.185 ;
        RECT 2702.950 1839.140 2703.270 1839.200 ;
        RECT 2721.900 1839.140 2722.040 1839.280 ;
        RECT 2702.950 1839.000 2722.040 1839.140 ;
        RECT 2702.030 1838.940 2702.350 1838.955 ;
        RECT 2702.950 1838.940 2703.270 1839.000 ;
        RECT 2697.430 1838.600 2697.750 1838.860 ;
        RECT 2700.205 1838.615 2700.495 1838.845 ;
        RECT 2701.165 1838.800 2701.455 1838.845 ;
        RECT 2704.395 1838.800 2704.685 1838.845 ;
        RECT 2701.165 1838.660 2704.685 1838.800 ;
        RECT 2701.165 1838.615 2701.455 1838.660 ;
        RECT 2704.395 1838.615 2704.685 1838.660 ;
        RECT 2700.280 1838.460 2700.420 1838.615 ;
        RECT 2702.490 1838.460 2702.810 1838.520 ;
        RECT 2700.280 1838.320 2702.810 1838.460 ;
        RECT 2702.490 1838.260 2702.810 1838.320 ;
        RECT 2703.870 1838.460 2704.190 1838.520 ;
        RECT 2706.185 1838.460 2706.475 1838.505 ;
        RECT 2703.870 1838.320 2706.475 1838.460 ;
        RECT 2703.870 1838.260 2704.190 1838.320 ;
        RECT 2706.185 1838.275 2706.475 1838.320 ;
        RECT 2697.905 1837.440 2698.195 1837.485 ;
        RECT 2702.030 1837.440 2702.350 1837.500 ;
        RECT 2697.905 1837.300 2702.350 1837.440 ;
        RECT 2697.905 1837.255 2698.195 1837.300 ;
        RECT 2702.030 1837.240 2702.350 1837.300 ;
        RECT 2694.670 1836.420 2694.990 1836.480 ;
        RECT 2696.985 1836.420 2697.275 1836.465 ;
        RECT 2694.670 1836.280 2697.275 1836.420 ;
        RECT 2694.670 1836.220 2694.990 1836.280 ;
        RECT 2696.985 1836.235 2697.275 1836.280 ;
        RECT 2604.590 1835.560 2604.910 1835.620 ;
        RECT 2677.270 1835.560 2677.590 1835.620 ;
        RECT 2604.590 1835.420 2677.590 1835.560 ;
        RECT 2604.590 1835.360 2604.910 1835.420 ;
        RECT 2677.270 1835.360 2677.590 1835.420 ;
        RECT 2698.370 1834.380 2698.660 1834.425 ;
        RECT 2703.890 1834.380 2704.180 1834.425 ;
        RECT 2704.810 1834.380 2705.100 1834.425 ;
        RECT 2698.370 1834.240 2705.100 1834.380 ;
        RECT 2698.370 1834.195 2698.660 1834.240 ;
        RECT 2703.890 1834.195 2704.180 1834.240 ;
        RECT 2704.810 1834.195 2705.100 1834.240 ;
        RECT 2696.970 1833.840 2697.290 1834.100 ;
        RECT 2697.890 1833.840 2698.210 1834.100 ;
        RECT 2699.290 1834.040 2699.580 1834.085 ;
        RECT 2701.130 1834.040 2701.420 1834.085 ;
        RECT 2699.290 1833.900 2701.420 1834.040 ;
        RECT 2699.290 1833.855 2699.580 1833.900 ;
        RECT 2701.130 1833.855 2701.420 1833.900 ;
        RECT 2702.950 1833.840 2703.270 1834.100 ;
        RECT 2703.475 1834.040 2703.765 1834.085 ;
        RECT 2705.315 1834.040 2705.605 1834.085 ;
        RECT 2703.475 1833.900 2705.605 1834.040 ;
        RECT 2703.475 1833.855 2703.765 1833.900 ;
        RECT 2705.315 1833.855 2705.605 1833.900 ;
        RECT 2698.810 1833.700 2699.130 1833.760 ;
        RECT 2702.030 1833.745 2702.350 1833.760 ;
        RECT 2701.585 1833.700 2701.875 1833.745 ;
        RECT 2698.810 1833.560 2701.875 1833.700 ;
        RECT 2698.810 1833.500 2699.130 1833.560 ;
        RECT 2701.585 1833.515 2701.875 1833.560 ;
        RECT 2702.030 1833.515 2702.460 1833.745 ;
        RECT 2702.030 1833.500 2702.350 1833.515 ;
        RECT 2700.205 1833.175 2700.495 1833.405 ;
        RECT 2701.165 1833.360 2701.455 1833.405 ;
        RECT 2704.395 1833.360 2704.685 1833.405 ;
        RECT 2701.165 1833.220 2704.685 1833.360 ;
        RECT 2701.165 1833.175 2701.455 1833.220 ;
        RECT 2704.395 1833.175 2704.685 1833.220 ;
        RECT 2698.350 1833.020 2698.670 1833.080 ;
        RECT 2700.280 1833.020 2700.420 1833.175 ;
        RECT 2702.490 1833.020 2702.810 1833.080 ;
        RECT 2698.350 1832.880 2702.810 1833.020 ;
        RECT 2698.350 1832.820 2698.670 1832.880 ;
        RECT 2702.490 1832.820 2702.810 1832.880 ;
        RECT 2706.170 1832.820 2706.490 1833.080 ;
        RECT 2697.905 1832.000 2698.195 1832.045 ;
        RECT 2702.030 1832.000 2702.350 1832.060 ;
        RECT 2706.170 1832.000 2706.490 1832.060 ;
        RECT 2697.905 1831.860 2702.350 1832.000 ;
        RECT 2697.905 1831.815 2698.195 1831.860 ;
        RECT 2702.030 1831.800 2702.350 1831.860 ;
        RECT 2703.960 1831.860 2706.490 1832.000 ;
        RECT 2697.890 1831.320 2698.210 1831.380 ;
        RECT 2701.570 1831.320 2701.890 1831.380 ;
        RECT 2703.960 1831.365 2704.100 1831.860 ;
        RECT 2706.170 1831.800 2706.490 1831.860 ;
        RECT 2697.890 1831.180 2703.640 1831.320 ;
        RECT 2697.890 1831.120 2698.210 1831.180 ;
        RECT 2701.570 1831.120 2701.890 1831.180 ;
        RECT 2694.670 1830.980 2694.990 1831.040 ;
        RECT 2696.985 1830.980 2697.275 1831.025 ;
        RECT 2694.670 1830.840 2697.275 1830.980 ;
        RECT 2703.500 1830.980 2703.640 1831.180 ;
        RECT 2703.885 1831.135 2704.175 1831.365 ;
        RECT 2704.345 1831.135 2704.635 1831.365 ;
        RECT 2704.420 1830.980 2704.560 1831.135 ;
        RECT 2703.500 1830.840 2704.560 1830.980 ;
        RECT 2694.670 1830.780 2694.990 1830.840 ;
        RECT 2696.985 1830.795 2697.275 1830.840 ;
        RECT 2703.425 1830.640 2703.715 1830.685 ;
        RECT 2703.870 1830.640 2704.190 1830.700 ;
        RECT 2703.425 1830.500 2704.190 1830.640 ;
        RECT 2703.425 1830.455 2703.715 1830.500 ;
        RECT 2703.870 1830.440 2704.190 1830.500 ;
        RECT 2701.570 1830.100 2701.890 1830.360 ;
        RECT 2576.990 1828.760 2577.310 1828.820 ;
        RECT 2677.270 1828.760 2677.590 1828.820 ;
        RECT 2576.990 1828.620 2677.590 1828.760 ;
        RECT 2576.990 1828.560 2577.310 1828.620 ;
        RECT 2677.270 1828.560 2677.590 1828.620 ;
        RECT 2697.430 1826.560 2697.750 1826.620 ;
        RECT 2697.905 1826.560 2698.195 1826.605 ;
        RECT 2697.430 1826.420 2698.195 1826.560 ;
        RECT 2697.430 1826.360 2697.750 1826.420 ;
        RECT 2697.905 1826.375 2698.195 1826.420 ;
        RECT 2694.670 1825.540 2694.990 1825.600 ;
        RECT 2696.985 1825.540 2697.275 1825.585 ;
        RECT 2694.670 1825.400 2697.275 1825.540 ;
        RECT 2694.670 1825.340 2694.990 1825.400 ;
        RECT 2696.985 1825.355 2697.275 1825.400 ;
        RECT 2701.570 1819.900 2701.890 1820.160 ;
        RECT 2702.505 1820.100 2702.795 1820.145 ;
        RECT 2703.870 1820.100 2704.190 1820.160 ;
        RECT 2731.470 1820.100 2731.790 1820.160 ;
        RECT 2702.505 1819.960 2731.790 1820.100 ;
        RECT 2702.505 1819.915 2702.795 1819.960 ;
        RECT 2703.870 1819.900 2704.190 1819.960 ;
        RECT 2731.470 1819.900 2731.790 1819.960 ;
        RECT 2702.030 1819.220 2702.350 1819.480 ;
        RECT 2697.905 1818.400 2698.195 1818.445 ;
        RECT 2698.810 1818.400 2699.130 1818.460 ;
        RECT 2697.905 1818.260 2699.130 1818.400 ;
        RECT 2697.905 1818.215 2698.195 1818.260 ;
        RECT 2698.810 1818.200 2699.130 1818.260 ;
        RECT 2702.030 1818.200 2702.350 1818.460 ;
        RECT 2703.870 1818.200 2704.190 1818.460 ;
        RECT 2694.670 1817.720 2694.990 1817.780 ;
        RECT 2702.120 1817.765 2702.260 1818.200 ;
        RECT 2703.960 1817.765 2704.100 1818.200 ;
        RECT 2696.985 1817.720 2697.275 1817.765 ;
        RECT 2694.670 1817.580 2697.275 1817.720 ;
        RECT 2694.670 1817.520 2694.990 1817.580 ;
        RECT 2696.985 1817.535 2697.275 1817.580 ;
        RECT 2702.045 1817.535 2702.335 1817.765 ;
        RECT 2703.885 1817.535 2704.175 1817.765 ;
        RECT 2704.790 1817.180 2705.110 1817.440 ;
        RECT 2702.490 1816.840 2702.810 1817.100 ;
        RECT 2702.490 1815.680 2702.810 1815.740 ;
        RECT 2702.490 1815.540 2724.570 1815.680 ;
        RECT 2702.490 1815.480 2702.810 1815.540 ;
        RECT 2724.430 1814.660 2724.570 1815.540 ;
        RECT 2725.505 1814.660 2725.795 1814.705 ;
        RECT 2724.430 1814.520 2725.795 1814.660 ;
        RECT 2725.505 1814.475 2725.795 1814.520 ;
        RECT 2694.670 1812.280 2694.990 1812.340 ;
        RECT 2696.985 1812.280 2697.275 1812.325 ;
        RECT 2694.670 1812.140 2697.275 1812.280 ;
        RECT 2694.670 1812.080 2694.990 1812.140 ;
        RECT 2696.985 1812.095 2697.275 1812.140 ;
        RECT 2697.430 1811.260 2697.750 1811.320 ;
        RECT 2697.905 1811.260 2698.195 1811.305 ;
        RECT 2697.430 1811.120 2698.195 1811.260 ;
        RECT 2697.430 1811.060 2697.750 1811.120 ;
        RECT 2697.905 1811.075 2698.195 1811.120 ;
        RECT 2611.490 1808.020 2611.810 1808.080 ;
        RECT 2677.270 1808.020 2677.590 1808.080 ;
        RECT 2611.490 1807.880 2677.590 1808.020 ;
        RECT 2611.490 1807.820 2611.810 1807.880 ;
        RECT 2677.270 1807.820 2677.590 1807.880 ;
        RECT 2697.890 1806.640 2698.210 1806.900 ;
        RECT 2698.350 1806.640 2698.670 1806.900 ;
        RECT 2697.430 1806.300 2697.750 1806.560 ;
        RECT 2697.980 1806.500 2698.120 1806.640 ;
        RECT 2702.030 1806.500 2702.350 1806.560 ;
        RECT 2697.980 1806.360 2702.350 1806.500 ;
        RECT 2702.030 1806.300 2702.350 1806.360 ;
        RECT 2523.545 1805.780 2523.865 1806.040 ;
        RECT 2699.285 1805.820 2699.575 1805.865 ;
        RECT 2702.950 1805.820 2703.270 1805.880 ;
        RECT 2699.285 1805.680 2703.270 1805.820 ;
        RECT 2699.285 1805.635 2699.575 1805.680 ;
        RECT 2702.950 1805.620 2703.270 1805.680 ;
        RECT 2694.670 1803.780 2694.990 1803.840 ;
        RECT 2696.985 1803.780 2697.275 1803.825 ;
        RECT 2694.670 1803.640 2697.275 1803.780 ;
        RECT 2694.670 1803.580 2694.990 1803.640 ;
        RECT 2696.985 1803.595 2697.275 1803.640 ;
        RECT 2697.890 1802.900 2698.210 1803.160 ;
        RECT 2697.890 1802.080 2698.210 1802.140 ;
        RECT 2698.825 1802.080 2699.115 1802.125 ;
        RECT 2697.890 1801.940 2699.115 1802.080 ;
        RECT 2697.890 1801.880 2698.210 1801.940 ;
        RECT 2698.825 1801.895 2699.115 1801.940 ;
        RECT 2700.665 1802.080 2700.955 1802.125 ;
        RECT 2701.585 1802.080 2701.875 1802.125 ;
        RECT 2700.665 1801.940 2701.875 1802.080 ;
        RECT 2700.665 1801.895 2700.955 1801.940 ;
        RECT 2701.585 1801.895 2701.875 1801.940 ;
        RECT 2702.030 1801.880 2702.350 1802.140 ;
        RECT 2702.950 1801.880 2703.270 1802.140 ;
        RECT 2703.410 1801.880 2703.730 1802.140 ;
        RECT 2698.350 1801.740 2698.670 1801.800 ;
        RECT 2697.980 1801.600 2698.670 1801.740 ;
        RECT 2697.980 1801.105 2698.120 1801.600 ;
        RECT 2698.350 1801.540 2698.670 1801.600 ;
        RECT 2702.120 1801.445 2702.260 1801.880 ;
        RECT 2702.045 1801.215 2702.335 1801.445 ;
        RECT 2702.490 1801.200 2702.810 1801.460 ;
        RECT 2703.040 1801.445 2703.180 1801.880 ;
        RECT 2702.965 1801.215 2703.255 1801.445 ;
        RECT 2697.905 1800.875 2698.195 1801.105 ;
        RECT 2698.350 1800.860 2698.670 1801.120 ;
        RECT 2702.580 1801.060 2702.720 1801.200 ;
        RECT 2703.425 1801.060 2703.715 1801.105 ;
        RECT 2702.580 1800.920 2703.715 1801.060 ;
        RECT 2703.425 1800.875 2703.715 1800.920 ;
        RECT 2702.490 1800.180 2702.810 1800.440 ;
        RECT 2698.810 1799.160 2699.130 1799.420 ;
        RECT 2699.745 1799.360 2700.035 1799.405 ;
        RECT 2702.490 1799.360 2702.810 1799.420 ;
        RECT 2699.745 1799.220 2702.810 1799.360 ;
        RECT 2699.745 1799.175 2700.035 1799.220 ;
        RECT 2702.490 1799.160 2702.810 1799.220 ;
        RECT 2696.985 1799.020 2697.275 1799.065 ;
        RECT 2697.430 1799.020 2697.750 1799.080 ;
        RECT 2696.985 1798.880 2697.750 1799.020 ;
        RECT 2698.900 1799.020 2699.040 1799.160 ;
        RECT 2702.030 1799.020 2702.350 1799.080 ;
        RECT 2698.900 1798.880 2702.350 1799.020 ;
        RECT 2696.985 1798.835 2697.275 1798.880 ;
        RECT 2697.430 1798.820 2697.750 1798.880 ;
        RECT 2702.030 1798.820 2702.350 1798.880 ;
        RECT 2523.545 1798.250 2523.865 1798.510 ;
        RECT 2698.810 1797.460 2699.130 1797.720 ;
        RECT 2697.905 1796.640 2698.195 1796.685 ;
        RECT 2698.810 1796.640 2699.130 1796.700 ;
        RECT 2697.905 1796.500 2699.130 1796.640 ;
        RECT 2697.905 1796.455 2698.195 1796.500 ;
        RECT 2698.810 1796.440 2699.130 1796.500 ;
        RECT 2694.670 1795.960 2694.990 1796.020 ;
        RECT 2696.985 1795.960 2697.275 1796.005 ;
        RECT 2694.670 1795.820 2697.275 1795.960 ;
        RECT 2694.670 1795.760 2694.990 1795.820 ;
        RECT 2696.985 1795.775 2697.275 1795.820 ;
        RECT 2700.205 1793.240 2700.495 1793.285 ;
        RECT 2701.570 1793.240 2701.890 1793.300 ;
        RECT 2700.205 1793.100 2701.890 1793.240 ;
        RECT 2700.205 1793.055 2700.495 1793.100 ;
        RECT 2701.570 1793.040 2701.890 1793.100 ;
        RECT 2698.365 1792.900 2698.655 1792.945 ;
        RECT 2699.730 1792.900 2700.050 1792.960 ;
        RECT 2698.365 1792.760 2700.050 1792.900 ;
        RECT 2698.365 1792.715 2698.655 1792.760 ;
        RECT 2699.730 1792.700 2700.050 1792.760 ;
        RECT 2700.665 1792.900 2700.955 1792.945 ;
        RECT 2703.410 1792.900 2703.730 1792.960 ;
        RECT 2700.665 1792.760 2703.730 1792.900 ;
        RECT 2700.665 1792.715 2700.955 1792.760 ;
        RECT 2703.410 1792.700 2703.730 1792.760 ;
        RECT 2696.970 1792.560 2697.290 1792.620 ;
        RECT 2702.030 1792.560 2702.350 1792.620 ;
        RECT 2523.545 1792.270 2523.865 1792.530 ;
        RECT 2696.970 1792.420 2702.350 1792.560 ;
        RECT 2696.970 1792.360 2697.290 1792.420 ;
        RECT 2702.030 1792.360 2702.350 1792.420 ;
        RECT 2698.810 1792.020 2699.130 1792.280 ;
        RECT 2699.270 1792.020 2699.590 1792.280 ;
        RECT 2701.585 1792.220 2701.875 1792.265 ;
        RECT 2703.870 1792.220 2704.190 1792.280 ;
        RECT 2701.585 1792.080 2704.190 1792.220 ;
        RECT 2701.585 1792.035 2701.875 1792.080 ;
        RECT 2703.870 1792.020 2704.190 1792.080 ;
        RECT 2698.810 1791.200 2699.130 1791.260 ;
        RECT 2701.125 1791.200 2701.415 1791.245 ;
        RECT 2698.810 1791.060 2701.415 1791.200 ;
        RECT 2698.810 1791.000 2699.130 1791.060 ;
        RECT 2701.125 1791.015 2701.415 1791.060 ;
        RECT 2699.730 1790.860 2700.050 1790.920 ;
        RECT 2697.520 1790.720 2699.500 1790.860 ;
        RECT 2697.520 1790.580 2697.660 1790.720 ;
        RECT 2697.430 1790.320 2697.750 1790.580 ;
        RECT 2697.890 1790.320 2698.210 1790.580 ;
        RECT 2369.490 1790.060 2369.780 1790.290 ;
        RECT 2377.005 1790.060 2377.295 1790.290 ;
        RECT 2382.620 1790.060 2382.910 1790.290 ;
        RECT 2369.550 1789.610 2369.720 1790.060 ;
        RECT 2377.065 1789.715 2377.235 1790.060 ;
        RECT 2369.460 1789.320 2369.810 1789.610 ;
        RECT 2376.965 1789.345 2377.335 1789.715 ;
        RECT 2382.680 1789.580 2382.850 1790.060 ;
        RECT 2384.410 1790.030 2384.705 1790.290 ;
        RECT 2385.400 1790.030 2385.695 1790.290 ;
        RECT 2392.265 1790.060 2392.555 1790.290 ;
        RECT 2397.880 1790.060 2398.170 1790.290 ;
        RECT 2383.590 1789.580 2383.940 1789.610 ;
        RECT 2382.680 1789.550 2383.940 1789.580 ;
        RECT 2382.620 1789.410 2383.940 1789.550 ;
        RECT 2377.005 1789.320 2377.295 1789.345 ;
        RECT 2382.620 1789.320 2382.910 1789.410 ;
        RECT 2383.590 1789.320 2383.940 1789.410 ;
        RECT 2377.635 1789.180 2377.985 1789.245 ;
        RECT 2383.075 1789.180 2383.400 1789.270 ;
        RECT 2377.435 1789.150 2377.985 1789.180 ;
        RECT 2383.050 1789.150 2383.400 1789.180 ;
        RECT 2377.265 1789.145 2377.985 1789.150 ;
        RECT 2382.880 1789.145 2383.400 1789.150 ;
        RECT 2377.265 1788.980 2383.400 1789.145 ;
        RECT 2377.325 1788.975 2383.400 1788.980 ;
        RECT 2377.435 1788.950 2377.985 1788.975 ;
        RECT 2383.050 1788.950 2383.400 1788.975 ;
        RECT 2377.635 1788.895 2377.985 1788.950 ;
        RECT 2383.075 1788.945 2383.400 1788.950 ;
        RECT 2384.470 1788.930 2384.640 1790.030 ;
        RECT 2385.460 1789.300 2385.630 1790.030 ;
        RECT 2392.325 1789.715 2392.495 1790.060 ;
        RECT 2392.225 1789.345 2392.595 1789.715 ;
        RECT 2397.940 1789.580 2398.110 1790.060 ;
        RECT 2399.670 1790.030 2399.965 1790.290 ;
        RECT 2400.660 1790.030 2400.955 1790.290 ;
        RECT 2407.525 1790.060 2407.815 1790.290 ;
        RECT 2413.140 1790.060 2413.430 1790.290 ;
        RECT 2398.850 1789.580 2399.200 1789.610 ;
        RECT 2397.940 1789.550 2399.200 1789.580 ;
        RECT 2397.880 1789.410 2399.200 1789.550 ;
        RECT 2392.265 1789.320 2392.555 1789.345 ;
        RECT 2397.880 1789.320 2398.170 1789.410 ;
        RECT 2398.850 1789.320 2399.200 1789.410 ;
        RECT 2385.455 1788.950 2385.805 1789.300 ;
        RECT 2392.895 1789.180 2393.245 1789.255 ;
        RECT 2398.335 1789.180 2398.660 1789.270 ;
        RECT 2392.695 1789.150 2393.245 1789.180 ;
        RECT 2398.310 1789.150 2398.660 1789.180 ;
        RECT 2392.525 1789.145 2393.245 1789.150 ;
        RECT 2398.140 1789.145 2398.660 1789.150 ;
        RECT 2392.525 1788.980 2398.660 1789.145 ;
        RECT 2392.585 1788.975 2398.660 1788.980 ;
        RECT 2392.695 1788.950 2393.245 1788.975 ;
        RECT 2398.310 1788.950 2398.660 1788.975 ;
        RECT 2385.455 1788.930 2385.750 1788.950 ;
        RECT 2384.410 1788.925 2384.640 1788.930 ;
        RECT 2369.085 1788.790 2369.435 1788.865 ;
        RECT 2382.275 1788.820 2382.595 1788.835 ;
        RECT 2382.250 1788.790 2382.595 1788.820 ;
        RECT 2368.945 1788.620 2369.435 1788.790 ;
        RECT 2382.075 1788.620 2382.595 1788.790 ;
        RECT 2384.410 1788.690 2384.700 1788.925 ;
        RECT 2385.400 1788.865 2385.750 1788.930 ;
        RECT 2392.895 1788.905 2393.245 1788.950 ;
        RECT 2398.335 1788.945 2398.660 1788.950 ;
        RECT 2399.730 1788.930 2399.900 1790.030 ;
        RECT 2400.720 1789.305 2400.890 1790.030 ;
        RECT 2407.585 1789.715 2407.755 1790.060 ;
        RECT 2407.485 1789.345 2407.855 1789.715 ;
        RECT 2413.200 1789.580 2413.370 1790.060 ;
        RECT 2414.930 1790.030 2415.225 1790.290 ;
        RECT 2415.920 1790.030 2416.215 1790.290 ;
        RECT 2422.785 1790.060 2423.075 1790.290 ;
        RECT 2428.400 1790.060 2428.690 1790.290 ;
        RECT 2414.110 1789.580 2414.460 1789.610 ;
        RECT 2413.200 1789.550 2414.460 1789.580 ;
        RECT 2413.140 1789.410 2414.460 1789.550 ;
        RECT 2407.525 1789.320 2407.815 1789.345 ;
        RECT 2413.140 1789.320 2413.430 1789.410 ;
        RECT 2414.110 1789.320 2414.460 1789.410 ;
        RECT 2400.710 1788.950 2401.065 1789.305 ;
        RECT 2408.155 1789.180 2408.505 1789.255 ;
        RECT 2413.595 1789.180 2413.920 1789.270 ;
        RECT 2407.955 1789.150 2408.505 1789.180 ;
        RECT 2413.570 1789.150 2413.920 1789.180 ;
        RECT 2407.785 1789.145 2408.505 1789.150 ;
        RECT 2413.400 1789.145 2413.920 1789.150 ;
        RECT 2407.785 1788.980 2413.920 1789.145 ;
        RECT 2407.845 1788.975 2413.920 1788.980 ;
        RECT 2407.955 1788.950 2408.505 1788.975 ;
        RECT 2413.570 1788.950 2413.920 1788.975 ;
        RECT 2400.710 1788.930 2401.010 1788.950 ;
        RECT 2399.670 1788.925 2399.900 1788.930 ;
        RECT 2385.400 1788.690 2385.690 1788.865 ;
        RECT 2397.535 1788.820 2397.855 1788.835 ;
        RECT 2397.510 1788.790 2397.855 1788.820 ;
        RECT 2397.335 1788.620 2397.855 1788.790 ;
        RECT 2399.670 1788.690 2399.960 1788.925 ;
        RECT 2400.660 1788.860 2401.010 1788.930 ;
        RECT 2408.155 1788.905 2408.505 1788.950 ;
        RECT 2413.595 1788.945 2413.920 1788.950 ;
        RECT 2414.990 1788.930 2415.160 1790.030 ;
        RECT 2415.980 1789.300 2416.150 1790.030 ;
        RECT 2422.845 1789.715 2423.015 1790.060 ;
        RECT 2422.745 1789.345 2423.115 1789.715 ;
        RECT 2428.460 1789.580 2428.630 1790.060 ;
        RECT 2430.190 1790.030 2430.485 1790.290 ;
        RECT 2431.180 1790.030 2431.475 1790.290 ;
        RECT 2438.045 1790.060 2438.335 1790.290 ;
        RECT 2443.660 1790.060 2443.950 1790.290 ;
        RECT 2429.370 1789.580 2429.720 1789.610 ;
        RECT 2428.460 1789.550 2429.720 1789.580 ;
        RECT 2428.400 1789.410 2429.720 1789.550 ;
        RECT 2422.785 1789.320 2423.075 1789.345 ;
        RECT 2428.400 1789.320 2428.690 1789.410 ;
        RECT 2429.370 1789.320 2429.720 1789.410 ;
        RECT 2415.930 1788.950 2416.280 1789.300 ;
        RECT 2423.420 1789.180 2423.770 1789.255 ;
        RECT 2428.855 1789.180 2429.180 1789.270 ;
        RECT 2423.215 1789.150 2423.770 1789.180 ;
        RECT 2428.830 1789.150 2429.180 1789.180 ;
        RECT 2423.045 1789.145 2423.770 1789.150 ;
        RECT 2428.660 1789.145 2429.180 1789.150 ;
        RECT 2423.045 1788.980 2429.180 1789.145 ;
        RECT 2423.105 1788.975 2429.180 1788.980 ;
        RECT 2423.215 1788.950 2423.770 1788.975 ;
        RECT 2428.830 1788.950 2429.180 1788.975 ;
        RECT 2415.930 1788.930 2416.270 1788.950 ;
        RECT 2414.930 1788.925 2415.160 1788.930 ;
        RECT 2400.660 1788.690 2400.950 1788.860 ;
        RECT 2412.795 1788.820 2413.115 1788.835 ;
        RECT 2412.770 1788.790 2413.115 1788.820 ;
        RECT 2412.595 1788.620 2413.115 1788.790 ;
        RECT 2414.930 1788.690 2415.220 1788.925 ;
        RECT 2415.920 1788.860 2416.270 1788.930 ;
        RECT 2423.420 1788.905 2423.770 1788.950 ;
        RECT 2428.855 1788.945 2429.180 1788.950 ;
        RECT 2430.250 1788.930 2430.420 1790.030 ;
        RECT 2431.240 1789.300 2431.410 1790.030 ;
        RECT 2438.105 1789.715 2438.275 1790.060 ;
        RECT 2438.005 1789.345 2438.375 1789.715 ;
        RECT 2443.720 1789.580 2443.890 1790.060 ;
        RECT 2445.450 1790.030 2445.745 1790.290 ;
        RECT 2446.440 1790.030 2446.735 1790.290 ;
        RECT 2699.360 1790.225 2699.500 1790.720 ;
        RECT 2699.730 1790.720 2700.880 1790.860 ;
        RECT 2699.730 1790.660 2700.050 1790.720 ;
        RECT 2444.630 1789.580 2444.980 1789.610 ;
        RECT 2443.720 1789.550 2444.980 1789.580 ;
        RECT 2443.660 1789.410 2444.980 1789.550 ;
        RECT 2438.045 1789.320 2438.335 1789.345 ;
        RECT 2443.660 1789.320 2443.950 1789.410 ;
        RECT 2444.630 1789.320 2444.980 1789.410 ;
        RECT 2431.190 1788.950 2431.540 1789.300 ;
        RECT 2438.675 1789.180 2439.025 1789.255 ;
        RECT 2444.115 1789.180 2444.440 1789.270 ;
        RECT 2438.475 1789.150 2439.025 1789.180 ;
        RECT 2444.090 1789.150 2444.440 1789.180 ;
        RECT 2438.305 1789.145 2439.025 1789.150 ;
        RECT 2443.920 1789.145 2444.440 1789.150 ;
        RECT 2438.305 1788.980 2444.440 1789.145 ;
        RECT 2438.365 1788.975 2444.440 1788.980 ;
        RECT 2438.475 1788.950 2439.025 1788.975 ;
        RECT 2444.090 1788.950 2444.440 1788.975 ;
        RECT 2431.190 1788.930 2431.530 1788.950 ;
        RECT 2430.190 1788.925 2430.420 1788.930 ;
        RECT 2415.920 1788.690 2416.210 1788.860 ;
        RECT 2428.055 1788.820 2428.375 1788.835 ;
        RECT 2428.030 1788.790 2428.375 1788.820 ;
        RECT 2427.855 1788.620 2428.375 1788.790 ;
        RECT 2430.190 1788.690 2430.480 1788.925 ;
        RECT 2431.180 1788.860 2431.530 1788.930 ;
        RECT 2438.675 1788.905 2439.025 1788.950 ;
        RECT 2444.115 1788.945 2444.440 1788.950 ;
        RECT 2445.510 1788.930 2445.680 1790.030 ;
        RECT 2446.475 1789.995 2446.735 1790.030 ;
        RECT 2699.285 1789.995 2699.575 1790.225 ;
        RECT 2446.475 1789.915 2446.795 1789.995 ;
        RECT 2446.475 1789.565 2446.825 1789.915 ;
        RECT 2446.500 1788.930 2446.670 1789.565 ;
        RECT 2696.970 1789.500 2697.290 1789.560 ;
        RECT 2698.365 1789.500 2698.655 1789.545 ;
        RECT 2696.970 1789.360 2698.655 1789.500 ;
        RECT 2699.360 1789.500 2699.500 1789.995 ;
        RECT 2700.740 1789.885 2700.880 1790.720 ;
        RECT 2702.030 1790.320 2702.350 1790.580 ;
        RECT 2702.490 1790.320 2702.810 1790.580 ;
        RECT 2702.965 1790.335 2703.255 1790.565 ;
        RECT 2703.040 1790.180 2703.180 1790.335 ;
        RECT 2702.580 1790.040 2703.180 1790.180 ;
        RECT 2700.665 1789.655 2700.955 1789.885 ;
        RECT 2702.580 1789.500 2702.720 1790.040 ;
        RECT 2699.360 1789.360 2702.720 1789.500 ;
        RECT 2696.970 1789.300 2697.290 1789.360 ;
        RECT 2698.365 1789.315 2698.655 1789.360 ;
        RECT 2445.450 1788.925 2445.680 1788.930 ;
        RECT 2446.440 1788.925 2446.670 1788.930 ;
        RECT 2431.180 1788.690 2431.470 1788.860 ;
        RECT 2443.315 1788.820 2443.635 1788.835 ;
        RECT 2443.290 1788.790 2443.635 1788.820 ;
        RECT 2443.115 1788.620 2443.635 1788.790 ;
        RECT 2445.450 1788.690 2445.740 1788.925 ;
        RECT 2446.440 1788.690 2446.730 1788.925 ;
        RECT 2369.085 1788.575 2369.435 1788.620 ;
        RECT 2382.250 1788.590 2382.595 1788.620 ;
        RECT 2397.510 1788.590 2397.855 1788.620 ;
        RECT 2412.770 1788.590 2413.115 1788.620 ;
        RECT 2428.030 1788.590 2428.375 1788.620 ;
        RECT 2443.290 1788.590 2443.635 1788.620 ;
        RECT 2382.275 1788.545 2382.595 1788.590 ;
        RECT 2397.535 1788.545 2397.855 1788.590 ;
        RECT 2412.795 1788.545 2413.115 1788.590 ;
        RECT 2428.055 1788.545 2428.375 1788.590 ;
        RECT 2443.315 1788.545 2443.635 1788.590 ;
        RECT 2697.905 1788.480 2698.195 1788.525 ;
        RECT 2698.350 1788.480 2698.670 1788.540 ;
        RECT 2697.905 1788.340 2698.670 1788.480 ;
        RECT 2697.905 1788.295 2698.195 1788.340 ;
        RECT 2698.350 1788.280 2698.670 1788.340 ;
        RECT 2698.810 1788.480 2699.130 1788.540 ;
        RECT 2699.285 1788.480 2699.575 1788.525 ;
        RECT 2698.810 1788.340 2699.575 1788.480 ;
        RECT 2698.810 1788.280 2699.130 1788.340 ;
        RECT 2699.285 1788.295 2699.575 1788.340 ;
        RECT 2694.670 1787.460 2694.990 1787.520 ;
        RECT 2696.985 1787.460 2697.275 1787.505 ;
        RECT 2694.670 1787.320 2697.275 1787.460 ;
        RECT 2694.670 1787.260 2694.990 1787.320 ;
        RECT 2696.985 1787.275 2697.275 1787.320 ;
        RECT 2697.430 1787.460 2697.750 1787.520 ;
        RECT 2698.825 1787.460 2699.115 1787.505 ;
        RECT 2697.430 1787.320 2699.115 1787.460 ;
        RECT 2697.430 1787.260 2697.750 1787.320 ;
        RECT 2698.825 1787.275 2699.115 1787.320 ;
        RECT 2699.730 1787.260 2700.050 1787.520 ;
        RECT 2523.545 1786.325 2523.865 1786.585 ;
        RECT 2699.730 1785.760 2700.050 1785.820 ;
        RECT 2700.665 1785.760 2700.955 1785.805 ;
        RECT 2699.730 1785.620 2700.955 1785.760 ;
        RECT 2699.730 1785.560 2700.050 1785.620 ;
        RECT 2700.665 1785.575 2700.955 1785.620 ;
        RECT 2373.665 1784.895 2373.955 1785.105 ;
        RECT 2372.775 1784.875 2373.955 1784.895 ;
        RECT 2371.755 1784.585 2372.075 1784.845 ;
        RECT 2372.775 1784.825 2373.875 1784.875 ;
        RECT 2374.605 1784.865 2374.925 1785.125 ;
        RECT 2375.205 1785.105 2375.525 1785.125 ;
        RECT 2375.105 1784.875 2375.525 1785.105 ;
        RECT 2375.205 1784.865 2375.525 1784.875 ;
        RECT 2376.765 1785.105 2377.100 1785.125 ;
        RECT 2376.765 1784.875 2377.290 1785.105 ;
        RECT 2378.945 1785.065 2379.235 1785.105 ;
        RECT 2379.375 1785.065 2379.695 1785.125 ;
        RECT 2378.945 1784.925 2379.695 1785.065 ;
        RECT 2378.945 1784.875 2379.235 1784.925 ;
        RECT 2376.765 1784.865 2377.100 1784.875 ;
        RECT 2379.375 1784.865 2379.695 1784.925 ;
        RECT 2388.925 1784.895 2389.215 1785.105 ;
        RECT 2388.035 1784.875 2389.215 1784.895 ;
        RECT 2372.705 1784.755 2373.875 1784.825 ;
        RECT 2372.705 1784.595 2372.995 1784.755 ;
        RECT 2375.135 1784.585 2375.305 1784.685 ;
        RECT 2377.515 1784.585 2377.835 1784.845 ;
        RECT 2387.015 1784.585 2387.335 1784.845 ;
        RECT 2388.035 1784.825 2389.135 1784.875 ;
        RECT 2389.865 1784.865 2390.185 1785.125 ;
        RECT 2390.465 1785.105 2390.785 1785.125 ;
        RECT 2390.365 1784.875 2390.785 1785.105 ;
        RECT 2390.465 1784.865 2390.785 1784.875 ;
        RECT 2392.025 1785.105 2392.360 1785.125 ;
        RECT 2392.025 1784.875 2392.550 1785.105 ;
        RECT 2394.205 1785.065 2394.495 1785.105 ;
        RECT 2394.635 1785.065 2394.955 1785.125 ;
        RECT 2394.205 1784.925 2394.955 1785.065 ;
        RECT 2394.205 1784.875 2394.495 1784.925 ;
        RECT 2392.025 1784.865 2392.360 1784.875 ;
        RECT 2394.635 1784.865 2394.955 1784.925 ;
        RECT 2404.185 1784.895 2404.475 1785.105 ;
        RECT 2403.295 1784.875 2404.475 1784.895 ;
        RECT 2387.965 1784.755 2389.135 1784.825 ;
        RECT 2387.965 1784.595 2388.255 1784.755 ;
        RECT 2390.395 1784.585 2390.565 1784.685 ;
        RECT 2392.775 1784.585 2393.095 1784.845 ;
        RECT 2402.275 1784.585 2402.595 1784.845 ;
        RECT 2403.295 1784.825 2404.395 1784.875 ;
        RECT 2405.125 1784.865 2405.445 1785.125 ;
        RECT 2405.725 1785.105 2406.045 1785.125 ;
        RECT 2405.625 1784.875 2406.045 1785.105 ;
        RECT 2405.725 1784.865 2406.045 1784.875 ;
        RECT 2407.285 1785.105 2407.620 1785.125 ;
        RECT 2407.285 1784.875 2407.810 1785.105 ;
        RECT 2409.465 1785.065 2409.755 1785.105 ;
        RECT 2409.895 1785.065 2410.215 1785.125 ;
        RECT 2409.465 1784.925 2410.215 1785.065 ;
        RECT 2409.465 1784.875 2409.755 1784.925 ;
        RECT 2407.285 1784.865 2407.620 1784.875 ;
        RECT 2409.895 1784.865 2410.215 1784.925 ;
        RECT 2419.445 1784.895 2419.735 1785.105 ;
        RECT 2418.555 1784.875 2419.735 1784.895 ;
        RECT 2403.225 1784.755 2404.395 1784.825 ;
        RECT 2403.225 1784.595 2403.515 1784.755 ;
        RECT 2405.655 1784.585 2405.825 1784.685 ;
        RECT 2408.035 1784.585 2408.355 1784.845 ;
        RECT 2417.535 1784.585 2417.855 1784.845 ;
        RECT 2418.555 1784.825 2419.655 1784.875 ;
        RECT 2420.385 1784.865 2420.705 1785.125 ;
        RECT 2420.985 1785.105 2421.305 1785.125 ;
        RECT 2420.885 1784.875 2421.305 1785.105 ;
        RECT 2420.985 1784.865 2421.305 1784.875 ;
        RECT 2422.545 1785.105 2422.880 1785.125 ;
        RECT 2422.545 1784.875 2423.070 1785.105 ;
        RECT 2424.725 1785.065 2425.015 1785.105 ;
        RECT 2425.155 1785.065 2425.475 1785.125 ;
        RECT 2424.725 1784.925 2425.475 1785.065 ;
        RECT 2424.725 1784.875 2425.015 1784.925 ;
        RECT 2422.545 1784.865 2422.880 1784.875 ;
        RECT 2425.155 1784.865 2425.475 1784.925 ;
        RECT 2434.705 1784.895 2434.995 1785.105 ;
        RECT 2433.815 1784.875 2434.995 1784.895 ;
        RECT 2418.485 1784.755 2419.655 1784.825 ;
        RECT 2418.485 1784.595 2418.775 1784.755 ;
        RECT 2420.915 1784.585 2421.085 1784.685 ;
        RECT 2423.295 1784.585 2423.615 1784.845 ;
        RECT 2432.795 1784.585 2433.115 1784.845 ;
        RECT 2433.815 1784.825 2434.915 1784.875 ;
        RECT 2435.645 1784.865 2435.965 1785.125 ;
        RECT 2436.245 1785.105 2436.565 1785.125 ;
        RECT 2436.145 1784.875 2436.565 1785.105 ;
        RECT 2436.245 1784.865 2436.565 1784.875 ;
        RECT 2437.805 1785.105 2438.140 1785.125 ;
        RECT 2437.805 1784.875 2438.330 1785.105 ;
        RECT 2439.985 1785.065 2440.275 1785.105 ;
        RECT 2440.415 1785.065 2440.735 1785.125 ;
        RECT 2439.985 1784.925 2440.735 1785.065 ;
        RECT 2439.985 1784.875 2440.275 1784.925 ;
        RECT 2437.805 1784.865 2438.140 1784.875 ;
        RECT 2440.415 1784.865 2440.735 1784.925 ;
        RECT 2698.810 1784.880 2699.130 1785.140 ;
        RECT 2433.745 1784.755 2434.915 1784.825 ;
        RECT 2433.745 1784.595 2434.035 1784.755 ;
        RECT 2436.175 1784.585 2436.345 1784.685 ;
        RECT 2438.555 1784.585 2438.875 1784.845 ;
        RECT 2696.970 1784.740 2697.290 1784.800 ;
        RECT 2697.445 1784.740 2697.735 1784.785 ;
        RECT 2696.970 1784.600 2697.735 1784.740 ;
        RECT 2374.125 1784.545 2374.445 1784.565 ;
        RECT 2373.185 1784.505 2373.475 1784.545 ;
        RECT 2373.185 1784.315 2373.635 1784.505 ;
        RECT 2372.445 1784.025 2372.765 1784.285 ;
        RECT 2372.925 1783.745 2373.245 1784.005 ;
        RECT 2373.495 1783.985 2373.635 1784.315 ;
        RECT 2374.125 1784.315 2374.675 1784.545 ;
        RECT 2374.815 1784.445 2376.995 1784.585 ;
        RECT 2389.385 1784.545 2389.705 1784.565 ;
        RECT 2374.815 1784.365 2376.115 1784.445 ;
        RECT 2374.125 1784.305 2374.445 1784.315 ;
        RECT 2374.815 1784.085 2375.155 1784.365 ;
        RECT 2375.825 1784.315 2376.115 1784.365 ;
        RECT 2374.865 1784.035 2375.155 1784.085 ;
        RECT 2376.285 1784.025 2376.605 1784.285 ;
        RECT 2373.495 1783.845 2373.755 1783.985 ;
        RECT 2371.755 1783.185 2372.075 1783.445 ;
        RECT 2373.615 1783.425 2373.755 1783.845 ;
        RECT 2373.905 1783.945 2374.195 1783.985 ;
        RECT 2374.365 1783.945 2374.685 1784.005 ;
        RECT 2373.905 1783.805 2374.685 1783.945 ;
        RECT 2373.905 1783.755 2374.195 1783.805 ;
        RECT 2374.365 1783.745 2374.685 1783.805 ;
        RECT 2375.345 1783.755 2375.635 1783.985 ;
        RECT 2375.495 1783.505 2375.635 1783.755 ;
        RECT 2375.805 1783.745 2376.125 1784.005 ;
        RECT 2376.855 1783.805 2376.995 1784.445 ;
        RECT 2378.705 1784.505 2378.995 1784.545 ;
        RECT 2388.445 1784.505 2388.735 1784.545 ;
        RECT 2378.705 1784.365 2379.275 1784.505 ;
        RECT 2377.335 1784.285 2378.435 1784.365 ;
        RECT 2378.705 1784.315 2378.995 1784.365 ;
        RECT 2377.145 1784.265 2378.435 1784.285 ;
        RECT 2379.135 1784.265 2379.395 1784.365 ;
        RECT 2377.145 1784.225 2378.515 1784.265 ;
        RECT 2379.135 1784.225 2379.475 1784.265 ;
        RECT 2377.145 1784.035 2377.555 1784.225 ;
        RECT 2378.225 1784.035 2378.515 1784.225 ;
        RECT 2379.185 1784.035 2379.475 1784.225 ;
        RECT 2377.145 1784.025 2377.465 1784.035 ;
        RECT 2377.745 1783.805 2378.035 1783.985 ;
        RECT 2376.855 1783.755 2378.035 1783.805 ;
        RECT 2376.855 1783.705 2377.955 1783.755 ;
        RECT 2378.685 1783.745 2379.005 1784.005 ;
        RECT 2380.670 1783.995 2381.010 1784.345 ;
        RECT 2388.445 1784.315 2388.895 1784.505 ;
        RECT 2385.170 1784.265 2385.490 1784.280 ;
        RECT 2385.170 1784.035 2385.685 1784.265 ;
        RECT 2385.170 1784.020 2385.490 1784.035 ;
        RECT 2387.705 1784.025 2388.025 1784.285 ;
        RECT 2376.785 1783.665 2377.955 1783.705 ;
        RECT 2375.495 1783.445 2375.795 1783.505 ;
        RECT 2376.785 1783.455 2377.075 1783.665 ;
        RECT 2380.760 1783.490 2380.930 1783.995 ;
        RECT 2382.275 1783.875 2382.595 1783.980 ;
        RECT 2382.250 1783.860 2382.595 1783.875 ;
        RECT 2382.240 1783.845 2382.595 1783.860 ;
        RECT 2382.075 1783.675 2382.595 1783.845 ;
        RECT 2382.250 1783.660 2382.595 1783.675 ;
        RECT 2382.250 1783.645 2382.540 1783.660 ;
        RECT 2383.050 1783.490 2383.400 1783.610 ;
        RECT 2384.410 1783.540 2384.700 1783.775 ;
        RECT 2385.395 1783.540 2385.685 1783.775 ;
        RECT 2388.185 1783.745 2388.505 1784.005 ;
        RECT 2388.755 1783.985 2388.895 1784.315 ;
        RECT 2389.385 1784.315 2389.935 1784.545 ;
        RECT 2390.075 1784.445 2392.255 1784.585 ;
        RECT 2404.645 1784.545 2404.965 1784.565 ;
        RECT 2390.075 1784.365 2391.375 1784.445 ;
        RECT 2389.385 1784.305 2389.705 1784.315 ;
        RECT 2390.075 1784.085 2390.415 1784.365 ;
        RECT 2391.085 1784.315 2391.375 1784.365 ;
        RECT 2390.125 1784.035 2390.415 1784.085 ;
        RECT 2391.545 1784.025 2391.865 1784.285 ;
        RECT 2388.755 1783.845 2389.015 1783.985 ;
        RECT 2384.410 1783.535 2384.640 1783.540 ;
        RECT 2385.395 1783.535 2385.625 1783.540 ;
        RECT 2373.615 1783.385 2373.955 1783.425 ;
        RECT 2374.485 1783.385 2374.805 1783.445 ;
        RECT 2373.615 1783.245 2374.805 1783.385 ;
        RECT 2373.665 1783.195 2373.955 1783.245 ;
        RECT 2374.485 1783.185 2374.805 1783.245 ;
        RECT 2374.955 1783.185 2375.355 1783.445 ;
        RECT 2375.495 1783.385 2375.885 1783.445 ;
        RECT 2376.285 1783.425 2376.605 1783.445 ;
        RECT 2376.065 1783.385 2376.605 1783.425 ;
        RECT 2375.495 1783.365 2376.605 1783.385 ;
        RECT 2375.565 1783.245 2376.605 1783.365 ;
        RECT 2375.565 1783.185 2375.885 1783.245 ;
        RECT 2376.065 1783.195 2376.605 1783.245 ;
        RECT 2376.285 1783.185 2376.605 1783.195 ;
        RECT 2377.515 1783.385 2377.835 1783.445 ;
        RECT 2377.985 1783.385 2378.275 1783.425 ;
        RECT 2377.515 1783.245 2378.275 1783.385 ;
        RECT 2377.515 1783.185 2377.835 1783.245 ;
        RECT 2377.985 1783.195 2378.275 1783.245 ;
        RECT 2378.945 1783.385 2379.235 1783.425 ;
        RECT 2379.375 1783.385 2379.695 1783.445 ;
        RECT 2378.945 1783.245 2379.695 1783.385 ;
        RECT 2380.760 1783.320 2383.400 1783.490 ;
        RECT 2382.880 1783.315 2383.400 1783.320 ;
        RECT 2383.050 1783.260 2383.400 1783.315 ;
        RECT 2378.945 1783.195 2379.235 1783.245 ;
        RECT 2379.375 1783.185 2379.695 1783.245 ;
        RECT 2382.620 1783.120 2382.910 1783.145 ;
        RECT 2383.590 1783.120 2383.940 1783.145 ;
        RECT 2382.620 1782.950 2383.940 1783.120 ;
        RECT 2382.620 1782.915 2382.910 1782.950 ;
        RECT 2382.680 1782.405 2382.850 1782.915 ;
        RECT 2383.590 1782.855 2383.940 1782.950 ;
        RECT 2384.470 1782.435 2384.640 1783.535 ;
        RECT 2385.455 1782.435 2385.625 1783.535 ;
        RECT 2387.015 1783.185 2387.335 1783.445 ;
        RECT 2388.875 1783.425 2389.015 1783.845 ;
        RECT 2389.165 1783.945 2389.455 1783.985 ;
        RECT 2389.625 1783.945 2389.945 1784.005 ;
        RECT 2389.165 1783.805 2389.945 1783.945 ;
        RECT 2389.165 1783.755 2389.455 1783.805 ;
        RECT 2389.625 1783.745 2389.945 1783.805 ;
        RECT 2390.605 1783.755 2390.895 1783.985 ;
        RECT 2390.755 1783.505 2390.895 1783.755 ;
        RECT 2391.065 1783.745 2391.385 1784.005 ;
        RECT 2392.115 1783.805 2392.255 1784.445 ;
        RECT 2393.965 1784.505 2394.255 1784.545 ;
        RECT 2403.705 1784.505 2403.995 1784.545 ;
        RECT 2393.965 1784.365 2394.535 1784.505 ;
        RECT 2392.595 1784.285 2393.695 1784.365 ;
        RECT 2393.965 1784.315 2394.255 1784.365 ;
        RECT 2392.405 1784.265 2393.695 1784.285 ;
        RECT 2394.395 1784.265 2394.655 1784.365 ;
        RECT 2392.405 1784.225 2393.775 1784.265 ;
        RECT 2394.395 1784.225 2394.735 1784.265 ;
        RECT 2392.405 1784.035 2392.815 1784.225 ;
        RECT 2393.485 1784.035 2393.775 1784.225 ;
        RECT 2394.445 1784.035 2394.735 1784.225 ;
        RECT 2392.405 1784.025 2392.725 1784.035 ;
        RECT 2393.005 1783.805 2393.295 1783.985 ;
        RECT 2392.115 1783.755 2393.295 1783.805 ;
        RECT 2392.115 1783.705 2393.215 1783.755 ;
        RECT 2393.945 1783.745 2394.265 1784.005 ;
        RECT 2395.930 1783.995 2396.270 1784.345 ;
        RECT 2403.705 1784.315 2404.155 1784.505 ;
        RECT 2400.810 1784.265 2401.130 1784.280 ;
        RECT 2400.655 1784.035 2401.130 1784.265 ;
        RECT 2400.810 1784.020 2401.130 1784.035 ;
        RECT 2402.965 1784.025 2403.285 1784.285 ;
        RECT 2392.045 1783.665 2393.215 1783.705 ;
        RECT 2390.755 1783.445 2391.055 1783.505 ;
        RECT 2392.045 1783.455 2392.335 1783.665 ;
        RECT 2396.020 1783.490 2396.190 1783.995 ;
        RECT 2397.535 1783.875 2397.855 1783.980 ;
        RECT 2397.510 1783.860 2397.855 1783.875 ;
        RECT 2397.500 1783.845 2397.855 1783.860 ;
        RECT 2397.335 1783.675 2397.855 1783.845 ;
        RECT 2397.510 1783.660 2397.855 1783.675 ;
        RECT 2397.510 1783.645 2397.800 1783.660 ;
        RECT 2398.310 1783.490 2398.660 1783.610 ;
        RECT 2399.670 1783.540 2399.960 1783.775 ;
        RECT 2400.655 1783.540 2400.945 1783.775 ;
        RECT 2403.445 1783.745 2403.765 1784.005 ;
        RECT 2404.015 1783.985 2404.155 1784.315 ;
        RECT 2404.645 1784.315 2405.195 1784.545 ;
        RECT 2405.335 1784.445 2407.515 1784.585 ;
        RECT 2419.905 1784.545 2420.225 1784.565 ;
        RECT 2405.335 1784.365 2406.635 1784.445 ;
        RECT 2404.645 1784.305 2404.965 1784.315 ;
        RECT 2405.335 1784.085 2405.675 1784.365 ;
        RECT 2406.345 1784.315 2406.635 1784.365 ;
        RECT 2405.385 1784.035 2405.675 1784.085 ;
        RECT 2406.805 1784.025 2407.125 1784.285 ;
        RECT 2404.015 1783.845 2404.275 1783.985 ;
        RECT 2399.670 1783.535 2399.900 1783.540 ;
        RECT 2400.655 1783.535 2400.885 1783.540 ;
        RECT 2388.875 1783.385 2389.215 1783.425 ;
        RECT 2389.745 1783.385 2390.065 1783.445 ;
        RECT 2388.875 1783.245 2390.065 1783.385 ;
        RECT 2388.925 1783.195 2389.215 1783.245 ;
        RECT 2389.745 1783.185 2390.065 1783.245 ;
        RECT 2390.215 1783.185 2390.615 1783.445 ;
        RECT 2390.755 1783.385 2391.145 1783.445 ;
        RECT 2391.545 1783.425 2391.865 1783.445 ;
        RECT 2391.325 1783.385 2391.865 1783.425 ;
        RECT 2390.755 1783.365 2391.865 1783.385 ;
        RECT 2390.825 1783.245 2391.865 1783.365 ;
        RECT 2390.825 1783.185 2391.145 1783.245 ;
        RECT 2391.325 1783.195 2391.865 1783.245 ;
        RECT 2391.545 1783.185 2391.865 1783.195 ;
        RECT 2392.775 1783.385 2393.095 1783.445 ;
        RECT 2393.245 1783.385 2393.535 1783.425 ;
        RECT 2392.775 1783.245 2393.535 1783.385 ;
        RECT 2392.775 1783.185 2393.095 1783.245 ;
        RECT 2393.245 1783.195 2393.535 1783.245 ;
        RECT 2394.205 1783.385 2394.495 1783.425 ;
        RECT 2394.635 1783.385 2394.955 1783.445 ;
        RECT 2394.205 1783.245 2394.955 1783.385 ;
        RECT 2396.020 1783.320 2398.660 1783.490 ;
        RECT 2398.140 1783.315 2398.660 1783.320 ;
        RECT 2398.310 1783.260 2398.660 1783.315 ;
        RECT 2394.205 1783.195 2394.495 1783.245 ;
        RECT 2394.635 1783.185 2394.955 1783.245 ;
        RECT 2397.880 1783.120 2398.170 1783.145 ;
        RECT 2398.850 1783.120 2399.200 1783.145 ;
        RECT 2397.880 1782.950 2399.200 1783.120 ;
        RECT 2397.880 1782.915 2398.170 1782.950 ;
        RECT 2382.620 1782.175 2382.910 1782.405 ;
        RECT 2384.410 1782.175 2384.705 1782.435 ;
        RECT 2385.395 1782.175 2385.690 1782.435 ;
        RECT 2397.940 1782.405 2398.110 1782.915 ;
        RECT 2398.850 1782.855 2399.200 1782.950 ;
        RECT 2399.730 1782.435 2399.900 1783.535 ;
        RECT 2400.715 1782.435 2400.885 1783.535 ;
        RECT 2402.275 1783.185 2402.595 1783.445 ;
        RECT 2404.135 1783.425 2404.275 1783.845 ;
        RECT 2404.425 1783.945 2404.715 1783.985 ;
        RECT 2404.885 1783.945 2405.205 1784.005 ;
        RECT 2404.425 1783.805 2405.205 1783.945 ;
        RECT 2404.425 1783.755 2404.715 1783.805 ;
        RECT 2404.885 1783.745 2405.205 1783.805 ;
        RECT 2405.865 1783.755 2406.155 1783.985 ;
        RECT 2406.015 1783.505 2406.155 1783.755 ;
        RECT 2406.325 1783.745 2406.645 1784.005 ;
        RECT 2407.375 1783.805 2407.515 1784.445 ;
        RECT 2409.225 1784.505 2409.515 1784.545 ;
        RECT 2418.965 1784.505 2419.255 1784.545 ;
        RECT 2409.225 1784.365 2409.795 1784.505 ;
        RECT 2407.855 1784.285 2408.955 1784.365 ;
        RECT 2409.225 1784.315 2409.515 1784.365 ;
        RECT 2407.665 1784.265 2408.955 1784.285 ;
        RECT 2409.655 1784.265 2409.915 1784.365 ;
        RECT 2407.665 1784.225 2409.035 1784.265 ;
        RECT 2409.655 1784.225 2409.995 1784.265 ;
        RECT 2407.665 1784.035 2408.075 1784.225 ;
        RECT 2408.745 1784.035 2409.035 1784.225 ;
        RECT 2409.705 1784.035 2409.995 1784.225 ;
        RECT 2407.665 1784.025 2407.985 1784.035 ;
        RECT 2408.265 1783.805 2408.555 1783.985 ;
        RECT 2407.375 1783.755 2408.555 1783.805 ;
        RECT 2407.375 1783.705 2408.475 1783.755 ;
        RECT 2409.205 1783.745 2409.525 1784.005 ;
        RECT 2411.190 1783.995 2411.530 1784.345 ;
        RECT 2418.965 1784.315 2419.415 1784.505 ;
        RECT 2418.225 1784.025 2418.545 1784.285 ;
        RECT 2407.305 1783.665 2408.475 1783.705 ;
        RECT 2406.015 1783.445 2406.315 1783.505 ;
        RECT 2407.305 1783.455 2407.595 1783.665 ;
        RECT 2411.280 1783.490 2411.450 1783.995 ;
        RECT 2412.795 1783.875 2413.115 1783.980 ;
        RECT 2412.770 1783.860 2413.115 1783.875 ;
        RECT 2412.760 1783.845 2413.115 1783.860 ;
        RECT 2412.595 1783.675 2413.115 1783.845 ;
        RECT 2412.770 1783.660 2413.115 1783.675 ;
        RECT 2412.770 1783.645 2413.060 1783.660 ;
        RECT 2413.570 1783.490 2413.920 1783.610 ;
        RECT 2414.930 1783.540 2415.220 1783.775 ;
        RECT 2415.915 1783.540 2416.205 1783.775 ;
        RECT 2418.705 1783.745 2419.025 1784.005 ;
        RECT 2419.275 1783.985 2419.415 1784.315 ;
        RECT 2419.905 1784.315 2420.455 1784.545 ;
        RECT 2420.595 1784.445 2422.775 1784.585 ;
        RECT 2435.165 1784.545 2435.485 1784.565 ;
        RECT 2420.595 1784.365 2421.895 1784.445 ;
        RECT 2419.905 1784.305 2420.225 1784.315 ;
        RECT 2420.595 1784.085 2420.935 1784.365 ;
        RECT 2421.605 1784.315 2421.895 1784.365 ;
        RECT 2420.645 1784.035 2420.935 1784.085 ;
        RECT 2422.065 1784.025 2422.385 1784.285 ;
        RECT 2419.275 1783.845 2419.535 1783.985 ;
        RECT 2414.930 1783.535 2415.160 1783.540 ;
        RECT 2415.915 1783.535 2416.145 1783.540 ;
        RECT 2404.135 1783.385 2404.475 1783.425 ;
        RECT 2405.005 1783.385 2405.325 1783.445 ;
        RECT 2404.135 1783.245 2405.325 1783.385 ;
        RECT 2404.185 1783.195 2404.475 1783.245 ;
        RECT 2405.005 1783.185 2405.325 1783.245 ;
        RECT 2405.475 1783.185 2405.875 1783.445 ;
        RECT 2406.015 1783.385 2406.405 1783.445 ;
        RECT 2406.805 1783.425 2407.125 1783.445 ;
        RECT 2406.585 1783.385 2407.125 1783.425 ;
        RECT 2406.015 1783.365 2407.125 1783.385 ;
        RECT 2406.085 1783.245 2407.125 1783.365 ;
        RECT 2406.085 1783.185 2406.405 1783.245 ;
        RECT 2406.585 1783.195 2407.125 1783.245 ;
        RECT 2406.805 1783.185 2407.125 1783.195 ;
        RECT 2408.035 1783.385 2408.355 1783.445 ;
        RECT 2408.505 1783.385 2408.795 1783.425 ;
        RECT 2408.035 1783.245 2408.795 1783.385 ;
        RECT 2408.035 1783.185 2408.355 1783.245 ;
        RECT 2408.505 1783.195 2408.795 1783.245 ;
        RECT 2409.465 1783.385 2409.755 1783.425 ;
        RECT 2409.895 1783.385 2410.215 1783.445 ;
        RECT 2409.465 1783.245 2410.215 1783.385 ;
        RECT 2411.280 1783.320 2413.920 1783.490 ;
        RECT 2413.400 1783.315 2413.920 1783.320 ;
        RECT 2413.570 1783.260 2413.920 1783.315 ;
        RECT 2409.465 1783.195 2409.755 1783.245 ;
        RECT 2409.895 1783.185 2410.215 1783.245 ;
        RECT 2413.140 1783.120 2413.430 1783.145 ;
        RECT 2414.110 1783.120 2414.460 1783.145 ;
        RECT 2413.140 1782.950 2414.460 1783.120 ;
        RECT 2413.140 1782.915 2413.430 1782.950 ;
        RECT 2397.880 1782.175 2398.170 1782.405 ;
        RECT 2399.670 1782.175 2399.965 1782.435 ;
        RECT 2400.655 1782.175 2400.950 1782.435 ;
        RECT 2413.200 1782.405 2413.370 1782.915 ;
        RECT 2414.110 1782.855 2414.460 1782.950 ;
        RECT 2414.990 1782.435 2415.160 1783.535 ;
        RECT 2415.975 1782.435 2416.145 1783.535 ;
        RECT 2417.535 1783.185 2417.855 1783.445 ;
        RECT 2419.395 1783.425 2419.535 1783.845 ;
        RECT 2419.685 1783.945 2419.975 1783.985 ;
        RECT 2420.145 1783.945 2420.465 1784.005 ;
        RECT 2419.685 1783.805 2420.465 1783.945 ;
        RECT 2419.685 1783.755 2419.975 1783.805 ;
        RECT 2420.145 1783.745 2420.465 1783.805 ;
        RECT 2421.125 1783.755 2421.415 1783.985 ;
        RECT 2421.275 1783.505 2421.415 1783.755 ;
        RECT 2421.585 1783.745 2421.905 1784.005 ;
        RECT 2422.635 1783.805 2422.775 1784.445 ;
        RECT 2424.485 1784.505 2424.775 1784.545 ;
        RECT 2434.225 1784.505 2434.515 1784.545 ;
        RECT 2424.485 1784.365 2425.055 1784.505 ;
        RECT 2423.115 1784.285 2424.215 1784.365 ;
        RECT 2424.485 1784.315 2424.775 1784.365 ;
        RECT 2422.925 1784.265 2424.215 1784.285 ;
        RECT 2424.915 1784.265 2425.175 1784.365 ;
        RECT 2422.925 1784.225 2424.295 1784.265 ;
        RECT 2424.915 1784.225 2425.255 1784.265 ;
        RECT 2422.925 1784.035 2423.335 1784.225 ;
        RECT 2424.005 1784.035 2424.295 1784.225 ;
        RECT 2424.965 1784.035 2425.255 1784.225 ;
        RECT 2422.925 1784.025 2423.245 1784.035 ;
        RECT 2423.525 1783.805 2423.815 1783.985 ;
        RECT 2422.635 1783.755 2423.815 1783.805 ;
        RECT 2422.635 1783.705 2423.735 1783.755 ;
        RECT 2424.465 1783.745 2424.785 1784.005 ;
        RECT 2426.450 1783.995 2426.790 1784.345 ;
        RECT 2434.225 1784.315 2434.675 1784.505 ;
        RECT 2433.485 1784.025 2433.805 1784.285 ;
        RECT 2422.565 1783.665 2423.735 1783.705 ;
        RECT 2421.275 1783.445 2421.575 1783.505 ;
        RECT 2422.565 1783.455 2422.855 1783.665 ;
        RECT 2426.540 1783.490 2426.710 1783.995 ;
        RECT 2428.055 1783.875 2428.375 1783.980 ;
        RECT 2428.030 1783.860 2428.375 1783.875 ;
        RECT 2428.020 1783.845 2428.375 1783.860 ;
        RECT 2427.855 1783.675 2428.375 1783.845 ;
        RECT 2428.030 1783.660 2428.375 1783.675 ;
        RECT 2428.030 1783.645 2428.320 1783.660 ;
        RECT 2428.830 1783.490 2429.180 1783.610 ;
        RECT 2430.190 1783.540 2430.480 1783.775 ;
        RECT 2431.175 1783.540 2431.465 1783.775 ;
        RECT 2433.965 1783.745 2434.285 1784.005 ;
        RECT 2434.535 1783.985 2434.675 1784.315 ;
        RECT 2435.165 1784.315 2435.715 1784.545 ;
        RECT 2435.855 1784.445 2438.035 1784.585 ;
        RECT 2435.855 1784.365 2437.155 1784.445 ;
        RECT 2435.165 1784.305 2435.485 1784.315 ;
        RECT 2435.855 1784.085 2436.195 1784.365 ;
        RECT 2436.865 1784.315 2437.155 1784.365 ;
        RECT 2435.905 1784.035 2436.195 1784.085 ;
        RECT 2437.325 1784.025 2437.645 1784.285 ;
        RECT 2434.535 1783.845 2434.795 1783.985 ;
        RECT 2430.190 1783.535 2430.420 1783.540 ;
        RECT 2431.175 1783.535 2431.405 1783.540 ;
        RECT 2419.395 1783.385 2419.735 1783.425 ;
        RECT 2420.265 1783.385 2420.585 1783.445 ;
        RECT 2419.395 1783.245 2420.585 1783.385 ;
        RECT 2419.445 1783.195 2419.735 1783.245 ;
        RECT 2420.265 1783.185 2420.585 1783.245 ;
        RECT 2420.735 1783.185 2421.135 1783.445 ;
        RECT 2421.275 1783.385 2421.665 1783.445 ;
        RECT 2422.065 1783.425 2422.385 1783.445 ;
        RECT 2421.845 1783.385 2422.385 1783.425 ;
        RECT 2421.275 1783.365 2422.385 1783.385 ;
        RECT 2421.345 1783.245 2422.385 1783.365 ;
        RECT 2421.345 1783.185 2421.665 1783.245 ;
        RECT 2421.845 1783.195 2422.385 1783.245 ;
        RECT 2422.065 1783.185 2422.385 1783.195 ;
        RECT 2423.295 1783.385 2423.615 1783.445 ;
        RECT 2423.765 1783.385 2424.055 1783.425 ;
        RECT 2423.295 1783.245 2424.055 1783.385 ;
        RECT 2423.295 1783.185 2423.615 1783.245 ;
        RECT 2423.765 1783.195 2424.055 1783.245 ;
        RECT 2424.725 1783.385 2425.015 1783.425 ;
        RECT 2425.155 1783.385 2425.475 1783.445 ;
        RECT 2424.725 1783.245 2425.475 1783.385 ;
        RECT 2426.540 1783.320 2429.180 1783.490 ;
        RECT 2428.660 1783.315 2429.180 1783.320 ;
        RECT 2428.830 1783.260 2429.180 1783.315 ;
        RECT 2424.725 1783.195 2425.015 1783.245 ;
        RECT 2425.155 1783.185 2425.475 1783.245 ;
        RECT 2428.400 1783.120 2428.690 1783.145 ;
        RECT 2429.370 1783.120 2429.720 1783.145 ;
        RECT 2428.400 1782.950 2429.720 1783.120 ;
        RECT 2428.400 1782.915 2428.690 1782.950 ;
        RECT 2413.140 1782.175 2413.430 1782.405 ;
        RECT 2414.930 1782.175 2415.225 1782.435 ;
        RECT 2415.915 1782.175 2416.310 1782.435 ;
        RECT 2428.460 1782.405 2428.630 1782.915 ;
        RECT 2429.370 1782.855 2429.720 1782.950 ;
        RECT 2430.250 1782.435 2430.420 1783.535 ;
        RECT 2431.235 1782.435 2431.405 1783.535 ;
        RECT 2432.795 1783.185 2433.115 1783.445 ;
        RECT 2434.655 1783.425 2434.795 1783.845 ;
        RECT 2434.945 1783.945 2435.235 1783.985 ;
        RECT 2435.405 1783.945 2435.725 1784.005 ;
        RECT 2434.945 1783.805 2435.725 1783.945 ;
        RECT 2434.945 1783.755 2435.235 1783.805 ;
        RECT 2435.405 1783.745 2435.725 1783.805 ;
        RECT 2436.385 1783.755 2436.675 1783.985 ;
        RECT 2436.535 1783.505 2436.675 1783.755 ;
        RECT 2436.845 1783.745 2437.165 1784.005 ;
        RECT 2437.895 1783.805 2438.035 1784.445 ;
        RECT 2439.745 1784.505 2440.035 1784.545 ;
        RECT 2696.970 1784.540 2697.290 1784.600 ;
        RECT 2697.445 1784.555 2697.735 1784.600 ;
        RECT 2698.350 1784.540 2698.670 1784.800 ;
        RECT 2439.745 1784.365 2440.315 1784.505 ;
        RECT 2438.375 1784.285 2439.475 1784.365 ;
        RECT 2439.745 1784.315 2440.035 1784.365 ;
        RECT 2438.185 1784.265 2439.475 1784.285 ;
        RECT 2440.175 1784.265 2440.435 1784.365 ;
        RECT 2438.185 1784.225 2439.555 1784.265 ;
        RECT 2440.175 1784.225 2440.515 1784.265 ;
        RECT 2438.185 1784.035 2438.595 1784.225 ;
        RECT 2439.265 1784.035 2439.555 1784.225 ;
        RECT 2440.225 1784.035 2440.515 1784.225 ;
        RECT 2438.185 1784.025 2438.505 1784.035 ;
        RECT 2438.785 1783.805 2439.075 1783.985 ;
        RECT 2437.895 1783.755 2439.075 1783.805 ;
        RECT 2437.895 1783.705 2438.995 1783.755 ;
        RECT 2439.725 1783.745 2440.045 1784.005 ;
        RECT 2441.710 1783.995 2442.050 1784.345 ;
        RECT 2437.825 1783.665 2438.995 1783.705 ;
        RECT 2436.535 1783.445 2436.835 1783.505 ;
        RECT 2437.825 1783.455 2438.115 1783.665 ;
        RECT 2441.800 1783.490 2441.970 1783.995 ;
        RECT 2443.315 1783.875 2443.635 1783.980 ;
        RECT 2443.290 1783.860 2443.635 1783.875 ;
        RECT 2443.280 1783.845 2443.635 1783.860 ;
        RECT 2443.115 1783.675 2443.635 1783.845 ;
        RECT 2443.290 1783.660 2443.635 1783.675 ;
        RECT 2443.290 1783.645 2443.580 1783.660 ;
        RECT 2444.090 1783.490 2444.440 1783.610 ;
        RECT 2445.450 1783.540 2445.740 1783.775 ;
        RECT 2446.435 1783.540 2446.725 1783.775 ;
        RECT 2445.450 1783.535 2445.680 1783.540 ;
        RECT 2446.435 1783.535 2446.665 1783.540 ;
        RECT 2434.655 1783.385 2434.995 1783.425 ;
        RECT 2435.525 1783.385 2435.845 1783.445 ;
        RECT 2434.655 1783.245 2435.845 1783.385 ;
        RECT 2434.705 1783.195 2434.995 1783.245 ;
        RECT 2435.525 1783.185 2435.845 1783.245 ;
        RECT 2435.995 1783.185 2436.395 1783.445 ;
        RECT 2436.535 1783.385 2436.925 1783.445 ;
        RECT 2437.325 1783.425 2437.645 1783.445 ;
        RECT 2437.105 1783.385 2437.645 1783.425 ;
        RECT 2436.535 1783.365 2437.645 1783.385 ;
        RECT 2436.605 1783.245 2437.645 1783.365 ;
        RECT 2436.605 1783.185 2436.925 1783.245 ;
        RECT 2437.105 1783.195 2437.645 1783.245 ;
        RECT 2437.325 1783.185 2437.645 1783.195 ;
        RECT 2438.555 1783.385 2438.875 1783.445 ;
        RECT 2439.025 1783.385 2439.315 1783.425 ;
        RECT 2438.555 1783.245 2439.315 1783.385 ;
        RECT 2438.555 1783.185 2438.875 1783.245 ;
        RECT 2439.025 1783.195 2439.315 1783.245 ;
        RECT 2439.985 1783.385 2440.275 1783.425 ;
        RECT 2440.415 1783.385 2440.735 1783.445 ;
        RECT 2439.985 1783.245 2440.735 1783.385 ;
        RECT 2441.800 1783.320 2444.440 1783.490 ;
        RECT 2443.920 1783.315 2444.440 1783.320 ;
        RECT 2444.090 1783.260 2444.440 1783.315 ;
        RECT 2439.985 1783.195 2440.275 1783.245 ;
        RECT 2440.415 1783.185 2440.735 1783.245 ;
        RECT 2443.660 1783.120 2443.950 1783.145 ;
        RECT 2444.630 1783.120 2444.980 1783.145 ;
        RECT 2443.660 1782.950 2444.980 1783.120 ;
        RECT 2443.660 1782.915 2443.950 1782.950 ;
        RECT 2428.400 1782.175 2428.690 1782.405 ;
        RECT 2430.190 1782.175 2430.485 1782.435 ;
        RECT 2431.170 1782.175 2431.490 1782.435 ;
        RECT 2443.720 1782.405 2443.890 1782.915 ;
        RECT 2444.630 1782.855 2444.980 1782.950 ;
        RECT 2445.510 1782.435 2445.680 1783.535 ;
        RECT 2446.495 1782.435 2446.665 1783.535 ;
        RECT 2697.890 1782.840 2698.210 1783.100 ;
        RECT 2443.660 1782.175 2443.950 1782.405 ;
        RECT 2445.450 1782.175 2445.745 1782.435 ;
        RECT 2446.435 1782.180 2446.730 1782.435 ;
        RECT 2460.610 1782.180 2460.930 1782.240 ;
        RECT 2446.435 1782.175 2460.930 1782.180 ;
        RECT 2446.440 1782.040 2460.930 1782.175 ;
        RECT 2460.610 1781.980 2460.930 1782.040 ;
        RECT 2694.670 1782.020 2694.990 1782.080 ;
        RECT 2696.985 1782.020 2697.275 1782.065 ;
        RECT 2694.670 1781.880 2697.275 1782.020 ;
        RECT 2694.670 1781.820 2694.990 1781.880 ;
        RECT 2696.985 1781.835 2697.275 1781.880 ;
        RECT 2523.545 1780.680 2523.865 1780.940 ;
        RECT 2697.905 1777.600 2698.195 1777.645 ;
        RECT 2698.810 1777.600 2699.130 1777.660 ;
        RECT 2697.905 1777.460 2699.130 1777.600 ;
        RECT 2697.905 1777.415 2698.195 1777.460 ;
        RECT 2698.810 1777.400 2699.130 1777.460 ;
        RECT 2694.670 1776.580 2694.990 1776.640 ;
        RECT 2696.985 1776.580 2697.275 1776.625 ;
        RECT 2694.670 1776.440 2697.275 1776.580 ;
        RECT 2694.670 1776.380 2694.990 1776.440 ;
        RECT 2696.985 1776.395 2697.275 1776.440 ;
        RECT 2415.990 1773.340 2416.310 1773.400 ;
        RECT 2604.590 1773.340 2604.910 1773.400 ;
        RECT 2415.990 1773.200 2604.910 1773.340 ;
        RECT 2415.990 1773.140 2416.310 1773.200 ;
        RECT 2604.590 1773.140 2604.910 1773.200 ;
        RECT 2400.810 1773.000 2401.130 1773.060 ;
        RECT 2583.890 1773.000 2584.210 1773.060 ;
        RECT 2400.810 1772.860 2584.210 1773.000 ;
        RECT 2400.810 1772.800 2401.130 1772.860 ;
        RECT 2583.890 1772.800 2584.210 1772.860 ;
        RECT 2385.630 1772.660 2385.950 1772.720 ;
        RECT 2480.390 1772.660 2480.710 1772.720 ;
        RECT 2385.630 1772.520 2480.710 1772.660 ;
        RECT 2385.630 1772.460 2385.950 1772.520 ;
        RECT 2480.390 1772.460 2480.710 1772.520 ;
        RECT 2698.350 1772.160 2698.670 1772.220 ;
        RECT 2699.285 1772.160 2699.575 1772.205 ;
        RECT 2698.350 1772.020 2699.575 1772.160 ;
        RECT 2698.350 1771.960 2698.670 1772.020 ;
        RECT 2699.285 1771.975 2699.575 1772.020 ;
        RECT 2702.490 1771.960 2702.810 1772.220 ;
        RECT 2697.905 1771.820 2698.195 1771.865 ;
        RECT 2702.580 1771.820 2702.720 1771.960 ;
        RECT 2697.905 1771.680 2702.720 1771.820 ;
        RECT 2697.905 1771.635 2698.195 1771.680 ;
        RECT 2694.670 1771.140 2694.990 1771.200 ;
        RECT 2696.985 1771.140 2697.275 1771.185 ;
        RECT 2694.670 1771.000 2697.275 1771.140 ;
        RECT 2694.670 1770.940 2694.990 1771.000 ;
        RECT 2696.985 1770.955 2697.275 1771.000 ;
        RECT 2698.350 1770.940 2698.670 1771.200 ;
        RECT 2523.545 1769.210 2523.865 1769.470 ;
        RECT 2431.170 1768.240 2431.490 1768.300 ;
        RECT 2431.170 1768.100 2449.570 1768.240 ;
        RECT 2431.170 1768.040 2431.490 1768.100 ;
        RECT 2449.430 1766.540 2449.570 1768.100 ;
        RECT 2625.290 1766.540 2625.610 1766.600 ;
        RECT 2449.430 1766.400 2625.610 1766.540 ;
        RECT 2625.290 1766.340 2625.610 1766.400 ;
        RECT 2359.910 1710.045 2360.200 1710.275 ;
        RECT 2363.140 1710.045 2363.430 1710.275 ;
        RECT 2374.365 1710.050 2374.655 1710.280 ;
        RECT 2359.970 1709.590 2360.140 1710.045 ;
        RECT 2363.200 1709.675 2363.370 1710.045 ;
        RECT 2359.890 1709.310 2360.230 1709.590 ;
        RECT 2359.910 1709.305 2360.200 1709.310 ;
        RECT 2363.100 1709.305 2363.470 1709.675 ;
        RECT 2374.425 1709.575 2374.595 1710.050 ;
        RECT 2376.155 1710.020 2376.450 1710.280 ;
        RECT 2377.145 1710.020 2377.440 1710.280 ;
        RECT 2379.725 1710.045 2380.015 1710.275 ;
        RECT 2390.950 1710.050 2391.240 1710.280 ;
        RECT 2375.335 1709.575 2375.685 1709.600 ;
        RECT 2374.425 1709.540 2375.685 1709.575 ;
        RECT 2374.365 1709.405 2375.685 1709.540 ;
        RECT 2374.365 1709.310 2374.655 1709.405 ;
        RECT 2375.335 1709.310 2375.685 1709.405 ;
        RECT 2363.600 1709.165 2363.940 1709.195 ;
        RECT 2374.820 1709.170 2375.145 1709.265 ;
        RECT 2363.570 1709.135 2363.940 1709.165 ;
        RECT 2374.795 1709.140 2375.145 1709.170 ;
        RECT 2363.400 1708.965 2363.940 1709.135 ;
        RECT 2374.625 1708.970 2375.145 1709.140 ;
        RECT 2363.570 1708.935 2363.940 1708.965 ;
        RECT 2374.795 1708.940 2375.145 1708.970 ;
        RECT 2363.600 1708.915 2363.940 1708.935 ;
        RECT 2376.215 1708.920 2376.385 1710.020 ;
        RECT 2377.205 1709.270 2377.375 1710.020 ;
        RECT 2379.785 1709.675 2379.955 1710.045 ;
        RECT 2379.685 1709.305 2380.055 1709.675 ;
        RECT 2391.010 1709.575 2391.180 1710.050 ;
        RECT 2392.740 1710.020 2393.035 1710.280 ;
        RECT 2393.730 1710.020 2394.025 1710.280 ;
        RECT 2396.310 1710.050 2396.600 1710.280 ;
        RECT 2407.535 1710.055 2407.825 1710.285 ;
        RECT 2391.920 1709.575 2392.270 1709.600 ;
        RECT 2391.010 1709.540 2392.270 1709.575 ;
        RECT 2390.950 1709.405 2392.270 1709.540 ;
        RECT 2390.950 1709.310 2391.240 1709.405 ;
        RECT 2391.920 1709.310 2392.270 1709.405 ;
        RECT 2377.205 1708.945 2377.535 1709.270 ;
        RECT 2380.185 1709.165 2380.525 1709.195 ;
        RECT 2391.405 1709.170 2391.730 1709.265 ;
        RECT 2380.155 1709.135 2380.525 1709.165 ;
        RECT 2391.380 1709.140 2391.730 1709.170 ;
        RECT 2379.985 1708.965 2380.525 1709.135 ;
        RECT 2391.210 1708.970 2391.730 1709.140 ;
        RECT 2377.205 1708.920 2377.495 1708.945 ;
        RECT 2380.155 1708.935 2380.525 1708.965 ;
        RECT 2391.380 1708.940 2391.730 1708.970 ;
        RECT 2376.155 1708.915 2376.385 1708.920 ;
        RECT 2359.505 1708.775 2359.845 1708.850 ;
        RECT 2374.020 1708.810 2374.340 1708.890 ;
        RECT 2373.995 1708.780 2374.340 1708.810 ;
        RECT 2359.365 1708.605 2359.845 1708.775 ;
        RECT 2373.820 1708.610 2374.340 1708.780 ;
        RECT 2376.155 1708.680 2376.445 1708.915 ;
        RECT 2377.145 1708.805 2377.495 1708.920 ;
        RECT 2380.185 1708.915 2380.525 1708.935 ;
        RECT 2392.800 1708.920 2392.970 1710.020 ;
        RECT 2393.790 1709.270 2393.960 1710.020 ;
        RECT 2396.370 1709.680 2396.540 1710.050 ;
        RECT 2396.270 1709.310 2396.640 1709.680 ;
        RECT 2407.595 1709.580 2407.765 1710.055 ;
        RECT 2409.325 1710.025 2409.620 1710.285 ;
        RECT 2410.315 1710.025 2410.610 1710.285 ;
        RECT 2412.895 1710.055 2413.185 1710.285 ;
        RECT 2424.120 1710.060 2424.410 1710.290 ;
        RECT 2408.505 1709.580 2408.855 1709.605 ;
        RECT 2407.595 1709.545 2408.855 1709.580 ;
        RECT 2407.535 1709.410 2408.855 1709.545 ;
        RECT 2407.535 1709.315 2407.825 1709.410 ;
        RECT 2408.505 1709.315 2408.855 1709.410 ;
        RECT 2393.790 1708.945 2394.120 1709.270 ;
        RECT 2396.800 1709.200 2397.080 1709.230 ;
        RECT 2396.770 1709.170 2397.110 1709.200 ;
        RECT 2407.990 1709.175 2408.315 1709.270 ;
        RECT 2396.740 1709.140 2397.110 1709.170 ;
        RECT 2407.965 1709.145 2408.315 1709.175 ;
        RECT 2396.570 1708.970 2397.110 1709.140 ;
        RECT 2407.795 1708.975 2408.315 1709.145 ;
        RECT 2393.790 1708.920 2394.080 1708.945 ;
        RECT 2392.740 1708.915 2392.970 1708.920 ;
        RECT 2390.605 1708.810 2390.925 1708.890 ;
        RECT 2377.145 1708.680 2377.435 1708.805 ;
        RECT 2390.580 1708.780 2390.925 1708.810 ;
        RECT 2390.405 1708.610 2390.925 1708.780 ;
        RECT 2392.740 1708.680 2393.030 1708.915 ;
        RECT 2393.730 1708.815 2394.080 1708.920 ;
        RECT 2396.740 1708.885 2397.110 1708.970 ;
        RECT 2407.965 1708.945 2408.315 1708.975 ;
        RECT 2409.385 1708.925 2409.555 1710.025 ;
        RECT 2410.375 1709.275 2410.545 1710.025 ;
        RECT 2412.955 1709.685 2413.125 1710.055 ;
        RECT 2412.855 1709.315 2413.225 1709.685 ;
        RECT 2424.180 1709.585 2424.350 1710.060 ;
        RECT 2425.910 1710.030 2426.205 1710.290 ;
        RECT 2426.900 1710.030 2427.195 1710.290 ;
        RECT 2429.475 1710.055 2429.765 1710.285 ;
        RECT 2440.700 1710.060 2440.990 1710.290 ;
        RECT 2425.090 1709.585 2425.440 1709.610 ;
        RECT 2424.180 1709.550 2425.440 1709.585 ;
        RECT 2424.120 1709.415 2425.440 1709.550 ;
        RECT 2424.120 1709.320 2424.410 1709.415 ;
        RECT 2425.090 1709.320 2425.440 1709.415 ;
        RECT 2410.375 1708.950 2410.705 1709.275 ;
        RECT 2413.355 1709.175 2413.695 1709.205 ;
        RECT 2424.575 1709.180 2424.900 1709.275 ;
        RECT 2413.325 1709.145 2413.695 1709.175 ;
        RECT 2424.550 1709.150 2424.900 1709.180 ;
        RECT 2413.155 1708.975 2413.695 1709.145 ;
        RECT 2424.380 1708.980 2424.900 1709.150 ;
        RECT 2410.375 1708.925 2410.665 1708.950 ;
        RECT 2413.325 1708.945 2413.695 1708.975 ;
        RECT 2424.550 1708.950 2424.900 1708.980 ;
        RECT 2413.355 1708.925 2413.695 1708.945 ;
        RECT 2425.970 1708.930 2426.140 1710.030 ;
        RECT 2426.960 1709.280 2427.130 1710.030 ;
        RECT 2429.535 1709.685 2429.705 1710.055 ;
        RECT 2429.435 1709.315 2429.805 1709.685 ;
        RECT 2440.760 1709.585 2440.930 1710.060 ;
        RECT 2442.490 1710.030 2442.785 1710.290 ;
        RECT 2443.480 1710.030 2443.775 1710.290 ;
        RECT 2441.670 1709.585 2442.020 1709.610 ;
        RECT 2440.760 1709.550 2442.020 1709.585 ;
        RECT 2440.700 1709.415 2442.020 1709.550 ;
        RECT 2440.700 1709.320 2440.990 1709.415 ;
        RECT 2441.670 1709.320 2442.020 1709.415 ;
        RECT 2426.960 1708.955 2427.290 1709.280 ;
        RECT 2429.935 1709.175 2430.275 1709.205 ;
        RECT 2441.155 1709.180 2441.480 1709.275 ;
        RECT 2429.905 1709.145 2430.275 1709.175 ;
        RECT 2441.130 1709.150 2441.480 1709.180 ;
        RECT 2429.735 1708.975 2430.275 1709.145 ;
        RECT 2440.960 1708.980 2441.480 1709.150 ;
        RECT 2426.960 1708.930 2427.250 1708.955 ;
        RECT 2429.905 1708.945 2430.275 1708.975 ;
        RECT 2441.130 1708.950 2441.480 1708.980 ;
        RECT 2425.910 1708.925 2426.140 1708.930 ;
        RECT 2409.325 1708.920 2409.555 1708.925 ;
        RECT 2407.190 1708.815 2407.510 1708.895 ;
        RECT 2393.730 1708.680 2394.020 1708.815 ;
        RECT 2407.165 1708.785 2407.510 1708.815 ;
        RECT 2406.990 1708.615 2407.510 1708.785 ;
        RECT 2409.325 1708.685 2409.615 1708.920 ;
        RECT 2410.315 1708.820 2410.665 1708.925 ;
        RECT 2423.775 1708.820 2424.095 1708.900 ;
        RECT 2410.315 1708.685 2410.605 1708.820 ;
        RECT 2423.750 1708.790 2424.095 1708.820 ;
        RECT 2423.575 1708.620 2424.095 1708.790 ;
        RECT 2425.910 1708.690 2426.200 1708.925 ;
        RECT 2426.900 1708.815 2427.250 1708.930 ;
        RECT 2429.935 1708.925 2430.275 1708.945 ;
        RECT 2442.550 1708.930 2442.720 1710.030 ;
        RECT 2443.510 1710.000 2443.775 1710.030 ;
        RECT 2443.510 1709.585 2443.835 1710.000 ;
        RECT 2443.540 1708.930 2443.710 1709.585 ;
        RECT 2442.490 1708.925 2442.720 1708.930 ;
        RECT 2443.480 1708.925 2443.710 1708.930 ;
        RECT 2440.355 1708.820 2440.675 1708.900 ;
        RECT 2426.900 1708.690 2427.190 1708.815 ;
        RECT 2440.330 1708.790 2440.675 1708.820 ;
        RECT 2440.155 1708.620 2440.675 1708.790 ;
        RECT 2442.490 1708.690 2442.780 1708.925 ;
        RECT 2443.480 1708.690 2443.770 1708.925 ;
        RECT 2359.505 1708.570 2359.845 1708.605 ;
        RECT 2373.995 1708.580 2374.340 1708.610 ;
        RECT 2390.580 1708.580 2390.925 1708.610 ;
        RECT 2407.165 1708.585 2407.510 1708.615 ;
        RECT 2423.750 1708.590 2424.095 1708.620 ;
        RECT 2440.330 1708.590 2440.675 1708.620 ;
        RECT 2374.020 1708.565 2374.340 1708.580 ;
        RECT 2390.605 1708.565 2390.925 1708.580 ;
        RECT 2407.190 1708.570 2407.510 1708.585 ;
        RECT 2423.775 1708.575 2424.095 1708.590 ;
        RECT 2440.355 1708.575 2440.675 1708.590 ;
        RECT 2367.280 1707.325 2367.570 1707.365 ;
        RECT 2367.950 1707.325 2368.270 1707.385 ;
        RECT 2367.280 1707.185 2368.270 1707.325 ;
        RECT 2367.280 1707.135 2367.570 1707.185 ;
        RECT 2367.950 1707.125 2368.270 1707.185 ;
        RECT 2368.970 1707.125 2369.290 1707.385 ;
        RECT 2369.660 1707.135 2369.950 1707.365 ;
        RECT 2370.330 1707.325 2370.650 1707.385 ;
        RECT 2383.865 1707.325 2384.155 1707.365 ;
        RECT 2384.535 1707.325 2384.855 1707.385 ;
        RECT 2370.330 1707.185 2370.920 1707.325 ;
        RECT 2383.865 1707.185 2384.855 1707.325 ;
        RECT 2368.040 1706.985 2368.180 1707.125 ;
        RECT 2369.740 1706.985 2369.880 1707.135 ;
        RECT 2370.330 1707.125 2370.650 1707.185 ;
        RECT 2383.865 1707.135 2384.155 1707.185 ;
        RECT 2384.535 1707.125 2384.855 1707.185 ;
        RECT 2385.555 1707.125 2385.875 1707.385 ;
        RECT 2386.245 1707.135 2386.535 1707.365 ;
        RECT 2386.915 1707.325 2387.235 1707.385 ;
        RECT 2400.450 1707.330 2400.740 1707.370 ;
        RECT 2401.120 1707.330 2401.440 1707.390 ;
        RECT 2386.915 1707.185 2387.505 1707.325 ;
        RECT 2400.450 1707.190 2401.440 1707.330 ;
        RECT 2368.040 1706.845 2369.880 1706.985 ;
        RECT 2384.625 1706.985 2384.765 1707.125 ;
        RECT 2386.325 1706.985 2386.465 1707.135 ;
        RECT 2386.915 1707.125 2387.235 1707.185 ;
        RECT 2400.450 1707.140 2400.740 1707.190 ;
        RECT 2401.120 1707.130 2401.440 1707.190 ;
        RECT 2402.140 1707.130 2402.460 1707.390 ;
        RECT 2402.830 1707.140 2403.120 1707.370 ;
        RECT 2403.500 1707.330 2403.820 1707.390 ;
        RECT 2417.035 1707.335 2417.325 1707.375 ;
        RECT 2417.705 1707.335 2418.025 1707.395 ;
        RECT 2403.500 1707.190 2404.090 1707.330 ;
        RECT 2417.035 1707.195 2418.025 1707.335 ;
        RECT 2384.625 1706.845 2386.465 1706.985 ;
        RECT 2401.210 1706.990 2401.350 1707.130 ;
        RECT 2402.910 1706.990 2403.050 1707.140 ;
        RECT 2403.500 1707.130 2403.820 1707.190 ;
        RECT 2417.035 1707.145 2417.325 1707.195 ;
        RECT 2417.705 1707.135 2418.025 1707.195 ;
        RECT 2418.725 1707.135 2419.045 1707.395 ;
        RECT 2419.415 1707.145 2419.705 1707.375 ;
        RECT 2420.085 1707.335 2420.405 1707.395 ;
        RECT 2433.615 1707.335 2433.905 1707.375 ;
        RECT 2434.285 1707.335 2434.605 1707.395 ;
        RECT 2420.085 1707.195 2420.675 1707.335 ;
        RECT 2433.615 1707.195 2434.605 1707.335 ;
        RECT 2401.210 1706.850 2403.050 1706.990 ;
        RECT 2417.795 1706.995 2417.935 1707.135 ;
        RECT 2419.495 1706.995 2419.635 1707.145 ;
        RECT 2420.085 1707.135 2420.405 1707.195 ;
        RECT 2433.615 1707.145 2433.905 1707.195 ;
        RECT 2434.285 1707.135 2434.605 1707.195 ;
        RECT 2435.305 1707.135 2435.625 1707.395 ;
        RECT 2435.995 1707.145 2436.285 1707.375 ;
        RECT 2436.665 1707.335 2436.985 1707.395 ;
        RECT 2436.665 1707.195 2437.255 1707.335 ;
        RECT 2417.795 1706.855 2419.635 1706.995 ;
        RECT 2434.375 1706.995 2434.515 1707.135 ;
        RECT 2436.075 1706.995 2436.215 1707.145 ;
        RECT 2436.665 1707.135 2436.985 1707.195 ;
        RECT 2434.375 1706.855 2436.215 1706.995 ;
        RECT 2365.580 1706.305 2365.870 1706.345 ;
        RECT 2368.290 1706.305 2368.610 1706.365 ;
        RECT 2365.580 1706.165 2368.610 1706.305 ;
        RECT 2365.580 1706.115 2365.870 1706.165 ;
        RECT 2368.290 1706.105 2368.610 1706.165 ;
        RECT 2371.020 1706.105 2371.670 1706.365 ;
        RECT 2382.165 1706.305 2382.455 1706.345 ;
        RECT 2384.875 1706.305 2385.195 1706.365 ;
        RECT 2382.165 1706.165 2385.195 1706.305 ;
        RECT 2382.165 1706.115 2382.455 1706.165 ;
        RECT 2384.875 1706.105 2385.195 1706.165 ;
        RECT 2387.605 1706.105 2388.255 1706.365 ;
        RECT 2398.750 1706.310 2399.040 1706.350 ;
        RECT 2401.460 1706.310 2401.780 1706.370 ;
        RECT 2398.750 1706.170 2401.780 1706.310 ;
        RECT 2398.750 1706.120 2399.040 1706.170 ;
        RECT 2401.460 1706.110 2401.780 1706.170 ;
        RECT 2404.190 1706.110 2404.840 1706.370 ;
        RECT 2415.335 1706.315 2415.625 1706.355 ;
        RECT 2418.045 1706.315 2418.365 1706.375 ;
        RECT 2415.335 1706.175 2418.365 1706.315 ;
        RECT 2415.335 1706.125 2415.625 1706.175 ;
        RECT 2418.045 1706.115 2418.365 1706.175 ;
        RECT 2420.775 1706.115 2421.425 1706.375 ;
        RECT 2431.915 1706.315 2432.205 1706.355 ;
        RECT 2434.625 1706.315 2434.945 1706.375 ;
        RECT 2431.915 1706.175 2434.945 1706.315 ;
        RECT 2431.915 1706.125 2432.205 1706.175 ;
        RECT 2434.625 1706.115 2434.945 1706.175 ;
        RECT 2437.355 1706.115 2438.005 1706.375 ;
        RECT 2366.770 1705.285 2367.060 1705.325 ;
        RECT 2368.980 1705.285 2369.270 1705.325 ;
        RECT 2369.650 1705.285 2369.970 1705.345 ;
        RECT 2366.770 1705.145 2369.970 1705.285 ;
        RECT 2366.770 1705.095 2367.060 1705.145 ;
        RECT 2368.980 1705.095 2369.270 1705.145 ;
        RECT 2369.650 1705.085 2369.970 1705.145 ;
        RECT 2383.355 1705.285 2383.645 1705.325 ;
        RECT 2385.565 1705.285 2385.855 1705.325 ;
        RECT 2386.235 1705.285 2386.555 1705.345 ;
        RECT 2383.355 1705.145 2386.555 1705.285 ;
        RECT 2383.355 1705.095 2383.645 1705.145 ;
        RECT 2385.565 1705.095 2385.855 1705.145 ;
        RECT 2386.235 1705.085 2386.555 1705.145 ;
        RECT 2399.940 1705.290 2400.230 1705.330 ;
        RECT 2402.150 1705.290 2402.440 1705.330 ;
        RECT 2402.820 1705.290 2403.140 1705.350 ;
        RECT 2399.940 1705.150 2403.140 1705.290 ;
        RECT 2399.940 1705.100 2400.230 1705.150 ;
        RECT 2402.150 1705.100 2402.440 1705.150 ;
        RECT 2402.820 1705.090 2403.140 1705.150 ;
        RECT 2416.525 1705.295 2416.815 1705.335 ;
        RECT 2418.735 1705.295 2419.025 1705.335 ;
        RECT 2419.405 1705.295 2419.725 1705.355 ;
        RECT 2416.525 1705.155 2419.725 1705.295 ;
        RECT 2416.525 1705.105 2416.815 1705.155 ;
        RECT 2418.735 1705.105 2419.025 1705.155 ;
        RECT 2419.405 1705.095 2419.725 1705.155 ;
        RECT 2433.105 1705.295 2433.395 1705.335 ;
        RECT 2435.315 1705.295 2435.605 1705.335 ;
        RECT 2435.985 1705.295 2436.305 1705.355 ;
        RECT 2433.105 1705.155 2436.305 1705.295 ;
        RECT 2433.105 1705.105 2433.395 1705.155 ;
        RECT 2435.315 1705.105 2435.605 1705.155 ;
        RECT 2435.985 1705.095 2436.305 1705.155 ;
        RECT 2368.970 1704.605 2369.290 1704.665 ;
        RECT 2370.940 1704.605 2371.230 1704.645 ;
        RECT 2385.555 1704.605 2385.875 1704.665 ;
        RECT 2387.525 1704.605 2387.815 1704.645 ;
        RECT 2402.140 1704.610 2402.460 1704.670 ;
        RECT 2404.110 1704.610 2404.400 1704.650 ;
        RECT 2418.725 1704.615 2419.045 1704.675 ;
        RECT 2420.695 1704.615 2420.985 1704.655 ;
        RECT 2435.305 1704.615 2435.625 1704.675 ;
        RECT 2437.275 1704.615 2437.565 1704.655 ;
        RECT 2368.970 1704.465 2371.235 1704.605 ;
        RECT 2385.555 1704.465 2387.820 1704.605 ;
        RECT 2402.140 1704.470 2404.405 1704.610 ;
        RECT 2418.725 1704.475 2420.990 1704.615 ;
        RECT 2435.305 1704.475 2437.570 1704.615 ;
        RECT 2368.970 1704.405 2369.290 1704.465 ;
        RECT 2370.940 1704.415 2371.230 1704.465 ;
        RECT 2385.555 1704.405 2385.875 1704.465 ;
        RECT 2387.525 1704.415 2387.815 1704.465 ;
        RECT 2402.140 1704.410 2402.460 1704.470 ;
        RECT 2404.110 1704.420 2404.400 1704.470 ;
        RECT 2418.725 1704.415 2419.045 1704.475 ;
        RECT 2420.695 1704.425 2420.985 1704.475 ;
        RECT 2435.305 1704.415 2435.625 1704.475 ;
        RECT 2437.275 1704.425 2437.565 1704.475 ;
        RECT 2410.470 1704.365 2410.790 1704.380 ;
        RECT 2364.610 1704.265 2364.900 1704.305 ;
        RECT 2367.345 1704.265 2368.215 1704.295 ;
        RECT 2369.650 1704.265 2369.970 1704.325 ;
        RECT 2371.350 1704.265 2371.670 1704.325 ;
        RECT 2364.610 1704.155 2369.970 1704.265 ;
        RECT 2364.610 1704.125 2367.485 1704.155 ;
        RECT 2368.075 1704.125 2369.970 1704.155 ;
        RECT 2371.070 1704.125 2371.670 1704.265 ;
        RECT 2364.610 1704.075 2364.900 1704.125 ;
        RECT 2369.650 1704.065 2369.970 1704.125 ;
        RECT 2371.350 1704.065 2371.670 1704.125 ;
        RECT 2381.195 1704.265 2381.485 1704.305 ;
        RECT 2383.930 1704.265 2384.800 1704.295 ;
        RECT 2386.235 1704.265 2386.555 1704.325 ;
        RECT 2387.935 1704.265 2388.255 1704.325 ;
        RECT 2381.195 1704.155 2386.555 1704.265 ;
        RECT 2381.195 1704.125 2384.070 1704.155 ;
        RECT 2384.660 1704.125 2386.555 1704.155 ;
        RECT 2387.655 1704.125 2388.255 1704.265 ;
        RECT 2381.195 1704.075 2381.485 1704.125 ;
        RECT 2386.235 1704.065 2386.555 1704.125 ;
        RECT 2387.935 1704.065 2388.255 1704.125 ;
        RECT 2397.780 1704.270 2398.070 1704.310 ;
        RECT 2400.515 1704.270 2401.385 1704.300 ;
        RECT 2402.820 1704.270 2403.140 1704.330 ;
        RECT 2404.520 1704.270 2404.840 1704.330 ;
        RECT 2397.780 1704.160 2403.140 1704.270 ;
        RECT 2397.780 1704.130 2400.655 1704.160 ;
        RECT 2401.245 1704.130 2403.140 1704.160 ;
        RECT 2404.240 1704.130 2404.840 1704.270 ;
        RECT 2410.315 1704.135 2410.790 1704.365 ;
        RECT 2397.780 1704.080 2398.070 1704.130 ;
        RECT 2402.820 1704.070 2403.140 1704.130 ;
        RECT 2404.520 1704.070 2404.840 1704.130 ;
        RECT 2410.470 1704.120 2410.790 1704.135 ;
        RECT 2414.365 1704.275 2414.655 1704.315 ;
        RECT 2417.100 1704.275 2417.970 1704.305 ;
        RECT 2419.405 1704.275 2419.725 1704.335 ;
        RECT 2421.105 1704.275 2421.425 1704.335 ;
        RECT 2414.365 1704.165 2419.725 1704.275 ;
        RECT 2414.365 1704.135 2417.240 1704.165 ;
        RECT 2417.830 1704.135 2419.725 1704.165 ;
        RECT 2420.825 1704.135 2421.425 1704.275 ;
        RECT 2414.365 1704.085 2414.655 1704.135 ;
        RECT 2419.405 1704.075 2419.725 1704.135 ;
        RECT 2421.105 1704.075 2421.425 1704.135 ;
        RECT 2430.945 1704.275 2431.235 1704.315 ;
        RECT 2433.680 1704.275 2434.550 1704.305 ;
        RECT 2435.985 1704.275 2436.305 1704.335 ;
        RECT 2437.685 1704.275 2438.005 1704.335 ;
        RECT 2430.945 1704.165 2436.305 1704.275 ;
        RECT 2430.945 1704.135 2433.820 1704.165 ;
        RECT 2434.410 1704.135 2436.305 1704.165 ;
        RECT 2437.405 1704.135 2438.005 1704.275 ;
        RECT 2430.945 1704.085 2431.235 1704.135 ;
        RECT 2435.985 1704.075 2436.305 1704.135 ;
        RECT 2437.685 1704.075 2438.005 1704.135 ;
        RECT 2367.610 1703.965 2367.930 1703.975 ;
        RECT 2366.940 1703.735 2367.230 1703.965 ;
        RECT 2367.610 1703.925 2368.070 1703.965 ;
        RECT 2368.290 1703.925 2368.610 1703.985 ;
        RECT 2369.740 1703.925 2369.880 1704.065 ;
        RECT 2367.610 1703.785 2368.090 1703.925 ;
        RECT 2368.290 1703.785 2368.880 1703.925 ;
        RECT 2369.740 1703.785 2370.220 1703.925 ;
        RECT 2374.020 1703.880 2374.340 1703.980 ;
        RECT 2384.195 1703.965 2384.515 1703.975 ;
        RECT 2373.995 1703.860 2374.340 1703.880 ;
        RECT 2367.610 1703.735 2368.070 1703.785 ;
        RECT 2367.020 1703.535 2367.160 1703.735 ;
        RECT 2367.610 1703.715 2367.930 1703.735 ;
        RECT 2368.290 1703.725 2368.610 1703.785 ;
        RECT 2369.340 1703.665 2369.600 1703.695 ;
        RECT 2369.310 1703.645 2369.630 1703.665 ;
        RECT 2370.080 1703.645 2370.220 1703.785 ;
        RECT 2373.705 1703.690 2374.340 1703.860 ;
        RECT 2373.820 1703.680 2374.340 1703.690 ;
        RECT 2373.995 1703.660 2374.340 1703.680 ;
        RECT 2373.995 1703.650 2374.285 1703.660 ;
        RECT 2369.210 1703.535 2369.630 1703.645 ;
        RECT 2367.020 1703.405 2369.630 1703.535 ;
        RECT 2370.000 1703.415 2370.290 1703.645 ;
        RECT 2372.350 1703.490 2372.675 1703.615 ;
        RECT 2374.795 1703.490 2375.145 1703.610 ;
        RECT 2376.155 1703.545 2376.445 1703.780 ;
        RECT 2377.145 1703.545 2377.435 1703.780 ;
        RECT 2383.525 1703.735 2383.815 1703.965 ;
        RECT 2384.195 1703.925 2384.655 1703.965 ;
        RECT 2384.875 1703.925 2385.195 1703.985 ;
        RECT 2386.325 1703.925 2386.465 1704.065 ;
        RECT 2384.195 1703.785 2384.675 1703.925 ;
        RECT 2384.875 1703.785 2385.465 1703.925 ;
        RECT 2386.325 1703.785 2386.805 1703.925 ;
        RECT 2390.605 1703.880 2390.925 1703.980 ;
        RECT 2400.780 1703.970 2401.100 1703.980 ;
        RECT 2390.580 1703.860 2390.925 1703.880 ;
        RECT 2384.195 1703.735 2384.655 1703.785 ;
        RECT 2376.155 1703.540 2376.385 1703.545 ;
        RECT 2377.145 1703.540 2377.375 1703.545 ;
        RECT 2367.020 1703.395 2369.270 1703.405 ;
        RECT 2372.350 1703.320 2375.145 1703.490 ;
        RECT 2372.350 1703.290 2372.675 1703.320 ;
        RECT 2374.795 1703.260 2375.145 1703.320 ;
        RECT 2374.365 1703.120 2374.655 1703.150 ;
        RECT 2375.335 1703.120 2375.685 1703.150 ;
        RECT 2374.365 1702.950 2375.685 1703.120 ;
        RECT 2374.365 1702.920 2374.655 1702.950 ;
        RECT 2374.425 1702.410 2374.595 1702.920 ;
        RECT 2375.335 1702.860 2375.685 1702.950 ;
        RECT 2376.215 1702.440 2376.385 1703.540 ;
        RECT 2377.205 1702.440 2377.375 1703.540 ;
        RECT 2383.605 1703.535 2383.745 1703.735 ;
        RECT 2384.195 1703.715 2384.515 1703.735 ;
        RECT 2384.875 1703.725 2385.195 1703.785 ;
        RECT 2385.925 1703.665 2386.185 1703.695 ;
        RECT 2385.895 1703.645 2386.215 1703.665 ;
        RECT 2386.665 1703.645 2386.805 1703.785 ;
        RECT 2390.290 1703.690 2390.925 1703.860 ;
        RECT 2390.405 1703.680 2390.925 1703.690 ;
        RECT 2390.580 1703.660 2390.925 1703.680 ;
        RECT 2390.580 1703.650 2390.870 1703.660 ;
        RECT 2385.795 1703.535 2386.215 1703.645 ;
        RECT 2383.605 1703.405 2386.215 1703.535 ;
        RECT 2386.585 1703.415 2386.875 1703.645 ;
        RECT 2388.935 1703.490 2389.260 1703.615 ;
        RECT 2391.380 1703.490 2391.730 1703.610 ;
        RECT 2392.740 1703.545 2393.030 1703.780 ;
        RECT 2393.730 1703.545 2394.020 1703.780 ;
        RECT 2400.110 1703.740 2400.400 1703.970 ;
        RECT 2400.780 1703.930 2401.240 1703.970 ;
        RECT 2401.460 1703.930 2401.780 1703.990 ;
        RECT 2402.910 1703.930 2403.050 1704.070 ;
        RECT 2400.780 1703.790 2401.260 1703.930 ;
        RECT 2401.460 1703.790 2402.050 1703.930 ;
        RECT 2402.910 1703.790 2403.390 1703.930 ;
        RECT 2407.190 1703.885 2407.510 1703.985 ;
        RECT 2417.365 1703.975 2417.685 1703.985 ;
        RECT 2407.165 1703.865 2407.510 1703.885 ;
        RECT 2400.780 1703.740 2401.240 1703.790 ;
        RECT 2392.740 1703.540 2392.970 1703.545 ;
        RECT 2393.730 1703.540 2393.960 1703.545 ;
        RECT 2383.605 1703.395 2385.855 1703.405 ;
        RECT 2388.935 1703.320 2391.730 1703.490 ;
        RECT 2388.935 1703.290 2389.260 1703.320 ;
        RECT 2391.380 1703.260 2391.730 1703.320 ;
        RECT 2390.950 1703.120 2391.240 1703.150 ;
        RECT 2391.920 1703.120 2392.270 1703.150 ;
        RECT 2390.950 1702.950 2392.270 1703.120 ;
        RECT 2390.950 1702.920 2391.240 1702.950 ;
        RECT 2374.365 1702.180 2374.655 1702.410 ;
        RECT 2376.155 1702.180 2376.450 1702.440 ;
        RECT 2377.145 1702.180 2377.440 1702.440 ;
        RECT 2391.010 1702.410 2391.180 1702.920 ;
        RECT 2391.920 1702.860 2392.270 1702.950 ;
        RECT 2392.800 1702.440 2392.970 1703.540 ;
        RECT 2393.790 1702.440 2393.960 1703.540 ;
        RECT 2400.190 1703.540 2400.330 1703.740 ;
        RECT 2400.780 1703.720 2401.100 1703.740 ;
        RECT 2401.460 1703.730 2401.780 1703.790 ;
        RECT 2402.510 1703.670 2402.770 1703.700 ;
        RECT 2402.480 1703.650 2402.800 1703.670 ;
        RECT 2403.250 1703.650 2403.390 1703.790 ;
        RECT 2406.875 1703.695 2407.510 1703.865 ;
        RECT 2406.990 1703.685 2407.510 1703.695 ;
        RECT 2407.165 1703.665 2407.510 1703.685 ;
        RECT 2407.165 1703.655 2407.455 1703.665 ;
        RECT 2402.380 1703.540 2402.800 1703.650 ;
        RECT 2400.190 1703.410 2402.800 1703.540 ;
        RECT 2403.170 1703.420 2403.460 1703.650 ;
        RECT 2405.520 1703.495 2405.845 1703.620 ;
        RECT 2407.965 1703.495 2408.315 1703.615 ;
        RECT 2409.325 1703.550 2409.615 1703.785 ;
        RECT 2410.315 1703.550 2410.605 1703.785 ;
        RECT 2416.695 1703.745 2416.985 1703.975 ;
        RECT 2417.365 1703.935 2417.825 1703.975 ;
        RECT 2418.045 1703.935 2418.365 1703.995 ;
        RECT 2419.495 1703.935 2419.635 1704.075 ;
        RECT 2417.365 1703.795 2417.845 1703.935 ;
        RECT 2418.045 1703.795 2418.635 1703.935 ;
        RECT 2419.495 1703.795 2419.975 1703.935 ;
        RECT 2423.775 1703.890 2424.095 1703.990 ;
        RECT 2433.945 1703.975 2434.265 1703.985 ;
        RECT 2423.750 1703.870 2424.095 1703.890 ;
        RECT 2417.365 1703.745 2417.825 1703.795 ;
        RECT 2409.325 1703.545 2409.555 1703.550 ;
        RECT 2410.315 1703.545 2410.545 1703.550 ;
        RECT 2400.190 1703.400 2402.440 1703.410 ;
        RECT 2405.520 1703.325 2408.315 1703.495 ;
        RECT 2405.520 1703.295 2405.845 1703.325 ;
        RECT 2407.965 1703.265 2408.315 1703.325 ;
        RECT 2407.535 1703.125 2407.825 1703.155 ;
        RECT 2408.505 1703.125 2408.855 1703.155 ;
        RECT 2407.535 1702.955 2408.855 1703.125 ;
        RECT 2407.535 1702.925 2407.825 1702.955 ;
        RECT 2390.950 1702.180 2391.240 1702.410 ;
        RECT 2392.740 1702.180 2393.035 1702.440 ;
        RECT 2393.730 1702.180 2394.025 1702.440 ;
        RECT 2407.595 1702.415 2407.765 1702.925 ;
        RECT 2408.505 1702.865 2408.855 1702.955 ;
        RECT 2409.385 1702.445 2409.555 1703.545 ;
        RECT 2410.375 1702.445 2410.545 1703.545 ;
        RECT 2416.775 1703.545 2416.915 1703.745 ;
        RECT 2417.365 1703.725 2417.685 1703.745 ;
        RECT 2418.045 1703.735 2418.365 1703.795 ;
        RECT 2419.095 1703.675 2419.355 1703.705 ;
        RECT 2419.065 1703.655 2419.385 1703.675 ;
        RECT 2419.835 1703.655 2419.975 1703.795 ;
        RECT 2423.460 1703.700 2424.095 1703.870 ;
        RECT 2423.575 1703.690 2424.095 1703.700 ;
        RECT 2423.750 1703.670 2424.095 1703.690 ;
        RECT 2423.750 1703.660 2424.040 1703.670 ;
        RECT 2418.965 1703.545 2419.385 1703.655 ;
        RECT 2416.775 1703.415 2419.385 1703.545 ;
        RECT 2419.755 1703.425 2420.045 1703.655 ;
        RECT 2422.105 1703.500 2422.430 1703.625 ;
        RECT 2424.550 1703.500 2424.900 1703.620 ;
        RECT 2425.910 1703.555 2426.200 1703.790 ;
        RECT 2426.900 1703.555 2427.190 1703.790 ;
        RECT 2433.275 1703.745 2433.565 1703.975 ;
        RECT 2433.945 1703.935 2434.405 1703.975 ;
        RECT 2434.625 1703.935 2434.945 1703.995 ;
        RECT 2436.075 1703.935 2436.215 1704.075 ;
        RECT 2433.945 1703.795 2434.425 1703.935 ;
        RECT 2434.625 1703.795 2435.215 1703.935 ;
        RECT 2436.075 1703.795 2436.555 1703.935 ;
        RECT 2440.355 1703.890 2440.675 1703.990 ;
        RECT 2440.330 1703.870 2440.675 1703.890 ;
        RECT 2433.945 1703.745 2434.405 1703.795 ;
        RECT 2425.910 1703.550 2426.140 1703.555 ;
        RECT 2426.900 1703.550 2427.130 1703.555 ;
        RECT 2416.775 1703.405 2419.025 1703.415 ;
        RECT 2422.105 1703.330 2424.900 1703.500 ;
        RECT 2422.105 1703.300 2422.430 1703.330 ;
        RECT 2424.550 1703.270 2424.900 1703.330 ;
        RECT 2424.120 1703.130 2424.410 1703.160 ;
        RECT 2425.090 1703.130 2425.440 1703.160 ;
        RECT 2424.120 1702.960 2425.440 1703.130 ;
        RECT 2424.120 1702.930 2424.410 1702.960 ;
        RECT 2407.535 1702.185 2407.825 1702.415 ;
        RECT 2409.325 1702.185 2409.620 1702.445 ;
        RECT 2410.315 1702.185 2410.610 1702.445 ;
        RECT 2424.180 1702.420 2424.350 1702.930 ;
        RECT 2425.090 1702.870 2425.440 1702.960 ;
        RECT 2425.970 1702.450 2426.140 1703.550 ;
        RECT 2426.960 1702.450 2427.130 1703.550 ;
        RECT 2433.355 1703.545 2433.495 1703.745 ;
        RECT 2433.945 1703.725 2434.265 1703.745 ;
        RECT 2434.625 1703.735 2434.945 1703.795 ;
        RECT 2435.675 1703.675 2435.935 1703.705 ;
        RECT 2435.645 1703.655 2435.965 1703.675 ;
        RECT 2436.415 1703.655 2436.555 1703.795 ;
        RECT 2440.040 1703.700 2440.675 1703.870 ;
        RECT 2440.155 1703.690 2440.675 1703.700 ;
        RECT 2440.330 1703.670 2440.675 1703.690 ;
        RECT 2440.330 1703.660 2440.620 1703.670 ;
        RECT 2435.545 1703.545 2435.965 1703.655 ;
        RECT 2433.355 1703.415 2435.965 1703.545 ;
        RECT 2436.335 1703.425 2436.625 1703.655 ;
        RECT 2438.685 1703.500 2439.010 1703.625 ;
        RECT 2441.130 1703.500 2441.480 1703.620 ;
        RECT 2442.490 1703.555 2442.780 1703.790 ;
        RECT 2443.480 1703.555 2443.770 1703.790 ;
        RECT 2442.490 1703.550 2442.720 1703.555 ;
        RECT 2443.480 1703.550 2443.710 1703.555 ;
        RECT 2433.355 1703.405 2435.605 1703.415 ;
        RECT 2438.685 1703.330 2441.480 1703.500 ;
        RECT 2438.685 1703.300 2439.010 1703.330 ;
        RECT 2441.130 1703.270 2441.480 1703.330 ;
        RECT 2440.700 1703.130 2440.990 1703.160 ;
        RECT 2441.670 1703.130 2442.020 1703.160 ;
        RECT 2440.700 1702.960 2442.020 1703.130 ;
        RECT 2440.700 1702.930 2440.990 1702.960 ;
        RECT 2424.120 1702.190 2424.410 1702.420 ;
        RECT 2425.910 1702.190 2426.205 1702.450 ;
        RECT 2426.900 1702.390 2427.195 1702.450 ;
        RECT 2427.950 1702.390 2428.270 1702.450 ;
        RECT 2440.760 1702.420 2440.930 1702.930 ;
        RECT 2441.670 1702.870 2442.020 1702.960 ;
        RECT 2442.550 1702.450 2442.720 1703.550 ;
        RECT 2443.540 1702.450 2443.710 1703.550 ;
        RECT 2426.900 1702.250 2428.270 1702.390 ;
        RECT 2426.900 1702.190 2427.195 1702.250 ;
        RECT 2427.950 1702.190 2428.270 1702.250 ;
        RECT 2440.700 1702.190 2440.990 1702.420 ;
        RECT 2442.490 1702.190 2442.785 1702.450 ;
        RECT 2443.480 1702.320 2443.775 1702.450 ;
        RECT 2443.480 1702.190 2443.820 1702.320 ;
        RECT 2377.350 1701.985 2377.670 1702.000 ;
        RECT 2393.910 1701.985 2394.230 1702.000 ;
        RECT 2377.150 1701.755 2377.670 1701.985 ;
        RECT 2393.735 1701.755 2394.230 1701.985 ;
        RECT 2443.680 1701.940 2443.820 1702.190 ;
        RECT 2461.070 1701.940 2461.390 1702.000 ;
        RECT 2443.680 1701.800 2461.390 1701.940 ;
        RECT 2377.350 1701.740 2377.670 1701.755 ;
        RECT 2393.910 1701.740 2394.230 1701.755 ;
        RECT 2461.070 1701.740 2461.390 1701.800 ;
        RECT 2377.350 1696.980 2377.670 1697.240 ;
        RECT 2393.910 1697.180 2394.230 1697.240 ;
        RECT 2681.870 1697.180 2682.190 1697.240 ;
        RECT 2393.910 1697.040 2682.190 1697.180 ;
        RECT 2393.910 1696.980 2394.230 1697.040 ;
        RECT 2681.870 1696.980 2682.190 1697.040 ;
        RECT 2377.440 1696.500 2377.580 1696.980 ;
        RECT 2410.470 1696.840 2410.790 1696.900 ;
        RECT 2576.990 1696.840 2577.310 1696.900 ;
        RECT 2410.470 1696.700 2577.310 1696.840 ;
        RECT 2410.470 1696.640 2410.790 1696.700 ;
        RECT 2576.990 1696.640 2577.310 1696.700 ;
        RECT 2487.290 1696.500 2487.610 1696.560 ;
        RECT 2377.440 1696.360 2487.610 1696.500 ;
        RECT 2487.290 1696.300 2487.610 1696.360 ;
        RECT 2618.390 1690.380 2618.710 1690.440 ;
        RECT 2677.270 1690.380 2677.590 1690.440 ;
        RECT 2618.390 1690.240 2677.590 1690.380 ;
        RECT 2618.390 1690.180 2618.710 1690.240 ;
        RECT 2677.270 1690.180 2677.590 1690.240 ;
        RECT 2695.590 1676.480 2695.910 1676.540 ;
        RECT 2698.810 1676.480 2699.130 1676.540 ;
        RECT 2700.205 1676.480 2700.495 1676.525 ;
        RECT 2695.590 1676.340 2698.120 1676.480 ;
        RECT 2695.590 1676.280 2695.910 1676.340 ;
        RECT 2697.980 1676.140 2698.120 1676.340 ;
        RECT 2698.810 1676.340 2700.495 1676.480 ;
        RECT 2698.810 1676.280 2699.130 1676.340 ;
        RECT 2700.205 1676.295 2700.495 1676.340 ;
        RECT 2702.490 1676.480 2702.810 1676.540 ;
        RECT 2709.865 1676.480 2710.155 1676.525 ;
        RECT 2702.490 1676.340 2710.155 1676.480 ;
        RECT 2702.490 1676.280 2702.810 1676.340 ;
        RECT 2709.865 1676.295 2710.155 1676.340 ;
        RECT 2697.980 1676.000 2701.340 1676.140 ;
        RECT 2695.130 1675.800 2695.450 1675.860 ;
        RECT 2701.200 1675.845 2701.340 1676.000 ;
        RECT 2699.745 1675.800 2700.035 1675.845 ;
        RECT 2695.130 1675.660 2700.035 1675.800 ;
        RECT 2695.130 1675.600 2695.450 1675.660 ;
        RECT 2699.745 1675.615 2700.035 1675.660 ;
        RECT 2701.125 1675.615 2701.415 1675.845 ;
        RECT 2698.365 1675.460 2698.655 1675.505 ;
        RECT 2701.570 1675.460 2701.890 1675.520 ;
        RECT 2698.365 1675.320 2701.890 1675.460 ;
        RECT 2698.365 1675.275 2698.655 1675.320 ;
        RECT 2701.570 1675.260 2701.890 1675.320 ;
        RECT 2721.810 1674.920 2722.130 1675.180 ;
        RECT 2698.350 1674.780 2698.670 1674.840 ;
        RECT 2698.825 1674.780 2699.115 1674.825 ;
        RECT 2698.350 1674.640 2699.115 1674.780 ;
        RECT 2698.350 1674.580 2698.670 1674.640 ;
        RECT 2698.825 1674.595 2699.115 1674.640 ;
        RECT 2731.470 1674.580 2731.790 1674.840 ;
        RECT 2694.670 1672.740 2694.990 1672.800 ;
        RECT 2696.985 1672.740 2697.275 1672.785 ;
        RECT 2694.670 1672.600 2697.275 1672.740 ;
        RECT 2694.670 1672.540 2694.990 1672.600 ;
        RECT 2696.985 1672.555 2697.275 1672.600 ;
        RECT 2697.890 1671.860 2698.210 1672.120 ;
        RECT 2694.670 1664.920 2694.990 1664.980 ;
        RECT 2696.985 1664.920 2697.275 1664.965 ;
        RECT 2694.670 1664.780 2697.275 1664.920 ;
        RECT 2694.670 1664.720 2694.990 1664.780 ;
        RECT 2696.985 1664.735 2697.275 1664.780 ;
        RECT 2696.970 1663.900 2697.290 1663.960 ;
        RECT 2697.905 1663.900 2698.195 1663.945 ;
        RECT 2696.970 1663.760 2698.195 1663.900 ;
        RECT 2696.970 1663.700 2697.290 1663.760 ;
        RECT 2697.905 1663.715 2698.195 1663.760 ;
        RECT 2625.290 1662.840 2625.610 1662.900 ;
        RECT 2677.270 1662.840 2677.590 1662.900 ;
        RECT 2625.290 1662.700 2677.590 1662.840 ;
        RECT 2625.290 1662.640 2625.610 1662.700 ;
        RECT 2677.270 1662.640 2677.590 1662.700 ;
        RECT 2697.430 1662.200 2697.750 1662.260 ;
        RECT 2698.350 1662.200 2698.670 1662.260 ;
        RECT 2697.430 1662.060 2698.670 1662.200 ;
        RECT 2697.430 1662.000 2697.750 1662.060 ;
        RECT 2698.350 1662.000 2698.670 1662.060 ;
        RECT 2698.370 1659.820 2698.660 1659.865 ;
        RECT 2703.890 1659.820 2704.180 1659.865 ;
        RECT 2704.810 1659.820 2705.100 1659.865 ;
        RECT 2698.370 1659.680 2705.100 1659.820 ;
        RECT 2698.370 1659.635 2698.660 1659.680 ;
        RECT 2703.890 1659.635 2704.180 1659.680 ;
        RECT 2704.810 1659.635 2705.100 1659.680 ;
        RECT 2696.985 1659.480 2697.275 1659.525 ;
        RECT 2697.430 1659.480 2697.750 1659.540 ;
        RECT 2696.985 1659.340 2697.750 1659.480 ;
        RECT 2696.985 1659.295 2697.275 1659.340 ;
        RECT 2697.430 1659.280 2697.750 1659.340 ;
        RECT 2697.890 1659.280 2698.210 1659.540 ;
        RECT 2699.290 1659.480 2699.580 1659.525 ;
        RECT 2701.130 1659.480 2701.420 1659.525 ;
        RECT 2699.290 1659.340 2701.420 1659.480 ;
        RECT 2699.290 1659.295 2699.580 1659.340 ;
        RECT 2701.130 1659.295 2701.420 1659.340 ;
        RECT 2703.475 1659.480 2703.765 1659.525 ;
        RECT 2705.315 1659.480 2705.605 1659.525 ;
        RECT 2703.475 1659.340 2705.605 1659.480 ;
        RECT 2703.475 1659.295 2703.765 1659.340 ;
        RECT 2705.315 1659.295 2705.605 1659.340 ;
        RECT 2721.810 1659.280 2722.130 1659.540 ;
        RECT 2702.030 1659.185 2702.350 1659.200 ;
        RECT 2701.585 1659.140 2701.875 1659.185 ;
        RECT 2697.520 1659.000 2701.875 1659.140 ;
        RECT 2697.520 1658.860 2697.660 1659.000 ;
        RECT 2701.585 1658.955 2701.875 1659.000 ;
        RECT 2702.030 1658.955 2702.460 1659.185 ;
        RECT 2702.950 1659.140 2703.270 1659.200 ;
        RECT 2721.900 1659.140 2722.040 1659.280 ;
        RECT 2702.950 1659.000 2722.040 1659.140 ;
        RECT 2702.030 1658.940 2702.350 1658.955 ;
        RECT 2702.950 1658.940 2703.270 1659.000 ;
        RECT 2697.430 1658.600 2697.750 1658.860 ;
        RECT 2700.205 1658.615 2700.495 1658.845 ;
        RECT 2701.165 1658.800 2701.455 1658.845 ;
        RECT 2704.395 1658.800 2704.685 1658.845 ;
        RECT 2701.165 1658.660 2704.685 1658.800 ;
        RECT 2701.165 1658.615 2701.455 1658.660 ;
        RECT 2704.395 1658.615 2704.685 1658.660 ;
        RECT 2700.280 1658.460 2700.420 1658.615 ;
        RECT 2702.490 1658.460 2702.810 1658.520 ;
        RECT 2700.280 1658.320 2702.810 1658.460 ;
        RECT 2702.490 1658.260 2702.810 1658.320 ;
        RECT 2703.870 1658.460 2704.190 1658.520 ;
        RECT 2706.185 1658.460 2706.475 1658.505 ;
        RECT 2703.870 1658.320 2706.475 1658.460 ;
        RECT 2703.870 1658.260 2704.190 1658.320 ;
        RECT 2706.185 1658.275 2706.475 1658.320 ;
        RECT 2697.905 1657.440 2698.195 1657.485 ;
        RECT 2702.030 1657.440 2702.350 1657.500 ;
        RECT 2697.905 1657.300 2702.350 1657.440 ;
        RECT 2697.905 1657.255 2698.195 1657.300 ;
        RECT 2702.030 1657.240 2702.350 1657.300 ;
        RECT 2694.670 1656.420 2694.990 1656.480 ;
        RECT 2696.985 1656.420 2697.275 1656.465 ;
        RECT 2694.670 1656.280 2697.275 1656.420 ;
        RECT 2694.670 1656.220 2694.990 1656.280 ;
        RECT 2696.985 1656.235 2697.275 1656.280 ;
        RECT 2428.410 1656.040 2428.730 1656.100 ;
        RECT 2677.270 1656.040 2677.590 1656.100 ;
        RECT 2428.410 1655.900 2677.590 1656.040 ;
        RECT 2428.410 1655.840 2428.730 1655.900 ;
        RECT 2677.270 1655.840 2677.590 1655.900 ;
        RECT 2698.370 1654.380 2698.660 1654.425 ;
        RECT 2703.890 1654.380 2704.180 1654.425 ;
        RECT 2704.810 1654.380 2705.100 1654.425 ;
        RECT 2698.370 1654.240 2705.100 1654.380 ;
        RECT 2698.370 1654.195 2698.660 1654.240 ;
        RECT 2703.890 1654.195 2704.180 1654.240 ;
        RECT 2704.810 1654.195 2705.100 1654.240 ;
        RECT 2696.970 1653.840 2697.290 1654.100 ;
        RECT 2697.890 1653.840 2698.210 1654.100 ;
        RECT 2699.290 1654.040 2699.580 1654.085 ;
        RECT 2701.130 1654.040 2701.420 1654.085 ;
        RECT 2699.290 1653.900 2701.420 1654.040 ;
        RECT 2699.290 1653.855 2699.580 1653.900 ;
        RECT 2701.130 1653.855 2701.420 1653.900 ;
        RECT 2702.950 1653.840 2703.270 1654.100 ;
        RECT 2703.475 1654.040 2703.765 1654.085 ;
        RECT 2705.315 1654.040 2705.605 1654.085 ;
        RECT 2703.475 1653.900 2705.605 1654.040 ;
        RECT 2703.475 1653.855 2703.765 1653.900 ;
        RECT 2705.315 1653.855 2705.605 1653.900 ;
        RECT 2698.810 1653.700 2699.130 1653.760 ;
        RECT 2702.030 1653.745 2702.350 1653.760 ;
        RECT 2701.585 1653.700 2701.875 1653.745 ;
        RECT 2698.810 1653.560 2701.875 1653.700 ;
        RECT 2698.810 1653.500 2699.130 1653.560 ;
        RECT 2701.585 1653.515 2701.875 1653.560 ;
        RECT 2702.030 1653.515 2702.460 1653.745 ;
        RECT 2702.030 1653.500 2702.350 1653.515 ;
        RECT 2700.205 1653.175 2700.495 1653.405 ;
        RECT 2701.165 1653.360 2701.455 1653.405 ;
        RECT 2704.395 1653.360 2704.685 1653.405 ;
        RECT 2701.165 1653.220 2704.685 1653.360 ;
        RECT 2701.165 1653.175 2701.455 1653.220 ;
        RECT 2704.395 1653.175 2704.685 1653.220 ;
        RECT 2698.350 1653.020 2698.670 1653.080 ;
        RECT 2700.280 1653.020 2700.420 1653.175 ;
        RECT 2702.490 1653.020 2702.810 1653.080 ;
        RECT 2698.350 1652.880 2702.810 1653.020 ;
        RECT 2698.350 1652.820 2698.670 1652.880 ;
        RECT 2702.490 1652.820 2702.810 1652.880 ;
        RECT 2706.170 1652.820 2706.490 1653.080 ;
        RECT 2697.905 1652.000 2698.195 1652.045 ;
        RECT 2702.030 1652.000 2702.350 1652.060 ;
        RECT 2706.170 1652.000 2706.490 1652.060 ;
        RECT 2697.905 1651.860 2702.350 1652.000 ;
        RECT 2697.905 1651.815 2698.195 1651.860 ;
        RECT 2702.030 1651.800 2702.350 1651.860 ;
        RECT 2703.960 1651.860 2706.490 1652.000 ;
        RECT 2697.890 1651.320 2698.210 1651.380 ;
        RECT 2701.570 1651.320 2701.890 1651.380 ;
        RECT 2703.960 1651.365 2704.100 1651.860 ;
        RECT 2706.170 1651.800 2706.490 1651.860 ;
        RECT 2697.890 1651.180 2703.640 1651.320 ;
        RECT 2697.890 1651.120 2698.210 1651.180 ;
        RECT 2701.570 1651.120 2701.890 1651.180 ;
        RECT 2694.670 1650.980 2694.990 1651.040 ;
        RECT 2696.985 1650.980 2697.275 1651.025 ;
        RECT 2694.670 1650.840 2697.275 1650.980 ;
        RECT 2703.500 1650.980 2703.640 1651.180 ;
        RECT 2703.885 1651.135 2704.175 1651.365 ;
        RECT 2704.345 1651.135 2704.635 1651.365 ;
        RECT 2704.420 1650.980 2704.560 1651.135 ;
        RECT 2703.500 1650.840 2704.560 1650.980 ;
        RECT 2694.670 1650.780 2694.990 1650.840 ;
        RECT 2696.985 1650.795 2697.275 1650.840 ;
        RECT 2703.425 1650.640 2703.715 1650.685 ;
        RECT 2703.870 1650.640 2704.190 1650.700 ;
        RECT 2703.425 1650.500 2704.190 1650.640 ;
        RECT 2703.425 1650.455 2703.715 1650.500 ;
        RECT 2703.870 1650.440 2704.190 1650.500 ;
        RECT 2701.570 1650.100 2701.890 1650.360 ;
        RECT 2697.430 1646.560 2697.750 1646.620 ;
        RECT 2697.905 1646.560 2698.195 1646.605 ;
        RECT 2697.430 1646.420 2698.195 1646.560 ;
        RECT 2697.430 1646.360 2697.750 1646.420 ;
        RECT 2697.905 1646.375 2698.195 1646.420 ;
        RECT 2694.670 1645.540 2694.990 1645.600 ;
        RECT 2696.985 1645.540 2697.275 1645.585 ;
        RECT 2694.670 1645.400 2697.275 1645.540 ;
        RECT 2694.670 1645.340 2694.990 1645.400 ;
        RECT 2696.985 1645.355 2697.275 1645.400 ;
        RECT 2701.570 1639.900 2701.890 1640.160 ;
        RECT 2702.505 1640.100 2702.795 1640.145 ;
        RECT 2703.870 1640.100 2704.190 1640.160 ;
        RECT 2731.470 1640.100 2731.790 1640.160 ;
        RECT 2702.505 1639.960 2731.790 1640.100 ;
        RECT 2702.505 1639.915 2702.795 1639.960 ;
        RECT 2703.870 1639.900 2704.190 1639.960 ;
        RECT 2731.470 1639.900 2731.790 1639.960 ;
        RECT 2702.030 1639.220 2702.350 1639.480 ;
        RECT 2697.905 1638.400 2698.195 1638.445 ;
        RECT 2698.810 1638.400 2699.130 1638.460 ;
        RECT 2697.905 1638.260 2699.130 1638.400 ;
        RECT 2697.905 1638.215 2698.195 1638.260 ;
        RECT 2698.810 1638.200 2699.130 1638.260 ;
        RECT 2702.030 1638.200 2702.350 1638.460 ;
        RECT 2703.870 1638.200 2704.190 1638.460 ;
        RECT 2694.670 1637.720 2694.990 1637.780 ;
        RECT 2702.120 1637.765 2702.260 1638.200 ;
        RECT 2703.960 1637.765 2704.100 1638.200 ;
        RECT 2696.985 1637.720 2697.275 1637.765 ;
        RECT 2694.670 1637.580 2697.275 1637.720 ;
        RECT 2694.670 1637.520 2694.990 1637.580 ;
        RECT 2696.985 1637.535 2697.275 1637.580 ;
        RECT 2702.045 1637.535 2702.335 1637.765 ;
        RECT 2703.885 1637.535 2704.175 1637.765 ;
        RECT 2704.790 1637.180 2705.110 1637.440 ;
        RECT 2702.490 1636.840 2702.810 1637.100 ;
        RECT 2702.490 1635.680 2702.810 1635.740 ;
        RECT 2702.490 1635.540 2724.570 1635.680 ;
        RECT 2702.490 1635.480 2702.810 1635.540 ;
        RECT 2724.430 1634.660 2724.570 1635.540 ;
        RECT 2725.505 1634.660 2725.795 1634.705 ;
        RECT 2724.430 1634.520 2725.795 1634.660 ;
        RECT 2725.505 1634.475 2725.795 1634.520 ;
        RECT 2694.670 1632.280 2694.990 1632.340 ;
        RECT 2696.985 1632.280 2697.275 1632.325 ;
        RECT 2694.670 1632.140 2697.275 1632.280 ;
        RECT 2694.670 1632.080 2694.990 1632.140 ;
        RECT 2696.985 1632.095 2697.275 1632.140 ;
        RECT 2697.430 1631.260 2697.750 1631.320 ;
        RECT 2697.905 1631.260 2698.195 1631.305 ;
        RECT 2697.430 1631.120 2698.195 1631.260 ;
        RECT 2697.430 1631.060 2697.750 1631.120 ;
        RECT 2697.905 1631.075 2698.195 1631.120 ;
        RECT 2618.390 1628.500 2618.710 1628.560 ;
        RECT 2677.270 1628.500 2677.590 1628.560 ;
        RECT 2618.390 1628.360 2677.590 1628.500 ;
        RECT 2618.390 1628.300 2618.710 1628.360 ;
        RECT 2677.270 1628.300 2677.590 1628.360 ;
        RECT 2697.890 1626.640 2698.210 1626.900 ;
        RECT 2698.350 1626.640 2698.670 1626.900 ;
        RECT 2697.430 1626.300 2697.750 1626.560 ;
        RECT 2697.980 1626.500 2698.120 1626.640 ;
        RECT 2702.030 1626.500 2702.350 1626.560 ;
        RECT 2697.980 1626.360 2702.350 1626.500 ;
        RECT 2702.030 1626.300 2702.350 1626.360 ;
        RECT 2699.285 1625.820 2699.575 1625.865 ;
        RECT 2702.950 1625.820 2703.270 1625.880 ;
        RECT 2699.285 1625.680 2703.270 1625.820 ;
        RECT 2699.285 1625.635 2699.575 1625.680 ;
        RECT 2702.950 1625.620 2703.270 1625.680 ;
        RECT 2523.545 1624.645 2523.865 1624.905 ;
        RECT 2694.670 1623.780 2694.990 1623.840 ;
        RECT 2696.985 1623.780 2697.275 1623.825 ;
        RECT 2694.670 1623.640 2697.275 1623.780 ;
        RECT 2694.670 1623.580 2694.990 1623.640 ;
        RECT 2696.985 1623.595 2697.275 1623.640 ;
        RECT 2697.890 1622.900 2698.210 1623.160 ;
        RECT 2697.890 1622.080 2698.210 1622.140 ;
        RECT 2698.825 1622.080 2699.115 1622.125 ;
        RECT 2697.890 1621.940 2699.115 1622.080 ;
        RECT 2697.890 1621.880 2698.210 1621.940 ;
        RECT 2698.825 1621.895 2699.115 1621.940 ;
        RECT 2700.665 1622.080 2700.955 1622.125 ;
        RECT 2701.585 1622.080 2701.875 1622.125 ;
        RECT 2700.665 1621.940 2701.875 1622.080 ;
        RECT 2700.665 1621.895 2700.955 1621.940 ;
        RECT 2701.585 1621.895 2701.875 1621.940 ;
        RECT 2702.030 1621.880 2702.350 1622.140 ;
        RECT 2702.950 1621.880 2703.270 1622.140 ;
        RECT 2703.410 1621.880 2703.730 1622.140 ;
        RECT 2698.350 1621.740 2698.670 1621.800 ;
        RECT 2697.980 1621.600 2698.670 1621.740 ;
        RECT 2697.980 1621.105 2698.120 1621.600 ;
        RECT 2698.350 1621.540 2698.670 1621.600 ;
        RECT 2702.120 1621.445 2702.260 1621.880 ;
        RECT 2702.045 1621.215 2702.335 1621.445 ;
        RECT 2702.490 1621.200 2702.810 1621.460 ;
        RECT 2703.040 1621.445 2703.180 1621.880 ;
        RECT 2702.965 1621.215 2703.255 1621.445 ;
        RECT 2697.905 1620.875 2698.195 1621.105 ;
        RECT 2698.350 1620.860 2698.670 1621.120 ;
        RECT 2702.580 1621.060 2702.720 1621.200 ;
        RECT 2703.425 1621.060 2703.715 1621.105 ;
        RECT 2702.580 1620.920 2703.715 1621.060 ;
        RECT 2703.425 1620.875 2703.715 1620.920 ;
        RECT 2702.490 1620.180 2702.810 1620.440 ;
        RECT 2698.810 1619.160 2699.130 1619.420 ;
        RECT 2699.745 1619.360 2700.035 1619.405 ;
        RECT 2702.490 1619.360 2702.810 1619.420 ;
        RECT 2699.745 1619.220 2702.810 1619.360 ;
        RECT 2699.745 1619.175 2700.035 1619.220 ;
        RECT 2702.490 1619.160 2702.810 1619.220 ;
        RECT 2696.985 1619.020 2697.275 1619.065 ;
        RECT 2697.430 1619.020 2697.750 1619.080 ;
        RECT 2696.985 1618.880 2697.750 1619.020 ;
        RECT 2698.900 1619.020 2699.040 1619.160 ;
        RECT 2702.030 1619.020 2702.350 1619.080 ;
        RECT 2698.900 1618.880 2702.350 1619.020 ;
        RECT 2696.985 1618.835 2697.275 1618.880 ;
        RECT 2697.430 1618.820 2697.750 1618.880 ;
        RECT 2702.030 1618.820 2702.350 1618.880 ;
        RECT 2523.545 1618.230 2523.865 1618.490 ;
        RECT 2698.810 1617.460 2699.130 1617.720 ;
        RECT 2697.905 1616.640 2698.195 1616.685 ;
        RECT 2698.810 1616.640 2699.130 1616.700 ;
        RECT 2697.905 1616.500 2699.130 1616.640 ;
        RECT 2697.905 1616.455 2698.195 1616.500 ;
        RECT 2698.810 1616.440 2699.130 1616.500 ;
        RECT 2694.670 1615.960 2694.990 1616.020 ;
        RECT 2696.985 1615.960 2697.275 1616.005 ;
        RECT 2694.670 1615.820 2697.275 1615.960 ;
        RECT 2694.670 1615.760 2694.990 1615.820 ;
        RECT 2696.985 1615.775 2697.275 1615.820 ;
        RECT 2700.205 1613.240 2700.495 1613.285 ;
        RECT 2701.570 1613.240 2701.890 1613.300 ;
        RECT 2700.205 1613.100 2701.890 1613.240 ;
        RECT 2700.205 1613.055 2700.495 1613.100 ;
        RECT 2701.570 1613.040 2701.890 1613.100 ;
        RECT 2698.365 1612.900 2698.655 1612.945 ;
        RECT 2699.730 1612.900 2700.050 1612.960 ;
        RECT 2698.365 1612.760 2700.050 1612.900 ;
        RECT 2698.365 1612.715 2698.655 1612.760 ;
        RECT 2699.730 1612.700 2700.050 1612.760 ;
        RECT 2700.665 1612.900 2700.955 1612.945 ;
        RECT 2703.410 1612.900 2703.730 1612.960 ;
        RECT 2700.665 1612.760 2703.730 1612.900 ;
        RECT 2700.665 1612.715 2700.955 1612.760 ;
        RECT 2703.410 1612.700 2703.730 1612.760 ;
        RECT 2696.970 1612.560 2697.290 1612.620 ;
        RECT 2702.030 1612.560 2702.350 1612.620 ;
        RECT 2696.970 1612.420 2702.350 1612.560 ;
        RECT 2696.970 1612.360 2697.290 1612.420 ;
        RECT 2702.030 1612.360 2702.350 1612.420 ;
        RECT 2698.810 1612.020 2699.130 1612.280 ;
        RECT 2699.270 1612.020 2699.590 1612.280 ;
        RECT 2701.585 1612.220 2701.875 1612.265 ;
        RECT 2703.870 1612.220 2704.190 1612.280 ;
        RECT 2701.585 1612.080 2704.190 1612.220 ;
        RECT 2701.585 1612.035 2701.875 1612.080 ;
        RECT 2703.870 1612.020 2704.190 1612.080 ;
        RECT 2698.810 1611.200 2699.130 1611.260 ;
        RECT 2701.125 1611.200 2701.415 1611.245 ;
        RECT 2698.810 1611.060 2701.415 1611.200 ;
        RECT 2698.810 1611.000 2699.130 1611.060 ;
        RECT 2701.125 1611.015 2701.415 1611.060 ;
        RECT 2699.730 1610.860 2700.050 1610.920 ;
        RECT 2697.520 1610.720 2699.500 1610.860 ;
        RECT 2697.520 1610.580 2697.660 1610.720 ;
        RECT 2697.430 1610.320 2697.750 1610.580 ;
        RECT 2697.890 1610.320 2698.210 1610.580 ;
        RECT 2359.540 1610.055 2359.830 1610.285 ;
        RECT 2362.950 1610.055 2363.240 1610.285 ;
        RECT 2374.635 1610.055 2374.925 1610.285 ;
        RECT 2359.600 1609.590 2359.770 1610.055 ;
        RECT 2363.010 1609.690 2363.180 1610.055 ;
        RECT 2359.510 1609.310 2359.850 1609.590 ;
        RECT 2362.915 1609.320 2363.285 1609.690 ;
        RECT 2374.695 1609.575 2374.865 1610.055 ;
        RECT 2376.425 1610.025 2376.720 1610.285 ;
        RECT 2377.415 1610.025 2377.710 1610.285 ;
        RECT 2380.170 1610.055 2380.460 1610.285 ;
        RECT 2391.855 1610.055 2392.145 1610.285 ;
        RECT 2376.055 1609.650 2376.285 1609.675 ;
        RECT 2376.025 1609.575 2376.315 1609.650 ;
        RECT 2374.695 1609.545 2376.315 1609.575 ;
        RECT 2374.635 1609.405 2376.315 1609.545 ;
        RECT 2362.950 1609.315 2363.240 1609.320 ;
        RECT 2374.635 1609.315 2374.925 1609.405 ;
        RECT 2376.025 1609.355 2376.315 1609.405 ;
        RECT 2376.055 1609.325 2376.285 1609.355 ;
        RECT 2375.090 1609.175 2375.415 1609.265 ;
        RECT 2363.380 1609.145 2363.670 1609.175 ;
        RECT 2375.065 1609.145 2375.415 1609.175 ;
        RECT 2363.210 1609.140 2363.670 1609.145 ;
        RECT 2363.210 1608.975 2363.700 1609.140 ;
        RECT 2374.895 1608.975 2375.415 1609.145 ;
        RECT 2363.360 1608.860 2363.700 1608.975 ;
        RECT 2375.065 1608.945 2375.415 1608.975 ;
        RECT 2375.090 1608.940 2375.415 1608.945 ;
        RECT 2376.485 1608.925 2376.655 1610.025 ;
        RECT 2377.475 1609.270 2377.645 1610.025 ;
        RECT 2380.230 1609.690 2380.400 1610.055 ;
        RECT 2380.135 1609.320 2380.505 1609.690 ;
        RECT 2391.915 1609.575 2392.085 1610.055 ;
        RECT 2393.645 1610.025 2393.940 1610.285 ;
        RECT 2394.635 1610.025 2394.930 1610.285 ;
        RECT 2397.390 1610.060 2397.680 1610.290 ;
        RECT 2409.075 1610.060 2409.365 1610.290 ;
        RECT 2393.275 1609.650 2393.505 1609.675 ;
        RECT 2393.245 1609.575 2393.535 1609.650 ;
        RECT 2391.915 1609.545 2393.535 1609.575 ;
        RECT 2391.855 1609.405 2393.535 1609.545 ;
        RECT 2380.170 1609.315 2380.460 1609.320 ;
        RECT 2391.855 1609.315 2392.145 1609.405 ;
        RECT 2393.245 1609.355 2393.535 1609.405 ;
        RECT 2393.275 1609.325 2393.505 1609.355 ;
        RECT 2377.475 1608.945 2377.805 1609.270 ;
        RECT 2392.310 1609.175 2392.635 1609.265 ;
        RECT 2380.600 1609.145 2380.890 1609.175 ;
        RECT 2392.285 1609.145 2392.635 1609.175 ;
        RECT 2380.430 1609.140 2380.890 1609.145 ;
        RECT 2380.430 1608.975 2380.920 1609.140 ;
        RECT 2392.115 1608.975 2392.635 1609.145 ;
        RECT 2377.475 1608.925 2377.765 1608.945 ;
        RECT 2376.425 1608.920 2376.655 1608.925 ;
        RECT 2359.135 1608.785 2359.475 1608.850 ;
        RECT 2374.290 1608.815 2374.610 1608.890 ;
        RECT 2374.265 1608.785 2374.610 1608.815 ;
        RECT 2358.995 1608.615 2359.475 1608.785 ;
        RECT 2374.090 1608.615 2374.610 1608.785 ;
        RECT 2376.425 1608.685 2376.715 1608.920 ;
        RECT 2377.415 1608.855 2377.765 1608.925 ;
        RECT 2380.580 1608.860 2380.920 1608.975 ;
        RECT 2392.285 1608.945 2392.635 1608.975 ;
        RECT 2392.310 1608.940 2392.635 1608.945 ;
        RECT 2393.705 1608.925 2393.875 1610.025 ;
        RECT 2394.695 1609.270 2394.865 1610.025 ;
        RECT 2397.450 1609.695 2397.620 1610.060 ;
        RECT 2397.355 1609.325 2397.725 1609.695 ;
        RECT 2409.135 1609.580 2409.305 1610.060 ;
        RECT 2410.865 1610.030 2411.160 1610.290 ;
        RECT 2411.855 1610.030 2412.150 1610.290 ;
        RECT 2414.610 1610.055 2414.900 1610.285 ;
        RECT 2426.295 1610.055 2426.585 1610.285 ;
        RECT 2410.495 1609.655 2410.725 1609.680 ;
        RECT 2410.465 1609.580 2410.755 1609.655 ;
        RECT 2409.135 1609.550 2410.755 1609.580 ;
        RECT 2409.075 1609.410 2410.755 1609.550 ;
        RECT 2397.390 1609.320 2397.680 1609.325 ;
        RECT 2409.075 1609.320 2409.365 1609.410 ;
        RECT 2410.465 1609.360 2410.755 1609.410 ;
        RECT 2410.495 1609.330 2410.725 1609.360 ;
        RECT 2394.695 1608.945 2395.025 1609.270 ;
        RECT 2409.530 1609.180 2409.855 1609.270 ;
        RECT 2397.820 1609.150 2398.110 1609.180 ;
        RECT 2409.505 1609.150 2409.855 1609.180 ;
        RECT 2397.650 1609.145 2398.110 1609.150 ;
        RECT 2397.650 1608.980 2398.140 1609.145 ;
        RECT 2409.335 1608.980 2409.855 1609.150 ;
        RECT 2394.695 1608.925 2394.985 1608.945 ;
        RECT 2393.645 1608.920 2393.875 1608.925 ;
        RECT 2377.415 1608.685 2377.705 1608.855 ;
        RECT 2391.510 1608.815 2391.830 1608.890 ;
        RECT 2391.485 1608.785 2391.830 1608.815 ;
        RECT 2391.310 1608.615 2391.830 1608.785 ;
        RECT 2393.645 1608.685 2393.935 1608.920 ;
        RECT 2394.635 1608.855 2394.985 1608.925 ;
        RECT 2397.800 1608.865 2398.140 1608.980 ;
        RECT 2409.505 1608.950 2409.855 1608.980 ;
        RECT 2409.530 1608.945 2409.855 1608.950 ;
        RECT 2410.925 1608.930 2411.095 1610.030 ;
        RECT 2411.915 1609.275 2412.085 1610.030 ;
        RECT 2414.670 1609.690 2414.840 1610.055 ;
        RECT 2414.575 1609.320 2414.945 1609.690 ;
        RECT 2426.355 1609.575 2426.525 1610.055 ;
        RECT 2428.085 1610.025 2428.380 1610.285 ;
        RECT 2429.075 1610.025 2429.370 1610.285 ;
        RECT 2431.830 1610.055 2432.120 1610.285 ;
        RECT 2443.515 1610.055 2443.805 1610.285 ;
        RECT 2427.715 1609.650 2427.945 1609.675 ;
        RECT 2427.685 1609.575 2427.975 1609.650 ;
        RECT 2426.355 1609.545 2427.975 1609.575 ;
        RECT 2426.295 1609.405 2427.975 1609.545 ;
        RECT 2414.610 1609.315 2414.900 1609.320 ;
        RECT 2426.295 1609.315 2426.585 1609.405 ;
        RECT 2427.685 1609.355 2427.975 1609.405 ;
        RECT 2427.715 1609.325 2427.945 1609.355 ;
        RECT 2411.915 1608.950 2412.245 1609.275 ;
        RECT 2426.750 1609.175 2427.075 1609.265 ;
        RECT 2415.040 1609.145 2415.330 1609.175 ;
        RECT 2426.725 1609.145 2427.075 1609.175 ;
        RECT 2414.870 1609.140 2415.330 1609.145 ;
        RECT 2414.870 1608.975 2415.360 1609.140 ;
        RECT 2426.555 1608.975 2427.075 1609.145 ;
        RECT 2411.915 1608.930 2412.205 1608.950 ;
        RECT 2410.865 1608.925 2411.095 1608.930 ;
        RECT 2394.635 1608.685 2394.925 1608.855 ;
        RECT 2408.730 1608.820 2409.050 1608.895 ;
        RECT 2408.705 1608.790 2409.050 1608.820 ;
        RECT 2408.530 1608.620 2409.050 1608.790 ;
        RECT 2410.865 1608.690 2411.155 1608.925 ;
        RECT 2411.855 1608.860 2412.205 1608.930 ;
        RECT 2415.020 1608.860 2415.360 1608.975 ;
        RECT 2426.725 1608.945 2427.075 1608.975 ;
        RECT 2426.750 1608.940 2427.075 1608.945 ;
        RECT 2428.145 1608.925 2428.315 1610.025 ;
        RECT 2429.135 1609.270 2429.305 1610.025 ;
        RECT 2431.890 1609.690 2432.060 1610.055 ;
        RECT 2431.795 1609.320 2432.165 1609.690 ;
        RECT 2443.575 1609.575 2443.745 1610.055 ;
        RECT 2445.305 1610.025 2445.600 1610.285 ;
        RECT 2446.295 1610.025 2446.590 1610.285 ;
        RECT 2699.360 1610.225 2699.500 1610.720 ;
        RECT 2699.730 1610.720 2700.880 1610.860 ;
        RECT 2699.730 1610.660 2700.050 1610.720 ;
        RECT 2444.935 1609.650 2445.165 1609.675 ;
        RECT 2444.905 1609.575 2445.195 1609.650 ;
        RECT 2443.575 1609.545 2445.195 1609.575 ;
        RECT 2443.515 1609.405 2445.195 1609.545 ;
        RECT 2431.830 1609.315 2432.120 1609.320 ;
        RECT 2443.515 1609.315 2443.805 1609.405 ;
        RECT 2444.905 1609.355 2445.195 1609.405 ;
        RECT 2444.935 1609.325 2445.165 1609.355 ;
        RECT 2429.135 1608.945 2429.465 1609.270 ;
        RECT 2443.970 1609.175 2444.295 1609.265 ;
        RECT 2432.260 1609.145 2432.550 1609.175 ;
        RECT 2443.945 1609.145 2444.295 1609.175 ;
        RECT 2432.090 1609.140 2432.550 1609.145 ;
        RECT 2432.090 1608.975 2432.580 1609.140 ;
        RECT 2443.775 1608.975 2444.295 1609.145 ;
        RECT 2429.135 1608.925 2429.425 1608.945 ;
        RECT 2428.085 1608.920 2428.315 1608.925 ;
        RECT 2411.855 1608.690 2412.145 1608.860 ;
        RECT 2425.950 1608.815 2426.270 1608.890 ;
        RECT 2425.925 1608.785 2426.270 1608.815 ;
        RECT 2359.135 1608.570 2359.475 1608.615 ;
        RECT 2374.265 1608.585 2374.610 1608.615 ;
        RECT 2391.485 1608.585 2391.830 1608.615 ;
        RECT 2408.705 1608.590 2409.050 1608.620 ;
        RECT 2425.750 1608.615 2426.270 1608.785 ;
        RECT 2428.085 1608.685 2428.375 1608.920 ;
        RECT 2429.075 1608.850 2429.425 1608.925 ;
        RECT 2432.240 1608.860 2432.580 1608.975 ;
        RECT 2443.945 1608.945 2444.295 1608.975 ;
        RECT 2443.970 1608.940 2444.295 1608.945 ;
        RECT 2445.365 1608.925 2445.535 1610.025 ;
        RECT 2446.325 1610.000 2446.590 1610.025 ;
        RECT 2446.325 1609.585 2446.650 1610.000 ;
        RECT 2699.285 1609.995 2699.575 1610.225 ;
        RECT 2446.355 1608.925 2446.525 1609.585 ;
        RECT 2696.970 1609.500 2697.290 1609.560 ;
        RECT 2698.365 1609.500 2698.655 1609.545 ;
        RECT 2696.970 1609.360 2698.655 1609.500 ;
        RECT 2699.360 1609.500 2699.500 1609.995 ;
        RECT 2700.740 1609.885 2700.880 1610.720 ;
        RECT 2702.030 1610.320 2702.350 1610.580 ;
        RECT 2702.490 1610.320 2702.810 1610.580 ;
        RECT 2702.965 1610.335 2703.255 1610.565 ;
        RECT 2703.040 1610.180 2703.180 1610.335 ;
        RECT 2702.580 1610.040 2703.180 1610.180 ;
        RECT 2700.665 1609.655 2700.955 1609.885 ;
        RECT 2702.580 1609.500 2702.720 1610.040 ;
        RECT 2699.360 1609.360 2702.720 1609.500 ;
        RECT 2696.970 1609.300 2697.290 1609.360 ;
        RECT 2698.365 1609.315 2698.655 1609.360 ;
        RECT 2445.305 1608.920 2445.535 1608.925 ;
        RECT 2446.295 1608.920 2446.525 1608.925 ;
        RECT 2429.075 1608.685 2429.365 1608.850 ;
        RECT 2443.170 1608.815 2443.490 1608.890 ;
        RECT 2443.145 1608.785 2443.490 1608.815 ;
        RECT 2442.970 1608.615 2443.490 1608.785 ;
        RECT 2445.305 1608.685 2445.595 1608.920 ;
        RECT 2446.295 1608.685 2446.585 1608.920 ;
        RECT 2374.290 1608.565 2374.610 1608.585 ;
        RECT 2391.510 1608.565 2391.830 1608.585 ;
        RECT 2408.730 1608.570 2409.050 1608.590 ;
        RECT 2425.925 1608.585 2426.270 1608.615 ;
        RECT 2443.145 1608.585 2443.490 1608.615 ;
        RECT 2425.950 1608.565 2426.270 1608.585 ;
        RECT 2443.170 1608.565 2443.490 1608.585 ;
        RECT 2697.905 1608.480 2698.195 1608.525 ;
        RECT 2698.350 1608.480 2698.670 1608.540 ;
        RECT 2697.905 1608.340 2698.670 1608.480 ;
        RECT 2697.905 1608.295 2698.195 1608.340 ;
        RECT 2698.350 1608.280 2698.670 1608.340 ;
        RECT 2698.810 1608.480 2699.130 1608.540 ;
        RECT 2699.285 1608.480 2699.575 1608.525 ;
        RECT 2698.810 1608.340 2699.575 1608.480 ;
        RECT 2698.810 1608.280 2699.130 1608.340 ;
        RECT 2699.285 1608.295 2699.575 1608.340 ;
        RECT 2366.650 1608.005 2366.940 1608.050 ;
        RECT 2367.655 1608.005 2367.975 1608.035 ;
        RECT 2369.015 1608.005 2369.335 1608.050 ;
        RECT 2366.650 1607.865 2368.565 1608.005 ;
        RECT 2366.650 1607.820 2366.940 1607.865 ;
        RECT 2367.650 1607.835 2367.980 1607.865 ;
        RECT 2367.655 1607.775 2367.975 1607.835 ;
        RECT 2368.425 1607.650 2368.565 1607.865 ;
        RECT 2369.015 1607.865 2369.610 1608.005 ;
        RECT 2369.015 1607.790 2369.335 1607.865 ;
        RECT 2370.390 1607.805 2371.035 1608.050 ;
        RECT 2383.870 1608.005 2384.160 1608.050 ;
        RECT 2384.875 1608.005 2385.195 1608.035 ;
        RECT 2386.235 1608.005 2386.555 1608.050 ;
        RECT 2383.870 1607.865 2385.785 1608.005 ;
        RECT 2383.870 1607.820 2384.160 1607.865 ;
        RECT 2384.870 1607.835 2385.200 1607.865 ;
        RECT 2370.715 1607.775 2371.035 1607.805 ;
        RECT 2384.875 1607.775 2385.195 1607.835 ;
        RECT 2385.645 1607.650 2385.785 1607.865 ;
        RECT 2386.235 1607.865 2386.830 1608.005 ;
        RECT 2386.235 1607.790 2386.555 1607.865 ;
        RECT 2387.610 1607.805 2388.255 1608.050 ;
        RECT 2401.090 1608.010 2401.380 1608.055 ;
        RECT 2402.095 1608.010 2402.415 1608.040 ;
        RECT 2403.455 1608.010 2403.775 1608.055 ;
        RECT 2401.090 1607.870 2403.005 1608.010 ;
        RECT 2401.090 1607.825 2401.380 1607.870 ;
        RECT 2402.090 1607.840 2402.420 1607.870 ;
        RECT 2387.935 1607.775 2388.255 1607.805 ;
        RECT 2402.095 1607.780 2402.415 1607.840 ;
        RECT 2402.865 1607.655 2403.005 1607.870 ;
        RECT 2403.455 1607.870 2404.050 1608.010 ;
        RECT 2403.455 1607.795 2403.775 1607.870 ;
        RECT 2404.830 1607.810 2405.475 1608.055 ;
        RECT 2418.310 1608.005 2418.600 1608.050 ;
        RECT 2419.315 1608.005 2419.635 1608.035 ;
        RECT 2420.675 1608.005 2420.995 1608.050 ;
        RECT 2418.310 1607.865 2420.225 1608.005 ;
        RECT 2418.310 1607.820 2418.600 1607.865 ;
        RECT 2419.310 1607.835 2419.640 1607.865 ;
        RECT 2405.155 1607.780 2405.475 1607.810 ;
        RECT 2419.315 1607.775 2419.635 1607.835 ;
        RECT 2368.425 1607.510 2370.435 1607.650 ;
        RECT 2385.645 1607.510 2387.655 1607.650 ;
        RECT 2402.865 1607.515 2404.875 1607.655 ;
        RECT 2370.295 1607.370 2370.435 1607.510 ;
        RECT 2387.515 1607.370 2387.655 1607.510 ;
        RECT 2404.735 1607.375 2404.875 1607.515 ;
        RECT 2420.085 1607.650 2420.225 1607.865 ;
        RECT 2420.675 1607.865 2421.270 1608.005 ;
        RECT 2420.675 1607.790 2420.995 1607.865 ;
        RECT 2422.050 1607.805 2422.695 1608.050 ;
        RECT 2435.530 1608.005 2435.820 1608.050 ;
        RECT 2436.535 1608.005 2436.855 1608.035 ;
        RECT 2437.895 1608.005 2438.215 1608.050 ;
        RECT 2435.530 1607.865 2437.445 1608.005 ;
        RECT 2435.530 1607.820 2435.820 1607.865 ;
        RECT 2436.530 1607.835 2436.860 1607.865 ;
        RECT 2422.375 1607.775 2422.695 1607.805 ;
        RECT 2436.535 1607.775 2436.855 1607.835 ;
        RECT 2437.305 1607.650 2437.445 1607.865 ;
        RECT 2437.895 1607.865 2438.490 1608.005 ;
        RECT 2437.895 1607.790 2438.215 1607.865 ;
        RECT 2439.270 1607.805 2439.915 1608.050 ;
        RECT 2439.595 1607.775 2439.915 1607.805 ;
        RECT 2420.085 1607.510 2422.095 1607.650 ;
        RECT 2437.305 1607.510 2439.315 1607.650 ;
        RECT 2368.340 1607.125 2368.985 1607.370 ;
        RECT 2368.665 1607.110 2368.985 1607.125 ;
        RECT 2369.695 1607.110 2370.015 1607.370 ;
        RECT 2370.220 1607.140 2370.510 1607.370 ;
        RECT 2371.070 1607.140 2371.360 1607.370 ;
        RECT 2369.785 1606.970 2369.925 1607.110 ;
        RECT 2371.145 1606.970 2371.285 1607.140 ;
        RECT 2385.560 1607.125 2386.205 1607.370 ;
        RECT 2385.885 1607.110 2386.205 1607.125 ;
        RECT 2386.915 1607.110 2387.235 1607.370 ;
        RECT 2387.440 1607.140 2387.730 1607.370 ;
        RECT 2388.290 1607.140 2388.580 1607.370 ;
        RECT 2369.785 1606.830 2371.285 1606.970 ;
        RECT 2387.005 1606.970 2387.145 1607.110 ;
        RECT 2388.365 1606.970 2388.505 1607.140 ;
        RECT 2402.780 1607.130 2403.425 1607.375 ;
        RECT 2403.105 1607.115 2403.425 1607.130 ;
        RECT 2404.135 1607.115 2404.455 1607.375 ;
        RECT 2404.660 1607.145 2404.950 1607.375 ;
        RECT 2405.510 1607.145 2405.800 1607.375 ;
        RECT 2421.955 1607.370 2422.095 1607.510 ;
        RECT 2439.175 1607.370 2439.315 1607.510 ;
        RECT 2694.670 1607.460 2694.990 1607.520 ;
        RECT 2696.985 1607.460 2697.275 1607.505 ;
        RECT 2387.005 1606.830 2388.505 1606.970 ;
        RECT 2404.225 1606.975 2404.365 1607.115 ;
        RECT 2405.585 1606.975 2405.725 1607.145 ;
        RECT 2420.000 1607.125 2420.645 1607.370 ;
        RECT 2420.325 1607.110 2420.645 1607.125 ;
        RECT 2421.355 1607.110 2421.675 1607.370 ;
        RECT 2421.880 1607.140 2422.170 1607.370 ;
        RECT 2422.730 1607.140 2423.020 1607.370 ;
        RECT 2404.225 1606.835 2405.725 1606.975 ;
        RECT 2421.445 1606.970 2421.585 1607.110 ;
        RECT 2422.805 1606.970 2422.945 1607.140 ;
        RECT 2437.220 1607.125 2437.865 1607.370 ;
        RECT 2437.545 1607.110 2437.865 1607.125 ;
        RECT 2438.575 1607.110 2438.895 1607.370 ;
        RECT 2439.100 1607.140 2439.390 1607.370 ;
        RECT 2439.950 1607.140 2440.240 1607.370 ;
        RECT 2694.670 1607.320 2697.275 1607.460 ;
        RECT 2694.670 1607.260 2694.990 1607.320 ;
        RECT 2696.985 1607.275 2697.275 1607.320 ;
        RECT 2697.430 1607.460 2697.750 1607.520 ;
        RECT 2698.825 1607.460 2699.115 1607.505 ;
        RECT 2697.430 1607.320 2699.115 1607.460 ;
        RECT 2697.430 1607.260 2697.750 1607.320 ;
        RECT 2698.825 1607.275 2699.115 1607.320 ;
        RECT 2699.730 1607.260 2700.050 1607.520 ;
        RECT 2421.445 1606.830 2422.945 1606.970 ;
        RECT 2438.665 1606.970 2438.805 1607.110 ;
        RECT 2440.025 1606.970 2440.165 1607.140 ;
        RECT 2438.665 1606.830 2440.165 1606.970 ;
        RECT 2365.615 1606.305 2365.935 1606.365 ;
        RECT 2365.340 1606.165 2365.935 1606.305 ;
        RECT 2365.615 1606.105 2365.935 1606.165 ;
        RECT 2367.890 1606.305 2368.180 1606.350 ;
        RECT 2370.035 1606.305 2370.355 1606.365 ;
        RECT 2382.835 1606.305 2383.155 1606.365 ;
        RECT 2367.890 1606.165 2370.355 1606.305 ;
        RECT 2382.560 1606.165 2383.155 1606.305 ;
        RECT 2367.890 1606.120 2368.180 1606.165 ;
        RECT 2370.035 1606.105 2370.355 1606.165 ;
        RECT 2382.835 1606.105 2383.155 1606.165 ;
        RECT 2385.110 1606.305 2385.400 1606.350 ;
        RECT 2387.255 1606.305 2387.575 1606.365 ;
        RECT 2400.055 1606.310 2400.375 1606.370 ;
        RECT 2385.110 1606.165 2387.575 1606.305 ;
        RECT 2399.780 1606.170 2400.375 1606.310 ;
        RECT 2385.110 1606.120 2385.400 1606.165 ;
        RECT 2387.255 1606.105 2387.575 1606.165 ;
        RECT 2400.055 1606.110 2400.375 1606.170 ;
        RECT 2402.330 1606.310 2402.620 1606.355 ;
        RECT 2404.475 1606.310 2404.795 1606.370 ;
        RECT 2402.330 1606.170 2404.795 1606.310 ;
        RECT 2417.275 1606.305 2417.595 1606.365 ;
        RECT 2402.330 1606.125 2402.620 1606.170 ;
        RECT 2404.475 1606.110 2404.795 1606.170 ;
        RECT 2417.000 1606.165 2417.595 1606.305 ;
        RECT 2417.275 1606.105 2417.595 1606.165 ;
        RECT 2419.550 1606.305 2419.840 1606.350 ;
        RECT 2421.695 1606.305 2422.015 1606.365 ;
        RECT 2434.495 1606.305 2434.815 1606.365 ;
        RECT 2419.550 1606.165 2422.015 1606.305 ;
        RECT 2434.220 1606.165 2434.815 1606.305 ;
        RECT 2419.550 1606.120 2419.840 1606.165 ;
        RECT 2421.695 1606.105 2422.015 1606.165 ;
        RECT 2434.495 1606.105 2434.815 1606.165 ;
        RECT 2436.770 1606.305 2437.060 1606.350 ;
        RECT 2438.915 1606.305 2439.235 1606.365 ;
        RECT 2436.770 1606.165 2439.235 1606.305 ;
        RECT 2436.770 1606.120 2437.060 1606.165 ;
        RECT 2438.915 1606.105 2439.235 1606.165 ;
        RECT 2699.730 1605.760 2700.050 1605.820 ;
        RECT 2700.665 1605.760 2700.955 1605.805 ;
        RECT 2699.730 1605.620 2700.955 1605.760 ;
        RECT 2699.730 1605.560 2700.050 1605.620 ;
        RECT 2700.665 1605.575 2700.955 1605.620 ;
        RECT 2366.990 1605.285 2367.280 1605.330 ;
        RECT 2369.355 1605.285 2369.675 1605.345 ;
        RECT 2366.990 1605.145 2369.675 1605.285 ;
        RECT 2366.990 1605.100 2367.280 1605.145 ;
        RECT 2369.355 1605.085 2369.675 1605.145 ;
        RECT 2370.035 1605.285 2370.355 1605.345 ;
        RECT 2371.070 1605.285 2371.360 1605.330 ;
        RECT 2370.035 1605.145 2371.360 1605.285 ;
        RECT 2370.035 1605.085 2370.355 1605.145 ;
        RECT 2371.070 1605.100 2371.360 1605.145 ;
        RECT 2384.210 1605.285 2384.500 1605.330 ;
        RECT 2386.575 1605.285 2386.895 1605.345 ;
        RECT 2384.210 1605.145 2386.895 1605.285 ;
        RECT 2384.210 1605.100 2384.500 1605.145 ;
        RECT 2386.575 1605.085 2386.895 1605.145 ;
        RECT 2387.255 1605.285 2387.575 1605.345 ;
        RECT 2388.290 1605.285 2388.580 1605.330 ;
        RECT 2387.255 1605.145 2388.580 1605.285 ;
        RECT 2387.255 1605.085 2387.575 1605.145 ;
        RECT 2388.290 1605.100 2388.580 1605.145 ;
        RECT 2401.430 1605.290 2401.720 1605.335 ;
        RECT 2403.795 1605.290 2404.115 1605.350 ;
        RECT 2401.430 1605.150 2404.115 1605.290 ;
        RECT 2401.430 1605.105 2401.720 1605.150 ;
        RECT 2403.795 1605.090 2404.115 1605.150 ;
        RECT 2404.475 1605.290 2404.795 1605.350 ;
        RECT 2405.510 1605.290 2405.800 1605.335 ;
        RECT 2404.475 1605.150 2405.800 1605.290 ;
        RECT 2404.475 1605.090 2404.795 1605.150 ;
        RECT 2405.510 1605.105 2405.800 1605.150 ;
        RECT 2418.650 1605.285 2418.940 1605.330 ;
        RECT 2421.015 1605.285 2421.335 1605.345 ;
        RECT 2418.650 1605.145 2421.335 1605.285 ;
        RECT 2418.650 1605.100 2418.940 1605.145 ;
        RECT 2421.015 1605.085 2421.335 1605.145 ;
        RECT 2421.695 1605.285 2422.015 1605.345 ;
        RECT 2422.730 1605.285 2423.020 1605.330 ;
        RECT 2421.695 1605.145 2423.020 1605.285 ;
        RECT 2421.695 1605.085 2422.015 1605.145 ;
        RECT 2422.730 1605.100 2423.020 1605.145 ;
        RECT 2435.870 1605.285 2436.160 1605.330 ;
        RECT 2438.235 1605.285 2438.555 1605.345 ;
        RECT 2435.870 1605.145 2438.555 1605.285 ;
        RECT 2435.870 1605.100 2436.160 1605.145 ;
        RECT 2438.235 1605.085 2438.555 1605.145 ;
        RECT 2438.915 1605.285 2439.235 1605.345 ;
        RECT 2439.950 1605.285 2440.240 1605.330 ;
        RECT 2438.915 1605.145 2440.240 1605.285 ;
        RECT 2438.915 1605.085 2439.235 1605.145 ;
        RECT 2439.950 1605.100 2440.240 1605.145 ;
        RECT 2365.120 1604.945 2365.410 1604.990 ;
        RECT 2367.995 1604.945 2368.315 1605.005 ;
        RECT 2365.120 1604.805 2368.315 1604.945 ;
        RECT 2365.120 1604.760 2365.410 1604.805 ;
        RECT 2365.615 1604.265 2365.935 1604.325 ;
        RECT 2367.575 1604.315 2367.715 1604.805 ;
        RECT 2367.995 1604.745 2368.315 1604.805 ;
        RECT 2382.340 1604.945 2382.630 1604.990 ;
        RECT 2385.215 1604.945 2385.535 1605.005 ;
        RECT 2382.340 1604.805 2385.535 1604.945 ;
        RECT 2382.340 1604.760 2382.630 1604.805 ;
        RECT 2369.015 1604.605 2369.335 1604.665 ;
        RECT 2368.740 1604.465 2369.335 1604.605 ;
        RECT 2369.015 1604.405 2369.335 1604.465 ;
        RECT 2366.990 1604.270 2367.280 1604.315 ;
        RECT 2365.340 1604.125 2365.935 1604.265 ;
        RECT 2365.615 1604.065 2365.935 1604.125 ;
        RECT 2366.385 1604.130 2367.280 1604.270 ;
        RECT 2366.385 1603.985 2366.525 1604.130 ;
        RECT 2366.990 1604.085 2367.280 1604.130 ;
        RECT 2367.500 1604.085 2367.790 1604.315 ;
        RECT 2368.335 1604.265 2368.655 1604.325 ;
        RECT 2370.715 1604.265 2371.035 1604.325 ;
        RECT 2382.835 1604.265 2383.155 1604.325 ;
        RECT 2384.795 1604.315 2384.935 1604.805 ;
        RECT 2385.215 1604.745 2385.535 1604.805 ;
        RECT 2399.560 1604.950 2399.850 1604.995 ;
        RECT 2402.435 1604.950 2402.755 1605.010 ;
        RECT 2399.560 1604.810 2402.755 1604.950 ;
        RECT 2399.560 1604.765 2399.850 1604.810 ;
        RECT 2386.235 1604.605 2386.555 1604.665 ;
        RECT 2385.960 1604.465 2386.555 1604.605 ;
        RECT 2386.235 1604.405 2386.555 1604.465 ;
        RECT 2384.210 1604.270 2384.500 1604.315 ;
        RECT 2368.060 1604.125 2368.655 1604.265 ;
        RECT 2370.440 1604.125 2371.035 1604.265 ;
        RECT 2382.560 1604.125 2383.155 1604.265 ;
        RECT 2368.335 1604.065 2368.655 1604.125 ;
        RECT 2370.715 1604.065 2371.035 1604.125 ;
        RECT 2382.835 1604.065 2383.155 1604.125 ;
        RECT 2383.605 1604.130 2384.500 1604.270 ;
        RECT 2383.605 1603.985 2383.745 1604.130 ;
        RECT 2384.210 1604.085 2384.500 1604.130 ;
        RECT 2384.720 1604.085 2385.010 1604.315 ;
        RECT 2385.555 1604.265 2385.875 1604.325 ;
        RECT 2387.935 1604.265 2388.255 1604.325 ;
        RECT 2400.055 1604.270 2400.375 1604.330 ;
        RECT 2402.015 1604.320 2402.155 1604.810 ;
        RECT 2402.435 1604.750 2402.755 1604.810 ;
        RECT 2416.780 1604.945 2417.070 1604.990 ;
        RECT 2419.655 1604.945 2419.975 1605.005 ;
        RECT 2416.780 1604.805 2419.975 1604.945 ;
        RECT 2416.780 1604.760 2417.070 1604.805 ;
        RECT 2403.455 1604.610 2403.775 1604.670 ;
        RECT 2403.180 1604.470 2403.775 1604.610 ;
        RECT 2403.455 1604.410 2403.775 1604.470 ;
        RECT 2401.430 1604.275 2401.720 1604.320 ;
        RECT 2385.280 1604.125 2385.875 1604.265 ;
        RECT 2387.660 1604.125 2388.255 1604.265 ;
        RECT 2399.780 1604.130 2400.375 1604.270 ;
        RECT 2385.555 1604.065 2385.875 1604.125 ;
        RECT 2387.935 1604.065 2388.255 1604.125 ;
        RECT 2400.055 1604.070 2400.375 1604.130 ;
        RECT 2400.825 1604.135 2401.720 1604.275 ;
        RECT 2400.825 1603.990 2400.965 1604.135 ;
        RECT 2401.430 1604.090 2401.720 1604.135 ;
        RECT 2401.940 1604.090 2402.230 1604.320 ;
        RECT 2402.775 1604.270 2403.095 1604.330 ;
        RECT 2405.155 1604.270 2405.475 1604.330 ;
        RECT 2402.500 1604.130 2403.095 1604.270 ;
        RECT 2404.880 1604.130 2405.475 1604.270 ;
        RECT 2417.275 1604.265 2417.595 1604.325 ;
        RECT 2419.235 1604.315 2419.375 1604.805 ;
        RECT 2419.655 1604.745 2419.975 1604.805 ;
        RECT 2434.000 1604.945 2434.290 1604.990 ;
        RECT 2436.875 1604.945 2437.195 1605.005 ;
        RECT 2434.000 1604.805 2437.195 1604.945 ;
        RECT 2698.810 1604.880 2699.130 1605.140 ;
        RECT 2434.000 1604.760 2434.290 1604.805 ;
        RECT 2420.675 1604.605 2420.995 1604.665 ;
        RECT 2420.400 1604.465 2420.995 1604.605 ;
        RECT 2420.675 1604.405 2420.995 1604.465 ;
        RECT 2418.650 1604.270 2418.940 1604.315 ;
        RECT 2402.775 1604.070 2403.095 1604.130 ;
        RECT 2405.155 1604.070 2405.475 1604.130 ;
        RECT 2417.000 1604.125 2417.595 1604.265 ;
        RECT 2417.275 1604.065 2417.595 1604.125 ;
        RECT 2418.045 1604.130 2418.940 1604.270 ;
        RECT 2366.295 1603.725 2366.615 1603.985 ;
        RECT 2374.290 1603.875 2374.610 1603.980 ;
        RECT 2374.265 1603.860 2374.610 1603.875 ;
        RECT 2367.655 1603.800 2367.975 1603.815 ;
        RECT 2367.655 1603.755 2368.160 1603.800 ;
        RECT 2367.565 1603.615 2368.160 1603.755 ;
        RECT 2373.975 1603.690 2374.610 1603.860 ;
        RECT 2374.090 1603.675 2374.610 1603.690 ;
        RECT 2374.265 1603.660 2374.610 1603.675 ;
        RECT 2374.265 1603.645 2374.555 1603.660 ;
        RECT 2367.655 1603.570 2368.160 1603.615 ;
        RECT 2367.655 1603.555 2367.975 1603.570 ;
        RECT 2372.620 1603.290 2372.945 1603.615 ;
        RECT 2375.065 1603.485 2375.415 1603.610 ;
        RECT 2376.425 1603.540 2376.715 1603.775 ;
        RECT 2377.410 1603.540 2377.700 1603.775 ;
        RECT 2383.515 1603.725 2383.835 1603.985 ;
        RECT 2391.510 1603.875 2391.830 1603.980 ;
        RECT 2391.485 1603.860 2391.830 1603.875 ;
        RECT 2384.875 1603.800 2385.195 1603.815 ;
        RECT 2384.875 1603.755 2385.380 1603.800 ;
        RECT 2384.785 1603.615 2385.380 1603.755 ;
        RECT 2391.195 1603.690 2391.830 1603.860 ;
        RECT 2391.310 1603.675 2391.830 1603.690 ;
        RECT 2391.485 1603.660 2391.830 1603.675 ;
        RECT 2391.485 1603.645 2391.775 1603.660 ;
        RECT 2384.875 1603.570 2385.380 1603.615 ;
        RECT 2384.875 1603.555 2385.195 1603.570 ;
        RECT 2376.425 1603.535 2376.655 1603.540 ;
        RECT 2377.410 1603.535 2377.640 1603.540 ;
        RECT 2374.895 1603.315 2375.415 1603.485 ;
        RECT 2375.065 1603.260 2375.415 1603.315 ;
        RECT 2376.030 1603.205 2376.260 1603.235 ;
        RECT 2374.635 1603.120 2374.925 1603.145 ;
        RECT 2376.000 1603.120 2376.290 1603.205 ;
        RECT 2374.635 1602.950 2376.290 1603.120 ;
        RECT 2374.635 1602.915 2374.925 1602.950 ;
        RECT 2374.695 1602.405 2374.865 1602.915 ;
        RECT 2376.000 1602.910 2376.290 1602.950 ;
        RECT 2376.030 1602.885 2376.260 1602.910 ;
        RECT 2376.485 1602.435 2376.655 1603.535 ;
        RECT 2377.470 1602.435 2377.640 1603.535 ;
        RECT 2389.840 1603.290 2390.165 1603.615 ;
        RECT 2392.285 1603.485 2392.635 1603.610 ;
        RECT 2393.645 1603.540 2393.935 1603.775 ;
        RECT 2394.630 1603.540 2394.920 1603.775 ;
        RECT 2400.735 1603.730 2401.055 1603.990 ;
        RECT 2418.045 1603.985 2418.185 1604.130 ;
        RECT 2418.650 1604.085 2418.940 1604.130 ;
        RECT 2419.160 1604.085 2419.450 1604.315 ;
        RECT 2419.995 1604.265 2420.315 1604.325 ;
        RECT 2422.375 1604.265 2422.695 1604.325 ;
        RECT 2434.495 1604.265 2434.815 1604.325 ;
        RECT 2436.455 1604.315 2436.595 1604.805 ;
        RECT 2436.875 1604.745 2437.195 1604.805 ;
        RECT 2696.970 1604.740 2697.290 1604.800 ;
        RECT 2697.445 1604.740 2697.735 1604.785 ;
        RECT 2437.895 1604.605 2438.215 1604.665 ;
        RECT 2437.620 1604.465 2438.215 1604.605 ;
        RECT 2696.970 1604.600 2697.735 1604.740 ;
        RECT 2696.970 1604.540 2697.290 1604.600 ;
        RECT 2697.445 1604.555 2697.735 1604.600 ;
        RECT 2698.350 1604.540 2698.670 1604.800 ;
        RECT 2437.895 1604.405 2438.215 1604.465 ;
        RECT 2435.870 1604.270 2436.160 1604.315 ;
        RECT 2419.720 1604.125 2420.315 1604.265 ;
        RECT 2422.100 1604.125 2422.695 1604.265 ;
        RECT 2434.220 1604.125 2434.815 1604.265 ;
        RECT 2419.995 1604.065 2420.315 1604.125 ;
        RECT 2422.375 1604.065 2422.695 1604.125 ;
        RECT 2434.495 1604.065 2434.815 1604.125 ;
        RECT 2435.265 1604.130 2436.160 1604.270 ;
        RECT 2435.265 1603.985 2435.405 1604.130 ;
        RECT 2435.870 1604.085 2436.160 1604.130 ;
        RECT 2436.380 1604.085 2436.670 1604.315 ;
        RECT 2437.215 1604.265 2437.535 1604.325 ;
        RECT 2439.595 1604.265 2439.915 1604.325 ;
        RECT 2436.940 1604.125 2437.535 1604.265 ;
        RECT 2439.320 1604.125 2439.915 1604.265 ;
        RECT 2437.215 1604.065 2437.535 1604.125 ;
        RECT 2439.595 1604.065 2439.915 1604.125 ;
        RECT 2408.730 1603.880 2409.050 1603.985 ;
        RECT 2408.705 1603.865 2409.050 1603.880 ;
        RECT 2402.095 1603.805 2402.415 1603.820 ;
        RECT 2402.095 1603.760 2402.600 1603.805 ;
        RECT 2402.005 1603.620 2402.600 1603.760 ;
        RECT 2408.415 1603.695 2409.050 1603.865 ;
        RECT 2408.530 1603.680 2409.050 1603.695 ;
        RECT 2408.705 1603.665 2409.050 1603.680 ;
        RECT 2408.705 1603.650 2408.995 1603.665 ;
        RECT 2402.095 1603.575 2402.600 1603.620 ;
        RECT 2402.095 1603.560 2402.415 1603.575 ;
        RECT 2393.645 1603.535 2393.875 1603.540 ;
        RECT 2394.630 1603.535 2394.860 1603.540 ;
        RECT 2392.115 1603.315 2392.635 1603.485 ;
        RECT 2392.285 1603.260 2392.635 1603.315 ;
        RECT 2393.250 1603.205 2393.480 1603.235 ;
        RECT 2391.855 1603.120 2392.145 1603.145 ;
        RECT 2393.220 1603.120 2393.510 1603.205 ;
        RECT 2391.855 1602.950 2393.510 1603.120 ;
        RECT 2391.855 1602.915 2392.145 1602.950 ;
        RECT 2374.635 1602.175 2374.925 1602.405 ;
        RECT 2376.425 1602.175 2376.720 1602.435 ;
        RECT 2377.350 1602.175 2377.705 1602.435 ;
        RECT 2391.915 1602.405 2392.085 1602.915 ;
        RECT 2393.220 1602.910 2393.510 1602.950 ;
        RECT 2393.250 1602.885 2393.480 1602.910 ;
        RECT 2393.705 1602.435 2393.875 1603.535 ;
        RECT 2394.690 1602.435 2394.860 1603.535 ;
        RECT 2407.060 1603.295 2407.385 1603.620 ;
        RECT 2409.505 1603.490 2409.855 1603.615 ;
        RECT 2410.865 1603.545 2411.155 1603.780 ;
        RECT 2411.850 1603.545 2412.140 1603.780 ;
        RECT 2417.955 1603.725 2418.275 1603.985 ;
        RECT 2425.950 1603.875 2426.270 1603.980 ;
        RECT 2425.925 1603.860 2426.270 1603.875 ;
        RECT 2419.315 1603.800 2419.635 1603.815 ;
        RECT 2419.315 1603.755 2419.820 1603.800 ;
        RECT 2419.225 1603.615 2419.820 1603.755 ;
        RECT 2425.635 1603.690 2426.270 1603.860 ;
        RECT 2425.750 1603.675 2426.270 1603.690 ;
        RECT 2425.925 1603.660 2426.270 1603.675 ;
        RECT 2425.925 1603.645 2426.215 1603.660 ;
        RECT 2419.315 1603.570 2419.820 1603.615 ;
        RECT 2419.315 1603.555 2419.635 1603.570 ;
        RECT 2410.865 1603.540 2411.095 1603.545 ;
        RECT 2411.850 1603.540 2412.080 1603.545 ;
        RECT 2409.335 1603.320 2409.855 1603.490 ;
        RECT 2409.505 1603.265 2409.855 1603.320 ;
        RECT 2410.470 1603.210 2410.700 1603.240 ;
        RECT 2409.075 1603.125 2409.365 1603.150 ;
        RECT 2410.440 1603.125 2410.730 1603.210 ;
        RECT 2409.075 1602.955 2410.730 1603.125 ;
        RECT 2409.075 1602.920 2409.365 1602.955 ;
        RECT 2391.855 1602.175 2392.145 1602.405 ;
        RECT 2393.645 1602.175 2393.940 1602.435 ;
        RECT 2394.630 1602.175 2394.925 1602.435 ;
        RECT 2409.135 1602.410 2409.305 1602.920 ;
        RECT 2410.440 1602.915 2410.730 1602.955 ;
        RECT 2410.470 1602.890 2410.700 1602.915 ;
        RECT 2410.925 1602.440 2411.095 1603.540 ;
        RECT 2411.910 1602.440 2412.080 1603.540 ;
        RECT 2424.280 1603.290 2424.605 1603.615 ;
        RECT 2426.725 1603.485 2427.075 1603.610 ;
        RECT 2428.085 1603.540 2428.375 1603.775 ;
        RECT 2429.070 1603.540 2429.360 1603.775 ;
        RECT 2435.175 1603.725 2435.495 1603.985 ;
        RECT 2443.170 1603.875 2443.490 1603.980 ;
        RECT 2443.145 1603.860 2443.490 1603.875 ;
        RECT 2436.535 1603.800 2436.855 1603.815 ;
        RECT 2436.535 1603.755 2437.040 1603.800 ;
        RECT 2436.445 1603.615 2437.040 1603.755 ;
        RECT 2442.855 1603.690 2443.490 1603.860 ;
        RECT 2442.970 1603.675 2443.490 1603.690 ;
        RECT 2443.145 1603.660 2443.490 1603.675 ;
        RECT 2443.145 1603.645 2443.435 1603.660 ;
        RECT 2436.535 1603.570 2437.040 1603.615 ;
        RECT 2436.535 1603.555 2436.855 1603.570 ;
        RECT 2428.085 1603.535 2428.315 1603.540 ;
        RECT 2429.070 1603.535 2429.300 1603.540 ;
        RECT 2426.555 1603.315 2427.075 1603.485 ;
        RECT 2426.725 1603.260 2427.075 1603.315 ;
        RECT 2427.690 1603.205 2427.920 1603.235 ;
        RECT 2426.295 1603.120 2426.585 1603.145 ;
        RECT 2427.660 1603.120 2427.950 1603.205 ;
        RECT 2426.295 1602.950 2427.950 1603.120 ;
        RECT 2426.295 1602.915 2426.585 1602.950 ;
        RECT 2409.075 1602.180 2409.365 1602.410 ;
        RECT 2410.865 1602.180 2411.160 1602.440 ;
        RECT 2411.850 1602.380 2412.145 1602.440 ;
        RECT 2426.355 1602.405 2426.525 1602.915 ;
        RECT 2427.660 1602.910 2427.950 1602.950 ;
        RECT 2427.690 1602.885 2427.920 1602.910 ;
        RECT 2428.145 1602.435 2428.315 1603.535 ;
        RECT 2429.130 1603.370 2429.300 1603.535 ;
        RECT 2429.130 1603.200 2429.310 1603.370 ;
        RECT 2441.500 1603.290 2441.825 1603.615 ;
        RECT 2443.945 1603.485 2444.295 1603.610 ;
        RECT 2445.305 1603.540 2445.595 1603.775 ;
        RECT 2446.290 1603.540 2446.580 1603.775 ;
        RECT 2445.305 1603.535 2445.535 1603.540 ;
        RECT 2446.290 1603.535 2446.520 1603.540 ;
        RECT 2443.775 1603.315 2444.295 1603.485 ;
        RECT 2443.945 1603.260 2444.295 1603.315 ;
        RECT 2444.910 1603.205 2445.140 1603.235 ;
        RECT 2429.130 1602.435 2429.300 1603.200 ;
        RECT 2443.515 1603.120 2443.805 1603.145 ;
        RECT 2444.880 1603.120 2445.170 1603.205 ;
        RECT 2443.515 1602.950 2445.170 1603.120 ;
        RECT 2443.515 1602.915 2443.805 1602.950 ;
        RECT 2411.850 1602.120 2412.170 1602.380 ;
        RECT 2426.295 1602.175 2426.585 1602.405 ;
        RECT 2428.085 1602.175 2428.380 1602.435 ;
        RECT 2429.070 1602.175 2429.365 1602.435 ;
        RECT 2443.575 1602.405 2443.745 1602.915 ;
        RECT 2444.880 1602.910 2445.170 1602.950 ;
        RECT 2444.910 1602.885 2445.140 1602.910 ;
        RECT 2445.365 1602.435 2445.535 1603.535 ;
        RECT 2446.350 1602.435 2446.520 1603.535 ;
        RECT 2697.890 1602.840 2698.210 1603.100 ;
        RECT 2443.515 1602.175 2443.805 1602.405 ;
        RECT 2445.305 1602.175 2445.600 1602.435 ;
        RECT 2446.290 1602.175 2446.585 1602.435 ;
        RECT 2394.635 1601.980 2394.925 1602.025 ;
        RECT 2395.290 1601.980 2395.610 1602.040 ;
        RECT 2394.635 1601.840 2395.610 1601.980 ;
        RECT 2394.635 1601.795 2394.925 1601.840 ;
        RECT 2395.290 1601.780 2395.610 1601.840 ;
        RECT 2429.075 1601.980 2429.365 1602.025 ;
        RECT 2429.790 1601.980 2430.110 1602.040 ;
        RECT 2429.075 1601.840 2430.110 1601.980 ;
        RECT 2446.440 1601.980 2446.580 1602.175 ;
        RECT 2461.530 1601.980 2461.850 1602.040 ;
        RECT 2446.440 1601.840 2461.850 1601.980 ;
        RECT 2429.075 1601.795 2429.365 1601.840 ;
        RECT 2429.790 1601.780 2430.110 1601.840 ;
        RECT 2461.530 1601.780 2461.850 1601.840 ;
        RECT 2694.670 1602.020 2694.990 1602.080 ;
        RECT 2696.985 1602.020 2697.275 1602.065 ;
        RECT 2694.670 1601.880 2697.275 1602.020 ;
        RECT 2694.670 1601.820 2694.990 1601.880 ;
        RECT 2696.985 1601.835 2697.275 1601.880 ;
        RECT 2697.905 1597.600 2698.195 1597.645 ;
        RECT 2698.810 1597.600 2699.130 1597.660 ;
        RECT 2697.905 1597.460 2699.130 1597.600 ;
        RECT 2697.905 1597.415 2698.195 1597.460 ;
        RECT 2698.810 1597.400 2699.130 1597.460 ;
        RECT 2694.670 1596.580 2694.990 1596.640 ;
        RECT 2696.985 1596.580 2697.275 1596.625 ;
        RECT 2694.670 1596.440 2697.275 1596.580 ;
        RECT 2694.670 1596.380 2694.990 1596.440 ;
        RECT 2696.985 1596.395 2697.275 1596.440 ;
        RECT 2377.350 1593.620 2377.670 1593.880 ;
        RECT 2395.290 1593.820 2395.610 1593.880 ;
        RECT 2681.410 1593.820 2681.730 1593.880 ;
        RECT 2395.290 1593.680 2681.730 1593.820 ;
        RECT 2395.290 1593.620 2395.610 1593.680 ;
        RECT 2681.410 1593.620 2681.730 1593.680 ;
        RECT 2377.440 1592.800 2377.580 1593.620 ;
        RECT 2411.850 1593.480 2412.170 1593.540 ;
        RECT 2682.790 1593.480 2683.110 1593.540 ;
        RECT 2411.850 1593.340 2683.110 1593.480 ;
        RECT 2411.850 1593.280 2412.170 1593.340 ;
        RECT 2682.790 1593.280 2683.110 1593.340 ;
        RECT 2429.790 1593.140 2430.110 1593.200 ;
        RECT 2680.030 1593.140 2680.350 1593.200 ;
        RECT 2429.790 1593.000 2680.350 1593.140 ;
        RECT 2429.790 1592.940 2430.110 1593.000 ;
        RECT 2680.030 1592.940 2680.350 1593.000 ;
        RECT 2494.190 1592.800 2494.510 1592.860 ;
        RECT 2377.440 1592.660 2494.510 1592.800 ;
        RECT 2494.190 1592.600 2494.510 1592.660 ;
        RECT 2698.350 1592.160 2698.670 1592.220 ;
        RECT 2699.285 1592.160 2699.575 1592.205 ;
        RECT 2698.350 1592.020 2699.575 1592.160 ;
        RECT 2698.350 1591.960 2698.670 1592.020 ;
        RECT 2699.285 1591.975 2699.575 1592.020 ;
        RECT 2702.490 1591.960 2702.810 1592.220 ;
        RECT 2697.905 1591.820 2698.195 1591.865 ;
        RECT 2702.580 1591.820 2702.720 1591.960 ;
        RECT 2697.905 1591.680 2702.720 1591.820 ;
        RECT 2697.905 1591.635 2698.195 1591.680 ;
        RECT 2694.670 1591.140 2694.990 1591.200 ;
        RECT 2696.985 1591.140 2697.275 1591.185 ;
        RECT 2694.670 1591.000 2697.275 1591.140 ;
        RECT 2694.670 1590.940 2694.990 1591.000 ;
        RECT 2696.985 1590.955 2697.275 1591.000 ;
        RECT 2698.350 1590.940 2698.670 1591.200 ;
        RECT 2523.545 1588.985 2523.865 1589.245 ;
        RECT 2523.545 1581.455 2523.865 1581.715 ;
        RECT 2523.545 1575.475 2523.865 1575.735 ;
        RECT 2523.545 1567.060 2523.865 1567.320 ;
        RECT 2359.540 1533.055 2359.830 1533.285 ;
        RECT 2368.120 1533.055 2368.410 1533.285 ;
        RECT 2373.735 1533.055 2374.025 1533.285 ;
        RECT 2359.600 1532.605 2359.770 1533.055 ;
        RECT 2368.180 1532.710 2368.350 1533.055 ;
        RECT 2359.510 1532.315 2359.860 1532.605 ;
        RECT 2368.100 1532.360 2368.470 1532.710 ;
        RECT 2373.795 1532.575 2373.965 1533.055 ;
        RECT 2375.525 1533.025 2375.820 1533.285 ;
        RECT 2374.705 1532.575 2375.055 1532.605 ;
        RECT 2373.795 1532.545 2375.055 1532.575 ;
        RECT 2373.735 1532.405 2375.055 1532.545 ;
        RECT 2368.100 1532.340 2368.410 1532.360 ;
        RECT 2368.120 1532.315 2368.410 1532.340 ;
        RECT 2373.735 1532.315 2374.025 1532.405 ;
        RECT 2374.705 1532.315 2375.055 1532.405 ;
        RECT 2368.550 1532.145 2368.840 1532.175 ;
        RECT 2368.380 1532.140 2368.840 1532.145 ;
        RECT 2369.585 1532.140 2369.935 1532.240 ;
        RECT 2374.190 1532.175 2374.515 1532.265 ;
        RECT 2374.165 1532.145 2374.515 1532.175 ;
        RECT 2373.995 1532.140 2374.515 1532.145 ;
        RECT 2368.380 1531.975 2374.515 1532.140 ;
        RECT 2368.550 1531.970 2374.515 1531.975 ;
        RECT 2368.550 1531.945 2368.840 1531.970 ;
        RECT 2369.585 1531.890 2369.935 1531.970 ;
        RECT 2374.165 1531.945 2374.515 1531.970 ;
        RECT 2374.190 1531.940 2374.515 1531.945 ;
        RECT 2375.585 1531.925 2375.755 1533.025 ;
        RECT 2376.520 1533.020 2376.815 1533.280 ;
        RECT 2384.445 1533.055 2384.735 1533.285 ;
        RECT 2390.060 1533.055 2390.350 1533.285 ;
        RECT 2376.580 1532.290 2376.750 1533.020 ;
        RECT 2384.505 1532.710 2384.675 1533.055 ;
        RECT 2384.425 1532.360 2384.795 1532.710 ;
        RECT 2390.120 1532.575 2390.290 1533.055 ;
        RECT 2391.850 1533.025 2392.145 1533.285 ;
        RECT 2391.030 1532.575 2391.380 1532.605 ;
        RECT 2390.120 1532.545 2391.380 1532.575 ;
        RECT 2390.060 1532.405 2391.380 1532.545 ;
        RECT 2384.425 1532.340 2384.735 1532.360 ;
        RECT 2384.445 1532.315 2384.735 1532.340 ;
        RECT 2390.060 1532.315 2390.350 1532.405 ;
        RECT 2391.030 1532.315 2391.380 1532.405 ;
        RECT 2375.525 1531.920 2375.755 1531.925 ;
        RECT 2376.570 1531.940 2376.920 1532.290 ;
        RECT 2385.075 1532.175 2385.425 1532.245 ;
        RECT 2390.515 1532.175 2390.840 1532.265 ;
        RECT 2384.875 1532.145 2385.425 1532.175 ;
        RECT 2390.490 1532.145 2390.840 1532.175 ;
        RECT 2384.705 1532.140 2385.425 1532.145 ;
        RECT 2390.320 1532.140 2390.840 1532.145 ;
        RECT 2384.705 1531.975 2390.840 1532.140 ;
        RECT 2384.875 1531.970 2390.840 1531.975 ;
        RECT 2384.875 1531.945 2385.425 1531.970 ;
        RECT 2390.490 1531.945 2390.840 1531.970 ;
        RECT 2376.570 1531.920 2376.870 1531.940 ;
        RECT 2359.135 1531.785 2359.485 1531.860 ;
        RECT 2373.390 1531.815 2373.710 1531.830 ;
        RECT 2373.365 1531.785 2373.710 1531.815 ;
        RECT 2358.995 1531.615 2359.485 1531.785 ;
        RECT 2373.190 1531.615 2373.710 1531.785 ;
        RECT 2375.525 1531.685 2375.815 1531.920 ;
        RECT 2376.520 1531.850 2376.870 1531.920 ;
        RECT 2385.075 1531.895 2385.425 1531.945 ;
        RECT 2390.515 1531.940 2390.840 1531.945 ;
        RECT 2391.910 1531.925 2392.080 1533.025 ;
        RECT 2392.845 1533.020 2393.140 1533.280 ;
        RECT 2400.770 1533.055 2401.060 1533.285 ;
        RECT 2406.385 1533.055 2406.675 1533.285 ;
        RECT 2392.905 1532.300 2393.075 1533.020 ;
        RECT 2400.830 1532.710 2401.000 1533.055 ;
        RECT 2400.750 1532.360 2401.120 1532.710 ;
        RECT 2406.445 1532.575 2406.615 1533.055 ;
        RECT 2408.175 1533.025 2408.470 1533.285 ;
        RECT 2407.355 1532.575 2407.705 1532.605 ;
        RECT 2406.445 1532.545 2407.705 1532.575 ;
        RECT 2406.385 1532.405 2407.705 1532.545 ;
        RECT 2400.750 1532.340 2401.060 1532.360 ;
        RECT 2400.770 1532.315 2401.060 1532.340 ;
        RECT 2406.385 1532.315 2406.675 1532.405 ;
        RECT 2407.355 1532.315 2407.705 1532.405 ;
        RECT 2391.850 1531.920 2392.080 1531.925 ;
        RECT 2392.890 1531.945 2393.245 1532.300 ;
        RECT 2401.400 1532.175 2401.750 1532.250 ;
        RECT 2406.840 1532.175 2407.165 1532.265 ;
        RECT 2401.200 1532.145 2401.750 1532.175 ;
        RECT 2406.815 1532.145 2407.165 1532.175 ;
        RECT 2401.030 1532.140 2401.750 1532.145 ;
        RECT 2406.645 1532.140 2407.165 1532.145 ;
        RECT 2401.030 1531.975 2407.165 1532.140 ;
        RECT 2401.200 1531.970 2407.165 1531.975 ;
        RECT 2401.200 1531.945 2401.750 1531.970 ;
        RECT 2406.815 1531.945 2407.165 1531.970 ;
        RECT 2392.890 1531.920 2393.195 1531.945 ;
        RECT 2376.520 1531.680 2376.810 1531.850 ;
        RECT 2389.715 1531.815 2390.035 1531.830 ;
        RECT 2389.690 1531.785 2390.035 1531.815 ;
        RECT 2389.515 1531.615 2390.035 1531.785 ;
        RECT 2391.850 1531.685 2392.140 1531.920 ;
        RECT 2392.845 1531.850 2393.195 1531.920 ;
        RECT 2401.400 1531.900 2401.750 1531.945 ;
        RECT 2406.840 1531.940 2407.165 1531.945 ;
        RECT 2408.235 1531.925 2408.405 1533.025 ;
        RECT 2409.170 1533.020 2409.465 1533.280 ;
        RECT 2417.095 1533.055 2417.385 1533.285 ;
        RECT 2422.710 1533.055 2423.000 1533.285 ;
        RECT 2409.230 1532.290 2409.400 1533.020 ;
        RECT 2417.155 1532.710 2417.325 1533.055 ;
        RECT 2417.075 1532.360 2417.445 1532.710 ;
        RECT 2422.770 1532.575 2422.940 1533.055 ;
        RECT 2424.500 1533.025 2424.795 1533.285 ;
        RECT 2423.680 1532.575 2424.030 1532.605 ;
        RECT 2422.770 1532.545 2424.030 1532.575 ;
        RECT 2422.710 1532.405 2424.030 1532.545 ;
        RECT 2417.075 1532.340 2417.385 1532.360 ;
        RECT 2417.095 1532.315 2417.385 1532.340 ;
        RECT 2422.710 1532.315 2423.000 1532.405 ;
        RECT 2423.680 1532.315 2424.030 1532.405 ;
        RECT 2408.175 1531.920 2408.405 1531.925 ;
        RECT 2409.175 1531.940 2409.525 1532.290 ;
        RECT 2417.725 1532.175 2418.075 1532.245 ;
        RECT 2423.165 1532.175 2423.490 1532.265 ;
        RECT 2417.525 1532.145 2418.075 1532.175 ;
        RECT 2423.140 1532.145 2423.490 1532.175 ;
        RECT 2417.355 1532.140 2418.075 1532.145 ;
        RECT 2422.970 1532.140 2423.490 1532.145 ;
        RECT 2417.355 1531.975 2423.490 1532.140 ;
        RECT 2417.525 1531.970 2423.490 1531.975 ;
        RECT 2417.525 1531.945 2418.075 1531.970 ;
        RECT 2423.140 1531.945 2423.490 1531.970 ;
        RECT 2409.175 1531.920 2409.520 1531.940 ;
        RECT 2392.845 1531.680 2393.135 1531.850 ;
        RECT 2406.040 1531.815 2406.360 1531.830 ;
        RECT 2406.015 1531.785 2406.360 1531.815 ;
        RECT 2405.840 1531.615 2406.360 1531.785 ;
        RECT 2408.175 1531.685 2408.465 1531.920 ;
        RECT 2409.170 1531.845 2409.520 1531.920 ;
        RECT 2417.725 1531.895 2418.075 1531.945 ;
        RECT 2423.165 1531.940 2423.490 1531.945 ;
        RECT 2424.560 1531.925 2424.730 1533.025 ;
        RECT 2425.495 1533.020 2425.790 1533.280 ;
        RECT 2433.420 1533.055 2433.710 1533.285 ;
        RECT 2439.035 1533.055 2439.325 1533.285 ;
        RECT 2425.555 1532.290 2425.725 1533.020 ;
        RECT 2433.480 1532.710 2433.650 1533.055 ;
        RECT 2433.400 1532.360 2433.770 1532.710 ;
        RECT 2439.095 1532.575 2439.265 1533.055 ;
        RECT 2440.825 1533.025 2441.120 1533.285 ;
        RECT 2440.005 1532.575 2440.355 1532.605 ;
        RECT 2439.095 1532.545 2440.355 1532.575 ;
        RECT 2439.035 1532.405 2440.355 1532.545 ;
        RECT 2433.400 1532.340 2433.710 1532.360 ;
        RECT 2433.420 1532.315 2433.710 1532.340 ;
        RECT 2439.035 1532.315 2439.325 1532.405 ;
        RECT 2440.005 1532.315 2440.355 1532.405 ;
        RECT 2424.500 1531.920 2424.730 1531.925 ;
        RECT 2425.500 1531.940 2425.850 1532.290 ;
        RECT 2434.055 1532.175 2434.405 1532.245 ;
        RECT 2439.490 1532.175 2439.815 1532.265 ;
        RECT 2433.850 1532.145 2434.405 1532.175 ;
        RECT 2439.465 1532.145 2439.815 1532.175 ;
        RECT 2433.680 1532.140 2434.405 1532.145 ;
        RECT 2439.295 1532.140 2439.815 1532.145 ;
        RECT 2433.680 1531.975 2439.815 1532.140 ;
        RECT 2433.850 1531.970 2439.815 1531.975 ;
        RECT 2433.850 1531.945 2434.405 1531.970 ;
        RECT 2439.465 1531.945 2439.815 1531.970 ;
        RECT 2425.500 1531.920 2425.845 1531.940 ;
        RECT 2409.170 1531.680 2409.460 1531.845 ;
        RECT 2422.365 1531.815 2422.685 1531.830 ;
        RECT 2422.340 1531.785 2422.685 1531.815 ;
        RECT 2422.165 1531.615 2422.685 1531.785 ;
        RECT 2424.500 1531.685 2424.790 1531.920 ;
        RECT 2425.495 1531.845 2425.845 1531.920 ;
        RECT 2434.055 1531.895 2434.405 1531.945 ;
        RECT 2439.490 1531.940 2439.815 1531.945 ;
        RECT 2440.885 1531.925 2441.055 1533.025 ;
        RECT 2441.820 1533.020 2442.115 1533.280 ;
        RECT 2441.850 1532.980 2442.115 1533.020 ;
        RECT 2441.850 1532.910 2442.175 1532.980 ;
        RECT 2441.850 1532.560 2442.200 1532.910 ;
        RECT 2440.825 1531.920 2441.055 1531.925 ;
        RECT 2441.880 1531.920 2442.050 1532.560 ;
        RECT 2425.495 1531.680 2425.785 1531.845 ;
        RECT 2438.690 1531.815 2439.010 1531.830 ;
        RECT 2438.665 1531.785 2439.010 1531.815 ;
        RECT 2438.490 1531.615 2439.010 1531.785 ;
        RECT 2440.825 1531.685 2441.115 1531.920 ;
        RECT 2441.820 1531.915 2442.050 1531.920 ;
        RECT 2441.820 1531.680 2442.110 1531.915 ;
        RECT 2359.135 1531.570 2359.485 1531.615 ;
        RECT 2373.365 1531.585 2373.710 1531.615 ;
        RECT 2389.690 1531.585 2390.035 1531.615 ;
        RECT 2406.015 1531.585 2406.360 1531.615 ;
        RECT 2422.340 1531.585 2422.685 1531.615 ;
        RECT 2438.665 1531.585 2439.010 1531.615 ;
        RECT 2373.390 1531.540 2373.710 1531.585 ;
        RECT 2389.715 1531.540 2390.035 1531.585 ;
        RECT 2406.040 1531.540 2406.360 1531.585 ;
        RECT 2422.365 1531.540 2422.685 1531.585 ;
        RECT 2438.690 1531.540 2439.010 1531.585 ;
        RECT 2362.285 1527.955 2362.575 1527.995 ;
        RECT 2362.985 1527.955 2363.305 1528.015 ;
        RECT 2362.285 1527.815 2363.305 1527.955 ;
        RECT 2362.285 1527.765 2362.615 1527.815 ;
        RECT 2362.985 1527.755 2363.305 1527.815 ;
        RECT 2368.125 1527.955 2368.415 1527.995 ;
        RECT 2368.125 1527.765 2368.455 1527.955 ;
        RECT 2363.485 1527.675 2363.775 1527.715 ;
        RECT 2364.705 1527.675 2365.025 1527.735 ;
        RECT 2365.545 1527.715 2365.865 1527.735 ;
        RECT 2365.545 1527.675 2365.975 1527.715 ;
        RECT 2363.485 1527.485 2363.935 1527.675 ;
        RECT 2361.785 1527.195 2362.105 1527.455 ;
        RECT 2362.745 1527.435 2363.065 1527.455 ;
        RECT 2362.745 1527.205 2363.295 1527.435 ;
        RECT 2363.795 1527.255 2363.935 1527.485 ;
        RECT 2364.705 1527.535 2365.975 1527.675 ;
        RECT 2364.705 1527.475 2365.025 1527.535 ;
        RECT 2365.545 1527.485 2365.975 1527.535 ;
        RECT 2365.545 1527.475 2365.865 1527.485 ;
        RECT 2362.745 1527.195 2363.065 1527.205 ;
        RECT 2361.875 1526.275 2362.015 1527.195 ;
        RECT 2363.435 1527.115 2363.935 1527.255 ;
        RECT 2364.245 1527.205 2364.535 1527.435 ;
        RECT 2362.745 1526.875 2363.065 1526.895 ;
        RECT 2362.745 1526.645 2363.295 1526.875 ;
        RECT 2362.745 1526.635 2363.065 1526.645 ;
        RECT 2363.435 1526.335 2363.575 1527.115 ;
        RECT 2364.315 1526.895 2364.455 1527.205 ;
        RECT 2365.515 1527.155 2368.095 1527.255 ;
        RECT 2365.445 1527.115 2368.175 1527.155 ;
        RECT 2365.445 1526.925 2366.105 1527.115 ;
        RECT 2367.885 1526.925 2368.175 1527.115 ;
        RECT 2365.785 1526.915 2366.105 1526.925 ;
        RECT 2363.965 1526.875 2364.455 1526.895 ;
        RECT 2363.725 1526.645 2364.455 1526.875 ;
        RECT 2363.965 1526.635 2364.455 1526.645 ;
        RECT 2364.945 1526.635 2365.265 1526.895 ;
        RECT 2366.785 1526.875 2367.105 1526.895 ;
        RECT 2366.785 1526.645 2367.215 1526.875 ;
        RECT 2366.785 1526.635 2367.105 1526.645 ;
        RECT 2367.385 1526.635 2367.705 1526.895 ;
        RECT 2362.285 1526.275 2362.575 1526.315 ;
        RECT 2361.875 1526.135 2362.575 1526.275 ;
        RECT 2362.285 1526.085 2362.575 1526.135 ;
        RECT 2363.225 1526.135 2363.575 1526.335 ;
        RECT 2364.315 1526.275 2364.455 1526.635 ;
        RECT 2365.425 1526.555 2365.745 1526.615 ;
        RECT 2368.315 1526.595 2368.455 1527.765 ;
        RECT 2369.125 1527.735 2369.415 1527.995 ;
        RECT 2378.610 1527.955 2378.900 1527.995 ;
        RECT 2379.310 1527.955 2379.630 1528.015 ;
        RECT 2378.610 1527.815 2379.630 1527.955 ;
        RECT 2378.610 1527.765 2378.940 1527.815 ;
        RECT 2379.310 1527.755 2379.630 1527.815 ;
        RECT 2384.450 1527.955 2384.740 1527.995 ;
        RECT 2384.450 1527.765 2384.780 1527.955 ;
        RECT 2369.105 1527.475 2369.425 1527.735 ;
        RECT 2379.810 1527.675 2380.100 1527.715 ;
        RECT 2381.030 1527.675 2381.350 1527.735 ;
        RECT 2381.870 1527.715 2382.190 1527.735 ;
        RECT 2381.870 1527.675 2382.300 1527.715 ;
        RECT 2379.810 1527.485 2380.260 1527.675 ;
        RECT 2378.110 1527.195 2378.430 1527.455 ;
        RECT 2379.070 1527.435 2379.390 1527.455 ;
        RECT 2379.070 1527.205 2379.620 1527.435 ;
        RECT 2380.120 1527.255 2380.260 1527.485 ;
        RECT 2381.030 1527.535 2382.300 1527.675 ;
        RECT 2381.030 1527.475 2381.350 1527.535 ;
        RECT 2381.870 1527.485 2382.300 1527.535 ;
        RECT 2381.870 1527.475 2382.190 1527.485 ;
        RECT 2379.070 1527.195 2379.390 1527.205 ;
        RECT 2369.225 1526.875 2369.545 1526.895 ;
        RECT 2373.390 1526.875 2373.710 1526.980 ;
        RECT 2369.225 1526.635 2369.695 1526.875 ;
        RECT 2369.845 1526.835 2370.135 1526.875 ;
        RECT 2373.365 1526.860 2373.710 1526.875 ;
        RECT 2373.360 1526.845 2373.710 1526.860 ;
        RECT 2369.845 1526.695 2370.295 1526.835 ;
        RECT 2369.845 1526.645 2370.775 1526.695 ;
        RECT 2373.190 1526.675 2373.710 1526.845 ;
        RECT 2373.365 1526.660 2373.710 1526.675 ;
        RECT 2373.365 1526.645 2373.655 1526.660 ;
        RECT 2365.925 1526.555 2366.215 1526.595 ;
        RECT 2368.315 1526.555 2368.655 1526.595 ;
        RECT 2365.425 1526.415 2366.215 1526.555 ;
        RECT 2365.425 1526.355 2365.745 1526.415 ;
        RECT 2365.925 1526.365 2366.215 1526.415 ;
        RECT 2367.955 1526.415 2368.655 1526.555 ;
        RECT 2367.955 1526.395 2368.095 1526.415 ;
        RECT 2366.495 1526.335 2368.095 1526.395 ;
        RECT 2368.365 1526.365 2368.655 1526.415 ;
        RECT 2369.555 1526.395 2369.695 1526.635 ;
        RECT 2370.155 1526.615 2370.775 1526.645 ;
        RECT 2370.155 1526.555 2370.865 1526.615 ;
        RECT 2364.725 1526.275 2365.015 1526.315 ;
        RECT 2364.315 1526.135 2365.015 1526.275 ;
        RECT 2363.225 1526.075 2363.545 1526.135 ;
        RECT 2364.725 1526.085 2365.015 1526.135 ;
        RECT 2366.405 1526.255 2368.095 1526.335 ;
        RECT 2368.845 1526.315 2369.165 1526.335 ;
        RECT 2366.405 1526.085 2366.975 1526.255 ;
        RECT 2368.845 1526.085 2369.415 1526.315 ;
        RECT 2369.555 1526.275 2369.815 1526.395 ;
        RECT 2370.545 1526.355 2370.865 1526.555 ;
        RECT 2374.165 1526.490 2374.515 1526.610 ;
        RECT 2375.525 1526.540 2375.815 1526.775 ;
        RECT 2376.515 1526.545 2376.805 1526.780 ;
        RECT 2376.515 1526.540 2376.745 1526.545 ;
        RECT 2375.525 1526.535 2375.755 1526.540 ;
        RECT 2371.860 1526.320 2374.515 1526.490 ;
        RECT 2370.085 1526.275 2370.375 1526.315 ;
        RECT 2369.555 1526.255 2370.375 1526.275 ;
        RECT 2369.675 1526.135 2370.375 1526.255 ;
        RECT 2370.085 1526.085 2370.375 1526.135 ;
        RECT 2371.860 1526.105 2372.030 1526.320 ;
        RECT 2373.995 1526.315 2374.515 1526.320 ;
        RECT 2374.165 1526.260 2374.515 1526.315 ;
        RECT 2373.735 1526.120 2374.025 1526.145 ;
        RECT 2374.705 1526.120 2375.055 1526.145 ;
        RECT 2366.405 1526.075 2366.725 1526.085 ;
        RECT 2368.845 1526.075 2369.165 1526.085 ;
        RECT 2371.770 1525.755 2372.110 1526.105 ;
        RECT 2373.735 1525.950 2375.055 1526.120 ;
        RECT 2373.735 1525.915 2374.025 1525.950 ;
        RECT 2373.795 1525.405 2373.965 1525.915 ;
        RECT 2374.705 1525.855 2375.055 1525.950 ;
        RECT 2375.585 1525.435 2375.755 1526.535 ;
        RECT 2376.575 1525.440 2376.745 1526.540 ;
        RECT 2378.200 1526.275 2378.340 1527.195 ;
        RECT 2379.760 1527.115 2380.260 1527.255 ;
        RECT 2380.570 1527.205 2380.860 1527.435 ;
        RECT 2379.070 1526.875 2379.390 1526.895 ;
        RECT 2379.070 1526.645 2379.620 1526.875 ;
        RECT 2379.070 1526.635 2379.390 1526.645 ;
        RECT 2379.760 1526.335 2379.900 1527.115 ;
        RECT 2380.640 1526.895 2380.780 1527.205 ;
        RECT 2381.840 1527.155 2384.420 1527.255 ;
        RECT 2381.770 1527.115 2384.500 1527.155 ;
        RECT 2381.770 1526.925 2382.430 1527.115 ;
        RECT 2384.210 1526.925 2384.500 1527.115 ;
        RECT 2382.110 1526.915 2382.430 1526.925 ;
        RECT 2380.290 1526.875 2380.780 1526.895 ;
        RECT 2380.050 1526.645 2380.780 1526.875 ;
        RECT 2380.290 1526.635 2380.780 1526.645 ;
        RECT 2381.270 1526.635 2381.590 1526.895 ;
        RECT 2383.110 1526.875 2383.430 1526.895 ;
        RECT 2383.110 1526.645 2383.540 1526.875 ;
        RECT 2383.110 1526.635 2383.430 1526.645 ;
        RECT 2383.710 1526.635 2384.030 1526.895 ;
        RECT 2378.610 1526.275 2378.900 1526.315 ;
        RECT 2378.200 1526.135 2378.900 1526.275 ;
        RECT 2378.610 1526.085 2378.900 1526.135 ;
        RECT 2379.550 1526.135 2379.900 1526.335 ;
        RECT 2380.640 1526.275 2380.780 1526.635 ;
        RECT 2381.750 1526.555 2382.070 1526.615 ;
        RECT 2384.640 1526.595 2384.780 1527.765 ;
        RECT 2385.450 1527.735 2385.740 1527.995 ;
        RECT 2394.935 1527.955 2395.225 1527.995 ;
        RECT 2395.635 1527.955 2395.955 1528.015 ;
        RECT 2394.935 1527.815 2395.955 1527.955 ;
        RECT 2394.935 1527.765 2395.265 1527.815 ;
        RECT 2395.635 1527.755 2395.955 1527.815 ;
        RECT 2400.775 1527.955 2401.065 1527.995 ;
        RECT 2400.775 1527.765 2401.105 1527.955 ;
        RECT 2385.430 1527.475 2385.750 1527.735 ;
        RECT 2396.135 1527.675 2396.425 1527.715 ;
        RECT 2397.355 1527.675 2397.675 1527.735 ;
        RECT 2398.195 1527.715 2398.515 1527.735 ;
        RECT 2398.195 1527.675 2398.625 1527.715 ;
        RECT 2396.135 1527.485 2396.585 1527.675 ;
        RECT 2392.990 1527.225 2393.310 1527.240 ;
        RECT 2392.840 1526.995 2393.310 1527.225 ;
        RECT 2394.435 1527.195 2394.755 1527.455 ;
        RECT 2395.395 1527.435 2395.715 1527.455 ;
        RECT 2395.395 1527.205 2395.945 1527.435 ;
        RECT 2396.445 1527.255 2396.585 1527.485 ;
        RECT 2397.355 1527.535 2398.625 1527.675 ;
        RECT 2397.355 1527.475 2397.675 1527.535 ;
        RECT 2398.195 1527.485 2398.625 1527.535 ;
        RECT 2398.195 1527.475 2398.515 1527.485 ;
        RECT 2395.395 1527.195 2395.715 1527.205 ;
        RECT 2392.990 1526.980 2393.310 1526.995 ;
        RECT 2385.550 1526.875 2385.870 1526.895 ;
        RECT 2389.715 1526.875 2390.035 1526.980 ;
        RECT 2385.550 1526.635 2386.020 1526.875 ;
        RECT 2386.170 1526.835 2386.460 1526.875 ;
        RECT 2389.690 1526.860 2390.035 1526.875 ;
        RECT 2389.685 1526.845 2390.035 1526.860 ;
        RECT 2386.170 1526.695 2386.620 1526.835 ;
        RECT 2386.170 1526.645 2387.100 1526.695 ;
        RECT 2389.515 1526.675 2390.035 1526.845 ;
        RECT 2389.690 1526.660 2390.035 1526.675 ;
        RECT 2389.690 1526.645 2389.980 1526.660 ;
        RECT 2382.250 1526.555 2382.540 1526.595 ;
        RECT 2384.640 1526.555 2384.980 1526.595 ;
        RECT 2381.750 1526.415 2382.540 1526.555 ;
        RECT 2381.750 1526.355 2382.070 1526.415 ;
        RECT 2382.250 1526.365 2382.540 1526.415 ;
        RECT 2384.280 1526.415 2384.980 1526.555 ;
        RECT 2384.280 1526.395 2384.420 1526.415 ;
        RECT 2382.820 1526.335 2384.420 1526.395 ;
        RECT 2384.690 1526.365 2384.980 1526.415 ;
        RECT 2385.880 1526.395 2386.020 1526.635 ;
        RECT 2386.480 1526.615 2387.100 1526.645 ;
        RECT 2386.480 1526.555 2387.190 1526.615 ;
        RECT 2381.050 1526.275 2381.340 1526.315 ;
        RECT 2380.640 1526.135 2381.340 1526.275 ;
        RECT 2379.550 1526.075 2379.870 1526.135 ;
        RECT 2381.050 1526.085 2381.340 1526.135 ;
        RECT 2382.730 1526.255 2384.420 1526.335 ;
        RECT 2385.170 1526.315 2385.490 1526.335 ;
        RECT 2382.730 1526.085 2383.300 1526.255 ;
        RECT 2385.170 1526.085 2385.740 1526.315 ;
        RECT 2385.880 1526.275 2386.140 1526.395 ;
        RECT 2386.870 1526.355 2387.190 1526.555 ;
        RECT 2390.490 1526.490 2390.840 1526.610 ;
        RECT 2391.850 1526.540 2392.140 1526.775 ;
        RECT 2392.840 1526.545 2393.130 1526.780 ;
        RECT 2392.840 1526.540 2393.070 1526.545 ;
        RECT 2391.850 1526.535 2392.080 1526.540 ;
        RECT 2388.185 1526.320 2390.840 1526.490 ;
        RECT 2386.410 1526.275 2386.700 1526.315 ;
        RECT 2385.880 1526.255 2386.700 1526.275 ;
        RECT 2386.000 1526.135 2386.700 1526.255 ;
        RECT 2386.410 1526.085 2386.700 1526.135 ;
        RECT 2388.185 1526.105 2388.355 1526.320 ;
        RECT 2390.320 1526.315 2390.840 1526.320 ;
        RECT 2390.490 1526.260 2390.840 1526.315 ;
        RECT 2390.060 1526.120 2390.350 1526.145 ;
        RECT 2391.030 1526.120 2391.380 1526.145 ;
        RECT 2382.730 1526.075 2383.050 1526.085 ;
        RECT 2385.170 1526.075 2385.490 1526.085 ;
        RECT 2388.095 1525.755 2388.435 1526.105 ;
        RECT 2390.060 1525.950 2391.380 1526.120 ;
        RECT 2390.060 1525.915 2390.350 1525.950 ;
        RECT 2373.735 1525.175 2374.025 1525.405 ;
        RECT 2375.525 1525.175 2375.820 1525.435 ;
        RECT 2376.430 1525.180 2376.810 1525.440 ;
        RECT 2390.120 1525.405 2390.290 1525.915 ;
        RECT 2391.030 1525.855 2391.380 1525.950 ;
        RECT 2391.910 1525.435 2392.080 1526.535 ;
        RECT 2392.900 1525.440 2393.070 1526.540 ;
        RECT 2394.525 1526.275 2394.665 1527.195 ;
        RECT 2396.085 1527.115 2396.585 1527.255 ;
        RECT 2396.895 1527.205 2397.185 1527.435 ;
        RECT 2395.395 1526.875 2395.715 1526.895 ;
        RECT 2395.395 1526.645 2395.945 1526.875 ;
        RECT 2395.395 1526.635 2395.715 1526.645 ;
        RECT 2396.085 1526.335 2396.225 1527.115 ;
        RECT 2396.965 1526.895 2397.105 1527.205 ;
        RECT 2398.165 1527.155 2400.745 1527.255 ;
        RECT 2398.095 1527.115 2400.825 1527.155 ;
        RECT 2398.095 1526.925 2398.755 1527.115 ;
        RECT 2400.535 1526.925 2400.825 1527.115 ;
        RECT 2398.435 1526.915 2398.755 1526.925 ;
        RECT 2396.615 1526.875 2397.105 1526.895 ;
        RECT 2396.375 1526.645 2397.105 1526.875 ;
        RECT 2396.615 1526.635 2397.105 1526.645 ;
        RECT 2397.595 1526.635 2397.915 1526.895 ;
        RECT 2399.435 1526.875 2399.755 1526.895 ;
        RECT 2399.435 1526.645 2399.865 1526.875 ;
        RECT 2399.435 1526.635 2399.755 1526.645 ;
        RECT 2400.035 1526.635 2400.355 1526.895 ;
        RECT 2394.935 1526.275 2395.225 1526.315 ;
        RECT 2394.525 1526.135 2395.225 1526.275 ;
        RECT 2394.935 1526.085 2395.225 1526.135 ;
        RECT 2395.875 1526.135 2396.225 1526.335 ;
        RECT 2396.965 1526.275 2397.105 1526.635 ;
        RECT 2398.075 1526.555 2398.395 1526.615 ;
        RECT 2400.965 1526.595 2401.105 1527.765 ;
        RECT 2401.775 1527.735 2402.065 1527.995 ;
        RECT 2411.260 1527.955 2411.550 1527.995 ;
        RECT 2411.960 1527.955 2412.280 1528.015 ;
        RECT 2411.260 1527.815 2412.280 1527.955 ;
        RECT 2411.260 1527.765 2411.590 1527.815 ;
        RECT 2411.960 1527.755 2412.280 1527.815 ;
        RECT 2417.100 1527.955 2417.390 1527.995 ;
        RECT 2417.100 1527.765 2417.430 1527.955 ;
        RECT 2401.755 1527.475 2402.075 1527.735 ;
        RECT 2412.460 1527.675 2412.750 1527.715 ;
        RECT 2413.680 1527.675 2414.000 1527.735 ;
        RECT 2414.520 1527.715 2414.840 1527.735 ;
        RECT 2414.520 1527.675 2414.950 1527.715 ;
        RECT 2412.460 1527.485 2412.910 1527.675 ;
        RECT 2410.760 1527.195 2411.080 1527.455 ;
        RECT 2411.720 1527.435 2412.040 1527.455 ;
        RECT 2411.720 1527.205 2412.270 1527.435 ;
        RECT 2412.770 1527.255 2412.910 1527.485 ;
        RECT 2413.680 1527.535 2414.950 1527.675 ;
        RECT 2413.680 1527.475 2414.000 1527.535 ;
        RECT 2414.520 1527.485 2414.950 1527.535 ;
        RECT 2414.520 1527.475 2414.840 1527.485 ;
        RECT 2411.720 1527.195 2412.040 1527.205 ;
        RECT 2401.875 1526.875 2402.195 1526.895 ;
        RECT 2406.040 1526.875 2406.360 1526.980 ;
        RECT 2401.875 1526.635 2402.345 1526.875 ;
        RECT 2402.495 1526.835 2402.785 1526.875 ;
        RECT 2406.015 1526.860 2406.360 1526.875 ;
        RECT 2406.010 1526.845 2406.360 1526.860 ;
        RECT 2402.495 1526.695 2402.945 1526.835 ;
        RECT 2402.495 1526.645 2403.425 1526.695 ;
        RECT 2405.840 1526.675 2406.360 1526.845 ;
        RECT 2406.015 1526.660 2406.360 1526.675 ;
        RECT 2406.015 1526.645 2406.305 1526.660 ;
        RECT 2398.575 1526.555 2398.865 1526.595 ;
        RECT 2400.965 1526.555 2401.305 1526.595 ;
        RECT 2398.075 1526.415 2398.865 1526.555 ;
        RECT 2398.075 1526.355 2398.395 1526.415 ;
        RECT 2398.575 1526.365 2398.865 1526.415 ;
        RECT 2400.605 1526.415 2401.305 1526.555 ;
        RECT 2400.605 1526.395 2400.745 1526.415 ;
        RECT 2399.145 1526.335 2400.745 1526.395 ;
        RECT 2401.015 1526.365 2401.305 1526.415 ;
        RECT 2402.205 1526.395 2402.345 1526.635 ;
        RECT 2402.805 1526.615 2403.425 1526.645 ;
        RECT 2402.805 1526.555 2403.515 1526.615 ;
        RECT 2397.375 1526.275 2397.665 1526.315 ;
        RECT 2396.965 1526.135 2397.665 1526.275 ;
        RECT 2395.875 1526.075 2396.195 1526.135 ;
        RECT 2397.375 1526.085 2397.665 1526.135 ;
        RECT 2399.055 1526.255 2400.745 1526.335 ;
        RECT 2401.495 1526.315 2401.815 1526.335 ;
        RECT 2399.055 1526.085 2399.625 1526.255 ;
        RECT 2401.495 1526.085 2402.065 1526.315 ;
        RECT 2402.205 1526.275 2402.465 1526.395 ;
        RECT 2403.195 1526.355 2403.515 1526.555 ;
        RECT 2406.815 1526.490 2407.165 1526.610 ;
        RECT 2408.175 1526.540 2408.465 1526.775 ;
        RECT 2409.165 1526.545 2409.455 1526.780 ;
        RECT 2409.165 1526.540 2409.395 1526.545 ;
        RECT 2408.175 1526.535 2408.405 1526.540 ;
        RECT 2404.510 1526.320 2407.165 1526.490 ;
        RECT 2402.735 1526.275 2403.025 1526.315 ;
        RECT 2402.205 1526.255 2403.025 1526.275 ;
        RECT 2402.325 1526.135 2403.025 1526.255 ;
        RECT 2402.735 1526.085 2403.025 1526.135 ;
        RECT 2404.510 1526.105 2404.680 1526.320 ;
        RECT 2406.645 1526.315 2407.165 1526.320 ;
        RECT 2406.815 1526.260 2407.165 1526.315 ;
        RECT 2406.385 1526.120 2406.675 1526.145 ;
        RECT 2407.355 1526.120 2407.705 1526.145 ;
        RECT 2399.055 1526.075 2399.375 1526.085 ;
        RECT 2401.495 1526.075 2401.815 1526.085 ;
        RECT 2404.420 1525.755 2404.760 1526.105 ;
        RECT 2406.385 1525.950 2407.705 1526.120 ;
        RECT 2406.385 1525.915 2406.675 1525.950 ;
        RECT 2390.060 1525.175 2390.350 1525.405 ;
        RECT 2391.850 1525.175 2392.145 1525.435 ;
        RECT 2392.840 1525.180 2393.135 1525.440 ;
        RECT 2406.445 1525.405 2406.615 1525.915 ;
        RECT 2407.355 1525.855 2407.705 1525.950 ;
        RECT 2408.235 1525.435 2408.405 1526.535 ;
        RECT 2409.225 1525.440 2409.395 1526.540 ;
        RECT 2410.850 1526.275 2410.990 1527.195 ;
        RECT 2412.410 1527.115 2412.910 1527.255 ;
        RECT 2413.220 1527.205 2413.510 1527.435 ;
        RECT 2411.720 1526.875 2412.040 1526.895 ;
        RECT 2411.720 1526.645 2412.270 1526.875 ;
        RECT 2411.720 1526.635 2412.040 1526.645 ;
        RECT 2412.410 1526.335 2412.550 1527.115 ;
        RECT 2413.290 1526.895 2413.430 1527.205 ;
        RECT 2414.490 1527.155 2417.070 1527.255 ;
        RECT 2414.420 1527.115 2417.150 1527.155 ;
        RECT 2414.420 1526.925 2415.080 1527.115 ;
        RECT 2416.860 1526.925 2417.150 1527.115 ;
        RECT 2414.760 1526.915 2415.080 1526.925 ;
        RECT 2412.940 1526.875 2413.430 1526.895 ;
        RECT 2412.700 1526.645 2413.430 1526.875 ;
        RECT 2412.940 1526.635 2413.430 1526.645 ;
        RECT 2413.920 1526.635 2414.240 1526.895 ;
        RECT 2415.760 1526.875 2416.080 1526.895 ;
        RECT 2415.760 1526.645 2416.190 1526.875 ;
        RECT 2415.760 1526.635 2416.080 1526.645 ;
        RECT 2416.360 1526.635 2416.680 1526.895 ;
        RECT 2411.260 1526.275 2411.550 1526.315 ;
        RECT 2410.850 1526.135 2411.550 1526.275 ;
        RECT 2411.260 1526.085 2411.550 1526.135 ;
        RECT 2412.200 1526.135 2412.550 1526.335 ;
        RECT 2413.290 1526.275 2413.430 1526.635 ;
        RECT 2414.400 1526.555 2414.720 1526.615 ;
        RECT 2417.290 1526.595 2417.430 1527.765 ;
        RECT 2418.100 1527.735 2418.390 1527.995 ;
        RECT 2427.585 1527.955 2427.875 1527.995 ;
        RECT 2428.285 1527.955 2428.605 1528.015 ;
        RECT 2427.585 1527.815 2428.605 1527.955 ;
        RECT 2427.585 1527.765 2427.915 1527.815 ;
        RECT 2428.285 1527.755 2428.605 1527.815 ;
        RECT 2433.425 1527.955 2433.715 1527.995 ;
        RECT 2433.425 1527.765 2433.755 1527.955 ;
        RECT 2418.080 1527.475 2418.400 1527.735 ;
        RECT 2428.785 1527.675 2429.075 1527.715 ;
        RECT 2430.005 1527.675 2430.325 1527.735 ;
        RECT 2430.845 1527.715 2431.165 1527.735 ;
        RECT 2430.845 1527.675 2431.275 1527.715 ;
        RECT 2428.785 1527.485 2429.235 1527.675 ;
        RECT 2425.650 1527.225 2425.970 1527.240 ;
        RECT 2425.490 1526.995 2425.970 1527.225 ;
        RECT 2427.085 1527.195 2427.405 1527.455 ;
        RECT 2428.045 1527.435 2428.365 1527.455 ;
        RECT 2428.045 1527.205 2428.595 1527.435 ;
        RECT 2429.095 1527.255 2429.235 1527.485 ;
        RECT 2430.005 1527.535 2431.275 1527.675 ;
        RECT 2430.005 1527.475 2430.325 1527.535 ;
        RECT 2430.845 1527.485 2431.275 1527.535 ;
        RECT 2430.845 1527.475 2431.165 1527.485 ;
        RECT 2428.045 1527.195 2428.365 1527.205 ;
        RECT 2425.650 1526.980 2425.970 1526.995 ;
        RECT 2418.200 1526.875 2418.520 1526.895 ;
        RECT 2422.365 1526.875 2422.685 1526.980 ;
        RECT 2418.200 1526.635 2418.670 1526.875 ;
        RECT 2418.820 1526.835 2419.110 1526.875 ;
        RECT 2422.340 1526.860 2422.685 1526.875 ;
        RECT 2422.335 1526.845 2422.685 1526.860 ;
        RECT 2418.820 1526.695 2419.270 1526.835 ;
        RECT 2418.820 1526.645 2419.750 1526.695 ;
        RECT 2422.165 1526.675 2422.685 1526.845 ;
        RECT 2422.340 1526.660 2422.685 1526.675 ;
        RECT 2422.340 1526.645 2422.630 1526.660 ;
        RECT 2414.900 1526.555 2415.190 1526.595 ;
        RECT 2417.290 1526.555 2417.630 1526.595 ;
        RECT 2414.400 1526.415 2415.190 1526.555 ;
        RECT 2414.400 1526.355 2414.720 1526.415 ;
        RECT 2414.900 1526.365 2415.190 1526.415 ;
        RECT 2416.930 1526.415 2417.630 1526.555 ;
        RECT 2416.930 1526.395 2417.070 1526.415 ;
        RECT 2415.470 1526.335 2417.070 1526.395 ;
        RECT 2417.340 1526.365 2417.630 1526.415 ;
        RECT 2418.530 1526.395 2418.670 1526.635 ;
        RECT 2419.130 1526.615 2419.750 1526.645 ;
        RECT 2419.130 1526.555 2419.840 1526.615 ;
        RECT 2413.700 1526.275 2413.990 1526.315 ;
        RECT 2413.290 1526.135 2413.990 1526.275 ;
        RECT 2412.200 1526.075 2412.520 1526.135 ;
        RECT 2413.700 1526.085 2413.990 1526.135 ;
        RECT 2415.380 1526.255 2417.070 1526.335 ;
        RECT 2417.820 1526.315 2418.140 1526.335 ;
        RECT 2415.380 1526.085 2415.950 1526.255 ;
        RECT 2417.820 1526.085 2418.390 1526.315 ;
        RECT 2418.530 1526.275 2418.790 1526.395 ;
        RECT 2419.520 1526.355 2419.840 1526.555 ;
        RECT 2423.140 1526.490 2423.490 1526.610 ;
        RECT 2424.500 1526.540 2424.790 1526.775 ;
        RECT 2425.490 1526.545 2425.780 1526.780 ;
        RECT 2425.490 1526.540 2425.720 1526.545 ;
        RECT 2424.500 1526.535 2424.730 1526.540 ;
        RECT 2420.835 1526.320 2423.490 1526.490 ;
        RECT 2419.060 1526.275 2419.350 1526.315 ;
        RECT 2418.530 1526.255 2419.350 1526.275 ;
        RECT 2418.650 1526.135 2419.350 1526.255 ;
        RECT 2419.060 1526.085 2419.350 1526.135 ;
        RECT 2420.835 1526.105 2421.005 1526.320 ;
        RECT 2422.970 1526.315 2423.490 1526.320 ;
        RECT 2423.140 1526.260 2423.490 1526.315 ;
        RECT 2422.710 1526.120 2423.000 1526.145 ;
        RECT 2423.680 1526.120 2424.030 1526.145 ;
        RECT 2415.380 1526.075 2415.700 1526.085 ;
        RECT 2417.820 1526.075 2418.140 1526.085 ;
        RECT 2420.745 1525.755 2421.085 1526.105 ;
        RECT 2422.710 1525.950 2424.030 1526.120 ;
        RECT 2422.710 1525.915 2423.000 1525.950 ;
        RECT 2406.385 1525.175 2406.675 1525.405 ;
        RECT 2408.175 1525.175 2408.470 1525.435 ;
        RECT 2409.090 1525.180 2409.460 1525.440 ;
        RECT 2422.770 1525.405 2422.940 1525.915 ;
        RECT 2423.680 1525.855 2424.030 1525.950 ;
        RECT 2424.560 1525.435 2424.730 1526.535 ;
        RECT 2425.550 1525.440 2425.720 1526.540 ;
        RECT 2427.175 1526.275 2427.315 1527.195 ;
        RECT 2428.735 1527.115 2429.235 1527.255 ;
        RECT 2429.545 1527.205 2429.835 1527.435 ;
        RECT 2428.045 1526.875 2428.365 1526.895 ;
        RECT 2428.045 1526.645 2428.595 1526.875 ;
        RECT 2428.045 1526.635 2428.365 1526.645 ;
        RECT 2428.735 1526.335 2428.875 1527.115 ;
        RECT 2429.615 1526.895 2429.755 1527.205 ;
        RECT 2430.815 1527.155 2433.395 1527.255 ;
        RECT 2430.745 1527.115 2433.475 1527.155 ;
        RECT 2430.745 1526.925 2431.405 1527.115 ;
        RECT 2433.185 1526.925 2433.475 1527.115 ;
        RECT 2431.085 1526.915 2431.405 1526.925 ;
        RECT 2429.265 1526.875 2429.755 1526.895 ;
        RECT 2429.025 1526.645 2429.755 1526.875 ;
        RECT 2429.265 1526.635 2429.755 1526.645 ;
        RECT 2430.245 1526.635 2430.565 1526.895 ;
        RECT 2432.085 1526.875 2432.405 1526.895 ;
        RECT 2432.085 1526.645 2432.515 1526.875 ;
        RECT 2432.085 1526.635 2432.405 1526.645 ;
        RECT 2432.685 1526.635 2433.005 1526.895 ;
        RECT 2427.585 1526.275 2427.875 1526.315 ;
        RECT 2427.175 1526.135 2427.875 1526.275 ;
        RECT 2427.585 1526.085 2427.875 1526.135 ;
        RECT 2428.525 1526.135 2428.875 1526.335 ;
        RECT 2429.615 1526.275 2429.755 1526.635 ;
        RECT 2430.725 1526.555 2431.045 1526.615 ;
        RECT 2433.615 1526.595 2433.755 1527.765 ;
        RECT 2434.425 1527.735 2434.715 1527.995 ;
        RECT 2434.405 1527.475 2434.725 1527.735 ;
        RECT 2434.525 1526.875 2434.845 1526.895 ;
        RECT 2438.690 1526.875 2439.010 1526.980 ;
        RECT 2434.525 1526.635 2434.995 1526.875 ;
        RECT 2435.145 1526.835 2435.435 1526.875 ;
        RECT 2438.665 1526.860 2439.010 1526.875 ;
        RECT 2438.660 1526.845 2439.010 1526.860 ;
        RECT 2435.145 1526.695 2435.595 1526.835 ;
        RECT 2435.145 1526.645 2436.075 1526.695 ;
        RECT 2438.490 1526.675 2439.010 1526.845 ;
        RECT 2438.665 1526.660 2439.010 1526.675 ;
        RECT 2438.665 1526.645 2438.955 1526.660 ;
        RECT 2431.225 1526.555 2431.515 1526.595 ;
        RECT 2433.615 1526.555 2433.955 1526.595 ;
        RECT 2430.725 1526.415 2431.515 1526.555 ;
        RECT 2430.725 1526.355 2431.045 1526.415 ;
        RECT 2431.225 1526.365 2431.515 1526.415 ;
        RECT 2433.255 1526.415 2433.955 1526.555 ;
        RECT 2433.255 1526.395 2433.395 1526.415 ;
        RECT 2431.795 1526.335 2433.395 1526.395 ;
        RECT 2433.665 1526.365 2433.955 1526.415 ;
        RECT 2434.855 1526.395 2434.995 1526.635 ;
        RECT 2435.455 1526.615 2436.075 1526.645 ;
        RECT 2435.455 1526.555 2436.165 1526.615 ;
        RECT 2430.025 1526.275 2430.315 1526.315 ;
        RECT 2429.615 1526.135 2430.315 1526.275 ;
        RECT 2428.525 1526.075 2428.845 1526.135 ;
        RECT 2430.025 1526.085 2430.315 1526.135 ;
        RECT 2431.705 1526.255 2433.395 1526.335 ;
        RECT 2434.145 1526.315 2434.465 1526.335 ;
        RECT 2431.705 1526.085 2432.275 1526.255 ;
        RECT 2434.145 1526.085 2434.715 1526.315 ;
        RECT 2434.855 1526.275 2435.115 1526.395 ;
        RECT 2435.845 1526.355 2436.165 1526.555 ;
        RECT 2439.465 1526.490 2439.815 1526.610 ;
        RECT 2440.825 1526.540 2441.115 1526.775 ;
        RECT 2441.815 1526.545 2442.105 1526.780 ;
        RECT 2441.815 1526.540 2442.045 1526.545 ;
        RECT 2440.825 1526.535 2441.055 1526.540 ;
        RECT 2437.160 1526.320 2439.815 1526.490 ;
        RECT 2435.385 1526.275 2435.675 1526.315 ;
        RECT 2434.855 1526.255 2435.675 1526.275 ;
        RECT 2434.975 1526.135 2435.675 1526.255 ;
        RECT 2435.385 1526.085 2435.675 1526.135 ;
        RECT 2437.160 1526.105 2437.330 1526.320 ;
        RECT 2439.295 1526.315 2439.815 1526.320 ;
        RECT 2439.465 1526.260 2439.815 1526.315 ;
        RECT 2439.035 1526.120 2439.325 1526.145 ;
        RECT 2440.005 1526.120 2440.355 1526.145 ;
        RECT 2431.705 1526.075 2432.025 1526.085 ;
        RECT 2434.145 1526.075 2434.465 1526.085 ;
        RECT 2437.070 1525.755 2437.410 1526.105 ;
        RECT 2439.035 1525.950 2440.355 1526.120 ;
        RECT 2439.035 1525.915 2439.325 1525.950 ;
        RECT 2422.710 1525.175 2423.000 1525.405 ;
        RECT 2424.500 1525.175 2424.795 1525.435 ;
        RECT 2425.490 1525.180 2425.785 1525.440 ;
        RECT 2439.095 1525.405 2439.265 1525.915 ;
        RECT 2440.005 1525.855 2440.355 1525.950 ;
        RECT 2440.885 1525.435 2441.055 1526.535 ;
        RECT 2441.875 1525.440 2442.045 1526.540 ;
        RECT 2439.035 1525.175 2439.325 1525.405 ;
        RECT 2440.825 1525.175 2441.120 1525.435 ;
        RECT 2441.815 1525.380 2442.110 1525.440 ;
        RECT 2441.815 1525.240 2443.360 1525.380 ;
        RECT 2441.815 1525.180 2442.110 1525.240 ;
        RECT 2443.220 1525.140 2443.360 1525.240 ;
        RECT 2452.790 1525.140 2453.110 1525.200 ;
        RECT 2443.220 1525.000 2453.110 1525.140 ;
        RECT 2452.790 1524.940 2453.110 1525.000 ;
        RECT 2425.280 1518.200 2426.340 1518.340 ;
        RECT 2376.430 1517.800 2376.750 1518.060 ;
        RECT 2392.990 1518.000 2393.310 1518.060 ;
        RECT 2409.090 1518.000 2409.410 1518.060 ;
        RECT 2425.280 1518.000 2425.420 1518.200 ;
        RECT 2392.990 1517.860 2401.270 1518.000 ;
        RECT 2392.990 1517.800 2393.310 1517.860 ;
        RECT 2376.520 1516.980 2376.660 1517.800 ;
        RECT 2401.130 1517.320 2401.270 1517.860 ;
        RECT 2409.090 1517.860 2425.420 1518.000 ;
        RECT 2409.090 1517.800 2409.410 1517.860 ;
        RECT 2425.650 1517.800 2425.970 1518.060 ;
        RECT 2426.200 1518.000 2426.340 1518.200 ;
        RECT 2682.330 1518.000 2682.650 1518.060 ;
        RECT 2426.200 1517.860 2682.650 1518.000 ;
        RECT 2682.330 1517.800 2682.650 1517.860 ;
        RECT 2425.740 1517.660 2425.880 1517.800 ;
        RECT 2683.250 1517.660 2683.570 1517.720 ;
        RECT 2425.740 1517.520 2683.570 1517.660 ;
        RECT 2683.250 1517.460 2683.570 1517.520 ;
        RECT 2590.790 1517.320 2591.110 1517.380 ;
        RECT 2401.130 1517.180 2591.110 1517.320 ;
        RECT 2590.790 1517.120 2591.110 1517.180 ;
        RECT 2501.090 1516.980 2501.410 1517.040 ;
        RECT 2376.520 1516.840 2501.410 1516.980 ;
        RECT 2501.090 1516.780 2501.410 1516.840 ;
        RECT 2459.690 1504.060 2460.010 1504.120 ;
        RECT 2677.270 1504.060 2677.590 1504.120 ;
        RECT 2459.690 1503.920 2677.590 1504.060 ;
        RECT 2459.690 1503.860 2460.010 1503.920 ;
        RECT 2677.270 1503.860 2677.590 1503.920 ;
        RECT 2460.150 1497.260 2460.470 1497.320 ;
        RECT 2677.270 1497.260 2677.590 1497.320 ;
        RECT 2460.150 1497.120 2677.590 1497.260 ;
        RECT 2460.150 1497.060 2460.470 1497.120 ;
        RECT 2677.270 1497.060 2677.590 1497.120 ;
        RECT 2695.590 1496.480 2695.910 1496.540 ;
        RECT 2698.810 1496.480 2699.130 1496.540 ;
        RECT 2700.205 1496.480 2700.495 1496.525 ;
        RECT 2695.590 1496.340 2698.120 1496.480 ;
        RECT 2695.590 1496.280 2695.910 1496.340 ;
        RECT 2697.980 1496.140 2698.120 1496.340 ;
        RECT 2698.810 1496.340 2700.495 1496.480 ;
        RECT 2698.810 1496.280 2699.130 1496.340 ;
        RECT 2700.205 1496.295 2700.495 1496.340 ;
        RECT 2702.490 1496.480 2702.810 1496.540 ;
        RECT 2709.865 1496.480 2710.155 1496.525 ;
        RECT 2702.490 1496.340 2710.155 1496.480 ;
        RECT 2702.490 1496.280 2702.810 1496.340 ;
        RECT 2709.865 1496.295 2710.155 1496.340 ;
        RECT 2697.980 1496.000 2701.340 1496.140 ;
        RECT 2695.130 1495.800 2695.450 1495.860 ;
        RECT 2701.200 1495.845 2701.340 1496.000 ;
        RECT 2699.745 1495.800 2700.035 1495.845 ;
        RECT 2695.130 1495.660 2700.035 1495.800 ;
        RECT 2695.130 1495.600 2695.450 1495.660 ;
        RECT 2699.745 1495.615 2700.035 1495.660 ;
        RECT 2701.125 1495.615 2701.415 1495.845 ;
        RECT 2698.365 1495.460 2698.655 1495.505 ;
        RECT 2701.570 1495.460 2701.890 1495.520 ;
        RECT 2698.365 1495.320 2701.890 1495.460 ;
        RECT 2698.365 1495.275 2698.655 1495.320 ;
        RECT 2701.570 1495.260 2701.890 1495.320 ;
        RECT 2721.810 1494.920 2722.130 1495.180 ;
        RECT 2698.350 1494.780 2698.670 1494.840 ;
        RECT 2698.825 1494.780 2699.115 1494.825 ;
        RECT 2698.350 1494.640 2699.115 1494.780 ;
        RECT 2698.350 1494.580 2698.670 1494.640 ;
        RECT 2698.825 1494.595 2699.115 1494.640 ;
        RECT 2731.470 1494.580 2731.790 1494.840 ;
        RECT 2694.670 1492.740 2694.990 1492.800 ;
        RECT 2696.985 1492.740 2697.275 1492.785 ;
        RECT 2694.670 1492.600 2697.275 1492.740 ;
        RECT 2694.670 1492.540 2694.990 1492.600 ;
        RECT 2696.985 1492.555 2697.275 1492.600 ;
        RECT 2697.890 1491.860 2698.210 1492.120 ;
        RECT 2453.710 1490.460 2454.030 1490.520 ;
        RECT 2677.270 1490.460 2677.590 1490.520 ;
        RECT 2453.710 1490.320 2677.590 1490.460 ;
        RECT 2453.710 1490.260 2454.030 1490.320 ;
        RECT 2677.270 1490.260 2677.590 1490.320 ;
        RECT 2694.670 1484.920 2694.990 1484.980 ;
        RECT 2696.985 1484.920 2697.275 1484.965 ;
        RECT 2694.670 1484.780 2697.275 1484.920 ;
        RECT 2694.670 1484.720 2694.990 1484.780 ;
        RECT 2696.985 1484.735 2697.275 1484.780 ;
        RECT 2696.970 1483.900 2697.290 1483.960 ;
        RECT 2697.905 1483.900 2698.195 1483.945 ;
        RECT 2696.970 1483.760 2698.195 1483.900 ;
        RECT 2696.970 1483.700 2697.290 1483.760 ;
        RECT 2697.905 1483.715 2698.195 1483.760 ;
        RECT 2460.610 1483.320 2460.930 1483.380 ;
        RECT 2677.730 1483.320 2678.050 1483.380 ;
        RECT 2460.610 1483.180 2678.050 1483.320 ;
        RECT 2460.610 1483.120 2460.930 1483.180 ;
        RECT 2677.730 1483.120 2678.050 1483.180 ;
        RECT 2466.590 1482.980 2466.910 1483.040 ;
        RECT 2677.270 1482.980 2677.590 1483.040 ;
        RECT 2466.590 1482.840 2677.590 1482.980 ;
        RECT 2466.590 1482.780 2466.910 1482.840 ;
        RECT 2677.270 1482.780 2677.590 1482.840 ;
        RECT 2697.430 1482.200 2697.750 1482.260 ;
        RECT 2698.350 1482.200 2698.670 1482.260 ;
        RECT 2697.430 1482.060 2698.670 1482.200 ;
        RECT 2697.430 1482.000 2697.750 1482.060 ;
        RECT 2698.350 1482.000 2698.670 1482.060 ;
        RECT 2698.370 1479.820 2698.660 1479.865 ;
        RECT 2703.890 1479.820 2704.180 1479.865 ;
        RECT 2704.810 1479.820 2705.100 1479.865 ;
        RECT 2698.370 1479.680 2705.100 1479.820 ;
        RECT 2698.370 1479.635 2698.660 1479.680 ;
        RECT 2703.890 1479.635 2704.180 1479.680 ;
        RECT 2704.810 1479.635 2705.100 1479.680 ;
        RECT 2696.985 1479.480 2697.275 1479.525 ;
        RECT 2697.430 1479.480 2697.750 1479.540 ;
        RECT 2696.985 1479.340 2697.750 1479.480 ;
        RECT 2696.985 1479.295 2697.275 1479.340 ;
        RECT 2697.430 1479.280 2697.750 1479.340 ;
        RECT 2697.890 1479.280 2698.210 1479.540 ;
        RECT 2699.290 1479.480 2699.580 1479.525 ;
        RECT 2701.130 1479.480 2701.420 1479.525 ;
        RECT 2699.290 1479.340 2701.420 1479.480 ;
        RECT 2699.290 1479.295 2699.580 1479.340 ;
        RECT 2701.130 1479.295 2701.420 1479.340 ;
        RECT 2703.475 1479.480 2703.765 1479.525 ;
        RECT 2705.315 1479.480 2705.605 1479.525 ;
        RECT 2703.475 1479.340 2705.605 1479.480 ;
        RECT 2703.475 1479.295 2703.765 1479.340 ;
        RECT 2705.315 1479.295 2705.605 1479.340 ;
        RECT 2721.810 1479.280 2722.130 1479.540 ;
        RECT 2702.030 1479.185 2702.350 1479.200 ;
        RECT 2701.585 1479.140 2701.875 1479.185 ;
        RECT 2697.520 1479.000 2701.875 1479.140 ;
        RECT 2697.520 1478.860 2697.660 1479.000 ;
        RECT 2701.585 1478.955 2701.875 1479.000 ;
        RECT 2702.030 1478.955 2702.460 1479.185 ;
        RECT 2702.950 1479.140 2703.270 1479.200 ;
        RECT 2721.900 1479.140 2722.040 1479.280 ;
        RECT 2702.950 1479.000 2722.040 1479.140 ;
        RECT 2702.030 1478.940 2702.350 1478.955 ;
        RECT 2702.950 1478.940 2703.270 1479.000 ;
        RECT 2697.430 1478.600 2697.750 1478.860 ;
        RECT 2700.205 1478.615 2700.495 1478.845 ;
        RECT 2701.165 1478.800 2701.455 1478.845 ;
        RECT 2704.395 1478.800 2704.685 1478.845 ;
        RECT 2701.165 1478.660 2704.685 1478.800 ;
        RECT 2701.165 1478.615 2701.455 1478.660 ;
        RECT 2704.395 1478.615 2704.685 1478.660 ;
        RECT 2700.280 1478.460 2700.420 1478.615 ;
        RECT 2702.490 1478.460 2702.810 1478.520 ;
        RECT 2700.280 1478.320 2702.810 1478.460 ;
        RECT 2702.490 1478.260 2702.810 1478.320 ;
        RECT 2703.870 1478.460 2704.190 1478.520 ;
        RECT 2706.185 1478.460 2706.475 1478.505 ;
        RECT 2703.870 1478.320 2706.475 1478.460 ;
        RECT 2703.870 1478.260 2704.190 1478.320 ;
        RECT 2706.185 1478.275 2706.475 1478.320 ;
        RECT 2697.905 1477.440 2698.195 1477.485 ;
        RECT 2702.030 1477.440 2702.350 1477.500 ;
        RECT 2697.905 1477.300 2702.350 1477.440 ;
        RECT 2697.905 1477.255 2698.195 1477.300 ;
        RECT 2702.030 1477.240 2702.350 1477.300 ;
        RECT 2461.070 1476.520 2461.390 1476.580 ;
        RECT 2677.270 1476.520 2677.590 1476.580 ;
        RECT 2461.070 1476.380 2677.590 1476.520 ;
        RECT 2461.070 1476.320 2461.390 1476.380 ;
        RECT 2677.270 1476.320 2677.590 1476.380 ;
        RECT 2694.670 1476.420 2694.990 1476.480 ;
        RECT 2696.985 1476.420 2697.275 1476.465 ;
        RECT 2694.670 1476.280 2697.275 1476.420 ;
        RECT 2694.670 1476.220 2694.990 1476.280 ;
        RECT 2696.985 1476.235 2697.275 1476.280 ;
        RECT 2698.370 1474.380 2698.660 1474.425 ;
        RECT 2703.890 1474.380 2704.180 1474.425 ;
        RECT 2704.810 1474.380 2705.100 1474.425 ;
        RECT 2698.370 1474.240 2705.100 1474.380 ;
        RECT 2698.370 1474.195 2698.660 1474.240 ;
        RECT 2703.890 1474.195 2704.180 1474.240 ;
        RECT 2704.810 1474.195 2705.100 1474.240 ;
        RECT 2696.970 1473.840 2697.290 1474.100 ;
        RECT 2697.890 1473.840 2698.210 1474.100 ;
        RECT 2699.290 1474.040 2699.580 1474.085 ;
        RECT 2701.130 1474.040 2701.420 1474.085 ;
        RECT 2699.290 1473.900 2701.420 1474.040 ;
        RECT 2699.290 1473.855 2699.580 1473.900 ;
        RECT 2701.130 1473.855 2701.420 1473.900 ;
        RECT 2702.950 1473.840 2703.270 1474.100 ;
        RECT 2703.475 1474.040 2703.765 1474.085 ;
        RECT 2705.315 1474.040 2705.605 1474.085 ;
        RECT 2703.475 1473.900 2705.605 1474.040 ;
        RECT 2703.475 1473.855 2703.765 1473.900 ;
        RECT 2705.315 1473.855 2705.605 1473.900 ;
        RECT 2698.810 1473.700 2699.130 1473.760 ;
        RECT 2702.030 1473.745 2702.350 1473.760 ;
        RECT 2701.585 1473.700 2701.875 1473.745 ;
        RECT 2698.810 1473.560 2701.875 1473.700 ;
        RECT 2698.810 1473.500 2699.130 1473.560 ;
        RECT 2701.585 1473.515 2701.875 1473.560 ;
        RECT 2702.030 1473.515 2702.460 1473.745 ;
        RECT 2702.030 1473.500 2702.350 1473.515 ;
        RECT 2700.205 1473.175 2700.495 1473.405 ;
        RECT 2701.165 1473.360 2701.455 1473.405 ;
        RECT 2704.395 1473.360 2704.685 1473.405 ;
        RECT 2701.165 1473.220 2704.685 1473.360 ;
        RECT 2701.165 1473.175 2701.455 1473.220 ;
        RECT 2704.395 1473.175 2704.685 1473.220 ;
        RECT 2698.350 1473.020 2698.670 1473.080 ;
        RECT 2700.280 1473.020 2700.420 1473.175 ;
        RECT 2702.490 1473.020 2702.810 1473.080 ;
        RECT 2698.350 1472.880 2702.810 1473.020 ;
        RECT 2698.350 1472.820 2698.670 1472.880 ;
        RECT 2702.490 1472.820 2702.810 1472.880 ;
        RECT 2706.170 1472.820 2706.490 1473.080 ;
        RECT 2697.905 1472.000 2698.195 1472.045 ;
        RECT 2702.030 1472.000 2702.350 1472.060 ;
        RECT 2706.170 1472.000 2706.490 1472.060 ;
        RECT 2697.905 1471.860 2702.350 1472.000 ;
        RECT 2697.905 1471.815 2698.195 1471.860 ;
        RECT 2702.030 1471.800 2702.350 1471.860 ;
        RECT 2703.960 1471.860 2706.490 1472.000 ;
        RECT 2697.890 1471.320 2698.210 1471.380 ;
        RECT 2701.570 1471.320 2701.890 1471.380 ;
        RECT 2703.960 1471.365 2704.100 1471.860 ;
        RECT 2706.170 1471.800 2706.490 1471.860 ;
        RECT 2697.890 1471.180 2703.640 1471.320 ;
        RECT 2697.890 1471.120 2698.210 1471.180 ;
        RECT 2701.570 1471.120 2701.890 1471.180 ;
        RECT 2694.670 1470.980 2694.990 1471.040 ;
        RECT 2696.985 1470.980 2697.275 1471.025 ;
        RECT 2694.670 1470.840 2697.275 1470.980 ;
        RECT 2703.500 1470.980 2703.640 1471.180 ;
        RECT 2703.885 1471.135 2704.175 1471.365 ;
        RECT 2704.345 1471.135 2704.635 1471.365 ;
        RECT 2704.420 1470.980 2704.560 1471.135 ;
        RECT 2703.500 1470.840 2704.560 1470.980 ;
        RECT 2694.670 1470.780 2694.990 1470.840 ;
        RECT 2696.985 1470.795 2697.275 1470.840 ;
        RECT 2703.425 1470.640 2703.715 1470.685 ;
        RECT 2703.870 1470.640 2704.190 1470.700 ;
        RECT 2703.425 1470.500 2704.190 1470.640 ;
        RECT 2703.425 1470.455 2703.715 1470.500 ;
        RECT 2703.870 1470.440 2704.190 1470.500 ;
        RECT 2701.570 1470.100 2701.890 1470.360 ;
        RECT 2461.530 1469.720 2461.850 1469.780 ;
        RECT 2677.730 1469.720 2678.050 1469.780 ;
        RECT 2461.530 1469.580 2678.050 1469.720 ;
        RECT 2461.530 1469.520 2461.850 1469.580 ;
        RECT 2677.730 1469.520 2678.050 1469.580 ;
        RECT 2697.430 1466.560 2697.750 1466.620 ;
        RECT 2697.905 1466.560 2698.195 1466.605 ;
        RECT 2697.430 1466.420 2698.195 1466.560 ;
        RECT 2697.430 1466.360 2697.750 1466.420 ;
        RECT 2697.905 1466.375 2698.195 1466.420 ;
        RECT 2694.670 1465.540 2694.990 1465.600 ;
        RECT 2696.985 1465.540 2697.275 1465.585 ;
        RECT 2694.670 1465.400 2697.275 1465.540 ;
        RECT 2694.670 1465.340 2694.990 1465.400 ;
        RECT 2696.985 1465.355 2697.275 1465.400 ;
        RECT 2452.790 1462.580 2453.110 1462.640 ;
        RECT 2677.270 1462.580 2677.590 1462.640 ;
        RECT 2452.790 1462.440 2677.590 1462.580 ;
        RECT 2452.790 1462.380 2453.110 1462.440 ;
        RECT 2677.270 1462.380 2677.590 1462.440 ;
        RECT 2701.570 1459.900 2701.890 1460.160 ;
        RECT 2702.505 1460.100 2702.795 1460.145 ;
        RECT 2703.870 1460.100 2704.190 1460.160 ;
        RECT 2731.470 1460.100 2731.790 1460.160 ;
        RECT 2702.505 1459.960 2731.790 1460.100 ;
        RECT 2702.505 1459.915 2702.795 1459.960 ;
        RECT 2703.870 1459.900 2704.190 1459.960 ;
        RECT 2731.470 1459.900 2731.790 1459.960 ;
        RECT 2702.030 1459.220 2702.350 1459.480 ;
        RECT 2697.905 1458.400 2698.195 1458.445 ;
        RECT 2698.810 1458.400 2699.130 1458.460 ;
        RECT 2697.905 1458.260 2699.130 1458.400 ;
        RECT 2697.905 1458.215 2698.195 1458.260 ;
        RECT 2698.810 1458.200 2699.130 1458.260 ;
        RECT 2702.030 1458.200 2702.350 1458.460 ;
        RECT 2703.870 1458.200 2704.190 1458.460 ;
        RECT 2694.670 1457.720 2694.990 1457.780 ;
        RECT 2702.120 1457.765 2702.260 1458.200 ;
        RECT 2703.960 1457.765 2704.100 1458.200 ;
        RECT 2696.985 1457.720 2697.275 1457.765 ;
        RECT 2694.670 1457.580 2697.275 1457.720 ;
        RECT 2694.670 1457.520 2694.990 1457.580 ;
        RECT 2696.985 1457.535 2697.275 1457.580 ;
        RECT 2702.045 1457.535 2702.335 1457.765 ;
        RECT 2703.885 1457.535 2704.175 1457.765 ;
        RECT 2704.790 1457.180 2705.110 1457.440 ;
        RECT 2702.490 1456.840 2702.810 1457.100 ;
        RECT 2702.490 1455.680 2702.810 1455.740 ;
        RECT 2702.490 1455.540 2724.570 1455.680 ;
        RECT 2702.490 1455.480 2702.810 1455.540 ;
        RECT 2724.430 1454.660 2724.570 1455.540 ;
        RECT 2725.505 1454.660 2725.795 1454.705 ;
        RECT 2724.430 1454.520 2725.795 1454.660 ;
        RECT 2725.505 1454.475 2725.795 1454.520 ;
        RECT 2694.670 1452.280 2694.990 1452.340 ;
        RECT 2696.985 1452.280 2697.275 1452.325 ;
        RECT 2694.670 1452.140 2697.275 1452.280 ;
        RECT 2694.670 1452.080 2694.990 1452.140 ;
        RECT 2696.985 1452.095 2697.275 1452.140 ;
        RECT 2697.430 1451.260 2697.750 1451.320 ;
        RECT 2697.905 1451.260 2698.195 1451.305 ;
        RECT 2697.430 1451.120 2698.195 1451.260 ;
        RECT 2697.430 1451.060 2697.750 1451.120 ;
        RECT 2697.905 1451.075 2698.195 1451.120 ;
        RECT 2464.750 1449.320 2465.070 1449.380 ;
        RECT 2677.270 1449.320 2677.590 1449.380 ;
        RECT 2464.750 1449.180 2677.590 1449.320 ;
        RECT 2464.750 1449.120 2465.070 1449.180 ;
        RECT 2677.270 1449.120 2677.590 1449.180 ;
        RECT 2697.890 1446.640 2698.210 1446.900 ;
        RECT 2698.350 1446.640 2698.670 1446.900 ;
        RECT 2697.430 1446.300 2697.750 1446.560 ;
        RECT 2697.980 1446.500 2698.120 1446.640 ;
        RECT 2702.030 1446.500 2702.350 1446.560 ;
        RECT 2697.980 1446.360 2702.350 1446.500 ;
        RECT 2702.030 1446.300 2702.350 1446.360 ;
        RECT 2699.285 1445.820 2699.575 1445.865 ;
        RECT 2702.950 1445.820 2703.270 1445.880 ;
        RECT 2699.285 1445.680 2703.270 1445.820 ;
        RECT 2699.285 1445.635 2699.575 1445.680 ;
        RECT 2702.950 1445.620 2703.270 1445.680 ;
        RECT 2694.670 1443.780 2694.990 1443.840 ;
        RECT 2696.985 1443.780 2697.275 1443.825 ;
        RECT 2694.670 1443.640 2697.275 1443.780 ;
        RECT 2694.670 1443.580 2694.990 1443.640 ;
        RECT 2696.985 1443.595 2697.275 1443.640 ;
        RECT 2697.890 1442.900 2698.210 1443.160 ;
        RECT 2459.690 1442.180 2460.010 1442.240 ;
        RECT 2677.270 1442.180 2677.590 1442.240 ;
        RECT 2459.690 1442.040 2677.590 1442.180 ;
        RECT 2459.690 1441.980 2460.010 1442.040 ;
        RECT 2677.270 1441.980 2677.590 1442.040 ;
        RECT 2697.890 1442.080 2698.210 1442.140 ;
        RECT 2698.825 1442.080 2699.115 1442.125 ;
        RECT 2697.890 1441.940 2699.115 1442.080 ;
        RECT 2697.890 1441.880 2698.210 1441.940 ;
        RECT 2698.825 1441.895 2699.115 1441.940 ;
        RECT 2700.665 1442.080 2700.955 1442.125 ;
        RECT 2701.585 1442.080 2701.875 1442.125 ;
        RECT 2700.665 1441.940 2701.875 1442.080 ;
        RECT 2700.665 1441.895 2700.955 1441.940 ;
        RECT 2701.585 1441.895 2701.875 1441.940 ;
        RECT 2702.030 1441.880 2702.350 1442.140 ;
        RECT 2702.950 1441.880 2703.270 1442.140 ;
        RECT 2703.410 1441.880 2703.730 1442.140 ;
        RECT 2698.350 1441.740 2698.670 1441.800 ;
        RECT 2697.980 1441.600 2698.670 1441.740 ;
        RECT 2697.980 1441.105 2698.120 1441.600 ;
        RECT 2698.350 1441.540 2698.670 1441.600 ;
        RECT 2702.120 1441.445 2702.260 1441.880 ;
        RECT 2702.045 1441.215 2702.335 1441.445 ;
        RECT 2702.490 1441.200 2702.810 1441.460 ;
        RECT 2703.040 1441.445 2703.180 1441.880 ;
        RECT 2702.965 1441.215 2703.255 1441.445 ;
        RECT 2697.905 1440.875 2698.195 1441.105 ;
        RECT 2698.350 1440.860 2698.670 1441.120 ;
        RECT 2702.580 1441.060 2702.720 1441.200 ;
        RECT 2703.425 1441.060 2703.715 1441.105 ;
        RECT 2702.580 1440.920 2703.715 1441.060 ;
        RECT 2703.425 1440.875 2703.715 1440.920 ;
        RECT 2702.490 1440.180 2702.810 1440.440 ;
        RECT 2698.810 1439.160 2699.130 1439.420 ;
        RECT 2699.745 1439.360 2700.035 1439.405 ;
        RECT 2702.490 1439.360 2702.810 1439.420 ;
        RECT 2699.745 1439.220 2702.810 1439.360 ;
        RECT 2699.745 1439.175 2700.035 1439.220 ;
        RECT 2702.490 1439.160 2702.810 1439.220 ;
        RECT 2696.985 1439.020 2697.275 1439.065 ;
        RECT 2697.430 1439.020 2697.750 1439.080 ;
        RECT 2696.985 1438.880 2697.750 1439.020 ;
        RECT 2698.900 1439.020 2699.040 1439.160 ;
        RECT 2702.030 1439.020 2702.350 1439.080 ;
        RECT 2698.900 1438.880 2702.350 1439.020 ;
        RECT 2696.985 1438.835 2697.275 1438.880 ;
        RECT 2697.430 1438.820 2697.750 1438.880 ;
        RECT 2702.030 1438.820 2702.350 1438.880 ;
        RECT 2523.545 1437.360 2523.865 1437.620 ;
        RECT 2698.810 1437.460 2699.130 1437.720 ;
        RECT 2697.905 1436.640 2698.195 1436.685 ;
        RECT 2698.810 1436.640 2699.130 1436.700 ;
        RECT 2697.905 1436.500 2699.130 1436.640 ;
        RECT 2697.905 1436.455 2698.195 1436.500 ;
        RECT 2698.810 1436.440 2699.130 1436.500 ;
        RECT 2694.670 1435.960 2694.990 1436.020 ;
        RECT 2696.985 1435.960 2697.275 1436.005 ;
        RECT 2694.670 1435.820 2697.275 1435.960 ;
        RECT 2694.670 1435.760 2694.990 1435.820 ;
        RECT 2696.985 1435.775 2697.275 1435.820 ;
        RECT 2359.540 1435.060 2359.830 1435.290 ;
        RECT 2370.355 1435.060 2370.645 1435.290 ;
        RECT 2375.970 1435.060 2376.260 1435.290 ;
        RECT 2359.600 1434.610 2359.770 1435.060 ;
        RECT 2370.415 1434.715 2370.585 1435.060 ;
        RECT 2359.510 1434.320 2359.860 1434.610 ;
        RECT 2370.315 1434.345 2370.695 1434.715 ;
        RECT 2376.030 1434.580 2376.200 1435.060 ;
        RECT 2377.760 1435.030 2378.055 1435.290 ;
        RECT 2377.390 1434.635 2377.620 1434.660 ;
        RECT 2377.360 1434.580 2377.650 1434.635 ;
        RECT 2376.030 1434.550 2377.650 1434.580 ;
        RECT 2375.970 1434.410 2377.650 1434.550 ;
        RECT 2370.355 1434.320 2370.645 1434.345 ;
        RECT 2375.970 1434.320 2376.260 1434.410 ;
        RECT 2377.360 1434.335 2377.650 1434.410 ;
        RECT 2377.390 1434.310 2377.620 1434.335 ;
        RECT 2370.990 1434.180 2371.340 1434.245 ;
        RECT 2376.425 1434.180 2376.750 1434.270 ;
        RECT 2370.785 1434.150 2371.340 1434.180 ;
        RECT 2376.400 1434.150 2376.750 1434.180 ;
        RECT 2370.615 1434.145 2371.340 1434.150 ;
        RECT 2376.230 1434.145 2376.750 1434.150 ;
        RECT 2370.615 1433.975 2376.750 1434.145 ;
        RECT 2370.785 1433.950 2371.340 1433.975 ;
        RECT 2376.400 1433.950 2376.750 1433.975 ;
        RECT 2370.990 1433.895 2371.340 1433.950 ;
        RECT 2376.425 1433.945 2376.750 1433.950 ;
        RECT 2377.820 1433.930 2377.990 1435.030 ;
        RECT 2378.755 1435.025 2379.050 1435.285 ;
        RECT 2388.915 1435.060 2389.205 1435.290 ;
        RECT 2394.530 1435.060 2394.820 1435.290 ;
        RECT 2378.815 1434.295 2378.985 1435.025 ;
        RECT 2388.975 1434.715 2389.145 1435.060 ;
        RECT 2388.875 1434.345 2389.255 1434.715 ;
        RECT 2394.590 1434.580 2394.760 1435.060 ;
        RECT 2396.320 1435.030 2396.615 1435.290 ;
        RECT 2395.950 1434.635 2396.180 1434.660 ;
        RECT 2395.920 1434.580 2396.210 1434.635 ;
        RECT 2394.590 1434.550 2396.210 1434.580 ;
        RECT 2394.530 1434.410 2396.210 1434.550 ;
        RECT 2388.915 1434.320 2389.205 1434.345 ;
        RECT 2394.530 1434.320 2394.820 1434.410 ;
        RECT 2395.920 1434.335 2396.210 1434.410 ;
        RECT 2395.950 1434.310 2396.180 1434.335 ;
        RECT 2377.760 1433.925 2377.990 1433.930 ;
        RECT 2378.805 1433.945 2379.155 1434.295 ;
        RECT 2389.550 1434.180 2389.900 1434.250 ;
        RECT 2394.985 1434.180 2395.310 1434.270 ;
        RECT 2389.345 1434.150 2389.900 1434.180 ;
        RECT 2394.960 1434.150 2395.310 1434.180 ;
        RECT 2389.175 1434.145 2389.900 1434.150 ;
        RECT 2394.790 1434.145 2395.310 1434.150 ;
        RECT 2389.175 1433.975 2395.310 1434.145 ;
        RECT 2389.345 1433.950 2389.900 1433.975 ;
        RECT 2394.960 1433.950 2395.310 1433.975 ;
        RECT 2378.805 1433.925 2379.105 1433.945 ;
        RECT 2359.135 1433.790 2359.485 1433.865 ;
        RECT 2375.625 1433.820 2375.945 1433.835 ;
        RECT 2375.600 1433.790 2375.945 1433.820 ;
        RECT 2358.995 1433.620 2359.485 1433.790 ;
        RECT 2375.425 1433.620 2375.945 1433.790 ;
        RECT 2377.760 1433.690 2378.050 1433.925 ;
        RECT 2378.755 1433.855 2379.105 1433.925 ;
        RECT 2389.550 1433.900 2389.900 1433.950 ;
        RECT 2394.985 1433.945 2395.310 1433.950 ;
        RECT 2396.380 1433.930 2396.550 1435.030 ;
        RECT 2397.315 1435.025 2397.610 1435.285 ;
        RECT 2407.475 1435.060 2407.765 1435.290 ;
        RECT 2413.090 1435.060 2413.380 1435.290 ;
        RECT 2397.375 1434.305 2397.545 1435.025 ;
        RECT 2407.535 1434.715 2407.705 1435.060 ;
        RECT 2407.435 1434.345 2407.815 1434.715 ;
        RECT 2413.150 1434.580 2413.320 1435.060 ;
        RECT 2414.880 1435.030 2415.175 1435.290 ;
        RECT 2414.510 1434.635 2414.740 1434.660 ;
        RECT 2414.480 1434.580 2414.770 1434.635 ;
        RECT 2413.150 1434.550 2414.770 1434.580 ;
        RECT 2413.090 1434.410 2414.770 1434.550 ;
        RECT 2407.475 1434.320 2407.765 1434.345 ;
        RECT 2413.090 1434.320 2413.380 1434.410 ;
        RECT 2414.480 1434.335 2414.770 1434.410 ;
        RECT 2414.510 1434.310 2414.740 1434.335 ;
        RECT 2396.320 1433.925 2396.550 1433.930 ;
        RECT 2397.360 1433.950 2397.715 1434.305 ;
        RECT 2408.105 1434.180 2408.455 1434.255 ;
        RECT 2413.545 1434.180 2413.870 1434.270 ;
        RECT 2407.905 1434.150 2408.455 1434.180 ;
        RECT 2413.520 1434.150 2413.870 1434.180 ;
        RECT 2407.735 1434.145 2408.455 1434.150 ;
        RECT 2413.350 1434.145 2413.870 1434.150 ;
        RECT 2407.735 1433.975 2413.870 1434.145 ;
        RECT 2407.905 1433.950 2408.455 1433.975 ;
        RECT 2413.520 1433.950 2413.870 1433.975 ;
        RECT 2397.360 1433.925 2397.665 1433.950 ;
        RECT 2378.755 1433.685 2379.045 1433.855 ;
        RECT 2394.185 1433.820 2394.505 1433.835 ;
        RECT 2394.160 1433.790 2394.505 1433.820 ;
        RECT 2393.985 1433.620 2394.505 1433.790 ;
        RECT 2396.320 1433.690 2396.610 1433.925 ;
        RECT 2397.315 1433.850 2397.665 1433.925 ;
        RECT 2408.105 1433.905 2408.455 1433.950 ;
        RECT 2413.545 1433.945 2413.870 1433.950 ;
        RECT 2414.940 1433.930 2415.110 1435.030 ;
        RECT 2415.875 1435.025 2416.170 1435.285 ;
        RECT 2426.035 1435.060 2426.325 1435.290 ;
        RECT 2431.650 1435.060 2431.940 1435.290 ;
        RECT 2415.935 1434.295 2416.105 1435.025 ;
        RECT 2426.095 1434.715 2426.265 1435.060 ;
        RECT 2425.995 1434.345 2426.375 1434.715 ;
        RECT 2431.710 1434.580 2431.880 1435.060 ;
        RECT 2433.440 1435.030 2433.735 1435.290 ;
        RECT 2433.070 1434.635 2433.300 1434.660 ;
        RECT 2433.040 1434.580 2433.330 1434.635 ;
        RECT 2431.710 1434.550 2433.330 1434.580 ;
        RECT 2431.650 1434.410 2433.330 1434.550 ;
        RECT 2426.035 1434.320 2426.325 1434.345 ;
        RECT 2431.650 1434.320 2431.940 1434.410 ;
        RECT 2433.040 1434.335 2433.330 1434.410 ;
        RECT 2433.070 1434.310 2433.300 1434.335 ;
        RECT 2414.880 1433.925 2415.110 1433.930 ;
        RECT 2415.880 1433.945 2416.230 1434.295 ;
        RECT 2426.665 1434.180 2427.015 1434.250 ;
        RECT 2432.105 1434.180 2432.430 1434.270 ;
        RECT 2426.465 1434.150 2427.015 1434.180 ;
        RECT 2432.080 1434.150 2432.430 1434.180 ;
        RECT 2426.295 1434.145 2427.015 1434.150 ;
        RECT 2431.910 1434.145 2432.430 1434.150 ;
        RECT 2426.295 1433.975 2432.430 1434.145 ;
        RECT 2426.465 1433.950 2427.015 1433.975 ;
        RECT 2432.080 1433.950 2432.430 1433.975 ;
        RECT 2415.880 1433.925 2416.225 1433.945 ;
        RECT 2397.315 1433.685 2397.605 1433.850 ;
        RECT 2412.745 1433.820 2413.065 1433.835 ;
        RECT 2412.720 1433.790 2413.065 1433.820 ;
        RECT 2412.545 1433.620 2413.065 1433.790 ;
        RECT 2414.880 1433.690 2415.170 1433.925 ;
        RECT 2415.875 1433.855 2416.225 1433.925 ;
        RECT 2426.665 1433.900 2427.015 1433.950 ;
        RECT 2432.105 1433.945 2432.430 1433.950 ;
        RECT 2433.500 1433.930 2433.670 1435.030 ;
        RECT 2434.435 1435.025 2434.730 1435.285 ;
        RECT 2444.595 1435.060 2444.885 1435.290 ;
        RECT 2450.210 1435.060 2450.500 1435.290 ;
        RECT 2434.495 1434.295 2434.665 1435.025 ;
        RECT 2444.655 1434.715 2444.825 1435.060 ;
        RECT 2444.555 1434.345 2444.935 1434.715 ;
        RECT 2450.270 1434.580 2450.440 1435.060 ;
        RECT 2452.000 1435.030 2452.295 1435.290 ;
        RECT 2451.630 1434.635 2451.860 1434.660 ;
        RECT 2451.600 1434.580 2451.890 1434.635 ;
        RECT 2450.270 1434.550 2451.890 1434.580 ;
        RECT 2450.210 1434.410 2451.890 1434.550 ;
        RECT 2444.595 1434.320 2444.885 1434.345 ;
        RECT 2450.210 1434.320 2450.500 1434.410 ;
        RECT 2451.600 1434.335 2451.890 1434.410 ;
        RECT 2451.630 1434.310 2451.860 1434.335 ;
        RECT 2433.440 1433.925 2433.670 1433.930 ;
        RECT 2434.440 1433.945 2434.790 1434.295 ;
        RECT 2445.225 1434.180 2445.575 1434.250 ;
        RECT 2450.665 1434.180 2450.990 1434.270 ;
        RECT 2445.025 1434.150 2445.575 1434.180 ;
        RECT 2450.640 1434.150 2450.990 1434.180 ;
        RECT 2444.855 1434.145 2445.575 1434.150 ;
        RECT 2450.470 1434.145 2450.990 1434.150 ;
        RECT 2444.855 1433.975 2450.990 1434.145 ;
        RECT 2445.025 1433.950 2445.575 1433.975 ;
        RECT 2450.640 1433.950 2450.990 1433.975 ;
        RECT 2434.440 1433.925 2434.785 1433.945 ;
        RECT 2415.875 1433.685 2416.165 1433.855 ;
        RECT 2431.305 1433.820 2431.625 1433.835 ;
        RECT 2431.280 1433.790 2431.625 1433.820 ;
        RECT 2431.105 1433.620 2431.625 1433.790 ;
        RECT 2433.440 1433.690 2433.730 1433.925 ;
        RECT 2434.435 1433.855 2434.785 1433.925 ;
        RECT 2445.225 1433.900 2445.575 1433.950 ;
        RECT 2450.665 1433.945 2450.990 1433.950 ;
        RECT 2452.060 1433.930 2452.230 1435.030 ;
        RECT 2452.995 1435.025 2453.290 1435.285 ;
        RECT 2453.025 1435.000 2453.290 1435.025 ;
        RECT 2453.025 1434.915 2453.350 1435.000 ;
        RECT 2453.025 1434.565 2453.375 1434.915 ;
        RECT 2452.000 1433.925 2452.230 1433.930 ;
        RECT 2453.055 1433.925 2453.225 1434.565 ;
        RECT 2434.435 1433.685 2434.725 1433.855 ;
        RECT 2449.865 1433.820 2450.185 1433.835 ;
        RECT 2449.840 1433.790 2450.185 1433.820 ;
        RECT 2449.665 1433.620 2450.185 1433.790 ;
        RECT 2452.000 1433.690 2452.290 1433.925 ;
        RECT 2452.995 1433.920 2453.225 1433.925 ;
        RECT 2452.995 1433.685 2453.285 1433.920 ;
        RECT 2359.135 1433.575 2359.485 1433.620 ;
        RECT 2375.600 1433.590 2375.945 1433.620 ;
        RECT 2394.160 1433.590 2394.505 1433.620 ;
        RECT 2412.720 1433.590 2413.065 1433.620 ;
        RECT 2431.280 1433.590 2431.625 1433.620 ;
        RECT 2449.840 1433.590 2450.185 1433.620 ;
        RECT 2375.625 1433.545 2375.945 1433.590 ;
        RECT 2394.185 1433.545 2394.505 1433.590 ;
        RECT 2412.745 1433.545 2413.065 1433.590 ;
        RECT 2431.305 1433.545 2431.625 1433.590 ;
        RECT 2449.865 1433.545 2450.185 1433.590 ;
        RECT 2700.205 1433.240 2700.495 1433.285 ;
        RECT 2701.570 1433.240 2701.890 1433.300 ;
        RECT 2700.205 1433.100 2701.890 1433.240 ;
        RECT 2700.205 1433.055 2700.495 1433.100 ;
        RECT 2701.570 1433.040 2701.890 1433.100 ;
        RECT 2698.365 1432.900 2698.655 1432.945 ;
        RECT 2699.730 1432.900 2700.050 1432.960 ;
        RECT 2698.365 1432.760 2700.050 1432.900 ;
        RECT 2698.365 1432.715 2698.655 1432.760 ;
        RECT 2699.730 1432.700 2700.050 1432.760 ;
        RECT 2700.665 1432.900 2700.955 1432.945 ;
        RECT 2703.410 1432.900 2703.730 1432.960 ;
        RECT 2700.665 1432.760 2703.730 1432.900 ;
        RECT 2700.665 1432.715 2700.955 1432.760 ;
        RECT 2703.410 1432.700 2703.730 1432.760 ;
        RECT 2696.970 1432.560 2697.290 1432.620 ;
        RECT 2702.030 1432.560 2702.350 1432.620 ;
        RECT 2696.970 1432.420 2702.350 1432.560 ;
        RECT 2696.970 1432.360 2697.290 1432.420 ;
        RECT 2702.030 1432.360 2702.350 1432.420 ;
        RECT 2698.810 1432.020 2699.130 1432.280 ;
        RECT 2699.270 1432.020 2699.590 1432.280 ;
        RECT 2701.585 1432.220 2701.875 1432.265 ;
        RECT 2703.870 1432.220 2704.190 1432.280 ;
        RECT 2701.585 1432.080 2704.190 1432.220 ;
        RECT 2701.585 1432.035 2701.875 1432.080 ;
        RECT 2703.870 1432.020 2704.190 1432.080 ;
        RECT 2523.545 1430.945 2523.865 1431.205 ;
        RECT 2698.810 1431.200 2699.130 1431.260 ;
        RECT 2701.125 1431.200 2701.415 1431.245 ;
        RECT 2698.810 1431.060 2701.415 1431.200 ;
        RECT 2698.810 1431.000 2699.130 1431.060 ;
        RECT 2701.125 1431.015 2701.415 1431.060 ;
        RECT 2699.730 1430.860 2700.050 1430.920 ;
        RECT 2697.520 1430.720 2699.500 1430.860 ;
        RECT 2697.520 1430.580 2697.660 1430.720 ;
        RECT 2697.430 1430.320 2697.750 1430.580 ;
        RECT 2697.890 1430.320 2698.210 1430.580 ;
        RECT 2699.360 1430.225 2699.500 1430.720 ;
        RECT 2699.730 1430.720 2700.880 1430.860 ;
        RECT 2699.730 1430.660 2700.050 1430.720 ;
        RECT 2366.550 1430.065 2366.870 1430.125 ;
        RECT 2361.790 1429.555 2362.110 1429.965 ;
        RECT 2366.550 1429.925 2367.620 1430.065 ;
        RECT 2364.800 1429.825 2365.900 1429.895 ;
        RECT 2366.550 1429.865 2366.870 1429.925 ;
        RECT 2364.730 1429.755 2365.980 1429.825 ;
        RECT 2364.730 1429.595 2365.020 1429.755 ;
        RECT 2365.690 1429.595 2365.980 1429.755 ;
        RECT 2361.870 1428.425 2362.030 1429.555 ;
        RECT 2362.750 1429.305 2363.070 1429.565 ;
        RECT 2363.870 1429.445 2364.190 1429.565 ;
        RECT 2365.210 1429.505 2365.500 1429.545 ;
        RECT 2363.870 1429.305 2364.700 1429.445 ;
        RECT 2365.210 1429.315 2365.540 1429.505 ;
        RECT 2364.490 1429.265 2364.700 1429.305 ;
        RECT 2364.490 1429.035 2364.780 1429.265 ;
        RECT 2362.270 1428.985 2362.590 1429.005 ;
        RECT 2362.270 1428.845 2363.220 1428.985 ;
        RECT 2363.680 1428.945 2363.970 1428.985 ;
        RECT 2362.270 1428.755 2362.820 1428.845 ;
        RECT 2363.080 1428.805 2363.220 1428.845 ;
        RECT 2363.580 1428.805 2363.970 1428.945 ;
        RECT 2363.080 1428.755 2363.970 1428.805 ;
        RECT 2362.270 1428.745 2362.590 1428.755 ;
        RECT 2363.080 1428.665 2363.720 1428.755 ;
        RECT 2361.810 1428.195 2362.100 1428.425 ;
        RECT 2362.750 1428.385 2363.070 1428.445 ;
        RECT 2364.710 1428.385 2365.030 1428.445 ;
        RECT 2365.400 1428.425 2365.540 1429.315 ;
        RECT 2366.190 1429.305 2366.510 1429.565 ;
        RECT 2366.910 1429.305 2367.230 1429.565 ;
        RECT 2367.480 1429.505 2367.620 1429.925 ;
        RECT 2368.110 1429.865 2368.430 1430.125 ;
        RECT 2368.650 1430.065 2368.940 1430.105 ;
        RECT 2369.110 1430.065 2369.430 1430.125 ;
        RECT 2368.650 1429.925 2369.430 1430.065 ;
        RECT 2368.650 1429.875 2368.940 1429.925 ;
        RECT 2369.110 1429.865 2369.430 1429.925 ;
        RECT 2369.590 1429.865 2369.910 1430.125 ;
        RECT 2370.070 1429.865 2370.390 1430.125 ;
        RECT 2371.070 1429.895 2371.390 1430.125 ;
        RECT 2385.110 1430.065 2385.430 1430.125 ;
        RECT 2371.070 1429.865 2372.500 1429.895 ;
        RECT 2371.160 1429.755 2372.500 1429.865 ;
        RECT 2368.650 1429.505 2368.940 1429.545 ;
        RECT 2367.480 1429.365 2368.940 1429.505 ;
        RECT 2368.650 1429.315 2368.940 1429.365 ;
        RECT 2370.590 1429.305 2370.910 1429.565 ;
        RECT 2371.160 1429.545 2371.300 1429.755 ;
        RECT 2371.090 1429.315 2371.380 1429.545 ;
        RECT 2371.810 1429.505 2372.100 1429.545 ;
        RECT 2371.810 1429.315 2372.140 1429.505 ;
        RECT 2370.090 1429.225 2370.380 1429.265 ;
        RECT 2370.590 1429.225 2370.820 1429.305 ;
        RECT 2370.090 1429.085 2370.820 1429.225 ;
        RECT 2370.090 1429.035 2370.380 1429.085 ;
        RECT 2365.930 1428.985 2366.250 1429.005 ;
        RECT 2365.690 1428.945 2366.250 1428.985 ;
        RECT 2366.930 1428.945 2367.220 1428.985 ;
        RECT 2365.690 1428.805 2367.220 1428.945 ;
        RECT 2365.690 1428.755 2366.250 1428.805 ;
        RECT 2366.930 1428.755 2367.220 1428.805 ;
        RECT 2367.410 1428.945 2367.700 1428.985 ;
        RECT 2367.410 1428.805 2368.340 1428.945 ;
        RECT 2367.410 1428.755 2367.700 1428.805 ;
        RECT 2365.930 1428.745 2366.250 1428.755 ;
        RECT 2362.750 1428.245 2365.030 1428.385 ;
        RECT 2362.750 1428.185 2363.070 1428.245 ;
        RECT 2364.710 1428.185 2365.030 1428.245 ;
        RECT 2365.210 1428.385 2365.540 1428.425 ;
        RECT 2366.190 1428.385 2366.510 1428.445 ;
        RECT 2366.910 1428.425 2367.230 1428.445 ;
        RECT 2365.210 1428.245 2366.510 1428.385 ;
        RECT 2365.210 1428.195 2365.500 1428.245 ;
        RECT 2366.190 1428.185 2366.510 1428.245 ;
        RECT 2366.690 1428.195 2367.230 1428.425 ;
        RECT 2366.910 1428.185 2367.230 1428.195 ;
        RECT 2367.630 1428.185 2367.950 1428.445 ;
        RECT 2368.200 1428.385 2368.340 1428.805 ;
        RECT 2368.630 1428.805 2368.950 1429.005 ;
        RECT 2371.330 1428.805 2371.620 1428.985 ;
        RECT 2368.630 1428.755 2371.620 1428.805 ;
        RECT 2368.630 1428.745 2371.540 1428.755 ;
        RECT 2368.720 1428.665 2371.540 1428.745 ;
        RECT 2372.000 1428.445 2372.140 1429.315 ;
        RECT 2372.360 1429.265 2372.500 1429.755 ;
        RECT 2374.020 1429.445 2374.360 1429.795 ;
        RECT 2380.350 1429.555 2380.670 1429.965 ;
        RECT 2385.110 1429.925 2386.180 1430.065 ;
        RECT 2383.360 1429.825 2384.460 1429.895 ;
        RECT 2385.110 1429.865 2385.430 1429.925 ;
        RECT 2383.290 1429.755 2384.540 1429.825 ;
        RECT 2383.290 1429.595 2383.580 1429.755 ;
        RECT 2384.250 1429.595 2384.540 1429.755 ;
        RECT 2372.290 1429.035 2372.580 1429.265 ;
        RECT 2374.110 1428.490 2374.280 1429.445 ;
        RECT 2375.625 1428.875 2375.945 1428.980 ;
        RECT 2375.600 1428.860 2375.945 1428.875 ;
        RECT 2375.595 1428.845 2375.945 1428.860 ;
        RECT 2375.425 1428.675 2375.945 1428.845 ;
        RECT 2375.600 1428.660 2375.945 1428.675 ;
        RECT 2375.600 1428.645 2375.890 1428.660 ;
        RECT 2376.400 1428.490 2376.750 1428.610 ;
        RECT 2377.760 1428.540 2378.050 1428.775 ;
        RECT 2378.750 1428.545 2379.040 1428.780 ;
        RECT 2378.750 1428.540 2378.980 1428.545 ;
        RECT 2377.760 1428.535 2377.990 1428.540 ;
        RECT 2368.870 1428.425 2369.190 1428.445 ;
        RECT 2368.650 1428.385 2369.190 1428.425 ;
        RECT 2368.200 1428.245 2369.190 1428.385 ;
        RECT 2368.650 1428.195 2369.190 1428.245 ;
        RECT 2368.870 1428.185 2369.190 1428.195 ;
        RECT 2369.470 1428.185 2370.150 1428.445 ;
        RECT 2370.590 1428.385 2370.910 1428.445 ;
        RECT 2371.090 1428.385 2371.380 1428.425 ;
        RECT 2370.590 1428.245 2371.380 1428.385 ;
        RECT 2372.000 1428.245 2372.350 1428.445 ;
        RECT 2374.110 1428.320 2376.750 1428.490 ;
        RECT 2376.230 1428.315 2376.750 1428.320 ;
        RECT 2376.400 1428.260 2376.750 1428.315 ;
        RECT 2370.590 1428.185 2370.910 1428.245 ;
        RECT 2371.090 1428.195 2371.380 1428.245 ;
        RECT 2372.030 1428.185 2372.350 1428.245 ;
        RECT 2377.390 1428.220 2377.620 1428.235 ;
        RECT 2375.970 1428.120 2376.260 1428.145 ;
        RECT 2377.360 1428.120 2377.655 1428.220 ;
        RECT 2375.970 1427.950 2377.655 1428.120 ;
        RECT 2375.970 1427.915 2376.260 1427.950 ;
        RECT 2376.030 1427.405 2376.200 1427.915 ;
        RECT 2377.360 1427.900 2377.655 1427.950 ;
        RECT 2377.390 1427.885 2377.620 1427.900 ;
        RECT 2377.820 1427.435 2377.990 1428.535 ;
        RECT 2378.810 1427.440 2378.980 1428.540 ;
        RECT 2380.430 1428.425 2380.590 1429.555 ;
        RECT 2381.310 1429.305 2381.630 1429.565 ;
        RECT 2382.430 1429.445 2382.750 1429.565 ;
        RECT 2383.770 1429.505 2384.060 1429.545 ;
        RECT 2382.430 1429.305 2383.260 1429.445 ;
        RECT 2383.770 1429.315 2384.100 1429.505 ;
        RECT 2383.050 1429.265 2383.260 1429.305 ;
        RECT 2383.050 1429.035 2383.340 1429.265 ;
        RECT 2380.830 1428.985 2381.150 1429.005 ;
        RECT 2380.830 1428.845 2381.780 1428.985 ;
        RECT 2382.240 1428.945 2382.530 1428.985 ;
        RECT 2380.830 1428.755 2381.380 1428.845 ;
        RECT 2381.640 1428.805 2381.780 1428.845 ;
        RECT 2382.140 1428.805 2382.530 1428.945 ;
        RECT 2381.640 1428.755 2382.530 1428.805 ;
        RECT 2380.830 1428.745 2381.150 1428.755 ;
        RECT 2381.640 1428.665 2382.280 1428.755 ;
        RECT 2380.370 1428.195 2380.660 1428.425 ;
        RECT 2381.310 1428.385 2381.630 1428.445 ;
        RECT 2383.270 1428.385 2383.590 1428.445 ;
        RECT 2383.960 1428.425 2384.100 1429.315 ;
        RECT 2384.750 1429.305 2385.070 1429.565 ;
        RECT 2385.470 1429.305 2385.790 1429.565 ;
        RECT 2386.040 1429.505 2386.180 1429.925 ;
        RECT 2386.670 1429.865 2386.990 1430.125 ;
        RECT 2387.210 1430.065 2387.500 1430.105 ;
        RECT 2387.670 1430.065 2387.990 1430.125 ;
        RECT 2387.210 1429.925 2387.990 1430.065 ;
        RECT 2387.210 1429.875 2387.500 1429.925 ;
        RECT 2387.670 1429.865 2387.990 1429.925 ;
        RECT 2388.150 1429.865 2388.470 1430.125 ;
        RECT 2388.630 1429.865 2388.950 1430.125 ;
        RECT 2389.630 1429.895 2389.950 1430.125 ;
        RECT 2403.670 1430.065 2403.990 1430.125 ;
        RECT 2389.630 1429.865 2391.060 1429.895 ;
        RECT 2389.720 1429.755 2391.060 1429.865 ;
        RECT 2387.210 1429.505 2387.500 1429.545 ;
        RECT 2386.040 1429.365 2387.500 1429.505 ;
        RECT 2387.210 1429.315 2387.500 1429.365 ;
        RECT 2389.150 1429.305 2389.470 1429.565 ;
        RECT 2389.720 1429.545 2389.860 1429.755 ;
        RECT 2389.650 1429.315 2389.940 1429.545 ;
        RECT 2390.370 1429.505 2390.660 1429.545 ;
        RECT 2390.370 1429.315 2390.700 1429.505 ;
        RECT 2388.650 1429.225 2388.940 1429.265 ;
        RECT 2389.150 1429.225 2389.380 1429.305 ;
        RECT 2388.650 1429.085 2389.380 1429.225 ;
        RECT 2388.650 1429.035 2388.940 1429.085 ;
        RECT 2384.490 1428.985 2384.810 1429.005 ;
        RECT 2384.250 1428.945 2384.810 1428.985 ;
        RECT 2385.490 1428.945 2385.780 1428.985 ;
        RECT 2384.250 1428.805 2385.780 1428.945 ;
        RECT 2384.250 1428.755 2384.810 1428.805 ;
        RECT 2385.490 1428.755 2385.780 1428.805 ;
        RECT 2385.970 1428.945 2386.260 1428.985 ;
        RECT 2385.970 1428.805 2386.900 1428.945 ;
        RECT 2385.970 1428.755 2386.260 1428.805 ;
        RECT 2384.490 1428.745 2384.810 1428.755 ;
        RECT 2381.310 1428.245 2383.590 1428.385 ;
        RECT 2381.310 1428.185 2381.630 1428.245 ;
        RECT 2383.270 1428.185 2383.590 1428.245 ;
        RECT 2383.770 1428.385 2384.100 1428.425 ;
        RECT 2384.750 1428.385 2385.070 1428.445 ;
        RECT 2385.470 1428.425 2385.790 1428.445 ;
        RECT 2383.770 1428.245 2385.070 1428.385 ;
        RECT 2383.770 1428.195 2384.060 1428.245 ;
        RECT 2384.750 1428.185 2385.070 1428.245 ;
        RECT 2385.250 1428.195 2385.790 1428.425 ;
        RECT 2385.470 1428.185 2385.790 1428.195 ;
        RECT 2386.190 1428.185 2386.510 1428.445 ;
        RECT 2386.760 1428.385 2386.900 1428.805 ;
        RECT 2387.190 1428.805 2387.510 1429.005 ;
        RECT 2389.890 1428.805 2390.180 1428.985 ;
        RECT 2387.190 1428.755 2390.180 1428.805 ;
        RECT 2387.190 1428.745 2390.100 1428.755 ;
        RECT 2387.280 1428.665 2390.100 1428.745 ;
        RECT 2390.560 1428.445 2390.700 1429.315 ;
        RECT 2390.920 1429.265 2391.060 1429.755 ;
        RECT 2392.580 1429.445 2392.920 1429.795 ;
        RECT 2398.910 1429.555 2399.230 1429.965 ;
        RECT 2403.670 1429.925 2404.740 1430.065 ;
        RECT 2401.920 1429.825 2403.020 1429.895 ;
        RECT 2403.670 1429.865 2403.990 1429.925 ;
        RECT 2401.850 1429.755 2403.100 1429.825 ;
        RECT 2401.850 1429.595 2402.140 1429.755 ;
        RECT 2402.810 1429.595 2403.100 1429.755 ;
        RECT 2390.850 1429.035 2391.140 1429.265 ;
        RECT 2392.670 1428.490 2392.840 1429.445 ;
        RECT 2397.130 1429.305 2397.450 1429.320 ;
        RECT 2397.130 1429.075 2397.600 1429.305 ;
        RECT 2397.130 1429.060 2397.450 1429.075 ;
        RECT 2394.185 1428.875 2394.505 1428.980 ;
        RECT 2394.160 1428.860 2394.505 1428.875 ;
        RECT 2394.155 1428.845 2394.505 1428.860 ;
        RECT 2393.985 1428.675 2394.505 1428.845 ;
        RECT 2394.160 1428.660 2394.505 1428.675 ;
        RECT 2394.160 1428.645 2394.450 1428.660 ;
        RECT 2394.960 1428.490 2395.310 1428.610 ;
        RECT 2396.320 1428.540 2396.610 1428.775 ;
        RECT 2397.310 1428.545 2397.600 1428.780 ;
        RECT 2397.310 1428.540 2397.540 1428.545 ;
        RECT 2396.320 1428.535 2396.550 1428.540 ;
        RECT 2387.430 1428.425 2387.750 1428.445 ;
        RECT 2387.210 1428.385 2387.750 1428.425 ;
        RECT 2386.760 1428.245 2387.750 1428.385 ;
        RECT 2387.210 1428.195 2387.750 1428.245 ;
        RECT 2387.430 1428.185 2387.750 1428.195 ;
        RECT 2388.030 1428.185 2388.710 1428.445 ;
        RECT 2389.150 1428.385 2389.470 1428.445 ;
        RECT 2389.650 1428.385 2389.940 1428.425 ;
        RECT 2389.150 1428.245 2389.940 1428.385 ;
        RECT 2390.560 1428.245 2390.910 1428.445 ;
        RECT 2392.670 1428.320 2395.310 1428.490 ;
        RECT 2394.790 1428.315 2395.310 1428.320 ;
        RECT 2394.960 1428.260 2395.310 1428.315 ;
        RECT 2389.150 1428.185 2389.470 1428.245 ;
        RECT 2389.650 1428.195 2389.940 1428.245 ;
        RECT 2390.590 1428.185 2390.910 1428.245 ;
        RECT 2395.950 1428.220 2396.180 1428.235 ;
        RECT 2394.530 1428.120 2394.820 1428.145 ;
        RECT 2395.920 1428.120 2396.215 1428.220 ;
        RECT 2394.530 1427.950 2396.215 1428.120 ;
        RECT 2394.530 1427.915 2394.820 1427.950 ;
        RECT 2375.970 1427.175 2376.260 1427.405 ;
        RECT 2377.760 1427.175 2378.055 1427.435 ;
        RECT 2378.730 1427.180 2379.050 1427.440 ;
        RECT 2394.590 1427.405 2394.760 1427.915 ;
        RECT 2395.920 1427.900 2396.215 1427.950 ;
        RECT 2395.950 1427.885 2396.180 1427.900 ;
        RECT 2396.380 1427.435 2396.550 1428.535 ;
        RECT 2397.370 1427.440 2397.540 1428.540 ;
        RECT 2398.990 1428.425 2399.150 1429.555 ;
        RECT 2399.870 1429.305 2400.190 1429.565 ;
        RECT 2400.990 1429.445 2401.310 1429.565 ;
        RECT 2402.330 1429.505 2402.620 1429.545 ;
        RECT 2400.990 1429.305 2401.820 1429.445 ;
        RECT 2402.330 1429.315 2402.660 1429.505 ;
        RECT 2401.610 1429.265 2401.820 1429.305 ;
        RECT 2401.610 1429.035 2401.900 1429.265 ;
        RECT 2399.390 1428.985 2399.710 1429.005 ;
        RECT 2399.390 1428.845 2400.340 1428.985 ;
        RECT 2400.800 1428.945 2401.090 1428.985 ;
        RECT 2399.390 1428.755 2399.940 1428.845 ;
        RECT 2400.200 1428.805 2400.340 1428.845 ;
        RECT 2400.700 1428.805 2401.090 1428.945 ;
        RECT 2400.200 1428.755 2401.090 1428.805 ;
        RECT 2399.390 1428.745 2399.710 1428.755 ;
        RECT 2400.200 1428.665 2400.840 1428.755 ;
        RECT 2398.930 1428.195 2399.220 1428.425 ;
        RECT 2399.870 1428.385 2400.190 1428.445 ;
        RECT 2401.830 1428.385 2402.150 1428.445 ;
        RECT 2402.520 1428.425 2402.660 1429.315 ;
        RECT 2403.310 1429.305 2403.630 1429.565 ;
        RECT 2404.030 1429.305 2404.350 1429.565 ;
        RECT 2404.600 1429.505 2404.740 1429.925 ;
        RECT 2405.230 1429.865 2405.550 1430.125 ;
        RECT 2405.770 1430.065 2406.060 1430.105 ;
        RECT 2406.230 1430.065 2406.550 1430.125 ;
        RECT 2405.770 1429.925 2406.550 1430.065 ;
        RECT 2405.770 1429.875 2406.060 1429.925 ;
        RECT 2406.230 1429.865 2406.550 1429.925 ;
        RECT 2406.710 1429.865 2407.030 1430.125 ;
        RECT 2407.190 1429.865 2407.510 1430.125 ;
        RECT 2408.190 1429.895 2408.510 1430.125 ;
        RECT 2422.230 1430.065 2422.550 1430.125 ;
        RECT 2408.190 1429.865 2409.620 1429.895 ;
        RECT 2408.280 1429.755 2409.620 1429.865 ;
        RECT 2405.770 1429.505 2406.060 1429.545 ;
        RECT 2404.600 1429.365 2406.060 1429.505 ;
        RECT 2405.770 1429.315 2406.060 1429.365 ;
        RECT 2407.710 1429.305 2408.030 1429.565 ;
        RECT 2408.280 1429.545 2408.420 1429.755 ;
        RECT 2408.210 1429.315 2408.500 1429.545 ;
        RECT 2408.930 1429.505 2409.220 1429.545 ;
        RECT 2408.930 1429.315 2409.260 1429.505 ;
        RECT 2407.210 1429.225 2407.500 1429.265 ;
        RECT 2407.710 1429.225 2407.940 1429.305 ;
        RECT 2407.210 1429.085 2407.940 1429.225 ;
        RECT 2407.210 1429.035 2407.500 1429.085 ;
        RECT 2403.050 1428.985 2403.370 1429.005 ;
        RECT 2402.810 1428.945 2403.370 1428.985 ;
        RECT 2404.050 1428.945 2404.340 1428.985 ;
        RECT 2402.810 1428.805 2404.340 1428.945 ;
        RECT 2402.810 1428.755 2403.370 1428.805 ;
        RECT 2404.050 1428.755 2404.340 1428.805 ;
        RECT 2404.530 1428.945 2404.820 1428.985 ;
        RECT 2404.530 1428.805 2405.460 1428.945 ;
        RECT 2404.530 1428.755 2404.820 1428.805 ;
        RECT 2403.050 1428.745 2403.370 1428.755 ;
        RECT 2399.870 1428.245 2402.150 1428.385 ;
        RECT 2399.870 1428.185 2400.190 1428.245 ;
        RECT 2401.830 1428.185 2402.150 1428.245 ;
        RECT 2402.330 1428.385 2402.660 1428.425 ;
        RECT 2403.310 1428.385 2403.630 1428.445 ;
        RECT 2404.030 1428.425 2404.350 1428.445 ;
        RECT 2402.330 1428.245 2403.630 1428.385 ;
        RECT 2402.330 1428.195 2402.620 1428.245 ;
        RECT 2403.310 1428.185 2403.630 1428.245 ;
        RECT 2403.810 1428.195 2404.350 1428.425 ;
        RECT 2404.030 1428.185 2404.350 1428.195 ;
        RECT 2404.750 1428.185 2405.070 1428.445 ;
        RECT 2405.320 1428.385 2405.460 1428.805 ;
        RECT 2405.750 1428.805 2406.070 1429.005 ;
        RECT 2408.450 1428.805 2408.740 1428.985 ;
        RECT 2405.750 1428.755 2408.740 1428.805 ;
        RECT 2405.750 1428.745 2408.660 1428.755 ;
        RECT 2405.840 1428.665 2408.660 1428.745 ;
        RECT 2409.120 1428.445 2409.260 1429.315 ;
        RECT 2409.480 1429.265 2409.620 1429.755 ;
        RECT 2411.140 1429.445 2411.480 1429.795 ;
        RECT 2417.470 1429.555 2417.790 1429.965 ;
        RECT 2422.230 1429.925 2423.300 1430.065 ;
        RECT 2420.480 1429.825 2421.580 1429.895 ;
        RECT 2422.230 1429.865 2422.550 1429.925 ;
        RECT 2420.410 1429.755 2421.660 1429.825 ;
        RECT 2420.410 1429.595 2420.700 1429.755 ;
        RECT 2421.370 1429.595 2421.660 1429.755 ;
        RECT 2409.410 1429.035 2409.700 1429.265 ;
        RECT 2411.230 1428.490 2411.400 1429.445 ;
        RECT 2412.745 1428.875 2413.065 1428.980 ;
        RECT 2412.720 1428.860 2413.065 1428.875 ;
        RECT 2412.715 1428.845 2413.065 1428.860 ;
        RECT 2412.545 1428.675 2413.065 1428.845 ;
        RECT 2412.720 1428.660 2413.065 1428.675 ;
        RECT 2412.720 1428.645 2413.010 1428.660 ;
        RECT 2413.520 1428.490 2413.870 1428.610 ;
        RECT 2414.880 1428.540 2415.170 1428.775 ;
        RECT 2415.870 1428.545 2416.160 1428.780 ;
        RECT 2415.870 1428.540 2416.100 1428.545 ;
        RECT 2414.880 1428.535 2415.110 1428.540 ;
        RECT 2405.990 1428.425 2406.310 1428.445 ;
        RECT 2405.770 1428.385 2406.310 1428.425 ;
        RECT 2405.320 1428.245 2406.310 1428.385 ;
        RECT 2405.770 1428.195 2406.310 1428.245 ;
        RECT 2405.990 1428.185 2406.310 1428.195 ;
        RECT 2406.590 1428.185 2407.270 1428.445 ;
        RECT 2407.710 1428.385 2408.030 1428.445 ;
        RECT 2408.210 1428.385 2408.500 1428.425 ;
        RECT 2407.710 1428.245 2408.500 1428.385 ;
        RECT 2409.120 1428.245 2409.470 1428.445 ;
        RECT 2411.230 1428.320 2413.870 1428.490 ;
        RECT 2413.350 1428.315 2413.870 1428.320 ;
        RECT 2413.520 1428.260 2413.870 1428.315 ;
        RECT 2407.710 1428.185 2408.030 1428.245 ;
        RECT 2408.210 1428.195 2408.500 1428.245 ;
        RECT 2409.150 1428.185 2409.470 1428.245 ;
        RECT 2414.510 1428.220 2414.740 1428.235 ;
        RECT 2413.090 1428.120 2413.380 1428.145 ;
        RECT 2414.480 1428.120 2414.775 1428.220 ;
        RECT 2413.090 1427.950 2414.775 1428.120 ;
        RECT 2413.090 1427.915 2413.380 1427.950 ;
        RECT 2394.530 1427.175 2394.820 1427.405 ;
        RECT 2396.320 1427.175 2396.615 1427.435 ;
        RECT 2397.310 1427.180 2397.605 1427.440 ;
        RECT 2413.150 1427.405 2413.320 1427.915 ;
        RECT 2414.480 1427.900 2414.775 1427.950 ;
        RECT 2414.510 1427.885 2414.740 1427.900 ;
        RECT 2414.940 1427.435 2415.110 1428.535 ;
        RECT 2415.930 1427.440 2416.100 1428.540 ;
        RECT 2417.550 1428.425 2417.710 1429.555 ;
        RECT 2418.430 1429.305 2418.750 1429.565 ;
        RECT 2419.550 1429.445 2419.870 1429.565 ;
        RECT 2420.890 1429.505 2421.180 1429.545 ;
        RECT 2419.550 1429.305 2420.380 1429.445 ;
        RECT 2420.890 1429.315 2421.220 1429.505 ;
        RECT 2420.170 1429.265 2420.380 1429.305 ;
        RECT 2420.170 1429.035 2420.460 1429.265 ;
        RECT 2417.950 1428.985 2418.270 1429.005 ;
        RECT 2417.950 1428.845 2418.900 1428.985 ;
        RECT 2419.360 1428.945 2419.650 1428.985 ;
        RECT 2417.950 1428.755 2418.500 1428.845 ;
        RECT 2418.760 1428.805 2418.900 1428.845 ;
        RECT 2419.260 1428.805 2419.650 1428.945 ;
        RECT 2418.760 1428.755 2419.650 1428.805 ;
        RECT 2417.950 1428.745 2418.270 1428.755 ;
        RECT 2418.760 1428.665 2419.400 1428.755 ;
        RECT 2417.490 1428.195 2417.780 1428.425 ;
        RECT 2418.430 1428.385 2418.750 1428.445 ;
        RECT 2420.390 1428.385 2420.710 1428.445 ;
        RECT 2421.080 1428.425 2421.220 1429.315 ;
        RECT 2421.870 1429.305 2422.190 1429.565 ;
        RECT 2422.590 1429.305 2422.910 1429.565 ;
        RECT 2423.160 1429.505 2423.300 1429.925 ;
        RECT 2423.790 1429.865 2424.110 1430.125 ;
        RECT 2424.330 1430.065 2424.620 1430.105 ;
        RECT 2424.790 1430.065 2425.110 1430.125 ;
        RECT 2424.330 1429.925 2425.110 1430.065 ;
        RECT 2424.330 1429.875 2424.620 1429.925 ;
        RECT 2424.790 1429.865 2425.110 1429.925 ;
        RECT 2425.270 1429.865 2425.590 1430.125 ;
        RECT 2425.750 1429.865 2426.070 1430.125 ;
        RECT 2426.750 1429.895 2427.070 1430.125 ;
        RECT 2440.790 1430.065 2441.110 1430.125 ;
        RECT 2426.750 1429.865 2428.180 1429.895 ;
        RECT 2426.840 1429.755 2428.180 1429.865 ;
        RECT 2424.330 1429.505 2424.620 1429.545 ;
        RECT 2423.160 1429.365 2424.620 1429.505 ;
        RECT 2424.330 1429.315 2424.620 1429.365 ;
        RECT 2426.270 1429.305 2426.590 1429.565 ;
        RECT 2426.840 1429.545 2426.980 1429.755 ;
        RECT 2426.770 1429.315 2427.060 1429.545 ;
        RECT 2427.490 1429.505 2427.780 1429.545 ;
        RECT 2427.490 1429.315 2427.820 1429.505 ;
        RECT 2425.770 1429.225 2426.060 1429.265 ;
        RECT 2426.270 1429.225 2426.500 1429.305 ;
        RECT 2425.770 1429.085 2426.500 1429.225 ;
        RECT 2425.770 1429.035 2426.060 1429.085 ;
        RECT 2421.610 1428.985 2421.930 1429.005 ;
        RECT 2421.370 1428.945 2421.930 1428.985 ;
        RECT 2422.610 1428.945 2422.900 1428.985 ;
        RECT 2421.370 1428.805 2422.900 1428.945 ;
        RECT 2421.370 1428.755 2421.930 1428.805 ;
        RECT 2422.610 1428.755 2422.900 1428.805 ;
        RECT 2423.090 1428.945 2423.380 1428.985 ;
        RECT 2423.090 1428.805 2424.020 1428.945 ;
        RECT 2423.090 1428.755 2423.380 1428.805 ;
        RECT 2421.610 1428.745 2421.930 1428.755 ;
        RECT 2418.430 1428.245 2420.710 1428.385 ;
        RECT 2418.430 1428.185 2418.750 1428.245 ;
        RECT 2420.390 1428.185 2420.710 1428.245 ;
        RECT 2420.890 1428.385 2421.220 1428.425 ;
        RECT 2421.870 1428.385 2422.190 1428.445 ;
        RECT 2422.590 1428.425 2422.910 1428.445 ;
        RECT 2420.890 1428.245 2422.190 1428.385 ;
        RECT 2420.890 1428.195 2421.180 1428.245 ;
        RECT 2421.870 1428.185 2422.190 1428.245 ;
        RECT 2422.370 1428.195 2422.910 1428.425 ;
        RECT 2422.590 1428.185 2422.910 1428.195 ;
        RECT 2423.310 1428.185 2423.630 1428.445 ;
        RECT 2423.880 1428.385 2424.020 1428.805 ;
        RECT 2424.310 1428.805 2424.630 1429.005 ;
        RECT 2427.010 1428.805 2427.300 1428.985 ;
        RECT 2424.310 1428.755 2427.300 1428.805 ;
        RECT 2424.310 1428.745 2427.220 1428.755 ;
        RECT 2424.400 1428.665 2427.220 1428.745 ;
        RECT 2427.680 1428.445 2427.820 1429.315 ;
        RECT 2428.040 1429.265 2428.180 1429.755 ;
        RECT 2429.700 1429.445 2430.040 1429.795 ;
        RECT 2436.030 1429.555 2436.350 1429.965 ;
        RECT 2440.790 1429.925 2441.860 1430.065 ;
        RECT 2439.040 1429.825 2440.140 1429.895 ;
        RECT 2440.790 1429.865 2441.110 1429.925 ;
        RECT 2438.970 1429.755 2440.220 1429.825 ;
        RECT 2438.970 1429.595 2439.260 1429.755 ;
        RECT 2439.930 1429.595 2440.220 1429.755 ;
        RECT 2427.970 1429.035 2428.260 1429.265 ;
        RECT 2429.790 1428.490 2429.960 1429.445 ;
        RECT 2431.305 1428.875 2431.625 1428.980 ;
        RECT 2431.280 1428.860 2431.625 1428.875 ;
        RECT 2431.275 1428.845 2431.625 1428.860 ;
        RECT 2431.105 1428.675 2431.625 1428.845 ;
        RECT 2431.280 1428.660 2431.625 1428.675 ;
        RECT 2431.280 1428.645 2431.570 1428.660 ;
        RECT 2432.080 1428.490 2432.430 1428.610 ;
        RECT 2433.440 1428.540 2433.730 1428.775 ;
        RECT 2434.430 1428.545 2434.720 1428.780 ;
        RECT 2434.430 1428.540 2434.660 1428.545 ;
        RECT 2433.440 1428.535 2433.670 1428.540 ;
        RECT 2424.550 1428.425 2424.870 1428.445 ;
        RECT 2424.330 1428.385 2424.870 1428.425 ;
        RECT 2423.880 1428.245 2424.870 1428.385 ;
        RECT 2424.330 1428.195 2424.870 1428.245 ;
        RECT 2424.550 1428.185 2424.870 1428.195 ;
        RECT 2425.150 1428.185 2425.830 1428.445 ;
        RECT 2426.270 1428.385 2426.590 1428.445 ;
        RECT 2426.770 1428.385 2427.060 1428.425 ;
        RECT 2426.270 1428.245 2427.060 1428.385 ;
        RECT 2427.680 1428.245 2428.030 1428.445 ;
        RECT 2429.790 1428.320 2432.430 1428.490 ;
        RECT 2431.910 1428.315 2432.430 1428.320 ;
        RECT 2432.080 1428.260 2432.430 1428.315 ;
        RECT 2426.270 1428.185 2426.590 1428.245 ;
        RECT 2426.770 1428.195 2427.060 1428.245 ;
        RECT 2427.710 1428.185 2428.030 1428.245 ;
        RECT 2433.070 1428.220 2433.300 1428.235 ;
        RECT 2431.650 1428.120 2431.940 1428.145 ;
        RECT 2433.040 1428.120 2433.335 1428.220 ;
        RECT 2431.650 1427.950 2433.335 1428.120 ;
        RECT 2431.650 1427.915 2431.940 1427.950 ;
        RECT 2413.090 1427.175 2413.380 1427.405 ;
        RECT 2414.880 1427.175 2415.175 1427.435 ;
        RECT 2415.870 1427.180 2416.310 1427.440 ;
        RECT 2431.710 1427.405 2431.880 1427.915 ;
        RECT 2433.040 1427.900 2433.335 1427.950 ;
        RECT 2433.070 1427.885 2433.300 1427.900 ;
        RECT 2433.500 1427.435 2433.670 1428.535 ;
        RECT 2434.490 1427.440 2434.660 1428.540 ;
        RECT 2436.110 1428.425 2436.270 1429.555 ;
        RECT 2436.990 1429.305 2437.310 1429.565 ;
        RECT 2438.110 1429.445 2438.430 1429.565 ;
        RECT 2439.450 1429.505 2439.740 1429.545 ;
        RECT 2438.110 1429.305 2438.940 1429.445 ;
        RECT 2439.450 1429.315 2439.780 1429.505 ;
        RECT 2438.730 1429.265 2438.940 1429.305 ;
        RECT 2438.730 1429.035 2439.020 1429.265 ;
        RECT 2436.510 1428.985 2436.830 1429.005 ;
        RECT 2436.510 1428.845 2437.460 1428.985 ;
        RECT 2437.920 1428.945 2438.210 1428.985 ;
        RECT 2436.510 1428.755 2437.060 1428.845 ;
        RECT 2437.320 1428.805 2437.460 1428.845 ;
        RECT 2437.820 1428.805 2438.210 1428.945 ;
        RECT 2437.320 1428.755 2438.210 1428.805 ;
        RECT 2436.510 1428.745 2436.830 1428.755 ;
        RECT 2437.320 1428.665 2437.960 1428.755 ;
        RECT 2436.050 1428.195 2436.340 1428.425 ;
        RECT 2436.990 1428.385 2437.310 1428.445 ;
        RECT 2438.950 1428.385 2439.270 1428.445 ;
        RECT 2439.640 1428.425 2439.780 1429.315 ;
        RECT 2440.430 1429.305 2440.750 1429.565 ;
        RECT 2441.150 1429.305 2441.470 1429.565 ;
        RECT 2441.720 1429.505 2441.860 1429.925 ;
        RECT 2442.350 1429.865 2442.670 1430.125 ;
        RECT 2442.890 1430.065 2443.180 1430.105 ;
        RECT 2443.350 1430.065 2443.670 1430.125 ;
        RECT 2442.890 1429.925 2443.670 1430.065 ;
        RECT 2442.890 1429.875 2443.180 1429.925 ;
        RECT 2443.350 1429.865 2443.670 1429.925 ;
        RECT 2443.830 1429.865 2444.150 1430.125 ;
        RECT 2444.310 1429.865 2444.630 1430.125 ;
        RECT 2445.310 1429.895 2445.630 1430.125 ;
        RECT 2699.285 1429.995 2699.575 1430.225 ;
        RECT 2452.990 1429.940 2453.280 1429.985 ;
        RECT 2445.310 1429.865 2446.740 1429.895 ;
        RECT 2445.400 1429.755 2446.740 1429.865 ;
        RECT 2452.990 1429.800 2454.400 1429.940 ;
        RECT 2442.890 1429.505 2443.180 1429.545 ;
        RECT 2441.720 1429.365 2443.180 1429.505 ;
        RECT 2442.890 1429.315 2443.180 1429.365 ;
        RECT 2444.830 1429.305 2445.150 1429.565 ;
        RECT 2445.400 1429.545 2445.540 1429.755 ;
        RECT 2445.330 1429.315 2445.620 1429.545 ;
        RECT 2446.050 1429.505 2446.340 1429.545 ;
        RECT 2446.050 1429.315 2446.380 1429.505 ;
        RECT 2444.330 1429.225 2444.620 1429.265 ;
        RECT 2444.830 1429.225 2445.060 1429.305 ;
        RECT 2444.330 1429.085 2445.060 1429.225 ;
        RECT 2444.330 1429.035 2444.620 1429.085 ;
        RECT 2440.170 1428.985 2440.490 1429.005 ;
        RECT 2439.930 1428.945 2440.490 1428.985 ;
        RECT 2441.170 1428.945 2441.460 1428.985 ;
        RECT 2439.930 1428.805 2441.460 1428.945 ;
        RECT 2439.930 1428.755 2440.490 1428.805 ;
        RECT 2441.170 1428.755 2441.460 1428.805 ;
        RECT 2441.650 1428.945 2441.940 1428.985 ;
        RECT 2441.650 1428.805 2442.580 1428.945 ;
        RECT 2441.650 1428.755 2441.940 1428.805 ;
        RECT 2440.170 1428.745 2440.490 1428.755 ;
        RECT 2436.990 1428.245 2439.270 1428.385 ;
        RECT 2436.990 1428.185 2437.310 1428.245 ;
        RECT 2438.950 1428.185 2439.270 1428.245 ;
        RECT 2439.450 1428.385 2439.780 1428.425 ;
        RECT 2440.430 1428.385 2440.750 1428.445 ;
        RECT 2441.150 1428.425 2441.470 1428.445 ;
        RECT 2439.450 1428.245 2440.750 1428.385 ;
        RECT 2439.450 1428.195 2439.740 1428.245 ;
        RECT 2440.430 1428.185 2440.750 1428.245 ;
        RECT 2440.930 1428.195 2441.470 1428.425 ;
        RECT 2441.150 1428.185 2441.470 1428.195 ;
        RECT 2441.870 1428.185 2442.190 1428.445 ;
        RECT 2442.440 1428.385 2442.580 1428.805 ;
        RECT 2442.870 1428.805 2443.190 1429.005 ;
        RECT 2445.570 1428.805 2445.860 1428.985 ;
        RECT 2442.870 1428.755 2445.860 1428.805 ;
        RECT 2442.870 1428.745 2445.780 1428.755 ;
        RECT 2442.960 1428.665 2445.780 1428.745 ;
        RECT 2446.240 1428.445 2446.380 1429.315 ;
        RECT 2446.600 1429.265 2446.740 1429.755 ;
        RECT 2448.260 1429.445 2448.600 1429.795 ;
        RECT 2452.990 1429.755 2453.280 1429.800 ;
        RECT 2446.530 1429.035 2446.820 1429.265 ;
        RECT 2448.350 1428.490 2448.520 1429.445 ;
        RECT 2449.865 1428.875 2450.185 1428.980 ;
        RECT 2449.840 1428.860 2450.185 1428.875 ;
        RECT 2449.835 1428.845 2450.185 1428.860 ;
        RECT 2449.665 1428.675 2450.185 1428.845 ;
        RECT 2449.840 1428.660 2450.185 1428.675 ;
        RECT 2449.840 1428.645 2450.130 1428.660 ;
        RECT 2450.640 1428.490 2450.990 1428.610 ;
        RECT 2452.000 1428.540 2452.290 1428.775 ;
        RECT 2452.990 1428.545 2453.280 1428.780 ;
        RECT 2452.990 1428.540 2453.220 1428.545 ;
        RECT 2452.000 1428.535 2452.230 1428.540 ;
        RECT 2443.110 1428.425 2443.430 1428.445 ;
        RECT 2442.890 1428.385 2443.430 1428.425 ;
        RECT 2442.440 1428.245 2443.430 1428.385 ;
        RECT 2442.890 1428.195 2443.430 1428.245 ;
        RECT 2443.110 1428.185 2443.430 1428.195 ;
        RECT 2443.710 1428.185 2444.390 1428.445 ;
        RECT 2444.830 1428.385 2445.150 1428.445 ;
        RECT 2445.330 1428.385 2445.620 1428.425 ;
        RECT 2444.830 1428.245 2445.620 1428.385 ;
        RECT 2446.240 1428.245 2446.590 1428.445 ;
        RECT 2448.350 1428.320 2450.990 1428.490 ;
        RECT 2450.470 1428.315 2450.990 1428.320 ;
        RECT 2450.640 1428.260 2450.990 1428.315 ;
        RECT 2444.830 1428.185 2445.150 1428.245 ;
        RECT 2445.330 1428.195 2445.620 1428.245 ;
        RECT 2446.270 1428.185 2446.590 1428.245 ;
        RECT 2451.630 1428.220 2451.860 1428.235 ;
        RECT 2450.210 1428.120 2450.500 1428.145 ;
        RECT 2451.600 1428.120 2451.895 1428.220 ;
        RECT 2450.210 1427.950 2451.895 1428.120 ;
        RECT 2450.210 1427.915 2450.500 1427.950 ;
        RECT 2431.650 1427.175 2431.940 1427.405 ;
        RECT 2433.440 1427.175 2433.735 1427.435 ;
        RECT 2434.390 1427.180 2434.725 1427.440 ;
        RECT 2450.270 1427.405 2450.440 1427.915 ;
        RECT 2451.600 1427.900 2451.895 1427.950 ;
        RECT 2451.630 1427.885 2451.860 1427.900 ;
        RECT 2452.060 1427.435 2452.230 1428.535 ;
        RECT 2453.050 1427.440 2453.220 1428.540 ;
        RECT 2454.260 1428.240 2454.400 1429.800 ;
        RECT 2696.970 1429.500 2697.290 1429.560 ;
        RECT 2698.365 1429.500 2698.655 1429.545 ;
        RECT 2696.970 1429.360 2698.655 1429.500 ;
        RECT 2699.360 1429.500 2699.500 1429.995 ;
        RECT 2700.740 1429.885 2700.880 1430.720 ;
        RECT 2702.030 1430.320 2702.350 1430.580 ;
        RECT 2702.490 1430.320 2702.810 1430.580 ;
        RECT 2702.965 1430.335 2703.255 1430.565 ;
        RECT 2703.040 1430.180 2703.180 1430.335 ;
        RECT 2702.580 1430.040 2703.180 1430.180 ;
        RECT 2700.665 1429.655 2700.955 1429.885 ;
        RECT 2702.580 1429.500 2702.720 1430.040 ;
        RECT 2699.360 1429.360 2702.720 1429.500 ;
        RECT 2696.970 1429.300 2697.290 1429.360 ;
        RECT 2698.365 1429.315 2698.655 1429.360 ;
        RECT 2697.905 1428.480 2698.195 1428.525 ;
        RECT 2698.350 1428.480 2698.670 1428.540 ;
        RECT 2697.905 1428.340 2698.670 1428.480 ;
        RECT 2464.750 1428.240 2465.070 1428.300 ;
        RECT 2697.905 1428.295 2698.195 1428.340 ;
        RECT 2698.350 1428.280 2698.670 1428.340 ;
        RECT 2698.810 1428.480 2699.130 1428.540 ;
        RECT 2699.285 1428.480 2699.575 1428.525 ;
        RECT 2698.810 1428.340 2699.575 1428.480 ;
        RECT 2698.810 1428.280 2699.130 1428.340 ;
        RECT 2699.285 1428.295 2699.575 1428.340 ;
        RECT 2454.260 1428.100 2465.070 1428.240 ;
        RECT 2464.750 1428.040 2465.070 1428.100 ;
        RECT 2694.670 1427.460 2694.990 1427.520 ;
        RECT 2696.985 1427.460 2697.275 1427.505 ;
        RECT 2450.210 1427.175 2450.500 1427.405 ;
        RECT 2452.000 1427.175 2452.295 1427.435 ;
        RECT 2452.990 1427.180 2453.285 1427.440 ;
        RECT 2694.670 1427.320 2697.275 1427.460 ;
        RECT 2694.670 1427.260 2694.990 1427.320 ;
        RECT 2696.985 1427.275 2697.275 1427.320 ;
        RECT 2697.430 1427.460 2697.750 1427.520 ;
        RECT 2698.825 1427.460 2699.115 1427.505 ;
        RECT 2697.430 1427.320 2699.115 1427.460 ;
        RECT 2697.430 1427.260 2697.750 1427.320 ;
        RECT 2698.825 1427.275 2699.115 1427.320 ;
        RECT 2699.730 1427.260 2700.050 1427.520 ;
        RECT 2699.730 1425.760 2700.050 1425.820 ;
        RECT 2700.665 1425.760 2700.955 1425.805 ;
        RECT 2699.730 1425.620 2700.955 1425.760 ;
        RECT 2699.730 1425.560 2700.050 1425.620 ;
        RECT 2700.665 1425.575 2700.955 1425.620 ;
        RECT 2698.810 1424.880 2699.130 1425.140 ;
        RECT 2696.970 1424.740 2697.290 1424.800 ;
        RECT 2697.445 1424.740 2697.735 1424.785 ;
        RECT 2696.970 1424.600 2697.735 1424.740 ;
        RECT 2696.970 1424.540 2697.290 1424.600 ;
        RECT 2697.445 1424.555 2697.735 1424.600 ;
        RECT 2698.350 1424.540 2698.670 1424.800 ;
        RECT 2697.890 1422.840 2698.210 1423.100 ;
        RECT 2694.670 1422.020 2694.990 1422.080 ;
        RECT 2696.985 1422.020 2697.275 1422.065 ;
        RECT 2694.670 1421.880 2697.275 1422.020 ;
        RECT 2694.670 1421.820 2694.990 1421.880 ;
        RECT 2696.985 1421.835 2697.275 1421.880 ;
        RECT 2378.730 1421.240 2379.050 1421.500 ;
        RECT 2397.130 1421.440 2397.450 1421.500 ;
        RECT 2680.490 1421.440 2680.810 1421.500 ;
        RECT 2397.130 1421.300 2680.810 1421.440 ;
        RECT 2397.130 1421.240 2397.450 1421.300 ;
        RECT 2680.490 1421.240 2680.810 1421.300 ;
        RECT 2378.820 1420.420 2378.960 1421.240 ;
        RECT 2415.990 1420.900 2416.310 1421.160 ;
        RECT 2611.490 1421.100 2611.810 1421.160 ;
        RECT 2428.730 1420.960 2611.810 1421.100 ;
        RECT 2416.080 1420.760 2416.220 1420.900 ;
        RECT 2428.730 1420.760 2428.870 1420.960 ;
        RECT 2611.490 1420.900 2611.810 1420.960 ;
        RECT 2416.080 1420.620 2428.870 1420.760 ;
        RECT 2434.390 1420.760 2434.710 1420.820 ;
        RECT 2618.390 1420.760 2618.710 1420.820 ;
        RECT 2434.390 1420.620 2618.710 1420.760 ;
        RECT 2434.390 1420.560 2434.710 1420.620 ;
        RECT 2618.390 1420.560 2618.710 1420.620 ;
        RECT 2507.990 1420.420 2508.310 1420.480 ;
        RECT 2378.820 1420.280 2508.310 1420.420 ;
        RECT 2507.990 1420.220 2508.310 1420.280 ;
        RECT 2697.905 1417.600 2698.195 1417.645 ;
        RECT 2698.810 1417.600 2699.130 1417.660 ;
        RECT 2697.905 1417.460 2699.130 1417.600 ;
        RECT 2697.905 1417.415 2698.195 1417.460 ;
        RECT 2698.810 1417.400 2699.130 1417.460 ;
        RECT 2523.545 1416.755 2523.865 1417.015 ;
        RECT 2694.670 1416.580 2694.990 1416.640 ;
        RECT 2696.985 1416.580 2697.275 1416.625 ;
        RECT 2694.670 1416.440 2697.275 1416.580 ;
        RECT 2694.670 1416.380 2694.990 1416.440 ;
        RECT 2696.985 1416.395 2697.275 1416.440 ;
        RECT 2698.350 1412.160 2698.670 1412.220 ;
        RECT 2699.285 1412.160 2699.575 1412.205 ;
        RECT 2698.350 1412.020 2699.575 1412.160 ;
        RECT 2698.350 1411.960 2698.670 1412.020 ;
        RECT 2699.285 1411.975 2699.575 1412.020 ;
        RECT 2702.490 1411.960 2702.810 1412.220 ;
        RECT 2697.905 1411.820 2698.195 1411.865 ;
        RECT 2702.580 1411.820 2702.720 1411.960 ;
        RECT 2697.905 1411.680 2702.720 1411.820 ;
        RECT 2697.905 1411.635 2698.195 1411.680 ;
        RECT 2694.670 1411.140 2694.990 1411.200 ;
        RECT 2696.985 1411.140 2697.275 1411.185 ;
        RECT 2694.670 1411.000 2697.275 1411.140 ;
        RECT 2694.670 1410.940 2694.990 1411.000 ;
        RECT 2696.985 1410.955 2697.275 1411.000 ;
        RECT 2698.350 1410.940 2698.670 1411.200 ;
        RECT 2523.545 1409.225 2523.865 1409.485 ;
        RECT 2523.545 1403.245 2523.865 1403.505 ;
        RECT 2523.545 1394.830 2523.865 1395.090 ;
        RECT 2369.540 1335.060 2369.830 1335.290 ;
        RECT 2377.055 1335.060 2377.345 1335.290 ;
        RECT 2382.670 1335.060 2382.960 1335.290 ;
        RECT 2369.600 1334.610 2369.770 1335.060 ;
        RECT 2377.115 1334.715 2377.285 1335.060 ;
        RECT 2369.510 1334.320 2369.860 1334.610 ;
        RECT 2377.015 1334.345 2377.385 1334.715 ;
        RECT 2382.730 1334.580 2382.900 1335.060 ;
        RECT 2384.460 1335.030 2384.755 1335.290 ;
        RECT 2385.450 1335.030 2385.745 1335.290 ;
        RECT 2392.315 1335.060 2392.605 1335.290 ;
        RECT 2397.930 1335.060 2398.220 1335.290 ;
        RECT 2384.090 1334.630 2384.320 1334.645 ;
        RECT 2384.045 1334.580 2384.355 1334.630 ;
        RECT 2382.730 1334.550 2384.355 1334.580 ;
        RECT 2382.670 1334.410 2384.355 1334.550 ;
        RECT 2377.055 1334.320 2377.345 1334.345 ;
        RECT 2382.670 1334.320 2382.960 1334.410 ;
        RECT 2384.045 1334.320 2384.355 1334.410 ;
        RECT 2384.090 1334.290 2384.320 1334.320 ;
        RECT 2377.685 1334.180 2378.035 1334.245 ;
        RECT 2383.125 1334.180 2383.450 1334.270 ;
        RECT 2377.485 1334.150 2378.035 1334.180 ;
        RECT 2383.100 1334.150 2383.450 1334.180 ;
        RECT 2377.315 1334.145 2378.035 1334.150 ;
        RECT 2382.930 1334.145 2383.450 1334.150 ;
        RECT 2377.315 1333.980 2383.450 1334.145 ;
        RECT 2377.375 1333.975 2383.450 1333.980 ;
        RECT 2377.485 1333.950 2378.035 1333.975 ;
        RECT 2383.100 1333.950 2383.450 1333.975 ;
        RECT 2377.685 1333.895 2378.035 1333.950 ;
        RECT 2383.125 1333.945 2383.450 1333.950 ;
        RECT 2384.520 1333.930 2384.690 1335.030 ;
        RECT 2385.510 1334.300 2385.680 1335.030 ;
        RECT 2392.375 1334.715 2392.545 1335.060 ;
        RECT 2392.275 1334.345 2392.645 1334.715 ;
        RECT 2397.990 1334.580 2398.160 1335.060 ;
        RECT 2399.720 1335.030 2400.015 1335.290 ;
        RECT 2400.710 1335.030 2401.005 1335.290 ;
        RECT 2407.575 1335.060 2407.865 1335.290 ;
        RECT 2413.190 1335.060 2413.480 1335.290 ;
        RECT 2399.350 1334.630 2399.580 1334.645 ;
        RECT 2399.305 1334.580 2399.615 1334.630 ;
        RECT 2397.990 1334.550 2399.615 1334.580 ;
        RECT 2397.930 1334.410 2399.615 1334.550 ;
        RECT 2392.315 1334.320 2392.605 1334.345 ;
        RECT 2397.930 1334.320 2398.220 1334.410 ;
        RECT 2399.305 1334.320 2399.615 1334.410 ;
        RECT 2385.505 1333.950 2385.855 1334.300 ;
        RECT 2399.350 1334.290 2399.580 1334.320 ;
        RECT 2392.945 1334.180 2393.295 1334.255 ;
        RECT 2398.385 1334.180 2398.710 1334.270 ;
        RECT 2392.745 1334.150 2393.295 1334.180 ;
        RECT 2398.360 1334.150 2398.710 1334.180 ;
        RECT 2392.575 1334.145 2393.295 1334.150 ;
        RECT 2398.190 1334.145 2398.710 1334.150 ;
        RECT 2392.575 1333.980 2398.710 1334.145 ;
        RECT 2392.635 1333.975 2398.710 1333.980 ;
        RECT 2392.745 1333.950 2393.295 1333.975 ;
        RECT 2398.360 1333.950 2398.710 1333.975 ;
        RECT 2385.505 1333.930 2385.800 1333.950 ;
        RECT 2384.460 1333.925 2384.690 1333.930 ;
        RECT 2369.135 1333.790 2369.485 1333.865 ;
        RECT 2382.325 1333.820 2382.645 1333.835 ;
        RECT 2382.300 1333.790 2382.645 1333.820 ;
        RECT 2368.995 1333.620 2369.485 1333.790 ;
        RECT 2382.125 1333.620 2382.645 1333.790 ;
        RECT 2384.460 1333.690 2384.750 1333.925 ;
        RECT 2385.450 1333.860 2385.800 1333.930 ;
        RECT 2392.945 1333.905 2393.295 1333.950 ;
        RECT 2398.385 1333.945 2398.710 1333.950 ;
        RECT 2399.780 1333.930 2399.950 1335.030 ;
        RECT 2400.770 1334.305 2400.940 1335.030 ;
        RECT 2407.635 1334.715 2407.805 1335.060 ;
        RECT 2407.535 1334.345 2407.905 1334.715 ;
        RECT 2413.250 1334.580 2413.420 1335.060 ;
        RECT 2414.980 1335.030 2415.275 1335.290 ;
        RECT 2415.970 1335.030 2416.265 1335.290 ;
        RECT 2422.835 1335.060 2423.125 1335.290 ;
        RECT 2428.450 1335.060 2428.740 1335.290 ;
        RECT 2414.610 1334.630 2414.840 1334.645 ;
        RECT 2414.565 1334.580 2414.875 1334.630 ;
        RECT 2413.250 1334.550 2414.875 1334.580 ;
        RECT 2413.190 1334.410 2414.875 1334.550 ;
        RECT 2407.575 1334.320 2407.865 1334.345 ;
        RECT 2413.190 1334.320 2413.480 1334.410 ;
        RECT 2414.565 1334.320 2414.875 1334.410 ;
        RECT 2400.760 1333.950 2401.115 1334.305 ;
        RECT 2414.610 1334.290 2414.840 1334.320 ;
        RECT 2408.205 1334.180 2408.555 1334.255 ;
        RECT 2413.645 1334.180 2413.970 1334.270 ;
        RECT 2408.005 1334.150 2408.555 1334.180 ;
        RECT 2413.620 1334.150 2413.970 1334.180 ;
        RECT 2407.835 1334.145 2408.555 1334.150 ;
        RECT 2413.450 1334.145 2413.970 1334.150 ;
        RECT 2407.835 1333.980 2413.970 1334.145 ;
        RECT 2407.895 1333.975 2413.970 1333.980 ;
        RECT 2408.005 1333.950 2408.555 1333.975 ;
        RECT 2413.620 1333.950 2413.970 1333.975 ;
        RECT 2400.760 1333.930 2401.060 1333.950 ;
        RECT 2399.720 1333.925 2399.950 1333.930 ;
        RECT 2385.450 1333.690 2385.740 1333.860 ;
        RECT 2397.585 1333.820 2397.905 1333.835 ;
        RECT 2397.560 1333.790 2397.905 1333.820 ;
        RECT 2397.385 1333.620 2397.905 1333.790 ;
        RECT 2399.720 1333.690 2400.010 1333.925 ;
        RECT 2400.710 1333.865 2401.060 1333.930 ;
        RECT 2408.205 1333.905 2408.555 1333.950 ;
        RECT 2413.645 1333.945 2413.970 1333.950 ;
        RECT 2415.040 1333.930 2415.210 1335.030 ;
        RECT 2416.030 1334.300 2416.200 1335.030 ;
        RECT 2422.895 1334.715 2423.065 1335.060 ;
        RECT 2422.795 1334.345 2423.165 1334.715 ;
        RECT 2428.510 1334.580 2428.680 1335.060 ;
        RECT 2430.240 1335.030 2430.535 1335.290 ;
        RECT 2431.230 1335.030 2431.525 1335.290 ;
        RECT 2438.095 1335.060 2438.385 1335.290 ;
        RECT 2443.710 1335.060 2444.000 1335.290 ;
        RECT 2429.870 1334.630 2430.100 1334.645 ;
        RECT 2429.825 1334.580 2430.135 1334.630 ;
        RECT 2428.510 1334.550 2430.135 1334.580 ;
        RECT 2428.450 1334.410 2430.135 1334.550 ;
        RECT 2422.835 1334.320 2423.125 1334.345 ;
        RECT 2428.450 1334.320 2428.740 1334.410 ;
        RECT 2429.825 1334.320 2430.135 1334.410 ;
        RECT 2415.980 1333.950 2416.330 1334.300 ;
        RECT 2429.870 1334.290 2430.100 1334.320 ;
        RECT 2423.470 1334.180 2423.820 1334.255 ;
        RECT 2428.905 1334.180 2429.230 1334.270 ;
        RECT 2423.265 1334.150 2423.820 1334.180 ;
        RECT 2428.880 1334.150 2429.230 1334.180 ;
        RECT 2423.095 1334.145 2423.820 1334.150 ;
        RECT 2428.710 1334.145 2429.230 1334.150 ;
        RECT 2423.095 1333.980 2429.230 1334.145 ;
        RECT 2423.155 1333.975 2429.230 1333.980 ;
        RECT 2423.265 1333.950 2423.820 1333.975 ;
        RECT 2428.880 1333.950 2429.230 1333.975 ;
        RECT 2415.980 1333.930 2416.320 1333.950 ;
        RECT 2414.980 1333.925 2415.210 1333.930 ;
        RECT 2400.710 1333.690 2401.000 1333.865 ;
        RECT 2412.845 1333.820 2413.165 1333.835 ;
        RECT 2412.820 1333.790 2413.165 1333.820 ;
        RECT 2412.645 1333.620 2413.165 1333.790 ;
        RECT 2414.980 1333.690 2415.270 1333.925 ;
        RECT 2415.970 1333.860 2416.320 1333.930 ;
        RECT 2423.470 1333.905 2423.820 1333.950 ;
        RECT 2428.905 1333.945 2429.230 1333.950 ;
        RECT 2430.300 1333.930 2430.470 1335.030 ;
        RECT 2431.290 1334.300 2431.460 1335.030 ;
        RECT 2438.155 1334.715 2438.325 1335.060 ;
        RECT 2438.055 1334.345 2438.425 1334.715 ;
        RECT 2443.770 1334.580 2443.940 1335.060 ;
        RECT 2445.500 1335.030 2445.795 1335.290 ;
        RECT 2446.490 1335.030 2446.785 1335.290 ;
        RECT 2445.130 1334.630 2445.360 1334.645 ;
        RECT 2445.085 1334.580 2445.395 1334.630 ;
        RECT 2443.770 1334.550 2445.395 1334.580 ;
        RECT 2443.710 1334.410 2445.395 1334.550 ;
        RECT 2438.095 1334.320 2438.385 1334.345 ;
        RECT 2443.710 1334.320 2444.000 1334.410 ;
        RECT 2445.085 1334.320 2445.395 1334.410 ;
        RECT 2431.240 1333.950 2431.590 1334.300 ;
        RECT 2445.130 1334.290 2445.360 1334.320 ;
        RECT 2438.725 1334.180 2439.075 1334.255 ;
        RECT 2444.165 1334.180 2444.490 1334.270 ;
        RECT 2438.525 1334.150 2439.075 1334.180 ;
        RECT 2444.140 1334.150 2444.490 1334.180 ;
        RECT 2438.355 1334.145 2439.075 1334.150 ;
        RECT 2443.970 1334.145 2444.490 1334.150 ;
        RECT 2438.355 1333.980 2444.490 1334.145 ;
        RECT 2438.415 1333.975 2444.490 1333.980 ;
        RECT 2438.525 1333.950 2439.075 1333.975 ;
        RECT 2444.140 1333.950 2444.490 1333.975 ;
        RECT 2431.240 1333.930 2431.580 1333.950 ;
        RECT 2430.240 1333.925 2430.470 1333.930 ;
        RECT 2415.970 1333.690 2416.260 1333.860 ;
        RECT 2428.105 1333.820 2428.425 1333.835 ;
        RECT 2428.080 1333.790 2428.425 1333.820 ;
        RECT 2427.905 1333.620 2428.425 1333.790 ;
        RECT 2430.240 1333.690 2430.530 1333.925 ;
        RECT 2431.230 1333.860 2431.580 1333.930 ;
        RECT 2438.725 1333.905 2439.075 1333.950 ;
        RECT 2444.165 1333.945 2444.490 1333.950 ;
        RECT 2445.560 1333.930 2445.730 1335.030 ;
        RECT 2446.525 1334.995 2446.785 1335.030 ;
        RECT 2446.525 1334.915 2446.845 1334.995 ;
        RECT 2446.525 1334.565 2446.875 1334.915 ;
        RECT 2446.550 1333.930 2446.720 1334.565 ;
        RECT 2445.500 1333.925 2445.730 1333.930 ;
        RECT 2446.490 1333.925 2446.720 1333.930 ;
        RECT 2431.230 1333.690 2431.520 1333.860 ;
        RECT 2443.365 1333.820 2443.685 1333.835 ;
        RECT 2443.340 1333.790 2443.685 1333.820 ;
        RECT 2443.165 1333.620 2443.685 1333.790 ;
        RECT 2445.500 1333.690 2445.790 1333.925 ;
        RECT 2446.490 1333.690 2446.780 1333.925 ;
        RECT 2369.135 1333.575 2369.485 1333.620 ;
        RECT 2382.300 1333.590 2382.645 1333.620 ;
        RECT 2397.560 1333.590 2397.905 1333.620 ;
        RECT 2412.820 1333.590 2413.165 1333.620 ;
        RECT 2428.080 1333.590 2428.425 1333.620 ;
        RECT 2443.340 1333.590 2443.685 1333.620 ;
        RECT 2382.325 1333.545 2382.645 1333.590 ;
        RECT 2397.585 1333.545 2397.905 1333.590 ;
        RECT 2412.845 1333.545 2413.165 1333.590 ;
        RECT 2428.105 1333.545 2428.425 1333.590 ;
        RECT 2443.365 1333.545 2443.685 1333.590 ;
        RECT 2373.715 1329.895 2374.005 1330.105 ;
        RECT 2372.825 1329.875 2374.005 1329.895 ;
        RECT 2371.805 1329.585 2372.125 1329.845 ;
        RECT 2372.825 1329.825 2373.925 1329.875 ;
        RECT 2374.655 1329.865 2374.975 1330.125 ;
        RECT 2375.255 1330.105 2375.575 1330.125 ;
        RECT 2375.155 1329.875 2375.575 1330.105 ;
        RECT 2375.255 1329.865 2375.575 1329.875 ;
        RECT 2376.815 1330.105 2377.150 1330.125 ;
        RECT 2376.815 1329.875 2377.340 1330.105 ;
        RECT 2378.995 1330.065 2379.285 1330.105 ;
        RECT 2379.425 1330.065 2379.745 1330.125 ;
        RECT 2378.995 1329.925 2379.745 1330.065 ;
        RECT 2378.995 1329.875 2379.285 1329.925 ;
        RECT 2376.815 1329.865 2377.150 1329.875 ;
        RECT 2379.425 1329.865 2379.745 1329.925 ;
        RECT 2388.975 1329.895 2389.265 1330.105 ;
        RECT 2388.085 1329.875 2389.265 1329.895 ;
        RECT 2372.755 1329.755 2373.925 1329.825 ;
        RECT 2372.755 1329.595 2373.045 1329.755 ;
        RECT 2375.185 1329.585 2375.355 1329.685 ;
        RECT 2377.565 1329.585 2377.885 1329.845 ;
        RECT 2387.065 1329.585 2387.385 1329.845 ;
        RECT 2388.085 1329.825 2389.185 1329.875 ;
        RECT 2389.915 1329.865 2390.235 1330.125 ;
        RECT 2390.515 1330.105 2390.835 1330.125 ;
        RECT 2390.415 1329.875 2390.835 1330.105 ;
        RECT 2390.515 1329.865 2390.835 1329.875 ;
        RECT 2392.075 1330.105 2392.410 1330.125 ;
        RECT 2392.075 1329.875 2392.600 1330.105 ;
        RECT 2394.255 1330.065 2394.545 1330.105 ;
        RECT 2394.685 1330.065 2395.005 1330.125 ;
        RECT 2394.255 1329.925 2395.005 1330.065 ;
        RECT 2394.255 1329.875 2394.545 1329.925 ;
        RECT 2392.075 1329.865 2392.410 1329.875 ;
        RECT 2394.685 1329.865 2395.005 1329.925 ;
        RECT 2404.235 1329.895 2404.525 1330.105 ;
        RECT 2403.345 1329.875 2404.525 1329.895 ;
        RECT 2388.015 1329.755 2389.185 1329.825 ;
        RECT 2388.015 1329.595 2388.305 1329.755 ;
        RECT 2390.445 1329.585 2390.615 1329.685 ;
        RECT 2392.825 1329.585 2393.145 1329.845 ;
        RECT 2402.325 1329.585 2402.645 1329.845 ;
        RECT 2403.345 1329.825 2404.445 1329.875 ;
        RECT 2405.175 1329.865 2405.495 1330.125 ;
        RECT 2405.775 1330.105 2406.095 1330.125 ;
        RECT 2405.675 1329.875 2406.095 1330.105 ;
        RECT 2405.775 1329.865 2406.095 1329.875 ;
        RECT 2407.335 1330.105 2407.670 1330.125 ;
        RECT 2407.335 1329.875 2407.860 1330.105 ;
        RECT 2409.515 1330.065 2409.805 1330.105 ;
        RECT 2409.945 1330.065 2410.265 1330.125 ;
        RECT 2409.515 1329.925 2410.265 1330.065 ;
        RECT 2409.515 1329.875 2409.805 1329.925 ;
        RECT 2407.335 1329.865 2407.670 1329.875 ;
        RECT 2409.945 1329.865 2410.265 1329.925 ;
        RECT 2419.495 1329.895 2419.785 1330.105 ;
        RECT 2418.605 1329.875 2419.785 1329.895 ;
        RECT 2403.275 1329.755 2404.445 1329.825 ;
        RECT 2403.275 1329.595 2403.565 1329.755 ;
        RECT 2405.705 1329.585 2405.875 1329.685 ;
        RECT 2408.085 1329.585 2408.405 1329.845 ;
        RECT 2417.585 1329.585 2417.905 1329.845 ;
        RECT 2418.605 1329.825 2419.705 1329.875 ;
        RECT 2420.435 1329.865 2420.755 1330.125 ;
        RECT 2421.035 1330.105 2421.355 1330.125 ;
        RECT 2420.935 1329.875 2421.355 1330.105 ;
        RECT 2421.035 1329.865 2421.355 1329.875 ;
        RECT 2422.595 1330.105 2422.930 1330.125 ;
        RECT 2422.595 1329.875 2423.120 1330.105 ;
        RECT 2424.775 1330.065 2425.065 1330.105 ;
        RECT 2425.205 1330.065 2425.525 1330.125 ;
        RECT 2424.775 1329.925 2425.525 1330.065 ;
        RECT 2424.775 1329.875 2425.065 1329.925 ;
        RECT 2422.595 1329.865 2422.930 1329.875 ;
        RECT 2425.205 1329.865 2425.525 1329.925 ;
        RECT 2434.755 1329.895 2435.045 1330.105 ;
        RECT 2433.865 1329.875 2435.045 1329.895 ;
        RECT 2418.535 1329.755 2419.705 1329.825 ;
        RECT 2418.535 1329.595 2418.825 1329.755 ;
        RECT 2420.965 1329.585 2421.135 1329.685 ;
        RECT 2423.345 1329.585 2423.665 1329.845 ;
        RECT 2432.845 1329.585 2433.165 1329.845 ;
        RECT 2433.865 1329.825 2434.965 1329.875 ;
        RECT 2435.695 1329.865 2436.015 1330.125 ;
        RECT 2436.295 1330.105 2436.615 1330.125 ;
        RECT 2436.195 1329.875 2436.615 1330.105 ;
        RECT 2436.295 1329.865 2436.615 1329.875 ;
        RECT 2437.855 1330.105 2438.190 1330.125 ;
        RECT 2437.855 1329.875 2438.380 1330.105 ;
        RECT 2440.035 1330.065 2440.325 1330.105 ;
        RECT 2440.465 1330.065 2440.785 1330.125 ;
        RECT 2440.035 1329.925 2440.785 1330.065 ;
        RECT 2459.690 1329.980 2460.010 1330.040 ;
        RECT 2440.035 1329.875 2440.325 1329.925 ;
        RECT 2437.855 1329.865 2438.190 1329.875 ;
        RECT 2440.465 1329.865 2440.785 1329.925 ;
        RECT 2433.795 1329.755 2434.965 1329.825 ;
        RECT 2433.795 1329.595 2434.085 1329.755 ;
        RECT 2436.225 1329.585 2436.395 1329.685 ;
        RECT 2438.605 1329.585 2438.925 1329.845 ;
        RECT 2446.440 1329.840 2460.010 1329.980 ;
        RECT 2374.175 1329.545 2374.495 1329.565 ;
        RECT 2373.235 1329.505 2373.525 1329.545 ;
        RECT 2373.235 1329.315 2373.685 1329.505 ;
        RECT 2372.495 1329.025 2372.815 1329.285 ;
        RECT 2372.975 1328.745 2373.295 1329.005 ;
        RECT 2373.545 1328.985 2373.685 1329.315 ;
        RECT 2374.175 1329.315 2374.725 1329.545 ;
        RECT 2374.865 1329.445 2377.045 1329.585 ;
        RECT 2389.435 1329.545 2389.755 1329.565 ;
        RECT 2374.865 1329.365 2376.165 1329.445 ;
        RECT 2374.175 1329.305 2374.495 1329.315 ;
        RECT 2374.865 1329.085 2375.205 1329.365 ;
        RECT 2375.875 1329.315 2376.165 1329.365 ;
        RECT 2374.915 1329.035 2375.205 1329.085 ;
        RECT 2376.335 1329.025 2376.655 1329.285 ;
        RECT 2373.545 1328.845 2373.805 1328.985 ;
        RECT 2371.805 1328.185 2372.125 1328.445 ;
        RECT 2373.665 1328.425 2373.805 1328.845 ;
        RECT 2373.955 1328.945 2374.245 1328.985 ;
        RECT 2374.415 1328.945 2374.735 1329.005 ;
        RECT 2373.955 1328.805 2374.735 1328.945 ;
        RECT 2373.955 1328.755 2374.245 1328.805 ;
        RECT 2374.415 1328.745 2374.735 1328.805 ;
        RECT 2375.395 1328.755 2375.685 1328.985 ;
        RECT 2375.545 1328.505 2375.685 1328.755 ;
        RECT 2375.855 1328.745 2376.175 1329.005 ;
        RECT 2376.905 1328.805 2377.045 1329.445 ;
        RECT 2378.755 1329.505 2379.045 1329.545 ;
        RECT 2388.495 1329.505 2388.785 1329.545 ;
        RECT 2378.755 1329.365 2379.325 1329.505 ;
        RECT 2377.385 1329.285 2378.485 1329.365 ;
        RECT 2378.755 1329.315 2379.045 1329.365 ;
        RECT 2377.195 1329.265 2378.485 1329.285 ;
        RECT 2379.185 1329.265 2379.445 1329.365 ;
        RECT 2385.630 1329.345 2385.950 1329.360 ;
        RECT 2377.195 1329.225 2378.565 1329.265 ;
        RECT 2379.185 1329.225 2379.525 1329.265 ;
        RECT 2377.195 1329.035 2377.605 1329.225 ;
        RECT 2378.275 1329.035 2378.565 1329.225 ;
        RECT 2379.235 1329.035 2379.525 1329.225 ;
        RECT 2377.195 1329.025 2377.515 1329.035 ;
        RECT 2377.795 1328.805 2378.085 1328.985 ;
        RECT 2376.905 1328.755 2378.085 1328.805 ;
        RECT 2376.905 1328.705 2378.005 1328.755 ;
        RECT 2378.735 1328.745 2379.055 1329.005 ;
        RECT 2380.720 1328.995 2381.060 1329.345 ;
        RECT 2385.445 1329.115 2385.950 1329.345 ;
        RECT 2388.495 1329.315 2388.945 1329.505 ;
        RECT 2385.630 1329.100 2385.950 1329.115 ;
        RECT 2387.755 1329.025 2388.075 1329.285 ;
        RECT 2376.835 1328.665 2378.005 1328.705 ;
        RECT 2375.545 1328.445 2375.845 1328.505 ;
        RECT 2376.835 1328.455 2377.125 1328.665 ;
        RECT 2380.810 1328.490 2380.980 1328.995 ;
        RECT 2382.325 1328.875 2382.645 1328.980 ;
        RECT 2382.300 1328.860 2382.645 1328.875 ;
        RECT 2382.290 1328.845 2382.645 1328.860 ;
        RECT 2382.125 1328.675 2382.645 1328.845 ;
        RECT 2382.300 1328.660 2382.645 1328.675 ;
        RECT 2382.300 1328.645 2382.590 1328.660 ;
        RECT 2383.100 1328.490 2383.450 1328.610 ;
        RECT 2384.460 1328.540 2384.750 1328.775 ;
        RECT 2385.445 1328.540 2385.735 1328.775 ;
        RECT 2388.235 1328.745 2388.555 1329.005 ;
        RECT 2388.805 1328.985 2388.945 1329.315 ;
        RECT 2389.435 1329.315 2389.985 1329.545 ;
        RECT 2390.125 1329.445 2392.305 1329.585 ;
        RECT 2404.695 1329.545 2405.015 1329.565 ;
        RECT 2390.125 1329.365 2391.425 1329.445 ;
        RECT 2389.435 1329.305 2389.755 1329.315 ;
        RECT 2390.125 1329.085 2390.465 1329.365 ;
        RECT 2391.135 1329.315 2391.425 1329.365 ;
        RECT 2390.175 1329.035 2390.465 1329.085 ;
        RECT 2391.595 1329.025 2391.915 1329.285 ;
        RECT 2388.805 1328.845 2389.065 1328.985 ;
        RECT 2384.460 1328.535 2384.690 1328.540 ;
        RECT 2385.445 1328.535 2385.675 1328.540 ;
        RECT 2373.665 1328.385 2374.005 1328.425 ;
        RECT 2374.535 1328.385 2374.855 1328.445 ;
        RECT 2373.665 1328.245 2374.855 1328.385 ;
        RECT 2373.715 1328.195 2374.005 1328.245 ;
        RECT 2374.535 1328.185 2374.855 1328.245 ;
        RECT 2375.005 1328.185 2375.405 1328.445 ;
        RECT 2375.545 1328.385 2375.935 1328.445 ;
        RECT 2376.335 1328.425 2376.655 1328.445 ;
        RECT 2376.115 1328.385 2376.655 1328.425 ;
        RECT 2375.545 1328.365 2376.655 1328.385 ;
        RECT 2375.615 1328.245 2376.655 1328.365 ;
        RECT 2375.615 1328.185 2375.935 1328.245 ;
        RECT 2376.115 1328.195 2376.655 1328.245 ;
        RECT 2376.335 1328.185 2376.655 1328.195 ;
        RECT 2377.565 1328.385 2377.885 1328.445 ;
        RECT 2378.035 1328.385 2378.325 1328.425 ;
        RECT 2377.565 1328.245 2378.325 1328.385 ;
        RECT 2377.565 1328.185 2377.885 1328.245 ;
        RECT 2378.035 1328.195 2378.325 1328.245 ;
        RECT 2378.995 1328.385 2379.285 1328.425 ;
        RECT 2379.425 1328.385 2379.745 1328.445 ;
        RECT 2378.995 1328.245 2379.745 1328.385 ;
        RECT 2380.810 1328.320 2383.450 1328.490 ;
        RECT 2382.930 1328.315 2383.450 1328.320 ;
        RECT 2383.100 1328.260 2383.450 1328.315 ;
        RECT 2378.995 1328.195 2379.285 1328.245 ;
        RECT 2379.425 1328.185 2379.745 1328.245 ;
        RECT 2384.090 1328.205 2384.320 1328.230 ;
        RECT 2382.670 1328.120 2382.960 1328.145 ;
        RECT 2384.060 1328.120 2384.350 1328.205 ;
        RECT 2382.670 1327.950 2384.350 1328.120 ;
        RECT 2382.670 1327.915 2382.960 1327.950 ;
        RECT 2382.730 1327.405 2382.900 1327.915 ;
        RECT 2384.060 1327.900 2384.350 1327.950 ;
        RECT 2384.090 1327.880 2384.320 1327.900 ;
        RECT 2384.520 1327.435 2384.690 1328.535 ;
        RECT 2385.505 1327.435 2385.675 1328.535 ;
        RECT 2387.065 1328.185 2387.385 1328.445 ;
        RECT 2388.925 1328.425 2389.065 1328.845 ;
        RECT 2389.215 1328.945 2389.505 1328.985 ;
        RECT 2389.675 1328.945 2389.995 1329.005 ;
        RECT 2389.215 1328.805 2389.995 1328.945 ;
        RECT 2389.215 1328.755 2389.505 1328.805 ;
        RECT 2389.675 1328.745 2389.995 1328.805 ;
        RECT 2390.655 1328.755 2390.945 1328.985 ;
        RECT 2390.805 1328.505 2390.945 1328.755 ;
        RECT 2391.115 1328.745 2391.435 1329.005 ;
        RECT 2392.165 1328.805 2392.305 1329.445 ;
        RECT 2394.015 1329.505 2394.305 1329.545 ;
        RECT 2403.755 1329.505 2404.045 1329.545 ;
        RECT 2394.015 1329.365 2394.585 1329.505 ;
        RECT 2392.645 1329.285 2393.745 1329.365 ;
        RECT 2394.015 1329.315 2394.305 1329.365 ;
        RECT 2392.455 1329.265 2393.745 1329.285 ;
        RECT 2394.445 1329.265 2394.705 1329.365 ;
        RECT 2392.455 1329.225 2393.825 1329.265 ;
        RECT 2394.445 1329.225 2394.785 1329.265 ;
        RECT 2392.455 1329.035 2392.865 1329.225 ;
        RECT 2393.535 1329.035 2393.825 1329.225 ;
        RECT 2394.495 1329.035 2394.785 1329.225 ;
        RECT 2392.455 1329.025 2392.775 1329.035 ;
        RECT 2393.055 1328.805 2393.345 1328.985 ;
        RECT 2392.165 1328.755 2393.345 1328.805 ;
        RECT 2392.165 1328.705 2393.265 1328.755 ;
        RECT 2393.995 1328.745 2394.315 1329.005 ;
        RECT 2395.980 1328.995 2396.320 1329.345 ;
        RECT 2403.755 1329.315 2404.205 1329.505 ;
        RECT 2403.015 1329.025 2403.335 1329.285 ;
        RECT 2392.095 1328.665 2393.265 1328.705 ;
        RECT 2390.805 1328.445 2391.105 1328.505 ;
        RECT 2392.095 1328.455 2392.385 1328.665 ;
        RECT 2396.070 1328.490 2396.240 1328.995 ;
        RECT 2397.585 1328.875 2397.905 1328.980 ;
        RECT 2397.560 1328.860 2397.905 1328.875 ;
        RECT 2397.550 1328.845 2397.905 1328.860 ;
        RECT 2397.385 1328.675 2397.905 1328.845 ;
        RECT 2397.560 1328.660 2397.905 1328.675 ;
        RECT 2397.560 1328.645 2397.850 1328.660 ;
        RECT 2398.360 1328.490 2398.710 1328.610 ;
        RECT 2399.720 1328.540 2400.010 1328.775 ;
        RECT 2400.705 1328.540 2400.995 1328.775 ;
        RECT 2403.495 1328.745 2403.815 1329.005 ;
        RECT 2404.065 1328.985 2404.205 1329.315 ;
        RECT 2404.695 1329.315 2405.245 1329.545 ;
        RECT 2405.385 1329.445 2407.565 1329.585 ;
        RECT 2419.955 1329.545 2420.275 1329.565 ;
        RECT 2405.385 1329.365 2406.685 1329.445 ;
        RECT 2404.695 1329.305 2405.015 1329.315 ;
        RECT 2405.385 1329.085 2405.725 1329.365 ;
        RECT 2406.395 1329.315 2406.685 1329.365 ;
        RECT 2405.435 1329.035 2405.725 1329.085 ;
        RECT 2406.855 1329.025 2407.175 1329.285 ;
        RECT 2404.065 1328.845 2404.325 1328.985 ;
        RECT 2399.720 1328.535 2399.950 1328.540 ;
        RECT 2400.705 1328.535 2400.935 1328.540 ;
        RECT 2388.925 1328.385 2389.265 1328.425 ;
        RECT 2389.795 1328.385 2390.115 1328.445 ;
        RECT 2388.925 1328.245 2390.115 1328.385 ;
        RECT 2388.975 1328.195 2389.265 1328.245 ;
        RECT 2389.795 1328.185 2390.115 1328.245 ;
        RECT 2390.265 1328.185 2390.665 1328.445 ;
        RECT 2390.805 1328.385 2391.195 1328.445 ;
        RECT 2391.595 1328.425 2391.915 1328.445 ;
        RECT 2391.375 1328.385 2391.915 1328.425 ;
        RECT 2390.805 1328.365 2391.915 1328.385 ;
        RECT 2390.875 1328.245 2391.915 1328.365 ;
        RECT 2390.875 1328.185 2391.195 1328.245 ;
        RECT 2391.375 1328.195 2391.915 1328.245 ;
        RECT 2391.595 1328.185 2391.915 1328.195 ;
        RECT 2392.825 1328.385 2393.145 1328.445 ;
        RECT 2393.295 1328.385 2393.585 1328.425 ;
        RECT 2392.825 1328.245 2393.585 1328.385 ;
        RECT 2392.825 1328.185 2393.145 1328.245 ;
        RECT 2393.295 1328.195 2393.585 1328.245 ;
        RECT 2394.255 1328.385 2394.545 1328.425 ;
        RECT 2394.685 1328.385 2395.005 1328.445 ;
        RECT 2394.255 1328.245 2395.005 1328.385 ;
        RECT 2396.070 1328.320 2398.710 1328.490 ;
        RECT 2398.190 1328.315 2398.710 1328.320 ;
        RECT 2398.360 1328.260 2398.710 1328.315 ;
        RECT 2394.255 1328.195 2394.545 1328.245 ;
        RECT 2394.685 1328.185 2395.005 1328.245 ;
        RECT 2399.350 1328.205 2399.580 1328.230 ;
        RECT 2397.930 1328.120 2398.220 1328.145 ;
        RECT 2399.320 1328.120 2399.610 1328.205 ;
        RECT 2397.930 1327.950 2399.610 1328.120 ;
        RECT 2397.930 1327.915 2398.220 1327.950 ;
        RECT 2382.670 1327.175 2382.960 1327.405 ;
        RECT 2384.460 1327.175 2384.755 1327.435 ;
        RECT 2385.445 1327.175 2385.740 1327.435 ;
        RECT 2397.990 1327.405 2398.160 1327.915 ;
        RECT 2399.320 1327.900 2399.610 1327.950 ;
        RECT 2399.350 1327.880 2399.580 1327.900 ;
        RECT 2399.780 1327.435 2399.950 1328.535 ;
        RECT 2400.765 1327.435 2400.935 1328.535 ;
        RECT 2402.325 1328.185 2402.645 1328.445 ;
        RECT 2404.185 1328.425 2404.325 1328.845 ;
        RECT 2404.475 1328.945 2404.765 1328.985 ;
        RECT 2404.935 1328.945 2405.255 1329.005 ;
        RECT 2404.475 1328.805 2405.255 1328.945 ;
        RECT 2404.475 1328.755 2404.765 1328.805 ;
        RECT 2404.935 1328.745 2405.255 1328.805 ;
        RECT 2405.915 1328.755 2406.205 1328.985 ;
        RECT 2406.065 1328.505 2406.205 1328.755 ;
        RECT 2406.375 1328.745 2406.695 1329.005 ;
        RECT 2407.425 1328.805 2407.565 1329.445 ;
        RECT 2409.275 1329.505 2409.565 1329.545 ;
        RECT 2419.015 1329.505 2419.305 1329.545 ;
        RECT 2409.275 1329.365 2409.845 1329.505 ;
        RECT 2407.905 1329.285 2409.005 1329.365 ;
        RECT 2409.275 1329.315 2409.565 1329.365 ;
        RECT 2407.715 1329.265 2409.005 1329.285 ;
        RECT 2409.705 1329.265 2409.965 1329.365 ;
        RECT 2407.715 1329.225 2409.085 1329.265 ;
        RECT 2409.705 1329.225 2410.045 1329.265 ;
        RECT 2407.715 1329.035 2408.125 1329.225 ;
        RECT 2408.795 1329.035 2409.085 1329.225 ;
        RECT 2409.755 1329.035 2410.045 1329.225 ;
        RECT 2407.715 1329.025 2408.035 1329.035 ;
        RECT 2408.315 1328.805 2408.605 1328.985 ;
        RECT 2407.425 1328.755 2408.605 1328.805 ;
        RECT 2407.425 1328.705 2408.525 1328.755 ;
        RECT 2409.255 1328.745 2409.575 1329.005 ;
        RECT 2411.240 1328.995 2411.580 1329.345 ;
        RECT 2419.015 1329.315 2419.465 1329.505 ;
        RECT 2418.275 1329.025 2418.595 1329.285 ;
        RECT 2407.355 1328.665 2408.525 1328.705 ;
        RECT 2406.065 1328.445 2406.365 1328.505 ;
        RECT 2407.355 1328.455 2407.645 1328.665 ;
        RECT 2411.330 1328.490 2411.500 1328.995 ;
        RECT 2412.845 1328.875 2413.165 1328.980 ;
        RECT 2412.820 1328.860 2413.165 1328.875 ;
        RECT 2412.810 1328.845 2413.165 1328.860 ;
        RECT 2412.645 1328.675 2413.165 1328.845 ;
        RECT 2412.820 1328.660 2413.165 1328.675 ;
        RECT 2412.820 1328.645 2413.110 1328.660 ;
        RECT 2413.620 1328.490 2413.970 1328.610 ;
        RECT 2414.980 1328.540 2415.270 1328.775 ;
        RECT 2415.965 1328.540 2416.255 1328.775 ;
        RECT 2418.755 1328.745 2419.075 1329.005 ;
        RECT 2419.325 1328.985 2419.465 1329.315 ;
        RECT 2419.955 1329.315 2420.505 1329.545 ;
        RECT 2420.645 1329.445 2422.825 1329.585 ;
        RECT 2435.215 1329.545 2435.535 1329.565 ;
        RECT 2420.645 1329.365 2421.945 1329.445 ;
        RECT 2419.955 1329.305 2420.275 1329.315 ;
        RECT 2420.645 1329.085 2420.985 1329.365 ;
        RECT 2421.655 1329.315 2421.945 1329.365 ;
        RECT 2420.695 1329.035 2420.985 1329.085 ;
        RECT 2422.115 1329.025 2422.435 1329.285 ;
        RECT 2419.325 1328.845 2419.585 1328.985 ;
        RECT 2414.980 1328.535 2415.210 1328.540 ;
        RECT 2415.965 1328.535 2416.195 1328.540 ;
        RECT 2404.185 1328.385 2404.525 1328.425 ;
        RECT 2405.055 1328.385 2405.375 1328.445 ;
        RECT 2404.185 1328.245 2405.375 1328.385 ;
        RECT 2404.235 1328.195 2404.525 1328.245 ;
        RECT 2405.055 1328.185 2405.375 1328.245 ;
        RECT 2405.525 1328.185 2405.925 1328.445 ;
        RECT 2406.065 1328.385 2406.455 1328.445 ;
        RECT 2406.855 1328.425 2407.175 1328.445 ;
        RECT 2406.635 1328.385 2407.175 1328.425 ;
        RECT 2406.065 1328.365 2407.175 1328.385 ;
        RECT 2406.135 1328.245 2407.175 1328.365 ;
        RECT 2406.135 1328.185 2406.455 1328.245 ;
        RECT 2406.635 1328.195 2407.175 1328.245 ;
        RECT 2406.855 1328.185 2407.175 1328.195 ;
        RECT 2408.085 1328.385 2408.405 1328.445 ;
        RECT 2408.555 1328.385 2408.845 1328.425 ;
        RECT 2408.085 1328.245 2408.845 1328.385 ;
        RECT 2408.085 1328.185 2408.405 1328.245 ;
        RECT 2408.555 1328.195 2408.845 1328.245 ;
        RECT 2409.515 1328.385 2409.805 1328.425 ;
        RECT 2409.945 1328.385 2410.265 1328.445 ;
        RECT 2409.515 1328.245 2410.265 1328.385 ;
        RECT 2411.330 1328.320 2413.970 1328.490 ;
        RECT 2413.450 1328.315 2413.970 1328.320 ;
        RECT 2413.620 1328.260 2413.970 1328.315 ;
        RECT 2409.515 1328.195 2409.805 1328.245 ;
        RECT 2409.945 1328.185 2410.265 1328.245 ;
        RECT 2414.610 1328.205 2414.840 1328.230 ;
        RECT 2413.190 1328.120 2413.480 1328.145 ;
        RECT 2414.580 1328.120 2414.870 1328.205 ;
        RECT 2413.190 1327.950 2414.870 1328.120 ;
        RECT 2413.190 1327.915 2413.480 1327.950 ;
        RECT 2397.930 1327.175 2398.220 1327.405 ;
        RECT 2399.720 1327.175 2400.015 1327.435 ;
        RECT 2400.705 1327.175 2401.130 1327.435 ;
        RECT 2413.250 1327.405 2413.420 1327.915 ;
        RECT 2414.580 1327.900 2414.870 1327.950 ;
        RECT 2414.610 1327.880 2414.840 1327.900 ;
        RECT 2415.040 1327.435 2415.210 1328.535 ;
        RECT 2416.025 1327.435 2416.195 1328.535 ;
        RECT 2417.585 1328.185 2417.905 1328.445 ;
        RECT 2419.445 1328.425 2419.585 1328.845 ;
        RECT 2419.735 1328.945 2420.025 1328.985 ;
        RECT 2420.195 1328.945 2420.515 1329.005 ;
        RECT 2419.735 1328.805 2420.515 1328.945 ;
        RECT 2419.735 1328.755 2420.025 1328.805 ;
        RECT 2420.195 1328.745 2420.515 1328.805 ;
        RECT 2421.175 1328.755 2421.465 1328.985 ;
        RECT 2421.325 1328.505 2421.465 1328.755 ;
        RECT 2421.635 1328.745 2421.955 1329.005 ;
        RECT 2422.685 1328.805 2422.825 1329.445 ;
        RECT 2424.535 1329.505 2424.825 1329.545 ;
        RECT 2434.275 1329.505 2434.565 1329.545 ;
        RECT 2424.535 1329.365 2425.105 1329.505 ;
        RECT 2423.165 1329.285 2424.265 1329.365 ;
        RECT 2424.535 1329.315 2424.825 1329.365 ;
        RECT 2422.975 1329.265 2424.265 1329.285 ;
        RECT 2424.965 1329.265 2425.225 1329.365 ;
        RECT 2422.975 1329.225 2424.345 1329.265 ;
        RECT 2424.965 1329.225 2425.305 1329.265 ;
        RECT 2422.975 1329.035 2423.385 1329.225 ;
        RECT 2424.055 1329.035 2424.345 1329.225 ;
        RECT 2425.015 1329.035 2425.305 1329.225 ;
        RECT 2422.975 1329.025 2423.295 1329.035 ;
        RECT 2423.575 1328.805 2423.865 1328.985 ;
        RECT 2422.685 1328.755 2423.865 1328.805 ;
        RECT 2422.685 1328.705 2423.785 1328.755 ;
        RECT 2424.515 1328.745 2424.835 1329.005 ;
        RECT 2426.500 1328.995 2426.840 1329.345 ;
        RECT 2434.275 1329.315 2434.725 1329.505 ;
        RECT 2433.535 1329.025 2433.855 1329.285 ;
        RECT 2422.615 1328.665 2423.785 1328.705 ;
        RECT 2421.325 1328.445 2421.625 1328.505 ;
        RECT 2422.615 1328.455 2422.905 1328.665 ;
        RECT 2426.590 1328.490 2426.760 1328.995 ;
        RECT 2428.105 1328.875 2428.425 1328.980 ;
        RECT 2428.080 1328.860 2428.425 1328.875 ;
        RECT 2428.070 1328.845 2428.425 1328.860 ;
        RECT 2427.905 1328.675 2428.425 1328.845 ;
        RECT 2428.080 1328.660 2428.425 1328.675 ;
        RECT 2428.080 1328.645 2428.370 1328.660 ;
        RECT 2428.880 1328.490 2429.230 1328.610 ;
        RECT 2430.240 1328.540 2430.530 1328.775 ;
        RECT 2431.225 1328.540 2431.515 1328.775 ;
        RECT 2434.015 1328.745 2434.335 1329.005 ;
        RECT 2434.585 1328.985 2434.725 1329.315 ;
        RECT 2435.215 1329.315 2435.765 1329.545 ;
        RECT 2435.905 1329.445 2438.085 1329.585 ;
        RECT 2435.905 1329.365 2437.205 1329.445 ;
        RECT 2435.215 1329.305 2435.535 1329.315 ;
        RECT 2435.905 1329.085 2436.245 1329.365 ;
        RECT 2436.915 1329.315 2437.205 1329.365 ;
        RECT 2435.955 1329.035 2436.245 1329.085 ;
        RECT 2437.375 1329.025 2437.695 1329.285 ;
        RECT 2434.585 1328.845 2434.845 1328.985 ;
        RECT 2430.240 1328.535 2430.470 1328.540 ;
        RECT 2431.225 1328.535 2431.455 1328.540 ;
        RECT 2419.445 1328.385 2419.785 1328.425 ;
        RECT 2420.315 1328.385 2420.635 1328.445 ;
        RECT 2419.445 1328.245 2420.635 1328.385 ;
        RECT 2419.495 1328.195 2419.785 1328.245 ;
        RECT 2420.315 1328.185 2420.635 1328.245 ;
        RECT 2420.785 1328.185 2421.185 1328.445 ;
        RECT 2421.325 1328.385 2421.715 1328.445 ;
        RECT 2422.115 1328.425 2422.435 1328.445 ;
        RECT 2421.895 1328.385 2422.435 1328.425 ;
        RECT 2421.325 1328.365 2422.435 1328.385 ;
        RECT 2421.395 1328.245 2422.435 1328.365 ;
        RECT 2421.395 1328.185 2421.715 1328.245 ;
        RECT 2421.895 1328.195 2422.435 1328.245 ;
        RECT 2422.115 1328.185 2422.435 1328.195 ;
        RECT 2423.345 1328.385 2423.665 1328.445 ;
        RECT 2423.815 1328.385 2424.105 1328.425 ;
        RECT 2423.345 1328.245 2424.105 1328.385 ;
        RECT 2423.345 1328.185 2423.665 1328.245 ;
        RECT 2423.815 1328.195 2424.105 1328.245 ;
        RECT 2424.775 1328.385 2425.065 1328.425 ;
        RECT 2425.205 1328.385 2425.525 1328.445 ;
        RECT 2424.775 1328.245 2425.525 1328.385 ;
        RECT 2426.590 1328.320 2429.230 1328.490 ;
        RECT 2428.710 1328.315 2429.230 1328.320 ;
        RECT 2428.880 1328.260 2429.230 1328.315 ;
        RECT 2424.775 1328.195 2425.065 1328.245 ;
        RECT 2425.205 1328.185 2425.525 1328.245 ;
        RECT 2429.870 1328.205 2430.100 1328.230 ;
        RECT 2428.450 1328.120 2428.740 1328.145 ;
        RECT 2429.840 1328.120 2430.130 1328.205 ;
        RECT 2428.450 1327.950 2430.130 1328.120 ;
        RECT 2428.450 1327.915 2428.740 1327.950 ;
        RECT 2413.190 1327.175 2413.480 1327.405 ;
        RECT 2414.980 1327.175 2415.275 1327.435 ;
        RECT 2415.965 1327.175 2416.310 1327.435 ;
        RECT 2428.510 1327.405 2428.680 1327.915 ;
        RECT 2429.840 1327.900 2430.130 1327.950 ;
        RECT 2429.870 1327.880 2430.100 1327.900 ;
        RECT 2430.300 1327.435 2430.470 1328.535 ;
        RECT 2431.285 1327.435 2431.455 1328.535 ;
        RECT 2432.845 1328.185 2433.165 1328.445 ;
        RECT 2434.705 1328.425 2434.845 1328.845 ;
        RECT 2434.995 1328.945 2435.285 1328.985 ;
        RECT 2435.455 1328.945 2435.775 1329.005 ;
        RECT 2434.995 1328.805 2435.775 1328.945 ;
        RECT 2434.995 1328.755 2435.285 1328.805 ;
        RECT 2435.455 1328.745 2435.775 1328.805 ;
        RECT 2436.435 1328.755 2436.725 1328.985 ;
        RECT 2436.585 1328.505 2436.725 1328.755 ;
        RECT 2436.895 1328.745 2437.215 1329.005 ;
        RECT 2437.945 1328.805 2438.085 1329.445 ;
        RECT 2439.795 1329.505 2440.085 1329.545 ;
        RECT 2439.795 1329.365 2440.365 1329.505 ;
        RECT 2438.425 1329.285 2439.525 1329.365 ;
        RECT 2439.795 1329.315 2440.085 1329.365 ;
        RECT 2438.235 1329.265 2439.525 1329.285 ;
        RECT 2440.225 1329.265 2440.485 1329.365 ;
        RECT 2438.235 1329.225 2439.605 1329.265 ;
        RECT 2440.225 1329.225 2440.565 1329.265 ;
        RECT 2438.235 1329.035 2438.645 1329.225 ;
        RECT 2439.315 1329.035 2439.605 1329.225 ;
        RECT 2440.275 1329.035 2440.565 1329.225 ;
        RECT 2438.235 1329.025 2438.555 1329.035 ;
        RECT 2438.835 1328.805 2439.125 1328.985 ;
        RECT 2437.945 1328.755 2439.125 1328.805 ;
        RECT 2437.945 1328.705 2439.045 1328.755 ;
        RECT 2439.775 1328.745 2440.095 1329.005 ;
        RECT 2441.760 1328.995 2442.100 1329.345 ;
        RECT 2437.875 1328.665 2439.045 1328.705 ;
        RECT 2436.585 1328.445 2436.885 1328.505 ;
        RECT 2437.875 1328.455 2438.165 1328.665 ;
        RECT 2441.850 1328.490 2442.020 1328.995 ;
        RECT 2443.365 1328.875 2443.685 1328.980 ;
        RECT 2443.340 1328.860 2443.685 1328.875 ;
        RECT 2443.330 1328.845 2443.685 1328.860 ;
        RECT 2443.165 1328.675 2443.685 1328.845 ;
        RECT 2446.440 1328.775 2446.580 1329.840 ;
        RECT 2459.690 1329.780 2460.010 1329.840 ;
        RECT 2443.340 1328.660 2443.685 1328.675 ;
        RECT 2443.340 1328.645 2443.630 1328.660 ;
        RECT 2444.140 1328.490 2444.490 1328.610 ;
        RECT 2445.500 1328.540 2445.790 1328.775 ;
        RECT 2446.440 1328.655 2446.775 1328.775 ;
        RECT 2446.485 1328.540 2446.775 1328.655 ;
        RECT 2445.500 1328.535 2445.730 1328.540 ;
        RECT 2446.485 1328.535 2446.715 1328.540 ;
        RECT 2434.705 1328.385 2435.045 1328.425 ;
        RECT 2435.575 1328.385 2435.895 1328.445 ;
        RECT 2434.705 1328.245 2435.895 1328.385 ;
        RECT 2434.755 1328.195 2435.045 1328.245 ;
        RECT 2435.575 1328.185 2435.895 1328.245 ;
        RECT 2436.045 1328.185 2436.445 1328.445 ;
        RECT 2436.585 1328.385 2436.975 1328.445 ;
        RECT 2437.375 1328.425 2437.695 1328.445 ;
        RECT 2437.155 1328.385 2437.695 1328.425 ;
        RECT 2436.585 1328.365 2437.695 1328.385 ;
        RECT 2436.655 1328.245 2437.695 1328.365 ;
        RECT 2436.655 1328.185 2436.975 1328.245 ;
        RECT 2437.155 1328.195 2437.695 1328.245 ;
        RECT 2437.375 1328.185 2437.695 1328.195 ;
        RECT 2438.605 1328.385 2438.925 1328.445 ;
        RECT 2439.075 1328.385 2439.365 1328.425 ;
        RECT 2438.605 1328.245 2439.365 1328.385 ;
        RECT 2438.605 1328.185 2438.925 1328.245 ;
        RECT 2439.075 1328.195 2439.365 1328.245 ;
        RECT 2440.035 1328.385 2440.325 1328.425 ;
        RECT 2440.465 1328.385 2440.785 1328.445 ;
        RECT 2440.035 1328.245 2440.785 1328.385 ;
        RECT 2441.850 1328.320 2444.490 1328.490 ;
        RECT 2443.970 1328.315 2444.490 1328.320 ;
        RECT 2444.140 1328.260 2444.490 1328.315 ;
        RECT 2440.035 1328.195 2440.325 1328.245 ;
        RECT 2440.465 1328.185 2440.785 1328.245 ;
        RECT 2445.130 1328.205 2445.360 1328.230 ;
        RECT 2443.710 1328.120 2444.000 1328.145 ;
        RECT 2445.100 1328.120 2445.390 1328.205 ;
        RECT 2443.710 1327.950 2445.390 1328.120 ;
        RECT 2443.710 1327.915 2444.000 1327.950 ;
        RECT 2428.450 1327.175 2428.740 1327.405 ;
        RECT 2430.240 1327.175 2430.535 1327.435 ;
        RECT 2431.170 1327.175 2431.520 1327.435 ;
        RECT 2443.770 1327.405 2443.940 1327.915 ;
        RECT 2445.100 1327.900 2445.390 1327.950 ;
        RECT 2445.130 1327.880 2445.360 1327.900 ;
        RECT 2445.560 1327.435 2445.730 1328.535 ;
        RECT 2446.545 1327.435 2446.715 1328.535 ;
        RECT 2443.710 1327.175 2444.000 1327.405 ;
        RECT 2445.500 1327.175 2445.795 1327.435 ;
        RECT 2446.485 1327.175 2446.780 1327.435 ;
        RECT 2473.580 1317.940 2474.640 1318.080 ;
        RECT 2385.630 1317.540 2385.950 1317.800 ;
        RECT 2400.810 1317.740 2401.130 1317.800 ;
        RECT 2400.810 1317.540 2401.270 1317.740 ;
        RECT 2415.990 1317.540 2416.310 1317.800 ;
        RECT 2431.170 1317.740 2431.490 1317.800 ;
        RECT 2473.580 1317.740 2473.720 1317.940 ;
        RECT 2431.170 1317.600 2473.720 1317.740 ;
        RECT 2474.500 1317.740 2474.640 1317.940 ;
        RECT 2475.330 1317.740 2475.650 1317.800 ;
        RECT 2680.950 1317.740 2681.270 1317.800 ;
        RECT 2474.500 1317.600 2475.100 1317.740 ;
        RECT 2431.170 1317.540 2431.490 1317.600 ;
        RECT 2385.720 1316.720 2385.860 1317.540 ;
        RECT 2401.130 1317.060 2401.270 1317.540 ;
        RECT 2416.080 1317.400 2416.220 1317.540 ;
        RECT 2473.950 1317.400 2474.270 1317.460 ;
        RECT 2416.080 1317.260 2474.270 1317.400 ;
        RECT 2474.960 1317.400 2475.100 1317.600 ;
        RECT 2475.330 1317.600 2681.270 1317.740 ;
        RECT 2475.330 1317.540 2475.650 1317.600 ;
        RECT 2680.950 1317.540 2681.270 1317.600 ;
        RECT 2681.870 1317.400 2682.190 1317.460 ;
        RECT 2474.960 1317.260 2682.190 1317.400 ;
        RECT 2473.950 1317.200 2474.270 1317.260 ;
        RECT 2681.870 1317.200 2682.190 1317.260 ;
        RECT 2597.690 1317.060 2598.010 1317.120 ;
        RECT 2401.130 1316.920 2598.010 1317.060 ;
        RECT 2597.690 1316.860 2598.010 1316.920 ;
        RECT 2514.890 1316.720 2515.210 1316.780 ;
        RECT 2385.720 1316.580 2515.210 1316.720 ;
        RECT 2514.890 1316.520 2515.210 1316.580 ;
      LAYER met2 ;
        RECT 2360.765 2255.285 2443.355 2255.290 ;
        RECT 2359.230 2255.120 2443.355 2255.285 ;
        RECT 2359.230 2255.115 2360.765 2255.120 ;
        RECT 2359.230 2253.875 2359.400 2255.115 ;
        RECT 2443.185 2254.910 2443.355 2255.120 ;
        RECT 2363.325 2254.720 2373.505 2254.890 ;
        RECT 2359.550 2254.510 2359.830 2254.615 ;
        RECT 2359.550 2254.340 2360.715 2254.510 ;
        RECT 2359.550 2254.275 2359.830 2254.340 ;
        RECT 2360.545 2254.145 2360.715 2254.340 ;
        RECT 2362.740 2254.305 2363.110 2254.675 ;
        RECT 2363.325 2254.225 2363.495 2254.720 ;
        RECT 2360.545 2254.140 2360.865 2254.145 ;
        RECT 2363.270 2254.140 2363.550 2254.225 ;
        RECT 2360.545 2253.970 2363.550 2254.140 ;
        RECT 2363.270 2253.885 2363.550 2253.970 ;
        RECT 2373.345 2254.200 2373.505 2254.720 ;
        RECT 2379.910 2254.720 2390.090 2254.890 ;
        RECT 2379.325 2254.305 2379.695 2254.675 ;
        RECT 2374.460 2254.200 2374.785 2254.265 ;
        RECT 2373.345 2254.030 2374.785 2254.200 ;
        RECT 2359.175 2253.535 2359.455 2253.875 ;
        RECT 2367.590 2252.415 2367.870 2252.440 ;
        RECT 2367.590 2252.095 2367.880 2252.415 ;
        RECT 2367.590 2252.065 2367.870 2252.095 ;
        RECT 2368.640 2252.065 2368.920 2252.440 ;
        RECT 2370.000 2252.325 2370.260 2252.415 ;
        RECT 2369.380 2252.185 2370.260 2252.325 ;
        RECT 2367.960 2251.045 2368.240 2251.420 ;
        RECT 2367.280 2248.655 2367.560 2249.035 ;
        RECT 2368.020 2249.015 2368.160 2251.045 ;
        RECT 2368.700 2250.285 2368.840 2252.065 ;
        RECT 2369.380 2250.400 2369.520 2252.185 ;
        RECT 2370.000 2252.095 2370.260 2252.185 ;
        RECT 2371.020 2251.075 2371.280 2251.395 ;
        RECT 2368.700 2250.145 2369.180 2250.285 ;
        RECT 2368.620 2249.345 2368.900 2249.720 ;
        RECT 2367.960 2248.695 2368.220 2249.015 ;
        RECT 2369.040 2248.695 2369.180 2250.145 ;
        RECT 2369.320 2250.025 2369.600 2250.400 ;
        RECT 2369.320 2249.005 2369.600 2249.380 ;
        RECT 2371.080 2249.355 2371.220 2251.075 ;
        RECT 2371.405 2249.695 2371.730 2249.805 ;
        RECT 2371.405 2249.510 2372.235 2249.695 ;
        RECT 2371.405 2249.480 2371.730 2249.510 ;
        RECT 2371.020 2249.035 2371.280 2249.355 ;
        RECT 2368.980 2248.355 2369.240 2248.695 ;
        RECT 2372.065 2248.615 2372.235 2249.510 ;
        RECT 2373.345 2248.860 2373.505 2254.030 ;
        RECT 2374.460 2253.940 2374.785 2254.030 ;
        RECT 2376.850 2254.145 2377.175 2254.270 ;
        RECT 2379.910 2254.225 2380.080 2254.720 ;
        RECT 2376.850 2254.140 2377.685 2254.145 ;
        RECT 2379.855 2254.140 2380.135 2254.225 ;
        RECT 2376.850 2253.975 2380.135 2254.140 ;
        RECT 2376.850 2253.945 2377.175 2253.975 ;
        RECT 2377.685 2253.970 2380.135 2253.975 ;
        RECT 2373.660 2253.565 2373.980 2253.890 ;
        RECT 2379.855 2253.885 2380.135 2253.970 ;
        RECT 2389.930 2254.200 2390.090 2254.720 ;
        RECT 2396.495 2254.720 2406.675 2254.890 ;
        RECT 2395.910 2254.280 2396.280 2254.675 ;
        RECT 2391.045 2254.200 2391.370 2254.265 ;
        RECT 2389.930 2254.030 2391.370 2254.200 ;
        RECT 2373.690 2253.330 2373.860 2253.565 ;
        RECT 2373.690 2253.155 2373.865 2253.330 ;
        RECT 2373.690 2252.980 2374.665 2253.155 ;
        RECT 2373.660 2248.860 2373.980 2248.980 ;
        RECT 2373.345 2248.690 2373.980 2248.860 ;
        RECT 2373.660 2248.660 2373.980 2248.690 ;
        RECT 2371.990 2248.290 2372.315 2248.615 ;
        RECT 2374.490 2248.610 2374.665 2252.980 ;
        RECT 2384.175 2252.415 2384.455 2252.440 ;
        RECT 2384.175 2252.095 2384.465 2252.415 ;
        RECT 2384.175 2252.065 2384.455 2252.095 ;
        RECT 2385.225 2252.065 2385.505 2252.440 ;
        RECT 2386.585 2252.325 2386.845 2252.415 ;
        RECT 2385.965 2252.185 2386.845 2252.325 ;
        RECT 2384.545 2251.045 2384.825 2251.420 ;
        RECT 2383.865 2248.655 2384.145 2249.035 ;
        RECT 2384.605 2249.015 2384.745 2251.045 ;
        RECT 2385.285 2250.285 2385.425 2252.065 ;
        RECT 2385.965 2250.400 2386.105 2252.185 ;
        RECT 2386.585 2252.095 2386.845 2252.185 ;
        RECT 2387.605 2251.075 2387.865 2251.395 ;
        RECT 2385.285 2250.145 2385.765 2250.285 ;
        RECT 2385.205 2249.345 2385.485 2249.720 ;
        RECT 2384.545 2248.695 2384.805 2249.015 ;
        RECT 2385.625 2248.695 2385.765 2250.145 ;
        RECT 2385.905 2250.025 2386.185 2250.400 ;
        RECT 2385.905 2249.005 2386.185 2249.380 ;
        RECT 2387.665 2249.355 2387.805 2251.075 ;
        RECT 2387.990 2249.695 2388.315 2249.805 ;
        RECT 2387.990 2249.510 2388.820 2249.695 ;
        RECT 2387.990 2249.480 2388.315 2249.510 ;
        RECT 2387.605 2249.035 2387.865 2249.355 ;
        RECT 2374.435 2248.260 2374.785 2248.610 ;
        RECT 2385.565 2248.355 2385.825 2248.695 ;
        RECT 2388.650 2248.615 2388.820 2249.510 ;
        RECT 2389.930 2248.860 2390.090 2254.030 ;
        RECT 2391.045 2253.940 2391.370 2254.030 ;
        RECT 2393.435 2254.145 2393.760 2254.270 ;
        RECT 2396.495 2254.225 2396.665 2254.720 ;
        RECT 2393.435 2254.140 2394.050 2254.145 ;
        RECT 2396.440 2254.140 2396.720 2254.225 ;
        RECT 2393.435 2253.975 2396.720 2254.140 ;
        RECT 2393.435 2253.945 2393.760 2253.975 ;
        RECT 2394.050 2253.970 2396.720 2253.975 ;
        RECT 2390.245 2253.565 2390.565 2253.890 ;
        RECT 2396.440 2253.885 2396.720 2253.970 ;
        RECT 2406.515 2254.200 2406.675 2254.720 ;
        RECT 2413.080 2254.720 2423.260 2254.890 ;
        RECT 2412.495 2254.280 2412.865 2254.675 ;
        RECT 2407.630 2254.200 2407.955 2254.265 ;
        RECT 2406.515 2254.030 2407.955 2254.200 ;
        RECT 2390.275 2253.330 2390.445 2253.565 ;
        RECT 2390.275 2253.155 2390.450 2253.330 ;
        RECT 2390.275 2252.980 2391.250 2253.155 ;
        RECT 2390.245 2248.860 2390.565 2248.980 ;
        RECT 2389.930 2248.690 2390.565 2248.860 ;
        RECT 2390.245 2248.660 2390.565 2248.690 ;
        RECT 2388.575 2248.290 2388.900 2248.615 ;
        RECT 2391.075 2248.610 2391.250 2252.980 ;
        RECT 2400.760 2252.415 2401.040 2252.440 ;
        RECT 2400.760 2252.095 2401.050 2252.415 ;
        RECT 2400.760 2252.065 2401.040 2252.095 ;
        RECT 2401.810 2252.065 2402.090 2252.440 ;
        RECT 2403.170 2252.325 2403.430 2252.415 ;
        RECT 2402.550 2252.185 2403.430 2252.325 ;
        RECT 2401.130 2251.045 2401.410 2251.420 ;
        RECT 2400.450 2248.655 2400.730 2249.035 ;
        RECT 2401.190 2249.015 2401.330 2251.045 ;
        RECT 2401.870 2250.285 2402.010 2252.065 ;
        RECT 2402.550 2250.400 2402.690 2252.185 ;
        RECT 2403.170 2252.095 2403.430 2252.185 ;
        RECT 2404.190 2251.075 2404.450 2251.395 ;
        RECT 2401.870 2250.145 2402.350 2250.285 ;
        RECT 2401.790 2249.345 2402.070 2249.720 ;
        RECT 2401.130 2248.695 2401.390 2249.015 ;
        RECT 2402.210 2248.695 2402.350 2250.145 ;
        RECT 2402.490 2250.025 2402.770 2250.400 ;
        RECT 2402.490 2249.005 2402.770 2249.380 ;
        RECT 2404.250 2249.355 2404.390 2251.075 ;
        RECT 2404.575 2249.695 2404.900 2249.805 ;
        RECT 2404.575 2249.510 2405.405 2249.695 ;
        RECT 2404.575 2249.480 2404.900 2249.510 ;
        RECT 2404.190 2249.035 2404.450 2249.355 ;
        RECT 2391.020 2248.260 2391.370 2248.610 ;
        RECT 2402.150 2248.355 2402.410 2248.695 ;
        RECT 2405.235 2248.615 2405.405 2249.510 ;
        RECT 2406.515 2248.860 2406.675 2254.030 ;
        RECT 2407.630 2253.940 2407.955 2254.030 ;
        RECT 2410.020 2254.145 2410.345 2254.270 ;
        RECT 2413.080 2254.225 2413.250 2254.720 ;
        RECT 2410.020 2254.140 2410.865 2254.145 ;
        RECT 2413.025 2254.140 2413.305 2254.225 ;
        RECT 2410.020 2253.975 2413.305 2254.140 ;
        RECT 2410.020 2253.945 2410.345 2253.975 ;
        RECT 2410.865 2253.970 2413.305 2253.975 ;
        RECT 2406.830 2253.565 2407.150 2253.890 ;
        RECT 2413.025 2253.885 2413.305 2253.970 ;
        RECT 2423.100 2254.200 2423.260 2254.720 ;
        RECT 2429.660 2254.720 2439.840 2254.890 ;
        RECT 2429.075 2254.650 2429.445 2254.675 ;
        RECT 2429.075 2254.305 2429.450 2254.650 ;
        RECT 2429.080 2254.280 2429.450 2254.305 ;
        RECT 2424.215 2254.200 2424.540 2254.265 ;
        RECT 2423.100 2254.030 2424.540 2254.200 ;
        RECT 2406.860 2253.330 2407.030 2253.565 ;
        RECT 2406.860 2253.155 2407.035 2253.330 ;
        RECT 2406.860 2252.980 2407.835 2253.155 ;
        RECT 2406.830 2248.860 2407.150 2248.980 ;
        RECT 2406.515 2248.690 2407.150 2248.860 ;
        RECT 2406.830 2248.660 2407.150 2248.690 ;
        RECT 2405.160 2248.290 2405.485 2248.615 ;
        RECT 2407.660 2248.610 2407.835 2252.980 ;
        RECT 2417.345 2252.415 2417.625 2252.440 ;
        RECT 2417.345 2252.095 2417.635 2252.415 ;
        RECT 2417.345 2252.065 2417.625 2252.095 ;
        RECT 2418.395 2252.065 2418.675 2252.440 ;
        RECT 2419.755 2252.325 2420.015 2252.415 ;
        RECT 2419.135 2252.185 2420.015 2252.325 ;
        RECT 2417.715 2251.045 2417.995 2251.420 ;
        RECT 2417.035 2248.655 2417.315 2249.035 ;
        RECT 2417.775 2249.015 2417.915 2251.045 ;
        RECT 2418.455 2250.285 2418.595 2252.065 ;
        RECT 2419.135 2250.400 2419.275 2252.185 ;
        RECT 2419.755 2252.095 2420.015 2252.185 ;
        RECT 2420.775 2251.075 2421.035 2251.395 ;
        RECT 2418.455 2250.145 2418.935 2250.285 ;
        RECT 2418.375 2249.345 2418.655 2249.720 ;
        RECT 2417.715 2248.695 2417.975 2249.015 ;
        RECT 2418.795 2248.695 2418.935 2250.145 ;
        RECT 2419.075 2250.025 2419.355 2250.400 ;
        RECT 2419.075 2249.005 2419.355 2249.380 ;
        RECT 2420.835 2249.355 2420.975 2251.075 ;
        RECT 2421.160 2249.695 2421.485 2249.805 ;
        RECT 2421.160 2249.510 2421.990 2249.695 ;
        RECT 2421.160 2249.480 2421.485 2249.510 ;
        RECT 2420.775 2249.035 2421.035 2249.355 ;
        RECT 2407.605 2248.260 2407.955 2248.610 ;
        RECT 2418.735 2248.355 2418.995 2248.695 ;
        RECT 2421.820 2248.615 2421.990 2249.510 ;
        RECT 2423.100 2248.860 2423.260 2254.030 ;
        RECT 2424.215 2253.940 2424.540 2254.030 ;
        RECT 2426.605 2254.145 2426.930 2254.270 ;
        RECT 2429.660 2254.225 2429.830 2254.720 ;
        RECT 2426.605 2254.140 2427.310 2254.145 ;
        RECT 2429.605 2254.140 2429.885 2254.225 ;
        RECT 2426.605 2253.975 2429.885 2254.140 ;
        RECT 2426.605 2253.945 2426.930 2253.975 ;
        RECT 2427.310 2253.970 2429.885 2253.975 ;
        RECT 2423.415 2253.565 2423.735 2253.890 ;
        RECT 2429.605 2253.885 2429.885 2253.970 ;
        RECT 2439.680 2254.200 2439.840 2254.720 ;
        RECT 2443.150 2254.585 2443.475 2254.910 ;
        RECT 2440.795 2254.200 2441.120 2254.265 ;
        RECT 2439.680 2254.030 2441.120 2254.200 ;
        RECT 2423.445 2253.330 2423.615 2253.565 ;
        RECT 2423.445 2253.155 2423.620 2253.330 ;
        RECT 2423.445 2252.980 2424.420 2253.155 ;
        RECT 2423.415 2248.860 2423.735 2248.980 ;
        RECT 2423.100 2248.690 2423.735 2248.860 ;
        RECT 2423.415 2248.660 2423.735 2248.690 ;
        RECT 2421.745 2248.290 2422.070 2248.615 ;
        RECT 2424.245 2248.610 2424.420 2252.980 ;
        RECT 2433.925 2252.415 2434.205 2252.440 ;
        RECT 2433.925 2252.095 2434.215 2252.415 ;
        RECT 2433.925 2252.065 2434.205 2252.095 ;
        RECT 2434.975 2252.065 2435.255 2252.440 ;
        RECT 2436.335 2252.325 2436.595 2252.415 ;
        RECT 2435.715 2252.185 2436.595 2252.325 ;
        RECT 2434.295 2251.045 2434.575 2251.420 ;
        RECT 2433.615 2248.655 2433.895 2249.035 ;
        RECT 2434.355 2249.015 2434.495 2251.045 ;
        RECT 2435.035 2250.285 2435.175 2252.065 ;
        RECT 2435.715 2250.400 2435.855 2252.185 ;
        RECT 2436.335 2252.095 2436.595 2252.185 ;
        RECT 2437.355 2251.075 2437.615 2251.395 ;
        RECT 2435.035 2250.145 2435.515 2250.285 ;
        RECT 2434.955 2249.345 2435.235 2249.720 ;
        RECT 2434.295 2248.695 2434.555 2249.015 ;
        RECT 2435.375 2248.695 2435.515 2250.145 ;
        RECT 2435.655 2250.025 2435.935 2250.400 ;
        RECT 2435.655 2249.005 2435.935 2249.380 ;
        RECT 2437.415 2249.355 2437.555 2251.075 ;
        RECT 2437.740 2249.695 2438.065 2249.805 ;
        RECT 2437.740 2249.510 2438.570 2249.695 ;
        RECT 2437.740 2249.480 2438.065 2249.510 ;
        RECT 2437.355 2249.035 2437.615 2249.355 ;
        RECT 2424.190 2248.260 2424.540 2248.610 ;
        RECT 2435.315 2248.355 2435.575 2248.695 ;
        RECT 2438.400 2248.615 2438.570 2249.510 ;
        RECT 2439.680 2248.860 2439.840 2254.030 ;
        RECT 2440.795 2253.940 2441.120 2254.030 ;
        RECT 2439.995 2253.565 2440.315 2253.890 ;
        RECT 2440.025 2253.330 2440.195 2253.565 ;
        RECT 2440.025 2253.155 2440.200 2253.330 ;
        RECT 2440.025 2252.980 2441.000 2253.155 ;
        RECT 2439.995 2248.860 2440.315 2248.980 ;
        RECT 2439.680 2248.690 2440.315 2248.860 ;
        RECT 2439.995 2248.660 2440.315 2248.690 ;
        RECT 2438.325 2248.290 2438.650 2248.615 ;
        RECT 2440.825 2248.610 2441.000 2252.980 ;
        RECT 2440.770 2248.260 2441.120 2248.610 ;
        RECT 2376.920 2247.150 2377.180 2247.470 ;
        RECT 2393.480 2247.150 2393.740 2247.470 ;
        RECT 2410.040 2247.150 2410.300 2247.470 ;
        RECT 2426.600 2247.150 2426.860 2247.470 ;
        RECT 2376.980 2228.690 2377.120 2247.150 ;
        RECT 2393.540 2231.410 2393.680 2247.150 ;
        RECT 2393.480 2231.090 2393.740 2231.410 ;
        RECT 2410.100 2229.370 2410.240 2247.150 ;
        RECT 2426.660 2229.370 2426.800 2247.150 ;
        RECT 2459.720 2246.730 2459.980 2247.050 ;
        RECT 2410.040 2229.050 2410.300 2229.370 ;
        RECT 2426.600 2229.050 2426.860 2229.370 ;
        RECT 2376.920 2228.370 2377.180 2228.690 ;
        RECT 2452.820 2214.770 2453.080 2215.090 ;
        RECT 2359.245 2163.065 2446.555 2163.235 ;
        RECT 2359.245 2161.880 2359.415 2163.065 ;
        RECT 2446.385 2162.910 2446.555 2163.065 ;
        RECT 2359.565 2162.515 2359.845 2162.620 ;
        RECT 2359.565 2162.345 2360.775 2162.515 ;
        RECT 2359.565 2162.280 2359.845 2162.345 ;
        RECT 2360.605 2162.140 2360.775 2162.345 ;
        RECT 2362.940 2162.310 2363.310 2162.680 ;
        RECT 2363.465 2162.650 2374.160 2162.820 ;
        RECT 2363.465 2162.170 2363.635 2162.650 ;
        RECT 2374.000 2162.200 2374.160 2162.650 ;
        RECT 2380.160 2162.310 2380.530 2162.680 ;
        RECT 2380.685 2162.650 2391.380 2162.820 ;
        RECT 2375.115 2162.200 2375.440 2162.265 ;
        RECT 2363.415 2162.140 2363.695 2162.170 ;
        RECT 2360.605 2161.970 2363.695 2162.140 ;
        RECT 2359.190 2161.540 2359.470 2161.880 ;
        RECT 2363.415 2161.830 2363.695 2161.970 ;
        RECT 2374.000 2162.030 2375.440 2162.200 ;
        RECT 2367.700 2160.725 2367.980 2161.095 ;
        RECT 2369.070 2161.050 2369.330 2161.095 ;
        RECT 2369.040 2160.805 2369.360 2161.050 ;
        RECT 2369.070 2160.760 2369.330 2160.805 ;
        RECT 2370.770 2160.760 2371.030 2161.095 ;
        RECT 2368.710 2160.065 2368.990 2160.435 ;
        RECT 2369.130 2159.645 2369.270 2160.760 ;
        RECT 2369.750 2160.065 2370.030 2160.435 ;
        RECT 2368.450 2159.505 2369.270 2159.645 ;
        RECT 2365.670 2159.075 2365.930 2159.395 ;
        RECT 2365.730 2157.355 2365.870 2159.075 ;
        RECT 2368.450 2158.800 2368.590 2159.505 ;
        RECT 2370.090 2159.075 2370.350 2159.395 ;
        RECT 2366.340 2158.430 2366.620 2158.800 ;
        RECT 2368.380 2158.430 2368.660 2158.800 ;
        RECT 2365.670 2157.035 2365.930 2157.355 ;
        RECT 2366.410 2157.015 2366.550 2158.430 ;
        RECT 2368.030 2157.690 2368.310 2158.060 ;
        RECT 2368.450 2157.355 2368.590 2158.430 ;
        RECT 2369.400 2158.030 2369.680 2158.400 ;
        RECT 2370.150 2158.375 2370.290 2159.075 ;
        RECT 2370.090 2158.055 2370.350 2158.375 ;
        RECT 2368.390 2157.035 2368.650 2157.355 ;
        RECT 2369.060 2157.350 2369.340 2157.720 ;
        RECT 2370.830 2157.355 2370.970 2160.760 ;
        RECT 2366.350 2156.695 2366.610 2157.015 ;
        RECT 2367.700 2156.500 2367.980 2156.870 ;
        RECT 2369.130 2156.815 2369.305 2157.350 ;
        RECT 2370.770 2157.035 2371.030 2157.355 ;
        RECT 2374.000 2156.860 2374.160 2162.030 ;
        RECT 2375.115 2161.940 2375.440 2162.030 ;
        RECT 2377.505 2162.145 2377.830 2162.270 ;
        RECT 2380.685 2162.170 2380.855 2162.650 ;
        RECT 2391.220 2162.200 2391.380 2162.650 ;
        RECT 2397.380 2162.310 2397.750 2162.680 ;
        RECT 2397.905 2162.650 2408.600 2162.820 ;
        RECT 2392.335 2162.200 2392.660 2162.265 ;
        RECT 2377.505 2162.140 2378.415 2162.145 ;
        RECT 2380.635 2162.140 2380.915 2162.170 ;
        RECT 2377.505 2161.975 2380.915 2162.140 ;
        RECT 2377.505 2161.945 2377.830 2161.975 ;
        RECT 2378.415 2161.970 2380.915 2161.975 ;
        RECT 2374.315 2161.565 2374.635 2161.890 ;
        RECT 2380.635 2161.830 2380.915 2161.970 ;
        RECT 2391.220 2162.030 2392.660 2162.200 ;
        RECT 2374.345 2161.330 2374.515 2161.565 ;
        RECT 2374.345 2161.155 2374.520 2161.330 ;
        RECT 2374.345 2160.980 2375.320 2161.155 ;
        RECT 2374.315 2156.860 2374.635 2156.980 ;
        RECT 2369.130 2156.640 2372.350 2156.815 ;
        RECT 2374.000 2156.690 2374.635 2156.860 ;
        RECT 2374.315 2156.660 2374.635 2156.690 ;
        RECT 2372.175 2156.490 2372.350 2156.640 ;
        RECT 2372.645 2156.490 2372.970 2156.615 ;
        RECT 2375.145 2156.610 2375.320 2160.980 ;
        RECT 2384.920 2160.725 2385.200 2161.095 ;
        RECT 2386.290 2161.050 2386.550 2161.095 ;
        RECT 2386.260 2160.805 2386.580 2161.050 ;
        RECT 2386.290 2160.760 2386.550 2160.805 ;
        RECT 2387.990 2160.760 2388.250 2161.095 ;
        RECT 2385.930 2160.065 2386.210 2160.435 ;
        RECT 2386.350 2159.645 2386.490 2160.760 ;
        RECT 2386.970 2160.065 2387.250 2160.435 ;
        RECT 2385.670 2159.505 2386.490 2159.645 ;
        RECT 2382.890 2159.075 2383.150 2159.395 ;
        RECT 2382.950 2157.355 2383.090 2159.075 ;
        RECT 2385.670 2158.800 2385.810 2159.505 ;
        RECT 2387.310 2159.075 2387.570 2159.395 ;
        RECT 2383.560 2158.430 2383.840 2158.800 ;
        RECT 2385.600 2158.430 2385.880 2158.800 ;
        RECT 2382.890 2157.035 2383.150 2157.355 ;
        RECT 2383.630 2157.015 2383.770 2158.430 ;
        RECT 2385.250 2157.690 2385.530 2158.060 ;
        RECT 2385.670 2157.355 2385.810 2158.430 ;
        RECT 2386.620 2158.030 2386.900 2158.400 ;
        RECT 2387.370 2158.375 2387.510 2159.075 ;
        RECT 2387.310 2158.055 2387.570 2158.375 ;
        RECT 2385.610 2157.035 2385.870 2157.355 ;
        RECT 2386.280 2157.350 2386.560 2157.720 ;
        RECT 2388.050 2157.355 2388.190 2160.760 ;
        RECT 2383.570 2156.695 2383.830 2157.015 ;
        RECT 2375.090 2156.490 2375.440 2156.610 ;
        RECT 2384.920 2156.500 2385.200 2156.870 ;
        RECT 2386.350 2156.815 2386.525 2157.350 ;
        RECT 2387.990 2157.035 2388.250 2157.355 ;
        RECT 2391.220 2156.860 2391.380 2162.030 ;
        RECT 2392.335 2161.940 2392.660 2162.030 ;
        RECT 2394.725 2162.145 2395.050 2162.270 ;
        RECT 2397.905 2162.170 2398.075 2162.650 ;
        RECT 2408.440 2162.200 2408.600 2162.650 ;
        RECT 2414.600 2162.310 2414.970 2162.680 ;
        RECT 2415.125 2162.650 2425.820 2162.820 ;
        RECT 2409.555 2162.200 2409.880 2162.265 ;
        RECT 2394.725 2162.140 2395.650 2162.145 ;
        RECT 2397.855 2162.140 2398.135 2162.170 ;
        RECT 2394.725 2161.975 2398.145 2162.140 ;
        RECT 2394.725 2161.945 2395.050 2161.975 ;
        RECT 2396.675 2161.970 2398.145 2161.975 ;
        RECT 2408.440 2162.030 2409.880 2162.200 ;
        RECT 2391.535 2161.565 2391.855 2161.890 ;
        RECT 2397.855 2161.830 2398.135 2161.970 ;
        RECT 2391.565 2161.330 2391.735 2161.565 ;
        RECT 2391.565 2161.155 2391.740 2161.330 ;
        RECT 2391.565 2160.980 2392.540 2161.155 ;
        RECT 2391.535 2156.860 2391.855 2156.980 ;
        RECT 2386.350 2156.640 2389.570 2156.815 ;
        RECT 2391.220 2156.690 2391.855 2156.860 ;
        RECT 2391.535 2156.660 2391.855 2156.690 ;
        RECT 2372.175 2156.320 2375.440 2156.490 ;
        RECT 2389.395 2156.490 2389.570 2156.640 ;
        RECT 2389.865 2156.490 2390.190 2156.615 ;
        RECT 2392.365 2156.610 2392.540 2160.980 ;
        RECT 2402.140 2160.725 2402.420 2161.095 ;
        RECT 2403.510 2161.050 2403.770 2161.095 ;
        RECT 2403.480 2160.805 2403.800 2161.050 ;
        RECT 2403.510 2160.760 2403.770 2160.805 ;
        RECT 2405.210 2160.760 2405.470 2161.095 ;
        RECT 2403.150 2160.065 2403.430 2160.435 ;
        RECT 2403.570 2159.645 2403.710 2160.760 ;
        RECT 2404.190 2160.065 2404.470 2160.435 ;
        RECT 2402.890 2159.505 2403.710 2159.645 ;
        RECT 2400.110 2159.075 2400.370 2159.395 ;
        RECT 2400.170 2157.355 2400.310 2159.075 ;
        RECT 2402.890 2158.800 2403.030 2159.505 ;
        RECT 2404.530 2159.075 2404.790 2159.395 ;
        RECT 2400.780 2158.430 2401.060 2158.800 ;
        RECT 2402.820 2158.430 2403.100 2158.800 ;
        RECT 2394.860 2156.970 2395.120 2157.290 ;
        RECT 2400.110 2157.035 2400.370 2157.355 ;
        RECT 2400.850 2157.015 2400.990 2158.430 ;
        RECT 2402.470 2157.690 2402.750 2158.060 ;
        RECT 2402.890 2157.355 2403.030 2158.430 ;
        RECT 2403.840 2158.030 2404.120 2158.400 ;
        RECT 2404.590 2158.375 2404.730 2159.075 ;
        RECT 2404.530 2158.055 2404.790 2158.375 ;
        RECT 2402.830 2157.035 2403.090 2157.355 ;
        RECT 2403.500 2157.350 2403.780 2157.720 ;
        RECT 2405.270 2157.355 2405.410 2160.760 ;
        RECT 2392.310 2156.490 2392.660 2156.610 ;
        RECT 2389.395 2156.320 2392.660 2156.490 ;
        RECT 2372.645 2156.290 2372.970 2156.320 ;
        RECT 2375.090 2156.260 2375.440 2156.320 ;
        RECT 2389.865 2156.290 2390.190 2156.320 ;
        RECT 2392.310 2156.260 2392.660 2156.320 ;
        RECT 2377.380 2155.145 2377.640 2155.465 ;
        RECT 2377.440 2145.730 2377.580 2155.145 ;
        RECT 2377.380 2145.410 2377.640 2145.730 ;
        RECT 2394.920 2139.805 2395.060 2156.970 ;
        RECT 2400.790 2156.695 2401.050 2157.015 ;
        RECT 2402.140 2156.500 2402.420 2156.870 ;
        RECT 2403.570 2156.815 2403.745 2157.350 ;
        RECT 2405.210 2157.035 2405.470 2157.355 ;
        RECT 2408.440 2156.860 2408.600 2162.030 ;
        RECT 2409.555 2161.940 2409.880 2162.030 ;
        RECT 2411.945 2162.145 2412.270 2162.270 ;
        RECT 2415.125 2162.170 2415.295 2162.650 ;
        RECT 2425.660 2162.200 2425.820 2162.650 ;
        RECT 2431.820 2162.310 2432.190 2162.680 ;
        RECT 2432.345 2162.650 2443.040 2162.820 ;
        RECT 2426.775 2162.200 2427.100 2162.265 ;
        RECT 2411.945 2162.140 2412.890 2162.145 ;
        RECT 2415.075 2162.140 2415.355 2162.170 ;
        RECT 2411.945 2161.975 2415.355 2162.140 ;
        RECT 2411.945 2161.945 2412.270 2161.975 ;
        RECT 2412.890 2161.970 2415.355 2161.975 ;
        RECT 2408.755 2161.565 2409.075 2161.890 ;
        RECT 2415.075 2161.830 2415.355 2161.970 ;
        RECT 2425.660 2162.030 2427.100 2162.200 ;
        RECT 2408.785 2161.330 2408.955 2161.565 ;
        RECT 2408.785 2161.155 2408.960 2161.330 ;
        RECT 2408.785 2160.980 2409.760 2161.155 ;
        RECT 2408.755 2156.860 2409.075 2156.980 ;
        RECT 2403.570 2156.640 2406.790 2156.815 ;
        RECT 2408.440 2156.690 2409.075 2156.860 ;
        RECT 2408.755 2156.660 2409.075 2156.690 ;
        RECT 2406.615 2156.490 2406.790 2156.640 ;
        RECT 2407.085 2156.490 2407.410 2156.615 ;
        RECT 2409.585 2156.610 2409.760 2160.980 ;
        RECT 2419.360 2160.725 2419.640 2161.095 ;
        RECT 2420.730 2161.050 2420.990 2161.095 ;
        RECT 2420.700 2160.805 2421.020 2161.050 ;
        RECT 2420.730 2160.760 2420.990 2160.805 ;
        RECT 2422.430 2160.760 2422.690 2161.095 ;
        RECT 2420.370 2160.065 2420.650 2160.435 ;
        RECT 2420.790 2159.645 2420.930 2160.760 ;
        RECT 2421.410 2160.065 2421.690 2160.435 ;
        RECT 2420.110 2159.505 2420.930 2159.645 ;
        RECT 2417.330 2159.075 2417.590 2159.395 ;
        RECT 2417.390 2157.355 2417.530 2159.075 ;
        RECT 2420.110 2158.800 2420.250 2159.505 ;
        RECT 2421.750 2159.075 2422.010 2159.395 ;
        RECT 2418.000 2158.430 2418.280 2158.800 ;
        RECT 2420.040 2158.430 2420.320 2158.800 ;
        RECT 2417.330 2157.035 2417.590 2157.355 ;
        RECT 2418.070 2157.015 2418.210 2158.430 ;
        RECT 2419.690 2157.690 2419.970 2158.060 ;
        RECT 2420.110 2157.355 2420.250 2158.430 ;
        RECT 2421.060 2158.030 2421.340 2158.400 ;
        RECT 2421.810 2158.375 2421.950 2159.075 ;
        RECT 2421.750 2158.055 2422.010 2158.375 ;
        RECT 2420.050 2157.035 2420.310 2157.355 ;
        RECT 2420.720 2157.350 2421.000 2157.720 ;
        RECT 2422.490 2157.355 2422.630 2160.760 ;
        RECT 2418.010 2156.695 2418.270 2157.015 ;
        RECT 2409.530 2156.490 2409.880 2156.610 ;
        RECT 2419.360 2156.500 2419.640 2156.870 ;
        RECT 2420.790 2156.815 2420.965 2157.350 ;
        RECT 2422.430 2157.035 2422.690 2157.355 ;
        RECT 2425.660 2156.860 2425.820 2162.030 ;
        RECT 2426.775 2161.940 2427.100 2162.030 ;
        RECT 2429.165 2162.145 2429.490 2162.270 ;
        RECT 2432.345 2162.170 2432.515 2162.650 ;
        RECT 2442.880 2162.200 2443.040 2162.650 ;
        RECT 2446.350 2162.585 2446.675 2162.910 ;
        RECT 2443.995 2162.200 2444.320 2162.265 ;
        RECT 2429.165 2162.140 2430.155 2162.145 ;
        RECT 2432.295 2162.140 2432.575 2162.170 ;
        RECT 2429.165 2161.975 2432.575 2162.140 ;
        RECT 2429.165 2161.945 2429.490 2161.975 ;
        RECT 2430.155 2161.970 2432.575 2161.975 ;
        RECT 2425.975 2161.565 2426.295 2161.890 ;
        RECT 2432.295 2161.830 2432.575 2161.970 ;
        RECT 2442.880 2162.030 2444.320 2162.200 ;
        RECT 2426.005 2161.330 2426.175 2161.565 ;
        RECT 2426.005 2161.155 2426.180 2161.330 ;
        RECT 2426.005 2160.980 2426.980 2161.155 ;
        RECT 2425.975 2156.860 2426.295 2156.980 ;
        RECT 2420.790 2156.640 2424.010 2156.815 ;
        RECT 2425.660 2156.690 2426.295 2156.860 ;
        RECT 2425.975 2156.660 2426.295 2156.690 ;
        RECT 2406.615 2156.320 2409.880 2156.490 ;
        RECT 2423.835 2156.490 2424.010 2156.640 ;
        RECT 2424.305 2156.490 2424.630 2156.615 ;
        RECT 2426.805 2156.610 2426.980 2160.980 ;
        RECT 2436.580 2160.725 2436.860 2161.095 ;
        RECT 2437.950 2161.050 2438.210 2161.095 ;
        RECT 2437.920 2160.805 2438.240 2161.050 ;
        RECT 2437.950 2160.760 2438.210 2160.805 ;
        RECT 2439.650 2160.760 2439.910 2161.095 ;
        RECT 2437.590 2160.065 2437.870 2160.435 ;
        RECT 2438.010 2159.645 2438.150 2160.760 ;
        RECT 2438.630 2160.065 2438.910 2160.435 ;
        RECT 2437.330 2159.505 2438.150 2159.645 ;
        RECT 2434.550 2159.075 2434.810 2159.395 ;
        RECT 2434.610 2157.355 2434.750 2159.075 ;
        RECT 2437.330 2158.800 2437.470 2159.505 ;
        RECT 2438.970 2159.075 2439.230 2159.395 ;
        RECT 2435.220 2158.430 2435.500 2158.800 ;
        RECT 2437.260 2158.430 2437.540 2158.800 ;
        RECT 2428.900 2156.970 2429.160 2157.290 ;
        RECT 2434.550 2157.035 2434.810 2157.355 ;
        RECT 2435.290 2157.015 2435.430 2158.430 ;
        RECT 2436.910 2157.690 2437.190 2158.060 ;
        RECT 2437.330 2157.355 2437.470 2158.430 ;
        RECT 2438.280 2158.030 2438.560 2158.400 ;
        RECT 2439.030 2158.375 2439.170 2159.075 ;
        RECT 2438.970 2158.055 2439.230 2158.375 ;
        RECT 2437.270 2157.035 2437.530 2157.355 ;
        RECT 2437.940 2157.350 2438.220 2157.720 ;
        RECT 2439.710 2157.355 2439.850 2160.760 ;
        RECT 2426.750 2156.490 2427.100 2156.610 ;
        RECT 2423.835 2156.320 2427.100 2156.490 ;
        RECT 2407.085 2156.290 2407.410 2156.320 ;
        RECT 2409.530 2156.260 2409.880 2156.320 ;
        RECT 2424.305 2156.290 2424.630 2156.320 ;
        RECT 2426.750 2156.260 2427.100 2156.320 ;
        RECT 2411.880 2155.145 2412.140 2155.465 ;
        RECT 2394.850 2139.435 2395.130 2139.805 ;
        RECT 2411.940 2139.270 2412.080 2155.145 ;
        RECT 2428.960 2139.805 2429.100 2156.970 ;
        RECT 2435.230 2156.695 2435.490 2157.015 ;
        RECT 2436.580 2156.500 2436.860 2156.870 ;
        RECT 2438.010 2156.815 2438.185 2157.350 ;
        RECT 2439.650 2157.035 2439.910 2157.355 ;
        RECT 2442.880 2156.860 2443.040 2162.030 ;
        RECT 2443.995 2161.940 2444.320 2162.030 ;
        RECT 2443.195 2161.565 2443.515 2161.890 ;
        RECT 2443.225 2161.330 2443.395 2161.565 ;
        RECT 2443.225 2161.155 2443.400 2161.330 ;
        RECT 2443.225 2160.980 2444.200 2161.155 ;
        RECT 2443.195 2156.860 2443.515 2156.980 ;
        RECT 2438.010 2156.640 2441.230 2156.815 ;
        RECT 2442.880 2156.690 2443.515 2156.860 ;
        RECT 2443.195 2156.660 2443.515 2156.690 ;
        RECT 2441.055 2156.490 2441.230 2156.640 ;
        RECT 2441.525 2156.490 2441.850 2156.615 ;
        RECT 2444.025 2156.610 2444.200 2160.980 ;
        RECT 2443.970 2156.490 2444.320 2156.610 ;
        RECT 2441.055 2156.320 2444.320 2156.490 ;
        RECT 2441.525 2156.290 2441.850 2156.320 ;
        RECT 2443.970 2156.260 2444.320 2156.320 ;
        RECT 2452.880 2145.730 2453.020 2214.770 ;
        RECT 2452.820 2145.410 2453.080 2145.730 ;
        RECT 2428.890 2139.435 2429.170 2139.805 ;
        RECT 2411.880 2138.950 2412.140 2139.270 ;
        RECT 2359.230 2058.685 2442.055 2058.855 ;
        RECT 2359.230 2056.890 2359.400 2058.685 ;
        RECT 2441.885 2057.910 2442.055 2058.685 ;
        RECT 2359.545 2057.515 2359.835 2057.635 ;
        RECT 2359.545 2057.510 2359.920 2057.515 ;
        RECT 2359.545 2057.335 2360.830 2057.510 ;
        RECT 2368.105 2057.340 2368.475 2057.710 ;
        RECT 2384.430 2057.340 2384.800 2057.710 ;
        RECT 2400.755 2057.340 2401.125 2057.710 ;
        RECT 2417.080 2057.340 2417.450 2057.710 ;
        RECT 2433.405 2057.340 2433.775 2057.710 ;
        RECT 2441.855 2057.560 2442.205 2057.910 ;
        RECT 2359.545 2057.285 2359.835 2057.335 ;
        RECT 2360.655 2057.145 2360.830 2057.335 ;
        RECT 2369.590 2057.145 2369.940 2057.240 ;
        RECT 2374.195 2057.200 2374.520 2057.265 ;
        RECT 2360.655 2056.970 2369.940 2057.145 ;
        RECT 2369.590 2056.890 2369.940 2056.970 ;
        RECT 2373.080 2057.030 2374.520 2057.200 ;
        RECT 2359.170 2056.540 2359.460 2056.890 ;
        RECT 2362.600 2053.295 2366.260 2053.435 ;
        RECT 2361.810 2052.245 2362.090 2052.620 ;
        RECT 2362.600 2052.615 2362.740 2053.295 ;
        RECT 2363.020 2053.065 2363.280 2053.155 ;
        RECT 2363.020 2052.925 2364.700 2053.065 ;
        RECT 2363.020 2052.835 2363.280 2052.925 ;
        RECT 2364.560 2052.875 2364.700 2052.925 ;
        RECT 2364.560 2052.645 2365.000 2052.875 ;
        RECT 2362.600 2052.365 2363.050 2052.615 ;
        RECT 2364.740 2052.555 2365.000 2052.645 ;
        RECT 2365.520 2052.555 2365.840 2052.875 ;
        RECT 2366.120 2052.615 2366.260 2053.295 ;
        RECT 2366.430 2053.065 2366.710 2053.180 ;
        RECT 2367.510 2053.065 2369.690 2053.175 ;
        RECT 2366.430 2053.015 2369.690 2053.065 ;
        RECT 2366.430 2052.925 2367.650 2053.015 ;
        RECT 2366.430 2052.805 2366.710 2052.925 ;
        RECT 2368.350 2052.615 2368.650 2052.620 ;
        RECT 2362.770 2052.245 2363.050 2052.365 ;
        RECT 2364.060 2052.060 2364.460 2052.225 ;
        RECT 2364.060 2052.035 2364.530 2052.060 ;
        RECT 2362.780 2051.945 2363.040 2052.035 ;
        RECT 2362.780 2051.805 2363.820 2051.945 ;
        RECT 2362.780 2051.715 2363.040 2051.805 ;
        RECT 2363.250 2051.125 2363.530 2051.500 ;
        RECT 2363.680 2051.155 2363.820 2051.805 ;
        RECT 2364.000 2051.715 2364.530 2052.035 ;
        RECT 2364.250 2051.685 2364.530 2051.715 ;
        RECT 2364.970 2051.685 2365.250 2052.060 ;
        RECT 2365.520 2051.755 2365.660 2052.555 ;
        RECT 2366.120 2052.505 2368.650 2052.615 ;
        RECT 2369.140 2052.555 2369.400 2052.875 ;
        RECT 2369.140 2052.505 2369.340 2052.555 ;
        RECT 2366.120 2052.475 2369.340 2052.505 ;
        RECT 2368.370 2052.365 2369.340 2052.475 ;
        RECT 2365.820 2052.225 2366.080 2052.315 ;
        RECT 2368.370 2052.245 2368.650 2052.365 ;
        RECT 2365.820 2052.060 2366.140 2052.225 ;
        RECT 2365.820 2051.995 2366.210 2052.060 ;
        RECT 2365.460 2051.435 2365.720 2051.755 ;
        RECT 2365.930 2051.685 2366.210 2051.995 ;
        RECT 2366.810 2051.685 2367.090 2052.060 ;
        RECT 2367.420 2051.715 2367.680 2052.035 ;
        RECT 2366.440 2051.155 2366.700 2051.475 ;
        RECT 2363.290 2050.735 2363.460 2051.125 ;
        RECT 2363.680 2051.015 2366.640 2051.155 ;
        RECT 2367.480 2051.015 2367.620 2051.715 ;
        RECT 2368.490 2051.685 2368.770 2052.055 ;
        RECT 2368.560 2051.015 2368.700 2051.685 ;
        RECT 2368.940 2051.475 2369.080 2052.365 ;
        RECT 2369.540 2052.035 2369.690 2053.015 ;
        RECT 2369.260 2051.895 2369.690 2052.035 ;
        RECT 2369.260 2051.715 2369.520 2051.895 ;
        RECT 2369.970 2051.665 2370.250 2051.895 ;
        RECT 2373.080 2051.825 2373.240 2057.030 ;
        RECT 2374.195 2056.940 2374.520 2057.030 ;
        RECT 2376.575 2057.170 2376.925 2057.290 ;
        RECT 2385.080 2057.170 2385.430 2057.245 ;
        RECT 2390.520 2057.200 2390.845 2057.265 ;
        RECT 2376.575 2056.970 2385.430 2057.170 ;
        RECT 2376.575 2056.940 2376.925 2056.970 ;
        RECT 2385.080 2056.895 2385.430 2056.970 ;
        RECT 2389.405 2057.030 2390.845 2057.200 ;
        RECT 2373.395 2056.505 2373.715 2056.830 ;
        RECT 2373.425 2056.330 2373.595 2056.505 ;
        RECT 2373.425 2056.155 2373.600 2056.330 ;
        RECT 2373.425 2055.980 2374.400 2056.155 ;
        RECT 2373.395 2051.825 2373.715 2051.945 ;
        RECT 2370.580 2051.665 2370.840 2051.755 ;
        RECT 2369.680 2051.525 2370.840 2051.665 ;
        RECT 2373.080 2051.655 2373.715 2051.825 ;
        RECT 2373.395 2051.625 2373.715 2051.655 ;
        RECT 2374.225 2051.610 2374.400 2055.980 ;
        RECT 2378.925 2053.295 2382.585 2053.435 ;
        RECT 2378.135 2052.245 2378.415 2052.620 ;
        RECT 2378.925 2052.615 2379.065 2053.295 ;
        RECT 2379.345 2053.065 2379.605 2053.155 ;
        RECT 2379.345 2052.925 2381.025 2053.065 ;
        RECT 2379.345 2052.835 2379.605 2052.925 ;
        RECT 2380.885 2052.875 2381.025 2052.925 ;
        RECT 2380.885 2052.645 2381.325 2052.875 ;
        RECT 2378.925 2052.365 2379.375 2052.615 ;
        RECT 2381.065 2052.555 2381.325 2052.645 ;
        RECT 2381.845 2052.555 2382.165 2052.875 ;
        RECT 2382.445 2052.615 2382.585 2053.295 ;
        RECT 2382.755 2053.065 2383.035 2053.180 ;
        RECT 2383.835 2053.065 2386.015 2053.175 ;
        RECT 2382.755 2053.015 2386.015 2053.065 ;
        RECT 2382.755 2052.925 2383.975 2053.015 ;
        RECT 2382.755 2052.805 2383.035 2052.925 ;
        RECT 2384.675 2052.615 2384.975 2052.620 ;
        RECT 2379.095 2052.245 2379.375 2052.365 ;
        RECT 2380.385 2052.060 2380.785 2052.225 ;
        RECT 2380.385 2052.035 2380.855 2052.060 ;
        RECT 2379.105 2051.945 2379.365 2052.035 ;
        RECT 2379.105 2051.805 2380.145 2051.945 ;
        RECT 2379.105 2051.715 2379.365 2051.805 ;
        RECT 2368.880 2051.155 2369.140 2051.475 ;
        RECT 2369.680 2051.015 2369.820 2051.525 ;
        RECT 2370.580 2051.435 2370.840 2051.525 ;
        RECT 2374.170 2051.260 2374.520 2051.610 ;
        RECT 2379.575 2051.125 2379.855 2051.500 ;
        RECT 2380.005 2051.155 2380.145 2051.805 ;
        RECT 2380.325 2051.715 2380.855 2052.035 ;
        RECT 2380.575 2051.685 2380.855 2051.715 ;
        RECT 2381.295 2051.685 2381.575 2052.060 ;
        RECT 2381.845 2051.755 2381.985 2052.555 ;
        RECT 2382.445 2052.505 2384.975 2052.615 ;
        RECT 2385.465 2052.555 2385.725 2052.875 ;
        RECT 2385.465 2052.505 2385.665 2052.555 ;
        RECT 2382.445 2052.475 2385.665 2052.505 ;
        RECT 2384.695 2052.365 2385.665 2052.475 ;
        RECT 2382.145 2052.225 2382.405 2052.315 ;
        RECT 2384.695 2052.245 2384.975 2052.365 ;
        RECT 2382.145 2052.060 2382.465 2052.225 ;
        RECT 2382.145 2051.995 2382.535 2052.060 ;
        RECT 2381.785 2051.435 2382.045 2051.755 ;
        RECT 2382.255 2051.685 2382.535 2051.995 ;
        RECT 2383.135 2051.685 2383.415 2052.060 ;
        RECT 2383.745 2051.715 2384.005 2052.035 ;
        RECT 2382.765 2051.155 2383.025 2051.475 ;
        RECT 2371.865 2051.105 2372.035 2051.110 ;
        RECT 2367.480 2050.875 2369.820 2051.015 ;
        RECT 2371.775 2050.755 2372.115 2051.105 ;
        RECT 2371.775 2050.735 2372.035 2050.755 ;
        RECT 2363.290 2050.565 2372.035 2050.735 ;
        RECT 2379.615 2050.735 2379.785 2051.125 ;
        RECT 2380.005 2051.015 2382.965 2051.155 ;
        RECT 2383.805 2051.015 2383.945 2051.715 ;
        RECT 2384.815 2051.685 2385.095 2052.055 ;
        RECT 2384.885 2051.015 2385.025 2051.685 ;
        RECT 2385.265 2051.475 2385.405 2052.365 ;
        RECT 2385.865 2052.035 2386.015 2053.015 ;
        RECT 2385.585 2051.895 2386.015 2052.035 ;
        RECT 2385.585 2051.715 2385.845 2051.895 ;
        RECT 2386.295 2051.665 2386.575 2051.895 ;
        RECT 2389.405 2051.825 2389.565 2057.030 ;
        RECT 2390.520 2056.940 2390.845 2057.030 ;
        RECT 2392.900 2057.175 2393.250 2057.295 ;
        RECT 2401.405 2057.175 2401.755 2057.250 ;
        RECT 2406.845 2057.200 2407.170 2057.265 ;
        RECT 2392.900 2056.975 2401.755 2057.175 ;
        RECT 2392.900 2056.945 2393.250 2056.975 ;
        RECT 2401.405 2056.900 2401.755 2056.975 ;
        RECT 2405.730 2057.030 2407.170 2057.200 ;
        RECT 2389.720 2056.505 2390.040 2056.830 ;
        RECT 2389.750 2056.330 2389.920 2056.505 ;
        RECT 2389.750 2056.155 2389.925 2056.330 ;
        RECT 2389.750 2055.980 2390.725 2056.155 ;
        RECT 2389.720 2051.825 2390.040 2051.945 ;
        RECT 2386.905 2051.665 2387.165 2051.755 ;
        RECT 2386.005 2051.525 2387.165 2051.665 ;
        RECT 2389.405 2051.655 2390.040 2051.825 ;
        RECT 2389.720 2051.625 2390.040 2051.655 ;
        RECT 2390.550 2051.610 2390.725 2055.980 ;
        RECT 2395.250 2053.295 2398.910 2053.435 ;
        RECT 2394.460 2052.245 2394.740 2052.620 ;
        RECT 2395.250 2052.615 2395.390 2053.295 ;
        RECT 2395.670 2053.065 2395.930 2053.155 ;
        RECT 2395.670 2052.925 2397.350 2053.065 ;
        RECT 2395.670 2052.835 2395.930 2052.925 ;
        RECT 2397.210 2052.875 2397.350 2052.925 ;
        RECT 2397.210 2052.645 2397.650 2052.875 ;
        RECT 2395.250 2052.365 2395.700 2052.615 ;
        RECT 2397.390 2052.555 2397.650 2052.645 ;
        RECT 2398.170 2052.555 2398.490 2052.875 ;
        RECT 2398.770 2052.615 2398.910 2053.295 ;
        RECT 2399.080 2053.065 2399.360 2053.180 ;
        RECT 2400.160 2053.065 2402.340 2053.175 ;
        RECT 2399.080 2053.015 2402.340 2053.065 ;
        RECT 2399.080 2052.925 2400.300 2053.015 ;
        RECT 2399.080 2052.805 2399.360 2052.925 ;
        RECT 2401.000 2052.615 2401.300 2052.620 ;
        RECT 2395.420 2052.245 2395.700 2052.365 ;
        RECT 2393.020 2051.910 2393.280 2052.230 ;
        RECT 2396.710 2052.060 2397.110 2052.225 ;
        RECT 2396.710 2052.035 2397.180 2052.060 ;
        RECT 2395.430 2051.945 2395.690 2052.035 ;
        RECT 2385.205 2051.155 2385.465 2051.475 ;
        RECT 2386.005 2051.015 2386.145 2051.525 ;
        RECT 2386.905 2051.435 2387.165 2051.525 ;
        RECT 2390.495 2051.260 2390.845 2051.610 ;
        RECT 2388.190 2051.105 2388.360 2051.110 ;
        RECT 2383.805 2050.875 2386.145 2051.015 ;
        RECT 2388.100 2050.755 2388.440 2051.105 ;
        RECT 2388.100 2050.735 2388.360 2050.755 ;
        RECT 2379.615 2050.565 2388.360 2050.735 ;
        RECT 2376.460 2050.150 2376.720 2050.470 ;
        RECT 2376.520 2042.370 2376.660 2050.150 ;
        RECT 2376.460 2042.050 2376.720 2042.370 ;
        RECT 2393.080 2035.570 2393.220 2051.910 ;
        RECT 2395.430 2051.805 2396.470 2051.945 ;
        RECT 2395.430 2051.715 2395.690 2051.805 ;
        RECT 2395.900 2051.125 2396.180 2051.500 ;
        RECT 2396.330 2051.155 2396.470 2051.805 ;
        RECT 2396.650 2051.715 2397.180 2052.035 ;
        RECT 2396.900 2051.685 2397.180 2051.715 ;
        RECT 2397.620 2051.685 2397.900 2052.060 ;
        RECT 2398.170 2051.755 2398.310 2052.555 ;
        RECT 2398.770 2052.505 2401.300 2052.615 ;
        RECT 2401.790 2052.555 2402.050 2052.875 ;
        RECT 2401.790 2052.505 2401.990 2052.555 ;
        RECT 2398.770 2052.475 2401.990 2052.505 ;
        RECT 2401.020 2052.365 2401.990 2052.475 ;
        RECT 2398.470 2052.225 2398.730 2052.315 ;
        RECT 2401.020 2052.245 2401.300 2052.365 ;
        RECT 2398.470 2052.060 2398.790 2052.225 ;
        RECT 2398.470 2051.995 2398.860 2052.060 ;
        RECT 2398.110 2051.435 2398.370 2051.755 ;
        RECT 2398.580 2051.685 2398.860 2051.995 ;
        RECT 2399.460 2051.685 2399.740 2052.060 ;
        RECT 2400.070 2051.715 2400.330 2052.035 ;
        RECT 2399.090 2051.155 2399.350 2051.475 ;
        RECT 2395.940 2050.735 2396.110 2051.125 ;
        RECT 2396.330 2051.015 2399.290 2051.155 ;
        RECT 2400.130 2051.015 2400.270 2051.715 ;
        RECT 2401.140 2051.685 2401.420 2052.055 ;
        RECT 2401.210 2051.015 2401.350 2051.685 ;
        RECT 2401.590 2051.475 2401.730 2052.365 ;
        RECT 2402.190 2052.035 2402.340 2053.015 ;
        RECT 2401.910 2051.895 2402.340 2052.035 ;
        RECT 2401.910 2051.715 2402.170 2051.895 ;
        RECT 2402.620 2051.665 2402.900 2051.895 ;
        RECT 2405.730 2051.825 2405.890 2057.030 ;
        RECT 2406.845 2056.940 2407.170 2057.030 ;
        RECT 2409.180 2057.170 2409.530 2057.290 ;
        RECT 2417.730 2057.170 2418.080 2057.245 ;
        RECT 2423.170 2057.200 2423.495 2057.265 ;
        RECT 2409.180 2056.970 2418.080 2057.170 ;
        RECT 2409.180 2056.940 2409.530 2056.970 ;
        RECT 2417.730 2056.895 2418.080 2056.970 ;
        RECT 2422.055 2057.030 2423.495 2057.200 ;
        RECT 2406.045 2056.505 2406.365 2056.830 ;
        RECT 2406.075 2056.330 2406.245 2056.505 ;
        RECT 2406.075 2056.155 2406.250 2056.330 ;
        RECT 2406.075 2055.980 2407.050 2056.155 ;
        RECT 2406.045 2051.825 2406.365 2051.945 ;
        RECT 2403.230 2051.665 2403.490 2051.755 ;
        RECT 2402.330 2051.525 2403.490 2051.665 ;
        RECT 2405.730 2051.655 2406.365 2051.825 ;
        RECT 2406.045 2051.625 2406.365 2051.655 ;
        RECT 2406.875 2051.610 2407.050 2055.980 ;
        RECT 2411.575 2053.295 2415.235 2053.435 ;
        RECT 2410.785 2052.245 2411.065 2052.620 ;
        RECT 2411.575 2052.615 2411.715 2053.295 ;
        RECT 2411.995 2053.065 2412.255 2053.155 ;
        RECT 2411.995 2052.925 2413.675 2053.065 ;
        RECT 2411.995 2052.835 2412.255 2052.925 ;
        RECT 2413.535 2052.875 2413.675 2052.925 ;
        RECT 2413.535 2052.645 2413.975 2052.875 ;
        RECT 2411.575 2052.365 2412.025 2052.615 ;
        RECT 2413.715 2052.555 2413.975 2052.645 ;
        RECT 2414.495 2052.555 2414.815 2052.875 ;
        RECT 2415.095 2052.615 2415.235 2053.295 ;
        RECT 2415.405 2053.065 2415.685 2053.180 ;
        RECT 2416.485 2053.065 2418.665 2053.175 ;
        RECT 2415.405 2053.015 2418.665 2053.065 ;
        RECT 2415.405 2052.925 2416.625 2053.015 ;
        RECT 2415.405 2052.805 2415.685 2052.925 ;
        RECT 2417.325 2052.615 2417.625 2052.620 ;
        RECT 2411.745 2052.245 2412.025 2052.365 ;
        RECT 2413.035 2052.060 2413.435 2052.225 ;
        RECT 2413.035 2052.035 2413.505 2052.060 ;
        RECT 2411.755 2051.945 2412.015 2052.035 ;
        RECT 2411.755 2051.805 2412.795 2051.945 ;
        RECT 2411.755 2051.715 2412.015 2051.805 ;
        RECT 2401.530 2051.155 2401.790 2051.475 ;
        RECT 2402.330 2051.015 2402.470 2051.525 ;
        RECT 2403.230 2051.435 2403.490 2051.525 ;
        RECT 2406.820 2051.260 2407.170 2051.610 ;
        RECT 2412.225 2051.125 2412.505 2051.500 ;
        RECT 2412.655 2051.155 2412.795 2051.805 ;
        RECT 2412.975 2051.715 2413.505 2052.035 ;
        RECT 2413.225 2051.685 2413.505 2051.715 ;
        RECT 2413.945 2051.685 2414.225 2052.060 ;
        RECT 2414.495 2051.755 2414.635 2052.555 ;
        RECT 2415.095 2052.505 2417.625 2052.615 ;
        RECT 2418.115 2052.555 2418.375 2052.875 ;
        RECT 2418.115 2052.505 2418.315 2052.555 ;
        RECT 2415.095 2052.475 2418.315 2052.505 ;
        RECT 2417.345 2052.365 2418.315 2052.475 ;
        RECT 2414.795 2052.225 2415.055 2052.315 ;
        RECT 2417.345 2052.245 2417.625 2052.365 ;
        RECT 2414.795 2052.060 2415.115 2052.225 ;
        RECT 2414.795 2051.995 2415.185 2052.060 ;
        RECT 2414.435 2051.435 2414.695 2051.755 ;
        RECT 2414.905 2051.685 2415.185 2051.995 ;
        RECT 2415.785 2051.685 2416.065 2052.060 ;
        RECT 2416.395 2051.715 2416.655 2052.035 ;
        RECT 2415.415 2051.155 2415.675 2051.475 ;
        RECT 2404.515 2051.105 2404.685 2051.110 ;
        RECT 2400.130 2050.875 2402.470 2051.015 ;
        RECT 2404.425 2050.755 2404.765 2051.105 ;
        RECT 2404.425 2050.735 2404.685 2050.755 ;
        RECT 2395.940 2050.565 2404.685 2050.735 ;
        RECT 2412.265 2050.735 2412.435 2051.125 ;
        RECT 2412.655 2051.015 2415.615 2051.155 ;
        RECT 2416.455 2051.015 2416.595 2051.715 ;
        RECT 2417.465 2051.685 2417.745 2052.055 ;
        RECT 2417.535 2051.015 2417.675 2051.685 ;
        RECT 2417.915 2051.475 2418.055 2052.365 ;
        RECT 2418.515 2052.035 2418.665 2053.015 ;
        RECT 2418.235 2051.895 2418.665 2052.035 ;
        RECT 2418.235 2051.715 2418.495 2051.895 ;
        RECT 2418.945 2051.665 2419.225 2051.895 ;
        RECT 2422.055 2051.825 2422.215 2057.030 ;
        RECT 2423.170 2056.940 2423.495 2057.030 ;
        RECT 2425.505 2057.170 2425.855 2057.290 ;
        RECT 2434.060 2057.170 2434.410 2057.245 ;
        RECT 2439.495 2057.200 2439.820 2057.265 ;
        RECT 2425.505 2056.970 2434.410 2057.170 ;
        RECT 2425.505 2056.940 2425.855 2056.970 ;
        RECT 2434.060 2056.895 2434.410 2056.970 ;
        RECT 2438.380 2057.030 2439.820 2057.200 ;
        RECT 2422.370 2056.505 2422.690 2056.830 ;
        RECT 2422.400 2056.330 2422.570 2056.505 ;
        RECT 2422.400 2056.155 2422.575 2056.330 ;
        RECT 2422.400 2055.980 2423.375 2056.155 ;
        RECT 2422.370 2051.825 2422.690 2051.945 ;
        RECT 2419.555 2051.665 2419.815 2051.755 ;
        RECT 2418.655 2051.525 2419.815 2051.665 ;
        RECT 2422.055 2051.655 2422.690 2051.825 ;
        RECT 2422.370 2051.625 2422.690 2051.655 ;
        RECT 2423.200 2051.610 2423.375 2055.980 ;
        RECT 2427.900 2053.295 2431.560 2053.435 ;
        RECT 2427.110 2052.245 2427.390 2052.620 ;
        RECT 2427.900 2052.615 2428.040 2053.295 ;
        RECT 2428.320 2053.065 2428.580 2053.155 ;
        RECT 2428.320 2052.925 2430.000 2053.065 ;
        RECT 2428.320 2052.835 2428.580 2052.925 ;
        RECT 2429.860 2052.875 2430.000 2052.925 ;
        RECT 2429.860 2052.645 2430.300 2052.875 ;
        RECT 2427.900 2052.365 2428.350 2052.615 ;
        RECT 2430.040 2052.555 2430.300 2052.645 ;
        RECT 2430.820 2052.555 2431.140 2052.875 ;
        RECT 2431.420 2052.615 2431.560 2053.295 ;
        RECT 2431.730 2053.065 2432.010 2053.180 ;
        RECT 2432.810 2053.065 2434.990 2053.175 ;
        RECT 2431.730 2053.015 2434.990 2053.065 ;
        RECT 2431.730 2052.925 2432.950 2053.015 ;
        RECT 2431.730 2052.805 2432.010 2052.925 ;
        RECT 2433.650 2052.615 2433.950 2052.620 ;
        RECT 2428.070 2052.245 2428.350 2052.365 ;
        RECT 2425.680 2051.910 2425.940 2052.230 ;
        RECT 2429.360 2052.060 2429.760 2052.225 ;
        RECT 2429.360 2052.035 2429.830 2052.060 ;
        RECT 2428.080 2051.945 2428.340 2052.035 ;
        RECT 2417.855 2051.155 2418.115 2051.475 ;
        RECT 2418.655 2051.015 2418.795 2051.525 ;
        RECT 2419.555 2051.435 2419.815 2051.525 ;
        RECT 2423.145 2051.260 2423.495 2051.610 ;
        RECT 2420.840 2051.105 2421.010 2051.110 ;
        RECT 2416.455 2050.875 2418.795 2051.015 ;
        RECT 2420.750 2050.755 2421.090 2051.105 ;
        RECT 2420.750 2050.735 2421.010 2050.755 ;
        RECT 2412.265 2050.565 2421.010 2050.735 ;
        RECT 2409.120 2050.150 2409.380 2050.470 ;
        RECT 2409.180 2035.765 2409.320 2050.150 ;
        RECT 2425.740 2035.765 2425.880 2051.910 ;
        RECT 2428.080 2051.805 2429.120 2051.945 ;
        RECT 2428.080 2051.715 2428.340 2051.805 ;
        RECT 2428.550 2051.125 2428.830 2051.500 ;
        RECT 2428.980 2051.155 2429.120 2051.805 ;
        RECT 2429.300 2051.715 2429.830 2052.035 ;
        RECT 2429.550 2051.685 2429.830 2051.715 ;
        RECT 2430.270 2051.685 2430.550 2052.060 ;
        RECT 2430.820 2051.755 2430.960 2052.555 ;
        RECT 2431.420 2052.505 2433.950 2052.615 ;
        RECT 2434.440 2052.555 2434.700 2052.875 ;
        RECT 2434.440 2052.505 2434.640 2052.555 ;
        RECT 2431.420 2052.475 2434.640 2052.505 ;
        RECT 2433.670 2052.365 2434.640 2052.475 ;
        RECT 2431.120 2052.225 2431.380 2052.315 ;
        RECT 2433.670 2052.245 2433.950 2052.365 ;
        RECT 2431.120 2052.060 2431.440 2052.225 ;
        RECT 2431.120 2051.995 2431.510 2052.060 ;
        RECT 2430.760 2051.435 2431.020 2051.755 ;
        RECT 2431.230 2051.685 2431.510 2051.995 ;
        RECT 2432.110 2051.685 2432.390 2052.060 ;
        RECT 2432.720 2051.715 2432.980 2052.035 ;
        RECT 2431.740 2051.155 2432.000 2051.475 ;
        RECT 2428.590 2050.735 2428.760 2051.125 ;
        RECT 2428.980 2051.015 2431.940 2051.155 ;
        RECT 2432.780 2051.015 2432.920 2051.715 ;
        RECT 2433.790 2051.685 2434.070 2052.055 ;
        RECT 2433.860 2051.015 2434.000 2051.685 ;
        RECT 2434.240 2051.475 2434.380 2052.365 ;
        RECT 2434.840 2052.035 2434.990 2053.015 ;
        RECT 2434.560 2051.895 2434.990 2052.035 ;
        RECT 2434.560 2051.715 2434.820 2051.895 ;
        RECT 2435.270 2051.665 2435.550 2051.895 ;
        RECT 2438.380 2051.825 2438.540 2057.030 ;
        RECT 2439.495 2056.940 2439.820 2057.030 ;
        RECT 2438.695 2056.505 2439.015 2056.830 ;
        RECT 2438.725 2056.330 2438.895 2056.505 ;
        RECT 2438.725 2056.155 2438.900 2056.330 ;
        RECT 2438.725 2055.980 2439.700 2056.155 ;
        RECT 2438.695 2051.825 2439.015 2051.945 ;
        RECT 2435.880 2051.665 2436.140 2051.755 ;
        RECT 2434.980 2051.525 2436.140 2051.665 ;
        RECT 2438.380 2051.655 2439.015 2051.825 ;
        RECT 2438.695 2051.625 2439.015 2051.655 ;
        RECT 2439.525 2051.610 2439.700 2055.980 ;
        RECT 2434.180 2051.155 2434.440 2051.475 ;
        RECT 2434.980 2051.015 2435.120 2051.525 ;
        RECT 2435.880 2051.435 2436.140 2051.525 ;
        RECT 2439.470 2051.260 2439.820 2051.610 ;
        RECT 2437.165 2051.105 2437.335 2051.110 ;
        RECT 2432.780 2050.875 2435.120 2051.015 ;
        RECT 2437.075 2050.755 2437.415 2051.105 ;
        RECT 2437.075 2050.735 2437.335 2050.755 ;
        RECT 2428.590 2050.565 2437.335 2050.735 ;
        RECT 2453.740 2049.870 2454.000 2050.190 ;
        RECT 2393.020 2035.250 2393.280 2035.570 ;
        RECT 2409.110 2035.395 2409.390 2035.765 ;
        RECT 2425.670 2035.395 2425.950 2035.765 ;
        RECT 2359.235 1953.690 2453.230 1953.860 ;
        RECT 2359.235 1951.895 2359.405 1953.690 ;
        RECT 2453.060 1952.915 2453.230 1953.690 ;
        RECT 2359.545 1952.515 2359.835 1952.640 ;
        RECT 2359.545 1952.510 2359.865 1952.515 ;
        RECT 2359.545 1952.340 2360.860 1952.510 ;
        RECT 2370.320 1952.345 2370.695 1952.715 ;
        RECT 2388.880 1952.345 2389.255 1952.715 ;
        RECT 2407.440 1952.345 2407.815 1952.715 ;
        RECT 2426.000 1952.345 2426.375 1952.715 ;
        RECT 2444.560 1952.345 2444.935 1952.715 ;
        RECT 2453.030 1952.565 2453.380 1952.915 ;
        RECT 2359.545 1952.290 2359.835 1952.340 ;
        RECT 2360.690 1952.145 2360.860 1952.340 ;
        RECT 2370.995 1952.145 2371.345 1952.245 ;
        RECT 2376.430 1952.205 2376.755 1952.270 ;
        RECT 2360.690 1951.975 2371.345 1952.145 ;
        RECT 2370.995 1951.895 2371.345 1951.975 ;
        RECT 2375.315 1952.035 2376.755 1952.205 ;
        RECT 2359.170 1951.545 2359.460 1951.895 ;
        RECT 2370.150 1948.430 2374.285 1948.620 ;
        RECT 2370.150 1948.180 2370.340 1948.430 ;
        RECT 2361.815 1947.805 2362.095 1948.180 ;
        RECT 2366.585 1947.835 2366.845 1948.155 ;
        RECT 2361.825 1947.555 2362.085 1947.805 ;
        RECT 2364.255 1947.595 2364.535 1947.620 ;
        RECT 2362.785 1947.275 2363.045 1947.595 ;
        RECT 2363.905 1947.505 2364.535 1947.595 ;
        RECT 2366.225 1947.505 2366.485 1947.595 ;
        RECT 2363.905 1947.365 2366.485 1947.505 ;
        RECT 2363.905 1947.275 2364.535 1947.365 ;
        RECT 2366.225 1947.275 2366.485 1947.365 ;
        RECT 2362.295 1946.685 2362.575 1947.060 ;
        RECT 2362.845 1946.475 2362.985 1947.275 ;
        RECT 2364.255 1947.245 2364.535 1947.275 ;
        RECT 2365.695 1947.035 2365.975 1947.060 ;
        RECT 2365.695 1946.715 2366.225 1947.035 ;
        RECT 2365.695 1946.685 2365.975 1946.715 ;
        RECT 2362.785 1946.155 2363.045 1946.475 ;
        RECT 2364.745 1946.385 2365.005 1946.475 ;
        RECT 2366.225 1946.385 2366.485 1946.475 ;
        RECT 2366.645 1946.385 2366.785 1947.835 ;
        RECT 2368.135 1947.805 2368.415 1948.180 ;
        RECT 2369.145 1947.835 2369.405 1948.155 ;
        RECT 2369.625 1947.835 2369.885 1948.155 ;
        RECT 2366.935 1947.245 2367.215 1947.620 ;
        RECT 2368.205 1947.615 2368.345 1947.805 ;
        RECT 2368.015 1947.505 2368.345 1947.615 ;
        RECT 2367.725 1947.365 2368.345 1947.505 ;
        RECT 2367.005 1946.475 2367.145 1947.245 ;
        RECT 2367.725 1946.475 2367.865 1947.365 ;
        RECT 2368.015 1947.245 2368.295 1947.365 ;
        RECT 2368.665 1946.945 2368.925 1947.035 ;
        RECT 2368.085 1946.805 2368.925 1946.945 ;
        RECT 2364.745 1946.245 2365.785 1946.385 ;
        RECT 2364.745 1946.155 2365.005 1946.245 ;
        RECT 2365.645 1946.005 2365.785 1946.245 ;
        RECT 2366.225 1946.245 2366.785 1946.385 ;
        RECT 2366.225 1946.155 2366.485 1946.245 ;
        RECT 2366.945 1946.155 2367.205 1946.475 ;
        RECT 2367.665 1946.155 2367.925 1946.475 ;
        RECT 2368.085 1946.005 2368.225 1946.805 ;
        RECT 2368.665 1946.715 2368.925 1946.805 ;
        RECT 2369.205 1946.475 2369.345 1947.835 ;
        RECT 2369.625 1947.785 2369.825 1947.835 ;
        RECT 2370.095 1947.805 2370.375 1948.180 ;
        RECT 2371.095 1947.805 2371.375 1948.180 ;
        RECT 2374.095 1947.795 2374.285 1948.430 ;
        RECT 2369.565 1947.615 2369.825 1947.785 ;
        RECT 2369.565 1947.245 2370.065 1947.615 ;
        RECT 2370.625 1947.275 2370.885 1947.595 ;
        RECT 2374.025 1947.445 2374.365 1947.795 ;
        RECT 2374.115 1947.440 2374.285 1947.445 ;
        RECT 2369.565 1946.475 2369.705 1947.245 ;
        RECT 2370.685 1946.475 2370.825 1947.275 ;
        RECT 2375.315 1946.860 2375.475 1952.035 ;
        RECT 2376.430 1951.945 2376.755 1952.035 ;
        RECT 2378.810 1952.175 2379.160 1952.295 ;
        RECT 2389.555 1952.175 2389.905 1952.250 ;
        RECT 2394.990 1952.205 2395.315 1952.270 ;
        RECT 2378.810 1951.975 2389.905 1952.175 ;
        RECT 2378.810 1951.945 2379.160 1951.975 ;
        RECT 2389.555 1951.900 2389.905 1951.975 ;
        RECT 2393.875 1952.035 2395.315 1952.205 ;
        RECT 2375.630 1951.510 2375.950 1951.835 ;
        RECT 2375.660 1951.335 2375.830 1951.510 ;
        RECT 2375.660 1951.160 2375.835 1951.335 ;
        RECT 2375.660 1950.985 2376.635 1951.160 ;
        RECT 2375.630 1946.860 2375.950 1946.980 ;
        RECT 2375.315 1946.690 2375.950 1946.860 ;
        RECT 2375.630 1946.660 2375.950 1946.690 ;
        RECT 2376.460 1946.610 2376.635 1950.985 ;
        RECT 2388.710 1948.430 2392.845 1948.620 ;
        RECT 2388.710 1948.180 2388.900 1948.430 ;
        RECT 2380.375 1947.805 2380.655 1948.180 ;
        RECT 2385.145 1947.835 2385.405 1948.155 ;
        RECT 2380.385 1947.555 2380.645 1947.805 ;
        RECT 2382.815 1947.595 2383.095 1947.620 ;
        RECT 2381.345 1947.275 2381.605 1947.595 ;
        RECT 2382.465 1947.505 2383.095 1947.595 ;
        RECT 2384.785 1947.505 2385.045 1947.595 ;
        RECT 2382.465 1947.365 2385.045 1947.505 ;
        RECT 2382.465 1947.275 2383.095 1947.365 ;
        RECT 2384.785 1947.275 2385.045 1947.365 ;
        RECT 2380.855 1946.685 2381.135 1947.060 ;
        RECT 2368.905 1946.245 2369.345 1946.475 ;
        RECT 2368.905 1946.155 2369.165 1946.245 ;
        RECT 2369.505 1946.155 2369.765 1946.475 ;
        RECT 2370.625 1946.155 2370.885 1946.475 ;
        RECT 2372.055 1946.125 2372.335 1946.500 ;
        RECT 2376.405 1946.260 2376.755 1946.610 ;
        RECT 2381.405 1946.475 2381.545 1947.275 ;
        RECT 2382.815 1947.245 2383.095 1947.275 ;
        RECT 2384.255 1947.035 2384.535 1947.060 ;
        RECT 2384.255 1946.715 2384.785 1947.035 ;
        RECT 2384.255 1946.685 2384.535 1946.715 ;
        RECT 2381.345 1946.155 2381.605 1946.475 ;
        RECT 2383.305 1946.385 2383.565 1946.475 ;
        RECT 2384.785 1946.385 2385.045 1946.475 ;
        RECT 2385.205 1946.385 2385.345 1947.835 ;
        RECT 2386.695 1947.805 2386.975 1948.180 ;
        RECT 2387.705 1947.835 2387.965 1948.155 ;
        RECT 2388.185 1947.835 2388.445 1948.155 ;
        RECT 2385.495 1947.245 2385.775 1947.620 ;
        RECT 2386.765 1947.615 2386.905 1947.805 ;
        RECT 2386.575 1947.505 2386.905 1947.615 ;
        RECT 2386.285 1947.365 2386.905 1947.505 ;
        RECT 2385.565 1946.475 2385.705 1947.245 ;
        RECT 2386.285 1946.475 2386.425 1947.365 ;
        RECT 2386.575 1947.245 2386.855 1947.365 ;
        RECT 2387.225 1946.945 2387.485 1947.035 ;
        RECT 2386.645 1946.805 2387.485 1946.945 ;
        RECT 2383.305 1946.245 2384.345 1946.385 ;
        RECT 2383.305 1946.155 2383.565 1946.245 ;
        RECT 2365.645 1945.865 2368.225 1946.005 ;
        RECT 2384.205 1946.005 2384.345 1946.245 ;
        RECT 2384.785 1946.245 2385.345 1946.385 ;
        RECT 2384.785 1946.155 2385.045 1946.245 ;
        RECT 2385.505 1946.155 2385.765 1946.475 ;
        RECT 2386.225 1946.155 2386.485 1946.475 ;
        RECT 2386.645 1946.005 2386.785 1946.805 ;
        RECT 2387.225 1946.715 2387.485 1946.805 ;
        RECT 2387.765 1946.475 2387.905 1947.835 ;
        RECT 2388.185 1947.785 2388.385 1947.835 ;
        RECT 2388.655 1947.805 2388.935 1948.180 ;
        RECT 2389.655 1947.805 2389.935 1948.180 ;
        RECT 2392.655 1947.795 2392.845 1948.430 ;
        RECT 2388.125 1947.615 2388.385 1947.785 ;
        RECT 2388.125 1947.245 2388.625 1947.615 ;
        RECT 2389.185 1947.275 2389.445 1947.595 ;
        RECT 2392.585 1947.445 2392.925 1947.795 ;
        RECT 2392.675 1947.440 2392.845 1947.445 ;
        RECT 2388.125 1946.475 2388.265 1947.245 ;
        RECT 2389.245 1946.475 2389.385 1947.275 ;
        RECT 2393.875 1946.860 2394.035 1952.035 ;
        RECT 2394.990 1951.945 2395.315 1952.035 ;
        RECT 2397.370 1952.180 2397.720 1952.300 ;
        RECT 2408.110 1952.180 2408.460 1952.255 ;
        RECT 2413.550 1952.205 2413.875 1952.270 ;
        RECT 2397.370 1951.980 2408.460 1952.180 ;
        RECT 2397.370 1951.950 2397.720 1951.980 ;
        RECT 2408.110 1951.905 2408.460 1951.980 ;
        RECT 2412.435 1952.035 2413.875 1952.205 ;
        RECT 2394.190 1951.510 2394.510 1951.835 ;
        RECT 2394.220 1951.335 2394.390 1951.510 ;
        RECT 2394.220 1951.160 2394.395 1951.335 ;
        RECT 2394.220 1950.985 2395.195 1951.160 ;
        RECT 2394.190 1946.860 2394.510 1946.980 ;
        RECT 2393.875 1946.690 2394.510 1946.860 ;
        RECT 2394.190 1946.660 2394.510 1946.690 ;
        RECT 2395.020 1946.610 2395.195 1950.985 ;
        RECT 2407.270 1948.430 2411.405 1948.620 ;
        RECT 2407.270 1948.180 2407.460 1948.430 ;
        RECT 2398.935 1947.805 2399.215 1948.180 ;
        RECT 2403.705 1947.835 2403.965 1948.155 ;
        RECT 2398.945 1947.555 2399.205 1947.805 ;
        RECT 2401.375 1947.595 2401.655 1947.620 ;
        RECT 2397.160 1947.190 2397.420 1947.510 ;
        RECT 2399.905 1947.275 2400.165 1947.595 ;
        RECT 2401.025 1947.505 2401.655 1947.595 ;
        RECT 2403.345 1947.505 2403.605 1947.595 ;
        RECT 2401.025 1947.365 2403.605 1947.505 ;
        RECT 2401.025 1947.275 2401.655 1947.365 ;
        RECT 2403.345 1947.275 2403.605 1947.365 ;
        RECT 2387.465 1946.245 2387.905 1946.475 ;
        RECT 2387.465 1946.155 2387.725 1946.245 ;
        RECT 2388.065 1946.155 2388.325 1946.475 ;
        RECT 2389.185 1946.155 2389.445 1946.475 ;
        RECT 2390.615 1946.125 2390.895 1946.500 ;
        RECT 2394.965 1946.260 2395.315 1946.610 ;
        RECT 2384.205 1945.865 2386.785 1946.005 ;
        RECT 2378.760 1945.150 2379.020 1945.470 ;
        RECT 2378.820 1939.010 2378.960 1945.150 ;
        RECT 2397.220 1939.010 2397.360 1947.190 ;
        RECT 2399.415 1946.685 2399.695 1947.060 ;
        RECT 2399.965 1946.475 2400.105 1947.275 ;
        RECT 2401.375 1947.245 2401.655 1947.275 ;
        RECT 2402.815 1947.035 2403.095 1947.060 ;
        RECT 2402.815 1946.715 2403.345 1947.035 ;
        RECT 2402.815 1946.685 2403.095 1946.715 ;
        RECT 2399.905 1946.155 2400.165 1946.475 ;
        RECT 2401.865 1946.385 2402.125 1946.475 ;
        RECT 2403.345 1946.385 2403.605 1946.475 ;
        RECT 2403.765 1946.385 2403.905 1947.835 ;
        RECT 2405.255 1947.805 2405.535 1948.180 ;
        RECT 2406.265 1947.835 2406.525 1948.155 ;
        RECT 2406.745 1947.835 2407.005 1948.155 ;
        RECT 2404.055 1947.245 2404.335 1947.620 ;
        RECT 2405.325 1947.615 2405.465 1947.805 ;
        RECT 2405.135 1947.505 2405.465 1947.615 ;
        RECT 2404.845 1947.365 2405.465 1947.505 ;
        RECT 2404.125 1946.475 2404.265 1947.245 ;
        RECT 2404.845 1946.475 2404.985 1947.365 ;
        RECT 2405.135 1947.245 2405.415 1947.365 ;
        RECT 2405.785 1946.945 2406.045 1947.035 ;
        RECT 2405.205 1946.805 2406.045 1946.945 ;
        RECT 2401.865 1946.245 2402.905 1946.385 ;
        RECT 2401.865 1946.155 2402.125 1946.245 ;
        RECT 2402.765 1946.005 2402.905 1946.245 ;
        RECT 2403.345 1946.245 2403.905 1946.385 ;
        RECT 2403.345 1946.155 2403.605 1946.245 ;
        RECT 2404.065 1946.155 2404.325 1946.475 ;
        RECT 2404.785 1946.155 2405.045 1946.475 ;
        RECT 2405.205 1946.005 2405.345 1946.805 ;
        RECT 2405.785 1946.715 2406.045 1946.805 ;
        RECT 2406.325 1946.475 2406.465 1947.835 ;
        RECT 2406.745 1947.785 2406.945 1947.835 ;
        RECT 2407.215 1947.805 2407.495 1948.180 ;
        RECT 2408.215 1947.805 2408.495 1948.180 ;
        RECT 2411.215 1947.795 2411.405 1948.430 ;
        RECT 2406.685 1947.615 2406.945 1947.785 ;
        RECT 2406.685 1947.245 2407.185 1947.615 ;
        RECT 2407.745 1947.275 2408.005 1947.595 ;
        RECT 2411.145 1947.445 2411.485 1947.795 ;
        RECT 2411.235 1947.440 2411.405 1947.445 ;
        RECT 2406.685 1946.475 2406.825 1947.245 ;
        RECT 2407.805 1946.475 2407.945 1947.275 ;
        RECT 2412.435 1946.860 2412.595 1952.035 ;
        RECT 2413.550 1951.945 2413.875 1952.035 ;
        RECT 2415.885 1952.175 2416.235 1952.295 ;
        RECT 2426.670 1952.175 2427.020 1952.250 ;
        RECT 2432.110 1952.205 2432.435 1952.270 ;
        RECT 2415.885 1951.975 2427.020 1952.175 ;
        RECT 2415.885 1951.945 2416.235 1951.975 ;
        RECT 2426.670 1951.900 2427.020 1951.975 ;
        RECT 2430.995 1952.035 2432.435 1952.205 ;
        RECT 2412.750 1951.510 2413.070 1951.835 ;
        RECT 2412.780 1951.335 2412.950 1951.510 ;
        RECT 2412.780 1951.160 2412.955 1951.335 ;
        RECT 2412.780 1950.985 2413.755 1951.160 ;
        RECT 2412.750 1946.860 2413.070 1946.980 ;
        RECT 2412.435 1946.690 2413.070 1946.860 ;
        RECT 2412.750 1946.660 2413.070 1946.690 ;
        RECT 2413.580 1946.610 2413.755 1950.985 ;
        RECT 2425.830 1948.430 2429.965 1948.620 ;
        RECT 2425.830 1948.180 2426.020 1948.430 ;
        RECT 2417.495 1947.805 2417.775 1948.180 ;
        RECT 2422.265 1947.835 2422.525 1948.155 ;
        RECT 2417.505 1947.555 2417.765 1947.805 ;
        RECT 2419.935 1947.595 2420.215 1947.620 ;
        RECT 2418.465 1947.275 2418.725 1947.595 ;
        RECT 2419.585 1947.505 2420.215 1947.595 ;
        RECT 2421.905 1947.505 2422.165 1947.595 ;
        RECT 2419.585 1947.365 2422.165 1947.505 ;
        RECT 2419.585 1947.275 2420.215 1947.365 ;
        RECT 2421.905 1947.275 2422.165 1947.365 ;
        RECT 2417.975 1946.685 2418.255 1947.060 ;
        RECT 2406.025 1946.245 2406.465 1946.475 ;
        RECT 2406.025 1946.155 2406.285 1946.245 ;
        RECT 2406.625 1946.155 2406.885 1946.475 ;
        RECT 2407.745 1946.155 2408.005 1946.475 ;
        RECT 2409.175 1946.125 2409.455 1946.500 ;
        RECT 2413.525 1946.260 2413.875 1946.610 ;
        RECT 2418.525 1946.475 2418.665 1947.275 ;
        RECT 2419.935 1947.245 2420.215 1947.275 ;
        RECT 2421.375 1947.035 2421.655 1947.060 ;
        RECT 2421.375 1946.715 2421.905 1947.035 ;
        RECT 2421.375 1946.685 2421.655 1946.715 ;
        RECT 2418.465 1946.155 2418.725 1946.475 ;
        RECT 2420.425 1946.385 2420.685 1946.475 ;
        RECT 2421.905 1946.385 2422.165 1946.475 ;
        RECT 2422.325 1946.385 2422.465 1947.835 ;
        RECT 2423.815 1947.805 2424.095 1948.180 ;
        RECT 2424.825 1947.835 2425.085 1948.155 ;
        RECT 2425.305 1947.835 2425.565 1948.155 ;
        RECT 2422.615 1947.245 2422.895 1947.620 ;
        RECT 2423.885 1947.615 2424.025 1947.805 ;
        RECT 2423.695 1947.505 2424.025 1947.615 ;
        RECT 2423.405 1947.365 2424.025 1947.505 ;
        RECT 2422.685 1946.475 2422.825 1947.245 ;
        RECT 2423.405 1946.475 2423.545 1947.365 ;
        RECT 2423.695 1947.245 2423.975 1947.365 ;
        RECT 2424.345 1946.945 2424.605 1947.035 ;
        RECT 2423.765 1946.805 2424.605 1946.945 ;
        RECT 2420.425 1946.245 2421.465 1946.385 ;
        RECT 2420.425 1946.155 2420.685 1946.245 ;
        RECT 2402.765 1945.865 2405.345 1946.005 ;
        RECT 2421.325 1946.005 2421.465 1946.245 ;
        RECT 2421.905 1946.245 2422.465 1946.385 ;
        RECT 2421.905 1946.155 2422.165 1946.245 ;
        RECT 2422.625 1946.155 2422.885 1946.475 ;
        RECT 2423.345 1946.155 2423.605 1946.475 ;
        RECT 2423.765 1946.005 2423.905 1946.805 ;
        RECT 2424.345 1946.715 2424.605 1946.805 ;
        RECT 2424.885 1946.475 2425.025 1947.835 ;
        RECT 2425.305 1947.785 2425.505 1947.835 ;
        RECT 2425.775 1947.805 2426.055 1948.180 ;
        RECT 2426.775 1947.805 2427.055 1948.180 ;
        RECT 2429.775 1947.795 2429.965 1948.430 ;
        RECT 2425.245 1947.615 2425.505 1947.785 ;
        RECT 2425.245 1947.245 2425.745 1947.615 ;
        RECT 2426.305 1947.275 2426.565 1947.595 ;
        RECT 2429.705 1947.445 2430.045 1947.795 ;
        RECT 2429.795 1947.440 2429.965 1947.445 ;
        RECT 2425.245 1946.475 2425.385 1947.245 ;
        RECT 2426.365 1946.475 2426.505 1947.275 ;
        RECT 2430.995 1946.860 2431.155 1952.035 ;
        RECT 2432.110 1951.945 2432.435 1952.035 ;
        RECT 2434.445 1952.175 2434.795 1952.295 ;
        RECT 2445.230 1952.175 2445.580 1952.250 ;
        RECT 2450.670 1952.205 2450.995 1952.270 ;
        RECT 2434.445 1951.975 2445.580 1952.175 ;
        RECT 2434.445 1951.945 2434.795 1951.975 ;
        RECT 2445.230 1951.900 2445.580 1951.975 ;
        RECT 2449.555 1952.035 2450.995 1952.205 ;
        RECT 2431.310 1951.510 2431.630 1951.835 ;
        RECT 2431.340 1951.335 2431.510 1951.510 ;
        RECT 2431.340 1951.160 2431.515 1951.335 ;
        RECT 2431.340 1950.985 2432.315 1951.160 ;
        RECT 2431.310 1946.860 2431.630 1946.980 ;
        RECT 2430.995 1946.690 2431.630 1946.860 ;
        RECT 2431.310 1946.660 2431.630 1946.690 ;
        RECT 2432.140 1946.610 2432.315 1950.985 ;
        RECT 2444.390 1948.430 2448.525 1948.620 ;
        RECT 2444.390 1948.180 2444.580 1948.430 ;
        RECT 2436.055 1947.805 2436.335 1948.180 ;
        RECT 2440.825 1947.835 2441.085 1948.155 ;
        RECT 2436.065 1947.555 2436.325 1947.805 ;
        RECT 2438.495 1947.595 2438.775 1947.620 ;
        RECT 2437.025 1947.275 2437.285 1947.595 ;
        RECT 2438.145 1947.505 2438.775 1947.595 ;
        RECT 2440.465 1947.505 2440.725 1947.595 ;
        RECT 2438.145 1947.365 2440.725 1947.505 ;
        RECT 2438.145 1947.275 2438.775 1947.365 ;
        RECT 2440.465 1947.275 2440.725 1947.365 ;
        RECT 2436.535 1946.685 2436.815 1947.060 ;
        RECT 2424.585 1946.245 2425.025 1946.475 ;
        RECT 2424.585 1946.155 2424.845 1946.245 ;
        RECT 2425.185 1946.155 2425.445 1946.475 ;
        RECT 2426.305 1946.155 2426.565 1946.475 ;
        RECT 2427.735 1946.125 2428.015 1946.500 ;
        RECT 2432.085 1946.260 2432.435 1946.610 ;
        RECT 2437.085 1946.475 2437.225 1947.275 ;
        RECT 2438.495 1947.245 2438.775 1947.275 ;
        RECT 2439.935 1947.035 2440.215 1947.060 ;
        RECT 2439.935 1946.715 2440.465 1947.035 ;
        RECT 2439.935 1946.685 2440.215 1946.715 ;
        RECT 2437.025 1946.155 2437.285 1946.475 ;
        RECT 2438.985 1946.385 2439.245 1946.475 ;
        RECT 2440.465 1946.385 2440.725 1946.475 ;
        RECT 2440.885 1946.385 2441.025 1947.835 ;
        RECT 2442.375 1947.805 2442.655 1948.180 ;
        RECT 2443.385 1947.835 2443.645 1948.155 ;
        RECT 2443.865 1947.835 2444.125 1948.155 ;
        RECT 2441.175 1947.245 2441.455 1947.620 ;
        RECT 2442.445 1947.615 2442.585 1947.805 ;
        RECT 2442.255 1947.505 2442.585 1947.615 ;
        RECT 2441.965 1947.365 2442.585 1947.505 ;
        RECT 2441.245 1946.475 2441.385 1947.245 ;
        RECT 2441.965 1946.475 2442.105 1947.365 ;
        RECT 2442.255 1947.245 2442.535 1947.365 ;
        RECT 2442.905 1946.945 2443.165 1947.035 ;
        RECT 2442.325 1946.805 2443.165 1946.945 ;
        RECT 2438.985 1946.245 2440.025 1946.385 ;
        RECT 2438.985 1946.155 2439.245 1946.245 ;
        RECT 2421.325 1945.865 2423.905 1946.005 ;
        RECT 2439.885 1946.005 2440.025 1946.245 ;
        RECT 2440.465 1946.245 2441.025 1946.385 ;
        RECT 2440.465 1946.155 2440.725 1946.245 ;
        RECT 2441.185 1946.155 2441.445 1946.475 ;
        RECT 2441.905 1946.155 2442.165 1946.475 ;
        RECT 2442.325 1946.005 2442.465 1946.805 ;
        RECT 2442.905 1946.715 2443.165 1946.805 ;
        RECT 2443.445 1946.475 2443.585 1947.835 ;
        RECT 2443.865 1947.785 2444.065 1947.835 ;
        RECT 2444.335 1947.805 2444.615 1948.180 ;
        RECT 2445.335 1947.805 2445.615 1948.180 ;
        RECT 2448.335 1947.795 2448.525 1948.430 ;
        RECT 2443.805 1947.615 2444.065 1947.785 ;
        RECT 2443.805 1947.245 2444.305 1947.615 ;
        RECT 2444.865 1947.275 2445.125 1947.595 ;
        RECT 2448.265 1947.445 2448.605 1947.795 ;
        RECT 2448.355 1947.440 2448.525 1947.445 ;
        RECT 2443.805 1946.475 2443.945 1947.245 ;
        RECT 2444.925 1946.475 2445.065 1947.275 ;
        RECT 2449.555 1946.860 2449.715 1952.035 ;
        RECT 2450.670 1951.945 2450.995 1952.035 ;
        RECT 2449.870 1951.510 2450.190 1951.835 ;
        RECT 2449.900 1951.335 2450.070 1951.510 ;
        RECT 2449.900 1951.160 2450.075 1951.335 ;
        RECT 2449.900 1950.985 2450.875 1951.160 ;
        RECT 2449.870 1946.860 2450.190 1946.980 ;
        RECT 2449.555 1946.690 2450.190 1946.860 ;
        RECT 2449.870 1946.660 2450.190 1946.690 ;
        RECT 2450.700 1946.610 2450.875 1950.985 ;
        RECT 2443.145 1946.245 2443.585 1946.475 ;
        RECT 2443.145 1946.155 2443.405 1946.245 ;
        RECT 2443.745 1946.155 2444.005 1946.475 ;
        RECT 2444.865 1946.155 2445.125 1946.475 ;
        RECT 2446.295 1946.125 2446.575 1946.500 ;
        RECT 2450.645 1946.260 2450.995 1946.610 ;
        RECT 2439.885 1945.865 2442.465 1946.005 ;
        RECT 2416.020 1945.150 2416.280 1945.470 ;
        RECT 2434.420 1945.150 2434.680 1945.470 ;
        RECT 2378.760 1938.690 2379.020 1939.010 ;
        RECT 2397.160 1938.690 2397.420 1939.010 ;
        RECT 2416.080 1932.210 2416.220 1945.150 ;
        RECT 2434.480 1932.405 2434.620 1945.150 ;
        RECT 2416.020 1931.890 2416.280 1932.210 ;
        RECT 2421.540 1931.890 2421.800 1932.210 ;
        RECT 2434.410 1932.035 2434.690 1932.405 ;
        RECT 2421.600 1849.250 2421.740 1931.890 ;
        RECT 2421.540 1848.930 2421.800 1849.250 ;
        RECT 2369.175 1790.690 2446.675 1790.860 ;
        RECT 2369.175 1788.895 2369.345 1790.690 ;
        RECT 2446.505 1789.915 2446.675 1790.690 ;
        RECT 2369.490 1789.530 2369.780 1789.640 ;
        RECT 2369.490 1789.525 2369.810 1789.530 ;
        RECT 2369.490 1789.355 2370.710 1789.525 ;
        RECT 2369.490 1789.290 2369.780 1789.355 ;
        RECT 2370.540 1789.145 2370.710 1789.355 ;
        RECT 2376.965 1789.345 2377.335 1789.715 ;
        RECT 2392.225 1789.345 2392.595 1789.715 ;
        RECT 2407.485 1789.345 2407.855 1789.715 ;
        RECT 2422.745 1789.345 2423.115 1789.715 ;
        RECT 2438.005 1789.345 2438.375 1789.715 ;
        RECT 2446.475 1789.565 2446.825 1789.915 ;
        RECT 2377.635 1789.145 2377.985 1789.245 ;
        RECT 2383.075 1789.205 2383.400 1789.270 ;
        RECT 2370.540 1788.975 2377.985 1789.145 ;
        RECT 2377.635 1788.895 2377.985 1788.975 ;
        RECT 2381.960 1789.035 2383.400 1789.205 ;
        RECT 2369.115 1788.545 2369.405 1788.895 ;
        RECT 2374.935 1785.305 2377.375 1785.445 ;
        RECT 2374.935 1785.155 2375.075 1785.305 ;
        RECT 2374.635 1785.065 2375.075 1785.155 ;
        RECT 2372.295 1784.925 2375.075 1785.065 ;
        RECT 2371.785 1784.785 2372.045 1784.875 ;
        RECT 2372.295 1784.785 2372.435 1784.925 ;
        RECT 2374.635 1784.835 2374.895 1784.925 ;
        RECT 2375.235 1784.835 2375.495 1785.155 ;
        RECT 2375.235 1784.785 2375.435 1784.835 ;
        RECT 2371.785 1784.645 2372.435 1784.785 ;
        RECT 2375.045 1784.645 2375.435 1784.785 ;
        RECT 2376.305 1784.775 2376.585 1785.155 ;
        RECT 2376.795 1784.835 2377.070 1785.155 ;
        RECT 2371.785 1784.555 2372.045 1784.645 ;
        RECT 2371.845 1783.475 2371.985 1784.555 ;
        RECT 2372.705 1784.505 2372.985 1784.620 ;
        RECT 2374.155 1784.505 2374.415 1784.595 ;
        RECT 2372.535 1784.365 2374.415 1784.505 ;
        RECT 2372.535 1784.315 2372.985 1784.365 ;
        RECT 2372.475 1784.245 2372.985 1784.315 ;
        RECT 2374.155 1784.275 2374.415 1784.365 ;
        RECT 2372.475 1784.055 2372.735 1784.245 ;
        RECT 2373.650 1784.055 2373.955 1784.060 ;
        RECT 2372.465 1783.685 2372.745 1784.055 ;
        RECT 2372.955 1783.945 2373.215 1784.035 ;
        RECT 2373.545 1783.945 2373.955 1784.055 ;
        RECT 2372.955 1783.805 2373.955 1783.945 ;
        RECT 2372.955 1783.715 2373.215 1783.805 ;
        RECT 2373.545 1783.685 2373.955 1783.805 ;
        RECT 2374.385 1783.685 2374.665 1784.060 ;
        RECT 2375.045 1783.525 2375.185 1784.645 ;
        RECT 2376.375 1784.315 2376.515 1784.775 ;
        RECT 2375.825 1783.685 2376.105 1784.155 ;
        RECT 2376.315 1784.055 2376.575 1784.315 ;
        RECT 2376.305 1783.685 2376.585 1784.055 ;
        RECT 2375.045 1783.475 2375.355 1783.525 ;
        RECT 2376.855 1783.515 2376.995 1784.835 ;
        RECT 2377.235 1784.315 2377.375 1785.305 ;
        RECT 2377.545 1784.555 2377.805 1784.875 ;
        RECT 2379.405 1784.835 2379.665 1785.155 ;
        RECT 2377.175 1783.995 2377.435 1784.315 ;
        RECT 2377.605 1783.515 2377.745 1784.555 ;
        RECT 2379.465 1784.055 2379.605 1784.835 ;
        RECT 2380.670 1784.265 2381.010 1784.345 ;
        RECT 2378.715 1783.945 2378.975 1784.035 ;
        RECT 2378.055 1783.805 2378.975 1783.945 ;
        RECT 2376.515 1783.495 2376.995 1783.515 ;
        RECT 2371.785 1783.155 2372.045 1783.475 ;
        RECT 2374.515 1783.385 2374.775 1783.475 ;
        RECT 2374.985 1783.445 2375.355 1783.475 ;
        RECT 2374.515 1783.155 2374.835 1783.385 ;
        RECT 2374.695 1783.005 2374.835 1783.155 ;
        RECT 2374.985 1783.150 2375.395 1783.445 ;
        RECT 2375.585 1783.155 2375.865 1783.495 ;
        RECT 2376.315 1783.245 2376.995 1783.495 ;
        RECT 2377.535 1783.445 2377.815 1783.515 ;
        RECT 2376.315 1783.145 2376.795 1783.245 ;
        RECT 2377.485 1783.185 2377.860 1783.445 ;
        RECT 2377.535 1783.145 2377.815 1783.185 ;
        RECT 2378.055 1783.005 2378.195 1783.805 ;
        RECT 2378.715 1783.715 2378.975 1783.805 ;
        RECT 2379.295 1783.685 2379.605 1784.055 ;
        RECT 2379.365 1783.500 2379.605 1783.685 ;
        RECT 2380.045 1784.065 2381.010 1784.265 ;
        RECT 2379.365 1783.435 2379.675 1783.500 ;
        RECT 2380.045 1783.435 2380.245 1784.065 ;
        RECT 2380.670 1783.995 2381.010 1784.065 ;
        RECT 2380.760 1783.990 2380.930 1783.995 ;
        RECT 2381.960 1783.860 2382.120 1789.035 ;
        RECT 2383.075 1788.945 2383.400 1789.035 ;
        RECT 2385.455 1789.180 2385.805 1789.300 ;
        RECT 2392.895 1789.180 2393.245 1789.255 ;
        RECT 2398.335 1789.205 2398.660 1789.270 ;
        RECT 2385.455 1788.980 2393.245 1789.180 ;
        RECT 2385.455 1788.950 2385.805 1788.980 ;
        RECT 2392.895 1788.905 2393.245 1788.980 ;
        RECT 2397.220 1789.035 2398.660 1789.205 ;
        RECT 2382.275 1788.510 2382.595 1788.835 ;
        RECT 2382.305 1788.335 2382.475 1788.510 ;
        RECT 2382.305 1788.160 2382.480 1788.335 ;
        RECT 2382.305 1787.985 2383.280 1788.160 ;
        RECT 2382.275 1783.860 2382.595 1783.980 ;
        RECT 2381.960 1783.690 2382.595 1783.860 ;
        RECT 2382.275 1783.660 2382.595 1783.690 ;
        RECT 2383.105 1783.610 2383.280 1787.985 ;
        RECT 2390.195 1785.305 2392.635 1785.445 ;
        RECT 2390.195 1785.155 2390.335 1785.305 ;
        RECT 2389.895 1785.065 2390.335 1785.155 ;
        RECT 2387.555 1784.925 2390.335 1785.065 ;
        RECT 2387.045 1784.785 2387.305 1784.875 ;
        RECT 2387.555 1784.785 2387.695 1784.925 ;
        RECT 2389.895 1784.835 2390.155 1784.925 ;
        RECT 2390.495 1784.835 2390.755 1785.155 ;
        RECT 2390.495 1784.785 2390.695 1784.835 ;
        RECT 2387.045 1784.645 2387.695 1784.785 ;
        RECT 2390.305 1784.645 2390.695 1784.785 ;
        RECT 2391.565 1784.775 2391.845 1785.155 ;
        RECT 2392.055 1784.835 2392.330 1785.155 ;
        RECT 2387.045 1784.555 2387.305 1784.645 ;
        RECT 2385.200 1783.990 2385.460 1784.310 ;
        RECT 2379.365 1783.245 2380.245 1783.435 ;
        RECT 2383.050 1783.260 2383.400 1783.610 ;
        RECT 2379.395 1783.235 2380.245 1783.245 ;
        RECT 2379.395 1783.125 2379.675 1783.235 ;
        RECT 2374.695 1782.865 2378.195 1783.005 ;
        RECT 2385.260 1773.370 2385.400 1783.990 ;
        RECT 2387.105 1783.475 2387.245 1784.555 ;
        RECT 2387.965 1784.505 2388.245 1784.620 ;
        RECT 2389.415 1784.505 2389.675 1784.595 ;
        RECT 2387.795 1784.365 2389.675 1784.505 ;
        RECT 2387.795 1784.315 2388.245 1784.365 ;
        RECT 2387.735 1784.245 2388.245 1784.315 ;
        RECT 2389.415 1784.275 2389.675 1784.365 ;
        RECT 2387.735 1784.055 2387.995 1784.245 ;
        RECT 2388.910 1784.055 2389.215 1784.060 ;
        RECT 2387.725 1783.685 2388.005 1784.055 ;
        RECT 2388.215 1783.945 2388.475 1784.035 ;
        RECT 2388.805 1783.945 2389.215 1784.055 ;
        RECT 2388.215 1783.805 2389.215 1783.945 ;
        RECT 2388.215 1783.715 2388.475 1783.805 ;
        RECT 2388.805 1783.685 2389.215 1783.805 ;
        RECT 2389.645 1783.685 2389.925 1784.060 ;
        RECT 2390.305 1783.525 2390.445 1784.645 ;
        RECT 2391.635 1784.315 2391.775 1784.775 ;
        RECT 2391.085 1783.685 2391.365 1784.155 ;
        RECT 2391.575 1784.055 2391.835 1784.315 ;
        RECT 2391.565 1783.685 2391.845 1784.055 ;
        RECT 2390.305 1783.475 2390.615 1783.525 ;
        RECT 2392.115 1783.515 2392.255 1784.835 ;
        RECT 2392.495 1784.315 2392.635 1785.305 ;
        RECT 2392.805 1784.555 2393.065 1784.875 ;
        RECT 2394.665 1784.835 2394.925 1785.155 ;
        RECT 2392.435 1783.995 2392.695 1784.315 ;
        RECT 2392.865 1783.515 2393.005 1784.555 ;
        RECT 2394.725 1784.055 2394.865 1784.835 ;
        RECT 2395.930 1784.265 2396.270 1784.345 ;
        RECT 2393.975 1783.945 2394.235 1784.035 ;
        RECT 2393.315 1783.805 2394.235 1783.945 ;
        RECT 2391.775 1783.495 2392.255 1783.515 ;
        RECT 2387.045 1783.155 2387.305 1783.475 ;
        RECT 2389.775 1783.385 2390.035 1783.475 ;
        RECT 2390.245 1783.445 2390.615 1783.475 ;
        RECT 2389.775 1783.155 2390.095 1783.385 ;
        RECT 2389.955 1783.005 2390.095 1783.155 ;
        RECT 2390.245 1783.150 2390.655 1783.445 ;
        RECT 2390.845 1783.155 2391.125 1783.495 ;
        RECT 2391.575 1783.245 2392.255 1783.495 ;
        RECT 2392.795 1783.445 2393.075 1783.515 ;
        RECT 2391.575 1783.145 2392.055 1783.245 ;
        RECT 2392.745 1783.185 2393.120 1783.445 ;
        RECT 2392.795 1783.145 2393.075 1783.185 ;
        RECT 2393.315 1783.005 2393.455 1783.805 ;
        RECT 2393.975 1783.715 2394.235 1783.805 ;
        RECT 2394.555 1783.685 2394.865 1784.055 ;
        RECT 2394.625 1783.500 2394.865 1783.685 ;
        RECT 2395.305 1784.065 2396.270 1784.265 ;
        RECT 2394.625 1783.435 2394.935 1783.500 ;
        RECT 2395.305 1783.435 2395.505 1784.065 ;
        RECT 2395.930 1783.995 2396.270 1784.065 ;
        RECT 2396.020 1783.990 2396.190 1783.995 ;
        RECT 2397.220 1783.860 2397.380 1789.035 ;
        RECT 2398.335 1788.945 2398.660 1789.035 ;
        RECT 2400.715 1789.180 2401.065 1789.300 ;
        RECT 2408.155 1789.180 2408.505 1789.255 ;
        RECT 2413.595 1789.205 2413.920 1789.270 ;
        RECT 2400.715 1788.980 2408.505 1789.180 ;
        RECT 2400.715 1788.950 2401.065 1788.980 ;
        RECT 2408.155 1788.905 2408.505 1788.980 ;
        RECT 2412.480 1789.035 2413.920 1789.205 ;
        RECT 2397.535 1788.510 2397.855 1788.835 ;
        RECT 2397.565 1788.335 2397.735 1788.510 ;
        RECT 2397.565 1788.160 2397.740 1788.335 ;
        RECT 2397.565 1787.985 2398.540 1788.160 ;
        RECT 2397.535 1783.860 2397.855 1783.980 ;
        RECT 2397.220 1783.690 2397.855 1783.860 ;
        RECT 2397.535 1783.660 2397.855 1783.690 ;
        RECT 2398.365 1783.610 2398.540 1787.985 ;
        RECT 2405.455 1785.305 2407.895 1785.445 ;
        RECT 2405.455 1785.155 2405.595 1785.305 ;
        RECT 2405.155 1785.065 2405.595 1785.155 ;
        RECT 2402.815 1784.925 2405.595 1785.065 ;
        RECT 2402.305 1784.785 2402.565 1784.875 ;
        RECT 2402.815 1784.785 2402.955 1784.925 ;
        RECT 2405.155 1784.835 2405.415 1784.925 ;
        RECT 2405.755 1784.835 2406.015 1785.155 ;
        RECT 2405.755 1784.785 2405.955 1784.835 ;
        RECT 2402.305 1784.645 2402.955 1784.785 ;
        RECT 2405.565 1784.645 2405.955 1784.785 ;
        RECT 2406.825 1784.775 2407.105 1785.155 ;
        RECT 2407.315 1784.835 2407.590 1785.155 ;
        RECT 2402.305 1784.555 2402.565 1784.645 ;
        RECT 2400.840 1783.990 2401.100 1784.310 ;
        RECT 2394.625 1783.245 2395.505 1783.435 ;
        RECT 2398.310 1783.260 2398.660 1783.610 ;
        RECT 2394.655 1783.235 2395.505 1783.245 ;
        RECT 2394.655 1783.125 2394.935 1783.235 ;
        RECT 2389.955 1782.865 2393.455 1783.005 ;
        RECT 2385.260 1773.230 2385.860 1773.370 ;
        RECT 2385.720 1772.750 2385.860 1773.230 ;
        RECT 2400.900 1773.090 2401.040 1783.990 ;
        RECT 2402.365 1783.475 2402.505 1784.555 ;
        RECT 2403.225 1784.505 2403.505 1784.620 ;
        RECT 2404.675 1784.505 2404.935 1784.595 ;
        RECT 2403.055 1784.365 2404.935 1784.505 ;
        RECT 2403.055 1784.315 2403.505 1784.365 ;
        RECT 2402.995 1784.245 2403.505 1784.315 ;
        RECT 2404.675 1784.275 2404.935 1784.365 ;
        RECT 2402.995 1784.055 2403.255 1784.245 ;
        RECT 2404.170 1784.055 2404.475 1784.060 ;
        RECT 2402.985 1783.685 2403.265 1784.055 ;
        RECT 2403.475 1783.945 2403.735 1784.035 ;
        RECT 2404.065 1783.945 2404.475 1784.055 ;
        RECT 2403.475 1783.805 2404.475 1783.945 ;
        RECT 2403.475 1783.715 2403.735 1783.805 ;
        RECT 2404.065 1783.685 2404.475 1783.805 ;
        RECT 2404.905 1783.685 2405.185 1784.060 ;
        RECT 2405.565 1783.525 2405.705 1784.645 ;
        RECT 2406.895 1784.315 2407.035 1784.775 ;
        RECT 2406.345 1783.685 2406.625 1784.155 ;
        RECT 2406.835 1784.055 2407.095 1784.315 ;
        RECT 2406.825 1783.685 2407.105 1784.055 ;
        RECT 2405.565 1783.475 2405.875 1783.525 ;
        RECT 2407.375 1783.515 2407.515 1784.835 ;
        RECT 2407.755 1784.315 2407.895 1785.305 ;
        RECT 2408.065 1784.555 2408.325 1784.875 ;
        RECT 2409.925 1784.835 2410.185 1785.155 ;
        RECT 2407.695 1783.995 2407.955 1784.315 ;
        RECT 2408.125 1783.515 2408.265 1784.555 ;
        RECT 2409.985 1784.055 2410.125 1784.835 ;
        RECT 2411.190 1784.265 2411.530 1784.345 ;
        RECT 2409.235 1783.945 2409.495 1784.035 ;
        RECT 2408.575 1783.805 2409.495 1783.945 ;
        RECT 2407.035 1783.495 2407.515 1783.515 ;
        RECT 2402.305 1783.155 2402.565 1783.475 ;
        RECT 2405.035 1783.385 2405.295 1783.475 ;
        RECT 2405.505 1783.445 2405.875 1783.475 ;
        RECT 2405.035 1783.155 2405.355 1783.385 ;
        RECT 2405.215 1783.005 2405.355 1783.155 ;
        RECT 2405.505 1783.150 2405.915 1783.445 ;
        RECT 2406.105 1783.155 2406.385 1783.495 ;
        RECT 2406.835 1783.245 2407.515 1783.495 ;
        RECT 2408.055 1783.445 2408.335 1783.515 ;
        RECT 2406.835 1783.145 2407.315 1783.245 ;
        RECT 2408.005 1783.185 2408.380 1783.445 ;
        RECT 2408.055 1783.145 2408.335 1783.185 ;
        RECT 2408.575 1783.005 2408.715 1783.805 ;
        RECT 2409.235 1783.715 2409.495 1783.805 ;
        RECT 2409.815 1783.685 2410.125 1784.055 ;
        RECT 2409.885 1783.500 2410.125 1783.685 ;
        RECT 2410.565 1784.065 2411.530 1784.265 ;
        RECT 2409.885 1783.435 2410.195 1783.500 ;
        RECT 2410.565 1783.435 2410.765 1784.065 ;
        RECT 2411.190 1783.995 2411.530 1784.065 ;
        RECT 2411.280 1783.990 2411.450 1783.995 ;
        RECT 2412.480 1783.860 2412.640 1789.035 ;
        RECT 2413.595 1788.945 2413.920 1789.035 ;
        RECT 2415.930 1789.180 2416.280 1789.300 ;
        RECT 2423.420 1789.180 2423.770 1789.255 ;
        RECT 2428.855 1789.205 2429.180 1789.270 ;
        RECT 2415.930 1788.980 2423.770 1789.180 ;
        RECT 2415.930 1788.950 2416.280 1788.980 ;
        RECT 2423.420 1788.905 2423.770 1788.980 ;
        RECT 2427.740 1789.035 2429.180 1789.205 ;
        RECT 2412.795 1788.510 2413.115 1788.835 ;
        RECT 2412.825 1788.335 2412.995 1788.510 ;
        RECT 2412.825 1788.160 2413.000 1788.335 ;
        RECT 2412.825 1787.985 2413.800 1788.160 ;
        RECT 2412.795 1783.860 2413.115 1783.980 ;
        RECT 2412.480 1783.690 2413.115 1783.860 ;
        RECT 2412.795 1783.660 2413.115 1783.690 ;
        RECT 2413.625 1783.610 2413.800 1787.985 ;
        RECT 2420.715 1785.305 2423.155 1785.445 ;
        RECT 2420.715 1785.155 2420.855 1785.305 ;
        RECT 2420.415 1785.065 2420.855 1785.155 ;
        RECT 2418.075 1784.925 2420.855 1785.065 ;
        RECT 2417.565 1784.785 2417.825 1784.875 ;
        RECT 2418.075 1784.785 2418.215 1784.925 ;
        RECT 2420.415 1784.835 2420.675 1784.925 ;
        RECT 2421.015 1784.835 2421.275 1785.155 ;
        RECT 2421.015 1784.785 2421.215 1784.835 ;
        RECT 2417.565 1784.645 2418.215 1784.785 ;
        RECT 2420.825 1784.645 2421.215 1784.785 ;
        RECT 2422.085 1784.775 2422.365 1785.155 ;
        RECT 2422.575 1784.835 2422.850 1785.155 ;
        RECT 2417.565 1784.555 2417.825 1784.645 ;
        RECT 2409.885 1783.245 2410.765 1783.435 ;
        RECT 2413.570 1783.260 2413.920 1783.610 ;
        RECT 2417.625 1783.475 2417.765 1784.555 ;
        RECT 2418.485 1784.505 2418.765 1784.620 ;
        RECT 2419.935 1784.505 2420.195 1784.595 ;
        RECT 2418.315 1784.365 2420.195 1784.505 ;
        RECT 2418.315 1784.315 2418.765 1784.365 ;
        RECT 2418.255 1784.245 2418.765 1784.315 ;
        RECT 2419.935 1784.275 2420.195 1784.365 ;
        RECT 2418.255 1784.055 2418.515 1784.245 ;
        RECT 2419.430 1784.055 2419.735 1784.060 ;
        RECT 2418.245 1783.685 2418.525 1784.055 ;
        RECT 2418.735 1783.945 2418.995 1784.035 ;
        RECT 2419.325 1783.945 2419.735 1784.055 ;
        RECT 2418.735 1783.805 2419.735 1783.945 ;
        RECT 2418.735 1783.715 2418.995 1783.805 ;
        RECT 2419.325 1783.685 2419.735 1783.805 ;
        RECT 2420.165 1783.685 2420.445 1784.060 ;
        RECT 2420.825 1783.525 2420.965 1784.645 ;
        RECT 2422.155 1784.315 2422.295 1784.775 ;
        RECT 2421.605 1783.685 2421.885 1784.155 ;
        RECT 2422.095 1784.055 2422.355 1784.315 ;
        RECT 2422.085 1783.685 2422.365 1784.055 ;
        RECT 2420.825 1783.475 2421.135 1783.525 ;
        RECT 2422.635 1783.515 2422.775 1784.835 ;
        RECT 2423.015 1784.315 2423.155 1785.305 ;
        RECT 2423.325 1784.555 2423.585 1784.875 ;
        RECT 2425.185 1784.835 2425.445 1785.155 ;
        RECT 2422.955 1783.995 2423.215 1784.315 ;
        RECT 2423.385 1783.515 2423.525 1784.555 ;
        RECT 2425.245 1784.055 2425.385 1784.835 ;
        RECT 2426.450 1784.265 2426.790 1784.345 ;
        RECT 2424.495 1783.945 2424.755 1784.035 ;
        RECT 2423.835 1783.805 2424.755 1783.945 ;
        RECT 2422.295 1783.495 2422.775 1783.515 ;
        RECT 2409.915 1783.235 2410.765 1783.245 ;
        RECT 2409.915 1783.125 2410.195 1783.235 ;
        RECT 2417.565 1783.155 2417.825 1783.475 ;
        RECT 2420.295 1783.385 2420.555 1783.475 ;
        RECT 2420.765 1783.445 2421.135 1783.475 ;
        RECT 2420.295 1783.155 2420.615 1783.385 ;
        RECT 2405.215 1782.865 2408.715 1783.005 ;
        RECT 2420.475 1783.005 2420.615 1783.155 ;
        RECT 2420.765 1783.150 2421.175 1783.445 ;
        RECT 2421.365 1783.155 2421.645 1783.495 ;
        RECT 2422.095 1783.245 2422.775 1783.495 ;
        RECT 2423.315 1783.445 2423.595 1783.515 ;
        RECT 2422.095 1783.145 2422.575 1783.245 ;
        RECT 2423.265 1783.185 2423.640 1783.445 ;
        RECT 2423.315 1783.145 2423.595 1783.185 ;
        RECT 2423.835 1783.005 2423.975 1783.805 ;
        RECT 2424.495 1783.715 2424.755 1783.805 ;
        RECT 2425.075 1783.685 2425.385 1784.055 ;
        RECT 2425.145 1783.500 2425.385 1783.685 ;
        RECT 2425.825 1784.065 2426.790 1784.265 ;
        RECT 2425.145 1783.435 2425.455 1783.500 ;
        RECT 2425.825 1783.435 2426.025 1784.065 ;
        RECT 2426.450 1783.995 2426.790 1784.065 ;
        RECT 2426.540 1783.990 2426.710 1783.995 ;
        RECT 2427.740 1783.860 2427.900 1789.035 ;
        RECT 2428.855 1788.945 2429.180 1789.035 ;
        RECT 2431.190 1789.180 2431.540 1789.300 ;
        RECT 2438.675 1789.180 2439.025 1789.255 ;
        RECT 2444.115 1789.205 2444.440 1789.270 ;
        RECT 2431.190 1788.980 2439.025 1789.180 ;
        RECT 2431.190 1788.950 2431.540 1788.980 ;
        RECT 2438.675 1788.905 2439.025 1788.980 ;
        RECT 2443.000 1789.035 2444.440 1789.205 ;
        RECT 2428.055 1788.510 2428.375 1788.835 ;
        RECT 2428.085 1788.335 2428.255 1788.510 ;
        RECT 2428.085 1788.160 2428.260 1788.335 ;
        RECT 2428.085 1787.985 2429.060 1788.160 ;
        RECT 2428.055 1783.860 2428.375 1783.980 ;
        RECT 2427.740 1783.690 2428.375 1783.860 ;
        RECT 2428.055 1783.660 2428.375 1783.690 ;
        RECT 2428.885 1783.610 2429.060 1787.985 ;
        RECT 2435.975 1785.305 2438.415 1785.445 ;
        RECT 2435.975 1785.155 2436.115 1785.305 ;
        RECT 2435.675 1785.065 2436.115 1785.155 ;
        RECT 2433.335 1784.925 2436.115 1785.065 ;
        RECT 2432.825 1784.785 2433.085 1784.875 ;
        RECT 2433.335 1784.785 2433.475 1784.925 ;
        RECT 2435.675 1784.835 2435.935 1784.925 ;
        RECT 2436.275 1784.835 2436.535 1785.155 ;
        RECT 2436.275 1784.785 2436.475 1784.835 ;
        RECT 2432.825 1784.645 2433.475 1784.785 ;
        RECT 2436.085 1784.645 2436.475 1784.785 ;
        RECT 2437.345 1784.775 2437.625 1785.155 ;
        RECT 2437.835 1784.835 2438.110 1785.155 ;
        RECT 2432.825 1784.555 2433.085 1784.645 ;
        RECT 2425.145 1783.245 2426.025 1783.435 ;
        RECT 2428.830 1783.260 2429.180 1783.610 ;
        RECT 2432.885 1783.475 2433.025 1784.555 ;
        RECT 2433.745 1784.505 2434.025 1784.620 ;
        RECT 2435.195 1784.505 2435.455 1784.595 ;
        RECT 2433.575 1784.365 2435.455 1784.505 ;
        RECT 2433.575 1784.315 2434.025 1784.365 ;
        RECT 2433.515 1784.245 2434.025 1784.315 ;
        RECT 2435.195 1784.275 2435.455 1784.365 ;
        RECT 2433.515 1784.055 2433.775 1784.245 ;
        RECT 2434.690 1784.055 2434.995 1784.060 ;
        RECT 2433.505 1783.685 2433.785 1784.055 ;
        RECT 2433.995 1783.945 2434.255 1784.035 ;
        RECT 2434.585 1783.945 2434.995 1784.055 ;
        RECT 2433.995 1783.805 2434.995 1783.945 ;
        RECT 2433.995 1783.715 2434.255 1783.805 ;
        RECT 2434.585 1783.685 2434.995 1783.805 ;
        RECT 2435.425 1783.685 2435.705 1784.060 ;
        RECT 2436.085 1783.525 2436.225 1784.645 ;
        RECT 2437.415 1784.315 2437.555 1784.775 ;
        RECT 2436.865 1783.685 2437.145 1784.155 ;
        RECT 2437.355 1784.055 2437.615 1784.315 ;
        RECT 2437.345 1783.685 2437.625 1784.055 ;
        RECT 2436.085 1783.475 2436.395 1783.525 ;
        RECT 2437.895 1783.515 2438.035 1784.835 ;
        RECT 2438.275 1784.315 2438.415 1785.305 ;
        RECT 2438.585 1784.555 2438.845 1784.875 ;
        RECT 2440.445 1784.835 2440.705 1785.155 ;
        RECT 2438.215 1783.995 2438.475 1784.315 ;
        RECT 2438.645 1783.515 2438.785 1784.555 ;
        RECT 2440.505 1784.055 2440.645 1784.835 ;
        RECT 2441.710 1784.265 2442.050 1784.345 ;
        RECT 2439.755 1783.945 2440.015 1784.035 ;
        RECT 2439.095 1783.805 2440.015 1783.945 ;
        RECT 2437.555 1783.495 2438.035 1783.515 ;
        RECT 2425.175 1783.235 2426.025 1783.245 ;
        RECT 2425.175 1783.125 2425.455 1783.235 ;
        RECT 2432.825 1783.155 2433.085 1783.475 ;
        RECT 2435.555 1783.385 2435.815 1783.475 ;
        RECT 2436.025 1783.445 2436.395 1783.475 ;
        RECT 2435.555 1783.155 2435.875 1783.385 ;
        RECT 2420.475 1782.865 2423.975 1783.005 ;
        RECT 2435.735 1783.005 2435.875 1783.155 ;
        RECT 2436.025 1783.150 2436.435 1783.445 ;
        RECT 2436.625 1783.155 2436.905 1783.495 ;
        RECT 2437.355 1783.245 2438.035 1783.495 ;
        RECT 2438.575 1783.445 2438.855 1783.515 ;
        RECT 2437.355 1783.145 2437.835 1783.245 ;
        RECT 2438.525 1783.185 2438.900 1783.445 ;
        RECT 2438.575 1783.145 2438.855 1783.185 ;
        RECT 2439.095 1783.005 2439.235 1783.805 ;
        RECT 2439.755 1783.715 2440.015 1783.805 ;
        RECT 2440.335 1783.685 2440.645 1784.055 ;
        RECT 2440.405 1783.500 2440.645 1783.685 ;
        RECT 2441.085 1784.065 2442.050 1784.265 ;
        RECT 2440.405 1783.435 2440.715 1783.500 ;
        RECT 2441.085 1783.435 2441.285 1784.065 ;
        RECT 2441.710 1783.995 2442.050 1784.065 ;
        RECT 2441.800 1783.990 2441.970 1783.995 ;
        RECT 2443.000 1783.860 2443.160 1789.035 ;
        RECT 2444.115 1788.945 2444.440 1789.035 ;
        RECT 2443.315 1788.510 2443.635 1788.835 ;
        RECT 2443.345 1788.335 2443.515 1788.510 ;
        RECT 2443.345 1788.160 2443.520 1788.335 ;
        RECT 2443.345 1787.985 2444.320 1788.160 ;
        RECT 2443.315 1783.860 2443.635 1783.980 ;
        RECT 2443.000 1783.690 2443.635 1783.860 ;
        RECT 2443.315 1783.660 2443.635 1783.690 ;
        RECT 2444.145 1783.610 2444.320 1787.985 ;
        RECT 2440.405 1783.245 2441.285 1783.435 ;
        RECT 2444.090 1783.260 2444.440 1783.610 ;
        RECT 2440.435 1783.235 2441.285 1783.245 ;
        RECT 2440.435 1783.125 2440.715 1783.235 ;
        RECT 2435.735 1782.865 2439.235 1783.005 ;
        RECT 2416.020 1782.145 2416.280 1782.465 ;
        RECT 2431.200 1782.145 2431.460 1782.465 ;
        RECT 2416.080 1773.430 2416.220 1782.145 ;
        RECT 2416.020 1773.110 2416.280 1773.430 ;
        RECT 2400.840 1772.770 2401.100 1773.090 ;
        RECT 2385.660 1772.430 2385.920 1772.750 ;
        RECT 2431.260 1768.330 2431.400 1782.145 ;
        RECT 2431.200 1768.010 2431.460 1768.330 ;
        RECT 2359.575 1710.065 2443.715 1710.235 ;
        RECT 2359.575 1708.880 2359.745 1710.065 ;
        RECT 2443.545 1709.910 2443.715 1710.065 ;
        RECT 2363.685 1709.705 2373.865 1709.875 ;
        RECT 2359.920 1709.515 2360.200 1709.620 ;
        RECT 2359.920 1709.345 2361.110 1709.515 ;
        RECT 2359.920 1709.280 2360.200 1709.345 ;
        RECT 2360.940 1709.140 2361.110 1709.345 ;
        RECT 2363.100 1709.305 2363.470 1709.675 ;
        RECT 2363.685 1709.225 2363.855 1709.705 ;
        RECT 2363.630 1709.140 2363.910 1709.225 ;
        RECT 2360.940 1708.970 2363.910 1709.140 ;
        RECT 2363.630 1708.885 2363.910 1708.970 ;
        RECT 2373.705 1709.200 2373.865 1709.705 ;
        RECT 2380.270 1709.705 2390.450 1709.875 ;
        RECT 2379.685 1709.305 2380.055 1709.675 ;
        RECT 2374.820 1709.200 2375.145 1709.265 ;
        RECT 2373.705 1709.030 2375.145 1709.200 ;
        RECT 2359.535 1708.540 2359.815 1708.880 ;
        RECT 2367.950 1707.415 2368.230 1707.440 ;
        RECT 2367.950 1707.095 2368.240 1707.415 ;
        RECT 2367.950 1707.065 2368.230 1707.095 ;
        RECT 2369.000 1707.065 2369.280 1707.440 ;
        RECT 2370.360 1707.325 2370.620 1707.415 ;
        RECT 2369.740 1707.185 2370.620 1707.325 ;
        RECT 2368.320 1706.045 2368.600 1706.420 ;
        RECT 2367.640 1703.655 2367.920 1704.035 ;
        RECT 2368.380 1704.015 2368.520 1706.045 ;
        RECT 2369.060 1705.285 2369.200 1707.065 ;
        RECT 2369.740 1705.400 2369.880 1707.185 ;
        RECT 2370.360 1707.095 2370.620 1707.185 ;
        RECT 2371.380 1706.075 2371.640 1706.395 ;
        RECT 2369.060 1705.145 2369.540 1705.285 ;
        RECT 2368.980 1704.345 2369.260 1704.720 ;
        RECT 2368.320 1703.695 2368.580 1704.015 ;
        RECT 2369.400 1703.695 2369.540 1705.145 ;
        RECT 2369.680 1705.025 2369.960 1705.400 ;
        RECT 2369.680 1704.005 2369.960 1704.380 ;
        RECT 2371.440 1704.355 2371.580 1706.075 ;
        RECT 2371.380 1704.035 2371.640 1704.355 ;
        RECT 2373.705 1703.860 2373.865 1709.030 ;
        RECT 2374.820 1708.940 2375.145 1709.030 ;
        RECT 2377.210 1709.145 2377.535 1709.270 ;
        RECT 2380.270 1709.225 2380.440 1709.705 ;
        RECT 2377.210 1709.140 2378.260 1709.145 ;
        RECT 2380.215 1709.140 2380.495 1709.225 ;
        RECT 2377.210 1708.975 2380.495 1709.140 ;
        RECT 2377.210 1708.945 2377.535 1708.975 ;
        RECT 2378.260 1708.970 2380.495 1708.975 ;
        RECT 2374.020 1708.565 2374.340 1708.890 ;
        RECT 2380.215 1708.885 2380.495 1708.970 ;
        RECT 2390.290 1709.200 2390.450 1709.705 ;
        RECT 2396.855 1709.710 2407.035 1709.880 ;
        RECT 2396.270 1709.280 2396.640 1709.680 ;
        RECT 2391.405 1709.200 2391.730 1709.265 ;
        RECT 2390.290 1709.030 2391.730 1709.200 ;
        RECT 2374.050 1708.330 2374.220 1708.565 ;
        RECT 2374.050 1708.155 2374.225 1708.330 ;
        RECT 2374.050 1707.980 2375.025 1708.155 ;
        RECT 2374.020 1703.860 2374.340 1703.980 ;
        RECT 2367.685 1703.070 2367.855 1703.655 ;
        RECT 2369.340 1703.355 2369.600 1703.695 ;
        RECT 2373.705 1703.690 2374.340 1703.860 ;
        RECT 2374.020 1703.660 2374.340 1703.690 ;
        RECT 2372.350 1703.290 2372.675 1703.615 ;
        RECT 2374.850 1703.610 2375.025 1707.980 ;
        RECT 2384.535 1707.415 2384.815 1707.440 ;
        RECT 2384.535 1707.095 2384.825 1707.415 ;
        RECT 2384.535 1707.065 2384.815 1707.095 ;
        RECT 2385.585 1707.065 2385.865 1707.440 ;
        RECT 2386.945 1707.325 2387.205 1707.415 ;
        RECT 2386.325 1707.185 2387.205 1707.325 ;
        RECT 2384.905 1706.045 2385.185 1706.420 ;
        RECT 2384.225 1703.655 2384.505 1704.035 ;
        RECT 2384.965 1704.015 2385.105 1706.045 ;
        RECT 2385.645 1705.285 2385.785 1707.065 ;
        RECT 2386.325 1705.400 2386.465 1707.185 ;
        RECT 2386.945 1707.095 2387.205 1707.185 ;
        RECT 2387.965 1706.075 2388.225 1706.395 ;
        RECT 2385.645 1705.145 2386.125 1705.285 ;
        RECT 2385.565 1704.345 2385.845 1704.720 ;
        RECT 2384.905 1703.695 2385.165 1704.015 ;
        RECT 2385.985 1703.695 2386.125 1705.145 ;
        RECT 2386.265 1705.025 2386.545 1705.400 ;
        RECT 2386.265 1704.005 2386.545 1704.380 ;
        RECT 2388.025 1704.355 2388.165 1706.075 ;
        RECT 2387.965 1704.035 2388.225 1704.355 ;
        RECT 2390.290 1703.860 2390.450 1709.030 ;
        RECT 2391.405 1708.940 2391.730 1709.030 ;
        RECT 2393.795 1709.145 2394.120 1709.270 ;
        RECT 2396.855 1709.230 2397.025 1709.710 ;
        RECT 2393.795 1709.140 2395.075 1709.145 ;
        RECT 2396.800 1709.140 2397.080 1709.230 ;
        RECT 2393.795 1708.975 2397.080 1709.140 ;
        RECT 2393.795 1708.945 2394.120 1708.975 ;
        RECT 2395.075 1708.970 2397.080 1708.975 ;
        RECT 2396.800 1708.890 2397.080 1708.970 ;
        RECT 2406.875 1709.205 2407.035 1709.710 ;
        RECT 2413.440 1709.715 2423.620 1709.885 ;
        RECT 2412.855 1709.280 2413.225 1709.685 ;
        RECT 2407.990 1709.205 2408.315 1709.270 ;
        RECT 2406.875 1709.035 2408.315 1709.205 ;
        RECT 2390.605 1708.565 2390.925 1708.890 ;
        RECT 2390.635 1708.330 2390.805 1708.565 ;
        RECT 2390.635 1708.155 2390.810 1708.330 ;
        RECT 2390.635 1707.980 2391.610 1708.155 ;
        RECT 2390.605 1703.860 2390.925 1703.980 ;
        RECT 2372.425 1703.070 2372.595 1703.290 ;
        RECT 2374.795 1703.260 2375.145 1703.610 ;
        RECT 2367.685 1702.900 2372.595 1703.070 ;
        RECT 2384.270 1703.070 2384.440 1703.655 ;
        RECT 2385.925 1703.355 2386.185 1703.695 ;
        RECT 2390.290 1703.690 2390.925 1703.860 ;
        RECT 2390.605 1703.660 2390.925 1703.690 ;
        RECT 2388.935 1703.290 2389.260 1703.615 ;
        RECT 2391.435 1703.610 2391.610 1707.980 ;
        RECT 2401.120 1707.420 2401.400 1707.445 ;
        RECT 2401.120 1707.100 2401.410 1707.420 ;
        RECT 2401.120 1707.070 2401.400 1707.100 ;
        RECT 2402.170 1707.070 2402.450 1707.445 ;
        RECT 2403.530 1707.330 2403.790 1707.420 ;
        RECT 2402.910 1707.190 2403.790 1707.330 ;
        RECT 2401.490 1706.050 2401.770 1706.425 ;
        RECT 2400.810 1703.660 2401.090 1704.040 ;
        RECT 2401.550 1704.020 2401.690 1706.050 ;
        RECT 2402.230 1705.290 2402.370 1707.070 ;
        RECT 2402.910 1705.405 2403.050 1707.190 ;
        RECT 2403.530 1707.100 2403.790 1707.190 ;
        RECT 2404.550 1706.080 2404.810 1706.400 ;
        RECT 2402.230 1705.150 2402.710 1705.290 ;
        RECT 2402.150 1704.350 2402.430 1704.725 ;
        RECT 2401.490 1703.700 2401.750 1704.020 ;
        RECT 2402.570 1703.700 2402.710 1705.150 ;
        RECT 2402.850 1705.030 2403.130 1705.405 ;
        RECT 2402.850 1704.010 2403.130 1704.385 ;
        RECT 2404.610 1704.360 2404.750 1706.080 ;
        RECT 2404.550 1704.040 2404.810 1704.360 ;
        RECT 2406.875 1703.865 2407.035 1709.035 ;
        RECT 2407.990 1708.945 2408.315 1709.035 ;
        RECT 2410.380 1709.150 2410.705 1709.275 ;
        RECT 2413.440 1709.235 2413.610 1709.715 ;
        RECT 2410.380 1709.140 2411.305 1709.150 ;
        RECT 2413.385 1709.140 2413.665 1709.235 ;
        RECT 2410.380 1708.980 2413.665 1709.140 ;
        RECT 2410.380 1708.950 2410.705 1708.980 ;
        RECT 2411.305 1708.970 2413.665 1708.980 ;
        RECT 2413.385 1708.895 2413.665 1708.970 ;
        RECT 2423.460 1709.210 2423.620 1709.715 ;
        RECT 2430.020 1709.715 2440.200 1709.885 ;
        RECT 2429.435 1709.660 2429.805 1709.685 ;
        RECT 2429.435 1709.315 2429.810 1709.660 ;
        RECT 2429.440 1709.280 2429.810 1709.315 ;
        RECT 2424.575 1709.210 2424.900 1709.275 ;
        RECT 2423.460 1709.040 2424.900 1709.210 ;
        RECT 2407.190 1708.570 2407.510 1708.895 ;
        RECT 2407.220 1708.335 2407.390 1708.570 ;
        RECT 2407.220 1708.160 2407.395 1708.335 ;
        RECT 2407.220 1707.985 2408.195 1708.160 ;
        RECT 2407.190 1703.865 2407.510 1703.985 ;
        RECT 2389.010 1703.070 2389.180 1703.290 ;
        RECT 2391.380 1703.260 2391.730 1703.610 ;
        RECT 2384.270 1702.900 2389.180 1703.070 ;
        RECT 2400.855 1703.075 2401.025 1703.660 ;
        RECT 2402.510 1703.360 2402.770 1703.700 ;
        RECT 2406.875 1703.695 2407.510 1703.865 ;
        RECT 2407.190 1703.665 2407.510 1703.695 ;
        RECT 2405.520 1703.295 2405.845 1703.620 ;
        RECT 2408.020 1703.615 2408.195 1707.985 ;
        RECT 2417.705 1707.425 2417.985 1707.450 ;
        RECT 2417.705 1707.105 2417.995 1707.425 ;
        RECT 2417.705 1707.075 2417.985 1707.105 ;
        RECT 2418.755 1707.075 2419.035 1707.450 ;
        RECT 2420.115 1707.335 2420.375 1707.425 ;
        RECT 2419.495 1707.195 2420.375 1707.335 ;
        RECT 2418.075 1706.055 2418.355 1706.430 ;
        RECT 2410.500 1704.090 2410.760 1704.410 ;
        RECT 2405.595 1703.075 2405.765 1703.295 ;
        RECT 2407.965 1703.265 2408.315 1703.615 ;
        RECT 2400.855 1702.905 2405.765 1703.075 ;
        RECT 2377.380 1701.710 2377.640 1702.030 ;
        RECT 2393.940 1701.710 2394.200 1702.030 ;
        RECT 2377.440 1697.270 2377.580 1701.710 ;
        RECT 2394.000 1697.270 2394.140 1701.710 ;
        RECT 2377.380 1696.950 2377.640 1697.270 ;
        RECT 2393.940 1696.950 2394.200 1697.270 ;
        RECT 2410.560 1696.930 2410.700 1704.090 ;
        RECT 2417.395 1703.665 2417.675 1704.045 ;
        RECT 2418.135 1704.025 2418.275 1706.055 ;
        RECT 2418.815 1705.295 2418.955 1707.075 ;
        RECT 2419.495 1705.410 2419.635 1707.195 ;
        RECT 2420.115 1707.105 2420.375 1707.195 ;
        RECT 2421.135 1706.085 2421.395 1706.405 ;
        RECT 2418.815 1705.155 2419.295 1705.295 ;
        RECT 2418.735 1704.355 2419.015 1704.730 ;
        RECT 2418.075 1703.705 2418.335 1704.025 ;
        RECT 2419.155 1703.705 2419.295 1705.155 ;
        RECT 2419.435 1705.035 2419.715 1705.410 ;
        RECT 2419.435 1704.015 2419.715 1704.390 ;
        RECT 2421.195 1704.365 2421.335 1706.085 ;
        RECT 2421.135 1704.045 2421.395 1704.365 ;
        RECT 2423.460 1703.870 2423.620 1709.040 ;
        RECT 2424.575 1708.950 2424.900 1709.040 ;
        RECT 2426.965 1709.155 2427.290 1709.280 ;
        RECT 2430.020 1709.235 2430.190 1709.715 ;
        RECT 2426.965 1709.140 2427.840 1709.155 ;
        RECT 2429.965 1709.140 2430.245 1709.235 ;
        RECT 2426.965 1708.985 2430.245 1709.140 ;
        RECT 2426.965 1708.955 2427.290 1708.985 ;
        RECT 2427.840 1708.970 2430.245 1708.985 ;
        RECT 2423.775 1708.575 2424.095 1708.900 ;
        RECT 2429.965 1708.895 2430.245 1708.970 ;
        RECT 2440.040 1709.210 2440.200 1709.715 ;
        RECT 2443.510 1709.585 2443.835 1709.910 ;
        RECT 2441.155 1709.210 2441.480 1709.275 ;
        RECT 2440.040 1709.040 2441.480 1709.210 ;
        RECT 2423.805 1708.340 2423.975 1708.575 ;
        RECT 2423.805 1708.165 2423.980 1708.340 ;
        RECT 2423.805 1707.990 2424.780 1708.165 ;
        RECT 2423.775 1703.870 2424.095 1703.990 ;
        RECT 2417.440 1703.080 2417.610 1703.665 ;
        RECT 2419.095 1703.365 2419.355 1703.705 ;
        RECT 2423.460 1703.700 2424.095 1703.870 ;
        RECT 2423.775 1703.670 2424.095 1703.700 ;
        RECT 2422.105 1703.300 2422.430 1703.625 ;
        RECT 2424.605 1703.620 2424.780 1707.990 ;
        RECT 2434.285 1707.425 2434.565 1707.450 ;
        RECT 2434.285 1707.105 2434.575 1707.425 ;
        RECT 2434.285 1707.075 2434.565 1707.105 ;
        RECT 2435.335 1707.075 2435.615 1707.450 ;
        RECT 2436.695 1707.335 2436.955 1707.425 ;
        RECT 2436.075 1707.195 2436.955 1707.335 ;
        RECT 2434.655 1706.055 2434.935 1706.430 ;
        RECT 2433.975 1703.665 2434.255 1704.045 ;
        RECT 2434.715 1704.025 2434.855 1706.055 ;
        RECT 2435.395 1705.295 2435.535 1707.075 ;
        RECT 2436.075 1705.410 2436.215 1707.195 ;
        RECT 2436.695 1707.105 2436.955 1707.195 ;
        RECT 2437.715 1706.085 2437.975 1706.405 ;
        RECT 2435.395 1705.155 2435.875 1705.295 ;
        RECT 2435.315 1704.355 2435.595 1704.730 ;
        RECT 2434.655 1703.705 2434.915 1704.025 ;
        RECT 2435.735 1703.705 2435.875 1705.155 ;
        RECT 2436.015 1705.035 2436.295 1705.410 ;
        RECT 2436.015 1704.015 2436.295 1704.390 ;
        RECT 2437.775 1704.365 2437.915 1706.085 ;
        RECT 2437.715 1704.045 2437.975 1704.365 ;
        RECT 2440.040 1703.870 2440.200 1709.040 ;
        RECT 2441.155 1708.950 2441.480 1709.040 ;
        RECT 2440.355 1708.575 2440.675 1708.900 ;
        RECT 2440.385 1708.340 2440.555 1708.575 ;
        RECT 2440.385 1708.165 2440.560 1708.340 ;
        RECT 2440.385 1707.990 2441.360 1708.165 ;
        RECT 2440.355 1703.870 2440.675 1703.990 ;
        RECT 2422.180 1703.080 2422.350 1703.300 ;
        RECT 2424.550 1703.270 2424.900 1703.620 ;
        RECT 2417.440 1702.910 2422.350 1703.080 ;
        RECT 2434.020 1703.080 2434.190 1703.665 ;
        RECT 2435.675 1703.365 2435.935 1703.705 ;
        RECT 2440.040 1703.700 2440.675 1703.870 ;
        RECT 2440.355 1703.670 2440.675 1703.700 ;
        RECT 2438.685 1703.300 2439.010 1703.625 ;
        RECT 2441.185 1703.620 2441.360 1707.990 ;
        RECT 2438.760 1703.080 2438.930 1703.300 ;
        RECT 2441.130 1703.270 2441.480 1703.620 ;
        RECT 2434.020 1702.910 2438.930 1703.080 ;
        RECT 2427.980 1702.160 2428.240 1702.480 ;
        RECT 2410.500 1696.610 2410.760 1696.930 ;
        RECT 2428.040 1676.770 2428.180 1702.160 ;
        RECT 2428.040 1676.630 2428.640 1676.770 ;
        RECT 2428.500 1656.130 2428.640 1676.630 ;
        RECT 2428.440 1655.810 2428.700 1656.130 ;
        RECT 2359.210 1610.055 2446.530 1610.225 ;
        RECT 2359.210 1608.880 2359.380 1610.055 ;
        RECT 2446.360 1609.910 2446.530 1610.055 ;
        RECT 2359.540 1609.515 2359.820 1609.620 ;
        RECT 2359.540 1609.345 2360.745 1609.515 ;
        RECT 2359.540 1609.280 2359.820 1609.345 ;
        RECT 2360.575 1609.140 2360.745 1609.345 ;
        RECT 2362.915 1609.320 2363.285 1609.690 ;
        RECT 2363.440 1609.550 2374.135 1609.720 ;
        RECT 2363.440 1609.170 2363.610 1609.550 ;
        RECT 2373.975 1609.200 2374.135 1609.550 ;
        RECT 2380.135 1609.320 2380.505 1609.690 ;
        RECT 2380.660 1609.550 2391.355 1609.720 ;
        RECT 2375.090 1609.200 2375.415 1609.265 ;
        RECT 2363.390 1609.140 2363.670 1609.170 ;
        RECT 2360.575 1608.970 2363.670 1609.140 ;
        RECT 2359.165 1608.540 2359.445 1608.880 ;
        RECT 2363.390 1608.830 2363.670 1608.970 ;
        RECT 2373.975 1609.030 2375.415 1609.200 ;
        RECT 2367.675 1607.725 2367.955 1608.095 ;
        RECT 2369.045 1608.050 2369.305 1608.095 ;
        RECT 2369.015 1607.805 2369.335 1608.050 ;
        RECT 2369.045 1607.760 2369.305 1607.805 ;
        RECT 2370.745 1607.760 2371.005 1608.095 ;
        RECT 2368.685 1607.065 2368.965 1607.435 ;
        RECT 2369.105 1606.645 2369.245 1607.760 ;
        RECT 2369.725 1607.065 2370.005 1607.435 ;
        RECT 2368.425 1606.505 2369.245 1606.645 ;
        RECT 2365.645 1606.075 2365.905 1606.395 ;
        RECT 2365.705 1604.355 2365.845 1606.075 ;
        RECT 2368.425 1605.800 2368.565 1606.505 ;
        RECT 2370.065 1606.075 2370.325 1606.395 ;
        RECT 2366.315 1605.430 2366.595 1605.800 ;
        RECT 2368.355 1605.430 2368.635 1605.800 ;
        RECT 2365.645 1604.035 2365.905 1604.355 ;
        RECT 2366.385 1604.015 2366.525 1605.430 ;
        RECT 2368.005 1604.690 2368.285 1605.060 ;
        RECT 2368.425 1604.355 2368.565 1605.430 ;
        RECT 2369.375 1605.030 2369.655 1605.400 ;
        RECT 2370.125 1605.375 2370.265 1606.075 ;
        RECT 2370.065 1605.055 2370.325 1605.375 ;
        RECT 2368.365 1604.035 2368.625 1604.355 ;
        RECT 2369.035 1604.350 2369.315 1604.720 ;
        RECT 2370.805 1604.355 2370.945 1607.760 ;
        RECT 2370.745 1604.035 2371.005 1604.355 ;
        RECT 2366.325 1603.695 2366.585 1604.015 ;
        RECT 2367.675 1603.815 2367.955 1603.870 ;
        RECT 2373.975 1603.860 2374.135 1609.030 ;
        RECT 2375.090 1608.940 2375.415 1609.030 ;
        RECT 2377.480 1609.145 2377.805 1609.270 ;
        RECT 2380.660 1609.170 2380.830 1609.550 ;
        RECT 2391.195 1609.200 2391.355 1609.550 ;
        RECT 2397.355 1609.325 2397.725 1609.695 ;
        RECT 2397.880 1609.555 2408.575 1609.725 ;
        RECT 2392.310 1609.200 2392.635 1609.265 ;
        RECT 2377.480 1609.140 2378.715 1609.145 ;
        RECT 2380.610 1609.140 2380.890 1609.170 ;
        RECT 2377.480 1608.975 2380.890 1609.140 ;
        RECT 2377.480 1608.945 2377.805 1608.975 ;
        RECT 2378.715 1608.970 2380.890 1608.975 ;
        RECT 2374.290 1608.565 2374.610 1608.890 ;
        RECT 2380.610 1608.830 2380.890 1608.970 ;
        RECT 2391.195 1609.030 2392.635 1609.200 ;
        RECT 2374.320 1608.330 2374.490 1608.565 ;
        RECT 2374.320 1608.155 2374.495 1608.330 ;
        RECT 2374.320 1607.980 2375.295 1608.155 ;
        RECT 2374.290 1603.860 2374.610 1603.980 ;
        RECT 2367.675 1603.640 2372.325 1603.815 ;
        RECT 2373.975 1603.690 2374.610 1603.860 ;
        RECT 2374.290 1603.660 2374.610 1603.690 ;
        RECT 2367.675 1603.500 2367.955 1603.640 ;
        RECT 2372.150 1603.490 2372.325 1603.640 ;
        RECT 2372.620 1603.490 2372.945 1603.615 ;
        RECT 2375.120 1603.610 2375.295 1607.980 ;
        RECT 2384.895 1607.725 2385.175 1608.095 ;
        RECT 2386.265 1608.050 2386.525 1608.095 ;
        RECT 2386.235 1607.805 2386.555 1608.050 ;
        RECT 2386.265 1607.760 2386.525 1607.805 ;
        RECT 2387.965 1607.760 2388.225 1608.095 ;
        RECT 2385.905 1607.065 2386.185 1607.435 ;
        RECT 2386.325 1606.645 2386.465 1607.760 ;
        RECT 2386.945 1607.065 2387.225 1607.435 ;
        RECT 2385.645 1606.505 2386.465 1606.645 ;
        RECT 2382.865 1606.075 2383.125 1606.395 ;
        RECT 2382.925 1604.355 2383.065 1606.075 ;
        RECT 2385.645 1605.800 2385.785 1606.505 ;
        RECT 2387.285 1606.075 2387.545 1606.395 ;
        RECT 2383.535 1605.430 2383.815 1605.800 ;
        RECT 2385.575 1605.430 2385.855 1605.800 ;
        RECT 2382.865 1604.035 2383.125 1604.355 ;
        RECT 2383.605 1604.015 2383.745 1605.430 ;
        RECT 2385.225 1604.690 2385.505 1605.060 ;
        RECT 2385.645 1604.355 2385.785 1605.430 ;
        RECT 2386.595 1605.030 2386.875 1605.400 ;
        RECT 2387.345 1605.375 2387.485 1606.075 ;
        RECT 2387.285 1605.055 2387.545 1605.375 ;
        RECT 2385.585 1604.035 2385.845 1604.355 ;
        RECT 2386.255 1604.350 2386.535 1604.720 ;
        RECT 2388.025 1604.355 2388.165 1607.760 ;
        RECT 2387.965 1604.035 2388.225 1604.355 ;
        RECT 2383.545 1603.695 2383.805 1604.015 ;
        RECT 2384.895 1603.815 2385.175 1603.870 ;
        RECT 2391.195 1603.860 2391.355 1609.030 ;
        RECT 2392.310 1608.940 2392.635 1609.030 ;
        RECT 2394.700 1609.145 2395.025 1609.270 ;
        RECT 2397.880 1609.175 2398.050 1609.555 ;
        RECT 2408.415 1609.205 2408.575 1609.555 ;
        RECT 2414.575 1609.320 2414.945 1609.690 ;
        RECT 2415.100 1609.550 2425.795 1609.720 ;
        RECT 2409.530 1609.205 2409.855 1609.270 ;
        RECT 2394.700 1609.140 2395.885 1609.145 ;
        RECT 2397.830 1609.140 2398.110 1609.175 ;
        RECT 2394.700 1608.975 2398.120 1609.140 ;
        RECT 2394.700 1608.945 2395.025 1608.975 ;
        RECT 2395.885 1608.970 2398.120 1608.975 ;
        RECT 2408.415 1609.035 2409.855 1609.205 ;
        RECT 2391.510 1608.565 2391.830 1608.890 ;
        RECT 2397.830 1608.835 2398.110 1608.970 ;
        RECT 2391.540 1608.330 2391.710 1608.565 ;
        RECT 2391.540 1608.155 2391.715 1608.330 ;
        RECT 2391.540 1607.980 2392.515 1608.155 ;
        RECT 2391.510 1603.860 2391.830 1603.980 ;
        RECT 2384.895 1603.640 2389.545 1603.815 ;
        RECT 2391.195 1603.690 2391.830 1603.860 ;
        RECT 2391.510 1603.660 2391.830 1603.690 ;
        RECT 2375.065 1603.490 2375.415 1603.610 ;
        RECT 2384.895 1603.500 2385.175 1603.640 ;
        RECT 2372.150 1603.320 2375.415 1603.490 ;
        RECT 2389.370 1603.490 2389.545 1603.640 ;
        RECT 2389.840 1603.490 2390.165 1603.615 ;
        RECT 2392.340 1603.610 2392.515 1607.980 ;
        RECT 2402.115 1607.730 2402.395 1608.100 ;
        RECT 2403.485 1608.055 2403.745 1608.100 ;
        RECT 2403.455 1607.810 2403.775 1608.055 ;
        RECT 2403.485 1607.765 2403.745 1607.810 ;
        RECT 2405.185 1607.765 2405.445 1608.100 ;
        RECT 2403.125 1607.070 2403.405 1607.440 ;
        RECT 2403.545 1606.650 2403.685 1607.765 ;
        RECT 2404.165 1607.070 2404.445 1607.440 ;
        RECT 2402.865 1606.510 2403.685 1606.650 ;
        RECT 2400.085 1606.080 2400.345 1606.400 ;
        RECT 2400.145 1604.360 2400.285 1606.080 ;
        RECT 2402.865 1605.805 2403.005 1606.510 ;
        RECT 2404.505 1606.080 2404.765 1606.400 ;
        RECT 2400.755 1605.435 2401.035 1605.805 ;
        RECT 2402.795 1605.435 2403.075 1605.805 ;
        RECT 2400.085 1604.040 2400.345 1604.360 ;
        RECT 2400.825 1604.020 2400.965 1605.435 ;
        RECT 2402.445 1604.695 2402.725 1605.065 ;
        RECT 2402.865 1604.360 2403.005 1605.435 ;
        RECT 2403.815 1605.035 2404.095 1605.405 ;
        RECT 2404.565 1605.380 2404.705 1606.080 ;
        RECT 2404.505 1605.060 2404.765 1605.380 ;
        RECT 2402.805 1604.040 2403.065 1604.360 ;
        RECT 2403.475 1604.355 2403.755 1604.725 ;
        RECT 2405.245 1604.360 2405.385 1607.765 ;
        RECT 2405.185 1604.040 2405.445 1604.360 ;
        RECT 2400.765 1603.700 2401.025 1604.020 ;
        RECT 2402.115 1603.820 2402.395 1603.875 ;
        RECT 2408.415 1603.865 2408.575 1609.035 ;
        RECT 2409.530 1608.945 2409.855 1609.035 ;
        RECT 2411.920 1609.150 2412.245 1609.275 ;
        RECT 2415.100 1609.170 2415.270 1609.550 ;
        RECT 2425.635 1609.200 2425.795 1609.550 ;
        RECT 2431.795 1609.320 2432.165 1609.690 ;
        RECT 2432.320 1609.550 2443.015 1609.720 ;
        RECT 2446.325 1609.585 2446.650 1609.910 ;
        RECT 2426.750 1609.200 2427.075 1609.265 ;
        RECT 2411.920 1609.145 2412.970 1609.150 ;
        RECT 2411.920 1609.140 2413.045 1609.145 ;
        RECT 2415.050 1609.140 2415.330 1609.170 ;
        RECT 2411.920 1608.980 2415.330 1609.140 ;
        RECT 2411.920 1608.950 2412.245 1608.980 ;
        RECT 2412.970 1608.975 2415.330 1608.980 ;
        RECT 2413.045 1608.970 2415.330 1608.975 ;
        RECT 2408.730 1608.570 2409.050 1608.895 ;
        RECT 2415.050 1608.830 2415.330 1608.970 ;
        RECT 2425.635 1609.030 2427.075 1609.200 ;
        RECT 2408.760 1608.335 2408.930 1608.570 ;
        RECT 2408.760 1608.160 2408.935 1608.335 ;
        RECT 2408.760 1607.985 2409.735 1608.160 ;
        RECT 2408.730 1603.865 2409.050 1603.985 ;
        RECT 2402.115 1603.645 2406.765 1603.820 ;
        RECT 2408.415 1603.695 2409.050 1603.865 ;
        RECT 2408.730 1603.665 2409.050 1603.695 ;
        RECT 2392.285 1603.490 2392.635 1603.610 ;
        RECT 2402.115 1603.505 2402.395 1603.645 ;
        RECT 2389.370 1603.320 2392.635 1603.490 ;
        RECT 2406.590 1603.495 2406.765 1603.645 ;
        RECT 2407.060 1603.495 2407.385 1603.620 ;
        RECT 2409.560 1603.615 2409.735 1607.985 ;
        RECT 2419.335 1607.725 2419.615 1608.095 ;
        RECT 2420.705 1608.050 2420.965 1608.095 ;
        RECT 2420.675 1607.805 2420.995 1608.050 ;
        RECT 2420.705 1607.760 2420.965 1607.805 ;
        RECT 2422.405 1607.760 2422.665 1608.095 ;
        RECT 2420.345 1607.065 2420.625 1607.435 ;
        RECT 2420.765 1606.645 2420.905 1607.760 ;
        RECT 2421.385 1607.065 2421.665 1607.435 ;
        RECT 2420.085 1606.505 2420.905 1606.645 ;
        RECT 2417.305 1606.075 2417.565 1606.395 ;
        RECT 2417.365 1604.355 2417.505 1606.075 ;
        RECT 2420.085 1605.800 2420.225 1606.505 ;
        RECT 2421.725 1606.075 2421.985 1606.395 ;
        RECT 2417.975 1605.430 2418.255 1605.800 ;
        RECT 2420.015 1605.430 2420.295 1605.800 ;
        RECT 2417.305 1604.035 2417.565 1604.355 ;
        RECT 2418.045 1604.015 2418.185 1605.430 ;
        RECT 2419.665 1604.690 2419.945 1605.060 ;
        RECT 2420.085 1604.355 2420.225 1605.430 ;
        RECT 2421.035 1605.030 2421.315 1605.400 ;
        RECT 2421.785 1605.375 2421.925 1606.075 ;
        RECT 2421.725 1605.055 2421.985 1605.375 ;
        RECT 2420.025 1604.035 2420.285 1604.355 ;
        RECT 2420.695 1604.350 2420.975 1604.720 ;
        RECT 2422.465 1604.355 2422.605 1607.760 ;
        RECT 2422.405 1604.035 2422.665 1604.355 ;
        RECT 2417.985 1603.695 2418.245 1604.015 ;
        RECT 2419.335 1603.815 2419.615 1603.870 ;
        RECT 2425.635 1603.860 2425.795 1609.030 ;
        RECT 2426.750 1608.940 2427.075 1609.030 ;
        RECT 2429.140 1609.145 2429.465 1609.270 ;
        RECT 2432.320 1609.170 2432.490 1609.550 ;
        RECT 2442.855 1609.200 2443.015 1609.550 ;
        RECT 2443.970 1609.200 2444.295 1609.265 ;
        RECT 2429.140 1609.140 2429.925 1609.145 ;
        RECT 2432.270 1609.140 2432.550 1609.170 ;
        RECT 2429.140 1608.975 2432.550 1609.140 ;
        RECT 2429.140 1608.945 2429.465 1608.975 ;
        RECT 2429.925 1608.970 2432.550 1608.975 ;
        RECT 2425.950 1608.565 2426.270 1608.890 ;
        RECT 2432.270 1608.830 2432.550 1608.970 ;
        RECT 2442.855 1609.030 2444.295 1609.200 ;
        RECT 2425.980 1608.330 2426.150 1608.565 ;
        RECT 2425.980 1608.155 2426.155 1608.330 ;
        RECT 2425.980 1607.980 2426.955 1608.155 ;
        RECT 2425.950 1603.860 2426.270 1603.980 ;
        RECT 2419.335 1603.640 2423.985 1603.815 ;
        RECT 2425.635 1603.690 2426.270 1603.860 ;
        RECT 2425.950 1603.660 2426.270 1603.690 ;
        RECT 2409.505 1603.495 2409.855 1603.615 ;
        RECT 2419.335 1603.500 2419.615 1603.640 ;
        RECT 2406.590 1603.325 2409.855 1603.495 ;
        RECT 2372.620 1603.290 2372.945 1603.320 ;
        RECT 2375.065 1603.260 2375.415 1603.320 ;
        RECT 2389.840 1603.290 2390.165 1603.320 ;
        RECT 2392.285 1603.260 2392.635 1603.320 ;
        RECT 2407.060 1603.295 2407.385 1603.325 ;
        RECT 2409.505 1603.265 2409.855 1603.325 ;
        RECT 2423.810 1603.490 2423.985 1603.640 ;
        RECT 2424.280 1603.490 2424.605 1603.615 ;
        RECT 2426.780 1603.610 2426.955 1607.980 ;
        RECT 2436.555 1607.725 2436.835 1608.095 ;
        RECT 2437.925 1608.050 2438.185 1608.095 ;
        RECT 2437.895 1607.805 2438.215 1608.050 ;
        RECT 2437.925 1607.760 2438.185 1607.805 ;
        RECT 2439.625 1607.760 2439.885 1608.095 ;
        RECT 2437.565 1607.065 2437.845 1607.435 ;
        RECT 2437.985 1606.645 2438.125 1607.760 ;
        RECT 2438.605 1607.065 2438.885 1607.435 ;
        RECT 2437.305 1606.505 2438.125 1606.645 ;
        RECT 2434.525 1606.075 2434.785 1606.395 ;
        RECT 2434.585 1604.355 2434.725 1606.075 ;
        RECT 2437.305 1605.800 2437.445 1606.505 ;
        RECT 2438.945 1606.075 2439.205 1606.395 ;
        RECT 2435.195 1605.430 2435.475 1605.800 ;
        RECT 2437.235 1605.430 2437.515 1605.800 ;
        RECT 2434.525 1604.035 2434.785 1604.355 ;
        RECT 2435.265 1604.015 2435.405 1605.430 ;
        RECT 2436.885 1604.690 2437.165 1605.060 ;
        RECT 2437.305 1604.355 2437.445 1605.430 ;
        RECT 2438.255 1605.030 2438.535 1605.400 ;
        RECT 2439.005 1605.375 2439.145 1606.075 ;
        RECT 2438.945 1605.055 2439.205 1605.375 ;
        RECT 2437.245 1604.035 2437.505 1604.355 ;
        RECT 2437.915 1604.350 2438.195 1604.720 ;
        RECT 2439.685 1604.355 2439.825 1607.760 ;
        RECT 2439.625 1604.035 2439.885 1604.355 ;
        RECT 2435.205 1603.695 2435.465 1604.015 ;
        RECT 2436.555 1603.815 2436.835 1603.870 ;
        RECT 2442.855 1603.860 2443.015 1609.030 ;
        RECT 2443.970 1608.940 2444.295 1609.030 ;
        RECT 2443.170 1608.565 2443.490 1608.890 ;
        RECT 2443.200 1608.330 2443.370 1608.565 ;
        RECT 2443.200 1608.155 2443.375 1608.330 ;
        RECT 2443.200 1607.980 2444.175 1608.155 ;
        RECT 2443.170 1603.860 2443.490 1603.980 ;
        RECT 2436.555 1603.640 2441.205 1603.815 ;
        RECT 2442.855 1603.690 2443.490 1603.860 ;
        RECT 2443.170 1603.660 2443.490 1603.690 ;
        RECT 2426.725 1603.490 2427.075 1603.610 ;
        RECT 2436.555 1603.500 2436.835 1603.640 ;
        RECT 2423.810 1603.320 2427.075 1603.490 ;
        RECT 2441.030 1603.490 2441.205 1603.640 ;
        RECT 2441.500 1603.490 2441.825 1603.615 ;
        RECT 2444.000 1603.610 2444.175 1607.980 ;
        RECT 2443.945 1603.490 2444.295 1603.610 ;
        RECT 2441.030 1603.320 2444.295 1603.490 ;
        RECT 2424.280 1603.290 2424.605 1603.320 ;
        RECT 2426.725 1603.260 2427.075 1603.320 ;
        RECT 2441.500 1603.290 2441.825 1603.320 ;
        RECT 2443.945 1603.260 2444.295 1603.320 ;
        RECT 2377.380 1602.145 2377.640 1602.465 ;
        RECT 2377.440 1593.910 2377.580 1602.145 ;
        RECT 2411.880 1602.090 2412.140 1602.410 ;
        RECT 2395.320 1601.750 2395.580 1602.070 ;
        RECT 2395.380 1593.910 2395.520 1601.750 ;
        RECT 2377.380 1593.590 2377.640 1593.910 ;
        RECT 2395.320 1593.590 2395.580 1593.910 ;
        RECT 2411.940 1593.570 2412.080 1602.090 ;
        RECT 2429.820 1601.750 2430.080 1602.070 ;
        RECT 2411.880 1593.250 2412.140 1593.570 ;
        RECT 2429.880 1593.230 2430.020 1601.750 ;
        RECT 2429.820 1592.910 2430.080 1593.230 ;
        RECT 2359.225 1533.685 2442.050 1533.855 ;
        RECT 2359.225 1531.890 2359.395 1533.685 ;
        RECT 2441.880 1532.910 2442.050 1533.685 ;
        RECT 2359.540 1532.510 2359.830 1532.635 ;
        RECT 2359.540 1532.505 2359.860 1532.510 ;
        RECT 2359.540 1532.335 2360.880 1532.505 ;
        RECT 2368.100 1532.340 2368.470 1532.710 ;
        RECT 2384.425 1532.340 2384.795 1532.710 ;
        RECT 2400.750 1532.340 2401.120 1532.710 ;
        RECT 2417.075 1532.340 2417.445 1532.710 ;
        RECT 2433.400 1532.340 2433.770 1532.710 ;
        RECT 2441.850 1532.560 2442.200 1532.910 ;
        RECT 2359.540 1532.285 2359.830 1532.335 ;
        RECT 2360.710 1532.140 2360.880 1532.335 ;
        RECT 2369.585 1532.140 2369.935 1532.240 ;
        RECT 2374.190 1532.200 2374.515 1532.265 ;
        RECT 2360.710 1531.970 2369.935 1532.140 ;
        RECT 2369.585 1531.890 2369.935 1531.970 ;
        RECT 2373.075 1532.030 2374.515 1532.200 ;
        RECT 2359.165 1531.540 2359.455 1531.890 ;
        RECT 2362.595 1528.185 2366.255 1528.325 ;
        RECT 2361.805 1527.135 2362.085 1527.510 ;
        RECT 2362.595 1527.505 2362.735 1528.185 ;
        RECT 2363.015 1527.955 2363.275 1528.045 ;
        RECT 2363.015 1527.815 2364.695 1527.955 ;
        RECT 2363.015 1527.725 2363.275 1527.815 ;
        RECT 2364.555 1527.765 2364.695 1527.815 ;
        RECT 2364.555 1527.535 2364.995 1527.765 ;
        RECT 2362.595 1527.255 2363.045 1527.505 ;
        RECT 2364.735 1527.445 2364.995 1527.535 ;
        RECT 2365.515 1527.445 2365.835 1527.765 ;
        RECT 2366.115 1527.505 2366.255 1528.185 ;
        RECT 2366.425 1527.955 2366.705 1528.070 ;
        RECT 2367.505 1527.955 2369.685 1528.065 ;
        RECT 2366.425 1527.905 2369.685 1527.955 ;
        RECT 2366.425 1527.815 2367.645 1527.905 ;
        RECT 2366.425 1527.695 2366.705 1527.815 ;
        RECT 2368.345 1527.505 2368.645 1527.510 ;
        RECT 2362.765 1527.135 2363.045 1527.255 ;
        RECT 2361.865 1525.515 2362.035 1527.135 ;
        RECT 2364.055 1526.950 2364.455 1527.115 ;
        RECT 2364.055 1526.925 2364.525 1526.950 ;
        RECT 2362.775 1526.835 2363.035 1526.925 ;
        RECT 2362.775 1526.695 2363.815 1526.835 ;
        RECT 2362.775 1526.605 2363.035 1526.695 ;
        RECT 2363.245 1526.015 2363.525 1526.390 ;
        RECT 2363.675 1526.045 2363.815 1526.695 ;
        RECT 2363.995 1526.605 2364.525 1526.925 ;
        RECT 2364.245 1526.575 2364.525 1526.605 ;
        RECT 2364.965 1526.575 2365.245 1526.950 ;
        RECT 2365.515 1526.645 2365.655 1527.445 ;
        RECT 2366.115 1527.395 2368.645 1527.505 ;
        RECT 2369.135 1527.445 2369.395 1527.765 ;
        RECT 2369.135 1527.395 2369.335 1527.445 ;
        RECT 2366.115 1527.365 2369.335 1527.395 ;
        RECT 2368.365 1527.255 2369.335 1527.365 ;
        RECT 2365.815 1527.115 2366.075 1527.205 ;
        RECT 2368.365 1527.135 2368.645 1527.255 ;
        RECT 2365.815 1526.950 2366.135 1527.115 ;
        RECT 2365.815 1526.885 2366.205 1526.950 ;
        RECT 2365.455 1526.325 2365.715 1526.645 ;
        RECT 2365.925 1526.575 2366.205 1526.885 ;
        RECT 2366.805 1526.575 2367.085 1526.950 ;
        RECT 2367.415 1526.605 2367.675 1526.925 ;
        RECT 2366.435 1526.045 2366.695 1526.365 ;
        RECT 2363.675 1525.905 2366.635 1526.045 ;
        RECT 2367.475 1525.905 2367.615 1526.605 ;
        RECT 2368.485 1526.575 2368.765 1526.945 ;
        RECT 2368.555 1525.905 2368.695 1526.575 ;
        RECT 2368.935 1526.365 2369.075 1527.255 ;
        RECT 2369.535 1526.925 2369.685 1527.905 ;
        RECT 2369.255 1526.785 2369.685 1526.925 ;
        RECT 2373.075 1526.860 2373.235 1532.030 ;
        RECT 2374.190 1531.940 2374.515 1532.030 ;
        RECT 2376.570 1532.170 2376.920 1532.290 ;
        RECT 2385.075 1532.170 2385.425 1532.245 ;
        RECT 2390.515 1532.200 2390.840 1532.265 ;
        RECT 2376.570 1531.970 2385.425 1532.170 ;
        RECT 2376.570 1531.940 2376.920 1531.970 ;
        RECT 2385.075 1531.895 2385.425 1531.970 ;
        RECT 2389.400 1532.030 2390.840 1532.200 ;
        RECT 2373.390 1531.505 2373.710 1531.830 ;
        RECT 2373.420 1531.330 2373.590 1531.505 ;
        RECT 2373.420 1531.155 2373.595 1531.330 ;
        RECT 2373.420 1530.980 2374.395 1531.155 ;
        RECT 2373.390 1526.860 2373.710 1526.980 ;
        RECT 2369.255 1526.605 2369.515 1526.785 ;
        RECT 2369.965 1526.555 2370.245 1526.785 ;
        RECT 2373.075 1526.690 2373.710 1526.860 ;
        RECT 2373.390 1526.660 2373.710 1526.690 ;
        RECT 2370.575 1526.555 2370.835 1526.645 ;
        RECT 2374.220 1526.610 2374.395 1530.980 ;
        RECT 2378.920 1528.185 2382.580 1528.325 ;
        RECT 2378.130 1527.135 2378.410 1527.510 ;
        RECT 2378.920 1527.505 2379.060 1528.185 ;
        RECT 2379.340 1527.955 2379.600 1528.045 ;
        RECT 2379.340 1527.815 2381.020 1527.955 ;
        RECT 2379.340 1527.725 2379.600 1527.815 ;
        RECT 2380.880 1527.765 2381.020 1527.815 ;
        RECT 2380.880 1527.535 2381.320 1527.765 ;
        RECT 2378.920 1527.255 2379.370 1527.505 ;
        RECT 2381.060 1527.445 2381.320 1527.535 ;
        RECT 2381.840 1527.445 2382.160 1527.765 ;
        RECT 2382.440 1527.505 2382.580 1528.185 ;
        RECT 2382.750 1527.955 2383.030 1528.070 ;
        RECT 2383.830 1527.955 2386.010 1528.065 ;
        RECT 2382.750 1527.905 2386.010 1527.955 ;
        RECT 2382.750 1527.815 2383.970 1527.905 ;
        RECT 2382.750 1527.695 2383.030 1527.815 ;
        RECT 2384.670 1527.505 2384.970 1527.510 ;
        RECT 2379.090 1527.135 2379.370 1527.255 ;
        RECT 2369.675 1526.415 2370.835 1526.555 ;
        RECT 2368.875 1526.045 2369.135 1526.365 ;
        RECT 2369.675 1525.905 2369.815 1526.415 ;
        RECT 2370.575 1526.325 2370.835 1526.415 ;
        RECT 2374.165 1526.260 2374.515 1526.610 ;
        RECT 2371.860 1526.105 2372.030 1526.110 ;
        RECT 2367.475 1525.765 2369.815 1525.905 ;
        RECT 2371.770 1525.755 2372.110 1526.105 ;
        RECT 2371.770 1525.515 2372.030 1525.755 ;
        RECT 2361.865 1525.355 2372.030 1525.515 ;
        RECT 2378.190 1525.515 2378.360 1527.135 ;
        RECT 2380.380 1526.950 2380.780 1527.115 ;
        RECT 2380.380 1526.925 2380.850 1526.950 ;
        RECT 2379.100 1526.835 2379.360 1526.925 ;
        RECT 2379.100 1526.695 2380.140 1526.835 ;
        RECT 2379.100 1526.605 2379.360 1526.695 ;
        RECT 2379.570 1526.015 2379.850 1526.390 ;
        RECT 2380.000 1526.045 2380.140 1526.695 ;
        RECT 2380.320 1526.605 2380.850 1526.925 ;
        RECT 2380.570 1526.575 2380.850 1526.605 ;
        RECT 2381.290 1526.575 2381.570 1526.950 ;
        RECT 2381.840 1526.645 2381.980 1527.445 ;
        RECT 2382.440 1527.395 2384.970 1527.505 ;
        RECT 2385.460 1527.445 2385.720 1527.765 ;
        RECT 2385.460 1527.395 2385.660 1527.445 ;
        RECT 2382.440 1527.365 2385.660 1527.395 ;
        RECT 2384.690 1527.255 2385.660 1527.365 ;
        RECT 2382.140 1527.115 2382.400 1527.205 ;
        RECT 2384.690 1527.135 2384.970 1527.255 ;
        RECT 2382.140 1526.950 2382.460 1527.115 ;
        RECT 2382.140 1526.885 2382.530 1526.950 ;
        RECT 2381.780 1526.325 2382.040 1526.645 ;
        RECT 2382.250 1526.575 2382.530 1526.885 ;
        RECT 2383.130 1526.575 2383.410 1526.950 ;
        RECT 2383.740 1526.605 2384.000 1526.925 ;
        RECT 2382.760 1526.045 2383.020 1526.365 ;
        RECT 2380.000 1525.905 2382.960 1526.045 ;
        RECT 2383.800 1525.905 2383.940 1526.605 ;
        RECT 2384.810 1526.575 2385.090 1526.945 ;
        RECT 2384.880 1525.905 2385.020 1526.575 ;
        RECT 2385.260 1526.365 2385.400 1527.255 ;
        RECT 2385.860 1526.925 2386.010 1527.905 ;
        RECT 2385.580 1526.785 2386.010 1526.925 ;
        RECT 2389.400 1526.860 2389.560 1532.030 ;
        RECT 2390.515 1531.940 2390.840 1532.030 ;
        RECT 2392.895 1532.175 2393.245 1532.295 ;
        RECT 2401.400 1532.175 2401.750 1532.250 ;
        RECT 2406.840 1532.200 2407.165 1532.265 ;
        RECT 2392.895 1531.975 2401.750 1532.175 ;
        RECT 2392.895 1531.945 2393.245 1531.975 ;
        RECT 2401.400 1531.900 2401.750 1531.975 ;
        RECT 2405.725 1532.030 2407.165 1532.200 ;
        RECT 2389.715 1531.505 2390.035 1531.830 ;
        RECT 2389.745 1531.330 2389.915 1531.505 ;
        RECT 2389.745 1531.155 2389.920 1531.330 ;
        RECT 2389.745 1530.980 2390.720 1531.155 ;
        RECT 2389.715 1526.860 2390.035 1526.980 ;
        RECT 2385.580 1526.605 2385.840 1526.785 ;
        RECT 2386.290 1526.555 2386.570 1526.785 ;
        RECT 2389.400 1526.690 2390.035 1526.860 ;
        RECT 2389.715 1526.660 2390.035 1526.690 ;
        RECT 2386.900 1526.555 2387.160 1526.645 ;
        RECT 2390.545 1526.610 2390.720 1530.980 ;
        RECT 2395.245 1528.185 2398.905 1528.325 ;
        RECT 2393.020 1526.950 2393.280 1527.270 ;
        RECT 2394.455 1527.135 2394.735 1527.510 ;
        RECT 2395.245 1527.505 2395.385 1528.185 ;
        RECT 2395.665 1527.955 2395.925 1528.045 ;
        RECT 2395.665 1527.815 2397.345 1527.955 ;
        RECT 2395.665 1527.725 2395.925 1527.815 ;
        RECT 2397.205 1527.765 2397.345 1527.815 ;
        RECT 2397.205 1527.535 2397.645 1527.765 ;
        RECT 2395.245 1527.255 2395.695 1527.505 ;
        RECT 2397.385 1527.445 2397.645 1527.535 ;
        RECT 2398.165 1527.445 2398.485 1527.765 ;
        RECT 2398.765 1527.505 2398.905 1528.185 ;
        RECT 2399.075 1527.955 2399.355 1528.070 ;
        RECT 2400.155 1527.955 2402.335 1528.065 ;
        RECT 2399.075 1527.905 2402.335 1527.955 ;
        RECT 2399.075 1527.815 2400.295 1527.905 ;
        RECT 2399.075 1527.695 2399.355 1527.815 ;
        RECT 2400.995 1527.505 2401.295 1527.510 ;
        RECT 2395.415 1527.135 2395.695 1527.255 ;
        RECT 2386.000 1526.415 2387.160 1526.555 ;
        RECT 2385.200 1526.045 2385.460 1526.365 ;
        RECT 2386.000 1525.905 2386.140 1526.415 ;
        RECT 2386.900 1526.325 2387.160 1526.415 ;
        RECT 2390.490 1526.260 2390.840 1526.610 ;
        RECT 2388.185 1526.105 2388.355 1526.110 ;
        RECT 2383.800 1525.765 2386.140 1525.905 ;
        RECT 2388.095 1525.755 2388.435 1526.105 ;
        RECT 2388.095 1525.515 2388.355 1525.755 ;
        RECT 2371.805 1525.350 2372.030 1525.355 ;
        RECT 2376.460 1525.150 2376.720 1525.470 ;
        RECT 2378.190 1525.355 2388.355 1525.515 ;
        RECT 2388.130 1525.350 2388.355 1525.355 ;
        RECT 2376.520 1518.090 2376.660 1525.150 ;
        RECT 2393.080 1518.090 2393.220 1526.950 ;
        RECT 2394.515 1525.515 2394.685 1527.135 ;
        RECT 2396.705 1526.950 2397.105 1527.115 ;
        RECT 2396.705 1526.925 2397.175 1526.950 ;
        RECT 2395.425 1526.835 2395.685 1526.925 ;
        RECT 2395.425 1526.695 2396.465 1526.835 ;
        RECT 2395.425 1526.605 2395.685 1526.695 ;
        RECT 2395.895 1526.015 2396.175 1526.390 ;
        RECT 2396.325 1526.045 2396.465 1526.695 ;
        RECT 2396.645 1526.605 2397.175 1526.925 ;
        RECT 2396.895 1526.575 2397.175 1526.605 ;
        RECT 2397.615 1526.575 2397.895 1526.950 ;
        RECT 2398.165 1526.645 2398.305 1527.445 ;
        RECT 2398.765 1527.395 2401.295 1527.505 ;
        RECT 2401.785 1527.445 2402.045 1527.765 ;
        RECT 2401.785 1527.395 2401.985 1527.445 ;
        RECT 2398.765 1527.365 2401.985 1527.395 ;
        RECT 2401.015 1527.255 2401.985 1527.365 ;
        RECT 2398.465 1527.115 2398.725 1527.205 ;
        RECT 2401.015 1527.135 2401.295 1527.255 ;
        RECT 2398.465 1526.950 2398.785 1527.115 ;
        RECT 2398.465 1526.885 2398.855 1526.950 ;
        RECT 2398.105 1526.325 2398.365 1526.645 ;
        RECT 2398.575 1526.575 2398.855 1526.885 ;
        RECT 2399.455 1526.575 2399.735 1526.950 ;
        RECT 2400.065 1526.605 2400.325 1526.925 ;
        RECT 2399.085 1526.045 2399.345 1526.365 ;
        RECT 2396.325 1525.905 2399.285 1526.045 ;
        RECT 2400.125 1525.905 2400.265 1526.605 ;
        RECT 2401.135 1526.575 2401.415 1526.945 ;
        RECT 2401.205 1525.905 2401.345 1526.575 ;
        RECT 2401.585 1526.365 2401.725 1527.255 ;
        RECT 2402.185 1526.925 2402.335 1527.905 ;
        RECT 2401.905 1526.785 2402.335 1526.925 ;
        RECT 2405.725 1526.860 2405.885 1532.030 ;
        RECT 2406.840 1531.940 2407.165 1532.030 ;
        RECT 2409.175 1532.170 2409.525 1532.290 ;
        RECT 2417.725 1532.170 2418.075 1532.245 ;
        RECT 2423.165 1532.200 2423.490 1532.265 ;
        RECT 2409.175 1531.970 2418.075 1532.170 ;
        RECT 2409.175 1531.940 2409.525 1531.970 ;
        RECT 2417.725 1531.895 2418.075 1531.970 ;
        RECT 2422.050 1532.030 2423.490 1532.200 ;
        RECT 2406.040 1531.505 2406.360 1531.830 ;
        RECT 2406.070 1531.330 2406.240 1531.505 ;
        RECT 2406.070 1531.155 2406.245 1531.330 ;
        RECT 2406.070 1530.980 2407.045 1531.155 ;
        RECT 2406.040 1526.860 2406.360 1526.980 ;
        RECT 2401.905 1526.605 2402.165 1526.785 ;
        RECT 2402.615 1526.555 2402.895 1526.785 ;
        RECT 2405.725 1526.690 2406.360 1526.860 ;
        RECT 2406.040 1526.660 2406.360 1526.690 ;
        RECT 2403.225 1526.555 2403.485 1526.645 ;
        RECT 2406.870 1526.610 2407.045 1530.980 ;
        RECT 2411.570 1528.185 2415.230 1528.325 ;
        RECT 2410.780 1527.135 2411.060 1527.510 ;
        RECT 2411.570 1527.505 2411.710 1528.185 ;
        RECT 2411.990 1527.955 2412.250 1528.045 ;
        RECT 2411.990 1527.815 2413.670 1527.955 ;
        RECT 2411.990 1527.725 2412.250 1527.815 ;
        RECT 2413.530 1527.765 2413.670 1527.815 ;
        RECT 2413.530 1527.535 2413.970 1527.765 ;
        RECT 2411.570 1527.255 2412.020 1527.505 ;
        RECT 2413.710 1527.445 2413.970 1527.535 ;
        RECT 2414.490 1527.445 2414.810 1527.765 ;
        RECT 2415.090 1527.505 2415.230 1528.185 ;
        RECT 2415.400 1527.955 2415.680 1528.070 ;
        RECT 2416.480 1527.955 2418.660 1528.065 ;
        RECT 2415.400 1527.905 2418.660 1527.955 ;
        RECT 2415.400 1527.815 2416.620 1527.905 ;
        RECT 2415.400 1527.695 2415.680 1527.815 ;
        RECT 2417.320 1527.505 2417.620 1527.510 ;
        RECT 2411.740 1527.135 2412.020 1527.255 ;
        RECT 2402.325 1526.415 2403.485 1526.555 ;
        RECT 2401.525 1526.045 2401.785 1526.365 ;
        RECT 2402.325 1525.905 2402.465 1526.415 ;
        RECT 2403.225 1526.325 2403.485 1526.415 ;
        RECT 2406.815 1526.260 2407.165 1526.610 ;
        RECT 2404.510 1526.105 2404.680 1526.110 ;
        RECT 2400.125 1525.765 2402.465 1525.905 ;
        RECT 2404.420 1525.755 2404.760 1526.105 ;
        RECT 2404.420 1525.515 2404.680 1525.755 ;
        RECT 2394.515 1525.355 2404.680 1525.515 ;
        RECT 2410.840 1525.515 2411.010 1527.135 ;
        RECT 2413.030 1526.950 2413.430 1527.115 ;
        RECT 2413.030 1526.925 2413.500 1526.950 ;
        RECT 2411.750 1526.835 2412.010 1526.925 ;
        RECT 2411.750 1526.695 2412.790 1526.835 ;
        RECT 2411.750 1526.605 2412.010 1526.695 ;
        RECT 2412.220 1526.015 2412.500 1526.390 ;
        RECT 2412.650 1526.045 2412.790 1526.695 ;
        RECT 2412.970 1526.605 2413.500 1526.925 ;
        RECT 2413.220 1526.575 2413.500 1526.605 ;
        RECT 2413.940 1526.575 2414.220 1526.950 ;
        RECT 2414.490 1526.645 2414.630 1527.445 ;
        RECT 2415.090 1527.395 2417.620 1527.505 ;
        RECT 2418.110 1527.445 2418.370 1527.765 ;
        RECT 2418.110 1527.395 2418.310 1527.445 ;
        RECT 2415.090 1527.365 2418.310 1527.395 ;
        RECT 2417.340 1527.255 2418.310 1527.365 ;
        RECT 2414.790 1527.115 2415.050 1527.205 ;
        RECT 2417.340 1527.135 2417.620 1527.255 ;
        RECT 2414.790 1526.950 2415.110 1527.115 ;
        RECT 2414.790 1526.885 2415.180 1526.950 ;
        RECT 2414.430 1526.325 2414.690 1526.645 ;
        RECT 2414.900 1526.575 2415.180 1526.885 ;
        RECT 2415.780 1526.575 2416.060 1526.950 ;
        RECT 2416.390 1526.605 2416.650 1526.925 ;
        RECT 2415.410 1526.045 2415.670 1526.365 ;
        RECT 2412.650 1525.905 2415.610 1526.045 ;
        RECT 2416.450 1525.905 2416.590 1526.605 ;
        RECT 2417.460 1526.575 2417.740 1526.945 ;
        RECT 2417.530 1525.905 2417.670 1526.575 ;
        RECT 2417.910 1526.365 2418.050 1527.255 ;
        RECT 2418.510 1526.925 2418.660 1527.905 ;
        RECT 2418.230 1526.785 2418.660 1526.925 ;
        RECT 2422.050 1526.860 2422.210 1532.030 ;
        RECT 2423.165 1531.940 2423.490 1532.030 ;
        RECT 2425.500 1532.170 2425.850 1532.290 ;
        RECT 2434.055 1532.170 2434.405 1532.245 ;
        RECT 2439.490 1532.200 2439.815 1532.265 ;
        RECT 2425.500 1531.970 2434.405 1532.170 ;
        RECT 2425.500 1531.940 2425.850 1531.970 ;
        RECT 2434.055 1531.895 2434.405 1531.970 ;
        RECT 2438.375 1532.030 2439.815 1532.200 ;
        RECT 2422.365 1531.505 2422.685 1531.830 ;
        RECT 2422.395 1531.330 2422.565 1531.505 ;
        RECT 2422.395 1531.155 2422.570 1531.330 ;
        RECT 2422.395 1530.980 2423.370 1531.155 ;
        RECT 2422.365 1526.860 2422.685 1526.980 ;
        RECT 2418.230 1526.605 2418.490 1526.785 ;
        RECT 2418.940 1526.555 2419.220 1526.785 ;
        RECT 2422.050 1526.690 2422.685 1526.860 ;
        RECT 2422.365 1526.660 2422.685 1526.690 ;
        RECT 2419.550 1526.555 2419.810 1526.645 ;
        RECT 2423.195 1526.610 2423.370 1530.980 ;
        RECT 2427.895 1528.185 2431.555 1528.325 ;
        RECT 2425.680 1526.950 2425.940 1527.270 ;
        RECT 2427.105 1527.135 2427.385 1527.510 ;
        RECT 2427.895 1527.505 2428.035 1528.185 ;
        RECT 2428.315 1527.955 2428.575 1528.045 ;
        RECT 2428.315 1527.815 2429.995 1527.955 ;
        RECT 2428.315 1527.725 2428.575 1527.815 ;
        RECT 2429.855 1527.765 2429.995 1527.815 ;
        RECT 2429.855 1527.535 2430.295 1527.765 ;
        RECT 2427.895 1527.255 2428.345 1527.505 ;
        RECT 2430.035 1527.445 2430.295 1527.535 ;
        RECT 2430.815 1527.445 2431.135 1527.765 ;
        RECT 2431.415 1527.505 2431.555 1528.185 ;
        RECT 2431.725 1527.955 2432.005 1528.070 ;
        RECT 2432.805 1527.955 2434.985 1528.065 ;
        RECT 2431.725 1527.905 2434.985 1527.955 ;
        RECT 2431.725 1527.815 2432.945 1527.905 ;
        RECT 2431.725 1527.695 2432.005 1527.815 ;
        RECT 2433.645 1527.505 2433.945 1527.510 ;
        RECT 2428.065 1527.135 2428.345 1527.255 ;
        RECT 2418.650 1526.415 2419.810 1526.555 ;
        RECT 2417.850 1526.045 2418.110 1526.365 ;
        RECT 2418.650 1525.905 2418.790 1526.415 ;
        RECT 2419.550 1526.325 2419.810 1526.415 ;
        RECT 2423.140 1526.260 2423.490 1526.610 ;
        RECT 2420.835 1526.105 2421.005 1526.110 ;
        RECT 2416.450 1525.765 2418.790 1525.905 ;
        RECT 2420.745 1525.755 2421.085 1526.105 ;
        RECT 2420.745 1525.515 2421.005 1525.755 ;
        RECT 2404.455 1525.350 2404.680 1525.355 ;
        RECT 2409.120 1525.150 2409.380 1525.470 ;
        RECT 2410.840 1525.355 2421.005 1525.515 ;
        RECT 2420.780 1525.350 2421.005 1525.355 ;
        RECT 2409.180 1518.090 2409.320 1525.150 ;
        RECT 2425.740 1518.090 2425.880 1526.950 ;
        RECT 2427.165 1525.515 2427.335 1527.135 ;
        RECT 2429.355 1526.950 2429.755 1527.115 ;
        RECT 2429.355 1526.925 2429.825 1526.950 ;
        RECT 2428.075 1526.835 2428.335 1526.925 ;
        RECT 2428.075 1526.695 2429.115 1526.835 ;
        RECT 2428.075 1526.605 2428.335 1526.695 ;
        RECT 2428.545 1526.015 2428.825 1526.390 ;
        RECT 2428.975 1526.045 2429.115 1526.695 ;
        RECT 2429.295 1526.605 2429.825 1526.925 ;
        RECT 2429.545 1526.575 2429.825 1526.605 ;
        RECT 2430.265 1526.575 2430.545 1526.950 ;
        RECT 2430.815 1526.645 2430.955 1527.445 ;
        RECT 2431.415 1527.395 2433.945 1527.505 ;
        RECT 2434.435 1527.445 2434.695 1527.765 ;
        RECT 2434.435 1527.395 2434.635 1527.445 ;
        RECT 2431.415 1527.365 2434.635 1527.395 ;
        RECT 2433.665 1527.255 2434.635 1527.365 ;
        RECT 2431.115 1527.115 2431.375 1527.205 ;
        RECT 2433.665 1527.135 2433.945 1527.255 ;
        RECT 2431.115 1526.950 2431.435 1527.115 ;
        RECT 2431.115 1526.885 2431.505 1526.950 ;
        RECT 2430.755 1526.325 2431.015 1526.645 ;
        RECT 2431.225 1526.575 2431.505 1526.885 ;
        RECT 2432.105 1526.575 2432.385 1526.950 ;
        RECT 2432.715 1526.605 2432.975 1526.925 ;
        RECT 2431.735 1526.045 2431.995 1526.365 ;
        RECT 2428.975 1525.905 2431.935 1526.045 ;
        RECT 2432.775 1525.905 2432.915 1526.605 ;
        RECT 2433.785 1526.575 2434.065 1526.945 ;
        RECT 2433.855 1525.905 2433.995 1526.575 ;
        RECT 2434.235 1526.365 2434.375 1527.255 ;
        RECT 2434.835 1526.925 2434.985 1527.905 ;
        RECT 2434.555 1526.785 2434.985 1526.925 ;
        RECT 2438.375 1526.860 2438.535 1532.030 ;
        RECT 2439.490 1531.940 2439.815 1532.030 ;
        RECT 2438.690 1531.505 2439.010 1531.830 ;
        RECT 2438.720 1531.330 2438.890 1531.505 ;
        RECT 2438.720 1531.155 2438.895 1531.330 ;
        RECT 2438.720 1530.980 2439.695 1531.155 ;
        RECT 2438.690 1526.860 2439.010 1526.980 ;
        RECT 2434.555 1526.605 2434.815 1526.785 ;
        RECT 2435.265 1526.555 2435.545 1526.785 ;
        RECT 2438.375 1526.690 2439.010 1526.860 ;
        RECT 2438.690 1526.660 2439.010 1526.690 ;
        RECT 2435.875 1526.555 2436.135 1526.645 ;
        RECT 2439.520 1526.610 2439.695 1530.980 ;
        RECT 2434.975 1526.415 2436.135 1526.555 ;
        RECT 2434.175 1526.045 2434.435 1526.365 ;
        RECT 2434.975 1525.905 2435.115 1526.415 ;
        RECT 2435.875 1526.325 2436.135 1526.415 ;
        RECT 2439.465 1526.260 2439.815 1526.610 ;
        RECT 2437.160 1526.105 2437.330 1526.110 ;
        RECT 2432.775 1525.765 2435.115 1525.905 ;
        RECT 2437.070 1525.755 2437.410 1526.105 ;
        RECT 2437.070 1525.515 2437.330 1525.755 ;
        RECT 2427.165 1525.355 2437.330 1525.515 ;
        RECT 2437.105 1525.350 2437.330 1525.355 ;
        RECT 2452.820 1524.910 2453.080 1525.230 ;
        RECT 2376.460 1517.770 2376.720 1518.090 ;
        RECT 2393.020 1517.770 2393.280 1518.090 ;
        RECT 2409.120 1517.770 2409.380 1518.090 ;
        RECT 2425.680 1517.770 2425.940 1518.090 ;
        RECT 2452.880 1462.670 2453.020 1524.910 ;
        RECT 2453.800 1490.550 2453.940 2049.870 ;
        RECT 2459.780 1504.150 2459.920 2246.730 ;
        RECT 2577.020 2229.390 2577.280 2229.710 ;
        RECT 2466.620 2207.970 2466.880 2208.290 ;
        RECT 2460.180 2154.930 2460.440 2155.250 ;
        RECT 2459.720 1503.830 2459.980 1504.150 ;
        RECT 2460.240 1497.350 2460.380 2154.930 ;
        RECT 2466.680 2042.370 2466.820 2207.970 ;
        RECT 2473.520 2201.170 2473.780 2201.490 ;
        RECT 2466.620 2042.050 2466.880 2042.370 ;
        RECT 2466.620 1947.190 2466.880 1947.510 ;
        RECT 2460.640 1781.950 2460.900 1782.270 ;
        RECT 2460.180 1497.030 2460.440 1497.350 ;
        RECT 2453.740 1490.230 2454.000 1490.550 ;
        RECT 2460.700 1483.410 2460.840 1781.950 ;
        RECT 2461.100 1701.710 2461.360 1702.030 ;
        RECT 2460.640 1483.090 2460.900 1483.410 ;
        RECT 2461.160 1476.610 2461.300 1701.710 ;
        RECT 2461.560 1601.750 2461.820 1602.070 ;
        RECT 2461.100 1476.290 2461.360 1476.610 ;
        RECT 2461.620 1469.810 2461.760 1601.750 ;
        RECT 2466.680 1483.070 2466.820 1947.190 ;
        RECT 2473.580 1938.670 2473.720 2201.170 ;
        RECT 2480.420 2194.370 2480.680 2194.690 ;
        RECT 2473.520 1938.350 2473.780 1938.670 ;
        RECT 2480.480 1772.750 2480.620 2194.370 ;
        RECT 2487.320 2187.230 2487.580 2187.550 ;
        RECT 2480.420 1772.430 2480.680 1772.750 ;
        RECT 2487.380 1696.590 2487.520 2187.230 ;
        RECT 2494.220 2180.430 2494.480 2180.750 ;
        RECT 2487.320 1696.270 2487.580 1696.590 ;
        RECT 2494.280 1592.890 2494.420 2180.430 ;
        RECT 2501.120 2173.630 2501.380 2173.950 ;
        RECT 2494.220 1592.570 2494.480 1592.890 ;
        RECT 2501.180 1517.070 2501.320 2173.630 ;
        RECT 2508.020 2166.490 2508.280 2166.810 ;
        RECT 2501.120 1516.750 2501.380 1517.070 ;
        RECT 2466.620 1482.750 2466.880 1483.070 ;
        RECT 2461.560 1469.490 2461.820 1469.810 ;
        RECT 2452.820 1462.350 2453.080 1462.670 ;
        RECT 2464.780 1449.090 2465.040 1449.410 ;
        RECT 2459.720 1441.950 2459.980 1442.270 ;
        RECT 2359.225 1435.690 2453.225 1435.860 ;
        RECT 2359.225 1433.895 2359.395 1435.690 ;
        RECT 2453.055 1434.915 2453.225 1435.690 ;
        RECT 2359.540 1434.520 2359.830 1434.640 ;
        RECT 2359.540 1434.515 2359.860 1434.520 ;
        RECT 2359.540 1434.345 2360.730 1434.515 ;
        RECT 2370.315 1434.345 2370.690 1434.715 ;
        RECT 2388.875 1434.345 2389.250 1434.715 ;
        RECT 2407.435 1434.345 2407.810 1434.715 ;
        RECT 2425.995 1434.345 2426.370 1434.715 ;
        RECT 2444.555 1434.345 2444.930 1434.715 ;
        RECT 2453.025 1434.565 2453.375 1434.915 ;
        RECT 2359.540 1434.290 2359.830 1434.345 ;
        RECT 2360.560 1434.145 2360.730 1434.345 ;
        RECT 2370.990 1434.145 2371.340 1434.245 ;
        RECT 2376.425 1434.205 2376.750 1434.270 ;
        RECT 2360.560 1433.975 2371.340 1434.145 ;
        RECT 2370.990 1433.895 2371.340 1433.975 ;
        RECT 2375.310 1434.035 2376.750 1434.205 ;
        RECT 2359.165 1433.545 2359.455 1433.895 ;
        RECT 2368.190 1430.430 2374.280 1430.620 ;
        RECT 2368.190 1430.180 2368.360 1430.430 ;
        RECT 2361.810 1429.805 2362.090 1430.180 ;
        RECT 2366.580 1429.835 2366.840 1430.155 ;
        RECT 2361.820 1429.555 2362.080 1429.805 ;
        RECT 2364.250 1429.595 2364.530 1429.620 ;
        RECT 2362.780 1429.275 2363.040 1429.595 ;
        RECT 2363.900 1429.505 2364.530 1429.595 ;
        RECT 2366.220 1429.505 2366.480 1429.595 ;
        RECT 2363.900 1429.365 2366.480 1429.505 ;
        RECT 2363.900 1429.275 2364.530 1429.365 ;
        RECT 2366.220 1429.275 2366.480 1429.365 ;
        RECT 2362.290 1428.685 2362.570 1429.060 ;
        RECT 2362.840 1428.475 2362.980 1429.275 ;
        RECT 2364.250 1429.245 2364.530 1429.275 ;
        RECT 2365.690 1429.035 2365.970 1429.060 ;
        RECT 2365.690 1428.715 2366.220 1429.035 ;
        RECT 2365.690 1428.685 2365.970 1428.715 ;
        RECT 2362.780 1428.155 2363.040 1428.475 ;
        RECT 2364.740 1428.385 2365.000 1428.475 ;
        RECT 2366.220 1428.385 2366.480 1428.475 ;
        RECT 2366.640 1428.385 2366.780 1429.835 ;
        RECT 2368.130 1429.805 2368.410 1430.180 ;
        RECT 2369.140 1429.835 2369.400 1430.155 ;
        RECT 2369.620 1429.835 2369.880 1430.155 ;
        RECT 2366.930 1429.245 2367.210 1429.620 ;
        RECT 2368.200 1429.615 2368.340 1429.805 ;
        RECT 2368.010 1429.505 2368.340 1429.615 ;
        RECT 2367.720 1429.365 2368.340 1429.505 ;
        RECT 2367.000 1428.475 2367.140 1429.245 ;
        RECT 2367.720 1428.475 2367.860 1429.365 ;
        RECT 2368.010 1429.245 2368.290 1429.365 ;
        RECT 2368.660 1428.945 2368.920 1429.035 ;
        RECT 2368.080 1428.805 2368.920 1428.945 ;
        RECT 2364.740 1428.245 2365.780 1428.385 ;
        RECT 2364.740 1428.155 2365.000 1428.245 ;
        RECT 2365.640 1428.005 2365.780 1428.245 ;
        RECT 2366.220 1428.245 2366.780 1428.385 ;
        RECT 2366.220 1428.155 2366.480 1428.245 ;
        RECT 2366.940 1428.155 2367.200 1428.475 ;
        RECT 2367.660 1428.155 2367.920 1428.475 ;
        RECT 2368.080 1428.005 2368.220 1428.805 ;
        RECT 2368.660 1428.715 2368.920 1428.805 ;
        RECT 2369.200 1428.475 2369.340 1429.835 ;
        RECT 2369.620 1429.785 2369.820 1429.835 ;
        RECT 2370.090 1429.805 2370.370 1430.180 ;
        RECT 2371.090 1429.805 2371.370 1430.180 ;
        RECT 2374.090 1429.795 2374.280 1430.430 ;
        RECT 2369.560 1429.615 2369.820 1429.785 ;
        RECT 2369.560 1429.245 2370.060 1429.615 ;
        RECT 2370.620 1429.275 2370.880 1429.595 ;
        RECT 2374.020 1429.445 2374.360 1429.795 ;
        RECT 2374.110 1429.440 2374.280 1429.445 ;
        RECT 2369.560 1428.475 2369.700 1429.245 ;
        RECT 2370.680 1428.475 2370.820 1429.275 ;
        RECT 2375.310 1428.860 2375.470 1434.035 ;
        RECT 2376.425 1433.945 2376.750 1434.035 ;
        RECT 2378.805 1434.175 2379.155 1434.295 ;
        RECT 2389.550 1434.175 2389.900 1434.250 ;
        RECT 2394.985 1434.205 2395.310 1434.270 ;
        RECT 2378.805 1433.975 2389.900 1434.175 ;
        RECT 2378.805 1433.945 2379.155 1433.975 ;
        RECT 2389.550 1433.900 2389.900 1433.975 ;
        RECT 2393.870 1434.035 2395.310 1434.205 ;
        RECT 2375.625 1433.510 2375.945 1433.835 ;
        RECT 2375.655 1433.335 2375.825 1433.510 ;
        RECT 2375.655 1433.160 2375.830 1433.335 ;
        RECT 2375.655 1432.985 2376.630 1433.160 ;
        RECT 2375.625 1428.860 2375.945 1428.980 ;
        RECT 2375.310 1428.690 2375.945 1428.860 ;
        RECT 2375.625 1428.660 2375.945 1428.690 ;
        RECT 2376.455 1428.610 2376.630 1432.985 ;
        RECT 2386.750 1430.430 2392.840 1430.620 ;
        RECT 2386.750 1430.180 2386.920 1430.430 ;
        RECT 2380.370 1429.805 2380.650 1430.180 ;
        RECT 2385.140 1429.835 2385.400 1430.155 ;
        RECT 2380.380 1429.555 2380.640 1429.805 ;
        RECT 2382.810 1429.595 2383.090 1429.620 ;
        RECT 2381.340 1429.275 2381.600 1429.595 ;
        RECT 2382.460 1429.505 2383.090 1429.595 ;
        RECT 2384.780 1429.505 2385.040 1429.595 ;
        RECT 2382.460 1429.365 2385.040 1429.505 ;
        RECT 2382.460 1429.275 2383.090 1429.365 ;
        RECT 2384.780 1429.275 2385.040 1429.365 ;
        RECT 2380.850 1428.685 2381.130 1429.060 ;
        RECT 2368.900 1428.245 2369.340 1428.475 ;
        RECT 2368.900 1428.155 2369.160 1428.245 ;
        RECT 2369.500 1428.155 2369.760 1428.475 ;
        RECT 2370.620 1428.155 2370.880 1428.475 ;
        RECT 2372.050 1428.125 2372.330 1428.500 ;
        RECT 2376.400 1428.260 2376.750 1428.610 ;
        RECT 2381.400 1428.475 2381.540 1429.275 ;
        RECT 2382.810 1429.245 2383.090 1429.275 ;
        RECT 2384.250 1429.035 2384.530 1429.060 ;
        RECT 2384.250 1428.715 2384.780 1429.035 ;
        RECT 2384.250 1428.685 2384.530 1428.715 ;
        RECT 2381.340 1428.155 2381.600 1428.475 ;
        RECT 2383.300 1428.385 2383.560 1428.475 ;
        RECT 2384.780 1428.385 2385.040 1428.475 ;
        RECT 2385.200 1428.385 2385.340 1429.835 ;
        RECT 2386.690 1429.805 2386.970 1430.180 ;
        RECT 2387.700 1429.835 2387.960 1430.155 ;
        RECT 2388.180 1429.835 2388.440 1430.155 ;
        RECT 2385.490 1429.245 2385.770 1429.620 ;
        RECT 2386.760 1429.615 2386.900 1429.805 ;
        RECT 2386.570 1429.505 2386.900 1429.615 ;
        RECT 2386.280 1429.365 2386.900 1429.505 ;
        RECT 2385.560 1428.475 2385.700 1429.245 ;
        RECT 2386.280 1428.475 2386.420 1429.365 ;
        RECT 2386.570 1429.245 2386.850 1429.365 ;
        RECT 2387.220 1428.945 2387.480 1429.035 ;
        RECT 2386.640 1428.805 2387.480 1428.945 ;
        RECT 2383.300 1428.245 2384.340 1428.385 ;
        RECT 2383.300 1428.155 2383.560 1428.245 ;
        RECT 2365.640 1427.865 2368.220 1428.005 ;
        RECT 2384.200 1428.005 2384.340 1428.245 ;
        RECT 2384.780 1428.245 2385.340 1428.385 ;
        RECT 2384.780 1428.155 2385.040 1428.245 ;
        RECT 2385.500 1428.155 2385.760 1428.475 ;
        RECT 2386.220 1428.155 2386.480 1428.475 ;
        RECT 2386.640 1428.005 2386.780 1428.805 ;
        RECT 2387.220 1428.715 2387.480 1428.805 ;
        RECT 2387.760 1428.475 2387.900 1429.835 ;
        RECT 2388.180 1429.785 2388.380 1429.835 ;
        RECT 2388.650 1429.805 2388.930 1430.180 ;
        RECT 2389.650 1429.805 2389.930 1430.180 ;
        RECT 2392.650 1429.795 2392.840 1430.430 ;
        RECT 2388.120 1429.615 2388.380 1429.785 ;
        RECT 2388.120 1429.245 2388.620 1429.615 ;
        RECT 2389.180 1429.275 2389.440 1429.595 ;
        RECT 2392.580 1429.445 2392.920 1429.795 ;
        RECT 2392.670 1429.440 2392.840 1429.445 ;
        RECT 2388.120 1428.475 2388.260 1429.245 ;
        RECT 2389.240 1428.475 2389.380 1429.275 ;
        RECT 2393.870 1428.860 2394.030 1434.035 ;
        RECT 2394.985 1433.945 2395.310 1434.035 ;
        RECT 2397.365 1434.180 2397.715 1434.300 ;
        RECT 2408.105 1434.180 2408.455 1434.255 ;
        RECT 2413.545 1434.205 2413.870 1434.270 ;
        RECT 2397.365 1433.980 2408.455 1434.180 ;
        RECT 2397.365 1433.950 2397.715 1433.980 ;
        RECT 2408.105 1433.905 2408.455 1433.980 ;
        RECT 2412.430 1434.035 2413.870 1434.205 ;
        RECT 2394.185 1433.510 2394.505 1433.835 ;
        RECT 2394.215 1433.335 2394.385 1433.510 ;
        RECT 2394.215 1433.160 2394.390 1433.335 ;
        RECT 2394.215 1432.985 2395.190 1433.160 ;
        RECT 2394.185 1428.860 2394.505 1428.980 ;
        RECT 2393.870 1428.690 2394.505 1428.860 ;
        RECT 2394.185 1428.660 2394.505 1428.690 ;
        RECT 2395.015 1428.610 2395.190 1432.985 ;
        RECT 2405.310 1430.430 2411.400 1430.620 ;
        RECT 2405.310 1430.180 2405.480 1430.430 ;
        RECT 2398.930 1429.805 2399.210 1430.180 ;
        RECT 2403.700 1429.835 2403.960 1430.155 ;
        RECT 2398.940 1429.555 2399.200 1429.805 ;
        RECT 2401.370 1429.595 2401.650 1429.620 ;
        RECT 2397.160 1429.030 2397.420 1429.350 ;
        RECT 2399.900 1429.275 2400.160 1429.595 ;
        RECT 2401.020 1429.505 2401.650 1429.595 ;
        RECT 2403.340 1429.505 2403.600 1429.595 ;
        RECT 2401.020 1429.365 2403.600 1429.505 ;
        RECT 2401.020 1429.275 2401.650 1429.365 ;
        RECT 2403.340 1429.275 2403.600 1429.365 ;
        RECT 2387.460 1428.245 2387.900 1428.475 ;
        RECT 2387.460 1428.155 2387.720 1428.245 ;
        RECT 2388.060 1428.155 2388.320 1428.475 ;
        RECT 2389.180 1428.155 2389.440 1428.475 ;
        RECT 2390.610 1428.125 2390.890 1428.500 ;
        RECT 2394.960 1428.260 2395.310 1428.610 ;
        RECT 2384.200 1427.865 2386.780 1428.005 ;
        RECT 2378.760 1427.150 2379.020 1427.470 ;
        RECT 2378.820 1421.530 2378.960 1427.150 ;
        RECT 2397.220 1421.530 2397.360 1429.030 ;
        RECT 2399.410 1428.685 2399.690 1429.060 ;
        RECT 2399.960 1428.475 2400.100 1429.275 ;
        RECT 2401.370 1429.245 2401.650 1429.275 ;
        RECT 2402.810 1429.035 2403.090 1429.060 ;
        RECT 2402.810 1428.715 2403.340 1429.035 ;
        RECT 2402.810 1428.685 2403.090 1428.715 ;
        RECT 2399.900 1428.155 2400.160 1428.475 ;
        RECT 2401.860 1428.385 2402.120 1428.475 ;
        RECT 2403.340 1428.385 2403.600 1428.475 ;
        RECT 2403.760 1428.385 2403.900 1429.835 ;
        RECT 2405.250 1429.805 2405.530 1430.180 ;
        RECT 2406.260 1429.835 2406.520 1430.155 ;
        RECT 2406.740 1429.835 2407.000 1430.155 ;
        RECT 2404.050 1429.245 2404.330 1429.620 ;
        RECT 2405.320 1429.615 2405.460 1429.805 ;
        RECT 2405.130 1429.505 2405.460 1429.615 ;
        RECT 2404.840 1429.365 2405.460 1429.505 ;
        RECT 2404.120 1428.475 2404.260 1429.245 ;
        RECT 2404.840 1428.475 2404.980 1429.365 ;
        RECT 2405.130 1429.245 2405.410 1429.365 ;
        RECT 2405.780 1428.945 2406.040 1429.035 ;
        RECT 2405.200 1428.805 2406.040 1428.945 ;
        RECT 2401.860 1428.245 2402.900 1428.385 ;
        RECT 2401.860 1428.155 2402.120 1428.245 ;
        RECT 2402.760 1428.005 2402.900 1428.245 ;
        RECT 2403.340 1428.245 2403.900 1428.385 ;
        RECT 2403.340 1428.155 2403.600 1428.245 ;
        RECT 2404.060 1428.155 2404.320 1428.475 ;
        RECT 2404.780 1428.155 2405.040 1428.475 ;
        RECT 2405.200 1428.005 2405.340 1428.805 ;
        RECT 2405.780 1428.715 2406.040 1428.805 ;
        RECT 2406.320 1428.475 2406.460 1429.835 ;
        RECT 2406.740 1429.785 2406.940 1429.835 ;
        RECT 2407.210 1429.805 2407.490 1430.180 ;
        RECT 2408.210 1429.805 2408.490 1430.180 ;
        RECT 2411.210 1429.795 2411.400 1430.430 ;
        RECT 2406.680 1429.615 2406.940 1429.785 ;
        RECT 2406.680 1429.245 2407.180 1429.615 ;
        RECT 2407.740 1429.275 2408.000 1429.595 ;
        RECT 2411.140 1429.445 2411.480 1429.795 ;
        RECT 2411.230 1429.440 2411.400 1429.445 ;
        RECT 2406.680 1428.475 2406.820 1429.245 ;
        RECT 2407.800 1428.475 2407.940 1429.275 ;
        RECT 2412.430 1428.860 2412.590 1434.035 ;
        RECT 2413.545 1433.945 2413.870 1434.035 ;
        RECT 2415.880 1434.175 2416.230 1434.295 ;
        RECT 2426.665 1434.175 2427.015 1434.250 ;
        RECT 2432.105 1434.205 2432.430 1434.270 ;
        RECT 2415.880 1433.975 2427.015 1434.175 ;
        RECT 2415.880 1433.945 2416.230 1433.975 ;
        RECT 2426.665 1433.900 2427.015 1433.975 ;
        RECT 2430.990 1434.035 2432.430 1434.205 ;
        RECT 2412.745 1433.510 2413.065 1433.835 ;
        RECT 2412.775 1433.335 2412.945 1433.510 ;
        RECT 2412.775 1433.160 2412.950 1433.335 ;
        RECT 2412.775 1432.985 2413.750 1433.160 ;
        RECT 2412.745 1428.860 2413.065 1428.980 ;
        RECT 2412.430 1428.690 2413.065 1428.860 ;
        RECT 2412.745 1428.660 2413.065 1428.690 ;
        RECT 2413.575 1428.610 2413.750 1432.985 ;
        RECT 2423.870 1430.430 2429.960 1430.620 ;
        RECT 2423.870 1430.180 2424.040 1430.430 ;
        RECT 2417.490 1429.805 2417.770 1430.180 ;
        RECT 2422.260 1429.835 2422.520 1430.155 ;
        RECT 2417.500 1429.555 2417.760 1429.805 ;
        RECT 2419.930 1429.595 2420.210 1429.620 ;
        RECT 2418.460 1429.275 2418.720 1429.595 ;
        RECT 2419.580 1429.505 2420.210 1429.595 ;
        RECT 2421.900 1429.505 2422.160 1429.595 ;
        RECT 2419.580 1429.365 2422.160 1429.505 ;
        RECT 2419.580 1429.275 2420.210 1429.365 ;
        RECT 2421.900 1429.275 2422.160 1429.365 ;
        RECT 2417.970 1428.685 2418.250 1429.060 ;
        RECT 2406.020 1428.245 2406.460 1428.475 ;
        RECT 2406.020 1428.155 2406.280 1428.245 ;
        RECT 2406.620 1428.155 2406.880 1428.475 ;
        RECT 2407.740 1428.155 2408.000 1428.475 ;
        RECT 2409.170 1428.125 2409.450 1428.500 ;
        RECT 2413.520 1428.260 2413.870 1428.610 ;
        RECT 2418.520 1428.475 2418.660 1429.275 ;
        RECT 2419.930 1429.245 2420.210 1429.275 ;
        RECT 2421.370 1429.035 2421.650 1429.060 ;
        RECT 2421.370 1428.715 2421.900 1429.035 ;
        RECT 2421.370 1428.685 2421.650 1428.715 ;
        RECT 2418.460 1428.155 2418.720 1428.475 ;
        RECT 2420.420 1428.385 2420.680 1428.475 ;
        RECT 2421.900 1428.385 2422.160 1428.475 ;
        RECT 2422.320 1428.385 2422.460 1429.835 ;
        RECT 2423.810 1429.805 2424.090 1430.180 ;
        RECT 2424.820 1429.835 2425.080 1430.155 ;
        RECT 2425.300 1429.835 2425.560 1430.155 ;
        RECT 2422.610 1429.245 2422.890 1429.620 ;
        RECT 2423.880 1429.615 2424.020 1429.805 ;
        RECT 2423.690 1429.505 2424.020 1429.615 ;
        RECT 2423.400 1429.365 2424.020 1429.505 ;
        RECT 2422.680 1428.475 2422.820 1429.245 ;
        RECT 2423.400 1428.475 2423.540 1429.365 ;
        RECT 2423.690 1429.245 2423.970 1429.365 ;
        RECT 2424.340 1428.945 2424.600 1429.035 ;
        RECT 2423.760 1428.805 2424.600 1428.945 ;
        RECT 2420.420 1428.245 2421.460 1428.385 ;
        RECT 2420.420 1428.155 2420.680 1428.245 ;
        RECT 2402.760 1427.865 2405.340 1428.005 ;
        RECT 2421.320 1428.005 2421.460 1428.245 ;
        RECT 2421.900 1428.245 2422.460 1428.385 ;
        RECT 2421.900 1428.155 2422.160 1428.245 ;
        RECT 2422.620 1428.155 2422.880 1428.475 ;
        RECT 2423.340 1428.155 2423.600 1428.475 ;
        RECT 2423.760 1428.005 2423.900 1428.805 ;
        RECT 2424.340 1428.715 2424.600 1428.805 ;
        RECT 2424.880 1428.475 2425.020 1429.835 ;
        RECT 2425.300 1429.785 2425.500 1429.835 ;
        RECT 2425.770 1429.805 2426.050 1430.180 ;
        RECT 2426.770 1429.805 2427.050 1430.180 ;
        RECT 2429.770 1429.795 2429.960 1430.430 ;
        RECT 2425.240 1429.615 2425.500 1429.785 ;
        RECT 2425.240 1429.245 2425.740 1429.615 ;
        RECT 2426.300 1429.275 2426.560 1429.595 ;
        RECT 2429.700 1429.445 2430.040 1429.795 ;
        RECT 2429.790 1429.440 2429.960 1429.445 ;
        RECT 2425.240 1428.475 2425.380 1429.245 ;
        RECT 2426.360 1428.475 2426.500 1429.275 ;
        RECT 2430.990 1428.860 2431.150 1434.035 ;
        RECT 2432.105 1433.945 2432.430 1434.035 ;
        RECT 2434.440 1434.175 2434.790 1434.295 ;
        RECT 2445.225 1434.175 2445.575 1434.250 ;
        RECT 2450.665 1434.205 2450.990 1434.270 ;
        RECT 2434.440 1433.975 2445.575 1434.175 ;
        RECT 2434.440 1433.945 2434.790 1433.975 ;
        RECT 2445.225 1433.900 2445.575 1433.975 ;
        RECT 2449.550 1434.035 2450.990 1434.205 ;
        RECT 2431.305 1433.510 2431.625 1433.835 ;
        RECT 2431.335 1433.335 2431.505 1433.510 ;
        RECT 2431.335 1433.160 2431.510 1433.335 ;
        RECT 2431.335 1432.985 2432.310 1433.160 ;
        RECT 2431.305 1428.860 2431.625 1428.980 ;
        RECT 2430.990 1428.690 2431.625 1428.860 ;
        RECT 2431.305 1428.660 2431.625 1428.690 ;
        RECT 2432.135 1428.610 2432.310 1432.985 ;
        RECT 2442.430 1430.430 2448.520 1430.620 ;
        RECT 2442.430 1430.180 2442.600 1430.430 ;
        RECT 2436.050 1429.805 2436.330 1430.180 ;
        RECT 2440.820 1429.835 2441.080 1430.155 ;
        RECT 2436.060 1429.555 2436.320 1429.805 ;
        RECT 2438.490 1429.595 2438.770 1429.620 ;
        RECT 2437.020 1429.275 2437.280 1429.595 ;
        RECT 2438.140 1429.505 2438.770 1429.595 ;
        RECT 2440.460 1429.505 2440.720 1429.595 ;
        RECT 2438.140 1429.365 2440.720 1429.505 ;
        RECT 2438.140 1429.275 2438.770 1429.365 ;
        RECT 2440.460 1429.275 2440.720 1429.365 ;
        RECT 2436.530 1428.685 2436.810 1429.060 ;
        RECT 2424.580 1428.245 2425.020 1428.475 ;
        RECT 2424.580 1428.155 2424.840 1428.245 ;
        RECT 2425.180 1428.155 2425.440 1428.475 ;
        RECT 2426.300 1428.155 2426.560 1428.475 ;
        RECT 2427.730 1428.125 2428.010 1428.500 ;
        RECT 2432.080 1428.260 2432.430 1428.610 ;
        RECT 2437.080 1428.475 2437.220 1429.275 ;
        RECT 2438.490 1429.245 2438.770 1429.275 ;
        RECT 2439.930 1429.035 2440.210 1429.060 ;
        RECT 2439.930 1428.715 2440.460 1429.035 ;
        RECT 2439.930 1428.685 2440.210 1428.715 ;
        RECT 2437.020 1428.155 2437.280 1428.475 ;
        RECT 2438.980 1428.385 2439.240 1428.475 ;
        RECT 2440.460 1428.385 2440.720 1428.475 ;
        RECT 2440.880 1428.385 2441.020 1429.835 ;
        RECT 2442.370 1429.805 2442.650 1430.180 ;
        RECT 2443.380 1429.835 2443.640 1430.155 ;
        RECT 2443.860 1429.835 2444.120 1430.155 ;
        RECT 2441.170 1429.245 2441.450 1429.620 ;
        RECT 2442.440 1429.615 2442.580 1429.805 ;
        RECT 2442.250 1429.505 2442.580 1429.615 ;
        RECT 2441.960 1429.365 2442.580 1429.505 ;
        RECT 2441.240 1428.475 2441.380 1429.245 ;
        RECT 2441.960 1428.475 2442.100 1429.365 ;
        RECT 2442.250 1429.245 2442.530 1429.365 ;
        RECT 2442.900 1428.945 2443.160 1429.035 ;
        RECT 2442.320 1428.805 2443.160 1428.945 ;
        RECT 2438.980 1428.245 2440.020 1428.385 ;
        RECT 2438.980 1428.155 2439.240 1428.245 ;
        RECT 2421.320 1427.865 2423.900 1428.005 ;
        RECT 2439.880 1428.005 2440.020 1428.245 ;
        RECT 2440.460 1428.245 2441.020 1428.385 ;
        RECT 2440.460 1428.155 2440.720 1428.245 ;
        RECT 2441.180 1428.155 2441.440 1428.475 ;
        RECT 2441.900 1428.155 2442.160 1428.475 ;
        RECT 2442.320 1428.005 2442.460 1428.805 ;
        RECT 2442.900 1428.715 2443.160 1428.805 ;
        RECT 2443.440 1428.475 2443.580 1429.835 ;
        RECT 2443.860 1429.785 2444.060 1429.835 ;
        RECT 2444.330 1429.805 2444.610 1430.180 ;
        RECT 2445.330 1429.805 2445.610 1430.180 ;
        RECT 2448.330 1429.795 2448.520 1430.430 ;
        RECT 2443.800 1429.615 2444.060 1429.785 ;
        RECT 2443.800 1429.245 2444.300 1429.615 ;
        RECT 2444.860 1429.275 2445.120 1429.595 ;
        RECT 2448.260 1429.445 2448.600 1429.795 ;
        RECT 2448.350 1429.440 2448.520 1429.445 ;
        RECT 2443.800 1428.475 2443.940 1429.245 ;
        RECT 2444.920 1428.475 2445.060 1429.275 ;
        RECT 2449.550 1428.860 2449.710 1434.035 ;
        RECT 2450.665 1433.945 2450.990 1434.035 ;
        RECT 2449.865 1433.510 2450.185 1433.835 ;
        RECT 2449.895 1433.335 2450.065 1433.510 ;
        RECT 2449.895 1433.160 2450.070 1433.335 ;
        RECT 2449.895 1432.985 2450.870 1433.160 ;
        RECT 2449.865 1428.860 2450.185 1428.980 ;
        RECT 2449.550 1428.690 2450.185 1428.860 ;
        RECT 2449.865 1428.660 2450.185 1428.690 ;
        RECT 2450.695 1428.610 2450.870 1432.985 ;
        RECT 2443.140 1428.245 2443.580 1428.475 ;
        RECT 2443.140 1428.155 2443.400 1428.245 ;
        RECT 2443.740 1428.155 2444.000 1428.475 ;
        RECT 2444.860 1428.155 2445.120 1428.475 ;
        RECT 2446.290 1428.125 2446.570 1428.500 ;
        RECT 2450.640 1428.260 2450.990 1428.610 ;
        RECT 2439.880 1427.865 2442.460 1428.005 ;
        RECT 2416.020 1427.150 2416.280 1427.470 ;
        RECT 2434.420 1427.150 2434.680 1427.470 ;
        RECT 2378.760 1421.210 2379.020 1421.530 ;
        RECT 2397.160 1421.210 2397.420 1421.530 ;
        RECT 2416.080 1421.190 2416.220 1427.150 ;
        RECT 2416.020 1420.870 2416.280 1421.190 ;
        RECT 2434.480 1420.850 2434.620 1427.150 ;
        RECT 2434.420 1420.530 2434.680 1420.850 ;
        RECT 2369.230 1335.690 2446.725 1335.860 ;
        RECT 2369.230 1333.895 2369.400 1335.690 ;
        RECT 2446.555 1334.915 2446.725 1335.690 ;
        RECT 2369.540 1334.515 2369.830 1334.640 ;
        RECT 2369.540 1334.510 2369.860 1334.515 ;
        RECT 2369.540 1334.340 2370.795 1334.510 ;
        RECT 2377.015 1334.345 2377.385 1334.715 ;
        RECT 2392.275 1334.345 2392.645 1334.715 ;
        RECT 2407.535 1334.345 2407.905 1334.715 ;
        RECT 2422.795 1334.345 2423.165 1334.715 ;
        RECT 2438.055 1334.345 2438.425 1334.715 ;
        RECT 2446.525 1334.565 2446.875 1334.915 ;
        RECT 2369.540 1334.290 2369.830 1334.340 ;
        RECT 2370.625 1334.145 2370.795 1334.340 ;
        RECT 2377.685 1334.145 2378.035 1334.245 ;
        RECT 2383.125 1334.205 2383.450 1334.270 ;
        RECT 2370.625 1333.975 2378.035 1334.145 ;
        RECT 2377.685 1333.895 2378.035 1333.975 ;
        RECT 2382.010 1334.035 2383.450 1334.205 ;
        RECT 2369.165 1333.545 2369.455 1333.895 ;
        RECT 2374.985 1330.305 2377.425 1330.445 ;
        RECT 2374.985 1330.155 2375.125 1330.305 ;
        RECT 2374.685 1330.065 2375.125 1330.155 ;
        RECT 2372.345 1329.925 2375.125 1330.065 ;
        RECT 2371.835 1329.785 2372.095 1329.875 ;
        RECT 2372.345 1329.785 2372.485 1329.925 ;
        RECT 2374.685 1329.835 2374.945 1329.925 ;
        RECT 2375.285 1329.835 2375.545 1330.155 ;
        RECT 2375.285 1329.785 2375.485 1329.835 ;
        RECT 2371.835 1329.645 2372.485 1329.785 ;
        RECT 2375.095 1329.645 2375.485 1329.785 ;
        RECT 2376.355 1329.775 2376.635 1330.155 ;
        RECT 2376.845 1329.835 2377.120 1330.155 ;
        RECT 2371.835 1329.555 2372.095 1329.645 ;
        RECT 2371.895 1328.475 2372.035 1329.555 ;
        RECT 2372.755 1329.505 2373.035 1329.620 ;
        RECT 2374.205 1329.505 2374.465 1329.595 ;
        RECT 2372.585 1329.365 2374.465 1329.505 ;
        RECT 2372.585 1329.315 2373.035 1329.365 ;
        RECT 2372.525 1329.245 2373.035 1329.315 ;
        RECT 2374.205 1329.275 2374.465 1329.365 ;
        RECT 2372.525 1329.055 2372.785 1329.245 ;
        RECT 2373.700 1329.055 2374.005 1329.060 ;
        RECT 2372.515 1328.685 2372.795 1329.055 ;
        RECT 2373.005 1328.945 2373.265 1329.035 ;
        RECT 2373.595 1328.945 2374.005 1329.055 ;
        RECT 2373.005 1328.805 2374.005 1328.945 ;
        RECT 2373.005 1328.715 2373.265 1328.805 ;
        RECT 2373.595 1328.685 2374.005 1328.805 ;
        RECT 2374.435 1328.685 2374.715 1329.060 ;
        RECT 2375.095 1328.525 2375.235 1329.645 ;
        RECT 2376.425 1329.315 2376.565 1329.775 ;
        RECT 2375.875 1328.685 2376.155 1329.155 ;
        RECT 2376.365 1329.055 2376.625 1329.315 ;
        RECT 2376.355 1328.685 2376.635 1329.055 ;
        RECT 2375.095 1328.475 2375.405 1328.525 ;
        RECT 2376.905 1328.515 2377.045 1329.835 ;
        RECT 2377.285 1329.315 2377.425 1330.305 ;
        RECT 2377.595 1329.555 2377.855 1329.875 ;
        RECT 2379.455 1329.835 2379.715 1330.155 ;
        RECT 2377.225 1328.995 2377.485 1329.315 ;
        RECT 2377.655 1328.515 2377.795 1329.555 ;
        RECT 2379.515 1329.055 2379.655 1329.835 ;
        RECT 2380.750 1329.345 2381.040 1329.360 ;
        RECT 2378.765 1328.945 2379.025 1329.035 ;
        RECT 2378.105 1328.805 2379.025 1328.945 ;
        RECT 2376.565 1328.495 2377.045 1328.515 ;
        RECT 2371.835 1328.155 2372.095 1328.475 ;
        RECT 2374.565 1328.385 2374.825 1328.475 ;
        RECT 2375.035 1328.445 2375.405 1328.475 ;
        RECT 2374.565 1328.155 2374.885 1328.385 ;
        RECT 2374.745 1328.005 2374.885 1328.155 ;
        RECT 2375.035 1328.150 2375.445 1328.445 ;
        RECT 2375.635 1328.155 2375.915 1328.495 ;
        RECT 2376.365 1328.245 2377.045 1328.495 ;
        RECT 2377.585 1328.445 2377.865 1328.515 ;
        RECT 2376.365 1328.145 2376.845 1328.245 ;
        RECT 2377.535 1328.185 2377.910 1328.445 ;
        RECT 2377.585 1328.145 2377.865 1328.185 ;
        RECT 2378.105 1328.005 2378.245 1328.805 ;
        RECT 2378.765 1328.715 2379.025 1328.805 ;
        RECT 2379.345 1328.685 2379.655 1329.055 ;
        RECT 2380.720 1328.995 2381.060 1329.345 ;
        RECT 2380.750 1328.980 2381.040 1328.995 ;
        RECT 2382.010 1328.860 2382.170 1334.035 ;
        RECT 2383.125 1333.945 2383.450 1334.035 ;
        RECT 2385.505 1334.180 2385.855 1334.300 ;
        RECT 2392.945 1334.180 2393.295 1334.255 ;
        RECT 2398.385 1334.205 2398.710 1334.270 ;
        RECT 2385.505 1333.980 2393.295 1334.180 ;
        RECT 2385.505 1333.950 2385.855 1333.980 ;
        RECT 2392.945 1333.905 2393.295 1333.980 ;
        RECT 2397.270 1334.035 2398.710 1334.205 ;
        RECT 2382.325 1333.510 2382.645 1333.835 ;
        RECT 2382.355 1333.335 2382.525 1333.510 ;
        RECT 2382.355 1333.160 2382.530 1333.335 ;
        RECT 2382.355 1332.985 2383.330 1333.160 ;
        RECT 2382.325 1328.860 2382.645 1328.980 ;
        RECT 2382.010 1328.690 2382.645 1328.860 ;
        RECT 2379.415 1328.500 2379.655 1328.685 ;
        RECT 2382.325 1328.660 2382.645 1328.690 ;
        RECT 2383.155 1328.610 2383.330 1332.985 ;
        RECT 2390.245 1330.305 2392.685 1330.445 ;
        RECT 2390.245 1330.155 2390.385 1330.305 ;
        RECT 2389.945 1330.065 2390.385 1330.155 ;
        RECT 2387.605 1329.925 2390.385 1330.065 ;
        RECT 2387.095 1329.785 2387.355 1329.875 ;
        RECT 2387.605 1329.785 2387.745 1329.925 ;
        RECT 2389.945 1329.835 2390.205 1329.925 ;
        RECT 2390.545 1329.835 2390.805 1330.155 ;
        RECT 2390.545 1329.785 2390.745 1329.835 ;
        RECT 2387.095 1329.645 2387.745 1329.785 ;
        RECT 2390.355 1329.645 2390.745 1329.785 ;
        RECT 2391.615 1329.775 2391.895 1330.155 ;
        RECT 2392.105 1329.835 2392.380 1330.155 ;
        RECT 2387.095 1329.555 2387.355 1329.645 ;
        RECT 2385.660 1329.070 2385.920 1329.390 ;
        RECT 2379.415 1328.435 2379.725 1328.500 ;
        RECT 2379.415 1328.245 2379.730 1328.435 ;
        RECT 2383.100 1328.260 2383.450 1328.610 ;
        RECT 2379.445 1328.235 2379.730 1328.245 ;
        RECT 2379.445 1328.125 2379.725 1328.235 ;
        RECT 2374.745 1327.865 2378.245 1328.005 ;
        RECT 2385.720 1317.830 2385.860 1329.070 ;
        RECT 2387.155 1328.475 2387.295 1329.555 ;
        RECT 2388.015 1329.505 2388.295 1329.620 ;
        RECT 2389.465 1329.505 2389.725 1329.595 ;
        RECT 2387.845 1329.365 2389.725 1329.505 ;
        RECT 2387.845 1329.315 2388.295 1329.365 ;
        RECT 2387.785 1329.245 2388.295 1329.315 ;
        RECT 2389.465 1329.275 2389.725 1329.365 ;
        RECT 2387.785 1329.055 2388.045 1329.245 ;
        RECT 2388.960 1329.055 2389.265 1329.060 ;
        RECT 2387.775 1328.685 2388.055 1329.055 ;
        RECT 2388.265 1328.945 2388.525 1329.035 ;
        RECT 2388.855 1328.945 2389.265 1329.055 ;
        RECT 2388.265 1328.805 2389.265 1328.945 ;
        RECT 2388.265 1328.715 2388.525 1328.805 ;
        RECT 2388.855 1328.685 2389.265 1328.805 ;
        RECT 2389.695 1328.685 2389.975 1329.060 ;
        RECT 2390.355 1328.525 2390.495 1329.645 ;
        RECT 2391.685 1329.315 2391.825 1329.775 ;
        RECT 2391.135 1328.685 2391.415 1329.155 ;
        RECT 2391.625 1329.055 2391.885 1329.315 ;
        RECT 2391.615 1328.685 2391.895 1329.055 ;
        RECT 2390.355 1328.475 2390.665 1328.525 ;
        RECT 2392.165 1328.515 2392.305 1329.835 ;
        RECT 2392.545 1329.315 2392.685 1330.305 ;
        RECT 2392.855 1329.555 2393.115 1329.875 ;
        RECT 2394.715 1329.835 2394.975 1330.155 ;
        RECT 2392.485 1328.995 2392.745 1329.315 ;
        RECT 2392.915 1328.515 2393.055 1329.555 ;
        RECT 2394.775 1329.055 2394.915 1329.835 ;
        RECT 2396.010 1329.345 2396.300 1329.360 ;
        RECT 2394.025 1328.945 2394.285 1329.035 ;
        RECT 2393.365 1328.805 2394.285 1328.945 ;
        RECT 2391.825 1328.495 2392.305 1328.515 ;
        RECT 2387.095 1328.155 2387.355 1328.475 ;
        RECT 2389.825 1328.385 2390.085 1328.475 ;
        RECT 2390.295 1328.445 2390.665 1328.475 ;
        RECT 2389.825 1328.155 2390.145 1328.385 ;
        RECT 2390.005 1328.005 2390.145 1328.155 ;
        RECT 2390.295 1328.150 2390.705 1328.445 ;
        RECT 2390.895 1328.155 2391.175 1328.495 ;
        RECT 2391.625 1328.245 2392.305 1328.495 ;
        RECT 2392.845 1328.445 2393.125 1328.515 ;
        RECT 2391.625 1328.145 2392.105 1328.245 ;
        RECT 2392.795 1328.185 2393.170 1328.445 ;
        RECT 2392.845 1328.145 2393.125 1328.185 ;
        RECT 2393.365 1328.005 2393.505 1328.805 ;
        RECT 2394.025 1328.715 2394.285 1328.805 ;
        RECT 2394.605 1328.685 2394.915 1329.055 ;
        RECT 2395.980 1328.995 2396.320 1329.345 ;
        RECT 2396.010 1328.980 2396.300 1328.995 ;
        RECT 2397.270 1328.860 2397.430 1334.035 ;
        RECT 2398.385 1333.945 2398.710 1334.035 ;
        RECT 2400.765 1334.180 2401.115 1334.300 ;
        RECT 2408.205 1334.180 2408.555 1334.255 ;
        RECT 2413.645 1334.205 2413.970 1334.270 ;
        RECT 2400.765 1333.980 2408.555 1334.180 ;
        RECT 2400.765 1333.950 2401.115 1333.980 ;
        RECT 2408.205 1333.905 2408.555 1333.980 ;
        RECT 2412.530 1334.035 2413.970 1334.205 ;
        RECT 2397.585 1333.510 2397.905 1333.835 ;
        RECT 2397.615 1333.335 2397.785 1333.510 ;
        RECT 2397.615 1333.160 2397.790 1333.335 ;
        RECT 2397.615 1332.985 2398.590 1333.160 ;
        RECT 2397.585 1328.860 2397.905 1328.980 ;
        RECT 2397.270 1328.690 2397.905 1328.860 ;
        RECT 2394.675 1328.500 2394.915 1328.685 ;
        RECT 2397.585 1328.660 2397.905 1328.690 ;
        RECT 2398.415 1328.610 2398.590 1332.985 ;
        RECT 2405.505 1330.305 2407.945 1330.445 ;
        RECT 2405.505 1330.155 2405.645 1330.305 ;
        RECT 2405.205 1330.065 2405.645 1330.155 ;
        RECT 2402.865 1329.925 2405.645 1330.065 ;
        RECT 2402.355 1329.785 2402.615 1329.875 ;
        RECT 2402.865 1329.785 2403.005 1329.925 ;
        RECT 2405.205 1329.835 2405.465 1329.925 ;
        RECT 2405.805 1329.835 2406.065 1330.155 ;
        RECT 2405.805 1329.785 2406.005 1329.835 ;
        RECT 2402.355 1329.645 2403.005 1329.785 ;
        RECT 2405.615 1329.645 2406.005 1329.785 ;
        RECT 2406.875 1329.775 2407.155 1330.155 ;
        RECT 2407.365 1329.835 2407.640 1330.155 ;
        RECT 2402.355 1329.555 2402.615 1329.645 ;
        RECT 2394.675 1328.435 2394.985 1328.500 ;
        RECT 2394.675 1328.245 2394.990 1328.435 ;
        RECT 2398.360 1328.260 2398.710 1328.610 ;
        RECT 2402.415 1328.475 2402.555 1329.555 ;
        RECT 2403.275 1329.505 2403.555 1329.620 ;
        RECT 2404.725 1329.505 2404.985 1329.595 ;
        RECT 2403.105 1329.365 2404.985 1329.505 ;
        RECT 2403.105 1329.315 2403.555 1329.365 ;
        RECT 2403.045 1329.245 2403.555 1329.315 ;
        RECT 2404.725 1329.275 2404.985 1329.365 ;
        RECT 2403.045 1329.055 2403.305 1329.245 ;
        RECT 2404.220 1329.055 2404.525 1329.060 ;
        RECT 2403.035 1328.685 2403.315 1329.055 ;
        RECT 2403.525 1328.945 2403.785 1329.035 ;
        RECT 2404.115 1328.945 2404.525 1329.055 ;
        RECT 2403.525 1328.805 2404.525 1328.945 ;
        RECT 2403.525 1328.715 2403.785 1328.805 ;
        RECT 2404.115 1328.685 2404.525 1328.805 ;
        RECT 2404.955 1328.685 2405.235 1329.060 ;
        RECT 2405.615 1328.525 2405.755 1329.645 ;
        RECT 2406.945 1329.315 2407.085 1329.775 ;
        RECT 2406.395 1328.685 2406.675 1329.155 ;
        RECT 2406.885 1329.055 2407.145 1329.315 ;
        RECT 2406.875 1328.685 2407.155 1329.055 ;
        RECT 2405.615 1328.475 2405.925 1328.525 ;
        RECT 2407.425 1328.515 2407.565 1329.835 ;
        RECT 2407.805 1329.315 2407.945 1330.305 ;
        RECT 2408.115 1329.555 2408.375 1329.875 ;
        RECT 2409.975 1329.835 2410.235 1330.155 ;
        RECT 2407.745 1328.995 2408.005 1329.315 ;
        RECT 2408.175 1328.515 2408.315 1329.555 ;
        RECT 2410.035 1329.055 2410.175 1329.835 ;
        RECT 2411.270 1329.345 2411.560 1329.360 ;
        RECT 2409.285 1328.945 2409.545 1329.035 ;
        RECT 2408.625 1328.805 2409.545 1328.945 ;
        RECT 2407.085 1328.495 2407.565 1328.515 ;
        RECT 2394.705 1328.235 2394.990 1328.245 ;
        RECT 2394.705 1328.125 2394.985 1328.235 ;
        RECT 2402.355 1328.155 2402.615 1328.475 ;
        RECT 2405.085 1328.385 2405.345 1328.475 ;
        RECT 2405.555 1328.445 2405.925 1328.475 ;
        RECT 2405.085 1328.155 2405.405 1328.385 ;
        RECT 2390.005 1327.865 2393.505 1328.005 ;
        RECT 2405.265 1328.005 2405.405 1328.155 ;
        RECT 2405.555 1328.150 2405.965 1328.445 ;
        RECT 2406.155 1328.155 2406.435 1328.495 ;
        RECT 2406.885 1328.245 2407.565 1328.495 ;
        RECT 2408.105 1328.445 2408.385 1328.515 ;
        RECT 2406.885 1328.145 2407.365 1328.245 ;
        RECT 2408.055 1328.185 2408.430 1328.445 ;
        RECT 2408.105 1328.145 2408.385 1328.185 ;
        RECT 2408.625 1328.005 2408.765 1328.805 ;
        RECT 2409.285 1328.715 2409.545 1328.805 ;
        RECT 2409.865 1328.685 2410.175 1329.055 ;
        RECT 2411.240 1328.995 2411.580 1329.345 ;
        RECT 2411.270 1328.980 2411.560 1328.995 ;
        RECT 2412.530 1328.860 2412.690 1334.035 ;
        RECT 2413.645 1333.945 2413.970 1334.035 ;
        RECT 2415.980 1334.180 2416.330 1334.300 ;
        RECT 2423.470 1334.180 2423.820 1334.255 ;
        RECT 2428.905 1334.205 2429.230 1334.270 ;
        RECT 2415.980 1333.980 2423.820 1334.180 ;
        RECT 2415.980 1333.950 2416.330 1333.980 ;
        RECT 2423.470 1333.905 2423.820 1333.980 ;
        RECT 2427.790 1334.035 2429.230 1334.205 ;
        RECT 2412.845 1333.510 2413.165 1333.835 ;
        RECT 2412.875 1333.335 2413.045 1333.510 ;
        RECT 2412.875 1333.160 2413.050 1333.335 ;
        RECT 2412.875 1332.985 2413.850 1333.160 ;
        RECT 2412.845 1328.860 2413.165 1328.980 ;
        RECT 2412.530 1328.690 2413.165 1328.860 ;
        RECT 2409.935 1328.500 2410.175 1328.685 ;
        RECT 2412.845 1328.660 2413.165 1328.690 ;
        RECT 2413.675 1328.610 2413.850 1332.985 ;
        RECT 2420.765 1330.305 2423.205 1330.445 ;
        RECT 2420.765 1330.155 2420.905 1330.305 ;
        RECT 2420.465 1330.065 2420.905 1330.155 ;
        RECT 2418.125 1329.925 2420.905 1330.065 ;
        RECT 2417.615 1329.785 2417.875 1329.875 ;
        RECT 2418.125 1329.785 2418.265 1329.925 ;
        RECT 2420.465 1329.835 2420.725 1329.925 ;
        RECT 2421.065 1329.835 2421.325 1330.155 ;
        RECT 2421.065 1329.785 2421.265 1329.835 ;
        RECT 2417.615 1329.645 2418.265 1329.785 ;
        RECT 2420.875 1329.645 2421.265 1329.785 ;
        RECT 2422.135 1329.775 2422.415 1330.155 ;
        RECT 2422.625 1329.835 2422.900 1330.155 ;
        RECT 2417.615 1329.555 2417.875 1329.645 ;
        RECT 2409.935 1328.435 2410.245 1328.500 ;
        RECT 2409.935 1328.245 2410.250 1328.435 ;
        RECT 2413.620 1328.260 2413.970 1328.610 ;
        RECT 2417.675 1328.475 2417.815 1329.555 ;
        RECT 2418.535 1329.505 2418.815 1329.620 ;
        RECT 2419.985 1329.505 2420.245 1329.595 ;
        RECT 2418.365 1329.365 2420.245 1329.505 ;
        RECT 2418.365 1329.315 2418.815 1329.365 ;
        RECT 2418.305 1329.245 2418.815 1329.315 ;
        RECT 2419.985 1329.275 2420.245 1329.365 ;
        RECT 2418.305 1329.055 2418.565 1329.245 ;
        RECT 2419.480 1329.055 2419.785 1329.060 ;
        RECT 2418.295 1328.685 2418.575 1329.055 ;
        RECT 2418.785 1328.945 2419.045 1329.035 ;
        RECT 2419.375 1328.945 2419.785 1329.055 ;
        RECT 2418.785 1328.805 2419.785 1328.945 ;
        RECT 2418.785 1328.715 2419.045 1328.805 ;
        RECT 2419.375 1328.685 2419.785 1328.805 ;
        RECT 2420.215 1328.685 2420.495 1329.060 ;
        RECT 2420.875 1328.525 2421.015 1329.645 ;
        RECT 2422.205 1329.315 2422.345 1329.775 ;
        RECT 2421.655 1328.685 2421.935 1329.155 ;
        RECT 2422.145 1329.055 2422.405 1329.315 ;
        RECT 2422.135 1328.685 2422.415 1329.055 ;
        RECT 2420.875 1328.475 2421.185 1328.525 ;
        RECT 2422.685 1328.515 2422.825 1329.835 ;
        RECT 2423.065 1329.315 2423.205 1330.305 ;
        RECT 2423.375 1329.555 2423.635 1329.875 ;
        RECT 2425.235 1329.835 2425.495 1330.155 ;
        RECT 2423.005 1328.995 2423.265 1329.315 ;
        RECT 2423.435 1328.515 2423.575 1329.555 ;
        RECT 2425.295 1329.055 2425.435 1329.835 ;
        RECT 2426.530 1329.345 2426.820 1329.360 ;
        RECT 2424.545 1328.945 2424.805 1329.035 ;
        RECT 2423.885 1328.805 2424.805 1328.945 ;
        RECT 2422.345 1328.495 2422.825 1328.515 ;
        RECT 2409.965 1328.235 2410.250 1328.245 ;
        RECT 2409.965 1328.125 2410.245 1328.235 ;
        RECT 2417.615 1328.155 2417.875 1328.475 ;
        RECT 2420.345 1328.385 2420.605 1328.475 ;
        RECT 2420.815 1328.445 2421.185 1328.475 ;
        RECT 2420.345 1328.155 2420.665 1328.385 ;
        RECT 2405.265 1327.865 2408.765 1328.005 ;
        RECT 2420.525 1328.005 2420.665 1328.155 ;
        RECT 2420.815 1328.150 2421.225 1328.445 ;
        RECT 2421.415 1328.155 2421.695 1328.495 ;
        RECT 2422.145 1328.245 2422.825 1328.495 ;
        RECT 2423.365 1328.445 2423.645 1328.515 ;
        RECT 2422.145 1328.145 2422.625 1328.245 ;
        RECT 2423.315 1328.185 2423.690 1328.445 ;
        RECT 2423.365 1328.145 2423.645 1328.185 ;
        RECT 2423.885 1328.005 2424.025 1328.805 ;
        RECT 2424.545 1328.715 2424.805 1328.805 ;
        RECT 2425.125 1328.685 2425.435 1329.055 ;
        RECT 2426.500 1328.995 2426.840 1329.345 ;
        RECT 2426.530 1328.980 2426.820 1328.995 ;
        RECT 2427.790 1328.860 2427.950 1334.035 ;
        RECT 2428.905 1333.945 2429.230 1334.035 ;
        RECT 2431.240 1334.180 2431.590 1334.300 ;
        RECT 2438.725 1334.180 2439.075 1334.255 ;
        RECT 2444.165 1334.205 2444.490 1334.270 ;
        RECT 2431.240 1333.980 2439.075 1334.180 ;
        RECT 2431.240 1333.950 2431.590 1333.980 ;
        RECT 2438.725 1333.905 2439.075 1333.980 ;
        RECT 2443.050 1334.035 2444.490 1334.205 ;
        RECT 2428.105 1333.510 2428.425 1333.835 ;
        RECT 2428.135 1333.335 2428.305 1333.510 ;
        RECT 2428.135 1333.160 2428.310 1333.335 ;
        RECT 2428.135 1332.985 2429.110 1333.160 ;
        RECT 2428.105 1328.860 2428.425 1328.980 ;
        RECT 2427.790 1328.690 2428.425 1328.860 ;
        RECT 2425.195 1328.500 2425.435 1328.685 ;
        RECT 2428.105 1328.660 2428.425 1328.690 ;
        RECT 2428.935 1328.610 2429.110 1332.985 ;
        RECT 2436.025 1330.305 2438.465 1330.445 ;
        RECT 2436.025 1330.155 2436.165 1330.305 ;
        RECT 2435.725 1330.065 2436.165 1330.155 ;
        RECT 2433.385 1329.925 2436.165 1330.065 ;
        RECT 2432.875 1329.785 2433.135 1329.875 ;
        RECT 2433.385 1329.785 2433.525 1329.925 ;
        RECT 2435.725 1329.835 2435.985 1329.925 ;
        RECT 2436.325 1329.835 2436.585 1330.155 ;
        RECT 2436.325 1329.785 2436.525 1329.835 ;
        RECT 2432.875 1329.645 2433.525 1329.785 ;
        RECT 2436.135 1329.645 2436.525 1329.785 ;
        RECT 2437.395 1329.775 2437.675 1330.155 ;
        RECT 2437.885 1329.835 2438.160 1330.155 ;
        RECT 2432.875 1329.555 2433.135 1329.645 ;
        RECT 2425.195 1328.435 2425.505 1328.500 ;
        RECT 2425.195 1328.245 2425.510 1328.435 ;
        RECT 2428.880 1328.260 2429.230 1328.610 ;
        RECT 2432.935 1328.475 2433.075 1329.555 ;
        RECT 2433.795 1329.505 2434.075 1329.620 ;
        RECT 2435.245 1329.505 2435.505 1329.595 ;
        RECT 2433.625 1329.365 2435.505 1329.505 ;
        RECT 2433.625 1329.315 2434.075 1329.365 ;
        RECT 2433.565 1329.245 2434.075 1329.315 ;
        RECT 2435.245 1329.275 2435.505 1329.365 ;
        RECT 2433.565 1329.055 2433.825 1329.245 ;
        RECT 2434.740 1329.055 2435.045 1329.060 ;
        RECT 2433.555 1328.685 2433.835 1329.055 ;
        RECT 2434.045 1328.945 2434.305 1329.035 ;
        RECT 2434.635 1328.945 2435.045 1329.055 ;
        RECT 2434.045 1328.805 2435.045 1328.945 ;
        RECT 2434.045 1328.715 2434.305 1328.805 ;
        RECT 2434.635 1328.685 2435.045 1328.805 ;
        RECT 2435.475 1328.685 2435.755 1329.060 ;
        RECT 2436.135 1328.525 2436.275 1329.645 ;
        RECT 2437.465 1329.315 2437.605 1329.775 ;
        RECT 2436.915 1328.685 2437.195 1329.155 ;
        RECT 2437.405 1329.055 2437.665 1329.315 ;
        RECT 2437.395 1328.685 2437.675 1329.055 ;
        RECT 2436.135 1328.475 2436.445 1328.525 ;
        RECT 2437.945 1328.515 2438.085 1329.835 ;
        RECT 2438.325 1329.315 2438.465 1330.305 ;
        RECT 2438.635 1329.555 2438.895 1329.875 ;
        RECT 2440.495 1329.835 2440.755 1330.155 ;
        RECT 2438.265 1328.995 2438.525 1329.315 ;
        RECT 2438.695 1328.515 2438.835 1329.555 ;
        RECT 2440.555 1329.055 2440.695 1329.835 ;
        RECT 2441.790 1329.345 2442.080 1329.360 ;
        RECT 2439.805 1328.945 2440.065 1329.035 ;
        RECT 2439.145 1328.805 2440.065 1328.945 ;
        RECT 2437.605 1328.495 2438.085 1328.515 ;
        RECT 2425.225 1328.235 2425.510 1328.245 ;
        RECT 2425.225 1328.125 2425.505 1328.235 ;
        RECT 2432.875 1328.155 2433.135 1328.475 ;
        RECT 2435.605 1328.385 2435.865 1328.475 ;
        RECT 2436.075 1328.445 2436.445 1328.475 ;
        RECT 2435.605 1328.155 2435.925 1328.385 ;
        RECT 2420.525 1327.865 2424.025 1328.005 ;
        RECT 2435.785 1328.005 2435.925 1328.155 ;
        RECT 2436.075 1328.150 2436.485 1328.445 ;
        RECT 2436.675 1328.155 2436.955 1328.495 ;
        RECT 2437.405 1328.245 2438.085 1328.495 ;
        RECT 2438.625 1328.445 2438.905 1328.515 ;
        RECT 2437.405 1328.145 2437.885 1328.245 ;
        RECT 2438.575 1328.185 2438.950 1328.445 ;
        RECT 2438.625 1328.145 2438.905 1328.185 ;
        RECT 2439.145 1328.005 2439.285 1328.805 ;
        RECT 2439.805 1328.715 2440.065 1328.805 ;
        RECT 2440.385 1328.685 2440.695 1329.055 ;
        RECT 2441.760 1328.995 2442.100 1329.345 ;
        RECT 2441.790 1328.980 2442.080 1328.995 ;
        RECT 2443.050 1328.860 2443.210 1334.035 ;
        RECT 2444.165 1333.945 2444.490 1334.035 ;
        RECT 2443.365 1333.510 2443.685 1333.835 ;
        RECT 2443.395 1333.335 2443.565 1333.510 ;
        RECT 2443.395 1333.160 2443.570 1333.335 ;
        RECT 2443.395 1332.985 2444.370 1333.160 ;
        RECT 2443.365 1328.860 2443.685 1328.980 ;
        RECT 2443.050 1328.690 2443.685 1328.860 ;
        RECT 2440.455 1328.500 2440.695 1328.685 ;
        RECT 2443.365 1328.660 2443.685 1328.690 ;
        RECT 2444.195 1328.610 2444.370 1332.985 ;
        RECT 2459.780 1330.070 2459.920 1441.950 ;
        RECT 2464.840 1428.330 2464.980 1449.090 ;
        RECT 2464.780 1428.010 2465.040 1428.330 ;
        RECT 2508.080 1420.510 2508.220 2166.490 ;
        RECT 2514.920 2159.690 2515.180 2160.010 ;
        RECT 2508.020 1420.190 2508.280 1420.510 ;
        RECT 2459.720 1329.750 2459.980 1330.070 ;
        RECT 2440.455 1328.435 2440.765 1328.500 ;
        RECT 2440.455 1328.245 2440.770 1328.435 ;
        RECT 2444.140 1328.260 2444.490 1328.610 ;
        RECT 2440.485 1328.235 2440.770 1328.245 ;
        RECT 2440.485 1328.125 2440.765 1328.235 ;
        RECT 2435.785 1327.865 2439.285 1328.005 ;
        RECT 2400.840 1327.145 2401.100 1327.465 ;
        RECT 2416.020 1327.145 2416.280 1327.465 ;
        RECT 2431.200 1327.145 2431.460 1327.465 ;
        RECT 2400.900 1317.830 2401.040 1327.145 ;
        RECT 2416.080 1317.830 2416.220 1327.145 ;
        RECT 2431.260 1317.830 2431.400 1327.145 ;
        RECT 2385.660 1317.510 2385.920 1317.830 ;
        RECT 2400.840 1317.510 2401.100 1317.830 ;
        RECT 2416.020 1317.510 2416.280 1317.830 ;
        RECT 2431.200 1317.510 2431.460 1317.830 ;
        RECT 2475.360 1317.570 2475.620 1317.830 ;
        RECT 2474.040 1317.510 2475.620 1317.570 ;
        RECT 2474.040 1317.490 2475.560 1317.510 ;
        RECT 2473.980 1317.430 2475.560 1317.490 ;
        RECT 2473.980 1317.170 2474.240 1317.430 ;
        RECT 2514.980 1316.810 2515.120 2159.690 ;
        RECT 2523.560 2134.955 2523.840 2135.325 ;
        RECT 2523.560 2127.425 2523.840 2127.795 ;
        RECT 2523.560 2121.445 2523.840 2121.815 ;
        RECT 2523.560 2115.500 2523.840 2115.870 ;
        RECT 2523.560 2109.855 2523.840 2110.225 ;
        RECT 2523.560 2103.850 2523.840 2104.220 ;
        RECT 2577.080 2049.170 2577.220 2229.390 ;
        RECT 2618.420 2229.050 2618.680 2229.370 ;
        RECT 2604.620 2228.710 2604.880 2229.030 ;
        RECT 2577.020 2048.850 2577.280 2049.170 ;
        RECT 2577.020 2021.650 2577.280 2021.970 ;
        RECT 2523.560 1982.700 2523.840 1983.070 ;
        RECT 2523.560 1975.170 2523.840 1975.540 ;
        RECT 2523.560 1969.190 2523.840 1969.560 ;
        RECT 2523.560 1963.245 2523.840 1963.615 ;
        RECT 2523.560 1957.600 2523.840 1957.970 ;
        RECT 2523.560 1951.595 2523.840 1951.965 ;
        RECT 2577.080 1939.010 2577.220 2021.650 ;
        RECT 2583.920 2014.850 2584.180 2015.170 ;
        RECT 2577.020 1938.690 2577.280 1939.010 ;
        RECT 2577.020 1828.530 2577.280 1828.850 ;
        RECT 2523.560 1805.730 2523.840 1806.100 ;
        RECT 2523.560 1798.200 2523.840 1798.570 ;
        RECT 2523.560 1792.220 2523.840 1792.590 ;
        RECT 2523.560 1786.275 2523.840 1786.645 ;
        RECT 2523.560 1780.630 2523.840 1781.000 ;
        RECT 2523.560 1769.160 2523.840 1769.530 ;
        RECT 2577.080 1696.930 2577.220 1828.530 ;
        RECT 2583.980 1773.090 2584.120 2014.850 ;
        RECT 2590.820 1994.110 2591.080 1994.430 ;
        RECT 2583.920 1772.770 2584.180 1773.090 ;
        RECT 2577.020 1696.610 2577.280 1696.930 ;
        RECT 2523.560 1624.595 2523.840 1624.965 ;
        RECT 2523.560 1618.180 2523.840 1618.550 ;
        RECT 2523.560 1588.935 2523.840 1589.305 ;
        RECT 2523.560 1581.405 2523.840 1581.775 ;
        RECT 2523.560 1575.425 2523.840 1575.795 ;
        RECT 2523.560 1567.010 2523.840 1567.380 ;
        RECT 2590.880 1517.410 2591.020 1994.110 ;
        RECT 2597.720 1980.170 2597.980 1980.490 ;
        RECT 2590.820 1517.090 2591.080 1517.410 ;
        RECT 2523.560 1437.310 2523.840 1437.680 ;
        RECT 2523.560 1430.895 2523.840 1431.265 ;
        RECT 2523.560 1416.705 2523.840 1417.075 ;
        RECT 2523.560 1409.175 2523.840 1409.545 ;
        RECT 2523.560 1403.195 2523.840 1403.565 ;
        RECT 2523.560 1394.780 2523.840 1395.150 ;
        RECT 2597.780 1317.150 2597.920 1980.170 ;
        RECT 2604.680 1869.990 2604.820 2228.710 ;
        RECT 2611.520 2138.950 2611.780 2139.270 ;
        RECT 2604.620 1869.670 2604.880 1869.990 ;
        RECT 2611.580 1862.850 2611.720 2138.950 ;
        RECT 2611.520 1862.530 2611.780 1862.850 ;
        RECT 2604.620 1835.330 2604.880 1835.650 ;
        RECT 2604.680 1773.430 2604.820 1835.330 ;
        RECT 2611.520 1807.790 2611.780 1808.110 ;
        RECT 2604.620 1773.110 2604.880 1773.430 ;
        RECT 2611.580 1421.190 2611.720 1807.790 ;
        RECT 2618.480 1690.470 2618.620 2229.050 ;
        RECT 2677.300 2228.370 2677.560 2228.690 ;
        RECT 2677.360 2224.125 2677.500 2228.370 ;
        RECT 2677.290 2223.755 2677.570 2224.125 ;
        RECT 2695.150 2223.875 2695.430 2224.245 ;
        RECT 2677.290 2216.955 2677.570 2217.325 ;
        RECT 2677.360 2215.090 2677.500 2216.955 ;
        RECT 2695.220 2215.890 2695.360 2223.875 ;
        RECT 2695.610 2217.075 2695.890 2217.445 ;
        RECT 2695.680 2216.570 2695.820 2217.075 ;
        RECT 2695.620 2216.250 2695.880 2216.570 ;
        RECT 2698.840 2216.250 2699.100 2216.570 ;
        RECT 2702.520 2216.250 2702.780 2216.570 ;
        RECT 2695.160 2215.570 2695.420 2215.890 ;
        RECT 2677.300 2214.770 2677.560 2215.090 ;
        RECT 2698.380 2214.550 2698.640 2214.870 ;
        RECT 2694.700 2212.510 2694.960 2212.830 ;
        RECT 2698.440 2212.570 2698.580 2214.550 ;
        RECT 2694.760 2210.645 2694.900 2212.510 ;
        RECT 2697.520 2212.430 2698.580 2212.570 ;
        RECT 2677.290 2210.155 2677.570 2210.525 ;
        RECT 2694.690 2210.275 2694.970 2210.645 ;
        RECT 2677.360 2208.290 2677.500 2210.155 ;
        RECT 2677.300 2207.970 2677.560 2208.290 ;
        RECT 2694.700 2204.690 2694.960 2205.010 ;
        RECT 2694.760 2203.845 2694.900 2204.690 ;
        RECT 2677.290 2203.355 2677.570 2203.725 ;
        RECT 2694.690 2203.475 2694.970 2203.845 ;
        RECT 2697.000 2203.670 2697.260 2203.990 ;
        RECT 2697.520 2203.730 2697.660 2212.430 ;
        RECT 2697.920 2211.830 2698.180 2212.150 ;
        RECT 2697.980 2204.410 2698.120 2211.830 ;
        RECT 2697.980 2204.270 2698.580 2204.410 ;
        RECT 2677.360 2201.490 2677.500 2203.355 ;
        RECT 2677.300 2201.170 2677.560 2201.490 ;
        RECT 2677.290 2196.555 2677.570 2196.925 ;
        RECT 2694.690 2196.675 2694.970 2197.045 ;
        RECT 2677.360 2194.690 2677.500 2196.555 ;
        RECT 2694.760 2196.510 2694.900 2196.675 ;
        RECT 2694.700 2196.190 2694.960 2196.510 ;
        RECT 2677.300 2194.370 2677.560 2194.690 ;
        RECT 2697.060 2194.130 2697.200 2203.670 ;
        RECT 2697.520 2203.590 2698.120 2203.730 ;
        RECT 2697.460 2201.970 2697.720 2202.290 ;
        RECT 2697.520 2199.570 2697.660 2201.970 ;
        RECT 2697.980 2199.570 2698.120 2203.590 ;
        RECT 2698.440 2202.290 2698.580 2204.270 ;
        RECT 2698.380 2201.970 2698.640 2202.290 ;
        RECT 2697.460 2199.250 2697.720 2199.570 ;
        RECT 2697.920 2199.250 2698.180 2199.570 ;
        RECT 2697.460 2198.570 2697.720 2198.890 ;
        RECT 2697.000 2193.810 2697.260 2194.130 ;
        RECT 2694.700 2190.750 2694.960 2191.070 ;
        RECT 2694.760 2190.245 2694.900 2190.750 ;
        RECT 2677.290 2189.755 2677.570 2190.125 ;
        RECT 2694.690 2189.875 2694.970 2190.245 ;
        RECT 2677.360 2187.550 2677.500 2189.755 ;
        RECT 2677.300 2187.230 2677.560 2187.550 ;
        RECT 2697.520 2186.650 2697.660 2198.570 ;
        RECT 2698.900 2197.610 2699.040 2216.250 ;
        RECT 2701.600 2215.230 2701.860 2215.550 ;
        RECT 2697.980 2197.470 2699.040 2197.610 ;
        RECT 2697.980 2194.130 2698.120 2197.470 ;
        RECT 2697.920 2193.810 2698.180 2194.130 ;
        RECT 2698.840 2193.470 2699.100 2193.790 ;
        RECT 2698.380 2192.790 2698.640 2193.110 ;
        RECT 2697.920 2191.090 2698.180 2191.410 ;
        RECT 2697.460 2186.330 2697.720 2186.650 ;
        RECT 2694.700 2185.310 2694.960 2185.630 ;
        RECT 2694.760 2183.445 2694.900 2185.310 ;
        RECT 2677.290 2182.955 2677.570 2183.325 ;
        RECT 2694.690 2183.075 2694.970 2183.445 ;
        RECT 2677.360 2180.750 2677.500 2182.955 ;
        RECT 2677.300 2180.430 2677.560 2180.750 ;
        RECT 2694.700 2177.490 2694.960 2177.810 ;
        RECT 2694.760 2176.645 2694.900 2177.490 ;
        RECT 2677.290 2176.155 2677.570 2176.525 ;
        RECT 2694.690 2176.275 2694.970 2176.645 ;
        RECT 2677.360 2173.950 2677.500 2176.155 ;
        RECT 2677.300 2173.630 2677.560 2173.950 ;
        RECT 2694.700 2172.050 2694.960 2172.370 ;
        RECT 2694.760 2169.845 2694.900 2172.050 ;
        RECT 2697.460 2171.030 2697.720 2171.350 ;
        RECT 2677.290 2169.355 2677.570 2169.725 ;
        RECT 2694.690 2169.475 2694.970 2169.845 ;
        RECT 2677.360 2166.810 2677.500 2169.355 ;
        RECT 2677.300 2166.490 2677.560 2166.810 ;
        RECT 2697.520 2166.590 2697.660 2171.030 ;
        RECT 2697.980 2166.930 2698.120 2191.090 ;
        RECT 2698.440 2166.930 2698.580 2192.790 ;
        RECT 2698.900 2178.490 2699.040 2193.470 ;
        RECT 2701.660 2191.410 2701.800 2215.230 ;
        RECT 2702.060 2198.910 2702.320 2199.230 ;
        RECT 2702.120 2197.530 2702.260 2198.910 ;
        RECT 2702.580 2198.550 2702.720 2216.250 ;
        RECT 2721.840 2214.890 2722.100 2215.210 ;
        RECT 2721.900 2199.570 2722.040 2214.890 ;
        RECT 2731.500 2214.550 2731.760 2214.870 ;
        RECT 2721.840 2199.250 2722.100 2199.570 ;
        RECT 2702.980 2198.910 2703.240 2199.230 ;
        RECT 2702.520 2198.230 2702.780 2198.550 ;
        RECT 2702.060 2197.210 2702.320 2197.530 ;
        RECT 2702.060 2193.470 2702.320 2193.790 ;
        RECT 2702.120 2192.090 2702.260 2193.470 ;
        RECT 2702.580 2193.110 2702.720 2198.230 ;
        RECT 2703.040 2194.130 2703.180 2198.910 ;
        RECT 2703.900 2198.230 2704.160 2198.550 ;
        RECT 2702.980 2193.810 2703.240 2194.130 ;
        RECT 2702.520 2192.790 2702.780 2193.110 ;
        RECT 2702.060 2191.770 2702.320 2192.090 ;
        RECT 2701.600 2191.090 2701.860 2191.410 ;
        RECT 2701.600 2190.070 2701.860 2190.390 ;
        RECT 2701.660 2180.190 2701.800 2190.070 ;
        RECT 2701.600 2179.870 2701.860 2180.190 ;
        RECT 2702.060 2179.190 2702.320 2179.510 ;
        RECT 2702.120 2178.490 2702.260 2179.190 ;
        RECT 2698.840 2178.170 2699.100 2178.490 ;
        RECT 2702.060 2178.170 2702.320 2178.490 ;
        RECT 2702.520 2176.810 2702.780 2177.130 ;
        RECT 2702.580 2175.770 2702.720 2176.810 ;
        RECT 2702.520 2175.450 2702.780 2175.770 ;
        RECT 2697.920 2166.610 2698.180 2166.930 ;
        RECT 2698.380 2166.610 2698.640 2166.930 ;
        RECT 2697.460 2166.270 2697.720 2166.590 ;
        RECT 2694.700 2163.550 2694.960 2163.870 ;
        RECT 2697.980 2163.610 2698.120 2166.610 ;
        RECT 2694.760 2163.045 2694.900 2163.550 ;
        RECT 2697.520 2163.470 2698.120 2163.610 ;
        RECT 2677.290 2162.555 2677.570 2162.925 ;
        RECT 2694.690 2162.675 2694.970 2163.045 ;
        RECT 2677.360 2160.010 2677.500 2162.555 ;
        RECT 2677.300 2159.690 2677.560 2160.010 ;
        RECT 2697.520 2159.110 2697.660 2163.470 ;
        RECT 2697.920 2162.870 2698.180 2163.190 ;
        RECT 2697.980 2162.170 2698.120 2162.870 ;
        RECT 2697.920 2161.850 2698.180 2162.170 ;
        RECT 2698.440 2161.830 2698.580 2166.610 ;
        RECT 2702.060 2166.270 2702.320 2166.590 ;
        RECT 2703.040 2166.330 2703.180 2193.810 ;
        RECT 2703.960 2190.730 2704.100 2198.230 ;
        RECT 2706.200 2192.790 2706.460 2193.110 ;
        RECT 2706.260 2192.090 2706.400 2192.790 ;
        RECT 2706.200 2191.770 2706.460 2192.090 ;
        RECT 2703.900 2190.410 2704.160 2190.730 ;
        RECT 2731.560 2180.190 2731.700 2214.550 ;
        RECT 2703.900 2179.870 2704.160 2180.190 ;
        RECT 2731.500 2179.870 2731.760 2180.190 ;
        RECT 2703.960 2178.490 2704.100 2179.870 ;
        RECT 2703.900 2178.170 2704.160 2178.490 ;
        RECT 2704.820 2177.150 2705.080 2177.470 ;
        RECT 2704.880 2174.490 2705.020 2177.150 ;
        RECT 2702.120 2162.170 2702.260 2166.270 ;
        RECT 2702.580 2166.190 2703.180 2166.330 ;
        RECT 2703.960 2174.350 2705.020 2174.490 ;
        RECT 2702.060 2161.850 2702.320 2162.170 ;
        RECT 2698.380 2161.570 2698.640 2161.830 ;
        RECT 2698.380 2161.510 2699.040 2161.570 ;
        RECT 2698.440 2161.430 2699.040 2161.510 ;
        RECT 2702.580 2161.490 2702.720 2166.190 ;
        RECT 2702.980 2165.590 2703.240 2165.910 ;
        RECT 2703.040 2162.170 2703.180 2165.590 ;
        RECT 2702.980 2161.850 2703.240 2162.170 ;
        RECT 2703.440 2161.850 2703.700 2162.170 ;
        RECT 2698.380 2160.830 2698.640 2161.150 ;
        RECT 2697.460 2158.790 2697.720 2159.110 ;
        RECT 2694.690 2155.875 2694.970 2156.245 ;
        RECT 2694.700 2155.730 2694.960 2155.875 ;
        RECT 2697.000 2152.330 2697.260 2152.650 ;
        RECT 2697.060 2149.590 2697.200 2152.330 ;
        RECT 2697.520 2150.610 2697.660 2158.790 ;
        RECT 2697.460 2150.290 2697.720 2150.610 ;
        RECT 2697.920 2150.290 2698.180 2150.610 ;
        RECT 2694.690 2149.075 2694.970 2149.445 ;
        RECT 2697.000 2149.270 2697.260 2149.590 ;
        RECT 2694.760 2147.550 2694.900 2149.075 ;
        RECT 2694.700 2147.230 2694.960 2147.550 ;
        RECT 2697.060 2144.830 2697.200 2149.270 ;
        RECT 2697.520 2147.550 2697.660 2150.290 ;
        RECT 2697.460 2147.230 2697.720 2147.550 ;
        RECT 2697.000 2144.510 2697.260 2144.830 ;
        RECT 2697.980 2143.130 2698.120 2150.290 ;
        RECT 2698.440 2148.570 2698.580 2160.830 ;
        RECT 2698.900 2159.450 2699.040 2161.430 ;
        RECT 2702.520 2161.170 2702.780 2161.490 ;
        RECT 2702.580 2160.890 2702.720 2161.170 ;
        RECT 2701.660 2160.750 2702.720 2160.890 ;
        RECT 2698.840 2159.130 2699.100 2159.450 ;
        RECT 2698.840 2157.430 2699.100 2157.750 ;
        RECT 2698.900 2156.730 2699.040 2157.430 ;
        RECT 2698.840 2156.410 2699.100 2156.730 ;
        RECT 2701.660 2153.330 2701.800 2160.750 ;
        RECT 2702.520 2160.150 2702.780 2160.470 ;
        RECT 2702.580 2159.450 2702.720 2160.150 ;
        RECT 2702.520 2159.130 2702.780 2159.450 ;
        RECT 2702.060 2158.790 2702.320 2159.110 ;
        RECT 2701.600 2153.010 2701.860 2153.330 ;
        RECT 2699.760 2152.670 2700.020 2152.990 ;
        RECT 2698.840 2151.990 2699.100 2152.310 ;
        RECT 2699.300 2151.990 2699.560 2152.310 ;
        RECT 2698.900 2151.290 2699.040 2151.990 ;
        RECT 2698.840 2150.970 2699.100 2151.290 ;
        RECT 2699.360 2150.010 2699.500 2151.990 ;
        RECT 2699.820 2150.950 2699.960 2152.670 ;
        RECT 2702.120 2152.650 2702.260 2158.790 ;
        RECT 2703.500 2152.990 2703.640 2161.850 ;
        RECT 2703.440 2152.670 2703.700 2152.990 ;
        RECT 2702.060 2152.330 2702.320 2152.650 ;
        RECT 2699.760 2150.630 2700.020 2150.950 ;
        RECT 2702.120 2150.610 2702.260 2152.330 ;
        RECT 2703.960 2152.310 2704.100 2174.350 ;
        RECT 2703.900 2151.990 2704.160 2152.310 ;
        RECT 2702.060 2150.290 2702.320 2150.610 ;
        RECT 2702.520 2150.290 2702.780 2150.610 ;
        RECT 2698.900 2149.870 2699.500 2150.010 ;
        RECT 2698.900 2148.570 2699.040 2149.870 ;
        RECT 2698.380 2148.250 2698.640 2148.570 ;
        RECT 2698.840 2148.250 2699.100 2148.570 ;
        RECT 2699.760 2147.230 2700.020 2147.550 ;
        RECT 2699.820 2145.850 2699.960 2147.230 ;
        RECT 2699.760 2145.530 2700.020 2145.850 ;
        RECT 2698.840 2144.850 2699.100 2145.170 ;
        RECT 2698.380 2144.510 2698.640 2144.830 ;
        RECT 2697.920 2142.810 2698.180 2143.130 ;
        RECT 2694.690 2142.275 2694.970 2142.645 ;
        RECT 2694.760 2142.110 2694.900 2142.275 ;
        RECT 2694.700 2141.790 2694.960 2142.110 ;
        RECT 2694.700 2136.350 2694.960 2136.670 ;
        RECT 2694.760 2135.845 2694.900 2136.350 ;
        RECT 2694.690 2135.475 2694.970 2135.845 ;
        RECT 2698.440 2132.250 2698.580 2144.510 ;
        RECT 2698.900 2137.690 2699.040 2144.850 ;
        RECT 2698.840 2137.370 2699.100 2137.690 ;
        RECT 2702.580 2132.250 2702.720 2150.290 ;
        RECT 2698.380 2131.930 2698.640 2132.250 ;
        RECT 2702.520 2131.930 2702.780 2132.250 ;
        RECT 2694.700 2130.910 2694.960 2131.230 ;
        RECT 2698.380 2130.910 2698.640 2131.230 ;
        RECT 2694.760 2129.045 2694.900 2130.910 ;
        RECT 2694.690 2128.675 2694.970 2129.045 ;
        RECT 2698.440 2122.925 2698.580 2130.910 ;
        RECT 2698.370 2122.555 2698.650 2122.925 ;
        RECT 2677.300 2048.850 2677.560 2049.170 ;
        RECT 2677.360 2046.645 2677.500 2048.850 ;
        RECT 2677.290 2046.275 2677.570 2046.645 ;
        RECT 2695.150 2043.875 2695.430 2044.245 ;
        RECT 2695.220 2035.890 2695.360 2043.875 ;
        RECT 2695.610 2037.075 2695.890 2037.445 ;
        RECT 2695.680 2036.570 2695.820 2037.075 ;
        RECT 2695.620 2036.250 2695.880 2036.570 ;
        RECT 2698.840 2036.250 2699.100 2036.570 ;
        RECT 2702.520 2036.250 2702.780 2036.570 ;
        RECT 2695.160 2035.570 2695.420 2035.890 ;
        RECT 2677.300 2035.250 2677.560 2035.570 ;
        RECT 2677.360 2033.045 2677.500 2035.250 ;
        RECT 2698.380 2034.550 2698.640 2034.870 ;
        RECT 2677.290 2032.675 2677.570 2033.045 ;
        RECT 2694.700 2032.510 2694.960 2032.830 ;
        RECT 2698.440 2032.570 2698.580 2034.550 ;
        RECT 2694.760 2030.645 2694.900 2032.510 ;
        RECT 2697.520 2032.430 2698.580 2032.570 ;
        RECT 2694.690 2030.275 2694.970 2030.645 ;
        RECT 2694.700 2024.690 2694.960 2025.010 ;
        RECT 2694.760 2023.845 2694.900 2024.690 ;
        RECT 2694.690 2023.475 2694.970 2023.845 ;
        RECT 2697.000 2023.670 2697.260 2023.990 ;
        RECT 2697.520 2023.730 2697.660 2032.430 ;
        RECT 2697.920 2031.830 2698.180 2032.150 ;
        RECT 2697.980 2024.410 2698.120 2031.830 ;
        RECT 2697.980 2024.270 2698.580 2024.410 ;
        RECT 2677.290 2022.475 2677.570 2022.845 ;
        RECT 2677.360 2021.970 2677.500 2022.475 ;
        RECT 2677.300 2021.650 2677.560 2021.970 ;
        RECT 2694.690 2016.675 2694.970 2017.045 ;
        RECT 2694.760 2016.510 2694.900 2016.675 ;
        RECT 2694.700 2016.190 2694.960 2016.510 ;
        RECT 2677.290 2015.675 2677.570 2016.045 ;
        RECT 2677.360 2015.170 2677.500 2015.675 ;
        RECT 2677.300 2014.850 2677.560 2015.170 ;
        RECT 2697.060 2014.130 2697.200 2023.670 ;
        RECT 2697.520 2023.590 2698.120 2023.730 ;
        RECT 2697.460 2021.970 2697.720 2022.290 ;
        RECT 2697.520 2019.570 2697.660 2021.970 ;
        RECT 2697.980 2019.570 2698.120 2023.590 ;
        RECT 2698.440 2022.290 2698.580 2024.270 ;
        RECT 2698.380 2021.970 2698.640 2022.290 ;
        RECT 2697.460 2019.250 2697.720 2019.570 ;
        RECT 2697.920 2019.250 2698.180 2019.570 ;
        RECT 2697.460 2018.570 2697.720 2018.890 ;
        RECT 2697.000 2013.810 2697.260 2014.130 ;
        RECT 2694.700 2010.750 2694.960 2011.070 ;
        RECT 2694.760 2010.245 2694.900 2010.750 ;
        RECT 2694.690 2009.875 2694.970 2010.245 ;
        RECT 2681.890 2008.195 2682.170 2008.565 ;
        RECT 2681.430 2001.395 2681.710 2001.765 ;
        RECT 2677.290 1995.275 2677.570 1995.645 ;
        RECT 2677.360 1994.430 2677.500 1995.275 ;
        RECT 2677.300 1994.110 2677.560 1994.430 ;
        RECT 2680.510 1987.115 2680.790 1987.485 ;
        RECT 2677.290 1981.675 2677.570 1982.045 ;
        RECT 2677.360 1980.490 2677.500 1981.675 ;
        RECT 2677.300 1980.170 2677.560 1980.490 ;
        RECT 2677.300 1869.670 2677.560 1869.990 ;
        RECT 2677.360 1864.405 2677.500 1869.670 ;
        RECT 2677.290 1864.035 2677.570 1864.405 ;
        RECT 2677.300 1862.530 2677.560 1862.850 ;
        RECT 2677.360 1857.605 2677.500 1862.530 ;
        RECT 2677.290 1857.235 2677.570 1857.605 ;
        RECT 2677.300 1848.930 2677.560 1849.250 ;
        RECT 2677.360 1844.005 2677.500 1848.930 ;
        RECT 2677.290 1843.635 2677.570 1844.005 ;
        RECT 2677.290 1836.835 2677.570 1837.205 ;
        RECT 2677.360 1835.650 2677.500 1836.835 ;
        RECT 2677.300 1835.330 2677.560 1835.650 ;
        RECT 2677.290 1830.035 2677.570 1830.405 ;
        RECT 2677.360 1828.850 2677.500 1830.035 ;
        RECT 2677.300 1828.530 2677.560 1828.850 ;
        RECT 2677.290 1809.635 2677.570 1810.005 ;
        RECT 2677.360 1808.110 2677.500 1809.635 ;
        RECT 2677.300 1807.790 2677.560 1808.110 ;
        RECT 2625.320 1766.310 2625.580 1766.630 ;
        RECT 2618.420 1690.150 2618.680 1690.470 ;
        RECT 2625.380 1662.930 2625.520 1766.310 ;
        RECT 2677.300 1690.150 2677.560 1690.470 ;
        RECT 2677.360 1684.205 2677.500 1690.150 ;
        RECT 2677.290 1683.835 2677.570 1684.205 ;
        RECT 2625.320 1662.610 2625.580 1662.930 ;
        RECT 2677.300 1662.610 2677.560 1662.930 ;
        RECT 2677.360 1657.005 2677.500 1662.610 ;
        RECT 2677.290 1656.635 2677.570 1657.005 ;
        RECT 2677.300 1655.810 2677.560 1656.130 ;
        RECT 2677.360 1650.205 2677.500 1655.810 ;
        RECT 2677.290 1649.835 2677.570 1650.205 ;
        RECT 2680.050 1643.035 2680.330 1643.405 ;
        RECT 2677.290 1629.435 2677.570 1629.805 ;
        RECT 2677.360 1628.590 2677.500 1629.435 ;
        RECT 2618.420 1628.270 2618.680 1628.590 ;
        RECT 2677.300 1628.270 2677.560 1628.590 ;
        RECT 2611.520 1420.870 2611.780 1421.190 ;
        RECT 2618.480 1420.850 2618.620 1628.270 ;
        RECT 2680.120 1593.230 2680.260 1643.035 ;
        RECT 2680.060 1592.910 2680.320 1593.230 ;
        RECT 2677.300 1504.005 2677.560 1504.150 ;
        RECT 2677.290 1503.635 2677.570 1504.005 ;
        RECT 2677.300 1497.205 2677.560 1497.350 ;
        RECT 2677.290 1496.835 2677.570 1497.205 ;
        RECT 2677.300 1490.405 2677.560 1490.550 ;
        RECT 2677.290 1490.035 2677.570 1490.405 ;
        RECT 2677.290 1483.235 2677.570 1483.605 ;
        RECT 2677.360 1483.070 2677.500 1483.235 ;
        RECT 2677.760 1483.090 2678.020 1483.410 ;
        RECT 2677.300 1482.750 2677.560 1483.070 ;
        RECT 2677.820 1476.805 2677.960 1483.090 ;
        RECT 2677.300 1476.290 2677.560 1476.610 ;
        RECT 2677.750 1476.435 2678.030 1476.805 ;
        RECT 2677.360 1470.005 2677.500 1476.290 ;
        RECT 2677.290 1469.635 2677.570 1470.005 ;
        RECT 2677.760 1469.490 2678.020 1469.810 ;
        RECT 2677.820 1463.205 2677.960 1469.490 ;
        RECT 2677.750 1462.835 2678.030 1463.205 ;
        RECT 2677.300 1462.350 2677.560 1462.670 ;
        RECT 2677.360 1456.405 2677.500 1462.350 ;
        RECT 2677.290 1456.035 2677.570 1456.405 ;
        RECT 2677.290 1449.235 2677.570 1449.605 ;
        RECT 2677.300 1449.090 2677.560 1449.235 ;
        RECT 2677.290 1442.435 2677.570 1442.805 ;
        RECT 2677.360 1442.270 2677.500 1442.435 ;
        RECT 2677.300 1441.950 2677.560 1442.270 ;
        RECT 2680.580 1421.530 2680.720 1987.115 ;
        RECT 2680.970 1802.835 2681.250 1803.205 ;
        RECT 2680.520 1421.210 2680.780 1421.530 ;
        RECT 2618.420 1420.530 2618.680 1420.850 ;
        RECT 2681.040 1317.830 2681.180 1802.835 ;
        RECT 2681.500 1593.910 2681.640 2001.395 ;
        RECT 2681.960 1697.270 2682.100 2008.195 ;
        RECT 2697.520 2006.650 2697.660 2018.570 ;
        RECT 2698.900 2017.610 2699.040 2036.250 ;
        RECT 2701.600 2035.230 2701.860 2035.550 ;
        RECT 2697.980 2017.470 2699.040 2017.610 ;
        RECT 2697.980 2014.130 2698.120 2017.470 ;
        RECT 2697.920 2013.810 2698.180 2014.130 ;
        RECT 2698.840 2013.470 2699.100 2013.790 ;
        RECT 2698.380 2012.790 2698.640 2013.110 ;
        RECT 2697.920 2011.090 2698.180 2011.410 ;
        RECT 2697.460 2006.330 2697.720 2006.650 ;
        RECT 2694.700 2005.310 2694.960 2005.630 ;
        RECT 2694.760 2003.445 2694.900 2005.310 ;
        RECT 2694.690 2003.075 2694.970 2003.445 ;
        RECT 2694.700 1997.490 2694.960 1997.810 ;
        RECT 2694.760 1996.645 2694.900 1997.490 ;
        RECT 2694.690 1996.275 2694.970 1996.645 ;
        RECT 2694.700 1992.050 2694.960 1992.370 ;
        RECT 2694.760 1989.845 2694.900 1992.050 ;
        RECT 2697.460 1991.030 2697.720 1991.350 ;
        RECT 2694.690 1989.475 2694.970 1989.845 ;
        RECT 2697.520 1986.590 2697.660 1991.030 ;
        RECT 2697.980 1986.930 2698.120 2011.090 ;
        RECT 2698.440 1986.930 2698.580 2012.790 ;
        RECT 2698.900 1998.490 2699.040 2013.470 ;
        RECT 2701.660 2011.410 2701.800 2035.230 ;
        RECT 2702.060 2018.910 2702.320 2019.230 ;
        RECT 2702.120 2017.530 2702.260 2018.910 ;
        RECT 2702.580 2018.550 2702.720 2036.250 ;
        RECT 2721.840 2034.890 2722.100 2035.210 ;
        RECT 2721.900 2019.570 2722.040 2034.890 ;
        RECT 2731.500 2034.550 2731.760 2034.870 ;
        RECT 2721.840 2019.250 2722.100 2019.570 ;
        RECT 2702.980 2018.910 2703.240 2019.230 ;
        RECT 2702.520 2018.230 2702.780 2018.550 ;
        RECT 2702.060 2017.210 2702.320 2017.530 ;
        RECT 2702.060 2013.470 2702.320 2013.790 ;
        RECT 2702.120 2012.090 2702.260 2013.470 ;
        RECT 2702.580 2013.110 2702.720 2018.230 ;
        RECT 2703.040 2014.130 2703.180 2018.910 ;
        RECT 2703.900 2018.230 2704.160 2018.550 ;
        RECT 2702.980 2013.810 2703.240 2014.130 ;
        RECT 2702.520 2012.790 2702.780 2013.110 ;
        RECT 2702.060 2011.770 2702.320 2012.090 ;
        RECT 2701.600 2011.090 2701.860 2011.410 ;
        RECT 2701.600 2010.070 2701.860 2010.390 ;
        RECT 2701.660 2000.190 2701.800 2010.070 ;
        RECT 2701.600 1999.870 2701.860 2000.190 ;
        RECT 2702.060 1999.190 2702.320 1999.510 ;
        RECT 2702.120 1998.490 2702.260 1999.190 ;
        RECT 2698.840 1998.170 2699.100 1998.490 ;
        RECT 2702.060 1998.170 2702.320 1998.490 ;
        RECT 2702.520 1996.810 2702.780 1997.130 ;
        RECT 2702.580 1995.770 2702.720 1996.810 ;
        RECT 2702.520 1995.450 2702.780 1995.770 ;
        RECT 2697.920 1986.610 2698.180 1986.930 ;
        RECT 2698.380 1986.610 2698.640 1986.930 ;
        RECT 2697.460 1986.270 2697.720 1986.590 ;
        RECT 2694.700 1983.550 2694.960 1983.870 ;
        RECT 2697.980 1983.610 2698.120 1986.610 ;
        RECT 2694.760 1983.045 2694.900 1983.550 ;
        RECT 2697.520 1983.470 2698.120 1983.610 ;
        RECT 2694.690 1982.675 2694.970 1983.045 ;
        RECT 2697.520 1979.110 2697.660 1983.470 ;
        RECT 2697.920 1982.870 2698.180 1983.190 ;
        RECT 2697.980 1982.170 2698.120 1982.870 ;
        RECT 2697.920 1981.850 2698.180 1982.170 ;
        RECT 2698.440 1981.830 2698.580 1986.610 ;
        RECT 2702.060 1986.270 2702.320 1986.590 ;
        RECT 2703.040 1986.330 2703.180 2013.810 ;
        RECT 2703.960 2010.730 2704.100 2018.230 ;
        RECT 2706.200 2012.790 2706.460 2013.110 ;
        RECT 2706.260 2012.090 2706.400 2012.790 ;
        RECT 2706.200 2011.770 2706.460 2012.090 ;
        RECT 2703.900 2010.410 2704.160 2010.730 ;
        RECT 2731.560 2000.190 2731.700 2034.550 ;
        RECT 2703.900 1999.870 2704.160 2000.190 ;
        RECT 2731.500 1999.870 2731.760 2000.190 ;
        RECT 2703.960 1998.490 2704.100 1999.870 ;
        RECT 2703.900 1998.170 2704.160 1998.490 ;
        RECT 2704.820 1997.150 2705.080 1997.470 ;
        RECT 2704.880 1994.490 2705.020 1997.150 ;
        RECT 2702.120 1982.170 2702.260 1986.270 ;
        RECT 2702.580 1986.190 2703.180 1986.330 ;
        RECT 2703.960 1994.350 2705.020 1994.490 ;
        RECT 2702.060 1981.850 2702.320 1982.170 ;
        RECT 2698.380 1981.570 2698.640 1981.830 ;
        RECT 2698.380 1981.510 2699.040 1981.570 ;
        RECT 2698.440 1981.430 2699.040 1981.510 ;
        RECT 2702.580 1981.490 2702.720 1986.190 ;
        RECT 2702.980 1985.590 2703.240 1985.910 ;
        RECT 2703.040 1982.170 2703.180 1985.590 ;
        RECT 2702.980 1981.850 2703.240 1982.170 ;
        RECT 2703.440 1981.850 2703.700 1982.170 ;
        RECT 2698.380 1980.830 2698.640 1981.150 ;
        RECT 2697.460 1978.790 2697.720 1979.110 ;
        RECT 2694.690 1975.875 2694.970 1976.245 ;
        RECT 2694.700 1975.730 2694.960 1975.875 ;
        RECT 2697.000 1972.330 2697.260 1972.650 ;
        RECT 2697.060 1969.590 2697.200 1972.330 ;
        RECT 2697.520 1970.610 2697.660 1978.790 ;
        RECT 2697.460 1970.290 2697.720 1970.610 ;
        RECT 2697.920 1970.290 2698.180 1970.610 ;
        RECT 2694.690 1969.075 2694.970 1969.445 ;
        RECT 2697.000 1969.270 2697.260 1969.590 ;
        RECT 2694.760 1967.550 2694.900 1969.075 ;
        RECT 2694.700 1967.230 2694.960 1967.550 ;
        RECT 2697.060 1964.830 2697.200 1969.270 ;
        RECT 2697.520 1967.550 2697.660 1970.290 ;
        RECT 2697.460 1967.230 2697.720 1967.550 ;
        RECT 2697.000 1964.510 2697.260 1964.830 ;
        RECT 2697.980 1963.130 2698.120 1970.290 ;
        RECT 2698.440 1968.570 2698.580 1980.830 ;
        RECT 2698.900 1979.450 2699.040 1981.430 ;
        RECT 2702.520 1981.170 2702.780 1981.490 ;
        RECT 2702.580 1980.890 2702.720 1981.170 ;
        RECT 2701.660 1980.750 2702.720 1980.890 ;
        RECT 2698.840 1979.130 2699.100 1979.450 ;
        RECT 2698.840 1977.430 2699.100 1977.750 ;
        RECT 2698.900 1976.730 2699.040 1977.430 ;
        RECT 2698.840 1976.410 2699.100 1976.730 ;
        RECT 2701.660 1973.330 2701.800 1980.750 ;
        RECT 2702.520 1980.150 2702.780 1980.470 ;
        RECT 2702.580 1979.450 2702.720 1980.150 ;
        RECT 2702.520 1979.130 2702.780 1979.450 ;
        RECT 2702.060 1978.790 2702.320 1979.110 ;
        RECT 2701.600 1973.010 2701.860 1973.330 ;
        RECT 2699.760 1972.670 2700.020 1972.990 ;
        RECT 2698.840 1971.990 2699.100 1972.310 ;
        RECT 2699.300 1971.990 2699.560 1972.310 ;
        RECT 2698.900 1971.290 2699.040 1971.990 ;
        RECT 2698.840 1970.970 2699.100 1971.290 ;
        RECT 2699.360 1970.010 2699.500 1971.990 ;
        RECT 2699.820 1970.950 2699.960 1972.670 ;
        RECT 2702.120 1972.650 2702.260 1978.790 ;
        RECT 2703.500 1972.990 2703.640 1981.850 ;
        RECT 2703.440 1972.670 2703.700 1972.990 ;
        RECT 2702.060 1972.330 2702.320 1972.650 ;
        RECT 2699.760 1970.630 2700.020 1970.950 ;
        RECT 2702.120 1970.610 2702.260 1972.330 ;
        RECT 2703.960 1972.310 2704.100 1994.350 ;
        RECT 2703.900 1971.990 2704.160 1972.310 ;
        RECT 2702.060 1970.290 2702.320 1970.610 ;
        RECT 2702.520 1970.290 2702.780 1970.610 ;
        RECT 2698.900 1969.870 2699.500 1970.010 ;
        RECT 2698.900 1968.570 2699.040 1969.870 ;
        RECT 2698.380 1968.250 2698.640 1968.570 ;
        RECT 2698.840 1968.250 2699.100 1968.570 ;
        RECT 2699.760 1967.230 2700.020 1967.550 ;
        RECT 2699.820 1965.850 2699.960 1967.230 ;
        RECT 2699.760 1965.530 2700.020 1965.850 ;
        RECT 2698.840 1964.850 2699.100 1965.170 ;
        RECT 2698.380 1964.510 2698.640 1964.830 ;
        RECT 2697.920 1962.810 2698.180 1963.130 ;
        RECT 2694.690 1962.275 2694.970 1962.645 ;
        RECT 2694.760 1962.110 2694.900 1962.275 ;
        RECT 2694.700 1961.790 2694.960 1962.110 ;
        RECT 2694.700 1956.350 2694.960 1956.670 ;
        RECT 2694.760 1955.845 2694.900 1956.350 ;
        RECT 2694.690 1955.475 2694.970 1955.845 ;
        RECT 2698.440 1952.250 2698.580 1964.510 ;
        RECT 2698.900 1957.690 2699.040 1964.850 ;
        RECT 2698.840 1957.370 2699.100 1957.690 ;
        RECT 2702.580 1952.250 2702.720 1970.290 ;
        RECT 2698.380 1951.930 2698.640 1952.250 ;
        RECT 2702.520 1951.930 2702.780 1952.250 ;
        RECT 2694.700 1950.910 2694.960 1951.230 ;
        RECT 2698.380 1950.910 2698.640 1951.230 ;
        RECT 2694.760 1949.045 2694.900 1950.910 ;
        RECT 2694.690 1948.675 2694.970 1949.045 ;
        RECT 2698.440 1942.925 2698.580 1950.910 ;
        RECT 2698.370 1942.555 2698.650 1942.925 ;
        RECT 2695.150 1863.875 2695.430 1864.245 ;
        RECT 2695.220 1855.890 2695.360 1863.875 ;
        RECT 2695.610 1857.075 2695.890 1857.445 ;
        RECT 2695.680 1856.570 2695.820 1857.075 ;
        RECT 2695.620 1856.250 2695.880 1856.570 ;
        RECT 2698.840 1856.250 2699.100 1856.570 ;
        RECT 2702.520 1856.250 2702.780 1856.570 ;
        RECT 2695.160 1855.570 2695.420 1855.890 ;
        RECT 2698.380 1854.550 2698.640 1854.870 ;
        RECT 2694.700 1852.510 2694.960 1852.830 ;
        RECT 2698.440 1852.570 2698.580 1854.550 ;
        RECT 2694.760 1850.645 2694.900 1852.510 ;
        RECT 2697.520 1852.430 2698.580 1852.570 ;
        RECT 2694.690 1850.275 2694.970 1850.645 ;
        RECT 2694.700 1844.690 2694.960 1845.010 ;
        RECT 2694.760 1843.845 2694.900 1844.690 ;
        RECT 2694.690 1843.475 2694.970 1843.845 ;
        RECT 2697.000 1843.670 2697.260 1843.990 ;
        RECT 2697.520 1843.730 2697.660 1852.430 ;
        RECT 2697.920 1851.830 2698.180 1852.150 ;
        RECT 2697.980 1844.410 2698.120 1851.830 ;
        RECT 2697.980 1844.270 2698.580 1844.410 ;
        RECT 2694.690 1836.675 2694.970 1837.045 ;
        RECT 2694.760 1836.510 2694.900 1836.675 ;
        RECT 2694.700 1836.190 2694.960 1836.510 ;
        RECT 2697.060 1834.130 2697.200 1843.670 ;
        RECT 2697.520 1843.590 2698.120 1843.730 ;
        RECT 2697.460 1841.970 2697.720 1842.290 ;
        RECT 2697.520 1839.570 2697.660 1841.970 ;
        RECT 2697.980 1839.570 2698.120 1843.590 ;
        RECT 2698.440 1842.290 2698.580 1844.270 ;
        RECT 2698.380 1841.970 2698.640 1842.290 ;
        RECT 2697.460 1839.250 2697.720 1839.570 ;
        RECT 2697.920 1839.250 2698.180 1839.570 ;
        RECT 2697.460 1838.570 2697.720 1838.890 ;
        RECT 2697.000 1833.810 2697.260 1834.130 ;
        RECT 2694.700 1830.750 2694.960 1831.070 ;
        RECT 2694.760 1830.245 2694.900 1830.750 ;
        RECT 2694.690 1829.875 2694.970 1830.245 ;
        RECT 2697.520 1826.650 2697.660 1838.570 ;
        RECT 2698.900 1837.610 2699.040 1856.250 ;
        RECT 2701.600 1855.230 2701.860 1855.550 ;
        RECT 2697.980 1837.470 2699.040 1837.610 ;
        RECT 2697.980 1834.130 2698.120 1837.470 ;
        RECT 2697.920 1833.810 2698.180 1834.130 ;
        RECT 2698.840 1833.470 2699.100 1833.790 ;
        RECT 2698.380 1832.790 2698.640 1833.110 ;
        RECT 2697.920 1831.090 2698.180 1831.410 ;
        RECT 2697.460 1826.330 2697.720 1826.650 ;
        RECT 2694.700 1825.310 2694.960 1825.630 ;
        RECT 2682.810 1823.235 2683.090 1823.605 ;
        RECT 2694.760 1823.445 2694.900 1825.310 ;
        RECT 2682.350 1816.435 2682.630 1816.805 ;
        RECT 2681.900 1696.950 2682.160 1697.270 ;
        RECT 2681.890 1622.635 2682.170 1623.005 ;
        RECT 2681.440 1593.590 2681.700 1593.910 ;
        RECT 2680.980 1317.510 2681.240 1317.830 ;
        RECT 2681.960 1317.490 2682.100 1622.635 ;
        RECT 2682.420 1518.090 2682.560 1816.435 ;
        RECT 2682.880 1593.570 2683.020 1823.235 ;
        RECT 2694.690 1823.075 2694.970 1823.445 ;
        RECT 2694.700 1817.490 2694.960 1817.810 ;
        RECT 2694.760 1816.645 2694.900 1817.490 ;
        RECT 2694.690 1816.275 2694.970 1816.645 ;
        RECT 2694.700 1812.050 2694.960 1812.370 ;
        RECT 2694.760 1809.845 2694.900 1812.050 ;
        RECT 2697.460 1811.030 2697.720 1811.350 ;
        RECT 2694.690 1809.475 2694.970 1809.845 ;
        RECT 2697.520 1806.590 2697.660 1811.030 ;
        RECT 2697.980 1806.930 2698.120 1831.090 ;
        RECT 2698.440 1806.930 2698.580 1832.790 ;
        RECT 2698.900 1818.490 2699.040 1833.470 ;
        RECT 2701.660 1831.410 2701.800 1855.230 ;
        RECT 2702.060 1838.910 2702.320 1839.230 ;
        RECT 2702.120 1837.530 2702.260 1838.910 ;
        RECT 2702.580 1838.550 2702.720 1856.250 ;
        RECT 2721.840 1854.890 2722.100 1855.210 ;
        RECT 2721.900 1839.570 2722.040 1854.890 ;
        RECT 2731.500 1854.550 2731.760 1854.870 ;
        RECT 2721.840 1839.250 2722.100 1839.570 ;
        RECT 2702.980 1838.910 2703.240 1839.230 ;
        RECT 2702.520 1838.230 2702.780 1838.550 ;
        RECT 2702.060 1837.210 2702.320 1837.530 ;
        RECT 2702.060 1833.470 2702.320 1833.790 ;
        RECT 2702.120 1832.090 2702.260 1833.470 ;
        RECT 2702.580 1833.110 2702.720 1838.230 ;
        RECT 2703.040 1834.130 2703.180 1838.910 ;
        RECT 2703.900 1838.230 2704.160 1838.550 ;
        RECT 2702.980 1833.810 2703.240 1834.130 ;
        RECT 2702.520 1832.790 2702.780 1833.110 ;
        RECT 2702.060 1831.770 2702.320 1832.090 ;
        RECT 2701.600 1831.090 2701.860 1831.410 ;
        RECT 2701.600 1830.070 2701.860 1830.390 ;
        RECT 2701.660 1820.190 2701.800 1830.070 ;
        RECT 2701.600 1819.870 2701.860 1820.190 ;
        RECT 2702.060 1819.190 2702.320 1819.510 ;
        RECT 2702.120 1818.490 2702.260 1819.190 ;
        RECT 2698.840 1818.170 2699.100 1818.490 ;
        RECT 2702.060 1818.170 2702.320 1818.490 ;
        RECT 2702.520 1816.810 2702.780 1817.130 ;
        RECT 2702.580 1815.770 2702.720 1816.810 ;
        RECT 2702.520 1815.450 2702.780 1815.770 ;
        RECT 2697.920 1806.610 2698.180 1806.930 ;
        RECT 2698.380 1806.610 2698.640 1806.930 ;
        RECT 2697.460 1806.270 2697.720 1806.590 ;
        RECT 2694.700 1803.550 2694.960 1803.870 ;
        RECT 2697.980 1803.610 2698.120 1806.610 ;
        RECT 2694.760 1803.045 2694.900 1803.550 ;
        RECT 2697.520 1803.470 2698.120 1803.610 ;
        RECT 2694.690 1802.675 2694.970 1803.045 ;
        RECT 2697.520 1799.110 2697.660 1803.470 ;
        RECT 2697.920 1802.870 2698.180 1803.190 ;
        RECT 2697.980 1802.170 2698.120 1802.870 ;
        RECT 2697.920 1801.850 2698.180 1802.170 ;
        RECT 2698.440 1801.830 2698.580 1806.610 ;
        RECT 2702.060 1806.270 2702.320 1806.590 ;
        RECT 2703.040 1806.330 2703.180 1833.810 ;
        RECT 2703.960 1830.730 2704.100 1838.230 ;
        RECT 2706.200 1832.790 2706.460 1833.110 ;
        RECT 2706.260 1832.090 2706.400 1832.790 ;
        RECT 2706.200 1831.770 2706.460 1832.090 ;
        RECT 2703.900 1830.410 2704.160 1830.730 ;
        RECT 2731.560 1820.190 2731.700 1854.550 ;
        RECT 2703.900 1819.870 2704.160 1820.190 ;
        RECT 2731.500 1819.870 2731.760 1820.190 ;
        RECT 2703.960 1818.490 2704.100 1819.870 ;
        RECT 2703.900 1818.170 2704.160 1818.490 ;
        RECT 2704.820 1817.150 2705.080 1817.470 ;
        RECT 2704.880 1814.490 2705.020 1817.150 ;
        RECT 2702.120 1802.170 2702.260 1806.270 ;
        RECT 2702.580 1806.190 2703.180 1806.330 ;
        RECT 2703.960 1814.350 2705.020 1814.490 ;
        RECT 2702.060 1801.850 2702.320 1802.170 ;
        RECT 2698.380 1801.570 2698.640 1801.830 ;
        RECT 2698.380 1801.510 2699.040 1801.570 ;
        RECT 2698.440 1801.430 2699.040 1801.510 ;
        RECT 2702.580 1801.490 2702.720 1806.190 ;
        RECT 2702.980 1805.590 2703.240 1805.910 ;
        RECT 2703.040 1802.170 2703.180 1805.590 ;
        RECT 2702.980 1801.850 2703.240 1802.170 ;
        RECT 2703.440 1801.850 2703.700 1802.170 ;
        RECT 2698.380 1800.830 2698.640 1801.150 ;
        RECT 2697.460 1798.790 2697.720 1799.110 ;
        RECT 2694.690 1795.875 2694.970 1796.245 ;
        RECT 2694.700 1795.730 2694.960 1795.875 ;
        RECT 2697.000 1792.330 2697.260 1792.650 ;
        RECT 2697.060 1789.590 2697.200 1792.330 ;
        RECT 2697.520 1790.610 2697.660 1798.790 ;
        RECT 2697.460 1790.290 2697.720 1790.610 ;
        RECT 2697.920 1790.290 2698.180 1790.610 ;
        RECT 2694.690 1789.075 2694.970 1789.445 ;
        RECT 2697.000 1789.270 2697.260 1789.590 ;
        RECT 2694.760 1787.550 2694.900 1789.075 ;
        RECT 2694.700 1787.230 2694.960 1787.550 ;
        RECT 2697.060 1784.830 2697.200 1789.270 ;
        RECT 2697.520 1787.550 2697.660 1790.290 ;
        RECT 2697.460 1787.230 2697.720 1787.550 ;
        RECT 2697.000 1784.510 2697.260 1784.830 ;
        RECT 2697.980 1783.130 2698.120 1790.290 ;
        RECT 2698.440 1788.570 2698.580 1800.830 ;
        RECT 2698.900 1799.450 2699.040 1801.430 ;
        RECT 2702.520 1801.170 2702.780 1801.490 ;
        RECT 2702.580 1800.890 2702.720 1801.170 ;
        RECT 2701.660 1800.750 2702.720 1800.890 ;
        RECT 2698.840 1799.130 2699.100 1799.450 ;
        RECT 2698.840 1797.430 2699.100 1797.750 ;
        RECT 2698.900 1796.730 2699.040 1797.430 ;
        RECT 2698.840 1796.410 2699.100 1796.730 ;
        RECT 2701.660 1793.330 2701.800 1800.750 ;
        RECT 2702.520 1800.150 2702.780 1800.470 ;
        RECT 2702.580 1799.450 2702.720 1800.150 ;
        RECT 2702.520 1799.130 2702.780 1799.450 ;
        RECT 2702.060 1798.790 2702.320 1799.110 ;
        RECT 2701.600 1793.010 2701.860 1793.330 ;
        RECT 2699.760 1792.670 2700.020 1792.990 ;
        RECT 2698.840 1791.990 2699.100 1792.310 ;
        RECT 2699.300 1791.990 2699.560 1792.310 ;
        RECT 2698.900 1791.290 2699.040 1791.990 ;
        RECT 2698.840 1790.970 2699.100 1791.290 ;
        RECT 2699.360 1790.010 2699.500 1791.990 ;
        RECT 2699.820 1790.950 2699.960 1792.670 ;
        RECT 2702.120 1792.650 2702.260 1798.790 ;
        RECT 2703.500 1792.990 2703.640 1801.850 ;
        RECT 2703.440 1792.670 2703.700 1792.990 ;
        RECT 2702.060 1792.330 2702.320 1792.650 ;
        RECT 2699.760 1790.630 2700.020 1790.950 ;
        RECT 2702.120 1790.610 2702.260 1792.330 ;
        RECT 2703.960 1792.310 2704.100 1814.350 ;
        RECT 2703.900 1791.990 2704.160 1792.310 ;
        RECT 2702.060 1790.290 2702.320 1790.610 ;
        RECT 2702.520 1790.290 2702.780 1790.610 ;
        RECT 2698.900 1789.870 2699.500 1790.010 ;
        RECT 2698.900 1788.570 2699.040 1789.870 ;
        RECT 2698.380 1788.250 2698.640 1788.570 ;
        RECT 2698.840 1788.250 2699.100 1788.570 ;
        RECT 2699.760 1787.230 2700.020 1787.550 ;
        RECT 2699.820 1785.850 2699.960 1787.230 ;
        RECT 2699.760 1785.530 2700.020 1785.850 ;
        RECT 2698.840 1784.850 2699.100 1785.170 ;
        RECT 2698.380 1784.510 2698.640 1784.830 ;
        RECT 2697.920 1782.810 2698.180 1783.130 ;
        RECT 2694.690 1782.275 2694.970 1782.645 ;
        RECT 2694.760 1782.110 2694.900 1782.275 ;
        RECT 2694.700 1781.790 2694.960 1782.110 ;
        RECT 2694.700 1776.350 2694.960 1776.670 ;
        RECT 2694.760 1775.845 2694.900 1776.350 ;
        RECT 2694.690 1775.475 2694.970 1775.845 ;
        RECT 2698.440 1772.250 2698.580 1784.510 ;
        RECT 2698.900 1777.690 2699.040 1784.850 ;
        RECT 2698.840 1777.370 2699.100 1777.690 ;
        RECT 2702.580 1772.250 2702.720 1790.290 ;
        RECT 2698.380 1771.930 2698.640 1772.250 ;
        RECT 2702.520 1771.930 2702.780 1772.250 ;
        RECT 2694.700 1770.910 2694.960 1771.230 ;
        RECT 2698.380 1770.910 2698.640 1771.230 ;
        RECT 2694.760 1769.045 2694.900 1770.910 ;
        RECT 2694.690 1768.675 2694.970 1769.045 ;
        RECT 2698.440 1762.925 2698.580 1770.910 ;
        RECT 2698.370 1762.555 2698.650 1762.925 ;
        RECT 2695.150 1683.875 2695.430 1684.245 ;
        RECT 2695.220 1675.890 2695.360 1683.875 ;
        RECT 2695.610 1677.075 2695.890 1677.445 ;
        RECT 2695.680 1676.570 2695.820 1677.075 ;
        RECT 2695.620 1676.250 2695.880 1676.570 ;
        RECT 2698.840 1676.250 2699.100 1676.570 ;
        RECT 2702.520 1676.250 2702.780 1676.570 ;
        RECT 2695.160 1675.570 2695.420 1675.890 ;
        RECT 2698.380 1674.550 2698.640 1674.870 ;
        RECT 2694.700 1672.510 2694.960 1672.830 ;
        RECT 2698.440 1672.570 2698.580 1674.550 ;
        RECT 2694.760 1670.645 2694.900 1672.510 ;
        RECT 2697.520 1672.430 2698.580 1672.570 ;
        RECT 2694.690 1670.275 2694.970 1670.645 ;
        RECT 2694.700 1664.690 2694.960 1665.010 ;
        RECT 2694.760 1663.845 2694.900 1664.690 ;
        RECT 2694.690 1663.475 2694.970 1663.845 ;
        RECT 2697.000 1663.670 2697.260 1663.990 ;
        RECT 2697.520 1663.730 2697.660 1672.430 ;
        RECT 2697.920 1671.830 2698.180 1672.150 ;
        RECT 2697.980 1664.410 2698.120 1671.830 ;
        RECT 2697.980 1664.270 2698.580 1664.410 ;
        RECT 2694.690 1656.675 2694.970 1657.045 ;
        RECT 2694.760 1656.510 2694.900 1656.675 ;
        RECT 2694.700 1656.190 2694.960 1656.510 ;
        RECT 2697.060 1654.130 2697.200 1663.670 ;
        RECT 2697.520 1663.590 2698.120 1663.730 ;
        RECT 2697.460 1661.970 2697.720 1662.290 ;
        RECT 2697.520 1659.570 2697.660 1661.970 ;
        RECT 2697.980 1659.570 2698.120 1663.590 ;
        RECT 2698.440 1662.290 2698.580 1664.270 ;
        RECT 2698.380 1661.970 2698.640 1662.290 ;
        RECT 2697.460 1659.250 2697.720 1659.570 ;
        RECT 2697.920 1659.250 2698.180 1659.570 ;
        RECT 2697.460 1658.570 2697.720 1658.890 ;
        RECT 2697.000 1653.810 2697.260 1654.130 ;
        RECT 2694.700 1650.750 2694.960 1651.070 ;
        RECT 2694.760 1650.245 2694.900 1650.750 ;
        RECT 2694.690 1649.875 2694.970 1650.245 ;
        RECT 2697.520 1646.650 2697.660 1658.570 ;
        RECT 2698.900 1657.610 2699.040 1676.250 ;
        RECT 2701.600 1675.230 2701.860 1675.550 ;
        RECT 2697.980 1657.470 2699.040 1657.610 ;
        RECT 2697.980 1654.130 2698.120 1657.470 ;
        RECT 2697.920 1653.810 2698.180 1654.130 ;
        RECT 2698.840 1653.470 2699.100 1653.790 ;
        RECT 2698.380 1652.790 2698.640 1653.110 ;
        RECT 2697.920 1651.090 2698.180 1651.410 ;
        RECT 2697.460 1646.330 2697.720 1646.650 ;
        RECT 2694.700 1645.310 2694.960 1645.630 ;
        RECT 2694.760 1643.445 2694.900 1645.310 ;
        RECT 2694.690 1643.075 2694.970 1643.445 ;
        RECT 2694.700 1637.490 2694.960 1637.810 ;
        RECT 2694.760 1636.645 2694.900 1637.490 ;
        RECT 2683.270 1636.235 2683.550 1636.605 ;
        RECT 2694.690 1636.275 2694.970 1636.645 ;
        RECT 2682.820 1593.250 2683.080 1593.570 ;
        RECT 2682.360 1517.770 2682.620 1518.090 ;
        RECT 2683.340 1517.750 2683.480 1636.235 ;
        RECT 2694.700 1632.050 2694.960 1632.370 ;
        RECT 2694.760 1629.845 2694.900 1632.050 ;
        RECT 2697.460 1631.030 2697.720 1631.350 ;
        RECT 2694.690 1629.475 2694.970 1629.845 ;
        RECT 2697.520 1626.590 2697.660 1631.030 ;
        RECT 2697.980 1626.930 2698.120 1651.090 ;
        RECT 2698.440 1626.930 2698.580 1652.790 ;
        RECT 2698.900 1638.490 2699.040 1653.470 ;
        RECT 2701.660 1651.410 2701.800 1675.230 ;
        RECT 2702.060 1658.910 2702.320 1659.230 ;
        RECT 2702.120 1657.530 2702.260 1658.910 ;
        RECT 2702.580 1658.550 2702.720 1676.250 ;
        RECT 2721.840 1674.890 2722.100 1675.210 ;
        RECT 2721.900 1659.570 2722.040 1674.890 ;
        RECT 2731.500 1674.550 2731.760 1674.870 ;
        RECT 2721.840 1659.250 2722.100 1659.570 ;
        RECT 2702.980 1658.910 2703.240 1659.230 ;
        RECT 2702.520 1658.230 2702.780 1658.550 ;
        RECT 2702.060 1657.210 2702.320 1657.530 ;
        RECT 2702.060 1653.470 2702.320 1653.790 ;
        RECT 2702.120 1652.090 2702.260 1653.470 ;
        RECT 2702.580 1653.110 2702.720 1658.230 ;
        RECT 2703.040 1654.130 2703.180 1658.910 ;
        RECT 2703.900 1658.230 2704.160 1658.550 ;
        RECT 2702.980 1653.810 2703.240 1654.130 ;
        RECT 2702.520 1652.790 2702.780 1653.110 ;
        RECT 2702.060 1651.770 2702.320 1652.090 ;
        RECT 2701.600 1651.090 2701.860 1651.410 ;
        RECT 2701.600 1650.070 2701.860 1650.390 ;
        RECT 2701.660 1640.190 2701.800 1650.070 ;
        RECT 2701.600 1639.870 2701.860 1640.190 ;
        RECT 2702.060 1639.190 2702.320 1639.510 ;
        RECT 2702.120 1638.490 2702.260 1639.190 ;
        RECT 2698.840 1638.170 2699.100 1638.490 ;
        RECT 2702.060 1638.170 2702.320 1638.490 ;
        RECT 2702.520 1636.810 2702.780 1637.130 ;
        RECT 2702.580 1635.770 2702.720 1636.810 ;
        RECT 2702.520 1635.450 2702.780 1635.770 ;
        RECT 2697.920 1626.610 2698.180 1626.930 ;
        RECT 2698.380 1626.610 2698.640 1626.930 ;
        RECT 2697.460 1626.270 2697.720 1626.590 ;
        RECT 2694.700 1623.550 2694.960 1623.870 ;
        RECT 2697.980 1623.610 2698.120 1626.610 ;
        RECT 2694.760 1623.045 2694.900 1623.550 ;
        RECT 2697.520 1623.470 2698.120 1623.610 ;
        RECT 2694.690 1622.675 2694.970 1623.045 ;
        RECT 2697.520 1619.110 2697.660 1623.470 ;
        RECT 2697.920 1622.870 2698.180 1623.190 ;
        RECT 2697.980 1622.170 2698.120 1622.870 ;
        RECT 2697.920 1621.850 2698.180 1622.170 ;
        RECT 2698.440 1621.830 2698.580 1626.610 ;
        RECT 2702.060 1626.270 2702.320 1626.590 ;
        RECT 2703.040 1626.330 2703.180 1653.810 ;
        RECT 2703.960 1650.730 2704.100 1658.230 ;
        RECT 2706.200 1652.790 2706.460 1653.110 ;
        RECT 2706.260 1652.090 2706.400 1652.790 ;
        RECT 2706.200 1651.770 2706.460 1652.090 ;
        RECT 2703.900 1650.410 2704.160 1650.730 ;
        RECT 2731.560 1640.190 2731.700 1674.550 ;
        RECT 2703.900 1639.870 2704.160 1640.190 ;
        RECT 2731.500 1639.870 2731.760 1640.190 ;
        RECT 2703.960 1638.490 2704.100 1639.870 ;
        RECT 2703.900 1638.170 2704.160 1638.490 ;
        RECT 2704.820 1637.150 2705.080 1637.470 ;
        RECT 2704.880 1634.490 2705.020 1637.150 ;
        RECT 2702.120 1622.170 2702.260 1626.270 ;
        RECT 2702.580 1626.190 2703.180 1626.330 ;
        RECT 2703.960 1634.350 2705.020 1634.490 ;
        RECT 2702.060 1621.850 2702.320 1622.170 ;
        RECT 2698.380 1621.570 2698.640 1621.830 ;
        RECT 2698.380 1621.510 2699.040 1621.570 ;
        RECT 2698.440 1621.430 2699.040 1621.510 ;
        RECT 2702.580 1621.490 2702.720 1626.190 ;
        RECT 2702.980 1625.590 2703.240 1625.910 ;
        RECT 2703.040 1622.170 2703.180 1625.590 ;
        RECT 2702.980 1621.850 2703.240 1622.170 ;
        RECT 2703.440 1621.850 2703.700 1622.170 ;
        RECT 2698.380 1620.830 2698.640 1621.150 ;
        RECT 2697.460 1618.790 2697.720 1619.110 ;
        RECT 2694.690 1615.875 2694.970 1616.245 ;
        RECT 2694.700 1615.730 2694.960 1615.875 ;
        RECT 2697.000 1612.330 2697.260 1612.650 ;
        RECT 2697.060 1609.590 2697.200 1612.330 ;
        RECT 2697.520 1610.610 2697.660 1618.790 ;
        RECT 2697.460 1610.290 2697.720 1610.610 ;
        RECT 2697.920 1610.290 2698.180 1610.610 ;
        RECT 2694.690 1609.075 2694.970 1609.445 ;
        RECT 2697.000 1609.270 2697.260 1609.590 ;
        RECT 2694.760 1607.550 2694.900 1609.075 ;
        RECT 2694.700 1607.230 2694.960 1607.550 ;
        RECT 2697.060 1604.830 2697.200 1609.270 ;
        RECT 2697.520 1607.550 2697.660 1610.290 ;
        RECT 2697.460 1607.230 2697.720 1607.550 ;
        RECT 2697.000 1604.510 2697.260 1604.830 ;
        RECT 2697.980 1603.130 2698.120 1610.290 ;
        RECT 2698.440 1608.570 2698.580 1620.830 ;
        RECT 2698.900 1619.450 2699.040 1621.430 ;
        RECT 2702.520 1621.170 2702.780 1621.490 ;
        RECT 2702.580 1620.890 2702.720 1621.170 ;
        RECT 2701.660 1620.750 2702.720 1620.890 ;
        RECT 2698.840 1619.130 2699.100 1619.450 ;
        RECT 2698.840 1617.430 2699.100 1617.750 ;
        RECT 2698.900 1616.730 2699.040 1617.430 ;
        RECT 2698.840 1616.410 2699.100 1616.730 ;
        RECT 2701.660 1613.330 2701.800 1620.750 ;
        RECT 2702.520 1620.150 2702.780 1620.470 ;
        RECT 2702.580 1619.450 2702.720 1620.150 ;
        RECT 2702.520 1619.130 2702.780 1619.450 ;
        RECT 2702.060 1618.790 2702.320 1619.110 ;
        RECT 2701.600 1613.010 2701.860 1613.330 ;
        RECT 2699.760 1612.670 2700.020 1612.990 ;
        RECT 2698.840 1611.990 2699.100 1612.310 ;
        RECT 2699.300 1611.990 2699.560 1612.310 ;
        RECT 2698.900 1611.290 2699.040 1611.990 ;
        RECT 2698.840 1610.970 2699.100 1611.290 ;
        RECT 2699.360 1610.010 2699.500 1611.990 ;
        RECT 2699.820 1610.950 2699.960 1612.670 ;
        RECT 2702.120 1612.650 2702.260 1618.790 ;
        RECT 2703.500 1612.990 2703.640 1621.850 ;
        RECT 2703.440 1612.670 2703.700 1612.990 ;
        RECT 2702.060 1612.330 2702.320 1612.650 ;
        RECT 2699.760 1610.630 2700.020 1610.950 ;
        RECT 2702.120 1610.610 2702.260 1612.330 ;
        RECT 2703.960 1612.310 2704.100 1634.350 ;
        RECT 2703.900 1611.990 2704.160 1612.310 ;
        RECT 2702.060 1610.290 2702.320 1610.610 ;
        RECT 2702.520 1610.290 2702.780 1610.610 ;
        RECT 2698.900 1609.870 2699.500 1610.010 ;
        RECT 2698.900 1608.570 2699.040 1609.870 ;
        RECT 2698.380 1608.250 2698.640 1608.570 ;
        RECT 2698.840 1608.250 2699.100 1608.570 ;
        RECT 2699.760 1607.230 2700.020 1607.550 ;
        RECT 2699.820 1605.850 2699.960 1607.230 ;
        RECT 2699.760 1605.530 2700.020 1605.850 ;
        RECT 2698.840 1604.850 2699.100 1605.170 ;
        RECT 2698.380 1604.510 2698.640 1604.830 ;
        RECT 2697.920 1602.810 2698.180 1603.130 ;
        RECT 2694.690 1602.275 2694.970 1602.645 ;
        RECT 2694.760 1602.110 2694.900 1602.275 ;
        RECT 2694.700 1601.790 2694.960 1602.110 ;
        RECT 2694.700 1596.350 2694.960 1596.670 ;
        RECT 2694.760 1595.845 2694.900 1596.350 ;
        RECT 2694.690 1595.475 2694.970 1595.845 ;
        RECT 2698.440 1592.250 2698.580 1604.510 ;
        RECT 2698.900 1597.690 2699.040 1604.850 ;
        RECT 2698.840 1597.370 2699.100 1597.690 ;
        RECT 2702.580 1592.250 2702.720 1610.290 ;
        RECT 2698.380 1591.930 2698.640 1592.250 ;
        RECT 2702.520 1591.930 2702.780 1592.250 ;
        RECT 2694.700 1590.910 2694.960 1591.230 ;
        RECT 2698.380 1590.910 2698.640 1591.230 ;
        RECT 2694.760 1589.045 2694.900 1590.910 ;
        RECT 2694.690 1588.675 2694.970 1589.045 ;
        RECT 2698.440 1582.925 2698.580 1590.910 ;
        RECT 2698.370 1582.555 2698.650 1582.925 ;
        RECT 2683.280 1517.430 2683.540 1517.750 ;
        RECT 2695.150 1503.875 2695.430 1504.245 ;
        RECT 2695.220 1495.890 2695.360 1503.875 ;
        RECT 2695.610 1497.075 2695.890 1497.445 ;
        RECT 2695.680 1496.570 2695.820 1497.075 ;
        RECT 2695.620 1496.250 2695.880 1496.570 ;
        RECT 2698.840 1496.250 2699.100 1496.570 ;
        RECT 2702.520 1496.250 2702.780 1496.570 ;
        RECT 2695.160 1495.570 2695.420 1495.890 ;
        RECT 2698.380 1494.550 2698.640 1494.870 ;
        RECT 2694.700 1492.510 2694.960 1492.830 ;
        RECT 2698.440 1492.570 2698.580 1494.550 ;
        RECT 2694.760 1490.645 2694.900 1492.510 ;
        RECT 2697.520 1492.430 2698.580 1492.570 ;
        RECT 2694.690 1490.275 2694.970 1490.645 ;
        RECT 2694.700 1484.690 2694.960 1485.010 ;
        RECT 2694.760 1483.845 2694.900 1484.690 ;
        RECT 2694.690 1483.475 2694.970 1483.845 ;
        RECT 2697.000 1483.670 2697.260 1483.990 ;
        RECT 2697.520 1483.730 2697.660 1492.430 ;
        RECT 2697.920 1491.830 2698.180 1492.150 ;
        RECT 2697.980 1484.410 2698.120 1491.830 ;
        RECT 2697.980 1484.270 2698.580 1484.410 ;
        RECT 2694.690 1476.675 2694.970 1477.045 ;
        RECT 2694.760 1476.510 2694.900 1476.675 ;
        RECT 2694.700 1476.190 2694.960 1476.510 ;
        RECT 2697.060 1474.130 2697.200 1483.670 ;
        RECT 2697.520 1483.590 2698.120 1483.730 ;
        RECT 2697.460 1481.970 2697.720 1482.290 ;
        RECT 2697.520 1479.570 2697.660 1481.970 ;
        RECT 2697.980 1479.570 2698.120 1483.590 ;
        RECT 2698.440 1482.290 2698.580 1484.270 ;
        RECT 2698.380 1481.970 2698.640 1482.290 ;
        RECT 2697.460 1479.250 2697.720 1479.570 ;
        RECT 2697.920 1479.250 2698.180 1479.570 ;
        RECT 2697.460 1478.570 2697.720 1478.890 ;
        RECT 2697.000 1473.810 2697.260 1474.130 ;
        RECT 2694.700 1470.750 2694.960 1471.070 ;
        RECT 2694.760 1470.245 2694.900 1470.750 ;
        RECT 2694.690 1469.875 2694.970 1470.245 ;
        RECT 2697.520 1466.650 2697.660 1478.570 ;
        RECT 2698.900 1477.610 2699.040 1496.250 ;
        RECT 2701.600 1495.230 2701.860 1495.550 ;
        RECT 2697.980 1477.470 2699.040 1477.610 ;
        RECT 2697.980 1474.130 2698.120 1477.470 ;
        RECT 2697.920 1473.810 2698.180 1474.130 ;
        RECT 2698.840 1473.470 2699.100 1473.790 ;
        RECT 2698.380 1472.790 2698.640 1473.110 ;
        RECT 2697.920 1471.090 2698.180 1471.410 ;
        RECT 2697.460 1466.330 2697.720 1466.650 ;
        RECT 2694.700 1465.310 2694.960 1465.630 ;
        RECT 2694.760 1463.445 2694.900 1465.310 ;
        RECT 2694.690 1463.075 2694.970 1463.445 ;
        RECT 2694.700 1457.490 2694.960 1457.810 ;
        RECT 2694.760 1456.645 2694.900 1457.490 ;
        RECT 2694.690 1456.275 2694.970 1456.645 ;
        RECT 2694.700 1452.050 2694.960 1452.370 ;
        RECT 2694.760 1449.845 2694.900 1452.050 ;
        RECT 2697.460 1451.030 2697.720 1451.350 ;
        RECT 2694.690 1449.475 2694.970 1449.845 ;
        RECT 2697.520 1446.590 2697.660 1451.030 ;
        RECT 2697.980 1446.930 2698.120 1471.090 ;
        RECT 2698.440 1446.930 2698.580 1472.790 ;
        RECT 2698.900 1458.490 2699.040 1473.470 ;
        RECT 2701.660 1471.410 2701.800 1495.230 ;
        RECT 2702.060 1478.910 2702.320 1479.230 ;
        RECT 2702.120 1477.530 2702.260 1478.910 ;
        RECT 2702.580 1478.550 2702.720 1496.250 ;
        RECT 2721.840 1494.890 2722.100 1495.210 ;
        RECT 2721.900 1479.570 2722.040 1494.890 ;
        RECT 2731.500 1494.550 2731.760 1494.870 ;
        RECT 2721.840 1479.250 2722.100 1479.570 ;
        RECT 2702.980 1478.910 2703.240 1479.230 ;
        RECT 2702.520 1478.230 2702.780 1478.550 ;
        RECT 2702.060 1477.210 2702.320 1477.530 ;
        RECT 2702.060 1473.470 2702.320 1473.790 ;
        RECT 2702.120 1472.090 2702.260 1473.470 ;
        RECT 2702.580 1473.110 2702.720 1478.230 ;
        RECT 2703.040 1474.130 2703.180 1478.910 ;
        RECT 2703.900 1478.230 2704.160 1478.550 ;
        RECT 2702.980 1473.810 2703.240 1474.130 ;
        RECT 2702.520 1472.790 2702.780 1473.110 ;
        RECT 2702.060 1471.770 2702.320 1472.090 ;
        RECT 2701.600 1471.090 2701.860 1471.410 ;
        RECT 2701.600 1470.070 2701.860 1470.390 ;
        RECT 2701.660 1460.190 2701.800 1470.070 ;
        RECT 2701.600 1459.870 2701.860 1460.190 ;
        RECT 2702.060 1459.190 2702.320 1459.510 ;
        RECT 2702.120 1458.490 2702.260 1459.190 ;
        RECT 2698.840 1458.170 2699.100 1458.490 ;
        RECT 2702.060 1458.170 2702.320 1458.490 ;
        RECT 2702.520 1456.810 2702.780 1457.130 ;
        RECT 2702.580 1455.770 2702.720 1456.810 ;
        RECT 2702.520 1455.450 2702.780 1455.770 ;
        RECT 2697.920 1446.610 2698.180 1446.930 ;
        RECT 2698.380 1446.610 2698.640 1446.930 ;
        RECT 2697.460 1446.270 2697.720 1446.590 ;
        RECT 2694.700 1443.550 2694.960 1443.870 ;
        RECT 2697.980 1443.610 2698.120 1446.610 ;
        RECT 2694.760 1443.045 2694.900 1443.550 ;
        RECT 2697.520 1443.470 2698.120 1443.610 ;
        RECT 2694.690 1442.675 2694.970 1443.045 ;
        RECT 2697.520 1439.110 2697.660 1443.470 ;
        RECT 2697.920 1442.870 2698.180 1443.190 ;
        RECT 2697.980 1442.170 2698.120 1442.870 ;
        RECT 2697.920 1441.850 2698.180 1442.170 ;
        RECT 2698.440 1441.830 2698.580 1446.610 ;
        RECT 2702.060 1446.270 2702.320 1446.590 ;
        RECT 2703.040 1446.330 2703.180 1473.810 ;
        RECT 2703.960 1470.730 2704.100 1478.230 ;
        RECT 2706.200 1472.790 2706.460 1473.110 ;
        RECT 2706.260 1472.090 2706.400 1472.790 ;
        RECT 2706.200 1471.770 2706.460 1472.090 ;
        RECT 2703.900 1470.410 2704.160 1470.730 ;
        RECT 2731.560 1460.190 2731.700 1494.550 ;
        RECT 2703.900 1459.870 2704.160 1460.190 ;
        RECT 2731.500 1459.870 2731.760 1460.190 ;
        RECT 2703.960 1458.490 2704.100 1459.870 ;
        RECT 2703.900 1458.170 2704.160 1458.490 ;
        RECT 2704.820 1457.150 2705.080 1457.470 ;
        RECT 2704.880 1454.490 2705.020 1457.150 ;
        RECT 2702.120 1442.170 2702.260 1446.270 ;
        RECT 2702.580 1446.190 2703.180 1446.330 ;
        RECT 2703.960 1454.350 2705.020 1454.490 ;
        RECT 2702.060 1441.850 2702.320 1442.170 ;
        RECT 2698.380 1441.570 2698.640 1441.830 ;
        RECT 2698.380 1441.510 2699.040 1441.570 ;
        RECT 2698.440 1441.430 2699.040 1441.510 ;
        RECT 2702.580 1441.490 2702.720 1446.190 ;
        RECT 2702.980 1445.590 2703.240 1445.910 ;
        RECT 2703.040 1442.170 2703.180 1445.590 ;
        RECT 2702.980 1441.850 2703.240 1442.170 ;
        RECT 2703.440 1441.850 2703.700 1442.170 ;
        RECT 2698.380 1440.830 2698.640 1441.150 ;
        RECT 2697.460 1438.790 2697.720 1439.110 ;
        RECT 2694.690 1435.875 2694.970 1436.245 ;
        RECT 2694.700 1435.730 2694.960 1435.875 ;
        RECT 2697.000 1432.330 2697.260 1432.650 ;
        RECT 2697.060 1429.590 2697.200 1432.330 ;
        RECT 2697.520 1430.610 2697.660 1438.790 ;
        RECT 2697.460 1430.290 2697.720 1430.610 ;
        RECT 2697.920 1430.290 2698.180 1430.610 ;
        RECT 2694.690 1429.075 2694.970 1429.445 ;
        RECT 2697.000 1429.270 2697.260 1429.590 ;
        RECT 2694.760 1427.550 2694.900 1429.075 ;
        RECT 2694.700 1427.230 2694.960 1427.550 ;
        RECT 2697.060 1424.830 2697.200 1429.270 ;
        RECT 2697.520 1427.550 2697.660 1430.290 ;
        RECT 2697.460 1427.230 2697.720 1427.550 ;
        RECT 2697.000 1424.510 2697.260 1424.830 ;
        RECT 2697.980 1423.130 2698.120 1430.290 ;
        RECT 2698.440 1428.570 2698.580 1440.830 ;
        RECT 2698.900 1439.450 2699.040 1441.430 ;
        RECT 2702.520 1441.170 2702.780 1441.490 ;
        RECT 2702.580 1440.890 2702.720 1441.170 ;
        RECT 2701.660 1440.750 2702.720 1440.890 ;
        RECT 2698.840 1439.130 2699.100 1439.450 ;
        RECT 2698.840 1437.430 2699.100 1437.750 ;
        RECT 2698.900 1436.730 2699.040 1437.430 ;
        RECT 2698.840 1436.410 2699.100 1436.730 ;
        RECT 2701.660 1433.330 2701.800 1440.750 ;
        RECT 2702.520 1440.150 2702.780 1440.470 ;
        RECT 2702.580 1439.450 2702.720 1440.150 ;
        RECT 2702.520 1439.130 2702.780 1439.450 ;
        RECT 2702.060 1438.790 2702.320 1439.110 ;
        RECT 2701.600 1433.010 2701.860 1433.330 ;
        RECT 2699.760 1432.670 2700.020 1432.990 ;
        RECT 2698.840 1431.990 2699.100 1432.310 ;
        RECT 2699.300 1431.990 2699.560 1432.310 ;
        RECT 2698.900 1431.290 2699.040 1431.990 ;
        RECT 2698.840 1430.970 2699.100 1431.290 ;
        RECT 2699.360 1430.010 2699.500 1431.990 ;
        RECT 2699.820 1430.950 2699.960 1432.670 ;
        RECT 2702.120 1432.650 2702.260 1438.790 ;
        RECT 2703.500 1432.990 2703.640 1441.850 ;
        RECT 2703.440 1432.670 2703.700 1432.990 ;
        RECT 2702.060 1432.330 2702.320 1432.650 ;
        RECT 2699.760 1430.630 2700.020 1430.950 ;
        RECT 2702.120 1430.610 2702.260 1432.330 ;
        RECT 2703.960 1432.310 2704.100 1454.350 ;
        RECT 2703.900 1431.990 2704.160 1432.310 ;
        RECT 2702.060 1430.290 2702.320 1430.610 ;
        RECT 2702.520 1430.290 2702.780 1430.610 ;
        RECT 2698.900 1429.870 2699.500 1430.010 ;
        RECT 2698.900 1428.570 2699.040 1429.870 ;
        RECT 2698.380 1428.250 2698.640 1428.570 ;
        RECT 2698.840 1428.250 2699.100 1428.570 ;
        RECT 2699.760 1427.230 2700.020 1427.550 ;
        RECT 2699.820 1425.850 2699.960 1427.230 ;
        RECT 2699.760 1425.530 2700.020 1425.850 ;
        RECT 2698.840 1424.850 2699.100 1425.170 ;
        RECT 2698.380 1424.510 2698.640 1424.830 ;
        RECT 2697.920 1422.810 2698.180 1423.130 ;
        RECT 2694.690 1422.275 2694.970 1422.645 ;
        RECT 2694.760 1422.110 2694.900 1422.275 ;
        RECT 2694.700 1421.790 2694.960 1422.110 ;
        RECT 2694.700 1416.350 2694.960 1416.670 ;
        RECT 2694.760 1415.845 2694.900 1416.350 ;
        RECT 2694.690 1415.475 2694.970 1415.845 ;
        RECT 2698.440 1412.250 2698.580 1424.510 ;
        RECT 2698.900 1417.690 2699.040 1424.850 ;
        RECT 2698.840 1417.370 2699.100 1417.690 ;
        RECT 2702.580 1412.250 2702.720 1430.290 ;
        RECT 2698.380 1411.930 2698.640 1412.250 ;
        RECT 2702.520 1411.930 2702.780 1412.250 ;
        RECT 2694.700 1410.910 2694.960 1411.230 ;
        RECT 2698.380 1410.910 2698.640 1411.230 ;
        RECT 2694.760 1409.045 2694.900 1410.910 ;
        RECT 2694.690 1408.675 2694.970 1409.045 ;
        RECT 2698.440 1402.925 2698.580 1410.910 ;
        RECT 2698.370 1402.555 2698.650 1402.925 ;
        RECT 2681.900 1317.170 2682.160 1317.490 ;
        RECT 2597.720 1316.830 2597.980 1317.150 ;
        RECT 2514.920 1316.490 2515.180 1316.810 ;
      LAYER met3 ;
        RECT 2362.740 2254.615 2363.110 2254.675 ;
        RECT 2379.325 2254.615 2379.695 2254.675 ;
        RECT 2395.910 2254.615 2396.280 2254.675 ;
        RECT 2412.495 2254.615 2412.865 2254.675 ;
        RECT 2429.075 2254.615 2429.445 2254.675 ;
        RECT 2362.740 2254.315 2367.970 2254.615 ;
        RECT 2379.325 2254.315 2384.555 2254.615 ;
        RECT 2395.910 2254.315 2401.140 2254.615 ;
        RECT 2412.495 2254.315 2417.725 2254.615 ;
        RECT 2429.075 2254.315 2434.305 2254.615 ;
        RECT 2362.740 2254.305 2363.110 2254.315 ;
        RECT 2367.590 2252.425 2367.890 2254.315 ;
        RECT 2379.325 2254.305 2379.695 2254.315 ;
        RECT 2384.175 2252.425 2384.475 2254.315 ;
        RECT 2395.910 2254.305 2396.280 2254.315 ;
        RECT 2400.760 2252.425 2401.060 2254.315 ;
        RECT 2412.495 2254.305 2412.865 2254.315 ;
        RECT 2417.345 2252.425 2417.645 2254.315 ;
        RECT 2429.075 2254.305 2429.445 2254.315 ;
        RECT 2433.925 2252.425 2434.225 2254.315 ;
        RECT 2366.960 2252.410 2367.900 2252.425 ;
        RECT 2368.600 2252.410 2368.945 2252.420 ;
        RECT 2366.960 2252.405 2368.945 2252.410 ;
        RECT 2383.545 2252.410 2384.485 2252.425 ;
        RECT 2385.185 2252.410 2385.530 2252.420 ;
        RECT 2383.545 2252.405 2385.530 2252.410 ;
        RECT 2400.130 2252.410 2401.070 2252.425 ;
        RECT 2401.770 2252.410 2402.115 2252.420 ;
        RECT 2400.130 2252.405 2402.115 2252.410 ;
        RECT 2416.715 2252.410 2417.655 2252.425 ;
        RECT 2418.355 2252.410 2418.700 2252.420 ;
        RECT 2416.715 2252.405 2418.700 2252.410 ;
        RECT 2433.295 2252.410 2434.235 2252.425 ;
        RECT 2434.935 2252.410 2435.280 2252.420 ;
        RECT 2433.295 2252.405 2435.280 2252.410 ;
        RECT 2366.960 2252.110 2369.410 2252.405 ;
        RECT 2366.960 2252.105 2367.900 2252.110 ;
        RECT 2366.960 2250.390 2367.260 2252.105 ;
        RECT 2367.560 2252.075 2367.900 2252.105 ;
        RECT 2368.395 2252.105 2369.410 2252.110 ;
        RECT 2383.545 2252.110 2385.995 2252.405 ;
        RECT 2383.545 2252.105 2384.485 2252.110 ;
        RECT 2368.395 2252.095 2368.945 2252.105 ;
        RECT 2368.600 2252.085 2368.945 2252.095 ;
        RECT 2368.600 2252.075 2368.940 2252.085 ;
        RECT 2367.920 2251.385 2368.265 2251.400 ;
        RECT 2367.920 2251.085 2368.730 2251.385 ;
        RECT 2367.920 2251.055 2368.265 2251.085 ;
        RECT 2383.545 2250.390 2383.845 2252.105 ;
        RECT 2384.145 2252.075 2384.485 2252.105 ;
        RECT 2384.980 2252.105 2385.995 2252.110 ;
        RECT 2400.130 2252.110 2402.580 2252.405 ;
        RECT 2400.130 2252.105 2401.070 2252.110 ;
        RECT 2384.980 2252.095 2385.530 2252.105 ;
        RECT 2385.185 2252.085 2385.530 2252.095 ;
        RECT 2385.185 2252.075 2385.525 2252.085 ;
        RECT 2384.505 2251.385 2384.850 2251.400 ;
        RECT 2384.505 2251.085 2385.315 2251.385 ;
        RECT 2384.505 2251.055 2384.850 2251.085 ;
        RECT 2400.130 2250.390 2400.430 2252.105 ;
        RECT 2400.730 2252.075 2401.070 2252.105 ;
        RECT 2401.565 2252.105 2402.580 2252.110 ;
        RECT 2416.715 2252.110 2419.165 2252.405 ;
        RECT 2416.715 2252.105 2417.655 2252.110 ;
        RECT 2401.565 2252.095 2402.115 2252.105 ;
        RECT 2401.770 2252.085 2402.115 2252.095 ;
        RECT 2401.770 2252.075 2402.110 2252.085 ;
        RECT 2401.090 2251.385 2401.435 2251.400 ;
        RECT 2401.090 2251.085 2401.900 2251.385 ;
        RECT 2401.090 2251.055 2401.435 2251.085 ;
        RECT 2416.715 2250.390 2417.015 2252.105 ;
        RECT 2417.315 2252.075 2417.655 2252.105 ;
        RECT 2418.150 2252.105 2419.165 2252.110 ;
        RECT 2433.295 2252.110 2435.745 2252.405 ;
        RECT 2433.295 2252.105 2434.235 2252.110 ;
        RECT 2418.150 2252.095 2418.700 2252.105 ;
        RECT 2418.355 2252.085 2418.700 2252.095 ;
        RECT 2418.355 2252.075 2418.695 2252.085 ;
        RECT 2417.675 2251.385 2418.020 2251.400 ;
        RECT 2417.675 2251.085 2418.485 2251.385 ;
        RECT 2417.675 2251.055 2418.020 2251.085 ;
        RECT 2433.295 2250.390 2433.595 2252.105 ;
        RECT 2433.895 2252.075 2434.235 2252.105 ;
        RECT 2434.730 2252.105 2435.745 2252.110 ;
        RECT 2434.730 2252.095 2435.280 2252.105 ;
        RECT 2434.935 2252.085 2435.280 2252.095 ;
        RECT 2434.935 2252.075 2435.275 2252.085 ;
        RECT 2434.255 2251.385 2434.600 2251.400 ;
        RECT 2434.255 2251.085 2435.065 2251.385 ;
        RECT 2434.255 2251.055 2434.600 2251.085 ;
        RECT 2366.960 2250.385 2369.615 2250.390 ;
        RECT 2383.545 2250.385 2386.200 2250.390 ;
        RECT 2400.130 2250.385 2402.785 2250.390 ;
        RECT 2416.715 2250.385 2419.370 2250.390 ;
        RECT 2433.295 2250.385 2435.950 2250.390 ;
        RECT 2366.960 2250.365 2369.625 2250.385 ;
        RECT 2383.545 2250.365 2386.210 2250.385 ;
        RECT 2400.130 2250.365 2402.795 2250.385 ;
        RECT 2416.715 2250.365 2419.380 2250.385 ;
        RECT 2433.295 2250.365 2435.960 2250.385 ;
        RECT 2366.960 2250.065 2370.090 2250.365 ;
        RECT 2383.545 2250.065 2386.675 2250.365 ;
        RECT 2400.130 2250.065 2403.260 2250.365 ;
        RECT 2416.715 2250.065 2419.845 2250.365 ;
        RECT 2433.295 2250.065 2436.425 2250.365 ;
        RECT 2366.960 2250.060 2369.625 2250.065 ;
        RECT 2383.545 2250.060 2386.210 2250.065 ;
        RECT 2400.130 2250.060 2402.795 2250.065 ;
        RECT 2416.715 2250.060 2419.380 2250.065 ;
        RECT 2433.295 2250.060 2435.960 2250.065 ;
        RECT 2369.280 2250.035 2369.625 2250.060 ;
        RECT 2385.865 2250.035 2386.210 2250.060 ;
        RECT 2402.450 2250.035 2402.795 2250.060 ;
        RECT 2419.035 2250.035 2419.380 2250.060 ;
        RECT 2435.615 2250.035 2435.960 2250.060 ;
        RECT 2369.300 2249.995 2369.600 2250.035 ;
        RECT 2385.885 2249.995 2386.185 2250.035 ;
        RECT 2402.470 2249.995 2402.770 2250.035 ;
        RECT 2419.055 2249.995 2419.355 2250.035 ;
        RECT 2435.635 2249.995 2435.935 2250.035 ;
        RECT 2368.590 2249.685 2368.930 2249.705 ;
        RECT 2385.175 2249.685 2385.515 2249.705 ;
        RECT 2401.760 2249.685 2402.100 2249.705 ;
        RECT 2418.345 2249.685 2418.685 2249.705 ;
        RECT 2434.925 2249.685 2435.265 2249.705 ;
        RECT 2368.120 2249.385 2368.930 2249.685 ;
        RECT 2384.705 2249.385 2385.515 2249.685 ;
        RECT 2401.290 2249.385 2402.100 2249.685 ;
        RECT 2417.875 2249.385 2418.685 2249.685 ;
        RECT 2434.455 2249.385 2435.265 2249.685 ;
        RECT 2368.590 2249.355 2368.930 2249.385 ;
        RECT 2369.290 2249.355 2369.625 2249.360 ;
        RECT 2385.175 2249.355 2385.515 2249.385 ;
        RECT 2385.875 2249.355 2386.210 2249.360 ;
        RECT 2401.760 2249.355 2402.100 2249.385 ;
        RECT 2402.460 2249.355 2402.795 2249.360 ;
        RECT 2418.345 2249.355 2418.685 2249.385 ;
        RECT 2419.045 2249.355 2419.380 2249.360 ;
        RECT 2434.925 2249.355 2435.265 2249.385 ;
        RECT 2435.625 2249.355 2435.960 2249.360 ;
        RECT 2369.280 2249.345 2369.625 2249.355 ;
        RECT 2385.865 2249.345 2386.210 2249.355 ;
        RECT 2402.450 2249.345 2402.795 2249.355 ;
        RECT 2419.035 2249.345 2419.380 2249.355 ;
        RECT 2435.615 2249.345 2435.960 2249.355 ;
        RECT 2369.280 2249.045 2370.090 2249.345 ;
        RECT 2385.865 2249.045 2386.675 2249.345 ;
        RECT 2402.450 2249.045 2403.260 2249.345 ;
        RECT 2419.035 2249.045 2419.845 2249.345 ;
        RECT 2435.615 2249.045 2436.425 2249.345 ;
        RECT 2369.280 2249.025 2369.625 2249.045 ;
        RECT 2385.865 2249.025 2386.210 2249.045 ;
        RECT 2402.450 2249.025 2402.795 2249.045 ;
        RECT 2419.035 2249.025 2419.380 2249.045 ;
        RECT 2435.615 2249.025 2435.960 2249.045 ;
        RECT 2369.280 2249.015 2369.620 2249.025 ;
        RECT 2385.865 2249.015 2386.205 2249.025 ;
        RECT 2402.450 2249.015 2402.790 2249.025 ;
        RECT 2419.035 2249.015 2419.375 2249.025 ;
        RECT 2435.615 2249.015 2435.955 2249.025 ;
        RECT 2367.240 2249.005 2367.585 2249.015 ;
        RECT 2383.825 2249.005 2384.170 2249.015 ;
        RECT 2400.410 2249.005 2400.755 2249.015 ;
        RECT 2416.995 2249.005 2417.340 2249.015 ;
        RECT 2433.575 2249.005 2433.920 2249.015 ;
        RECT 2366.780 2248.705 2367.585 2249.005 ;
        RECT 2383.365 2248.705 2384.170 2249.005 ;
        RECT 2399.950 2248.705 2400.755 2249.005 ;
        RECT 2416.535 2248.705 2417.340 2249.005 ;
        RECT 2433.115 2248.705 2433.920 2249.005 ;
        RECT 2367.140 2248.695 2367.585 2248.705 ;
        RECT 2383.725 2248.695 2384.170 2248.705 ;
        RECT 2400.310 2248.695 2400.755 2248.705 ;
        RECT 2416.895 2248.695 2417.340 2248.705 ;
        RECT 2433.475 2248.695 2433.920 2248.705 ;
        RECT 2367.240 2248.675 2367.585 2248.695 ;
        RECT 2383.825 2248.675 2384.170 2248.695 ;
        RECT 2400.410 2248.675 2400.755 2248.695 ;
        RECT 2416.995 2248.675 2417.340 2248.695 ;
        RECT 2433.575 2248.675 2433.920 2248.695 ;
        RECT 2690.000 2224.210 2694.000 2224.360 ;
        RECT 2695.125 2224.210 2695.455 2224.225 ;
        RECT 2677.265 2224.090 2677.595 2224.105 ;
        RECT 2690.000 2224.090 2695.455 2224.210 ;
        RECT 2677.265 2223.910 2695.455 2224.090 ;
        RECT 2677.265 2223.790 2694.000 2223.910 ;
        RECT 2695.125 2223.895 2695.455 2223.910 ;
        RECT 2677.265 2223.775 2677.595 2223.790 ;
        RECT 2690.000 2223.760 2694.000 2223.790 ;
        RECT 2690.000 2217.410 2694.000 2217.560 ;
        RECT 2695.585 2217.410 2695.915 2217.425 ;
        RECT 2677.265 2217.290 2677.595 2217.305 ;
        RECT 2690.000 2217.290 2695.915 2217.410 ;
        RECT 2677.265 2217.110 2695.915 2217.290 ;
        RECT 2677.265 2216.990 2694.000 2217.110 ;
        RECT 2695.585 2217.095 2695.915 2217.110 ;
        RECT 2677.265 2216.975 2677.595 2216.990 ;
        RECT 2690.000 2216.960 2694.000 2216.990 ;
        RECT 2690.000 2210.610 2694.000 2210.760 ;
        RECT 2694.665 2210.610 2694.995 2210.625 ;
        RECT 2677.265 2210.490 2677.595 2210.505 ;
        RECT 2690.000 2210.490 2694.995 2210.610 ;
        RECT 2677.265 2210.310 2694.995 2210.490 ;
        RECT 2677.265 2210.190 2694.000 2210.310 ;
        RECT 2694.665 2210.295 2694.995 2210.310 ;
        RECT 2677.265 2210.175 2677.595 2210.190 ;
        RECT 2690.000 2210.160 2694.000 2210.190 ;
        RECT 2690.000 2203.810 2694.000 2203.960 ;
        RECT 2694.665 2203.810 2694.995 2203.825 ;
        RECT 2677.265 2203.690 2677.595 2203.705 ;
        RECT 2690.000 2203.690 2694.995 2203.810 ;
        RECT 2677.265 2203.510 2694.995 2203.690 ;
        RECT 2677.265 2203.390 2694.000 2203.510 ;
        RECT 2694.665 2203.495 2694.995 2203.510 ;
        RECT 2677.265 2203.375 2677.595 2203.390 ;
        RECT 2690.000 2203.360 2694.000 2203.390 ;
        RECT 2690.000 2197.010 2694.000 2197.160 ;
        RECT 2694.665 2197.010 2694.995 2197.025 ;
        RECT 2677.265 2196.890 2677.595 2196.905 ;
        RECT 2690.000 2196.890 2694.995 2197.010 ;
        RECT 2677.265 2196.710 2694.995 2196.890 ;
        RECT 2677.265 2196.590 2694.000 2196.710 ;
        RECT 2694.665 2196.695 2694.995 2196.710 ;
        RECT 2677.265 2196.575 2677.595 2196.590 ;
        RECT 2690.000 2196.560 2694.000 2196.590 ;
        RECT 2690.000 2190.210 2694.000 2190.360 ;
        RECT 2694.665 2190.210 2694.995 2190.225 ;
        RECT 2677.265 2190.090 2677.595 2190.105 ;
        RECT 2690.000 2190.090 2694.995 2190.210 ;
        RECT 2677.265 2189.910 2694.995 2190.090 ;
        RECT 2677.265 2189.790 2694.000 2189.910 ;
        RECT 2694.665 2189.895 2694.995 2189.910 ;
        RECT 2677.265 2189.775 2677.595 2189.790 ;
        RECT 2690.000 2189.760 2694.000 2189.790 ;
        RECT 2690.000 2183.410 2694.000 2183.560 ;
        RECT 2694.665 2183.410 2694.995 2183.425 ;
        RECT 2677.265 2183.290 2677.595 2183.305 ;
        RECT 2690.000 2183.290 2694.995 2183.410 ;
        RECT 2677.265 2183.110 2694.995 2183.290 ;
        RECT 2677.265 2182.990 2694.000 2183.110 ;
        RECT 2694.665 2183.095 2694.995 2183.110 ;
        RECT 2677.265 2182.975 2677.595 2182.990 ;
        RECT 2690.000 2182.960 2694.000 2182.990 ;
        RECT 2690.000 2176.610 2694.000 2176.760 ;
        RECT 2694.665 2176.610 2694.995 2176.625 ;
        RECT 2677.265 2176.490 2677.595 2176.505 ;
        RECT 2690.000 2176.490 2694.995 2176.610 ;
        RECT 2677.265 2176.310 2694.995 2176.490 ;
        RECT 2677.265 2176.190 2694.000 2176.310 ;
        RECT 2694.665 2176.295 2694.995 2176.310 ;
        RECT 2677.265 2176.175 2677.595 2176.190 ;
        RECT 2690.000 2176.160 2694.000 2176.190 ;
        RECT 2690.000 2169.810 2694.000 2169.960 ;
        RECT 2694.665 2169.810 2694.995 2169.825 ;
        RECT 2677.265 2169.690 2677.595 2169.705 ;
        RECT 2690.000 2169.690 2694.995 2169.810 ;
        RECT 2677.265 2169.510 2694.995 2169.690 ;
        RECT 2677.265 2169.390 2694.000 2169.510 ;
        RECT 2694.665 2169.495 2694.995 2169.510 ;
        RECT 2677.265 2169.375 2677.595 2169.390 ;
        RECT 2690.000 2169.360 2694.000 2169.390 ;
        RECT 2690.000 2163.010 2694.000 2163.160 ;
        RECT 2694.665 2163.010 2694.995 2163.025 ;
        RECT 2677.265 2162.890 2677.595 2162.905 ;
        RECT 2690.000 2162.890 2694.995 2163.010 ;
        RECT 2677.265 2162.710 2694.995 2162.890 ;
        RECT 2362.940 2162.620 2363.310 2162.680 ;
        RECT 2380.160 2162.620 2380.530 2162.680 ;
        RECT 2397.380 2162.620 2397.750 2162.680 ;
        RECT 2414.600 2162.620 2414.970 2162.680 ;
        RECT 2431.820 2162.620 2432.190 2162.680 ;
        RECT 2362.940 2162.320 2370.090 2162.620 ;
        RECT 2362.940 2162.310 2363.310 2162.320 ;
        RECT 2367.705 2161.090 2368.005 2162.320 ;
        RECT 2367.205 2160.790 2368.005 2161.090 ;
        RECT 2367.585 2160.745 2368.005 2160.790 ;
        RECT 2367.585 2160.720 2367.885 2160.745 ;
        RECT 2368.735 2160.430 2369.035 2162.320 ;
        RECT 2369.790 2160.465 2370.090 2162.320 ;
        RECT 2380.160 2162.320 2387.310 2162.620 ;
        RECT 2380.160 2162.310 2380.530 2162.320 ;
        RECT 2384.925 2161.090 2385.225 2162.320 ;
        RECT 2384.425 2160.790 2385.225 2161.090 ;
        RECT 2384.805 2160.745 2385.225 2160.790 ;
        RECT 2384.805 2160.720 2385.105 2160.745 ;
        RECT 2368.695 2160.415 2369.035 2160.430 ;
        RECT 2368.685 2160.400 2369.035 2160.415 ;
        RECT 2368.215 2160.100 2369.035 2160.400 ;
        RECT 2369.715 2160.400 2370.090 2160.465 ;
        RECT 2385.955 2160.430 2386.255 2162.320 ;
        RECT 2387.010 2160.465 2387.310 2162.320 ;
        RECT 2397.380 2162.320 2404.530 2162.620 ;
        RECT 2397.380 2162.310 2397.750 2162.320 ;
        RECT 2402.145 2161.090 2402.445 2162.320 ;
        RECT 2401.645 2160.790 2402.445 2161.090 ;
        RECT 2402.025 2160.745 2402.445 2160.790 ;
        RECT 2402.025 2160.720 2402.325 2160.745 ;
        RECT 2385.915 2160.415 2386.255 2160.430 ;
        RECT 2385.905 2160.400 2386.255 2160.415 ;
        RECT 2369.715 2160.100 2370.525 2160.400 ;
        RECT 2385.435 2160.100 2386.255 2160.400 ;
        RECT 2386.935 2160.400 2387.310 2160.465 ;
        RECT 2403.175 2160.430 2403.475 2162.320 ;
        RECT 2404.230 2160.465 2404.530 2162.320 ;
        RECT 2414.600 2162.320 2421.750 2162.620 ;
        RECT 2414.600 2162.310 2414.970 2162.320 ;
        RECT 2419.365 2161.090 2419.665 2162.320 ;
        RECT 2418.865 2160.790 2419.665 2161.090 ;
        RECT 2419.245 2160.745 2419.665 2160.790 ;
        RECT 2419.245 2160.720 2419.545 2160.745 ;
        RECT 2403.135 2160.415 2403.475 2160.430 ;
        RECT 2403.125 2160.400 2403.475 2160.415 ;
        RECT 2386.935 2160.100 2387.745 2160.400 ;
        RECT 2402.655 2160.100 2403.475 2160.400 ;
        RECT 2404.155 2160.400 2404.530 2160.465 ;
        RECT 2420.395 2160.430 2420.695 2162.320 ;
        RECT 2421.450 2160.465 2421.750 2162.320 ;
        RECT 2431.820 2162.320 2438.970 2162.620 ;
        RECT 2677.265 2162.590 2694.000 2162.710 ;
        RECT 2694.665 2162.695 2694.995 2162.710 ;
        RECT 2677.265 2162.575 2677.595 2162.590 ;
        RECT 2690.000 2162.560 2694.000 2162.590 ;
        RECT 2431.820 2162.310 2432.190 2162.320 ;
        RECT 2436.585 2161.090 2436.885 2162.320 ;
        RECT 2436.085 2160.790 2436.885 2161.090 ;
        RECT 2436.465 2160.745 2436.885 2160.790 ;
        RECT 2436.465 2160.720 2436.765 2160.745 ;
        RECT 2420.355 2160.415 2420.695 2160.430 ;
        RECT 2420.345 2160.400 2420.695 2160.415 ;
        RECT 2404.155 2160.100 2404.965 2160.400 ;
        RECT 2419.875 2160.100 2420.695 2160.400 ;
        RECT 2421.375 2160.400 2421.750 2160.465 ;
        RECT 2437.615 2160.430 2437.915 2162.320 ;
        RECT 2438.670 2160.465 2438.970 2162.320 ;
        RECT 2437.575 2160.415 2437.915 2160.430 ;
        RECT 2437.565 2160.400 2437.915 2160.415 ;
        RECT 2421.375 2160.100 2422.185 2160.400 ;
        RECT 2437.095 2160.100 2437.915 2160.400 ;
        RECT 2438.595 2160.400 2438.970 2160.465 ;
        RECT 2438.595 2160.100 2439.405 2160.400 ;
        RECT 2368.685 2160.085 2369.035 2160.100 ;
        RECT 2369.725 2160.085 2370.080 2160.100 ;
        RECT 2385.905 2160.085 2386.255 2160.100 ;
        RECT 2386.945 2160.085 2387.300 2160.100 ;
        RECT 2403.125 2160.085 2403.475 2160.100 ;
        RECT 2404.165 2160.085 2404.520 2160.100 ;
        RECT 2420.345 2160.085 2420.695 2160.100 ;
        RECT 2421.385 2160.085 2421.740 2160.100 ;
        RECT 2437.565 2160.085 2437.915 2160.100 ;
        RECT 2438.605 2160.085 2438.960 2160.100 ;
        RECT 2368.695 2160.080 2369.035 2160.085 ;
        RECT 2368.710 2160.040 2369.010 2160.080 ;
        RECT 2369.780 2160.060 2370.080 2160.085 ;
        RECT 2385.915 2160.080 2386.255 2160.085 ;
        RECT 2385.930 2160.040 2386.230 2160.080 ;
        RECT 2387.000 2160.060 2387.300 2160.085 ;
        RECT 2403.135 2160.080 2403.475 2160.085 ;
        RECT 2403.150 2160.040 2403.450 2160.080 ;
        RECT 2404.220 2160.060 2404.520 2160.085 ;
        RECT 2420.355 2160.080 2420.695 2160.085 ;
        RECT 2420.370 2160.040 2420.670 2160.080 ;
        RECT 2421.440 2160.060 2421.740 2160.085 ;
        RECT 2437.575 2160.080 2437.915 2160.085 ;
        RECT 2437.590 2160.040 2437.890 2160.080 ;
        RECT 2438.660 2160.060 2438.960 2160.085 ;
        RECT 2366.315 2158.765 2366.645 2158.780 ;
        RECT 2368.355 2158.765 2368.685 2158.780 ;
        RECT 2366.315 2158.465 2368.685 2158.765 ;
        RECT 2366.315 2158.450 2366.645 2158.465 ;
        RECT 2368.355 2158.450 2368.685 2158.465 ;
        RECT 2383.535 2158.765 2383.865 2158.780 ;
        RECT 2385.575 2158.765 2385.905 2158.780 ;
        RECT 2383.535 2158.465 2385.905 2158.765 ;
        RECT 2383.535 2158.450 2383.865 2158.465 ;
        RECT 2385.575 2158.450 2385.905 2158.465 ;
        RECT 2400.755 2158.765 2401.085 2158.780 ;
        RECT 2402.795 2158.765 2403.125 2158.780 ;
        RECT 2400.755 2158.465 2403.125 2158.765 ;
        RECT 2400.755 2158.450 2401.085 2158.465 ;
        RECT 2402.795 2158.450 2403.125 2158.465 ;
        RECT 2417.975 2158.765 2418.305 2158.780 ;
        RECT 2420.015 2158.765 2420.345 2158.780 ;
        RECT 2417.975 2158.465 2420.345 2158.765 ;
        RECT 2417.975 2158.450 2418.305 2158.465 ;
        RECT 2420.015 2158.450 2420.345 2158.465 ;
        RECT 2435.195 2158.765 2435.525 2158.780 ;
        RECT 2437.235 2158.765 2437.565 2158.780 ;
        RECT 2435.195 2158.465 2437.565 2158.765 ;
        RECT 2435.195 2158.450 2435.525 2158.465 ;
        RECT 2437.235 2158.450 2437.565 2158.465 ;
        RECT 2369.375 2158.365 2369.705 2158.380 ;
        RECT 2386.595 2158.365 2386.925 2158.380 ;
        RECT 2403.815 2158.365 2404.145 2158.380 ;
        RECT 2421.035 2158.365 2421.365 2158.380 ;
        RECT 2438.255 2158.365 2438.585 2158.380 ;
        RECT 2369.375 2158.065 2370.175 2158.365 ;
        RECT 2386.595 2158.065 2387.395 2158.365 ;
        RECT 2403.815 2158.065 2404.615 2158.365 ;
        RECT 2421.035 2158.065 2421.835 2158.365 ;
        RECT 2438.255 2158.065 2439.055 2158.365 ;
        RECT 2369.375 2158.050 2369.705 2158.065 ;
        RECT 2386.595 2158.050 2386.925 2158.065 ;
        RECT 2403.815 2158.050 2404.145 2158.065 ;
        RECT 2421.035 2158.050 2421.365 2158.065 ;
        RECT 2438.255 2158.050 2438.585 2158.065 ;
        RECT 2368.005 2158.025 2368.335 2158.040 ;
        RECT 2367.545 2157.725 2368.345 2158.025 ;
        RECT 2369.390 2158.020 2369.690 2158.050 ;
        RECT 2385.225 2158.025 2385.555 2158.040 ;
        RECT 2384.765 2157.725 2385.565 2158.025 ;
        RECT 2386.610 2158.020 2386.910 2158.050 ;
        RECT 2402.445 2158.025 2402.775 2158.040 ;
        RECT 2401.985 2157.725 2402.785 2158.025 ;
        RECT 2403.830 2158.020 2404.130 2158.050 ;
        RECT 2419.665 2158.025 2419.995 2158.040 ;
        RECT 2419.205 2157.725 2420.005 2158.025 ;
        RECT 2421.050 2158.020 2421.350 2158.050 ;
        RECT 2436.885 2158.025 2437.215 2158.040 ;
        RECT 2436.425 2157.725 2437.225 2158.025 ;
        RECT 2438.270 2158.020 2438.570 2158.050 ;
        RECT 2368.005 2157.710 2368.335 2157.725 ;
        RECT 2385.225 2157.710 2385.555 2157.725 ;
        RECT 2402.445 2157.710 2402.775 2157.725 ;
        RECT 2419.665 2157.710 2419.995 2157.725 ;
        RECT 2436.885 2157.710 2437.215 2157.725 ;
        RECT 2369.035 2157.685 2369.365 2157.700 ;
        RECT 2386.255 2157.685 2386.585 2157.700 ;
        RECT 2403.475 2157.685 2403.805 2157.700 ;
        RECT 2420.695 2157.685 2421.025 2157.700 ;
        RECT 2437.915 2157.685 2438.245 2157.700 ;
        RECT 2369.035 2157.385 2369.835 2157.685 ;
        RECT 2386.255 2157.385 2387.055 2157.685 ;
        RECT 2403.475 2157.385 2404.275 2157.685 ;
        RECT 2420.695 2157.385 2421.495 2157.685 ;
        RECT 2437.915 2157.385 2438.715 2157.685 ;
        RECT 2369.035 2157.370 2369.420 2157.385 ;
        RECT 2386.255 2157.370 2386.640 2157.385 ;
        RECT 2403.475 2157.370 2403.860 2157.385 ;
        RECT 2420.695 2157.370 2421.080 2157.385 ;
        RECT 2437.915 2157.370 2438.300 2157.385 ;
        RECT 2369.120 2157.360 2369.420 2157.370 ;
        RECT 2386.340 2157.360 2386.640 2157.370 ;
        RECT 2403.560 2157.360 2403.860 2157.370 ;
        RECT 2420.780 2157.360 2421.080 2157.370 ;
        RECT 2438.000 2157.360 2438.300 2157.370 ;
        RECT 2367.675 2156.835 2368.005 2156.850 ;
        RECT 2384.895 2156.835 2385.225 2156.850 ;
        RECT 2402.115 2156.835 2402.445 2156.850 ;
        RECT 2419.335 2156.835 2419.665 2156.850 ;
        RECT 2436.555 2156.835 2436.885 2156.850 ;
        RECT 2367.205 2156.535 2368.005 2156.835 ;
        RECT 2384.425 2156.535 2385.225 2156.835 ;
        RECT 2401.645 2156.535 2402.445 2156.835 ;
        RECT 2418.865 2156.535 2419.665 2156.835 ;
        RECT 2436.085 2156.535 2436.885 2156.835 ;
        RECT 2367.665 2156.530 2368.005 2156.535 ;
        RECT 2384.885 2156.530 2385.225 2156.535 ;
        RECT 2402.105 2156.530 2402.445 2156.535 ;
        RECT 2419.325 2156.530 2419.665 2156.535 ;
        RECT 2436.545 2156.530 2436.885 2156.535 ;
        RECT 2367.675 2156.520 2368.005 2156.530 ;
        RECT 2384.895 2156.520 2385.225 2156.530 ;
        RECT 2402.115 2156.520 2402.445 2156.530 ;
        RECT 2419.335 2156.520 2419.665 2156.530 ;
        RECT 2436.555 2156.520 2436.885 2156.530 ;
        RECT 2690.000 2156.270 2694.000 2156.360 ;
        RECT 2668.890 2156.210 2694.000 2156.270 ;
        RECT 2694.665 2156.210 2694.995 2156.225 ;
        RECT 2668.890 2155.940 2694.995 2156.210 ;
        RECT 2394.825 2139.770 2395.155 2139.785 ;
        RECT 2400.550 2139.770 2400.930 2139.780 ;
        RECT 2394.825 2139.470 2400.930 2139.770 ;
        RECT 2394.825 2139.455 2395.155 2139.470 ;
        RECT 2400.550 2139.460 2400.930 2139.470 ;
        RECT 2428.865 2139.770 2429.195 2139.785 ;
        RECT 2432.750 2139.770 2433.130 2139.780 ;
        RECT 2428.865 2139.470 2433.130 2139.770 ;
        RECT 2428.865 2139.455 2429.195 2139.470 ;
        RECT 2432.750 2139.460 2433.130 2139.470 ;
        RECT 2668.890 2135.305 2669.220 2155.940 ;
        RECT 2690.000 2155.910 2694.995 2155.940 ;
        RECT 2690.000 2155.760 2694.000 2155.910 ;
        RECT 2694.665 2155.895 2694.995 2155.910 ;
        RECT 2523.535 2134.975 2669.220 2135.305 ;
        RECT 2673.570 2149.560 2690.785 2149.680 ;
        RECT 2673.570 2149.410 2694.000 2149.560 ;
        RECT 2694.665 2149.410 2694.995 2149.425 ;
        RECT 2673.570 2149.350 2694.995 2149.410 ;
        RECT 2673.570 2127.775 2673.900 2149.350 ;
        RECT 2690.000 2149.110 2694.995 2149.350 ;
        RECT 2690.000 2148.960 2694.000 2149.110 ;
        RECT 2694.665 2149.095 2694.995 2149.110 ;
        RECT 2690.000 2142.655 2694.000 2142.760 ;
        RECT 2523.535 2127.445 2673.900 2127.775 ;
        RECT 2676.865 2142.610 2694.000 2142.655 ;
        RECT 2694.665 2142.610 2694.995 2142.625 ;
        RECT 2676.865 2142.325 2694.995 2142.610 ;
        RECT 2676.865 2121.795 2677.195 2142.325 ;
        RECT 2690.000 2142.310 2694.995 2142.325 ;
        RECT 2690.000 2142.160 2694.000 2142.310 ;
        RECT 2694.665 2142.295 2694.995 2142.310 ;
        RECT 2690.000 2135.935 2694.000 2135.960 ;
        RECT 2523.535 2121.465 2677.195 2121.795 ;
        RECT 2679.895 2135.810 2694.000 2135.935 ;
        RECT 2694.665 2135.810 2694.995 2135.825 ;
        RECT 2679.895 2135.605 2694.995 2135.810 ;
        RECT 2679.895 2115.850 2680.225 2135.605 ;
        RECT 2690.000 2135.510 2694.995 2135.605 ;
        RECT 2690.000 2135.360 2694.000 2135.510 ;
        RECT 2694.665 2135.495 2694.995 2135.510 ;
        RECT 2690.000 2129.090 2694.000 2129.160 ;
        RECT 2523.535 2115.520 2680.225 2115.850 ;
        RECT 2682.885 2129.010 2694.000 2129.090 ;
        RECT 2694.665 2129.010 2694.995 2129.025 ;
        RECT 2682.885 2128.760 2694.995 2129.010 ;
        RECT 2682.885 2110.205 2683.215 2128.760 ;
        RECT 2690.000 2128.710 2694.995 2128.760 ;
        RECT 2690.000 2128.560 2694.000 2128.710 ;
        RECT 2694.665 2128.695 2694.995 2128.710 ;
        RECT 2698.345 2122.890 2698.675 2122.905 ;
        RECT 2694.910 2122.590 2698.675 2122.890 ;
        RECT 2523.535 2109.875 2683.215 2110.205 ;
        RECT 2686.555 2122.360 2690.745 2122.410 ;
        RECT 2686.555 2122.210 2694.000 2122.360 ;
        RECT 2694.910 2122.210 2695.210 2122.590 ;
        RECT 2698.345 2122.575 2698.675 2122.590 ;
        RECT 2686.555 2122.080 2695.210 2122.210 ;
        RECT 2686.555 2104.200 2686.885 2122.080 ;
        RECT 2690.000 2121.910 2695.210 2122.080 ;
        RECT 2690.000 2121.760 2694.000 2121.910 ;
        RECT 2523.535 2103.870 2686.885 2104.200 ;
        RECT 2368.105 2057.675 2368.475 2057.710 ;
        RECT 2384.430 2057.675 2384.800 2057.710 ;
        RECT 2400.755 2057.675 2401.125 2057.710 ;
        RECT 2417.080 2057.675 2417.450 2057.710 ;
        RECT 2433.405 2057.675 2433.775 2057.710 ;
        RECT 2368.105 2057.375 2370.090 2057.675 ;
        RECT 2368.105 2057.340 2368.475 2057.375 ;
        RECT 2366.405 2053.145 2366.740 2053.165 ;
        RECT 2365.200 2052.845 2366.740 2053.145 ;
        RECT 2361.785 2051.865 2362.120 2052.600 ;
        RECT 2364.230 2052.040 2364.560 2052.435 ;
        RECT 2365.200 2052.040 2365.500 2052.845 ;
        RECT 2366.405 2052.825 2366.740 2052.845 ;
        RECT 2368.345 2052.275 2368.680 2052.600 ;
        RECT 2363.230 2051.470 2363.560 2051.875 ;
        RECT 2364.225 2051.705 2364.560 2052.040 ;
        RECT 2364.945 2051.725 2365.500 2052.040 ;
        RECT 2365.905 2051.875 2366.240 2052.040 ;
        RECT 2366.785 2051.875 2367.120 2052.040 ;
        RECT 2364.945 2051.705 2365.280 2051.725 ;
        RECT 2365.905 2051.710 2368.050 2051.875 ;
        RECT 2368.350 2051.865 2368.680 2052.275 ;
        RECT 2369.790 2051.875 2370.090 2057.375 ;
        RECT 2384.430 2057.375 2386.415 2057.675 ;
        RECT 2384.430 2057.340 2384.800 2057.375 ;
        RECT 2382.730 2053.145 2383.065 2053.165 ;
        RECT 2381.525 2052.845 2383.065 2053.145 ;
        RECT 2363.225 2051.145 2363.560 2051.470 ;
        RECT 2365.910 2051.575 2368.050 2051.710 ;
        RECT 2365.910 2051.305 2366.240 2051.575 ;
        RECT 2366.790 2051.305 2367.120 2051.575 ;
        RECT 2367.750 2051.565 2368.050 2051.575 ;
        RECT 2368.990 2051.575 2370.280 2051.875 ;
        RECT 2378.110 2051.865 2378.445 2052.600 ;
        RECT 2380.555 2052.040 2380.885 2052.435 ;
        RECT 2381.525 2052.040 2381.825 2052.845 ;
        RECT 2382.730 2052.825 2383.065 2052.845 ;
        RECT 2384.670 2052.275 2385.005 2052.600 ;
        RECT 2368.990 2051.565 2369.295 2051.575 ;
        RECT 2367.750 2051.275 2369.295 2051.565 ;
        RECT 2369.945 2051.525 2370.280 2051.575 ;
        RECT 2367.750 2051.260 2369.110 2051.275 ;
        RECT 2369.950 2051.145 2370.280 2051.525 ;
        RECT 2379.555 2051.470 2379.885 2051.875 ;
        RECT 2380.550 2051.705 2380.885 2052.040 ;
        RECT 2381.270 2051.725 2381.825 2052.040 ;
        RECT 2382.230 2051.875 2382.565 2052.040 ;
        RECT 2383.110 2051.875 2383.445 2052.040 ;
        RECT 2381.270 2051.705 2381.605 2051.725 ;
        RECT 2382.230 2051.710 2384.375 2051.875 ;
        RECT 2384.675 2051.865 2385.005 2052.275 ;
        RECT 2386.115 2051.875 2386.415 2057.375 ;
        RECT 2400.755 2057.375 2402.740 2057.675 ;
        RECT 2400.755 2057.340 2401.125 2057.375 ;
        RECT 2399.055 2053.145 2399.390 2053.165 ;
        RECT 2397.850 2052.845 2399.390 2053.145 ;
        RECT 2379.550 2051.145 2379.885 2051.470 ;
        RECT 2382.235 2051.575 2384.375 2051.710 ;
        RECT 2382.235 2051.305 2382.565 2051.575 ;
        RECT 2383.115 2051.305 2383.445 2051.575 ;
        RECT 2384.075 2051.565 2384.375 2051.575 ;
        RECT 2385.315 2051.575 2386.605 2051.875 ;
        RECT 2394.435 2051.865 2394.770 2052.600 ;
        RECT 2396.880 2052.040 2397.210 2052.435 ;
        RECT 2397.850 2052.040 2398.150 2052.845 ;
        RECT 2399.055 2052.825 2399.390 2052.845 ;
        RECT 2400.995 2052.275 2401.330 2052.600 ;
        RECT 2385.315 2051.565 2385.620 2051.575 ;
        RECT 2384.075 2051.275 2385.620 2051.565 ;
        RECT 2386.270 2051.525 2386.605 2051.575 ;
        RECT 2384.075 2051.260 2385.435 2051.275 ;
        RECT 2386.275 2051.145 2386.605 2051.525 ;
        RECT 2395.880 2051.470 2396.210 2051.875 ;
        RECT 2396.875 2051.705 2397.210 2052.040 ;
        RECT 2397.595 2051.725 2398.150 2052.040 ;
        RECT 2398.555 2051.875 2398.890 2052.040 ;
        RECT 2399.435 2051.875 2399.770 2052.040 ;
        RECT 2397.595 2051.705 2397.930 2051.725 ;
        RECT 2398.555 2051.710 2400.700 2051.875 ;
        RECT 2401.000 2051.865 2401.330 2052.275 ;
        RECT 2402.440 2051.875 2402.740 2057.375 ;
        RECT 2417.080 2057.375 2419.065 2057.675 ;
        RECT 2417.080 2057.340 2417.450 2057.375 ;
        RECT 2415.380 2053.145 2415.715 2053.165 ;
        RECT 2414.175 2052.845 2415.715 2053.145 ;
        RECT 2395.875 2051.145 2396.210 2051.470 ;
        RECT 2398.560 2051.575 2400.700 2051.710 ;
        RECT 2398.560 2051.305 2398.890 2051.575 ;
        RECT 2399.440 2051.305 2399.770 2051.575 ;
        RECT 2400.400 2051.565 2400.700 2051.575 ;
        RECT 2401.640 2051.575 2402.930 2051.875 ;
        RECT 2410.760 2051.865 2411.095 2052.600 ;
        RECT 2413.205 2052.040 2413.535 2052.435 ;
        RECT 2414.175 2052.040 2414.475 2052.845 ;
        RECT 2415.380 2052.825 2415.715 2052.845 ;
        RECT 2417.320 2052.275 2417.655 2052.600 ;
        RECT 2401.640 2051.565 2401.945 2051.575 ;
        RECT 2400.400 2051.275 2401.945 2051.565 ;
        RECT 2402.595 2051.525 2402.930 2051.575 ;
        RECT 2400.400 2051.260 2401.760 2051.275 ;
        RECT 2402.600 2051.145 2402.930 2051.525 ;
        RECT 2412.205 2051.470 2412.535 2051.875 ;
        RECT 2413.200 2051.705 2413.535 2052.040 ;
        RECT 2413.920 2051.725 2414.475 2052.040 ;
        RECT 2414.880 2051.875 2415.215 2052.040 ;
        RECT 2415.760 2051.875 2416.095 2052.040 ;
        RECT 2413.920 2051.705 2414.255 2051.725 ;
        RECT 2414.880 2051.710 2417.025 2051.875 ;
        RECT 2417.325 2051.865 2417.655 2052.275 ;
        RECT 2418.765 2051.875 2419.065 2057.375 ;
        RECT 2433.405 2057.375 2435.390 2057.675 ;
        RECT 2433.405 2057.340 2433.775 2057.375 ;
        RECT 2431.705 2053.145 2432.040 2053.165 ;
        RECT 2430.500 2052.845 2432.040 2053.145 ;
        RECT 2412.200 2051.145 2412.535 2051.470 ;
        RECT 2414.885 2051.575 2417.025 2051.710 ;
        RECT 2414.885 2051.305 2415.215 2051.575 ;
        RECT 2415.765 2051.305 2416.095 2051.575 ;
        RECT 2416.725 2051.565 2417.025 2051.575 ;
        RECT 2417.965 2051.575 2419.255 2051.875 ;
        RECT 2427.085 2051.865 2427.420 2052.600 ;
        RECT 2429.530 2052.040 2429.860 2052.435 ;
        RECT 2430.500 2052.040 2430.800 2052.845 ;
        RECT 2431.705 2052.825 2432.040 2052.845 ;
        RECT 2433.645 2052.275 2433.980 2052.600 ;
        RECT 2417.965 2051.565 2418.270 2051.575 ;
        RECT 2416.725 2051.275 2418.270 2051.565 ;
        RECT 2418.920 2051.525 2419.255 2051.575 ;
        RECT 2416.725 2051.260 2418.085 2051.275 ;
        RECT 2418.925 2051.145 2419.255 2051.525 ;
        RECT 2428.530 2051.470 2428.860 2051.875 ;
        RECT 2429.525 2051.705 2429.860 2052.040 ;
        RECT 2430.245 2051.725 2430.800 2052.040 ;
        RECT 2431.205 2051.875 2431.540 2052.040 ;
        RECT 2432.085 2051.875 2432.420 2052.040 ;
        RECT 2430.245 2051.705 2430.580 2051.725 ;
        RECT 2431.205 2051.710 2433.350 2051.875 ;
        RECT 2433.650 2051.865 2433.980 2052.275 ;
        RECT 2435.090 2051.875 2435.390 2057.375 ;
        RECT 2428.525 2051.145 2428.860 2051.470 ;
        RECT 2431.210 2051.575 2433.350 2051.710 ;
        RECT 2431.210 2051.305 2431.540 2051.575 ;
        RECT 2432.090 2051.305 2432.420 2051.575 ;
        RECT 2433.050 2051.565 2433.350 2051.575 ;
        RECT 2434.290 2051.575 2435.580 2051.875 ;
        RECT 2434.290 2051.565 2434.595 2051.575 ;
        RECT 2433.050 2051.275 2434.595 2051.565 ;
        RECT 2435.245 2051.525 2435.580 2051.575 ;
        RECT 2433.050 2051.260 2434.410 2051.275 ;
        RECT 2435.250 2051.145 2435.580 2051.525 ;
        RECT 2677.265 2046.610 2677.595 2046.625 ;
        RECT 2677.265 2046.310 2690.690 2046.610 ;
        RECT 2677.265 2046.295 2677.595 2046.310 ;
        RECT 2690.390 2044.360 2690.690 2046.310 ;
        RECT 2690.000 2044.210 2694.000 2044.360 ;
        RECT 2695.125 2044.210 2695.455 2044.225 ;
        RECT 2690.000 2043.910 2695.455 2044.210 ;
        RECT 2690.000 2043.760 2694.000 2043.910 ;
        RECT 2695.125 2043.895 2695.455 2043.910 ;
        RECT 2400.550 2037.770 2400.930 2037.780 ;
        RECT 2400.550 2037.560 2690.690 2037.770 ;
        RECT 2400.550 2037.470 2694.000 2037.560 ;
        RECT 2400.550 2037.460 2400.930 2037.470 ;
        RECT 2690.000 2037.410 2694.000 2037.470 ;
        RECT 2695.585 2037.410 2695.915 2037.425 ;
        RECT 2690.000 2037.110 2695.915 2037.410 ;
        RECT 2690.000 2036.960 2694.000 2037.110 ;
        RECT 2695.585 2037.095 2695.915 2037.110 ;
        RECT 2409.085 2035.730 2409.415 2035.745 ;
        RECT 2414.350 2035.730 2414.730 2035.740 ;
        RECT 2409.085 2035.430 2414.730 2035.730 ;
        RECT 2409.085 2035.415 2409.415 2035.430 ;
        RECT 2414.350 2035.420 2414.730 2035.430 ;
        RECT 2425.645 2035.730 2425.975 2035.745 ;
        RECT 2428.150 2035.730 2428.530 2035.740 ;
        RECT 2425.645 2035.430 2428.530 2035.730 ;
        RECT 2425.645 2035.415 2425.975 2035.430 ;
        RECT 2428.150 2035.420 2428.530 2035.430 ;
        RECT 2677.265 2033.010 2677.595 2033.025 ;
        RECT 2677.265 2032.710 2690.690 2033.010 ;
        RECT 2677.265 2032.695 2677.595 2032.710 ;
        RECT 2690.390 2030.760 2690.690 2032.710 ;
        RECT 2690.000 2030.610 2694.000 2030.760 ;
        RECT 2694.665 2030.610 2694.995 2030.625 ;
        RECT 2690.000 2030.310 2694.995 2030.610 ;
        RECT 2690.000 2030.160 2694.000 2030.310 ;
        RECT 2694.665 2030.295 2694.995 2030.310 ;
        RECT 2690.000 2023.810 2694.000 2023.960 ;
        RECT 2694.665 2023.810 2694.995 2023.825 ;
        RECT 2690.000 2023.510 2694.995 2023.810 ;
        RECT 2690.000 2023.360 2694.000 2023.510 ;
        RECT 2694.665 2023.495 2694.995 2023.510 ;
        RECT 2677.265 2022.810 2677.595 2022.825 ;
        RECT 2690.390 2022.810 2690.690 2023.360 ;
        RECT 2677.265 2022.510 2690.690 2022.810 ;
        RECT 2677.265 2022.495 2677.595 2022.510 ;
        RECT 2690.000 2017.010 2694.000 2017.160 ;
        RECT 2694.665 2017.010 2694.995 2017.025 ;
        RECT 2690.000 2016.710 2694.995 2017.010 ;
        RECT 2690.000 2016.560 2694.000 2016.710 ;
        RECT 2694.665 2016.695 2694.995 2016.710 ;
        RECT 2677.265 2016.010 2677.595 2016.025 ;
        RECT 2690.390 2016.010 2690.690 2016.560 ;
        RECT 2677.265 2015.710 2690.690 2016.010 ;
        RECT 2677.265 2015.695 2677.595 2015.710 ;
        RECT 2690.000 2010.210 2694.000 2010.360 ;
        RECT 2694.665 2010.210 2694.995 2010.225 ;
        RECT 2690.000 2009.910 2694.995 2010.210 ;
        RECT 2690.000 2009.760 2694.000 2009.910 ;
        RECT 2694.665 2009.895 2694.995 2009.910 ;
        RECT 2681.865 2008.530 2682.195 2008.545 ;
        RECT 2690.390 2008.530 2690.690 2009.760 ;
        RECT 2681.865 2008.230 2690.690 2008.530 ;
        RECT 2681.865 2008.215 2682.195 2008.230 ;
        RECT 2690.000 2003.410 2694.000 2003.560 ;
        RECT 2694.665 2003.410 2694.995 2003.425 ;
        RECT 2690.000 2003.110 2694.995 2003.410 ;
        RECT 2690.000 2002.960 2694.000 2003.110 ;
        RECT 2694.665 2003.095 2694.995 2003.110 ;
        RECT 2681.405 2001.730 2681.735 2001.745 ;
        RECT 2690.390 2001.730 2690.690 2002.960 ;
        RECT 2681.405 2001.430 2690.690 2001.730 ;
        RECT 2681.405 2001.415 2681.735 2001.430 ;
        RECT 2690.000 1996.610 2694.000 1996.760 ;
        RECT 2694.665 1996.610 2694.995 1996.625 ;
        RECT 2690.000 1996.310 2694.995 1996.610 ;
        RECT 2690.000 1996.160 2694.000 1996.310 ;
        RECT 2694.665 1996.295 2694.995 1996.310 ;
        RECT 2677.265 1995.610 2677.595 1995.625 ;
        RECT 2690.390 1995.610 2690.690 1996.160 ;
        RECT 2677.265 1995.310 2690.690 1995.610 ;
        RECT 2677.265 1995.295 2677.595 1995.310 ;
        RECT 2690.000 1989.810 2694.000 1989.960 ;
        RECT 2694.665 1989.810 2694.995 1989.825 ;
        RECT 2690.000 1989.510 2694.995 1989.810 ;
        RECT 2690.000 1989.360 2694.000 1989.510 ;
        RECT 2694.665 1989.495 2694.995 1989.510 ;
        RECT 2680.485 1987.450 2680.815 1987.465 ;
        RECT 2690.390 1987.450 2690.690 1989.360 ;
        RECT 2680.485 1987.150 2690.690 1987.450 ;
        RECT 2680.485 1987.135 2680.815 1987.150 ;
        RECT 2523.535 1982.720 2672.715 1983.050 ;
        RECT 2672.385 1976.680 2672.715 1982.720 ;
        RECT 2690.000 1983.010 2694.000 1983.160 ;
        RECT 2694.665 1983.010 2694.995 1983.025 ;
        RECT 2690.000 1982.710 2694.995 1983.010 ;
        RECT 2690.000 1982.560 2694.000 1982.710 ;
        RECT 2694.665 1982.695 2694.995 1982.710 ;
        RECT 2677.265 1982.010 2677.595 1982.025 ;
        RECT 2690.390 1982.010 2690.690 1982.560 ;
        RECT 2677.265 1981.710 2690.690 1982.010 ;
        RECT 2677.265 1981.695 2677.595 1981.710 ;
        RECT 2672.385 1976.360 2690.700 1976.680 ;
        RECT 2672.385 1976.350 2694.000 1976.360 ;
        RECT 2690.000 1976.210 2694.000 1976.350 ;
        RECT 2694.665 1976.210 2694.995 1976.225 ;
        RECT 2690.000 1975.910 2694.995 1976.210 ;
        RECT 2690.000 1975.760 2694.000 1975.910 ;
        RECT 2694.665 1975.895 2694.995 1975.910 ;
        RECT 2523.535 1975.190 2670.765 1975.520 ;
        RECT 2670.435 1969.750 2670.765 1975.190 ;
        RECT 2670.435 1969.560 2690.840 1969.750 ;
        RECT 2523.535 1969.210 2667.785 1969.540 ;
        RECT 2670.435 1969.420 2694.000 1969.560 ;
        RECT 2523.535 1963.265 2664.705 1963.595 ;
        RECT 2523.535 1957.620 2661.325 1957.950 ;
        RECT 2370.320 1952.685 2370.695 1952.715 ;
        RECT 2388.880 1952.685 2389.255 1952.715 ;
        RECT 2407.440 1952.685 2407.815 1952.715 ;
        RECT 2426.000 1952.685 2426.375 1952.715 ;
        RECT 2444.560 1952.685 2444.935 1952.715 ;
        RECT 2370.320 1952.385 2371.325 1952.685 ;
        RECT 2370.320 1952.345 2370.695 1952.385 ;
        RECT 2371.025 1949.995 2371.325 1952.385 ;
        RECT 2388.880 1952.385 2389.885 1952.685 ;
        RECT 2388.880 1952.345 2389.255 1952.385 ;
        RECT 2389.585 1949.995 2389.885 1952.385 ;
        RECT 2407.440 1952.385 2408.445 1952.685 ;
        RECT 2407.440 1952.345 2407.815 1952.385 ;
        RECT 2408.145 1949.995 2408.445 1952.385 ;
        RECT 2426.000 1952.385 2427.005 1952.685 ;
        RECT 2426.000 1952.345 2426.375 1952.385 ;
        RECT 2426.705 1949.995 2427.005 1952.385 ;
        RECT 2444.560 1952.385 2445.565 1952.685 ;
        RECT 2444.560 1952.345 2444.935 1952.385 ;
        RECT 2445.265 1949.995 2445.565 1952.385 ;
        RECT 2523.535 1951.615 2657.150 1951.945 ;
        RECT 2361.190 1948.925 2371.325 1949.995 ;
        RECT 2379.750 1948.925 2389.885 1949.995 ;
        RECT 2398.310 1948.925 2408.445 1949.995 ;
        RECT 2416.870 1948.925 2427.005 1949.995 ;
        RECT 2435.430 1948.925 2445.565 1949.995 ;
        RECT 2360.800 1948.700 2371.325 1948.925 ;
        RECT 2379.360 1948.700 2389.885 1948.925 ;
        RECT 2397.920 1948.700 2408.445 1948.925 ;
        RECT 2416.480 1948.700 2427.005 1948.925 ;
        RECT 2435.040 1948.700 2445.565 1948.925 ;
        RECT 2360.800 1948.435 2361.640 1948.700 ;
        RECT 2361.190 1947.015 2361.490 1948.435 ;
        RECT 2361.790 1948.155 2362.120 1948.160 ;
        RECT 2361.790 1947.825 2362.525 1948.155 ;
        RECT 2361.790 1947.820 2362.115 1947.825 ;
        RECT 2364.265 1947.600 2364.565 1948.700 ;
        RECT 2364.230 1947.595 2364.565 1947.600 ;
        RECT 2364.230 1947.265 2364.965 1947.595 ;
        RECT 2364.230 1947.260 2364.560 1947.265 ;
        RECT 2365.700 1947.040 2366.000 1948.700 ;
        RECT 2379.360 1948.435 2380.200 1948.700 ;
        RECT 2371.075 1948.160 2371.395 1948.180 ;
        RECT 2368.110 1948.155 2368.445 1948.160 ;
        RECT 2370.075 1948.155 2370.400 1948.160 ;
        RECT 2371.075 1948.155 2371.400 1948.160 ;
        RECT 2368.110 1947.825 2368.845 1948.155 ;
        RECT 2369.815 1947.825 2370.545 1948.155 ;
        RECT 2370.845 1947.825 2371.405 1948.155 ;
        RECT 2368.110 1947.820 2368.445 1947.825 ;
        RECT 2370.075 1947.820 2370.400 1947.825 ;
        RECT 2366.910 1947.595 2367.235 1947.600 ;
        RECT 2366.910 1947.260 2367.465 1947.595 ;
        RECT 2362.125 1947.035 2362.645 1947.040 ;
        RECT 2365.670 1947.035 2366.000 1947.040 ;
        RECT 2362.125 1947.015 2362.855 1947.035 ;
        RECT 2361.190 1946.715 2362.855 1947.015 ;
        RECT 2362.125 1946.705 2362.855 1946.715 ;
        RECT 2365.670 1946.705 2366.405 1947.035 ;
        RECT 2365.670 1946.700 2365.995 1946.705 ;
        RECT 2367.165 1946.465 2367.465 1947.260 ;
        RECT 2370.845 1946.465 2371.145 1947.825 ;
        RECT 2379.750 1947.015 2380.050 1948.435 ;
        RECT 2380.350 1948.155 2380.680 1948.160 ;
        RECT 2380.350 1947.825 2381.085 1948.155 ;
        RECT 2380.350 1947.820 2380.675 1947.825 ;
        RECT 2382.825 1947.600 2383.125 1948.700 ;
        RECT 2382.790 1947.595 2383.125 1947.600 ;
        RECT 2382.790 1947.265 2383.525 1947.595 ;
        RECT 2382.790 1947.260 2383.120 1947.265 ;
        RECT 2384.260 1947.040 2384.560 1948.700 ;
        RECT 2397.920 1948.435 2398.760 1948.700 ;
        RECT 2389.635 1948.160 2389.955 1948.180 ;
        RECT 2386.670 1948.155 2387.005 1948.160 ;
        RECT 2388.635 1948.155 2388.960 1948.160 ;
        RECT 2389.635 1948.155 2389.960 1948.160 ;
        RECT 2386.670 1947.825 2387.405 1948.155 ;
        RECT 2388.375 1947.825 2389.105 1948.155 ;
        RECT 2389.405 1947.825 2389.965 1948.155 ;
        RECT 2386.670 1947.820 2387.005 1947.825 ;
        RECT 2388.635 1947.820 2388.960 1947.825 ;
        RECT 2385.470 1947.595 2385.795 1947.600 ;
        RECT 2385.470 1947.260 2386.025 1947.595 ;
        RECT 2380.685 1947.035 2381.205 1947.040 ;
        RECT 2384.230 1947.035 2384.560 1947.040 ;
        RECT 2380.685 1947.015 2381.415 1947.035 ;
        RECT 2379.750 1946.715 2381.415 1947.015 ;
        RECT 2380.685 1946.705 2381.415 1946.715 ;
        RECT 2384.230 1946.705 2384.965 1947.035 ;
        RECT 2384.230 1946.700 2384.555 1946.705 ;
        RECT 2367.165 1946.165 2371.145 1946.465 ;
        RECT 2372.030 1946.475 2372.355 1946.500 ;
        RECT 2372.030 1946.145 2372.765 1946.475 ;
        RECT 2385.725 1946.465 2386.025 1947.260 ;
        RECT 2389.405 1946.465 2389.705 1947.825 ;
        RECT 2398.310 1947.015 2398.610 1948.435 ;
        RECT 2398.910 1948.155 2399.240 1948.160 ;
        RECT 2398.910 1947.825 2399.645 1948.155 ;
        RECT 2398.910 1947.820 2399.235 1947.825 ;
        RECT 2401.385 1947.600 2401.685 1948.700 ;
        RECT 2401.350 1947.595 2401.685 1947.600 ;
        RECT 2401.350 1947.265 2402.085 1947.595 ;
        RECT 2401.350 1947.260 2401.680 1947.265 ;
        RECT 2402.820 1947.040 2403.120 1948.700 ;
        RECT 2416.480 1948.435 2417.320 1948.700 ;
        RECT 2408.195 1948.160 2408.515 1948.180 ;
        RECT 2405.230 1948.155 2405.565 1948.160 ;
        RECT 2407.195 1948.155 2407.520 1948.160 ;
        RECT 2408.195 1948.155 2408.520 1948.160 ;
        RECT 2405.230 1947.825 2405.965 1948.155 ;
        RECT 2406.935 1947.825 2407.665 1948.155 ;
        RECT 2407.965 1947.825 2408.525 1948.155 ;
        RECT 2405.230 1947.820 2405.565 1947.825 ;
        RECT 2407.195 1947.820 2407.520 1947.825 ;
        RECT 2404.030 1947.595 2404.355 1947.600 ;
        RECT 2404.030 1947.260 2404.585 1947.595 ;
        RECT 2399.245 1947.035 2399.765 1947.040 ;
        RECT 2402.790 1947.035 2403.120 1947.040 ;
        RECT 2399.245 1947.015 2399.975 1947.035 ;
        RECT 2398.310 1946.715 2399.975 1947.015 ;
        RECT 2399.245 1946.705 2399.975 1946.715 ;
        RECT 2402.790 1946.705 2403.525 1947.035 ;
        RECT 2402.790 1946.700 2403.115 1946.705 ;
        RECT 2385.725 1946.165 2389.705 1946.465 ;
        RECT 2390.590 1946.475 2390.915 1946.500 ;
        RECT 2390.590 1946.145 2391.325 1946.475 ;
        RECT 2404.285 1946.465 2404.585 1947.260 ;
        RECT 2407.965 1946.465 2408.265 1947.825 ;
        RECT 2416.870 1947.015 2417.170 1948.435 ;
        RECT 2417.470 1948.155 2417.800 1948.160 ;
        RECT 2417.470 1947.825 2418.205 1948.155 ;
        RECT 2417.470 1947.820 2417.795 1947.825 ;
        RECT 2419.945 1947.600 2420.245 1948.700 ;
        RECT 2419.910 1947.595 2420.245 1947.600 ;
        RECT 2419.910 1947.265 2420.645 1947.595 ;
        RECT 2419.910 1947.260 2420.240 1947.265 ;
        RECT 2421.380 1947.040 2421.680 1948.700 ;
        RECT 2435.040 1948.435 2435.880 1948.700 ;
        RECT 2426.755 1948.160 2427.075 1948.180 ;
        RECT 2423.790 1948.155 2424.125 1948.160 ;
        RECT 2425.755 1948.155 2426.080 1948.160 ;
        RECT 2426.755 1948.155 2427.080 1948.160 ;
        RECT 2423.790 1947.825 2424.525 1948.155 ;
        RECT 2425.495 1947.825 2426.225 1948.155 ;
        RECT 2426.525 1947.825 2427.085 1948.155 ;
        RECT 2423.790 1947.820 2424.125 1947.825 ;
        RECT 2425.755 1947.820 2426.080 1947.825 ;
        RECT 2422.590 1947.595 2422.915 1947.600 ;
        RECT 2422.590 1947.260 2423.145 1947.595 ;
        RECT 2417.805 1947.035 2418.325 1947.040 ;
        RECT 2421.350 1947.035 2421.680 1947.040 ;
        RECT 2417.805 1947.015 2418.535 1947.035 ;
        RECT 2416.870 1946.715 2418.535 1947.015 ;
        RECT 2417.805 1946.705 2418.535 1946.715 ;
        RECT 2421.350 1946.705 2422.085 1947.035 ;
        RECT 2421.350 1946.700 2421.675 1946.705 ;
        RECT 2404.285 1946.165 2408.265 1946.465 ;
        RECT 2409.150 1946.475 2409.475 1946.500 ;
        RECT 2409.150 1946.145 2409.885 1946.475 ;
        RECT 2422.845 1946.465 2423.145 1947.260 ;
        RECT 2426.525 1946.465 2426.825 1947.825 ;
        RECT 2435.430 1947.015 2435.730 1948.435 ;
        RECT 2436.030 1948.155 2436.360 1948.160 ;
        RECT 2436.030 1947.825 2436.765 1948.155 ;
        RECT 2436.030 1947.820 2436.355 1947.825 ;
        RECT 2438.505 1947.600 2438.805 1948.700 ;
        RECT 2438.470 1947.595 2438.805 1947.600 ;
        RECT 2438.470 1947.265 2439.205 1947.595 ;
        RECT 2438.470 1947.260 2438.800 1947.265 ;
        RECT 2439.940 1947.040 2440.240 1948.700 ;
        RECT 2445.315 1948.160 2445.635 1948.180 ;
        RECT 2442.350 1948.155 2442.685 1948.160 ;
        RECT 2444.315 1948.155 2444.640 1948.160 ;
        RECT 2445.315 1948.155 2445.640 1948.160 ;
        RECT 2442.350 1947.825 2443.085 1948.155 ;
        RECT 2444.055 1947.825 2444.785 1948.155 ;
        RECT 2445.085 1947.825 2445.645 1948.155 ;
        RECT 2442.350 1947.820 2442.685 1947.825 ;
        RECT 2444.315 1947.820 2444.640 1947.825 ;
        RECT 2441.150 1947.595 2441.475 1947.600 ;
        RECT 2441.150 1947.260 2441.705 1947.595 ;
        RECT 2436.365 1947.035 2436.885 1947.040 ;
        RECT 2439.910 1947.035 2440.240 1947.040 ;
        RECT 2436.365 1947.015 2437.095 1947.035 ;
        RECT 2435.430 1946.715 2437.095 1947.015 ;
        RECT 2436.365 1946.705 2437.095 1946.715 ;
        RECT 2439.910 1946.705 2440.645 1947.035 ;
        RECT 2439.910 1946.700 2440.235 1946.705 ;
        RECT 2422.845 1946.165 2426.825 1946.465 ;
        RECT 2427.710 1946.475 2428.035 1946.500 ;
        RECT 2427.710 1946.145 2428.445 1946.475 ;
        RECT 2441.405 1946.465 2441.705 1947.260 ;
        RECT 2445.085 1946.465 2445.385 1947.825 ;
        RECT 2441.405 1946.165 2445.385 1946.465 ;
        RECT 2446.270 1946.475 2446.595 1946.500 ;
        RECT 2446.270 1946.145 2447.005 1946.475 ;
        RECT 2372.030 1946.140 2372.355 1946.145 ;
        RECT 2390.590 1946.140 2390.915 1946.145 ;
        RECT 2409.150 1946.140 2409.475 1946.145 ;
        RECT 2427.710 1946.140 2428.035 1946.145 ;
        RECT 2446.270 1946.140 2446.595 1946.145 ;
        RECT 2656.820 1942.620 2657.150 1951.615 ;
        RECT 2660.995 1949.180 2661.325 1957.620 ;
        RECT 2664.375 1955.640 2664.705 1963.265 ;
        RECT 2667.455 1962.895 2667.785 1969.210 ;
        RECT 2690.000 1969.410 2694.000 1969.420 ;
        RECT 2694.665 1969.410 2694.995 1969.425 ;
        RECT 2690.000 1969.110 2694.995 1969.410 ;
        RECT 2690.000 1968.960 2694.000 1969.110 ;
        RECT 2694.665 1969.095 2694.995 1969.110 ;
        RECT 2667.455 1962.760 2691.835 1962.895 ;
        RECT 2667.455 1962.610 2694.000 1962.760 ;
        RECT 2694.665 1962.610 2694.995 1962.625 ;
        RECT 2667.455 1962.565 2694.995 1962.610 ;
        RECT 2690.000 1962.310 2694.995 1962.565 ;
        RECT 2690.000 1962.160 2694.000 1962.310 ;
        RECT 2694.665 1962.295 2694.995 1962.310 ;
        RECT 2690.000 1955.810 2694.000 1955.960 ;
        RECT 2694.665 1955.810 2694.995 1955.825 ;
        RECT 2690.000 1955.640 2694.995 1955.810 ;
        RECT 2664.375 1955.510 2694.995 1955.640 ;
        RECT 2664.375 1955.360 2694.000 1955.510 ;
        RECT 2694.665 1955.495 2694.995 1955.510 ;
        RECT 2664.375 1955.310 2691.140 1955.360 ;
        RECT 2660.995 1949.160 2691.240 1949.180 ;
        RECT 2660.995 1949.010 2694.000 1949.160 ;
        RECT 2694.665 1949.010 2694.995 1949.025 ;
        RECT 2660.995 1948.850 2694.995 1949.010 ;
        RECT 2690.000 1948.710 2694.995 1948.850 ;
        RECT 2690.000 1948.560 2694.000 1948.710 ;
        RECT 2694.665 1948.695 2694.995 1948.710 ;
        RECT 2698.345 1942.890 2698.675 1942.905 ;
        RECT 2656.820 1942.360 2690.940 1942.620 ;
        RECT 2694.910 1942.590 2698.675 1942.890 ;
        RECT 2656.820 1942.290 2694.000 1942.360 ;
        RECT 2690.000 1942.210 2694.000 1942.290 ;
        RECT 2694.910 1942.210 2695.210 1942.590 ;
        RECT 2698.345 1942.575 2698.675 1942.590 ;
        RECT 2690.000 1941.910 2695.210 1942.210 ;
        RECT 2690.000 1941.760 2694.000 1941.910 ;
        RECT 2433.670 1932.370 2434.050 1932.380 ;
        RECT 2434.385 1932.370 2434.715 1932.385 ;
        RECT 2433.670 1932.070 2434.715 1932.370 ;
        RECT 2433.670 1932.060 2434.050 1932.070 ;
        RECT 2434.385 1932.055 2434.715 1932.070 ;
        RECT 2677.265 1864.370 2677.595 1864.385 ;
        RECT 2677.265 1864.360 2690.540 1864.370 ;
        RECT 2677.265 1864.210 2694.000 1864.360 ;
        RECT 2695.125 1864.210 2695.455 1864.225 ;
        RECT 2677.265 1864.070 2695.455 1864.210 ;
        RECT 2677.265 1864.055 2677.595 1864.070 ;
        RECT 2690.000 1863.910 2695.455 1864.070 ;
        RECT 2690.000 1863.760 2694.000 1863.910 ;
        RECT 2695.125 1863.895 2695.455 1863.910 ;
        RECT 2677.265 1857.570 2677.595 1857.585 ;
        RECT 2677.265 1857.560 2690.540 1857.570 ;
        RECT 2677.265 1857.410 2694.000 1857.560 ;
        RECT 2695.585 1857.410 2695.915 1857.425 ;
        RECT 2677.265 1857.270 2695.915 1857.410 ;
        RECT 2677.265 1857.255 2677.595 1857.270 ;
        RECT 2690.000 1857.110 2695.915 1857.270 ;
        RECT 2690.000 1856.960 2694.000 1857.110 ;
        RECT 2695.585 1857.095 2695.915 1857.110 ;
        RECT 2414.350 1850.770 2414.730 1850.780 ;
        RECT 2414.350 1850.760 2690.540 1850.770 ;
        RECT 2414.350 1850.610 2694.000 1850.760 ;
        RECT 2694.665 1850.610 2694.995 1850.625 ;
        RECT 2414.350 1850.470 2694.995 1850.610 ;
        RECT 2414.350 1850.460 2414.730 1850.470 ;
        RECT 2690.000 1850.310 2694.995 1850.470 ;
        RECT 2690.000 1850.160 2694.000 1850.310 ;
        RECT 2694.665 1850.295 2694.995 1850.310 ;
        RECT 2677.265 1843.970 2677.595 1843.985 ;
        RECT 2677.265 1843.960 2690.540 1843.970 ;
        RECT 2677.265 1843.810 2694.000 1843.960 ;
        RECT 2694.665 1843.810 2694.995 1843.825 ;
        RECT 2677.265 1843.670 2694.995 1843.810 ;
        RECT 2677.265 1843.655 2677.595 1843.670 ;
        RECT 2690.000 1843.510 2694.995 1843.670 ;
        RECT 2690.000 1843.360 2694.000 1843.510 ;
        RECT 2694.665 1843.495 2694.995 1843.510 ;
        RECT 2677.265 1837.170 2677.595 1837.185 ;
        RECT 2677.265 1837.160 2690.540 1837.170 ;
        RECT 2677.265 1837.010 2694.000 1837.160 ;
        RECT 2694.665 1837.010 2694.995 1837.025 ;
        RECT 2677.265 1836.870 2694.995 1837.010 ;
        RECT 2677.265 1836.855 2677.595 1836.870 ;
        RECT 2690.000 1836.710 2694.995 1836.870 ;
        RECT 2690.000 1836.560 2694.000 1836.710 ;
        RECT 2694.665 1836.695 2694.995 1836.710 ;
        RECT 2677.265 1830.370 2677.595 1830.385 ;
        RECT 2677.265 1830.360 2690.540 1830.370 ;
        RECT 2677.265 1830.210 2694.000 1830.360 ;
        RECT 2694.665 1830.210 2694.995 1830.225 ;
        RECT 2677.265 1830.070 2694.995 1830.210 ;
        RECT 2677.265 1830.055 2677.595 1830.070 ;
        RECT 2690.000 1829.910 2694.995 1830.070 ;
        RECT 2690.000 1829.760 2694.000 1829.910 ;
        RECT 2694.665 1829.895 2694.995 1829.910 ;
        RECT 2682.785 1823.570 2683.115 1823.585 ;
        RECT 2682.785 1823.560 2690.540 1823.570 ;
        RECT 2682.785 1823.410 2694.000 1823.560 ;
        RECT 2694.665 1823.410 2694.995 1823.425 ;
        RECT 2682.785 1823.270 2694.995 1823.410 ;
        RECT 2682.785 1823.255 2683.115 1823.270 ;
        RECT 2690.000 1823.110 2694.995 1823.270 ;
        RECT 2690.000 1822.960 2694.000 1823.110 ;
        RECT 2694.665 1823.095 2694.995 1823.110 ;
        RECT 2682.325 1816.770 2682.655 1816.785 ;
        RECT 2682.325 1816.760 2690.540 1816.770 ;
        RECT 2682.325 1816.610 2694.000 1816.760 ;
        RECT 2694.665 1816.610 2694.995 1816.625 ;
        RECT 2682.325 1816.470 2694.995 1816.610 ;
        RECT 2682.325 1816.455 2682.655 1816.470 ;
        RECT 2690.000 1816.310 2694.995 1816.470 ;
        RECT 2690.000 1816.160 2694.000 1816.310 ;
        RECT 2694.665 1816.295 2694.995 1816.310 ;
        RECT 2677.265 1809.970 2677.595 1809.985 ;
        RECT 2677.265 1809.960 2690.540 1809.970 ;
        RECT 2677.265 1809.810 2694.000 1809.960 ;
        RECT 2694.665 1809.810 2694.995 1809.825 ;
        RECT 2677.265 1809.670 2694.995 1809.810 ;
        RECT 2677.265 1809.655 2677.595 1809.670 ;
        RECT 2690.000 1809.510 2694.995 1809.670 ;
        RECT 2690.000 1809.360 2694.000 1809.510 ;
        RECT 2694.665 1809.495 2694.995 1809.510 ;
        RECT 2523.535 1805.750 2677.370 1806.080 ;
        RECT 2523.535 1798.220 2673.170 1798.550 ;
        RECT 2523.535 1792.240 2670.050 1792.570 ;
        RECT 2376.965 1789.345 2377.335 1789.715 ;
        RECT 2392.225 1789.345 2392.595 1789.715 ;
        RECT 2407.485 1789.345 2407.855 1789.715 ;
        RECT 2422.745 1789.345 2423.115 1789.715 ;
        RECT 2438.005 1789.345 2438.375 1789.715 ;
        RECT 2377.000 1786.530 2377.300 1789.345 ;
        RECT 2392.260 1786.530 2392.560 1789.345 ;
        RECT 2407.520 1786.530 2407.820 1789.345 ;
        RECT 2422.780 1786.530 2423.080 1789.345 ;
        RECT 2438.040 1786.530 2438.340 1789.345 ;
        RECT 2376.995 1786.175 2377.300 1786.530 ;
        RECT 2392.255 1786.175 2392.560 1786.530 ;
        RECT 2407.515 1786.175 2407.820 1786.530 ;
        RECT 2422.775 1786.175 2423.080 1786.530 ;
        RECT 2438.035 1786.175 2438.340 1786.530 ;
        RECT 2523.535 1786.295 2665.850 1786.625 ;
        RECT 2376.995 1785.770 2377.295 1786.175 ;
        RECT 2392.255 1785.770 2392.555 1786.175 ;
        RECT 2407.515 1785.770 2407.815 1786.175 ;
        RECT 2422.775 1785.770 2423.075 1786.175 ;
        RECT 2438.035 1785.770 2438.335 1786.175 ;
        RECT 2372.765 1785.470 2377.295 1785.770 ;
        RECT 2388.025 1785.470 2392.555 1785.770 ;
        RECT 2403.285 1785.470 2407.815 1785.770 ;
        RECT 2418.545 1785.470 2423.075 1785.770 ;
        RECT 2433.805 1785.470 2438.335 1785.770 ;
        RECT 2372.765 1784.600 2373.065 1785.470 ;
        RECT 2375.560 1785.145 2375.860 1785.470 ;
        RECT 2376.285 1785.145 2376.615 1785.155 ;
        RECT 2374.375 1784.845 2376.615 1785.145 ;
        RECT 2372.685 1784.595 2373.065 1784.600 ;
        RECT 2372.455 1784.265 2373.185 1784.595 ;
        RECT 2373.645 1784.245 2373.965 1784.625 ;
        RECT 2373.645 1784.055 2373.975 1784.245 ;
        RECT 2374.375 1784.055 2374.675 1784.845 ;
        RECT 2375.560 1784.155 2375.860 1784.845 ;
        RECT 2376.275 1784.795 2376.615 1784.845 ;
        RECT 2388.025 1784.600 2388.325 1785.470 ;
        RECT 2390.820 1785.145 2391.120 1785.470 ;
        RECT 2391.545 1785.145 2391.875 1785.155 ;
        RECT 2389.635 1784.845 2391.875 1785.145 ;
        RECT 2387.945 1784.595 2388.325 1784.600 ;
        RECT 2387.715 1784.265 2388.445 1784.595 ;
        RECT 2388.905 1784.245 2389.225 1784.625 ;
        RECT 2373.645 1783.705 2373.980 1784.055 ;
        RECT 2374.355 1784.040 2374.675 1784.055 ;
        RECT 2374.355 1783.705 2374.695 1784.040 ;
        RECT 2375.355 1783.815 2376.135 1784.155 ;
        RECT 2375.560 1783.810 2376.135 1783.815 ;
        RECT 2375.795 1783.805 2376.135 1783.810 ;
        RECT 2375.805 1783.775 2376.135 1783.805 ;
        RECT 2388.905 1784.055 2389.235 1784.245 ;
        RECT 2389.635 1784.055 2389.935 1784.845 ;
        RECT 2390.820 1784.155 2391.120 1784.845 ;
        RECT 2391.535 1784.795 2391.875 1784.845 ;
        RECT 2403.285 1784.600 2403.585 1785.470 ;
        RECT 2406.080 1785.145 2406.380 1785.470 ;
        RECT 2406.805 1785.145 2407.135 1785.155 ;
        RECT 2404.895 1784.845 2407.135 1785.145 ;
        RECT 2403.205 1784.595 2403.585 1784.600 ;
        RECT 2402.975 1784.265 2403.705 1784.595 ;
        RECT 2404.165 1784.245 2404.485 1784.625 ;
        RECT 2388.905 1783.705 2389.240 1784.055 ;
        RECT 2389.615 1784.040 2389.935 1784.055 ;
        RECT 2389.615 1783.705 2389.955 1784.040 ;
        RECT 2390.615 1783.815 2391.395 1784.155 ;
        RECT 2390.820 1783.810 2391.395 1783.815 ;
        RECT 2391.055 1783.805 2391.395 1783.810 ;
        RECT 2391.065 1783.775 2391.395 1783.805 ;
        RECT 2404.165 1784.055 2404.495 1784.245 ;
        RECT 2404.895 1784.055 2405.195 1784.845 ;
        RECT 2406.080 1784.155 2406.380 1784.845 ;
        RECT 2406.795 1784.795 2407.135 1784.845 ;
        RECT 2418.545 1784.600 2418.845 1785.470 ;
        RECT 2421.340 1785.145 2421.640 1785.470 ;
        RECT 2422.065 1785.145 2422.395 1785.155 ;
        RECT 2420.155 1784.845 2422.395 1785.145 ;
        RECT 2418.465 1784.595 2418.845 1784.600 ;
        RECT 2418.235 1784.265 2418.965 1784.595 ;
        RECT 2419.425 1784.245 2419.745 1784.625 ;
        RECT 2404.165 1783.705 2404.500 1784.055 ;
        RECT 2404.875 1784.040 2405.195 1784.055 ;
        RECT 2404.875 1783.705 2405.215 1784.040 ;
        RECT 2405.875 1783.815 2406.655 1784.155 ;
        RECT 2406.080 1783.810 2406.655 1783.815 ;
        RECT 2406.315 1783.805 2406.655 1783.810 ;
        RECT 2406.325 1783.775 2406.655 1783.805 ;
        RECT 2419.425 1784.055 2419.755 1784.245 ;
        RECT 2420.155 1784.055 2420.455 1784.845 ;
        RECT 2421.340 1784.155 2421.640 1784.845 ;
        RECT 2422.055 1784.795 2422.395 1784.845 ;
        RECT 2433.805 1784.600 2434.105 1785.470 ;
        RECT 2436.600 1785.145 2436.900 1785.470 ;
        RECT 2437.325 1785.145 2437.655 1785.155 ;
        RECT 2435.415 1784.845 2437.655 1785.145 ;
        RECT 2433.725 1784.595 2434.105 1784.600 ;
        RECT 2433.495 1784.265 2434.225 1784.595 ;
        RECT 2434.685 1784.245 2435.005 1784.625 ;
        RECT 2419.425 1783.705 2419.760 1784.055 ;
        RECT 2420.135 1784.040 2420.455 1784.055 ;
        RECT 2420.135 1783.705 2420.475 1784.040 ;
        RECT 2421.135 1783.815 2421.915 1784.155 ;
        RECT 2421.340 1783.810 2421.915 1783.815 ;
        RECT 2421.575 1783.805 2421.915 1783.810 ;
        RECT 2421.585 1783.775 2421.915 1783.805 ;
        RECT 2434.685 1784.055 2435.015 1784.245 ;
        RECT 2435.415 1784.055 2435.715 1784.845 ;
        RECT 2436.600 1784.155 2436.900 1784.845 ;
        RECT 2437.315 1784.795 2437.655 1784.845 ;
        RECT 2434.685 1783.705 2435.020 1784.055 ;
        RECT 2435.395 1784.040 2435.715 1784.055 ;
        RECT 2435.395 1783.705 2435.735 1784.040 ;
        RECT 2436.395 1783.815 2437.175 1784.155 ;
        RECT 2436.600 1783.810 2437.175 1783.815 ;
        RECT 2436.835 1783.805 2437.175 1783.810 ;
        RECT 2436.845 1783.775 2437.175 1783.805 ;
        RECT 2374.925 1783.175 2375.655 1783.505 ;
        RECT 2376.470 1783.495 2376.820 1783.500 ;
        RECT 2374.925 1783.165 2375.405 1783.175 ;
        RECT 2376.470 1783.145 2377.205 1783.495 ;
        RECT 2377.505 1783.165 2378.245 1783.495 ;
        RECT 2379.365 1783.475 2379.725 1783.480 ;
        RECT 2377.505 1783.155 2377.835 1783.165 ;
        RECT 2379.205 1783.145 2379.935 1783.475 ;
        RECT 2390.185 1783.175 2390.915 1783.505 ;
        RECT 2391.730 1783.495 2392.080 1783.500 ;
        RECT 2390.185 1783.165 2390.665 1783.175 ;
        RECT 2391.730 1783.145 2392.465 1783.495 ;
        RECT 2392.765 1783.165 2393.505 1783.495 ;
        RECT 2394.625 1783.475 2394.985 1783.480 ;
        RECT 2392.765 1783.155 2393.095 1783.165 ;
        RECT 2394.465 1783.145 2395.195 1783.475 ;
        RECT 2405.445 1783.175 2406.175 1783.505 ;
        RECT 2406.990 1783.495 2407.340 1783.500 ;
        RECT 2405.445 1783.165 2405.925 1783.175 ;
        RECT 2406.990 1783.145 2407.725 1783.495 ;
        RECT 2408.025 1783.165 2408.765 1783.495 ;
        RECT 2409.885 1783.475 2410.245 1783.480 ;
        RECT 2408.025 1783.155 2408.355 1783.165 ;
        RECT 2409.725 1783.145 2410.455 1783.475 ;
        RECT 2420.705 1783.175 2421.435 1783.505 ;
        RECT 2422.250 1783.495 2422.600 1783.500 ;
        RECT 2420.705 1783.165 2421.185 1783.175 ;
        RECT 2422.250 1783.145 2422.985 1783.495 ;
        RECT 2423.285 1783.165 2424.025 1783.495 ;
        RECT 2425.145 1783.475 2425.505 1783.480 ;
        RECT 2423.285 1783.155 2423.615 1783.165 ;
        RECT 2424.985 1783.145 2425.715 1783.475 ;
        RECT 2435.965 1783.175 2436.695 1783.505 ;
        RECT 2437.510 1783.495 2437.860 1783.500 ;
        RECT 2435.965 1783.165 2436.445 1783.175 ;
        RECT 2437.510 1783.145 2438.245 1783.495 ;
        RECT 2438.545 1783.165 2439.285 1783.495 ;
        RECT 2440.405 1783.475 2440.765 1783.480 ;
        RECT 2438.545 1783.155 2438.875 1783.165 ;
        RECT 2440.245 1783.145 2440.975 1783.475 ;
        RECT 2376.470 1783.140 2376.820 1783.145 ;
        RECT 2379.365 1783.140 2379.725 1783.145 ;
        RECT 2391.730 1783.140 2392.080 1783.145 ;
        RECT 2394.625 1783.140 2394.985 1783.145 ;
        RECT 2406.990 1783.140 2407.340 1783.145 ;
        RECT 2409.885 1783.140 2410.245 1783.145 ;
        RECT 2422.250 1783.140 2422.600 1783.145 ;
        RECT 2425.145 1783.140 2425.505 1783.145 ;
        RECT 2437.510 1783.140 2437.860 1783.145 ;
        RECT 2440.405 1783.140 2440.765 1783.145 ;
        RECT 2523.535 1780.650 2662.610 1780.980 ;
        RECT 2523.535 1769.180 2657.930 1769.510 ;
        RECT 2657.600 1762.475 2657.930 1769.180 ;
        RECT 2662.280 1769.315 2662.610 1780.650 ;
        RECT 2665.520 1775.915 2665.850 1786.295 ;
        RECT 2669.720 1782.880 2670.050 1792.240 ;
        RECT 2672.840 1789.840 2673.170 1798.220 ;
        RECT 2677.040 1796.200 2677.370 1805.750 ;
        RECT 2680.945 1803.170 2681.275 1803.185 ;
        RECT 2680.945 1803.160 2690.540 1803.170 ;
        RECT 2680.945 1803.010 2694.000 1803.160 ;
        RECT 2694.665 1803.010 2694.995 1803.025 ;
        RECT 2680.945 1802.870 2694.995 1803.010 ;
        RECT 2680.945 1802.855 2681.275 1802.870 ;
        RECT 2690.000 1802.710 2694.995 1802.870 ;
        RECT 2690.000 1802.560 2694.000 1802.710 ;
        RECT 2694.665 1802.695 2694.995 1802.710 ;
        RECT 2690.000 1796.210 2694.000 1796.360 ;
        RECT 2694.665 1796.210 2694.995 1796.225 ;
        RECT 2690.000 1796.200 2694.995 1796.210 ;
        RECT 2677.040 1795.910 2694.995 1796.200 ;
        RECT 2677.040 1795.870 2694.000 1795.910 ;
        RECT 2694.665 1795.895 2694.995 1795.910 ;
        RECT 2690.000 1795.760 2694.000 1795.870 ;
        RECT 2672.840 1789.560 2691.055 1789.840 ;
        RECT 2672.840 1789.510 2694.000 1789.560 ;
        RECT 2690.000 1789.410 2694.000 1789.510 ;
        RECT 2694.665 1789.410 2694.995 1789.425 ;
        RECT 2690.000 1789.110 2694.995 1789.410 ;
        RECT 2690.000 1788.960 2694.000 1789.110 ;
        RECT 2694.665 1789.095 2694.995 1789.110 ;
        RECT 2669.720 1782.760 2691.175 1782.880 ;
        RECT 2669.720 1782.610 2694.000 1782.760 ;
        RECT 2694.665 1782.610 2694.995 1782.625 ;
        RECT 2669.720 1782.550 2694.995 1782.610 ;
        RECT 2690.000 1782.310 2694.995 1782.550 ;
        RECT 2690.000 1782.160 2694.000 1782.310 ;
        RECT 2694.665 1782.295 2694.995 1782.310 ;
        RECT 2690.000 1775.915 2694.000 1775.960 ;
        RECT 2665.520 1775.810 2694.000 1775.915 ;
        RECT 2694.665 1775.810 2694.995 1775.825 ;
        RECT 2665.520 1775.585 2694.995 1775.810 ;
        RECT 2690.000 1775.510 2694.995 1775.585 ;
        RECT 2690.000 1775.360 2694.000 1775.510 ;
        RECT 2694.665 1775.495 2694.995 1775.510 ;
        RECT 2662.280 1769.160 2691.535 1769.315 ;
        RECT 2662.280 1769.010 2694.000 1769.160 ;
        RECT 2694.665 1769.010 2694.995 1769.025 ;
        RECT 2662.280 1768.985 2694.995 1769.010 ;
        RECT 2690.000 1768.710 2694.995 1768.985 ;
        RECT 2690.000 1768.560 2694.000 1768.710 ;
        RECT 2694.665 1768.695 2694.995 1768.710 ;
        RECT 2698.345 1762.890 2698.675 1762.905 ;
        RECT 2694.910 1762.590 2698.675 1762.890 ;
        RECT 2657.600 1762.360 2691.415 1762.475 ;
        RECT 2657.600 1762.210 2694.000 1762.360 ;
        RECT 2694.910 1762.210 2695.210 1762.590 ;
        RECT 2698.345 1762.575 2698.675 1762.590 ;
        RECT 2657.600 1762.145 2695.210 1762.210 ;
        RECT 2690.000 1761.910 2695.210 1762.145 ;
        RECT 2690.000 1761.760 2694.000 1761.910 ;
        RECT 2363.100 1709.615 2363.470 1709.675 ;
        RECT 2379.685 1709.615 2380.055 1709.675 ;
        RECT 2396.270 1709.620 2396.640 1709.680 ;
        RECT 2412.855 1709.625 2413.225 1709.685 ;
        RECT 2429.435 1709.625 2429.805 1709.685 ;
        RECT 2363.100 1709.315 2368.255 1709.615 ;
        RECT 2379.685 1709.315 2384.840 1709.615 ;
        RECT 2396.270 1709.320 2401.425 1709.620 ;
        RECT 2412.855 1709.325 2418.010 1709.625 ;
        RECT 2429.435 1709.325 2434.590 1709.625 ;
        RECT 2363.100 1709.305 2363.470 1709.315 ;
        RECT 2367.950 1707.420 2368.250 1709.315 ;
        RECT 2379.685 1709.305 2380.055 1709.315 ;
        RECT 2384.535 1707.420 2384.835 1709.315 ;
        RECT 2396.270 1709.310 2396.640 1709.320 ;
        RECT 2401.120 1707.425 2401.420 1709.320 ;
        RECT 2412.855 1709.315 2413.225 1709.325 ;
        RECT 2417.705 1707.430 2418.005 1709.325 ;
        RECT 2429.435 1709.315 2429.805 1709.325 ;
        RECT 2434.285 1707.430 2434.585 1709.325 ;
        RECT 2367.320 1707.405 2368.260 1707.420 ;
        RECT 2368.960 1707.405 2369.305 1707.420 ;
        RECT 2383.905 1707.405 2384.845 1707.420 ;
        RECT 2385.545 1707.405 2385.890 1707.420 ;
        RECT 2400.490 1707.410 2401.430 1707.425 ;
        RECT 2402.130 1707.410 2402.475 1707.425 ;
        RECT 2417.075 1707.415 2418.015 1707.430 ;
        RECT 2418.715 1707.415 2419.060 1707.430 ;
        RECT 2433.655 1707.415 2434.595 1707.430 ;
        RECT 2435.295 1707.415 2435.640 1707.430 ;
        RECT 2367.320 1707.105 2369.770 1707.405 ;
        RECT 2383.905 1707.105 2386.355 1707.405 ;
        RECT 2400.490 1707.110 2402.940 1707.410 ;
        RECT 2417.075 1707.115 2419.525 1707.415 ;
        RECT 2433.655 1707.115 2436.105 1707.415 ;
        RECT 2367.320 1707.090 2369.305 1707.105 ;
        RECT 2367.320 1707.080 2368.260 1707.090 ;
        RECT 2367.320 1705.390 2367.620 1707.080 ;
        RECT 2367.920 1707.075 2368.260 1707.080 ;
        RECT 2368.960 1707.085 2369.305 1707.090 ;
        RECT 2383.905 1707.090 2385.890 1707.105 ;
        RECT 2368.960 1707.075 2369.300 1707.085 ;
        RECT 2383.905 1707.080 2384.845 1707.090 ;
        RECT 2368.280 1706.385 2368.625 1706.400 ;
        RECT 2368.280 1706.085 2369.090 1706.385 ;
        RECT 2368.280 1706.055 2368.625 1706.085 ;
        RECT 2383.905 1705.390 2384.205 1707.080 ;
        RECT 2384.505 1707.075 2384.845 1707.080 ;
        RECT 2385.545 1707.085 2385.890 1707.090 ;
        RECT 2400.490 1707.095 2402.475 1707.110 ;
        RECT 2400.490 1707.085 2401.430 1707.095 ;
        RECT 2385.545 1707.075 2385.885 1707.085 ;
        RECT 2384.865 1706.385 2385.210 1706.400 ;
        RECT 2384.865 1706.085 2385.675 1706.385 ;
        RECT 2384.865 1706.055 2385.210 1706.085 ;
        RECT 2400.490 1705.395 2400.790 1707.085 ;
        RECT 2401.090 1707.080 2401.430 1707.085 ;
        RECT 2402.130 1707.090 2402.475 1707.095 ;
        RECT 2417.075 1707.100 2419.060 1707.115 ;
        RECT 2417.075 1707.090 2418.015 1707.100 ;
        RECT 2402.130 1707.080 2402.470 1707.090 ;
        RECT 2401.450 1706.390 2401.795 1706.405 ;
        RECT 2401.450 1706.090 2402.260 1706.390 ;
        RECT 2401.450 1706.060 2401.795 1706.090 ;
        RECT 2417.075 1705.400 2417.375 1707.090 ;
        RECT 2417.675 1707.085 2418.015 1707.090 ;
        RECT 2418.715 1707.095 2419.060 1707.100 ;
        RECT 2433.655 1707.100 2435.640 1707.115 ;
        RECT 2418.715 1707.085 2419.055 1707.095 ;
        RECT 2433.655 1707.090 2434.595 1707.100 ;
        RECT 2418.035 1706.395 2418.380 1706.410 ;
        RECT 2418.035 1706.095 2418.845 1706.395 ;
        RECT 2418.035 1706.065 2418.380 1706.095 ;
        RECT 2433.655 1705.400 2433.955 1707.090 ;
        RECT 2434.255 1707.085 2434.595 1707.090 ;
        RECT 2435.295 1707.095 2435.640 1707.100 ;
        RECT 2435.295 1707.085 2435.635 1707.095 ;
        RECT 2434.615 1706.395 2434.960 1706.410 ;
        RECT 2434.615 1706.095 2435.425 1706.395 ;
        RECT 2434.615 1706.065 2434.960 1706.095 ;
        RECT 2417.075 1705.395 2419.730 1705.400 ;
        RECT 2433.655 1705.395 2436.310 1705.400 ;
        RECT 2400.490 1705.390 2403.145 1705.395 ;
        RECT 2367.320 1705.385 2369.975 1705.390 ;
        RECT 2383.905 1705.385 2386.560 1705.390 ;
        RECT 2367.320 1705.365 2369.985 1705.385 ;
        RECT 2383.905 1705.365 2386.570 1705.385 ;
        RECT 2400.490 1705.370 2403.155 1705.390 ;
        RECT 2417.075 1705.375 2419.740 1705.395 ;
        RECT 2433.655 1705.375 2436.320 1705.395 ;
        RECT 2367.320 1705.065 2370.450 1705.365 ;
        RECT 2383.905 1705.065 2387.035 1705.365 ;
        RECT 2400.490 1705.070 2403.620 1705.370 ;
        RECT 2417.075 1705.075 2420.205 1705.375 ;
        RECT 2433.655 1705.075 2436.785 1705.375 ;
        RECT 2417.075 1705.070 2419.740 1705.075 ;
        RECT 2433.655 1705.070 2436.320 1705.075 ;
        RECT 2400.490 1705.065 2403.155 1705.070 ;
        RECT 2367.320 1705.060 2369.985 1705.065 ;
        RECT 2383.905 1705.060 2386.570 1705.065 ;
        RECT 2369.640 1705.035 2369.985 1705.060 ;
        RECT 2386.225 1705.035 2386.570 1705.060 ;
        RECT 2402.810 1705.040 2403.155 1705.065 ;
        RECT 2419.395 1705.045 2419.740 1705.070 ;
        RECT 2435.975 1705.045 2436.320 1705.070 ;
        RECT 2369.660 1704.995 2369.960 1705.035 ;
        RECT 2386.245 1704.995 2386.545 1705.035 ;
        RECT 2402.830 1705.000 2403.130 1705.040 ;
        RECT 2419.415 1705.005 2419.715 1705.045 ;
        RECT 2435.995 1705.005 2436.295 1705.045 ;
        RECT 2368.950 1704.685 2369.290 1704.705 ;
        RECT 2385.535 1704.685 2385.875 1704.705 ;
        RECT 2402.120 1704.690 2402.460 1704.710 ;
        RECT 2418.705 1704.695 2419.045 1704.715 ;
        RECT 2435.285 1704.695 2435.625 1704.715 ;
        RECT 2368.480 1704.385 2369.290 1704.685 ;
        RECT 2385.065 1704.385 2385.875 1704.685 ;
        RECT 2401.650 1704.390 2402.460 1704.690 ;
        RECT 2418.235 1704.395 2419.045 1704.695 ;
        RECT 2434.815 1704.395 2435.625 1704.695 ;
        RECT 2368.950 1704.355 2369.290 1704.385 ;
        RECT 2369.650 1704.355 2369.985 1704.360 ;
        RECT 2385.535 1704.355 2385.875 1704.385 ;
        RECT 2402.120 1704.360 2402.460 1704.390 ;
        RECT 2418.705 1704.365 2419.045 1704.395 ;
        RECT 2419.405 1704.365 2419.740 1704.370 ;
        RECT 2435.285 1704.365 2435.625 1704.395 ;
        RECT 2435.985 1704.365 2436.320 1704.370 ;
        RECT 2402.820 1704.360 2403.155 1704.365 ;
        RECT 2386.235 1704.355 2386.570 1704.360 ;
        RECT 2369.640 1704.345 2369.985 1704.355 ;
        RECT 2386.225 1704.345 2386.570 1704.355 ;
        RECT 2402.810 1704.350 2403.155 1704.360 ;
        RECT 2419.395 1704.355 2419.740 1704.365 ;
        RECT 2435.975 1704.355 2436.320 1704.365 ;
        RECT 2369.640 1704.045 2370.450 1704.345 ;
        RECT 2386.225 1704.045 2387.035 1704.345 ;
        RECT 2402.810 1704.050 2403.620 1704.350 ;
        RECT 2419.395 1704.055 2420.205 1704.355 ;
        RECT 2435.975 1704.055 2436.785 1704.355 ;
        RECT 2369.640 1704.025 2369.985 1704.045 ;
        RECT 2386.225 1704.025 2386.570 1704.045 ;
        RECT 2402.810 1704.030 2403.155 1704.050 ;
        RECT 2419.395 1704.035 2419.740 1704.055 ;
        RECT 2435.975 1704.035 2436.320 1704.055 ;
        RECT 2369.640 1704.015 2369.980 1704.025 ;
        RECT 2386.225 1704.015 2386.565 1704.025 ;
        RECT 2402.810 1704.020 2403.150 1704.030 ;
        RECT 2419.395 1704.025 2419.735 1704.035 ;
        RECT 2435.975 1704.025 2436.315 1704.035 ;
        RECT 2367.600 1704.005 2367.945 1704.015 ;
        RECT 2384.185 1704.005 2384.530 1704.015 ;
        RECT 2400.770 1704.010 2401.115 1704.020 ;
        RECT 2417.355 1704.015 2417.700 1704.025 ;
        RECT 2433.935 1704.015 2434.280 1704.025 ;
        RECT 2367.140 1703.705 2367.945 1704.005 ;
        RECT 2383.725 1703.705 2384.530 1704.005 ;
        RECT 2400.310 1703.710 2401.115 1704.010 ;
        RECT 2416.895 1703.715 2417.700 1704.015 ;
        RECT 2433.475 1703.715 2434.280 1704.015 ;
        RECT 2367.500 1703.695 2367.945 1703.705 ;
        RECT 2384.085 1703.695 2384.530 1703.705 ;
        RECT 2400.670 1703.700 2401.115 1703.710 ;
        RECT 2417.255 1703.705 2417.700 1703.715 ;
        RECT 2433.835 1703.705 2434.280 1703.715 ;
        RECT 2367.600 1703.675 2367.945 1703.695 ;
        RECT 2384.185 1703.675 2384.530 1703.695 ;
        RECT 2400.770 1703.680 2401.115 1703.700 ;
        RECT 2417.355 1703.685 2417.700 1703.705 ;
        RECT 2433.935 1703.685 2434.280 1703.705 ;
        RECT 2690.000 1684.210 2694.000 1684.360 ;
        RECT 2695.125 1684.210 2695.455 1684.225 ;
        RECT 2677.265 1684.170 2677.595 1684.185 ;
        RECT 2690.000 1684.170 2695.455 1684.210 ;
        RECT 2677.265 1683.910 2695.455 1684.170 ;
        RECT 2677.265 1683.870 2694.000 1683.910 ;
        RECT 2695.125 1683.895 2695.455 1683.910 ;
        RECT 2677.265 1683.855 2677.595 1683.870 ;
        RECT 2690.000 1683.760 2694.000 1683.870 ;
        RECT 2690.000 1677.410 2694.000 1677.560 ;
        RECT 2695.585 1677.410 2695.915 1677.425 ;
        RECT 2432.750 1677.370 2433.130 1677.380 ;
        RECT 2690.000 1677.370 2695.915 1677.410 ;
        RECT 2432.750 1677.110 2695.915 1677.370 ;
        RECT 2432.750 1677.070 2694.000 1677.110 ;
        RECT 2695.585 1677.095 2695.915 1677.110 ;
        RECT 2432.750 1677.060 2433.130 1677.070 ;
        RECT 2690.000 1676.960 2694.000 1677.070 ;
        RECT 2690.000 1670.610 2694.000 1670.760 ;
        RECT 2694.665 1670.610 2694.995 1670.625 ;
        RECT 2428.150 1670.570 2428.530 1670.580 ;
        RECT 2690.000 1670.570 2694.995 1670.610 ;
        RECT 2428.150 1670.310 2694.995 1670.570 ;
        RECT 2428.150 1670.270 2694.000 1670.310 ;
        RECT 2694.665 1670.295 2694.995 1670.310 ;
        RECT 2428.150 1670.260 2428.530 1670.270 ;
        RECT 2690.000 1670.160 2694.000 1670.270 ;
        RECT 2690.000 1663.810 2694.000 1663.960 ;
        RECT 2694.665 1663.810 2694.995 1663.825 ;
        RECT 2433.670 1663.770 2434.050 1663.780 ;
        RECT 2690.000 1663.770 2694.995 1663.810 ;
        RECT 2433.670 1663.510 2694.995 1663.770 ;
        RECT 2433.670 1663.470 2694.000 1663.510 ;
        RECT 2694.665 1663.495 2694.995 1663.510 ;
        RECT 2433.670 1663.460 2434.050 1663.470 ;
        RECT 2690.000 1663.360 2694.000 1663.470 ;
        RECT 2690.000 1657.010 2694.000 1657.160 ;
        RECT 2694.665 1657.010 2694.995 1657.025 ;
        RECT 2677.265 1656.970 2677.595 1656.985 ;
        RECT 2690.000 1656.970 2694.995 1657.010 ;
        RECT 2677.265 1656.710 2694.995 1656.970 ;
        RECT 2677.265 1656.670 2694.000 1656.710 ;
        RECT 2694.665 1656.695 2694.995 1656.710 ;
        RECT 2677.265 1656.655 2677.595 1656.670 ;
        RECT 2690.000 1656.560 2694.000 1656.670 ;
        RECT 2690.000 1650.210 2694.000 1650.360 ;
        RECT 2694.665 1650.210 2694.995 1650.225 ;
        RECT 2677.265 1650.170 2677.595 1650.185 ;
        RECT 2690.000 1650.170 2694.995 1650.210 ;
        RECT 2677.265 1649.910 2694.995 1650.170 ;
        RECT 2677.265 1649.870 2694.000 1649.910 ;
        RECT 2694.665 1649.895 2694.995 1649.910 ;
        RECT 2677.265 1649.855 2677.595 1649.870 ;
        RECT 2690.000 1649.760 2694.000 1649.870 ;
        RECT 2690.000 1643.410 2694.000 1643.560 ;
        RECT 2694.665 1643.410 2694.995 1643.425 ;
        RECT 2680.025 1643.370 2680.355 1643.385 ;
        RECT 2690.000 1643.370 2694.995 1643.410 ;
        RECT 2680.025 1643.110 2694.995 1643.370 ;
        RECT 2680.025 1643.070 2694.000 1643.110 ;
        RECT 2694.665 1643.095 2694.995 1643.110 ;
        RECT 2680.025 1643.055 2680.355 1643.070 ;
        RECT 2690.000 1642.960 2694.000 1643.070 ;
        RECT 2690.000 1636.610 2694.000 1636.760 ;
        RECT 2694.665 1636.610 2694.995 1636.625 ;
        RECT 2683.245 1636.570 2683.575 1636.585 ;
        RECT 2690.000 1636.570 2694.995 1636.610 ;
        RECT 2683.245 1636.310 2694.995 1636.570 ;
        RECT 2683.245 1636.270 2694.000 1636.310 ;
        RECT 2694.665 1636.295 2694.995 1636.310 ;
        RECT 2683.245 1636.255 2683.575 1636.270 ;
        RECT 2690.000 1636.160 2694.000 1636.270 ;
        RECT 2690.000 1629.810 2694.000 1629.960 ;
        RECT 2694.665 1629.810 2694.995 1629.825 ;
        RECT 2677.265 1629.770 2677.595 1629.785 ;
        RECT 2690.000 1629.770 2694.995 1629.810 ;
        RECT 2677.265 1629.510 2694.995 1629.770 ;
        RECT 2677.265 1629.470 2694.000 1629.510 ;
        RECT 2694.665 1629.495 2694.995 1629.510 ;
        RECT 2677.265 1629.455 2677.595 1629.470 ;
        RECT 2690.000 1629.360 2694.000 1629.470 ;
        RECT 2523.535 1624.615 2678.820 1624.945 ;
        RECT 2523.535 1618.200 2674.980 1618.530 ;
        RECT 2674.650 1609.805 2674.980 1618.200 ;
        RECT 2678.490 1616.455 2678.820 1624.615 ;
        RECT 2690.000 1623.010 2694.000 1623.160 ;
        RECT 2694.665 1623.010 2694.995 1623.025 ;
        RECT 2681.865 1622.970 2682.195 1622.985 ;
        RECT 2690.000 1622.970 2694.995 1623.010 ;
        RECT 2681.865 1622.710 2694.995 1622.970 ;
        RECT 2681.865 1622.670 2694.000 1622.710 ;
        RECT 2694.665 1622.695 2694.995 1622.710 ;
        RECT 2681.865 1622.655 2682.195 1622.670 ;
        RECT 2690.000 1622.560 2694.000 1622.670 ;
        RECT 2678.490 1616.360 2690.625 1616.455 ;
        RECT 2678.490 1616.210 2694.000 1616.360 ;
        RECT 2694.665 1616.210 2694.995 1616.225 ;
        RECT 2678.490 1616.125 2694.995 1616.210 ;
        RECT 2690.000 1615.910 2694.995 1616.125 ;
        RECT 2690.000 1615.760 2694.000 1615.910 ;
        RECT 2694.665 1615.895 2694.995 1615.910 ;
        RECT 2362.915 1609.620 2363.285 1609.690 ;
        RECT 2380.135 1609.620 2380.505 1609.690 ;
        RECT 2397.355 1609.625 2397.725 1609.695 ;
        RECT 2362.915 1609.320 2370.065 1609.620 ;
        RECT 2380.135 1609.320 2387.285 1609.620 ;
        RECT 2397.355 1609.325 2404.505 1609.625 ;
        RECT 2367.680 1608.090 2367.980 1609.320 ;
        RECT 2367.180 1607.790 2367.980 1608.090 ;
        RECT 2367.560 1607.745 2367.980 1607.790 ;
        RECT 2368.710 1608.100 2369.015 1609.320 ;
        RECT 2367.560 1607.720 2367.860 1607.745 ;
        RECT 2368.710 1607.430 2369.010 1608.100 ;
        RECT 2369.765 1607.465 2370.065 1609.320 ;
        RECT 2384.900 1608.090 2385.200 1609.320 ;
        RECT 2384.400 1607.790 2385.200 1608.090 ;
        RECT 2384.780 1607.745 2385.200 1607.790 ;
        RECT 2385.930 1608.100 2386.235 1609.320 ;
        RECT 2384.780 1607.720 2385.080 1607.745 ;
        RECT 2368.670 1607.415 2369.010 1607.430 ;
        RECT 2368.660 1607.400 2369.010 1607.415 ;
        RECT 2368.190 1607.100 2369.010 1607.400 ;
        RECT 2369.690 1607.400 2370.065 1607.465 ;
        RECT 2385.930 1607.430 2386.230 1608.100 ;
        RECT 2386.985 1607.465 2387.285 1609.320 ;
        RECT 2402.120 1608.095 2402.420 1609.325 ;
        RECT 2401.620 1607.795 2402.420 1608.095 ;
        RECT 2402.000 1607.750 2402.420 1607.795 ;
        RECT 2403.150 1608.105 2403.455 1609.325 ;
        RECT 2402.000 1607.725 2402.300 1607.750 ;
        RECT 2385.890 1607.415 2386.230 1607.430 ;
        RECT 2385.880 1607.400 2386.230 1607.415 ;
        RECT 2369.690 1607.100 2370.500 1607.400 ;
        RECT 2385.410 1607.100 2386.230 1607.400 ;
        RECT 2386.910 1607.400 2387.285 1607.465 ;
        RECT 2403.150 1607.435 2403.450 1608.105 ;
        RECT 2404.205 1607.470 2404.505 1609.325 ;
        RECT 2414.575 1609.620 2414.945 1609.690 ;
        RECT 2431.795 1609.620 2432.165 1609.690 ;
        RECT 2414.575 1609.320 2421.725 1609.620 ;
        RECT 2431.795 1609.320 2438.945 1609.620 ;
        RECT 2674.650 1609.560 2691.175 1609.805 ;
        RECT 2674.650 1609.475 2694.000 1609.560 ;
        RECT 2419.340 1608.090 2419.640 1609.320 ;
        RECT 2418.840 1607.790 2419.640 1608.090 ;
        RECT 2419.220 1607.745 2419.640 1607.790 ;
        RECT 2420.370 1608.100 2420.675 1609.320 ;
        RECT 2419.220 1607.720 2419.520 1607.745 ;
        RECT 2403.110 1607.420 2403.450 1607.435 ;
        RECT 2403.100 1607.405 2403.450 1607.420 ;
        RECT 2386.910 1607.100 2387.720 1607.400 ;
        RECT 2402.630 1607.105 2403.450 1607.405 ;
        RECT 2404.130 1607.405 2404.505 1607.470 ;
        RECT 2420.370 1607.430 2420.670 1608.100 ;
        RECT 2421.425 1607.465 2421.725 1609.320 ;
        RECT 2436.560 1608.090 2436.860 1609.320 ;
        RECT 2436.060 1607.790 2436.860 1608.090 ;
        RECT 2436.440 1607.745 2436.860 1607.790 ;
        RECT 2437.590 1608.100 2437.895 1609.320 ;
        RECT 2436.440 1607.720 2436.740 1607.745 ;
        RECT 2420.330 1607.415 2420.670 1607.430 ;
        RECT 2404.130 1607.105 2404.940 1607.405 ;
        RECT 2420.320 1607.400 2420.670 1607.415 ;
        RECT 2368.660 1607.085 2369.010 1607.100 ;
        RECT 2369.700 1607.085 2370.055 1607.100 ;
        RECT 2385.880 1607.085 2386.230 1607.100 ;
        RECT 2386.920 1607.085 2387.275 1607.100 ;
        RECT 2403.100 1607.090 2403.450 1607.105 ;
        RECT 2404.140 1607.090 2404.495 1607.105 ;
        RECT 2419.850 1607.100 2420.670 1607.400 ;
        RECT 2421.350 1607.400 2421.725 1607.465 ;
        RECT 2437.590 1607.430 2437.890 1608.100 ;
        RECT 2438.645 1607.465 2438.945 1609.320 ;
        RECT 2690.000 1609.410 2694.000 1609.475 ;
        RECT 2694.665 1609.410 2694.995 1609.425 ;
        RECT 2690.000 1609.110 2694.995 1609.410 ;
        RECT 2690.000 1608.960 2694.000 1609.110 ;
        RECT 2694.665 1609.095 2694.995 1609.110 ;
        RECT 2437.550 1607.415 2437.890 1607.430 ;
        RECT 2437.540 1607.400 2437.890 1607.415 ;
        RECT 2421.350 1607.100 2422.160 1607.400 ;
        RECT 2437.070 1607.100 2437.890 1607.400 ;
        RECT 2438.570 1607.400 2438.945 1607.465 ;
        RECT 2438.570 1607.100 2439.380 1607.400 ;
        RECT 2403.110 1607.085 2403.450 1607.090 ;
        RECT 2368.670 1607.080 2369.010 1607.085 ;
        RECT 2368.685 1607.040 2368.985 1607.080 ;
        RECT 2369.755 1607.060 2370.055 1607.085 ;
        RECT 2385.890 1607.080 2386.230 1607.085 ;
        RECT 2385.905 1607.040 2386.205 1607.080 ;
        RECT 2386.975 1607.060 2387.275 1607.085 ;
        RECT 2403.125 1607.045 2403.425 1607.085 ;
        RECT 2404.195 1607.065 2404.495 1607.090 ;
        RECT 2420.320 1607.085 2420.670 1607.100 ;
        RECT 2421.360 1607.085 2421.715 1607.100 ;
        RECT 2437.540 1607.085 2437.890 1607.100 ;
        RECT 2438.580 1607.085 2438.935 1607.100 ;
        RECT 2420.330 1607.080 2420.670 1607.085 ;
        RECT 2420.345 1607.040 2420.645 1607.080 ;
        RECT 2421.415 1607.060 2421.715 1607.085 ;
        RECT 2437.550 1607.080 2437.890 1607.085 ;
        RECT 2437.565 1607.040 2437.865 1607.080 ;
        RECT 2438.635 1607.060 2438.935 1607.085 ;
        RECT 2366.290 1605.765 2366.620 1605.780 ;
        RECT 2368.330 1605.765 2368.660 1605.780 ;
        RECT 2366.290 1605.465 2368.660 1605.765 ;
        RECT 2366.290 1605.450 2366.620 1605.465 ;
        RECT 2368.330 1605.450 2368.660 1605.465 ;
        RECT 2383.510 1605.765 2383.840 1605.780 ;
        RECT 2385.550 1605.765 2385.880 1605.780 ;
        RECT 2383.510 1605.465 2385.880 1605.765 ;
        RECT 2383.510 1605.450 2383.840 1605.465 ;
        RECT 2385.550 1605.450 2385.880 1605.465 ;
        RECT 2400.730 1605.770 2401.060 1605.785 ;
        RECT 2402.770 1605.770 2403.100 1605.785 ;
        RECT 2400.730 1605.470 2403.100 1605.770 ;
        RECT 2400.730 1605.455 2401.060 1605.470 ;
        RECT 2402.770 1605.455 2403.100 1605.470 ;
        RECT 2417.950 1605.765 2418.280 1605.780 ;
        RECT 2419.990 1605.765 2420.320 1605.780 ;
        RECT 2417.950 1605.465 2420.320 1605.765 ;
        RECT 2417.950 1605.450 2418.280 1605.465 ;
        RECT 2419.990 1605.450 2420.320 1605.465 ;
        RECT 2435.170 1605.765 2435.500 1605.780 ;
        RECT 2437.210 1605.765 2437.540 1605.780 ;
        RECT 2435.170 1605.465 2437.540 1605.765 ;
        RECT 2435.170 1605.450 2435.500 1605.465 ;
        RECT 2437.210 1605.450 2437.540 1605.465 ;
        RECT 2369.350 1605.365 2369.680 1605.380 ;
        RECT 2386.570 1605.365 2386.900 1605.380 ;
        RECT 2403.790 1605.370 2404.120 1605.385 ;
        RECT 2369.350 1605.065 2370.150 1605.365 ;
        RECT 2386.570 1605.065 2387.370 1605.365 ;
        RECT 2403.790 1605.070 2404.590 1605.370 ;
        RECT 2421.010 1605.365 2421.340 1605.380 ;
        RECT 2438.230 1605.365 2438.560 1605.380 ;
        RECT 2369.350 1605.050 2369.680 1605.065 ;
        RECT 2386.570 1605.050 2386.900 1605.065 ;
        RECT 2403.790 1605.055 2404.120 1605.070 ;
        RECT 2421.010 1605.065 2421.810 1605.365 ;
        RECT 2438.230 1605.065 2439.030 1605.365 ;
        RECT 2367.980 1605.025 2368.310 1605.040 ;
        RECT 2367.520 1604.725 2368.320 1605.025 ;
        RECT 2369.365 1605.020 2369.665 1605.050 ;
        RECT 2385.200 1605.025 2385.530 1605.040 ;
        RECT 2384.740 1604.725 2385.540 1605.025 ;
        RECT 2386.585 1605.020 2386.885 1605.050 ;
        RECT 2402.420 1605.030 2402.750 1605.045 ;
        RECT 2401.960 1604.730 2402.760 1605.030 ;
        RECT 2403.805 1605.025 2404.105 1605.055 ;
        RECT 2421.010 1605.050 2421.340 1605.065 ;
        RECT 2438.230 1605.050 2438.560 1605.065 ;
        RECT 2419.640 1605.025 2419.970 1605.040 ;
        RECT 2367.980 1604.710 2368.310 1604.725 ;
        RECT 2385.200 1604.710 2385.530 1604.725 ;
        RECT 2402.420 1604.715 2402.750 1604.730 ;
        RECT 2419.180 1604.725 2419.980 1605.025 ;
        RECT 2421.025 1605.020 2421.325 1605.050 ;
        RECT 2436.860 1605.025 2437.190 1605.040 ;
        RECT 2436.400 1604.725 2437.200 1605.025 ;
        RECT 2438.245 1605.020 2438.545 1605.050 ;
        RECT 2419.640 1604.710 2419.970 1604.725 ;
        RECT 2436.860 1604.710 2437.190 1604.725 ;
        RECT 2369.010 1604.685 2369.340 1604.700 ;
        RECT 2386.230 1604.685 2386.560 1604.700 ;
        RECT 2403.450 1604.690 2403.780 1604.705 ;
        RECT 2369.010 1604.385 2369.810 1604.685 ;
        RECT 2386.230 1604.385 2387.030 1604.685 ;
        RECT 2403.450 1604.390 2404.250 1604.690 ;
        RECT 2420.670 1604.685 2421.000 1604.700 ;
        RECT 2437.890 1604.685 2438.220 1604.700 ;
        RECT 2369.010 1604.370 2369.395 1604.385 ;
        RECT 2386.230 1604.370 2386.615 1604.385 ;
        RECT 2403.450 1604.375 2403.835 1604.390 ;
        RECT 2369.095 1604.360 2369.395 1604.370 ;
        RECT 2386.315 1604.360 2386.615 1604.370 ;
        RECT 2403.535 1604.365 2403.835 1604.375 ;
        RECT 2420.670 1604.385 2421.470 1604.685 ;
        RECT 2437.890 1604.385 2438.690 1604.685 ;
        RECT 2420.670 1604.370 2421.055 1604.385 ;
        RECT 2437.890 1604.370 2438.275 1604.385 ;
        RECT 2420.755 1604.360 2421.055 1604.370 ;
        RECT 2437.975 1604.360 2438.275 1604.370 ;
        RECT 2367.650 1603.835 2367.980 1603.850 ;
        RECT 2384.870 1603.835 2385.200 1603.850 ;
        RECT 2402.090 1603.840 2402.420 1603.855 ;
        RECT 2367.180 1603.535 2367.980 1603.835 ;
        RECT 2384.400 1603.535 2385.200 1603.835 ;
        RECT 2401.620 1603.540 2402.420 1603.840 ;
        RECT 2419.310 1603.835 2419.640 1603.850 ;
        RECT 2436.530 1603.835 2436.860 1603.850 ;
        RECT 2402.080 1603.535 2402.420 1603.540 ;
        RECT 2418.840 1603.535 2419.640 1603.835 ;
        RECT 2436.060 1603.535 2436.860 1603.835 ;
        RECT 2367.640 1603.530 2367.980 1603.535 ;
        RECT 2384.860 1603.530 2385.200 1603.535 ;
        RECT 2367.650 1603.520 2367.980 1603.530 ;
        RECT 2384.870 1603.520 2385.200 1603.530 ;
        RECT 2402.090 1603.525 2402.420 1603.535 ;
        RECT 2419.300 1603.530 2419.640 1603.535 ;
        RECT 2436.520 1603.530 2436.860 1603.535 ;
        RECT 2419.310 1603.520 2419.640 1603.530 ;
        RECT 2436.530 1603.520 2436.860 1603.530 ;
        RECT 2690.000 1602.610 2694.000 1602.760 ;
        RECT 2694.665 1602.610 2694.995 1602.625 ;
        RECT 2690.000 1602.320 2694.995 1602.610 ;
        RECT 2666.230 1602.310 2694.995 1602.320 ;
        RECT 2666.230 1602.160 2694.000 1602.310 ;
        RECT 2694.665 1602.295 2694.995 1602.310 ;
        RECT 2666.230 1601.990 2690.795 1602.160 ;
        RECT 2666.230 1589.285 2666.560 1601.990 ;
        RECT 2523.535 1588.955 2666.560 1589.285 ;
        RECT 2670.115 1595.960 2690.640 1595.980 ;
        RECT 2670.115 1595.810 2694.000 1595.960 ;
        RECT 2694.665 1595.810 2694.995 1595.825 ;
        RECT 2670.115 1595.650 2694.995 1595.810 ;
        RECT 2670.115 1581.755 2670.445 1595.650 ;
        RECT 2690.000 1595.510 2694.995 1595.650 ;
        RECT 2690.000 1595.360 2694.000 1595.510 ;
        RECT 2694.665 1595.495 2694.995 1595.510 ;
        RECT 2690.000 1589.010 2694.000 1589.160 ;
        RECT 2694.665 1589.010 2694.995 1589.025 ;
        RECT 2690.000 1588.845 2694.995 1589.010 ;
        RECT 2523.535 1581.425 2670.445 1581.755 ;
        RECT 2672.900 1588.710 2694.995 1588.845 ;
        RECT 2672.900 1588.560 2694.000 1588.710 ;
        RECT 2694.665 1588.695 2694.995 1588.710 ;
        RECT 2672.900 1588.515 2691.165 1588.560 ;
        RECT 2672.900 1575.775 2673.230 1588.515 ;
        RECT 2698.345 1582.890 2698.675 1582.905 ;
        RECT 2694.910 1582.590 2698.675 1582.890 ;
        RECT 2690.000 1582.225 2694.000 1582.360 ;
        RECT 2523.535 1575.445 2673.230 1575.775 ;
        RECT 2678.125 1582.210 2694.000 1582.225 ;
        RECT 2694.910 1582.210 2695.210 1582.590 ;
        RECT 2698.345 1582.575 2698.675 1582.590 ;
        RECT 2678.125 1581.910 2695.210 1582.210 ;
        RECT 2678.125 1581.895 2694.000 1581.910 ;
        RECT 2678.125 1567.360 2678.455 1581.895 ;
        RECT 2690.000 1581.760 2694.000 1581.895 ;
        RECT 2523.535 1567.030 2678.455 1567.360 ;
        RECT 2368.100 1532.675 2368.470 1532.710 ;
        RECT 2384.425 1532.675 2384.795 1532.710 ;
        RECT 2400.750 1532.675 2401.120 1532.710 ;
        RECT 2417.075 1532.675 2417.445 1532.710 ;
        RECT 2433.400 1532.675 2433.770 1532.710 ;
        RECT 2368.100 1532.375 2370.085 1532.675 ;
        RECT 2368.100 1532.340 2368.470 1532.375 ;
        RECT 2366.400 1528.035 2366.735 1528.055 ;
        RECT 2365.195 1527.735 2366.735 1528.035 ;
        RECT 2361.780 1526.755 2362.115 1527.490 ;
        RECT 2364.225 1526.930 2364.555 1527.325 ;
        RECT 2365.195 1526.930 2365.495 1527.735 ;
        RECT 2366.400 1527.715 2366.735 1527.735 ;
        RECT 2368.340 1527.165 2368.675 1527.490 ;
        RECT 2363.225 1526.360 2363.555 1526.765 ;
        RECT 2364.220 1526.595 2364.555 1526.930 ;
        RECT 2364.940 1526.615 2365.495 1526.930 ;
        RECT 2365.900 1526.875 2366.235 1526.930 ;
        RECT 2366.780 1526.875 2367.115 1526.930 ;
        RECT 2364.940 1526.595 2365.275 1526.615 ;
        RECT 2365.900 1526.600 2368.045 1526.875 ;
        RECT 2368.345 1526.755 2368.675 1527.165 ;
        RECT 2369.785 1526.875 2370.085 1532.375 ;
        RECT 2384.425 1532.375 2386.410 1532.675 ;
        RECT 2384.425 1532.340 2384.795 1532.375 ;
        RECT 2382.725 1528.035 2383.060 1528.055 ;
        RECT 2381.520 1527.735 2383.060 1528.035 ;
        RECT 2363.220 1526.035 2363.555 1526.360 ;
        RECT 2365.905 1526.575 2368.045 1526.600 ;
        RECT 2365.905 1526.195 2366.235 1526.575 ;
        RECT 2366.785 1526.195 2367.115 1526.575 ;
        RECT 2367.745 1526.455 2368.045 1526.575 ;
        RECT 2368.985 1526.575 2370.275 1526.875 ;
        RECT 2378.105 1526.755 2378.440 1527.490 ;
        RECT 2380.550 1526.930 2380.880 1527.325 ;
        RECT 2381.520 1526.930 2381.820 1527.735 ;
        RECT 2382.725 1527.715 2383.060 1527.735 ;
        RECT 2384.665 1527.165 2385.000 1527.490 ;
        RECT 2368.985 1526.455 2369.290 1526.575 ;
        RECT 2367.745 1526.155 2369.290 1526.455 ;
        RECT 2369.940 1526.415 2370.275 1526.575 ;
        RECT 2369.945 1526.035 2370.275 1526.415 ;
        RECT 2379.550 1526.360 2379.880 1526.765 ;
        RECT 2380.545 1526.595 2380.880 1526.930 ;
        RECT 2381.265 1526.615 2381.820 1526.930 ;
        RECT 2382.225 1526.875 2382.560 1526.930 ;
        RECT 2383.105 1526.875 2383.440 1526.930 ;
        RECT 2381.265 1526.595 2381.600 1526.615 ;
        RECT 2382.225 1526.600 2384.370 1526.875 ;
        RECT 2384.670 1526.755 2385.000 1527.165 ;
        RECT 2386.110 1526.875 2386.410 1532.375 ;
        RECT 2400.750 1532.375 2402.735 1532.675 ;
        RECT 2400.750 1532.340 2401.120 1532.375 ;
        RECT 2399.050 1528.035 2399.385 1528.055 ;
        RECT 2397.845 1527.735 2399.385 1528.035 ;
        RECT 2379.545 1526.035 2379.880 1526.360 ;
        RECT 2382.230 1526.575 2384.370 1526.600 ;
        RECT 2382.230 1526.195 2382.560 1526.575 ;
        RECT 2383.110 1526.195 2383.440 1526.575 ;
        RECT 2384.070 1526.455 2384.370 1526.575 ;
        RECT 2385.310 1526.575 2386.600 1526.875 ;
        RECT 2394.430 1526.755 2394.765 1527.490 ;
        RECT 2396.875 1526.930 2397.205 1527.325 ;
        RECT 2397.845 1526.930 2398.145 1527.735 ;
        RECT 2399.050 1527.715 2399.385 1527.735 ;
        RECT 2400.990 1527.165 2401.325 1527.490 ;
        RECT 2385.310 1526.455 2385.615 1526.575 ;
        RECT 2384.070 1526.155 2385.615 1526.455 ;
        RECT 2386.265 1526.415 2386.600 1526.575 ;
        RECT 2386.270 1526.035 2386.600 1526.415 ;
        RECT 2395.875 1526.360 2396.205 1526.765 ;
        RECT 2396.870 1526.595 2397.205 1526.930 ;
        RECT 2397.590 1526.615 2398.145 1526.930 ;
        RECT 2398.550 1526.875 2398.885 1526.930 ;
        RECT 2399.430 1526.875 2399.765 1526.930 ;
        RECT 2397.590 1526.595 2397.925 1526.615 ;
        RECT 2398.550 1526.600 2400.695 1526.875 ;
        RECT 2400.995 1526.755 2401.325 1527.165 ;
        RECT 2402.435 1526.875 2402.735 1532.375 ;
        RECT 2417.075 1532.375 2419.060 1532.675 ;
        RECT 2417.075 1532.340 2417.445 1532.375 ;
        RECT 2415.375 1528.035 2415.710 1528.055 ;
        RECT 2414.170 1527.735 2415.710 1528.035 ;
        RECT 2395.870 1526.035 2396.205 1526.360 ;
        RECT 2398.555 1526.575 2400.695 1526.600 ;
        RECT 2398.555 1526.195 2398.885 1526.575 ;
        RECT 2399.435 1526.195 2399.765 1526.575 ;
        RECT 2400.395 1526.455 2400.695 1526.575 ;
        RECT 2401.635 1526.575 2402.925 1526.875 ;
        RECT 2410.755 1526.755 2411.090 1527.490 ;
        RECT 2413.200 1526.930 2413.530 1527.325 ;
        RECT 2414.170 1526.930 2414.470 1527.735 ;
        RECT 2415.375 1527.715 2415.710 1527.735 ;
        RECT 2417.315 1527.165 2417.650 1527.490 ;
        RECT 2401.635 1526.455 2401.940 1526.575 ;
        RECT 2400.395 1526.155 2401.940 1526.455 ;
        RECT 2402.590 1526.415 2402.925 1526.575 ;
        RECT 2402.595 1526.035 2402.925 1526.415 ;
        RECT 2412.200 1526.360 2412.530 1526.765 ;
        RECT 2413.195 1526.595 2413.530 1526.930 ;
        RECT 2413.915 1526.615 2414.470 1526.930 ;
        RECT 2414.875 1526.875 2415.210 1526.930 ;
        RECT 2415.755 1526.875 2416.090 1526.930 ;
        RECT 2413.915 1526.595 2414.250 1526.615 ;
        RECT 2414.875 1526.600 2417.020 1526.875 ;
        RECT 2417.320 1526.755 2417.650 1527.165 ;
        RECT 2418.760 1526.875 2419.060 1532.375 ;
        RECT 2433.400 1532.375 2435.385 1532.675 ;
        RECT 2433.400 1532.340 2433.770 1532.375 ;
        RECT 2431.700 1528.035 2432.035 1528.055 ;
        RECT 2430.495 1527.735 2432.035 1528.035 ;
        RECT 2412.195 1526.035 2412.530 1526.360 ;
        RECT 2414.880 1526.575 2417.020 1526.600 ;
        RECT 2414.880 1526.195 2415.210 1526.575 ;
        RECT 2415.760 1526.195 2416.090 1526.575 ;
        RECT 2416.720 1526.455 2417.020 1526.575 ;
        RECT 2417.960 1526.575 2419.250 1526.875 ;
        RECT 2427.080 1526.755 2427.415 1527.490 ;
        RECT 2429.525 1526.930 2429.855 1527.325 ;
        RECT 2430.495 1526.930 2430.795 1527.735 ;
        RECT 2431.700 1527.715 2432.035 1527.735 ;
        RECT 2433.640 1527.165 2433.975 1527.490 ;
        RECT 2417.960 1526.455 2418.265 1526.575 ;
        RECT 2416.720 1526.155 2418.265 1526.455 ;
        RECT 2418.915 1526.415 2419.250 1526.575 ;
        RECT 2418.920 1526.035 2419.250 1526.415 ;
        RECT 2428.525 1526.360 2428.855 1526.765 ;
        RECT 2429.520 1526.595 2429.855 1526.930 ;
        RECT 2430.240 1526.615 2430.795 1526.930 ;
        RECT 2431.200 1526.875 2431.535 1526.930 ;
        RECT 2432.080 1526.875 2432.415 1526.930 ;
        RECT 2430.240 1526.595 2430.575 1526.615 ;
        RECT 2431.200 1526.600 2433.345 1526.875 ;
        RECT 2433.645 1526.755 2433.975 1527.165 ;
        RECT 2435.085 1526.875 2435.385 1532.375 ;
        RECT 2428.520 1526.035 2428.855 1526.360 ;
        RECT 2431.205 1526.575 2433.345 1526.600 ;
        RECT 2431.205 1526.195 2431.535 1526.575 ;
        RECT 2432.085 1526.195 2432.415 1526.575 ;
        RECT 2433.045 1526.455 2433.345 1526.575 ;
        RECT 2434.285 1526.575 2435.575 1526.875 ;
        RECT 2434.285 1526.455 2434.590 1526.575 ;
        RECT 2433.045 1526.155 2434.590 1526.455 ;
        RECT 2435.240 1526.415 2435.575 1526.575 ;
        RECT 2435.245 1526.035 2435.575 1526.415 ;
        RECT 2690.000 1504.210 2694.000 1504.360 ;
        RECT 2695.125 1504.210 2695.455 1504.225 ;
        RECT 2677.265 1503.970 2677.595 1503.985 ;
        RECT 2690.000 1503.970 2695.455 1504.210 ;
        RECT 2677.265 1503.910 2695.455 1503.970 ;
        RECT 2677.265 1503.760 2694.000 1503.910 ;
        RECT 2695.125 1503.895 2695.455 1503.910 ;
        RECT 2677.265 1503.670 2690.540 1503.760 ;
        RECT 2677.265 1503.655 2677.595 1503.670 ;
        RECT 2690.000 1497.410 2694.000 1497.560 ;
        RECT 2695.585 1497.410 2695.915 1497.425 ;
        RECT 2677.265 1497.170 2677.595 1497.185 ;
        RECT 2690.000 1497.170 2695.915 1497.410 ;
        RECT 2677.265 1497.110 2695.915 1497.170 ;
        RECT 2677.265 1496.960 2694.000 1497.110 ;
        RECT 2695.585 1497.095 2695.915 1497.110 ;
        RECT 2677.265 1496.870 2690.540 1496.960 ;
        RECT 2677.265 1496.855 2677.595 1496.870 ;
        RECT 2690.000 1490.610 2694.000 1490.760 ;
        RECT 2694.665 1490.610 2694.995 1490.625 ;
        RECT 2677.265 1490.370 2677.595 1490.385 ;
        RECT 2690.000 1490.370 2694.995 1490.610 ;
        RECT 2677.265 1490.310 2694.995 1490.370 ;
        RECT 2677.265 1490.160 2694.000 1490.310 ;
        RECT 2694.665 1490.295 2694.995 1490.310 ;
        RECT 2677.265 1490.070 2690.540 1490.160 ;
        RECT 2677.265 1490.055 2677.595 1490.070 ;
        RECT 2690.000 1483.810 2694.000 1483.960 ;
        RECT 2694.665 1483.810 2694.995 1483.825 ;
        RECT 2677.265 1483.570 2677.595 1483.585 ;
        RECT 2690.000 1483.570 2694.995 1483.810 ;
        RECT 2677.265 1483.510 2694.995 1483.570 ;
        RECT 2677.265 1483.360 2694.000 1483.510 ;
        RECT 2694.665 1483.495 2694.995 1483.510 ;
        RECT 2677.265 1483.270 2690.540 1483.360 ;
        RECT 2677.265 1483.255 2677.595 1483.270 ;
        RECT 2690.000 1477.010 2694.000 1477.160 ;
        RECT 2694.665 1477.010 2694.995 1477.025 ;
        RECT 2677.725 1476.770 2678.055 1476.785 ;
        RECT 2690.000 1476.770 2694.995 1477.010 ;
        RECT 2677.725 1476.710 2694.995 1476.770 ;
        RECT 2677.725 1476.560 2694.000 1476.710 ;
        RECT 2694.665 1476.695 2694.995 1476.710 ;
        RECT 2677.725 1476.470 2690.540 1476.560 ;
        RECT 2677.725 1476.455 2678.055 1476.470 ;
        RECT 2690.000 1470.210 2694.000 1470.360 ;
        RECT 2694.665 1470.210 2694.995 1470.225 ;
        RECT 2677.265 1469.970 2677.595 1469.985 ;
        RECT 2690.000 1469.970 2694.995 1470.210 ;
        RECT 2677.265 1469.910 2694.995 1469.970 ;
        RECT 2677.265 1469.760 2694.000 1469.910 ;
        RECT 2694.665 1469.895 2694.995 1469.910 ;
        RECT 2677.265 1469.670 2690.540 1469.760 ;
        RECT 2677.265 1469.655 2677.595 1469.670 ;
        RECT 2690.000 1463.410 2694.000 1463.560 ;
        RECT 2694.665 1463.410 2694.995 1463.425 ;
        RECT 2677.725 1463.170 2678.055 1463.185 ;
        RECT 2690.000 1463.170 2694.995 1463.410 ;
        RECT 2677.725 1463.110 2694.995 1463.170 ;
        RECT 2677.725 1462.960 2694.000 1463.110 ;
        RECT 2694.665 1463.095 2694.995 1463.110 ;
        RECT 2677.725 1462.870 2690.540 1462.960 ;
        RECT 2677.725 1462.855 2678.055 1462.870 ;
        RECT 2690.000 1456.610 2694.000 1456.760 ;
        RECT 2694.665 1456.610 2694.995 1456.625 ;
        RECT 2677.265 1456.370 2677.595 1456.385 ;
        RECT 2690.000 1456.370 2694.995 1456.610 ;
        RECT 2677.265 1456.310 2694.995 1456.370 ;
        RECT 2677.265 1456.160 2694.000 1456.310 ;
        RECT 2694.665 1456.295 2694.995 1456.310 ;
        RECT 2677.265 1456.070 2690.540 1456.160 ;
        RECT 2677.265 1456.055 2677.595 1456.070 ;
        RECT 2690.000 1449.810 2694.000 1449.960 ;
        RECT 2694.665 1449.810 2694.995 1449.825 ;
        RECT 2677.265 1449.570 2677.595 1449.585 ;
        RECT 2690.000 1449.570 2694.995 1449.810 ;
        RECT 2677.265 1449.510 2694.995 1449.570 ;
        RECT 2677.265 1449.360 2694.000 1449.510 ;
        RECT 2694.665 1449.495 2694.995 1449.510 ;
        RECT 2677.265 1449.270 2690.540 1449.360 ;
        RECT 2677.265 1449.255 2677.595 1449.270 ;
        RECT 2690.000 1443.010 2694.000 1443.160 ;
        RECT 2694.665 1443.010 2694.995 1443.025 ;
        RECT 2677.265 1442.770 2677.595 1442.785 ;
        RECT 2690.000 1442.770 2694.995 1443.010 ;
        RECT 2677.265 1442.710 2694.995 1442.770 ;
        RECT 2677.265 1442.560 2694.000 1442.710 ;
        RECT 2694.665 1442.695 2694.995 1442.710 ;
        RECT 2677.265 1442.470 2690.540 1442.560 ;
        RECT 2677.265 1442.455 2677.595 1442.470 ;
        RECT 2523.535 1437.330 2690.720 1437.660 ;
        RECT 2690.390 1436.360 2690.720 1437.330 ;
        RECT 2690.000 1436.210 2694.000 1436.360 ;
        RECT 2694.665 1436.210 2694.995 1436.225 ;
        RECT 2690.000 1435.910 2694.995 1436.210 ;
        RECT 2690.000 1435.760 2694.000 1435.910 ;
        RECT 2694.665 1435.895 2694.995 1435.910 ;
        RECT 2370.315 1434.685 2370.690 1434.715 ;
        RECT 2388.875 1434.685 2389.250 1434.715 ;
        RECT 2407.435 1434.685 2407.810 1434.715 ;
        RECT 2425.995 1434.685 2426.370 1434.715 ;
        RECT 2444.555 1434.685 2444.930 1434.715 ;
        RECT 2370.315 1434.385 2371.320 1434.685 ;
        RECT 2370.315 1434.345 2370.690 1434.385 ;
        RECT 2371.020 1431.995 2371.320 1434.385 ;
        RECT 2388.875 1434.385 2389.880 1434.685 ;
        RECT 2388.875 1434.345 2389.250 1434.385 ;
        RECT 2389.580 1431.995 2389.880 1434.385 ;
        RECT 2407.435 1434.385 2408.440 1434.685 ;
        RECT 2407.435 1434.345 2407.810 1434.385 ;
        RECT 2408.140 1431.995 2408.440 1434.385 ;
        RECT 2425.995 1434.385 2427.000 1434.685 ;
        RECT 2425.995 1434.345 2426.370 1434.385 ;
        RECT 2426.700 1431.995 2427.000 1434.385 ;
        RECT 2444.555 1434.385 2445.560 1434.685 ;
        RECT 2444.555 1434.345 2444.930 1434.385 ;
        RECT 2445.260 1431.995 2445.560 1434.385 ;
        RECT 2361.185 1431.695 2371.320 1431.995 ;
        RECT 2379.745 1431.695 2389.880 1431.995 ;
        RECT 2398.305 1431.695 2408.440 1431.995 ;
        RECT 2416.865 1431.695 2427.000 1431.995 ;
        RECT 2435.425 1431.695 2445.560 1431.995 ;
        RECT 2361.185 1429.015 2361.485 1431.695 ;
        RECT 2361.785 1430.155 2362.110 1430.160 ;
        RECT 2361.785 1429.825 2362.520 1430.155 ;
        RECT 2361.785 1429.820 2362.110 1429.825 ;
        RECT 2364.260 1429.600 2364.560 1431.695 ;
        RECT 2364.225 1429.595 2364.560 1429.600 ;
        RECT 2364.225 1429.265 2364.960 1429.595 ;
        RECT 2364.225 1429.260 2364.555 1429.265 ;
        RECT 2365.695 1429.040 2365.995 1431.695 ;
        RECT 2368.105 1430.155 2368.435 1430.160 ;
        RECT 2370.070 1430.155 2370.395 1430.160 ;
        RECT 2371.075 1430.155 2371.395 1430.160 ;
        RECT 2368.105 1429.825 2368.840 1430.155 ;
        RECT 2369.810 1429.825 2370.540 1430.155 ;
        RECT 2370.840 1429.825 2371.400 1430.155 ;
        RECT 2368.105 1429.820 2368.435 1429.825 ;
        RECT 2370.070 1429.820 2370.395 1429.825 ;
        RECT 2366.905 1429.595 2367.225 1429.600 ;
        RECT 2366.905 1429.260 2367.460 1429.595 ;
        RECT 2362.120 1429.035 2362.640 1429.040 ;
        RECT 2365.665 1429.035 2365.995 1429.040 ;
        RECT 2362.120 1429.015 2362.850 1429.035 ;
        RECT 2361.185 1428.715 2362.850 1429.015 ;
        RECT 2362.120 1428.705 2362.850 1428.715 ;
        RECT 2365.665 1428.705 2366.400 1429.035 ;
        RECT 2365.665 1428.700 2365.990 1428.705 ;
        RECT 2367.160 1428.465 2367.460 1429.260 ;
        RECT 2370.840 1428.465 2371.140 1429.825 ;
        RECT 2379.745 1429.015 2380.045 1431.695 ;
        RECT 2380.345 1430.155 2380.670 1430.160 ;
        RECT 2380.345 1429.825 2381.080 1430.155 ;
        RECT 2380.345 1429.820 2380.670 1429.825 ;
        RECT 2382.820 1429.600 2383.120 1431.695 ;
        RECT 2382.785 1429.595 2383.120 1429.600 ;
        RECT 2382.785 1429.265 2383.520 1429.595 ;
        RECT 2382.785 1429.260 2383.115 1429.265 ;
        RECT 2384.255 1429.040 2384.555 1431.695 ;
        RECT 2386.665 1430.155 2386.995 1430.160 ;
        RECT 2388.630 1430.155 2388.955 1430.160 ;
        RECT 2389.635 1430.155 2389.955 1430.160 ;
        RECT 2386.665 1429.825 2387.400 1430.155 ;
        RECT 2388.370 1429.825 2389.100 1430.155 ;
        RECT 2389.400 1429.825 2389.960 1430.155 ;
        RECT 2386.665 1429.820 2386.995 1429.825 ;
        RECT 2388.630 1429.820 2388.955 1429.825 ;
        RECT 2385.465 1429.595 2385.785 1429.600 ;
        RECT 2385.465 1429.260 2386.020 1429.595 ;
        RECT 2380.680 1429.035 2381.200 1429.040 ;
        RECT 2384.225 1429.035 2384.555 1429.040 ;
        RECT 2380.680 1429.015 2381.410 1429.035 ;
        RECT 2379.745 1428.715 2381.410 1429.015 ;
        RECT 2380.680 1428.705 2381.410 1428.715 ;
        RECT 2384.225 1428.705 2384.960 1429.035 ;
        RECT 2384.225 1428.700 2384.550 1428.705 ;
        RECT 2367.160 1428.165 2371.140 1428.465 ;
        RECT 2372.025 1428.475 2372.350 1428.480 ;
        RECT 2372.025 1428.145 2372.760 1428.475 ;
        RECT 2385.720 1428.465 2386.020 1429.260 ;
        RECT 2389.400 1428.465 2389.700 1429.825 ;
        RECT 2398.305 1429.015 2398.605 1431.695 ;
        RECT 2398.905 1430.155 2399.230 1430.160 ;
        RECT 2398.905 1429.825 2399.640 1430.155 ;
        RECT 2398.905 1429.820 2399.230 1429.825 ;
        RECT 2401.380 1429.600 2401.680 1431.695 ;
        RECT 2401.345 1429.595 2401.680 1429.600 ;
        RECT 2401.345 1429.265 2402.080 1429.595 ;
        RECT 2401.345 1429.260 2401.675 1429.265 ;
        RECT 2402.815 1429.040 2403.115 1431.695 ;
        RECT 2405.225 1430.155 2405.555 1430.160 ;
        RECT 2407.190 1430.155 2407.515 1430.160 ;
        RECT 2408.195 1430.155 2408.515 1430.160 ;
        RECT 2405.225 1429.825 2405.960 1430.155 ;
        RECT 2406.930 1429.825 2407.660 1430.155 ;
        RECT 2407.960 1429.825 2408.520 1430.155 ;
        RECT 2405.225 1429.820 2405.555 1429.825 ;
        RECT 2407.190 1429.820 2407.515 1429.825 ;
        RECT 2404.025 1429.595 2404.345 1429.600 ;
        RECT 2404.025 1429.260 2404.580 1429.595 ;
        RECT 2399.240 1429.035 2399.760 1429.040 ;
        RECT 2402.785 1429.035 2403.115 1429.040 ;
        RECT 2399.240 1429.015 2399.970 1429.035 ;
        RECT 2398.305 1428.715 2399.970 1429.015 ;
        RECT 2399.240 1428.705 2399.970 1428.715 ;
        RECT 2402.785 1428.705 2403.520 1429.035 ;
        RECT 2402.785 1428.700 2403.110 1428.705 ;
        RECT 2385.720 1428.165 2389.700 1428.465 ;
        RECT 2390.585 1428.475 2390.910 1428.480 ;
        RECT 2390.585 1428.145 2391.320 1428.475 ;
        RECT 2404.280 1428.465 2404.580 1429.260 ;
        RECT 2407.960 1428.465 2408.260 1429.825 ;
        RECT 2416.865 1429.015 2417.165 1431.695 ;
        RECT 2417.465 1430.155 2417.790 1430.160 ;
        RECT 2417.465 1429.825 2418.200 1430.155 ;
        RECT 2417.465 1429.820 2417.790 1429.825 ;
        RECT 2419.940 1429.600 2420.240 1431.695 ;
        RECT 2419.905 1429.595 2420.240 1429.600 ;
        RECT 2419.905 1429.265 2420.640 1429.595 ;
        RECT 2419.905 1429.260 2420.235 1429.265 ;
        RECT 2421.375 1429.040 2421.675 1431.695 ;
        RECT 2423.785 1430.155 2424.115 1430.160 ;
        RECT 2425.750 1430.155 2426.075 1430.160 ;
        RECT 2426.755 1430.155 2427.075 1430.160 ;
        RECT 2423.785 1429.825 2424.520 1430.155 ;
        RECT 2425.490 1429.825 2426.220 1430.155 ;
        RECT 2426.520 1429.825 2427.080 1430.155 ;
        RECT 2423.785 1429.820 2424.115 1429.825 ;
        RECT 2425.750 1429.820 2426.075 1429.825 ;
        RECT 2422.585 1429.595 2422.905 1429.600 ;
        RECT 2422.585 1429.260 2423.140 1429.595 ;
        RECT 2417.800 1429.035 2418.320 1429.040 ;
        RECT 2421.345 1429.035 2421.675 1429.040 ;
        RECT 2417.800 1429.015 2418.530 1429.035 ;
        RECT 2416.865 1428.715 2418.530 1429.015 ;
        RECT 2417.800 1428.705 2418.530 1428.715 ;
        RECT 2421.345 1428.705 2422.080 1429.035 ;
        RECT 2421.345 1428.700 2421.670 1428.705 ;
        RECT 2404.280 1428.165 2408.260 1428.465 ;
        RECT 2409.145 1428.475 2409.470 1428.480 ;
        RECT 2409.145 1428.145 2409.880 1428.475 ;
        RECT 2422.840 1428.465 2423.140 1429.260 ;
        RECT 2426.520 1428.465 2426.820 1429.825 ;
        RECT 2435.425 1429.015 2435.725 1431.695 ;
        RECT 2436.025 1430.155 2436.350 1430.160 ;
        RECT 2436.025 1429.825 2436.760 1430.155 ;
        RECT 2436.025 1429.820 2436.350 1429.825 ;
        RECT 2438.500 1429.600 2438.800 1431.695 ;
        RECT 2438.465 1429.595 2438.800 1429.600 ;
        RECT 2438.465 1429.265 2439.200 1429.595 ;
        RECT 2438.465 1429.260 2438.795 1429.265 ;
        RECT 2439.935 1429.040 2440.235 1431.695 ;
        RECT 2523.535 1430.915 2691.085 1431.245 ;
        RECT 2442.345 1430.155 2442.675 1430.160 ;
        RECT 2444.310 1430.155 2444.635 1430.160 ;
        RECT 2445.315 1430.155 2445.635 1430.160 ;
        RECT 2442.345 1429.825 2443.080 1430.155 ;
        RECT 2444.050 1429.825 2444.780 1430.155 ;
        RECT 2445.080 1429.825 2445.640 1430.155 ;
        RECT 2442.345 1429.820 2442.675 1429.825 ;
        RECT 2444.310 1429.820 2444.635 1429.825 ;
        RECT 2441.145 1429.595 2441.465 1429.600 ;
        RECT 2441.145 1429.260 2441.700 1429.595 ;
        RECT 2436.360 1429.035 2436.880 1429.040 ;
        RECT 2439.905 1429.035 2440.235 1429.040 ;
        RECT 2436.360 1429.015 2437.090 1429.035 ;
        RECT 2435.425 1428.715 2437.090 1429.015 ;
        RECT 2436.360 1428.705 2437.090 1428.715 ;
        RECT 2439.905 1428.705 2440.640 1429.035 ;
        RECT 2439.905 1428.700 2440.230 1428.705 ;
        RECT 2422.840 1428.165 2426.820 1428.465 ;
        RECT 2427.705 1428.475 2428.030 1428.480 ;
        RECT 2427.705 1428.145 2428.440 1428.475 ;
        RECT 2441.400 1428.465 2441.700 1429.260 ;
        RECT 2445.080 1428.465 2445.380 1429.825 ;
        RECT 2690.755 1429.560 2691.085 1430.915 ;
        RECT 2690.000 1429.410 2694.000 1429.560 ;
        RECT 2694.665 1429.410 2694.995 1429.425 ;
        RECT 2690.000 1429.110 2694.995 1429.410 ;
        RECT 2690.000 1428.960 2694.000 1429.110 ;
        RECT 2694.665 1429.095 2694.995 1429.110 ;
        RECT 2441.400 1428.165 2445.380 1428.465 ;
        RECT 2446.265 1428.475 2446.590 1428.480 ;
        RECT 2446.265 1428.145 2447.000 1428.475 ;
        RECT 2372.025 1428.140 2372.350 1428.145 ;
        RECT 2390.585 1428.140 2390.910 1428.145 ;
        RECT 2409.145 1428.140 2409.470 1428.145 ;
        RECT 2427.705 1428.140 2428.030 1428.145 ;
        RECT 2446.265 1428.140 2446.590 1428.145 ;
        RECT 2670.405 1423.045 2690.330 1423.375 ;
        RECT 2670.405 1417.055 2670.735 1423.045 ;
        RECT 2690.000 1422.760 2690.330 1423.045 ;
        RECT 2690.000 1422.610 2694.000 1422.760 ;
        RECT 2694.665 1422.610 2694.995 1422.625 ;
        RECT 2690.000 1422.310 2694.995 1422.610 ;
        RECT 2690.000 1422.160 2694.000 1422.310 ;
        RECT 2694.665 1422.295 2694.995 1422.310 ;
        RECT 2523.535 1416.725 2670.735 1417.055 ;
        RECT 2672.730 1415.960 2690.610 1416.005 ;
        RECT 2672.730 1415.810 2694.000 1415.960 ;
        RECT 2694.665 1415.810 2694.995 1415.825 ;
        RECT 2672.730 1415.675 2694.995 1415.810 ;
        RECT 2672.730 1409.525 2673.060 1415.675 ;
        RECT 2690.000 1415.510 2694.995 1415.675 ;
        RECT 2690.000 1415.360 2694.000 1415.510 ;
        RECT 2694.665 1415.495 2694.995 1415.510 ;
        RECT 2523.535 1409.195 2673.060 1409.525 ;
        RECT 2690.000 1409.080 2694.000 1409.160 ;
        RECT 2676.470 1409.010 2694.000 1409.080 ;
        RECT 2694.665 1409.010 2694.995 1409.025 ;
        RECT 2676.470 1408.750 2694.995 1409.010 ;
        RECT 2676.470 1403.545 2676.800 1408.750 ;
        RECT 2690.000 1408.710 2694.995 1408.750 ;
        RECT 2690.000 1408.560 2694.000 1408.710 ;
        RECT 2694.665 1408.695 2694.995 1408.710 ;
        RECT 2523.535 1403.215 2676.800 1403.545 ;
        RECT 2698.345 1402.890 2698.675 1402.905 ;
        RECT 2694.910 1402.590 2698.675 1402.890 ;
        RECT 2690.000 1402.210 2694.000 1402.360 ;
        RECT 2694.910 1402.210 2695.210 1402.590 ;
        RECT 2698.345 1402.575 2698.675 1402.590 ;
        RECT 2690.000 1401.910 2695.210 1402.210 ;
        RECT 2690.000 1401.760 2694.000 1401.910 ;
        RECT 2691.075 1395.130 2691.405 1401.760 ;
        RECT 2523.535 1394.800 2691.405 1395.130 ;
        RECT 2377.015 1334.345 2377.385 1334.715 ;
        RECT 2392.275 1334.345 2392.645 1334.715 ;
        RECT 2407.535 1334.345 2407.905 1334.715 ;
        RECT 2422.795 1334.345 2423.165 1334.715 ;
        RECT 2438.055 1334.345 2438.425 1334.715 ;
        RECT 2377.050 1331.070 2377.350 1334.345 ;
        RECT 2392.310 1331.070 2392.610 1334.345 ;
        RECT 2407.570 1331.070 2407.870 1334.345 ;
        RECT 2422.830 1331.070 2423.130 1334.345 ;
        RECT 2438.090 1331.070 2438.390 1334.345 ;
        RECT 2372.815 1330.770 2377.350 1331.070 ;
        RECT 2388.075 1330.770 2392.610 1331.070 ;
        RECT 2403.335 1330.770 2407.870 1331.070 ;
        RECT 2418.595 1330.770 2423.130 1331.070 ;
        RECT 2433.855 1330.770 2438.390 1331.070 ;
        RECT 2372.815 1330.550 2375.910 1330.770 ;
        RECT 2372.815 1329.600 2373.115 1330.550 ;
        RECT 2375.610 1330.145 2375.910 1330.550 ;
        RECT 2388.075 1330.550 2391.170 1330.770 ;
        RECT 2376.335 1330.145 2376.665 1330.155 ;
        RECT 2374.425 1329.845 2376.665 1330.145 ;
        RECT 2372.735 1329.595 2373.115 1329.600 ;
        RECT 2372.505 1329.265 2373.235 1329.595 ;
        RECT 2373.695 1329.245 2374.015 1329.625 ;
        RECT 2373.695 1329.055 2374.025 1329.245 ;
        RECT 2374.425 1329.055 2374.725 1329.845 ;
        RECT 2375.610 1329.155 2375.910 1329.845 ;
        RECT 2376.325 1329.795 2376.665 1329.845 ;
        RECT 2388.075 1329.600 2388.375 1330.550 ;
        RECT 2390.870 1330.145 2391.170 1330.550 ;
        RECT 2403.335 1330.550 2406.430 1330.770 ;
        RECT 2391.595 1330.145 2391.925 1330.155 ;
        RECT 2389.685 1329.845 2391.925 1330.145 ;
        RECT 2387.995 1329.595 2388.375 1329.600 ;
        RECT 2373.695 1328.705 2374.030 1329.055 ;
        RECT 2374.405 1329.040 2374.725 1329.055 ;
        RECT 2374.405 1328.705 2374.745 1329.040 ;
        RECT 2375.405 1328.815 2376.185 1329.155 ;
        RECT 2375.610 1328.810 2376.185 1328.815 ;
        RECT 2375.845 1328.805 2376.185 1328.810 ;
        RECT 2375.855 1328.775 2376.185 1328.805 ;
        RECT 2380.720 1328.940 2381.080 1329.365 ;
        RECT 2387.765 1329.265 2388.495 1329.595 ;
        RECT 2388.955 1329.245 2389.275 1329.625 ;
        RECT 2388.955 1329.055 2389.285 1329.245 ;
        RECT 2389.685 1329.055 2389.985 1329.845 ;
        RECT 2390.870 1329.155 2391.170 1329.845 ;
        RECT 2391.585 1329.795 2391.925 1329.845 ;
        RECT 2403.335 1329.600 2403.635 1330.550 ;
        RECT 2406.130 1330.145 2406.430 1330.550 ;
        RECT 2418.595 1330.550 2421.690 1330.770 ;
        RECT 2406.855 1330.145 2407.185 1330.155 ;
        RECT 2404.945 1329.845 2407.185 1330.145 ;
        RECT 2403.255 1329.595 2403.635 1329.600 ;
        RECT 2374.975 1328.175 2375.705 1328.505 ;
        RECT 2376.520 1328.495 2376.870 1328.500 ;
        RECT 2374.975 1328.165 2375.455 1328.175 ;
        RECT 2375.130 1327.700 2375.430 1328.165 ;
        RECT 2376.520 1328.145 2377.255 1328.495 ;
        RECT 2377.555 1328.165 2378.295 1328.495 ;
        RECT 2379.415 1328.475 2379.775 1328.480 ;
        RECT 2377.555 1328.155 2377.885 1328.165 ;
        RECT 2379.255 1328.145 2379.985 1328.475 ;
        RECT 2376.520 1328.140 2376.870 1328.145 ;
        RECT 2379.415 1328.140 2379.775 1328.145 ;
        RECT 2380.720 1327.700 2381.060 1328.940 ;
        RECT 2388.955 1328.705 2389.290 1329.055 ;
        RECT 2389.665 1329.040 2389.985 1329.055 ;
        RECT 2389.665 1328.705 2390.005 1329.040 ;
        RECT 2390.665 1328.815 2391.445 1329.155 ;
        RECT 2390.870 1328.810 2391.445 1328.815 ;
        RECT 2391.105 1328.805 2391.445 1328.810 ;
        RECT 2391.115 1328.775 2391.445 1328.805 ;
        RECT 2395.980 1328.940 2396.340 1329.365 ;
        RECT 2403.025 1329.265 2403.755 1329.595 ;
        RECT 2404.215 1329.245 2404.535 1329.625 ;
        RECT 2404.215 1329.055 2404.545 1329.245 ;
        RECT 2404.945 1329.055 2405.245 1329.845 ;
        RECT 2406.130 1329.155 2406.430 1329.845 ;
        RECT 2406.845 1329.795 2407.185 1329.845 ;
        RECT 2418.595 1329.600 2418.895 1330.550 ;
        RECT 2421.390 1330.145 2421.690 1330.550 ;
        RECT 2433.855 1330.550 2436.950 1330.770 ;
        RECT 2422.115 1330.145 2422.445 1330.155 ;
        RECT 2420.205 1329.845 2422.445 1330.145 ;
        RECT 2418.515 1329.595 2418.895 1329.600 ;
        RECT 2390.235 1328.175 2390.965 1328.505 ;
        RECT 2391.780 1328.495 2392.130 1328.500 ;
        RECT 2390.235 1328.165 2390.715 1328.175 ;
        RECT 2375.130 1327.400 2381.060 1327.700 ;
        RECT 2390.390 1327.700 2390.690 1328.165 ;
        RECT 2391.780 1328.145 2392.515 1328.495 ;
        RECT 2392.815 1328.165 2393.555 1328.495 ;
        RECT 2394.675 1328.475 2395.035 1328.480 ;
        RECT 2392.815 1328.155 2393.145 1328.165 ;
        RECT 2394.515 1328.145 2395.245 1328.475 ;
        RECT 2391.780 1328.140 2392.130 1328.145 ;
        RECT 2394.675 1328.140 2395.035 1328.145 ;
        RECT 2395.980 1327.700 2396.320 1328.940 ;
        RECT 2404.215 1328.705 2404.550 1329.055 ;
        RECT 2404.925 1329.040 2405.245 1329.055 ;
        RECT 2404.925 1328.705 2405.265 1329.040 ;
        RECT 2405.925 1328.815 2406.705 1329.155 ;
        RECT 2406.130 1328.810 2406.705 1328.815 ;
        RECT 2406.365 1328.805 2406.705 1328.810 ;
        RECT 2406.375 1328.775 2406.705 1328.805 ;
        RECT 2411.240 1328.940 2411.600 1329.365 ;
        RECT 2418.285 1329.265 2419.015 1329.595 ;
        RECT 2419.475 1329.245 2419.795 1329.625 ;
        RECT 2419.475 1329.055 2419.805 1329.245 ;
        RECT 2420.205 1329.055 2420.505 1329.845 ;
        RECT 2421.390 1329.155 2421.690 1329.845 ;
        RECT 2422.105 1329.795 2422.445 1329.845 ;
        RECT 2433.855 1329.600 2434.155 1330.550 ;
        RECT 2436.650 1330.145 2436.950 1330.550 ;
        RECT 2437.375 1330.145 2437.705 1330.155 ;
        RECT 2435.465 1329.845 2437.705 1330.145 ;
        RECT 2433.775 1329.595 2434.155 1329.600 ;
        RECT 2405.495 1328.175 2406.225 1328.505 ;
        RECT 2407.040 1328.495 2407.390 1328.500 ;
        RECT 2405.495 1328.165 2405.975 1328.175 ;
        RECT 2390.390 1327.400 2396.320 1327.700 ;
        RECT 2405.650 1327.700 2405.950 1328.165 ;
        RECT 2407.040 1328.145 2407.775 1328.495 ;
        RECT 2408.075 1328.165 2408.815 1328.495 ;
        RECT 2409.935 1328.475 2410.295 1328.480 ;
        RECT 2408.075 1328.155 2408.405 1328.165 ;
        RECT 2409.775 1328.145 2410.505 1328.475 ;
        RECT 2407.040 1328.140 2407.390 1328.145 ;
        RECT 2409.935 1328.140 2410.295 1328.145 ;
        RECT 2411.240 1327.700 2411.580 1328.940 ;
        RECT 2419.475 1328.705 2419.810 1329.055 ;
        RECT 2420.185 1329.040 2420.505 1329.055 ;
        RECT 2420.185 1328.705 2420.525 1329.040 ;
        RECT 2421.185 1328.815 2421.965 1329.155 ;
        RECT 2421.390 1328.810 2421.965 1328.815 ;
        RECT 2421.625 1328.805 2421.965 1328.810 ;
        RECT 2421.635 1328.775 2421.965 1328.805 ;
        RECT 2426.500 1328.940 2426.860 1329.365 ;
        RECT 2433.545 1329.265 2434.275 1329.595 ;
        RECT 2434.735 1329.245 2435.055 1329.625 ;
        RECT 2434.735 1329.055 2435.065 1329.245 ;
        RECT 2435.465 1329.055 2435.765 1329.845 ;
        RECT 2436.650 1329.155 2436.950 1329.845 ;
        RECT 2437.365 1329.795 2437.705 1329.845 ;
        RECT 2420.755 1328.175 2421.485 1328.505 ;
        RECT 2422.300 1328.495 2422.650 1328.500 ;
        RECT 2420.755 1328.165 2421.235 1328.175 ;
        RECT 2405.650 1327.400 2411.580 1327.700 ;
        RECT 2420.910 1327.700 2421.210 1328.165 ;
        RECT 2422.300 1328.145 2423.035 1328.495 ;
        RECT 2423.335 1328.165 2424.075 1328.495 ;
        RECT 2425.195 1328.475 2425.555 1328.480 ;
        RECT 2423.335 1328.155 2423.665 1328.165 ;
        RECT 2425.035 1328.145 2425.765 1328.475 ;
        RECT 2422.300 1328.140 2422.650 1328.145 ;
        RECT 2425.195 1328.140 2425.555 1328.145 ;
        RECT 2426.500 1327.700 2426.840 1328.940 ;
        RECT 2434.735 1328.705 2435.070 1329.055 ;
        RECT 2435.445 1329.040 2435.765 1329.055 ;
        RECT 2435.445 1328.705 2435.785 1329.040 ;
        RECT 2436.445 1328.815 2437.225 1329.155 ;
        RECT 2436.650 1328.810 2437.225 1328.815 ;
        RECT 2436.885 1328.805 2437.225 1328.810 ;
        RECT 2436.895 1328.775 2437.225 1328.805 ;
        RECT 2441.760 1328.940 2442.120 1329.365 ;
        RECT 2436.015 1328.175 2436.745 1328.505 ;
        RECT 2437.560 1328.495 2437.910 1328.500 ;
        RECT 2436.015 1328.165 2436.495 1328.175 ;
        RECT 2420.910 1327.400 2426.840 1327.700 ;
        RECT 2436.170 1327.700 2436.470 1328.165 ;
        RECT 2437.560 1328.145 2438.295 1328.495 ;
        RECT 2438.595 1328.165 2439.335 1328.495 ;
        RECT 2440.455 1328.475 2440.815 1328.480 ;
        RECT 2438.595 1328.155 2438.925 1328.165 ;
        RECT 2440.295 1328.145 2441.025 1328.475 ;
        RECT 2437.560 1328.140 2437.910 1328.145 ;
        RECT 2440.455 1328.140 2440.815 1328.145 ;
        RECT 2441.760 1327.700 2442.100 1328.940 ;
        RECT 2436.170 1327.400 2442.100 1327.700 ;
      LAYER met4 ;
        RECT 2400.575 2139.455 2400.905 2139.785 ;
        RECT 2432.775 2139.455 2433.105 2139.785 ;
        RECT 2400.590 2037.785 2400.890 2139.455 ;
        RECT 2400.575 2037.455 2400.905 2037.785 ;
        RECT 2414.375 2035.415 2414.705 2035.745 ;
        RECT 2428.175 2035.415 2428.505 2035.745 ;
        RECT 2414.390 1850.785 2414.690 2035.415 ;
        RECT 2414.375 1850.455 2414.705 1850.785 ;
        RECT 2373.635 1784.265 2373.975 1784.600 ;
        RECT 2388.895 1784.265 2389.235 1784.600 ;
        RECT 2404.155 1784.265 2404.495 1784.600 ;
        RECT 2419.415 1784.265 2419.755 1784.600 ;
        RECT 2373.655 1784.095 2373.975 1784.265 ;
        RECT 2375.795 1784.095 2376.135 1784.135 ;
        RECT 2373.655 1783.795 2376.135 1784.095 ;
        RECT 2388.915 1784.095 2389.235 1784.265 ;
        RECT 2391.055 1784.095 2391.395 1784.135 ;
        RECT 2388.915 1783.795 2391.395 1784.095 ;
        RECT 2404.175 1784.095 2404.495 1784.265 ;
        RECT 2406.315 1784.095 2406.655 1784.135 ;
        RECT 2404.175 1783.795 2406.655 1784.095 ;
        RECT 2419.435 1784.095 2419.755 1784.265 ;
        RECT 2421.575 1784.095 2421.915 1784.135 ;
        RECT 2419.435 1783.795 2421.915 1784.095 ;
        RECT 2375.805 1783.775 2376.135 1783.795 ;
        RECT 2391.065 1783.775 2391.395 1783.795 ;
        RECT 2406.325 1783.775 2406.655 1783.795 ;
        RECT 2421.585 1783.775 2421.915 1783.795 ;
        RECT 2428.190 1670.585 2428.490 2035.415 ;
        RECT 2432.790 1677.385 2433.090 2139.455 ;
        RECT 2433.695 1932.055 2434.025 1932.385 ;
        RECT 2432.775 1677.055 2433.105 1677.385 ;
        RECT 2428.175 1670.255 2428.505 1670.585 ;
        RECT 2433.710 1663.785 2434.010 1932.055 ;
        RECT 2434.675 1784.265 2435.015 1784.600 ;
        RECT 2434.695 1784.095 2435.015 1784.265 ;
        RECT 2436.835 1784.095 2437.175 1784.135 ;
        RECT 2434.695 1783.795 2437.175 1784.095 ;
        RECT 2436.845 1783.775 2437.175 1783.795 ;
        RECT 2433.695 1663.455 2434.025 1663.785 ;
        RECT 2373.685 1329.265 2374.025 1329.600 ;
        RECT 2388.945 1329.265 2389.285 1329.600 ;
        RECT 2404.205 1329.265 2404.545 1329.600 ;
        RECT 2419.465 1329.265 2419.805 1329.600 ;
        RECT 2434.725 1329.265 2435.065 1329.600 ;
        RECT 2373.705 1329.095 2374.025 1329.265 ;
        RECT 2375.845 1329.095 2376.185 1329.135 ;
        RECT 2373.705 1328.795 2376.185 1329.095 ;
        RECT 2388.965 1329.095 2389.285 1329.265 ;
        RECT 2391.105 1329.095 2391.445 1329.135 ;
        RECT 2388.965 1328.795 2391.445 1329.095 ;
        RECT 2404.225 1329.095 2404.545 1329.265 ;
        RECT 2406.365 1329.095 2406.705 1329.135 ;
        RECT 2404.225 1328.795 2406.705 1329.095 ;
        RECT 2419.485 1329.095 2419.805 1329.265 ;
        RECT 2421.625 1329.095 2421.965 1329.135 ;
        RECT 2419.485 1328.795 2421.965 1329.095 ;
        RECT 2434.745 1329.095 2435.065 1329.265 ;
        RECT 2436.885 1329.095 2437.225 1329.135 ;
        RECT 2434.745 1328.795 2437.225 1329.095 ;
        RECT 2375.855 1328.775 2376.185 1328.795 ;
        RECT 2391.115 1328.775 2391.445 1328.795 ;
        RECT 2406.375 1328.775 2406.705 1328.795 ;
        RECT 2421.635 1328.775 2421.965 1328.795 ;
        RECT 2436.895 1328.775 2437.225 1328.795 ;
  END
END user_project_wrapper
END LIBRARY

