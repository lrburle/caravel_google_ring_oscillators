magic
tech sky130A
magscale 1 2
timestamp 1712673195
<< nwell >>
rect -38 260 1970 582
<< pwell >>
rect 32 -12 66 16
rect 28 -16 66 -12
rect 520 -16 554 16
rect 1008 -16 1042 16
rect 1496 -12 1530 16
rect 1496 -16 1534 -12
rect 28 -18 62 -16
rect 1500 -18 1534 -16
<< nmos >>
rect 116 46 146 176
rect 212 46 242 176
rect 308 46 338 176
rect 404 46 434 176
rect 604 46 634 176
rect 700 46 730 176
rect 796 46 826 176
rect 892 46 922 176
rect 1092 46 1122 176
rect 1188 46 1218 176
rect 1284 46 1314 176
rect 1380 46 1410 176
rect 1580 46 1610 176
rect 1676 46 1706 176
rect 1772 46 1802 176
<< pmos >>
rect 116 296 146 496
rect 212 296 242 496
rect 308 296 338 496
rect 404 296 434 496
rect 604 296 634 496
rect 700 296 730 496
rect 796 296 826 496
rect 892 296 922 496
rect 1092 296 1122 496
rect 1188 296 1218 496
rect 1284 296 1314 496
rect 1380 296 1410 496
rect 1580 296 1610 496
rect 1676 296 1706 496
rect 1772 296 1802 496
<< ndiff >>
rect 58 100 116 176
rect 58 66 66 100
rect 100 66 116 100
rect 58 46 116 66
rect 146 100 212 176
rect 146 66 162 100
rect 196 66 212 100
rect 146 46 212 66
rect 242 100 308 176
rect 242 66 258 100
rect 292 66 308 100
rect 242 46 308 66
rect 338 100 404 176
rect 338 66 354 100
rect 388 66 404 100
rect 338 46 404 66
rect 434 100 492 176
rect 434 66 450 100
rect 484 66 492 100
rect 434 46 492 66
rect 546 100 604 176
rect 546 66 554 100
rect 588 66 604 100
rect 546 46 604 66
rect 634 100 700 176
rect 634 66 650 100
rect 684 66 700 100
rect 634 46 700 66
rect 730 100 796 176
rect 730 66 746 100
rect 780 66 796 100
rect 730 46 796 66
rect 826 46 892 176
rect 922 168 980 176
rect 922 134 934 168
rect 968 134 980 168
rect 922 46 980 134
rect 1034 100 1092 176
rect 1034 66 1042 100
rect 1076 66 1092 100
rect 1034 46 1092 66
rect 1122 46 1188 176
rect 1218 100 1284 176
rect 1218 66 1234 100
rect 1268 66 1284 100
rect 1218 46 1284 66
rect 1314 46 1380 176
rect 1410 100 1468 176
rect 1410 66 1426 100
rect 1460 66 1468 100
rect 1410 46 1468 66
rect 1522 100 1580 176
rect 1522 66 1530 100
rect 1564 66 1580 100
rect 1522 46 1580 66
rect 1610 100 1676 176
rect 1610 66 1626 100
rect 1660 66 1676 100
rect 1610 46 1676 66
rect 1706 46 1772 176
rect 1802 100 1860 176
rect 1802 66 1818 100
rect 1852 66 1860 100
rect 1802 46 1860 66
<< pdiff >>
rect 58 378 116 496
rect 58 344 66 378
rect 100 344 116 378
rect 58 296 116 344
rect 146 296 212 496
rect 242 476 308 496
rect 242 442 258 476
rect 292 442 308 476
rect 242 296 308 442
rect 338 296 404 496
rect 434 378 492 496
rect 434 344 450 378
rect 484 344 492 378
rect 434 296 492 344
rect 546 378 604 496
rect 546 344 554 378
rect 588 344 604 378
rect 546 296 604 344
rect 634 296 700 496
rect 730 476 796 496
rect 730 442 746 476
rect 780 442 796 476
rect 730 296 796 442
rect 826 378 892 496
rect 826 344 842 378
rect 876 344 892 378
rect 826 296 892 344
rect 922 476 980 496
rect 922 442 938 476
rect 972 442 980 476
rect 922 296 980 442
rect 1034 378 1092 496
rect 1034 344 1042 378
rect 1076 344 1092 378
rect 1034 296 1092 344
rect 1122 476 1188 496
rect 1122 442 1138 476
rect 1172 442 1188 476
rect 1122 296 1188 442
rect 1218 378 1284 496
rect 1218 344 1234 378
rect 1268 344 1284 378
rect 1218 296 1284 344
rect 1314 446 1380 496
rect 1314 412 1330 446
rect 1364 412 1380 446
rect 1314 296 1380 412
rect 1410 378 1468 496
rect 1410 344 1426 378
rect 1460 344 1468 378
rect 1410 296 1468 344
rect 1522 446 1580 496
rect 1522 412 1530 446
rect 1564 412 1580 446
rect 1522 296 1580 412
rect 1610 476 1676 496
rect 1610 442 1626 476
rect 1660 442 1676 476
rect 1610 296 1676 442
rect 1706 378 1772 496
rect 1706 344 1722 378
rect 1756 344 1772 378
rect 1706 296 1772 344
rect 1802 476 1860 496
rect 1802 442 1818 476
rect 1852 442 1860 476
rect 1802 296 1860 442
<< ndiffc >>
rect 66 66 100 100
rect 162 66 196 100
rect 258 66 292 100
rect 354 66 388 100
rect 450 66 484 100
rect 554 66 588 100
rect 650 66 684 100
rect 746 66 780 100
rect 934 134 968 168
rect 1042 66 1076 100
rect 1234 66 1268 100
rect 1426 66 1460 100
rect 1530 66 1564 100
rect 1626 66 1660 100
rect 1818 66 1852 100
<< pdiffc >>
rect 66 344 100 378
rect 258 442 292 476
rect 450 344 484 378
rect 554 344 588 378
rect 746 442 780 476
rect 842 344 876 378
rect 938 442 972 476
rect 1042 344 1076 378
rect 1138 442 1172 476
rect 1234 344 1268 378
rect 1330 412 1364 446
rect 1426 344 1460 378
rect 1530 412 1564 446
rect 1626 442 1660 476
rect 1722 344 1756 378
rect 1818 442 1852 476
<< poly >>
rect 116 496 146 522
rect 212 496 242 522
rect 308 496 338 522
rect 404 496 434 522
rect 604 496 634 522
rect 700 496 730 522
rect 796 496 826 522
rect 892 496 922 522
rect 1092 496 1122 522
rect 1188 496 1218 522
rect 1284 496 1314 522
rect 1380 496 1410 522
rect 1580 496 1610 522
rect 1676 496 1706 522
rect 1772 496 1802 522
rect 116 264 146 296
rect 212 264 242 296
rect 308 264 338 296
rect 404 264 434 296
rect 604 264 634 296
rect 700 264 730 296
rect 796 264 826 296
rect 892 264 922 296
rect 1092 264 1122 296
rect 1188 264 1218 296
rect 1284 264 1314 296
rect 1380 264 1410 296
rect 1580 264 1610 296
rect 1676 264 1706 296
rect 1772 264 1802 296
rect 104 248 158 264
rect 104 214 114 248
rect 148 214 158 248
rect 104 198 158 214
rect 200 248 254 264
rect 200 214 210 248
rect 244 214 254 248
rect 200 198 254 214
rect 296 248 350 264
rect 296 214 306 248
rect 340 214 350 248
rect 296 198 350 214
rect 392 248 446 264
rect 392 214 402 248
rect 436 214 446 248
rect 392 198 446 214
rect 592 248 646 264
rect 592 214 602 248
rect 636 214 646 248
rect 592 198 646 214
rect 688 248 742 264
rect 688 214 698 248
rect 732 214 742 248
rect 688 198 742 214
rect 784 248 838 264
rect 784 214 794 248
rect 828 214 838 248
rect 784 198 838 214
rect 880 248 934 264
rect 880 214 890 248
rect 924 214 934 248
rect 880 198 934 214
rect 1080 248 1134 264
rect 1080 214 1090 248
rect 1124 214 1134 248
rect 1080 198 1134 214
rect 1176 248 1230 264
rect 1176 214 1186 248
rect 1220 214 1230 248
rect 1176 198 1230 214
rect 1272 248 1326 264
rect 1272 214 1282 248
rect 1316 214 1326 248
rect 1272 198 1326 214
rect 1368 248 1422 264
rect 1368 214 1378 248
rect 1412 214 1422 248
rect 1368 198 1422 214
rect 1568 248 1622 264
rect 1568 214 1578 248
rect 1612 214 1622 248
rect 1568 198 1622 214
rect 1664 248 1718 264
rect 1664 214 1674 248
rect 1708 214 1718 248
rect 1664 198 1718 214
rect 1760 248 1814 264
rect 1760 214 1770 248
rect 1804 214 1814 248
rect 1760 198 1814 214
rect 116 176 146 198
rect 212 176 242 198
rect 308 176 338 198
rect 404 176 434 198
rect 604 176 634 198
rect 700 176 730 198
rect 796 176 826 198
rect 892 176 922 198
rect 1092 176 1122 198
rect 1188 176 1218 198
rect 1284 176 1314 198
rect 1380 176 1410 198
rect 1580 176 1610 198
rect 1676 176 1706 198
rect 1772 176 1802 198
rect 116 20 146 46
rect 212 20 242 46
rect 308 20 338 46
rect 404 20 434 46
rect 604 20 634 46
rect 700 20 730 46
rect 796 20 826 46
rect 892 20 922 46
rect 1092 20 1122 46
rect 1188 20 1218 46
rect 1284 20 1314 46
rect 1380 20 1410 46
rect 1580 20 1610 46
rect 1676 20 1706 46
rect 1772 20 1802 46
<< polycont >>
rect 114 214 148 248
rect 210 214 244 248
rect 306 214 340 248
rect 402 214 436 248
rect 602 214 636 248
rect 698 214 732 248
rect 794 214 828 248
rect 890 214 924 248
rect 1090 214 1124 248
rect 1186 214 1220 248
rect 1282 214 1316 248
rect 1378 214 1412 248
rect 1578 214 1612 248
rect 1674 214 1708 248
rect 1770 214 1804 248
<< locali >>
rect 0 526 28 560
rect 62 526 120 560
rect 154 526 212 560
rect 246 526 304 560
rect 338 526 396 560
rect 430 526 488 560
rect 522 526 580 560
rect 614 526 672 560
rect 706 526 764 560
rect 798 526 856 560
rect 890 526 948 560
rect 982 526 1040 560
rect 1074 526 1132 560
rect 1166 526 1224 560
rect 1258 526 1316 560
rect 1350 526 1408 560
rect 1442 526 1500 560
rect 1534 526 1592 560
rect 1626 526 1684 560
rect 1718 526 1776 560
rect 1810 526 1868 560
rect 1902 526 1932 560
rect 258 476 292 526
rect 138 422 162 456
rect 258 426 292 442
rect 746 476 780 526
rect 746 426 780 442
rect 938 476 972 526
rect 938 426 972 442
rect 1138 476 1172 526
rect 1626 476 1660 526
rect 1138 426 1172 442
rect 1330 456 1364 462
rect 66 378 100 394
rect 138 248 172 422
rect 436 378 484 400
rect 436 366 450 378
rect 98 214 114 248
rect 148 214 172 248
rect 210 310 306 344
rect 450 328 484 344
rect 554 378 588 394
rect 626 366 650 400
rect 1330 396 1364 412
rect 1530 456 1564 462
rect 1626 426 1660 442
rect 1818 476 1852 526
rect 1818 426 1852 442
rect 1530 396 1564 412
rect 210 248 244 310
rect 210 198 244 214
rect 306 248 340 264
rect 626 248 660 366
rect 1026 344 1042 378
rect 1076 344 1234 378
rect 1268 362 1284 378
rect 1410 362 1426 378
rect 1268 344 1426 362
rect 1460 344 1476 378
rect 1706 344 1722 378
rect 1756 344 1772 378
rect 842 328 876 344
rect 1234 328 1460 344
rect 1554 310 1756 344
rect 386 214 402 248
rect 436 232 484 248
rect 436 214 450 232
rect 586 214 602 248
rect 636 214 660 248
rect 698 248 732 264
rect 794 248 828 254
rect 1186 248 1220 264
rect 874 214 890 248
rect 924 214 1090 248
rect 1124 214 1140 248
rect 794 198 828 214
rect 1282 248 1316 254
rect 1426 248 1460 254
rect 1362 214 1378 248
rect 1412 214 1460 248
rect 1554 264 1588 310
rect 1554 248 1612 264
rect 1554 214 1578 248
rect 1282 198 1316 214
rect 1674 248 1708 264
rect 1818 248 1852 254
rect 1754 214 1770 248
rect 1804 214 1852 248
rect 924 142 934 168
rect 890 134 934 142
rect 968 134 988 168
rect 1412 142 1460 176
rect 66 100 100 116
rect 66 16 100 66
rect 162 50 196 66
rect 258 100 292 116
rect 258 16 292 66
rect 354 50 388 66
rect 450 100 484 116
rect 450 16 484 66
rect 554 100 588 116
rect 554 16 588 66
rect 650 50 684 66
rect 746 100 780 116
rect 746 16 780 66
rect 1042 50 1076 66
rect 1234 100 1268 116
rect 1234 16 1268 66
rect 1426 100 1460 142
rect 1426 50 1460 66
rect 1530 50 1564 66
rect 1626 100 1660 116
rect 1756 86 1818 100
rect 1722 66 1818 86
rect 1852 66 1868 100
rect 1626 16 1660 66
rect 0 -18 28 16
rect 62 -18 120 16
rect 154 -18 212 16
rect 246 -18 304 16
rect 338 -18 396 16
rect 430 -18 488 16
rect 522 -18 580 16
rect 614 -18 672 16
rect 706 -18 764 16
rect 798 -18 856 16
rect 890 -18 948 16
rect 982 -18 1040 16
rect 1074 -18 1132 16
rect 1166 -18 1224 16
rect 1258 -18 1316 16
rect 1350 -18 1408 16
rect 1442 -18 1500 16
rect 1534 -18 1592 16
rect 1626 -18 1684 16
rect 1718 -18 1776 16
rect 1810 -18 1868 16
rect 1902 -18 1932 16
<< viali >>
rect 28 526 62 560
rect 120 526 154 560
rect 212 526 246 560
rect 304 526 338 560
rect 396 526 430 560
rect 488 526 522 560
rect 580 526 614 560
rect 672 526 706 560
rect 764 526 798 560
rect 856 526 890 560
rect 948 526 982 560
rect 1040 526 1074 560
rect 1132 526 1166 560
rect 1224 526 1258 560
rect 1316 526 1350 560
rect 1408 526 1442 560
rect 1500 526 1534 560
rect 1592 526 1626 560
rect 1684 526 1718 560
rect 1776 526 1810 560
rect 1868 526 1902 560
rect 162 422 196 456
rect 1330 446 1364 456
rect 1330 422 1364 446
rect 66 310 100 344
rect 402 366 436 400
rect 306 310 340 344
rect 554 310 588 344
rect 650 366 684 400
rect 842 378 876 400
rect 1530 446 1564 456
rect 1530 422 1564 446
rect 842 366 876 378
rect 306 214 340 232
rect 306 198 340 214
rect 450 198 484 232
rect 698 214 732 232
rect 698 198 732 214
rect 794 254 828 288
rect 1090 214 1124 232
rect 1186 214 1220 232
rect 1090 198 1124 214
rect 1186 198 1220 214
rect 1282 254 1316 288
rect 1426 254 1460 288
rect 1578 214 1612 232
rect 1578 198 1612 214
rect 1818 254 1852 288
rect 1674 214 1708 232
rect 1674 198 1708 214
rect 890 142 924 176
rect 1378 142 1412 176
rect 162 100 196 120
rect 162 86 196 100
rect 354 100 388 120
rect 354 86 388 100
rect 650 100 684 120
rect 650 86 684 100
rect 1042 100 1076 120
rect 1042 86 1076 100
rect 1530 100 1564 120
rect 1530 86 1564 100
rect 1722 86 1756 120
rect 28 -18 62 16
rect 120 -18 154 16
rect 212 -18 246 16
rect 304 -18 338 16
rect 396 -18 430 16
rect 488 -18 522 16
rect 580 -18 614 16
rect 672 -18 706 16
rect 764 -18 798 16
rect 856 -18 890 16
rect 948 -18 982 16
rect 1040 -18 1074 16
rect 1132 -18 1166 16
rect 1224 -18 1258 16
rect 1316 -18 1350 16
rect 1408 -18 1442 16
rect 1500 -18 1534 16
rect 1592 -18 1626 16
rect 1684 -18 1718 16
rect 1776 -18 1810 16
rect 1868 -18 1902 16
<< metal1 >>
rect 0 560 1932 592
rect 0 526 28 560
rect 62 526 120 560
rect 154 526 212 560
rect 246 526 304 560
rect 338 526 396 560
rect 430 526 488 560
rect 522 526 580 560
rect 614 526 672 560
rect 706 526 764 560
rect 798 526 856 560
rect 890 526 948 560
rect 982 526 1040 560
rect 1074 526 1132 560
rect 1166 526 1224 560
rect 1258 526 1316 560
rect 1350 526 1408 560
rect 1442 526 1500 560
rect 1534 526 1592 560
rect 1626 526 1684 560
rect 1718 526 1776 560
rect 1810 526 1868 560
rect 1902 526 1932 560
rect 0 520 1932 526
rect 150 456 208 462
rect 150 422 162 456
rect 196 454 208 456
rect 290 454 296 466
rect 196 426 296 454
rect 196 422 216 426
rect 150 416 216 422
rect 290 414 296 426
rect 348 414 354 466
rect 1318 456 1376 462
rect 1318 422 1330 456
rect 1364 454 1376 456
rect 1518 456 1576 462
rect 1364 422 1384 454
rect 1318 416 1384 422
rect 390 400 448 406
rect 390 366 402 400
rect 436 398 448 400
rect 436 366 480 398
rect 390 360 480 366
rect 50 302 56 354
rect 108 302 114 354
rect 242 302 248 354
rect 300 350 306 354
rect 300 344 352 350
rect 300 310 306 344
rect 340 310 352 344
rect 452 314 480 360
rect 634 358 640 410
rect 692 398 698 410
rect 802 398 808 410
rect 860 406 866 410
rect 860 400 888 406
rect 692 370 808 398
rect 692 358 698 370
rect 802 358 808 370
rect 876 366 888 400
rect 860 360 888 366
rect 860 358 866 360
rect 300 304 352 310
rect 300 302 306 304
rect 68 118 96 302
rect 380 286 480 314
rect 542 344 600 350
rect 542 310 554 344
rect 588 310 600 344
rect 542 304 600 310
rect 242 190 248 242
rect 300 238 306 242
rect 300 232 352 238
rect 300 198 306 232
rect 340 198 352 232
rect 300 192 352 198
rect 300 190 306 192
rect 380 130 408 286
rect 556 242 584 304
rect 796 298 1312 314
rect 796 294 856 298
rect 782 288 856 294
rect 782 254 794 288
rect 828 254 856 288
rect 782 248 856 254
rect 850 246 856 248
rect 908 294 1312 298
rect 908 288 1328 294
rect 908 286 1282 288
rect 908 246 914 286
rect 1270 254 1282 286
rect 1316 254 1328 288
rect 1270 248 1328 254
rect 486 238 492 242
rect 438 232 492 238
rect 438 198 450 232
rect 484 198 492 232
rect 438 192 492 198
rect 486 190 492 192
rect 544 190 584 242
rect 682 190 688 242
rect 740 190 746 242
rect 1050 190 1056 242
rect 1108 238 1114 242
rect 1108 232 1136 238
rect 1124 198 1136 232
rect 1108 192 1136 198
rect 1108 190 1114 192
rect 1170 190 1176 242
rect 1228 190 1234 242
rect 150 120 208 126
rect 150 118 162 120
rect 68 90 162 118
rect 150 86 162 90
rect 196 86 208 120
rect 150 80 208 86
rect 338 78 344 130
rect 396 90 408 130
rect 556 118 584 190
rect 778 134 784 186
rect 836 174 842 186
rect 1356 182 1384 416
rect 1518 422 1530 456
rect 1564 422 1576 456
rect 1518 410 1576 422
rect 1514 358 1520 410
rect 1572 358 1578 410
rect 1480 298 1800 314
rect 1480 294 1784 298
rect 1414 288 1784 294
rect 1836 294 1842 298
rect 1836 288 1864 294
rect 1414 254 1426 288
rect 1460 286 1784 288
rect 1460 258 1508 286
rect 1772 258 1784 286
rect 1460 254 1472 258
rect 1414 248 1472 254
rect 1778 246 1784 258
rect 1852 254 1864 288
rect 1836 248 1864 254
rect 1836 246 1842 248
rect 1538 190 1544 242
rect 1596 238 1602 242
rect 1596 232 1632 238
rect 1612 198 1632 232
rect 1596 190 1632 198
rect 1662 232 1720 238
rect 1662 198 1674 232
rect 1708 230 1720 232
rect 1708 202 1752 230
rect 1708 198 1848 202
rect 1662 192 1848 198
rect 878 176 936 182
rect 878 174 890 176
rect 836 146 890 174
rect 836 134 842 146
rect 878 142 890 146
rect 924 142 936 176
rect 1356 176 1424 182
rect 1356 174 1378 176
rect 1284 146 1378 174
rect 1284 142 1312 146
rect 878 136 936 142
rect 992 130 1312 142
rect 1366 142 1378 146
rect 1412 142 1424 176
rect 1366 136 1424 142
rect 1604 142 1632 190
rect 1724 186 1848 192
rect 1724 174 1808 186
rect 638 120 696 126
rect 638 118 650 120
rect 556 90 650 118
rect 396 78 402 90
rect 638 86 650 90
rect 684 86 696 120
rect 638 80 696 86
rect 974 78 980 130
rect 1032 120 1312 130
rect 1032 86 1042 120
rect 1076 114 1312 120
rect 1076 86 1088 114
rect 1032 80 1088 86
rect 1032 78 1038 80
rect 1462 78 1468 130
rect 1520 126 1526 130
rect 1520 120 1576 126
rect 1520 86 1530 120
rect 1564 86 1576 120
rect 1604 118 1656 142
rect 1802 134 1808 174
rect 1860 134 1866 186
rect 1710 120 1768 126
rect 1710 118 1722 120
rect 1604 114 1722 118
rect 1628 90 1722 114
rect 1520 80 1576 86
rect 1710 86 1722 90
rect 1756 86 1768 120
rect 1710 80 1768 86
rect 1520 78 1526 80
rect 0 16 1932 22
rect 0 -18 28 16
rect 62 -18 120 16
rect 154 -18 212 16
rect 246 -18 304 16
rect 338 -18 396 16
rect 430 -18 488 16
rect 522 -18 580 16
rect 614 -18 672 16
rect 706 -18 764 16
rect 798 -18 856 16
rect 890 -18 948 16
rect 982 -18 1040 16
rect 1074 -18 1132 16
rect 1166 -18 1224 16
rect 1258 -18 1316 16
rect 1350 -18 1408 16
rect 1442 -18 1500 16
rect 1534 -18 1592 16
rect 1626 -18 1684 16
rect 1718 -18 1776 16
rect 1810 -18 1868 16
rect 1902 -18 1932 16
rect 0 -48 1932 -18
<< via1 >>
rect 296 414 348 466
rect 56 344 108 354
rect 56 310 66 344
rect 66 310 100 344
rect 100 310 108 344
rect 56 302 108 310
rect 248 302 300 354
rect 640 400 692 410
rect 640 366 650 400
rect 650 366 684 400
rect 684 366 692 400
rect 808 400 860 410
rect 640 358 692 366
rect 808 366 842 400
rect 842 366 860 400
rect 808 358 860 366
rect 248 190 300 242
rect 856 246 908 298
rect 492 190 544 242
rect 688 232 740 242
rect 688 198 698 232
rect 698 198 732 232
rect 732 198 740 232
rect 688 190 740 198
rect 1056 232 1108 242
rect 1056 198 1090 232
rect 1090 198 1108 232
rect 1056 190 1108 198
rect 1176 232 1228 242
rect 1176 198 1186 232
rect 1186 198 1220 232
rect 1220 198 1228 232
rect 1176 190 1228 198
rect 344 120 396 130
rect 344 86 354 120
rect 354 86 388 120
rect 388 86 396 120
rect 784 134 836 186
rect 1520 358 1572 410
rect 1784 288 1836 298
rect 1784 254 1818 288
rect 1818 254 1836 288
rect 1784 246 1836 254
rect 1544 232 1596 242
rect 1544 198 1578 232
rect 1578 198 1596 232
rect 1544 190 1596 198
rect 344 78 396 86
rect 980 78 1032 130
rect 1468 78 1520 130
rect 1808 134 1860 186
<< metal2 >>
rect 212 500 944 528
rect 54 356 110 365
rect 212 364 240 500
rect 296 466 348 472
rect 348 426 632 454
rect 296 408 348 414
rect 604 416 632 426
rect 604 410 692 416
rect 604 370 640 410
rect 212 354 302 364
rect 212 314 248 354
rect 54 290 110 300
rect 246 302 248 314
rect 300 302 302 354
rect 640 352 692 358
rect 796 410 860 416
rect 796 358 808 410
rect 796 352 860 358
rect 916 364 944 500
rect 978 468 1034 477
rect 1194 454 1630 476
rect 1034 444 1630 454
rect 1034 426 1222 444
rect 978 402 1034 412
rect 1520 410 1572 416
rect 1362 364 1422 365
rect 916 356 1422 364
rect 246 290 302 302
rect 504 253 584 286
rect 504 248 598 253
rect 248 242 300 248
rect 492 244 598 248
rect 492 242 542 244
rect 300 202 456 230
rect 248 184 300 190
rect 342 132 398 141
rect 342 66 398 76
rect 428 72 456 202
rect 492 188 542 190
rect 492 184 598 188
rect 542 178 598 184
rect 686 244 742 253
rect 796 192 824 352
rect 916 336 1366 356
rect 856 298 908 304
rect 1520 352 1572 358
rect 1520 342 1560 352
rect 1422 314 1560 342
rect 1366 290 1422 300
rect 908 253 920 286
rect 908 246 934 253
rect 856 244 934 246
rect 856 240 878 244
rect 686 178 742 188
rect 784 186 836 192
rect 878 178 934 188
rect 1054 244 1110 253
rect 1054 178 1110 188
rect 1176 242 1228 248
rect 1176 184 1228 190
rect 784 128 836 134
rect 980 130 1032 136
rect 980 72 1032 78
rect 428 44 1020 72
rect 1188 44 1216 184
rect 1390 178 1446 252
rect 1404 44 1432 178
rect 1480 136 1508 314
rect 1600 248 1630 444
rect 1782 356 1838 365
rect 1782 298 1838 300
rect 1782 290 1784 298
rect 1544 242 1630 248
rect 1596 220 1630 242
rect 1836 290 1838 298
rect 1784 240 1836 246
rect 1544 184 1596 190
rect 1686 210 1742 220
rect 1628 154 1686 174
rect 1808 186 1860 192
rect 1742 154 1808 174
rect 1628 146 1808 154
rect 1468 130 1520 136
rect 1468 72 1520 78
rect 1628 44 1656 146
rect 1808 128 1860 134
rect 1188 16 1656 44
<< via2 >>
rect 54 354 110 356
rect 54 302 56 354
rect 56 302 108 354
rect 108 302 110 354
rect 54 300 110 302
rect 978 412 1034 468
rect 542 242 598 244
rect 342 130 398 132
rect 342 78 344 130
rect 344 78 396 130
rect 396 78 398 130
rect 342 76 398 78
rect 542 190 544 242
rect 544 190 598 242
rect 542 188 598 190
rect 686 242 742 244
rect 686 190 688 242
rect 688 190 740 242
rect 740 190 742 242
rect 1366 300 1422 356
rect 686 188 742 190
rect 878 188 934 244
rect 1054 242 1110 244
rect 1054 190 1056 242
rect 1056 190 1108 242
rect 1108 190 1110 242
rect 1054 188 1110 190
rect 1782 300 1838 356
rect 1686 154 1742 210
<< metal3 >>
rect 973 470 1040 474
rect 732 468 1040 470
rect 732 412 978 468
rect 1034 412 1040 468
rect 732 410 1040 412
rect 49 356 116 361
rect 49 300 54 356
rect 110 300 116 356
rect 49 214 116 300
rect 538 249 604 328
rect 732 249 792 410
rect 973 406 1040 410
rect 1361 356 1428 361
rect 1778 360 1844 440
rect 1361 300 1366 356
rect 1422 300 1428 356
rect 1361 296 1428 300
rect 537 244 604 249
rect 338 135 404 216
rect 537 188 542 244
rect 598 188 604 244
rect 537 182 604 188
rect 681 244 792 249
rect 681 188 686 244
rect 742 188 792 244
rect 681 186 792 188
rect 873 244 940 249
rect 873 188 878 244
rect 934 188 940 244
rect 681 182 748 186
rect 873 183 940 188
rect 1049 244 1116 249
rect 1049 188 1054 244
rect 1110 188 1116 244
rect 1362 214 1428 296
rect 1777 356 1844 360
rect 1777 300 1782 356
rect 1838 300 1844 356
rect 1777 294 1844 300
rect 1049 185 1116 188
rect 337 132 404 135
rect 337 76 342 132
rect 398 76 404 132
rect 874 102 940 183
rect 1050 102 1116 185
rect 1681 210 1748 216
rect 1681 154 1686 210
rect 1742 154 1748 210
rect 1681 146 1748 154
rect 337 70 404 76
rect 1682 70 1748 146
<< labels >>
flabel nwell s 1496 526 1530 560 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 1008 526 1042 560 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 520 526 554 560 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 32 526 66 560 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel pwell s 1496 -16 1530 16 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 1008 -16 1042 16 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 520 -16 554 16 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 32 -16 66 16 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel comment s 0 0 0 0 0 FreeSans 100 0 0 0 scs130hd_mpr2ea_8
rlabel metal3 s 1778 294 1844 440 4 B0
port 3 nsew
rlabel metal3 s 874 102 940 248 4 A1
port 4 nsew
rlabel metal3 s 50 214 116 360 4 R2
port 5 nsew
rlabel metal3 s 1682 70 1748 216 4 A0
port 6 nsew
rlabel metal3 s 1362 214 1428 360 4 R0
port 7 nsew
rlabel metal3 s 538 182 604 328 4 R3
port 8 nsew
rlabel metal3 s 1050 102 1116 248 4 B1
port 9 nsew
rlabel metal3 s 338 70 404 216 4 R1
port 10 nsew
flabel metal1 s 30 526 64 560 0 FreeSans 100 0 0 0 vpwr
port 11 nsew
flabel metal1 s 30 -16 64 16 0 FreeSans 100 0 0 0 vgnd
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 1932 544
<< end >>
