magic
tech sky130A
magscale 1 2
timestamp 1707852631
<< viali >>
rect 305066 490025 305100 490059
rect 297400 472481 297434 472515
rect 299182 471053 299216 471087
rect 302767 471053 302801 471087
rect 306352 471053 306386 471087
rect 313522 471053 313556 471087
rect 302488 428961 302522 428995
rect 296907 409445 296941 409479
rect 297354 388433 297388 388467
rect 303019 387005 303053 387039
rect 307801 366333 307835 366367
rect 296695 346477 296729 346511
rect 307808 345049 307842 345083
rect 301920 324037 301954 324071
rect 298986 282013 299020 282047
rect 302303 282013 302337 282047
rect 305620 282013 305654 282047
rect 299317 262429 299351 262463
rect 302484 261001 302518 261035
rect 302125 240465 302159 240499
rect 308655 240465 308689 240499
rect 297353 220473 297387 220507
rect 303019 219045 303053 219079
rect 296693 199325 296727 199359
<< metal1 >>
rect 296876 491656 297196 491662
rect 296876 491604 296882 491656
rect 296934 491604 296946 491656
rect 296998 491604 297010 491656
rect 297062 491604 297074 491656
rect 297126 491604 297138 491656
rect 297190 491604 297196 491656
rect 296876 491592 297196 491604
rect 296876 491540 296882 491592
rect 296934 491540 296946 491592
rect 296998 491540 297010 491592
rect 297062 491540 297074 491592
rect 297126 491540 297138 491592
rect 297190 491540 297196 491592
rect 296876 491528 297196 491540
rect 296876 491476 296882 491528
rect 296934 491476 296946 491528
rect 296998 491476 297010 491528
rect 297062 491476 297074 491528
rect 297126 491476 297138 491528
rect 297190 491476 297196 491528
rect 296876 491464 297196 491476
rect 296876 491412 296882 491464
rect 296934 491412 296946 491464
rect 296998 491412 297010 491464
rect 297062 491412 297074 491464
rect 297126 491412 297138 491464
rect 297190 491412 297196 491464
rect 296876 491400 297196 491412
rect 296876 491348 296882 491400
rect 296934 491348 296946 491400
rect 296998 491348 297010 491400
rect 297062 491348 297074 491400
rect 297126 491348 297138 491400
rect 297190 491348 297196 491400
rect 296876 491342 297196 491348
rect 303876 491656 304196 491662
rect 303876 491604 303882 491656
rect 303934 491604 303946 491656
rect 303998 491604 304010 491656
rect 304062 491604 304074 491656
rect 304126 491604 304138 491656
rect 304190 491604 304196 491656
rect 303876 491592 304196 491604
rect 303876 491540 303882 491592
rect 303934 491540 303946 491592
rect 303998 491540 304010 491592
rect 304062 491540 304074 491592
rect 304126 491540 304138 491592
rect 304190 491540 304196 491592
rect 303876 491528 304196 491540
rect 303876 491476 303882 491528
rect 303934 491476 303946 491528
rect 303998 491476 304010 491528
rect 304062 491476 304074 491528
rect 304126 491476 304138 491528
rect 304190 491476 304196 491528
rect 303876 491464 304196 491476
rect 303876 491412 303882 491464
rect 303934 491412 303946 491464
rect 303998 491412 304010 491464
rect 304062 491412 304074 491464
rect 304126 491412 304138 491464
rect 304190 491412 304196 491464
rect 303876 491400 304196 491412
rect 303876 491348 303882 491400
rect 303934 491348 303946 491400
rect 303998 491348 304010 491400
rect 304062 491348 304074 491400
rect 304126 491348 304138 491400
rect 304190 491348 304196 491400
rect 303876 491342 304196 491348
rect 310876 491656 311196 491662
rect 310876 491604 310882 491656
rect 310934 491604 310946 491656
rect 310998 491604 311010 491656
rect 311062 491604 311074 491656
rect 311126 491604 311138 491656
rect 311190 491604 311196 491656
rect 310876 491592 311196 491604
rect 310876 491540 310882 491592
rect 310934 491540 310946 491592
rect 310998 491540 311010 491592
rect 311062 491540 311074 491592
rect 311126 491540 311138 491592
rect 311190 491540 311196 491592
rect 310876 491528 311196 491540
rect 310876 491476 310882 491528
rect 310934 491476 310946 491528
rect 310998 491476 311010 491528
rect 311062 491476 311074 491528
rect 311126 491476 311138 491528
rect 311190 491476 311196 491528
rect 310876 491464 311196 491476
rect 310876 491412 310882 491464
rect 310934 491412 310946 491464
rect 310998 491412 311010 491464
rect 311062 491412 311074 491464
rect 311126 491412 311138 491464
rect 311190 491412 311196 491464
rect 310876 491400 311196 491412
rect 310876 491348 310882 491400
rect 310934 491348 310946 491400
rect 310998 491348 311010 491400
rect 311062 491348 311074 491400
rect 311126 491348 311138 491400
rect 311190 491348 311196 491400
rect 310876 491342 311196 491348
rect 296996 490859 297048 490865
rect 292482 490696 292488 490748
rect 292540 490736 292546 490748
rect 295168 490736 295196 490833
rect 296996 490801 297048 490807
rect 292540 490708 295196 490736
rect 292540 490696 292546 490708
rect 294874 490628 294880 490680
rect 294932 490668 294938 490680
rect 296990 490668 296996 490680
rect 294932 490640 296996 490668
rect 294932 490628 294938 490640
rect 296990 490628 296996 490640
rect 297048 490628 297054 490680
rect 295144 490548 295464 490576
rect 295144 490496 295150 490548
rect 295202 490496 295214 490548
rect 295266 490496 295278 490548
rect 295330 490496 295342 490548
rect 295394 490496 295406 490548
rect 295458 490496 295464 490548
rect 295144 490484 295464 490496
rect 295144 490432 295150 490484
rect 295202 490432 295214 490484
rect 295266 490432 295278 490484
rect 295330 490432 295342 490484
rect 295394 490432 295406 490484
rect 295458 490432 295464 490484
rect 295144 490420 295464 490432
rect 295144 490368 295150 490420
rect 295202 490368 295214 490420
rect 295266 490368 295278 490420
rect 295330 490368 295342 490420
rect 295394 490368 295406 490420
rect 295458 490368 295464 490420
rect 295144 490356 295464 490368
rect 295144 490304 295150 490356
rect 295202 490304 295214 490356
rect 295266 490304 295278 490356
rect 295330 490304 295342 490356
rect 295394 490304 295406 490356
rect 295458 490304 295464 490356
rect 295144 490276 295464 490304
rect 312078 490192 312084 490204
rect 307404 490164 312084 490192
rect 305086 490065 305092 490068
rect 305054 490059 305092 490065
rect 305054 490025 305066 490059
rect 305054 490019 305092 490025
rect 305086 490016 305092 490019
rect 305144 490016 305150 490068
rect 307404 489999 307432 490164
rect 312078 490152 312084 490164
rect 312136 490152 312142 490204
rect 298738 489744 298744 489796
rect 298796 489744 298802 489796
rect 308122 489676 308128 489728
rect 308180 489716 308186 489728
rect 308180 489688 308246 489716
rect 308180 489676 308186 489688
rect 301774 489603 301780 489655
rect 301832 489643 301838 489655
rect 311526 489643 311532 489655
rect 301832 489615 301898 489643
rect 311374 489615 311532 489643
rect 301832 489603 301838 489615
rect 311526 489603 311532 489615
rect 311584 489603 311590 489655
rect 303876 489484 304196 489490
rect 303876 489432 303882 489484
rect 303934 489432 303946 489484
rect 303998 489432 304010 489484
rect 304062 489432 304074 489484
rect 304126 489432 304138 489484
rect 304190 489432 304196 489484
rect 303876 489420 304196 489432
rect 303876 489368 303882 489420
rect 303934 489368 303946 489420
rect 303998 489368 304010 489420
rect 304062 489368 304074 489420
rect 304126 489368 304138 489420
rect 304190 489368 304196 489420
rect 303876 489356 304196 489368
rect 303876 489304 303882 489356
rect 303934 489304 303946 489356
rect 303998 489304 304010 489356
rect 304062 489304 304074 489356
rect 304126 489304 304138 489356
rect 304190 489304 304196 489356
rect 303876 489292 304196 489304
rect 303876 489240 303882 489292
rect 303934 489240 303946 489292
rect 303998 489240 304010 489292
rect 304062 489240 304074 489292
rect 304126 489240 304138 489292
rect 304190 489240 304196 489292
rect 303876 489228 304196 489240
rect 303876 489176 303882 489228
rect 303934 489176 303946 489228
rect 303998 489176 304010 489228
rect 304062 489176 304074 489228
rect 304126 489176 304138 489228
rect 304190 489176 304196 489228
rect 303876 489170 304196 489176
rect 310876 489484 311196 489490
rect 310876 489432 310882 489484
rect 310934 489432 310946 489484
rect 310998 489432 311010 489484
rect 311062 489432 311074 489484
rect 311126 489432 311138 489484
rect 311190 489432 311196 489484
rect 310876 489420 311196 489432
rect 310876 489368 310882 489420
rect 310934 489368 310946 489420
rect 310998 489368 311010 489420
rect 311062 489368 311074 489420
rect 311126 489368 311138 489420
rect 311190 489368 311196 489420
rect 310876 489356 311196 489368
rect 310876 489304 310882 489356
rect 310934 489304 310946 489356
rect 310998 489304 311010 489356
rect 311062 489304 311074 489356
rect 311126 489304 311138 489356
rect 311190 489304 311196 489356
rect 310876 489292 311196 489304
rect 310876 489240 310882 489292
rect 310934 489240 310946 489292
rect 310998 489240 311010 489292
rect 311062 489240 311074 489292
rect 311126 489240 311138 489292
rect 311190 489240 311196 489292
rect 310876 489228 311196 489240
rect 310876 489176 310882 489228
rect 310934 489176 310946 489228
rect 310998 489176 311010 489228
rect 311062 489176 311074 489228
rect 311126 489176 311138 489228
rect 311190 489176 311196 489228
rect 310876 489170 311196 489176
rect 296876 473116 297196 473122
rect 296876 473064 296882 473116
rect 296934 473064 296946 473116
rect 296998 473064 297010 473116
rect 297062 473064 297074 473116
rect 297126 473064 297138 473116
rect 297190 473064 297196 473116
rect 296876 473052 297196 473064
rect 296876 473000 296882 473052
rect 296934 473000 296946 473052
rect 296998 473000 297010 473052
rect 297062 473000 297074 473052
rect 297126 473000 297138 473052
rect 297190 473000 297196 473052
rect 296876 472988 297196 473000
rect 296876 472936 296882 472988
rect 296934 472936 296946 472988
rect 296998 472936 297010 472988
rect 297062 472936 297074 472988
rect 297126 472936 297138 472988
rect 297190 472936 297196 472988
rect 296876 472924 297196 472936
rect 296876 472872 296882 472924
rect 296934 472872 296946 472924
rect 296998 472872 297010 472924
rect 297062 472872 297074 472924
rect 297126 472872 297138 472924
rect 297190 472872 297196 472924
rect 296876 472860 297196 472872
rect 296876 472808 296882 472860
rect 296934 472808 296946 472860
rect 296998 472808 297010 472860
rect 297062 472808 297074 472860
rect 297126 472808 297138 472860
rect 297190 472808 297196 472860
rect 296876 472802 297196 472808
rect 303876 473116 304196 473122
rect 303876 473064 303882 473116
rect 303934 473064 303946 473116
rect 303998 473064 304010 473116
rect 304062 473064 304074 473116
rect 304126 473064 304138 473116
rect 304190 473064 304196 473116
rect 303876 473052 304196 473064
rect 303876 473000 303882 473052
rect 303934 473000 303946 473052
rect 303998 473000 304010 473052
rect 304062 473000 304074 473052
rect 304126 473000 304138 473052
rect 304190 473000 304196 473052
rect 303876 472988 304196 473000
rect 303876 472936 303882 472988
rect 303934 472936 303946 472988
rect 303998 472936 304010 472988
rect 304062 472936 304074 472988
rect 304126 472936 304138 472988
rect 304190 472936 304196 472988
rect 303876 472924 304196 472936
rect 303876 472872 303882 472924
rect 303934 472872 303946 472924
rect 303998 472872 304010 472924
rect 304062 472872 304074 472924
rect 304126 472872 304138 472924
rect 304190 472872 304196 472924
rect 303876 472860 304196 472872
rect 303876 472808 303882 472860
rect 303934 472808 303946 472860
rect 303998 472808 304010 472860
rect 304062 472808 304074 472860
rect 304126 472808 304138 472860
rect 304190 472808 304196 472860
rect 303876 472802 304196 472808
rect 310876 473116 311196 473122
rect 310876 473064 310882 473116
rect 310934 473064 310946 473116
rect 310998 473064 311010 473116
rect 311062 473064 311074 473116
rect 311126 473064 311138 473116
rect 311190 473064 311196 473116
rect 310876 473052 311196 473064
rect 310876 473000 310882 473052
rect 310934 473000 310946 473052
rect 310998 473000 311010 473052
rect 311062 473000 311074 473052
rect 311126 473000 311138 473052
rect 311190 473000 311196 473052
rect 310876 472988 311196 473000
rect 310876 472936 310882 472988
rect 310934 472936 310946 472988
rect 310998 472936 311010 472988
rect 311062 472936 311074 472988
rect 311126 472936 311138 472988
rect 311190 472936 311196 472988
rect 310876 472924 311196 472936
rect 310876 472872 310882 472924
rect 310934 472872 310946 472924
rect 310998 472872 311010 472924
rect 311062 472872 311074 472924
rect 311126 472872 311138 472924
rect 311190 472872 311196 472924
rect 310876 472860 311196 472872
rect 310876 472808 310882 472860
rect 310934 472808 310946 472860
rect 310998 472808 311010 472860
rect 311062 472808 311074 472860
rect 311126 472808 311138 472860
rect 311190 472808 311196 472860
rect 310876 472802 311196 472808
rect 294874 472540 294880 472592
rect 294932 472580 294938 472592
rect 295242 472580 295248 472592
rect 294932 472552 295248 472580
rect 294932 472540 294938 472552
rect 295242 472540 295248 472552
rect 295300 472580 295306 472592
rect 295300 472552 297404 472580
rect 295300 472540 295306 472552
rect 297376 472521 297404 472552
rect 297376 472515 297446 472521
rect 297376 472484 297400 472515
rect 297388 472481 297400 472484
rect 297434 472481 297446 472515
rect 297388 472475 297446 472481
rect 292482 472336 292488 472388
rect 292540 472376 292546 472388
rect 292540 472348 295104 472376
rect 292540 472336 292546 472348
rect 295076 472307 295104 472348
rect 309140 472319 309192 472325
rect 295076 472279 295182 472307
rect 309140 472261 309192 472267
rect 302144 472015 302464 472036
rect 302144 471963 302150 472015
rect 302202 471963 302214 472015
rect 302266 471963 302278 472015
rect 302330 471963 302342 472015
rect 302394 471963 302406 472015
rect 302458 471963 302464 472015
rect 302144 471951 302464 471963
rect 302144 471899 302150 471951
rect 302202 471899 302214 471951
rect 302266 471899 302278 471951
rect 302330 471899 302342 471951
rect 302394 471899 302406 471951
rect 302458 471899 302464 471951
rect 302144 471887 302464 471899
rect 302144 471835 302150 471887
rect 302202 471835 302214 471887
rect 302266 471835 302278 471887
rect 302330 471835 302342 471887
rect 302394 471835 302406 471887
rect 302458 471835 302464 471887
rect 302144 471823 302464 471835
rect 302144 471771 302150 471823
rect 302202 471771 302214 471823
rect 302266 471771 302278 471823
rect 302330 471771 302342 471823
rect 302394 471771 302406 471823
rect 302458 471771 302464 471823
rect 302144 471759 302464 471771
rect 302144 471707 302150 471759
rect 302202 471707 302214 471759
rect 302266 471707 302278 471759
rect 302330 471707 302342 471759
rect 302394 471707 302406 471759
rect 302458 471707 302464 471759
rect 302144 471686 302464 471707
rect 309144 472015 309464 472036
rect 309144 471963 309150 472015
rect 309202 471963 309214 472015
rect 309266 471963 309278 472015
rect 309330 471963 309342 472015
rect 309394 471963 309406 472015
rect 309458 471963 309464 472015
rect 309144 471951 309464 471963
rect 309144 471899 309150 471951
rect 309202 471899 309214 471951
rect 309266 471899 309278 471951
rect 309330 471899 309342 471951
rect 309394 471899 309406 471951
rect 309458 471899 309464 471951
rect 309144 471887 309464 471899
rect 309144 471835 309150 471887
rect 309202 471835 309214 471887
rect 309266 471835 309278 471887
rect 309330 471835 309342 471887
rect 309394 471835 309406 471887
rect 309458 471835 309464 471887
rect 309144 471823 309464 471835
rect 309144 471771 309150 471823
rect 309202 471771 309214 471823
rect 309266 471771 309278 471823
rect 309330 471771 309342 471823
rect 309394 471771 309406 471823
rect 309458 471771 309464 471823
rect 309144 471759 309464 471771
rect 309144 471707 309150 471759
rect 309202 471707 309214 471759
rect 309266 471707 309278 471759
rect 309330 471707 309342 471759
rect 309394 471707 309406 471759
rect 309458 471707 309464 471759
rect 309144 471686 309464 471707
rect 313734 471248 313740 471300
rect 313792 471248 313798 471300
rect 313752 471096 313780 471248
rect 299170 471087 299228 471093
rect 299170 471053 299182 471087
rect 299216 471084 299228 471087
rect 299290 471084 299296 471096
rect 299216 471056 299296 471084
rect 299216 471053 299228 471056
rect 299170 471047 299228 471053
rect 299290 471044 299296 471056
rect 299348 471044 299354 471096
rect 302755 471087 302813 471093
rect 302755 471053 302767 471087
rect 302801 471084 302813 471087
rect 302878 471084 302884 471096
rect 302801 471056 302884 471084
rect 302801 471053 302813 471056
rect 302755 471047 302813 471053
rect 302878 471044 302884 471056
rect 302936 471044 302942 471096
rect 306340 471087 306398 471093
rect 306340 471053 306352 471087
rect 306386 471084 306398 471087
rect 306466 471084 306472 471096
rect 306386 471056 306472 471084
rect 306386 471053 306398 471056
rect 306340 471047 306398 471053
rect 306466 471044 306472 471056
rect 306524 471044 306530 471096
rect 313510 471087 313568 471093
rect 313510 471053 313522 471087
rect 313556 471084 313568 471087
rect 313642 471084 313648 471096
rect 313556 471056 313648 471084
rect 313556 471053 313568 471056
rect 313510 471047 313568 471053
rect 313642 471044 313648 471056
rect 313700 471044 313706 471096
rect 313734 471044 313740 471096
rect 313792 471044 313798 471096
rect 296876 452076 297196 452091
rect 296876 452024 296882 452076
rect 296934 452024 296946 452076
rect 296998 452024 297010 452076
rect 297062 452024 297074 452076
rect 297126 452024 297138 452076
rect 297190 452024 297196 452076
rect 296876 452012 297196 452024
rect 296876 451960 296882 452012
rect 296934 451960 296946 452012
rect 296998 451960 297010 452012
rect 297062 451960 297074 452012
rect 297126 451960 297138 452012
rect 297190 451960 297196 452012
rect 296876 451948 297196 451960
rect 296876 451896 296882 451948
rect 296934 451896 296946 451948
rect 296998 451896 297010 451948
rect 297062 451896 297074 451948
rect 297126 451896 297138 451948
rect 297190 451896 297196 451948
rect 296876 451884 297196 451896
rect 296876 451832 296882 451884
rect 296934 451832 296946 451884
rect 296998 451832 297010 451884
rect 297062 451832 297074 451884
rect 297126 451832 297138 451884
rect 297190 451832 297196 451884
rect 296876 451820 297196 451832
rect 296876 451768 296882 451820
rect 296934 451768 296946 451820
rect 296998 451768 297010 451820
rect 297062 451768 297074 451820
rect 297126 451768 297138 451820
rect 297190 451768 297196 451820
rect 296876 451756 297196 451768
rect 296876 451704 296882 451756
rect 296934 451704 296946 451756
rect 296998 451704 297010 451756
rect 297062 451704 297074 451756
rect 297126 451704 297138 451756
rect 297190 451704 297196 451756
rect 296876 451692 297196 451704
rect 296876 451640 296882 451692
rect 296934 451640 296946 451692
rect 296998 451640 297010 451692
rect 297062 451640 297074 451692
rect 297126 451640 297138 451692
rect 297190 451640 297196 451692
rect 296876 451628 297196 451640
rect 296876 451576 296882 451628
rect 296934 451576 296946 451628
rect 296998 451576 297010 451628
rect 297062 451576 297074 451628
rect 297126 451576 297138 451628
rect 297190 451576 297196 451628
rect 296876 451564 297196 451576
rect 296876 451512 296882 451564
rect 296934 451512 296946 451564
rect 296998 451512 297010 451564
rect 297062 451512 297074 451564
rect 297126 451512 297138 451564
rect 297190 451512 297196 451564
rect 296876 451500 297196 451512
rect 296876 451448 296882 451500
rect 296934 451448 296946 451500
rect 296998 451448 297010 451500
rect 297062 451448 297074 451500
rect 297126 451448 297138 451500
rect 297190 451448 297196 451500
rect 296876 451436 297196 451448
rect 296876 451384 296882 451436
rect 296934 451384 296946 451436
rect 296998 451384 297010 451436
rect 297062 451384 297074 451436
rect 297126 451384 297138 451436
rect 297190 451384 297196 451436
rect 292482 451324 292488 451376
rect 292540 451324 292546 451376
rect 296876 451372 297196 451384
rect 292500 451296 292528 451324
rect 296876 451320 296882 451372
rect 296934 451320 296946 451372
rect 296998 451320 297010 451372
rect 297062 451320 297074 451372
rect 297126 451320 297138 451372
rect 297190 451320 297196 451372
rect 296876 451308 297196 451320
rect 292500 451276 295012 451296
rect 292500 451268 295274 451276
rect 294984 451248 295274 451268
rect 295628 451249 295918 451277
rect 296876 451256 296882 451308
rect 296934 451256 296946 451308
rect 296998 451256 297010 451308
rect 297062 451256 297074 451308
rect 297126 451256 297138 451308
rect 297190 451256 297196 451308
rect 295242 451120 295248 451172
rect 295300 451160 295306 451172
rect 295628 451160 295656 451249
rect 296876 451241 297196 451256
rect 303876 452076 304196 452091
rect 303876 452024 303882 452076
rect 303934 452024 303946 452076
rect 303998 452024 304010 452076
rect 304062 452024 304074 452076
rect 304126 452024 304138 452076
rect 304190 452024 304196 452076
rect 303876 452012 304196 452024
rect 303876 451960 303882 452012
rect 303934 451960 303946 452012
rect 303998 451960 304010 452012
rect 304062 451960 304074 452012
rect 304126 451960 304138 452012
rect 304190 451960 304196 452012
rect 303876 451948 304196 451960
rect 303876 451896 303882 451948
rect 303934 451896 303946 451948
rect 303998 451896 304010 451948
rect 304062 451896 304074 451948
rect 304126 451896 304138 451948
rect 304190 451896 304196 451948
rect 303876 451884 304196 451896
rect 303876 451832 303882 451884
rect 303934 451832 303946 451884
rect 303998 451832 304010 451884
rect 304062 451832 304074 451884
rect 304126 451832 304138 451884
rect 304190 451832 304196 451884
rect 303876 451820 304196 451832
rect 303876 451768 303882 451820
rect 303934 451768 303946 451820
rect 303998 451768 304010 451820
rect 304062 451768 304074 451820
rect 304126 451768 304138 451820
rect 304190 451768 304196 451820
rect 303876 451756 304196 451768
rect 303876 451704 303882 451756
rect 303934 451704 303946 451756
rect 303998 451704 304010 451756
rect 304062 451704 304074 451756
rect 304126 451704 304138 451756
rect 304190 451704 304196 451756
rect 303876 451692 304196 451704
rect 303876 451640 303882 451692
rect 303934 451640 303946 451692
rect 303998 451640 304010 451692
rect 304062 451640 304074 451692
rect 304126 451640 304138 451692
rect 304190 451640 304196 451692
rect 303876 451628 304196 451640
rect 303876 451576 303882 451628
rect 303934 451576 303946 451628
rect 303998 451576 304010 451628
rect 304062 451576 304074 451628
rect 304126 451576 304138 451628
rect 304190 451576 304196 451628
rect 303876 451564 304196 451576
rect 303876 451512 303882 451564
rect 303934 451512 303946 451564
rect 303998 451512 304010 451564
rect 304062 451512 304074 451564
rect 304126 451512 304138 451564
rect 304190 451512 304196 451564
rect 303876 451500 304196 451512
rect 303876 451448 303882 451500
rect 303934 451448 303946 451500
rect 303998 451448 304010 451500
rect 304062 451448 304074 451500
rect 304126 451448 304138 451500
rect 304190 451448 304196 451500
rect 303876 451436 304196 451448
rect 303876 451384 303882 451436
rect 303934 451384 303946 451436
rect 303998 451384 304010 451436
rect 304062 451384 304074 451436
rect 304126 451384 304138 451436
rect 304190 451384 304196 451436
rect 303876 451372 304196 451384
rect 303876 451320 303882 451372
rect 303934 451320 303946 451372
rect 303998 451320 304010 451372
rect 304062 451320 304074 451372
rect 304126 451320 304138 451372
rect 304190 451320 304196 451372
rect 303876 451308 304196 451320
rect 303876 451256 303882 451308
rect 303934 451256 303946 451308
rect 303998 451256 304010 451308
rect 304062 451256 304074 451308
rect 304126 451256 304138 451308
rect 304190 451256 304196 451308
rect 303876 451241 304196 451256
rect 310876 452076 311098 452091
rect 310876 452024 310897 452076
rect 310949 452024 310961 452076
rect 311013 452024 311025 452076
rect 311077 452024 311098 452076
rect 310876 452012 311098 452024
rect 310876 451960 310897 452012
rect 310949 451960 310961 452012
rect 311013 451960 311025 452012
rect 311077 451960 311098 452012
rect 310876 451948 311098 451960
rect 310876 451896 310897 451948
rect 310949 451896 310961 451948
rect 311013 451896 311025 451948
rect 311077 451896 311098 451948
rect 310876 451884 311098 451896
rect 310876 451832 310897 451884
rect 310949 451832 310961 451884
rect 311013 451832 311025 451884
rect 311077 451832 311098 451884
rect 310876 451820 311098 451832
rect 310876 451768 310897 451820
rect 310949 451768 310961 451820
rect 311013 451768 311025 451820
rect 311077 451768 311098 451820
rect 310876 451756 311098 451768
rect 310876 451704 310897 451756
rect 310949 451704 310961 451756
rect 311013 451704 311025 451756
rect 311077 451704 311098 451756
rect 310876 451692 311098 451704
rect 310876 451640 310897 451692
rect 310949 451640 310961 451692
rect 311013 451640 311025 451692
rect 311077 451640 311098 451692
rect 310876 451628 311098 451640
rect 310876 451576 310897 451628
rect 310949 451576 310961 451628
rect 311013 451576 311025 451628
rect 311077 451576 311098 451628
rect 310876 451564 311098 451576
rect 310876 451512 310897 451564
rect 310949 451512 310961 451564
rect 311013 451512 311025 451564
rect 311077 451512 311098 451564
rect 310876 451500 311098 451512
rect 310876 451448 310897 451500
rect 310949 451448 310961 451500
rect 311013 451448 311025 451500
rect 311077 451448 311098 451500
rect 310876 451436 311098 451448
rect 310876 451384 310897 451436
rect 310949 451384 310961 451436
rect 311013 451384 311025 451436
rect 311077 451384 311098 451436
rect 310876 451372 311098 451384
rect 310876 451320 310897 451372
rect 310949 451320 310961 451372
rect 311013 451320 311025 451372
rect 311077 451320 311098 451372
rect 310876 451308 311098 451320
rect 310876 451256 310897 451308
rect 310949 451256 310961 451308
rect 311013 451256 311025 451308
rect 311077 451256 311098 451308
rect 310876 451241 311098 451256
rect 295300 451132 295656 451160
rect 295300 451120 295306 451132
rect 312998 450548 313004 450560
rect 311374 450520 313004 450548
rect 312998 450508 313004 450520
rect 313056 450508 313062 450560
rect 306190 450480 306196 450492
rect 305012 450452 306196 450480
rect 305012 450443 305040 450452
rect 300854 450372 300860 450424
rect 300912 450412 300918 450424
rect 301424 450412 301452 450429
rect 304750 450415 305040 450443
rect 306190 450440 306196 450452
rect 306248 450440 306254 450492
rect 300912 450384 301452 450412
rect 300912 450372 300918 450384
rect 310876 450191 311136 450218
rect 310876 450139 310884 450191
rect 310936 450139 310948 450191
rect 311000 450139 311012 450191
rect 311064 450139 311076 450191
rect 311128 450139 311136 450191
rect 310876 450127 311136 450139
rect 310876 450075 310884 450127
rect 310936 450075 310948 450127
rect 311000 450075 311012 450127
rect 311064 450075 311076 450127
rect 311128 450075 311136 450127
rect 310876 450063 311136 450075
rect 310876 450011 310884 450063
rect 310936 450011 310948 450063
rect 311000 450011 311012 450063
rect 311064 450011 311076 450063
rect 311128 450011 311136 450063
rect 310876 449999 311136 450011
rect 310876 449947 310884 449999
rect 310936 449947 310948 449999
rect 311000 449947 311012 449999
rect 311064 449947 311076 449999
rect 311128 449947 311136 449999
rect 310876 449935 311136 449947
rect 310876 449883 310884 449935
rect 310936 449883 310948 449935
rect 311000 449883 311012 449935
rect 311064 449883 311076 449935
rect 311128 449883 311136 449935
rect 310876 449871 311136 449883
rect 310876 449819 310884 449871
rect 310936 449819 310948 449871
rect 311000 449819 311012 449871
rect 311064 449819 311076 449871
rect 311128 449819 311136 449871
rect 310876 449807 311136 449819
rect 310876 449755 310884 449807
rect 310936 449755 310948 449807
rect 311000 449755 311012 449807
rect 311064 449755 311076 449807
rect 311128 449755 311136 449807
rect 310876 449743 311136 449755
rect 310876 449691 310884 449743
rect 310936 449691 310948 449743
rect 311000 449691 311012 449743
rect 311064 449691 311076 449743
rect 311128 449691 311136 449743
rect 310876 449679 311136 449691
rect 310876 449627 310884 449679
rect 310936 449627 310948 449679
rect 311000 449627 311012 449679
rect 311064 449627 311076 449679
rect 311128 449627 311136 449679
rect 310876 449600 311136 449627
rect 292482 430244 292488 430296
rect 292540 430284 292546 430296
rect 295892 430289 295944 430295
rect 292540 430277 295012 430284
rect 292540 430256 295274 430277
rect 292540 430244 292546 430256
rect 294984 430249 295274 430256
rect 312446 430284 312452 430296
rect 312018 430256 312452 430284
rect 312446 430244 312452 430256
rect 312504 430284 312510 430296
rect 312814 430284 312820 430296
rect 312504 430256 312820 430284
rect 312504 430244 312510 430256
rect 312814 430244 312820 430256
rect 312872 430244 312878 430296
rect 295892 430231 295944 430237
rect 309144 430000 309454 430007
rect 309144 429948 309177 430000
rect 309229 429948 309241 430000
rect 309293 429948 309305 430000
rect 309357 429948 309369 430000
rect 309421 429948 309454 430000
rect 309144 429936 309454 429948
rect 309144 429884 309177 429936
rect 309229 429884 309241 429936
rect 309293 429884 309305 429936
rect 309357 429884 309369 429936
rect 309421 429884 309454 429936
rect 309144 429872 309454 429884
rect 309144 429820 309177 429872
rect 309229 429820 309241 429872
rect 309293 429820 309305 429872
rect 309357 429820 309369 429872
rect 309421 429820 309454 429872
rect 309144 429808 309454 429820
rect 309144 429756 309177 429808
rect 309229 429756 309241 429808
rect 309293 429756 309305 429808
rect 309357 429756 309369 429808
rect 309421 429756 309454 429808
rect 309144 429744 309454 429756
rect 309144 429692 309177 429744
rect 309229 429692 309241 429744
rect 309293 429692 309305 429744
rect 309357 429692 309369 429744
rect 309421 429692 309454 429744
rect 309144 429685 309454 429692
rect 301688 429455 301740 429461
rect 301688 429397 301740 429403
rect 301700 429208 301728 429397
rect 301682 429156 301688 429208
rect 301740 429156 301746 429208
rect 299020 429084 299072 429090
rect 312998 429072 313004 429084
rect 299020 429026 299072 429032
rect 305914 429020 305920 429072
rect 305972 429020 305978 429072
rect 312846 429044 313004 429072
rect 312998 429032 313004 429044
rect 313056 429032 313062 429084
rect 302510 429001 302516 429004
rect 302476 428995 302516 429001
rect 302476 428961 302488 428995
rect 302476 428955 302516 428961
rect 302510 428952 302516 428955
rect 302568 428952 302574 429004
rect 526990 421336 526996 421388
rect 527048 421376 527054 421388
rect 529198 421376 529204 421388
rect 527048 421348 529204 421376
rect 527048 421336 527054 421348
rect 529198 421336 529204 421348
rect 529256 421336 529262 421388
rect 296876 410086 297196 410092
rect 296876 410034 296882 410086
rect 296934 410034 296946 410086
rect 296998 410034 297010 410086
rect 297062 410034 297074 410086
rect 297126 410034 297138 410086
rect 297190 410034 297196 410086
rect 296876 410022 297196 410034
rect 296876 409970 296882 410022
rect 296934 409970 296946 410022
rect 296998 409970 297010 410022
rect 297062 409970 297074 410022
rect 297126 409970 297138 410022
rect 297190 409970 297196 410022
rect 296876 409958 297196 409970
rect 296876 409906 296882 409958
rect 296934 409906 296946 409958
rect 296998 409906 297010 409958
rect 297062 409906 297074 409958
rect 297126 409906 297138 409958
rect 297190 409906 297196 409958
rect 296876 409894 297196 409906
rect 296876 409842 296882 409894
rect 296934 409842 296946 409894
rect 296998 409842 297010 409894
rect 297062 409842 297074 409894
rect 297126 409842 297138 409894
rect 297190 409842 297196 409894
rect 296876 409830 297196 409842
rect 296876 409778 296882 409830
rect 296934 409778 296946 409830
rect 296998 409778 297010 409830
rect 297062 409778 297074 409830
rect 297126 409778 297138 409830
rect 297190 409778 297196 409830
rect 296876 409772 297196 409778
rect 303876 410086 304196 410092
rect 303876 410034 303882 410086
rect 303934 410034 303946 410086
rect 303998 410034 304010 410086
rect 304062 410034 304074 410086
rect 304126 410034 304138 410086
rect 304190 410034 304196 410086
rect 303876 410022 304196 410034
rect 303876 409970 303882 410022
rect 303934 409970 303946 410022
rect 303998 409970 304010 410022
rect 304062 409970 304074 410022
rect 304126 409970 304138 410022
rect 304190 409970 304196 410022
rect 303876 409958 304196 409970
rect 303876 409906 303882 409958
rect 303934 409906 303946 409958
rect 303998 409906 304010 409958
rect 304062 409906 304074 409958
rect 304126 409906 304138 409958
rect 304190 409906 304196 409958
rect 303876 409894 304196 409906
rect 303876 409842 303882 409894
rect 303934 409842 303946 409894
rect 303998 409842 304010 409894
rect 304062 409842 304074 409894
rect 304126 409842 304138 409894
rect 304190 409842 304196 409894
rect 303876 409830 304196 409842
rect 303876 409778 303882 409830
rect 303934 409778 303946 409830
rect 303998 409778 304010 409830
rect 304062 409778 304074 409830
rect 304126 409778 304138 409830
rect 304190 409778 304196 409830
rect 303876 409772 304196 409778
rect 310876 410086 311196 410092
rect 310876 410034 310882 410086
rect 310934 410034 310946 410086
rect 310998 410034 311010 410086
rect 311062 410034 311074 410086
rect 311126 410034 311138 410086
rect 311190 410034 311196 410086
rect 310876 410022 311196 410034
rect 310876 409970 310882 410022
rect 310934 409970 310946 410022
rect 310998 409970 311010 410022
rect 311062 409970 311074 410022
rect 311126 409970 311138 410022
rect 311190 409970 311196 410022
rect 310876 409958 311196 409970
rect 310876 409906 310882 409958
rect 310934 409906 310946 409958
rect 310998 409906 311010 409958
rect 311062 409906 311074 409958
rect 311126 409906 311138 409958
rect 311190 409906 311196 409958
rect 310876 409894 311196 409906
rect 310876 409842 310882 409894
rect 310934 409842 310946 409894
rect 310998 409842 311010 409894
rect 311062 409842 311074 409894
rect 311126 409842 311138 409894
rect 311190 409842 311196 409894
rect 310876 409830 311196 409842
rect 310876 409778 310882 409830
rect 310934 409778 310946 409830
rect 310998 409778 311010 409830
rect 311062 409778 311074 409830
rect 311126 409778 311138 409830
rect 311190 409778 311196 409830
rect 310876 409772 311196 409778
rect 295242 409504 295248 409556
rect 295300 409544 295306 409556
rect 295300 409516 296944 409544
rect 295300 409504 295306 409516
rect 296916 409485 296944 409516
rect 296895 409479 296953 409485
rect 296895 409445 296907 409479
rect 296941 409445 296953 409479
rect 296895 409439 296953 409445
rect 292482 409232 292488 409284
rect 292540 409272 292546 409284
rect 292540 409244 295196 409272
rect 292540 409232 292546 409244
rect 302144 409000 302464 409006
rect 302144 408948 302150 409000
rect 302202 408948 302214 409000
rect 302266 408948 302278 409000
rect 302330 408948 302342 409000
rect 302394 408948 302406 409000
rect 302458 408948 302464 409000
rect 302144 408936 302464 408948
rect 302144 408884 302150 408936
rect 302202 408884 302214 408936
rect 302266 408884 302278 408936
rect 302330 408884 302342 408936
rect 302394 408884 302406 408936
rect 302458 408884 302464 408936
rect 302144 408872 302464 408884
rect 302144 408820 302150 408872
rect 302202 408820 302214 408872
rect 302266 408820 302278 408872
rect 302330 408820 302342 408872
rect 302394 408820 302406 408872
rect 302458 408820 302464 408872
rect 302144 408808 302464 408820
rect 302144 408756 302150 408808
rect 302202 408756 302214 408808
rect 302266 408756 302278 408808
rect 302330 408756 302342 408808
rect 302394 408756 302406 408808
rect 302458 408756 302464 408808
rect 302144 408744 302464 408756
rect 302144 408692 302150 408744
rect 302202 408692 302214 408744
rect 302266 408692 302278 408744
rect 302330 408692 302342 408744
rect 302394 408692 302406 408744
rect 302458 408692 302464 408744
rect 302144 408686 302464 408692
rect 313274 408456 313280 408468
rect 311098 408428 313280 408456
rect 313274 408416 313280 408428
rect 313332 408456 313338 408468
rect 314562 408456 314568 408468
rect 313332 408428 314568 408456
rect 313332 408416 313338 408428
rect 314562 408416 314568 408428
rect 314620 408416 314626 408468
rect 311912 408048 311940 408059
rect 312170 408048 312176 408060
rect 311912 408020 312176 408048
rect 312170 408008 312176 408020
rect 312228 408008 312234 408060
rect 310876 407914 311196 407920
rect 310876 407862 310882 407914
rect 310934 407862 310946 407914
rect 310998 407862 311010 407914
rect 311062 407862 311074 407914
rect 311126 407862 311138 407914
rect 311190 407862 311196 407914
rect 310876 407850 311196 407862
rect 310876 407798 310882 407850
rect 310934 407798 310946 407850
rect 310998 407798 311010 407850
rect 311062 407798 311074 407850
rect 311126 407798 311138 407850
rect 311190 407798 311196 407850
rect 310876 407786 311196 407798
rect 310876 407734 310882 407786
rect 310934 407734 310946 407786
rect 310998 407734 311010 407786
rect 311062 407734 311074 407786
rect 311126 407734 311138 407786
rect 311190 407734 311196 407786
rect 310876 407722 311196 407734
rect 310876 407670 310882 407722
rect 310934 407670 310946 407722
rect 310998 407670 311010 407722
rect 311062 407670 311074 407722
rect 311126 407670 311138 407722
rect 311190 407670 311196 407722
rect 310876 407658 311196 407670
rect 310876 407606 310882 407658
rect 310934 407606 310946 407658
rect 310998 407606 311010 407658
rect 311062 407606 311074 407658
rect 311126 407606 311138 407658
rect 311190 407606 311196 407658
rect 310876 407600 311196 407606
rect 316862 404336 316868 404388
rect 316920 404376 316926 404388
rect 514754 404376 514760 404388
rect 316920 404348 514760 404376
rect 316920 404336 316926 404348
rect 514754 404336 514760 404348
rect 514812 404336 514818 404388
rect 296876 389087 297196 389093
rect 296876 389035 296882 389087
rect 296934 389035 296946 389087
rect 296998 389035 297010 389087
rect 297062 389035 297074 389087
rect 297126 389035 297138 389087
rect 297190 389035 297196 389087
rect 296876 389023 297196 389035
rect 296876 388971 296882 389023
rect 296934 388971 296946 389023
rect 296998 388971 297010 389023
rect 297062 388971 297074 389023
rect 297126 388971 297138 389023
rect 297190 388971 297196 389023
rect 296876 388959 297196 388971
rect 296876 388907 296882 388959
rect 296934 388907 296946 388959
rect 296998 388907 297010 388959
rect 297062 388907 297074 388959
rect 297126 388907 297138 388959
rect 297190 388907 297196 388959
rect 296876 388895 297196 388907
rect 296876 388843 296882 388895
rect 296934 388843 296946 388895
rect 296998 388843 297010 388895
rect 297062 388843 297074 388895
rect 297126 388843 297138 388895
rect 297190 388843 297196 388895
rect 296876 388831 297196 388843
rect 296876 388779 296882 388831
rect 296934 388779 296946 388831
rect 296998 388779 297010 388831
rect 297062 388779 297074 388831
rect 297126 388779 297138 388831
rect 297190 388779 297196 388831
rect 296876 388773 297196 388779
rect 303876 389087 304196 389093
rect 303876 389035 303882 389087
rect 303934 389035 303946 389087
rect 303998 389035 304010 389087
rect 304062 389035 304074 389087
rect 304126 389035 304138 389087
rect 304190 389035 304196 389087
rect 303876 389023 304196 389035
rect 303876 388971 303882 389023
rect 303934 388971 303946 389023
rect 303998 388971 304010 389023
rect 304062 388971 304074 389023
rect 304126 388971 304138 389023
rect 304190 388971 304196 389023
rect 303876 388959 304196 388971
rect 303876 388907 303882 388959
rect 303934 388907 303946 388959
rect 303998 388907 304010 388959
rect 304062 388907 304074 388959
rect 304126 388907 304138 388959
rect 304190 388907 304196 388959
rect 303876 388895 304196 388907
rect 303876 388843 303882 388895
rect 303934 388843 303946 388895
rect 303998 388843 304010 388895
rect 304062 388843 304074 388895
rect 304126 388843 304138 388895
rect 304190 388843 304196 388895
rect 303876 388831 304196 388843
rect 303876 388779 303882 388831
rect 303934 388779 303946 388831
rect 303998 388779 304010 388831
rect 304062 388779 304074 388831
rect 304126 388779 304138 388831
rect 304190 388779 304196 388831
rect 303876 388773 304196 388779
rect 310876 389087 311196 389093
rect 310876 389035 310882 389087
rect 310934 389035 310946 389087
rect 310998 389035 311010 389087
rect 311062 389035 311074 389087
rect 311126 389035 311138 389087
rect 311190 389035 311196 389087
rect 310876 389023 311196 389035
rect 310876 388971 310882 389023
rect 310934 388971 310946 389023
rect 310998 388971 311010 389023
rect 311062 388971 311074 389023
rect 311126 388971 311138 389023
rect 311190 388971 311196 389023
rect 310876 388959 311196 388971
rect 310876 388907 310882 388959
rect 310934 388907 310946 388959
rect 310998 388907 311010 388959
rect 311062 388907 311074 388959
rect 311126 388907 311138 388959
rect 311190 388907 311196 388959
rect 310876 388895 311196 388907
rect 310876 388843 310882 388895
rect 310934 388843 310946 388895
rect 310998 388843 311010 388895
rect 311062 388843 311074 388895
rect 311126 388843 311138 388895
rect 311190 388843 311196 388895
rect 310876 388831 311196 388843
rect 310876 388779 310882 388831
rect 310934 388779 310946 388831
rect 310998 388779 311010 388831
rect 311062 388779 311074 388831
rect 311126 388779 311138 388831
rect 311190 388779 311196 388831
rect 310876 388773 311196 388779
rect 295058 388492 295064 388544
rect 295116 388532 295122 388544
rect 295116 388504 297404 388532
rect 295116 388492 295122 388504
rect 292482 388424 292488 388476
rect 292540 388464 292546 388476
rect 297376 388473 297404 388504
rect 297342 388467 297404 388473
rect 292540 388436 295196 388464
rect 292540 388424 292546 388436
rect 295168 388264 295196 388436
rect 297342 388433 297354 388467
rect 297388 388436 297404 388467
rect 297388 388433 297400 388436
rect 297342 388427 297400 388433
rect 301590 388238 301596 388290
rect 301648 388238 301654 388290
rect 295144 388004 295464 388010
rect 295144 387952 295150 388004
rect 295202 387952 295214 388004
rect 295266 387952 295278 388004
rect 295330 387952 295342 388004
rect 295394 387952 295406 388004
rect 295458 387952 295464 388004
rect 295144 387940 295464 387952
rect 295144 387888 295150 387940
rect 295202 387888 295214 387940
rect 295266 387888 295278 387940
rect 295330 387888 295342 387940
rect 295394 387888 295406 387940
rect 295458 387888 295464 387940
rect 295144 387876 295464 387888
rect 295144 387824 295150 387876
rect 295202 387824 295214 387876
rect 295266 387824 295278 387876
rect 295330 387824 295342 387876
rect 295394 387824 295406 387876
rect 295458 387824 295464 387876
rect 295144 387812 295464 387824
rect 295144 387760 295150 387812
rect 295202 387760 295214 387812
rect 295266 387760 295278 387812
rect 295330 387760 295342 387812
rect 295394 387760 295406 387812
rect 295458 387760 295464 387812
rect 295144 387748 295464 387760
rect 295144 387696 295150 387748
rect 295202 387696 295214 387748
rect 295266 387696 295278 387748
rect 295330 387696 295342 387748
rect 295394 387696 295406 387748
rect 295458 387696 295464 387748
rect 295144 387690 295464 387696
rect 302144 387999 302464 388005
rect 302144 387947 302150 387999
rect 302202 387947 302214 387999
rect 302266 387947 302278 387999
rect 302330 387947 302342 387999
rect 302394 387947 302406 387999
rect 302458 387947 302464 387999
rect 302144 387935 302464 387947
rect 302144 387883 302150 387935
rect 302202 387883 302214 387935
rect 302266 387883 302278 387935
rect 302330 387883 302342 387935
rect 302394 387883 302406 387935
rect 302458 387883 302464 387935
rect 302144 387871 302464 387883
rect 302144 387819 302150 387871
rect 302202 387819 302214 387871
rect 302266 387819 302278 387871
rect 302330 387819 302342 387871
rect 302394 387819 302406 387871
rect 302458 387819 302464 387871
rect 302144 387807 302464 387819
rect 302144 387755 302150 387807
rect 302202 387755 302214 387807
rect 302266 387755 302278 387807
rect 302330 387755 302342 387807
rect 302394 387755 302406 387807
rect 302458 387755 302464 387807
rect 302144 387743 302464 387755
rect 302144 387691 302150 387743
rect 302202 387691 302214 387743
rect 302266 387691 302278 387743
rect 302330 387691 302342 387743
rect 302394 387691 302406 387743
rect 302458 387691 302464 387743
rect 302144 387685 302464 387691
rect 309144 387999 309464 388005
rect 309144 387947 309150 387999
rect 309202 387947 309214 387999
rect 309266 387947 309278 387999
rect 309330 387947 309342 387999
rect 309394 387947 309406 387999
rect 309458 387947 309464 387999
rect 309144 387935 309464 387947
rect 309144 387883 309150 387935
rect 309202 387883 309214 387935
rect 309266 387883 309278 387935
rect 309330 387883 309342 387935
rect 309394 387883 309406 387935
rect 309458 387883 309464 387935
rect 309144 387871 309464 387883
rect 309144 387819 309150 387871
rect 309202 387819 309214 387871
rect 309266 387819 309278 387871
rect 309330 387819 309342 387871
rect 309394 387819 309406 387871
rect 309458 387819 309464 387871
rect 309144 387807 309464 387819
rect 309144 387755 309150 387807
rect 309202 387755 309214 387807
rect 309266 387755 309278 387807
rect 309330 387755 309342 387807
rect 309394 387755 309406 387807
rect 309458 387755 309464 387807
rect 309144 387743 309464 387755
rect 309144 387691 309150 387743
rect 309202 387691 309214 387743
rect 309266 387691 309278 387743
rect 309330 387691 309342 387743
rect 309394 387691 309406 387743
rect 309458 387691 309464 387743
rect 309144 387685 309464 387691
rect 311040 387461 311046 387513
rect 311098 387461 311104 387513
rect 303963 387396 304021 387407
rect 303963 387344 303966 387396
rect 304018 387344 304021 387396
rect 303963 387333 304021 387344
rect 299296 387085 299348 387091
rect 306748 387085 306800 387091
rect 299296 387027 299348 387033
rect 303007 387039 303065 387045
rect 303007 387005 303019 387039
rect 303053 387036 303065 387039
rect 303154 387036 303160 387048
rect 303053 387008 303160 387036
rect 303053 387005 303065 387008
rect 303007 386999 303065 387005
rect 303154 386996 303160 387008
rect 303212 386996 303218 387048
rect 306748 387027 306800 387033
rect 310428 387085 310480 387091
rect 310428 387027 310480 387033
rect 295058 374688 295064 374740
rect 295116 374688 295122 374740
rect 295076 374536 295104 374688
rect 295058 374484 295064 374536
rect 295116 374484 295122 374536
rect 294966 370744 294972 370796
rect 295024 370784 295030 370796
rect 295242 370784 295248 370796
rect 295024 370756 295248 370784
rect 295024 370744 295030 370756
rect 295242 370744 295248 370756
rect 295300 370744 295306 370796
rect 292482 367412 292488 367464
rect 292540 367452 292546 367464
rect 292540 367424 295196 367452
rect 292540 367412 292546 367424
rect 295168 367264 295196 367424
rect 296720 367290 296772 367296
rect 296720 367232 296772 367238
rect 299756 367290 299808 367296
rect 299756 367232 299808 367238
rect 295058 367140 295064 367192
rect 295116 367180 295122 367192
rect 296714 367180 296720 367192
rect 295116 367152 296720 367180
rect 295116 367140 295122 367152
rect 296714 367140 296720 367152
rect 296772 367140 296778 367192
rect 307050 366432 307156 366443
rect 307662 366432 307668 366444
rect 307050 366415 307668 366432
rect 307128 366404 307668 366415
rect 307662 366392 307668 366404
rect 307720 366392 307726 366444
rect 307789 366367 307847 366373
rect 307789 366333 307801 366367
rect 307835 366364 307847 366367
rect 307938 366364 307944 366376
rect 307835 366336 307944 366364
rect 307835 366333 307847 366336
rect 307789 366327 307847 366333
rect 307938 366324 307944 366336
rect 307996 366324 308002 366376
rect 298652 366084 298704 366090
rect 298652 366026 298704 366032
rect 301688 366084 301740 366090
rect 301688 366026 301740 366032
rect 304724 366084 304776 366090
rect 304724 366026 304776 366032
rect 313918 364352 313924 364404
rect 313976 364392 313982 364404
rect 514754 364392 514760 364404
rect 313976 364364 514760 364392
rect 313976 364352 313982 364364
rect 514754 364352 514760 364364
rect 514812 364352 514818 364404
rect 310514 347148 310520 347200
rect 310572 347188 310578 347200
rect 311434 347188 311440 347200
rect 310572 347160 311440 347188
rect 310572 347148 310578 347160
rect 311434 347148 311440 347160
rect 311492 347148 311498 347200
rect 296876 347087 297196 347093
rect 296876 347035 296882 347087
rect 296934 347035 296946 347087
rect 296998 347035 297010 347087
rect 297062 347035 297074 347087
rect 297126 347035 297138 347087
rect 297190 347035 297196 347087
rect 296876 347023 297196 347035
rect 296876 346971 296882 347023
rect 296934 346971 296946 347023
rect 296998 346971 297010 347023
rect 297062 346971 297074 347023
rect 297126 346971 297138 347023
rect 297190 346971 297196 347023
rect 296876 346959 297196 346971
rect 296876 346907 296882 346959
rect 296934 346907 296946 346959
rect 296998 346907 297010 346959
rect 297062 346907 297074 346959
rect 297126 346907 297138 346959
rect 297190 346907 297196 346959
rect 296876 346895 297196 346907
rect 296876 346843 296882 346895
rect 296934 346843 296946 346895
rect 296998 346843 297010 346895
rect 297062 346843 297074 346895
rect 297126 346843 297138 346895
rect 297190 346843 297196 346895
rect 296876 346831 297196 346843
rect 296876 346779 296882 346831
rect 296934 346779 296946 346831
rect 296998 346779 297010 346831
rect 297062 346779 297074 346831
rect 297126 346779 297138 346831
rect 297190 346779 297196 346831
rect 296876 346773 297196 346779
rect 303876 347087 304196 347093
rect 303876 347035 303882 347087
rect 303934 347035 303946 347087
rect 303998 347035 304010 347087
rect 304062 347035 304074 347087
rect 304126 347035 304138 347087
rect 304190 347035 304196 347087
rect 303876 347023 304196 347035
rect 303876 346971 303882 347023
rect 303934 346971 303946 347023
rect 303998 346971 304010 347023
rect 304062 346971 304074 347023
rect 304126 346971 304138 347023
rect 304190 346971 304196 347023
rect 303876 346959 304196 346971
rect 303876 346907 303882 346959
rect 303934 346907 303946 346959
rect 303998 346907 304010 346959
rect 304062 346907 304074 346959
rect 304126 346907 304138 346959
rect 304190 346907 304196 346959
rect 303876 346895 304196 346907
rect 303876 346843 303882 346895
rect 303934 346843 303946 346895
rect 303998 346843 304010 346895
rect 304062 346843 304074 346895
rect 304126 346843 304138 346895
rect 304190 346843 304196 346895
rect 303876 346831 304196 346843
rect 303876 346779 303882 346831
rect 303934 346779 303946 346831
rect 303998 346779 304010 346831
rect 304062 346779 304074 346831
rect 304126 346779 304138 346831
rect 304190 346779 304196 346831
rect 303876 346773 304196 346779
rect 295150 346468 295156 346520
rect 295208 346508 295214 346520
rect 296683 346511 296741 346517
rect 296683 346508 296695 346511
rect 295208 346480 296695 346508
rect 295208 346468 295214 346480
rect 296683 346477 296695 346480
rect 296729 346477 296741 346511
rect 296683 346471 296741 346477
rect 292482 346332 292488 346384
rect 292540 346332 292546 346384
rect 292500 346304 292528 346332
rect 292500 346278 295012 346304
rect 292500 346276 295274 346278
rect 294984 346250 295274 346276
rect 302144 345985 302464 346007
rect 302144 345933 302150 345985
rect 302202 345933 302214 345985
rect 302266 345933 302278 345985
rect 302330 345933 302342 345985
rect 302394 345933 302406 345985
rect 302458 345933 302464 345985
rect 302144 345921 302464 345933
rect 302144 345869 302150 345921
rect 302202 345869 302214 345921
rect 302266 345869 302278 345921
rect 302330 345869 302342 345921
rect 302394 345869 302406 345921
rect 302458 345869 302464 345921
rect 302144 345857 302464 345869
rect 302144 345805 302150 345857
rect 302202 345805 302214 345857
rect 302266 345805 302278 345857
rect 302330 345805 302342 345857
rect 302394 345805 302406 345857
rect 302458 345805 302464 345857
rect 302144 345793 302464 345805
rect 302144 345741 302150 345793
rect 302202 345741 302214 345793
rect 302266 345741 302278 345793
rect 302330 345741 302342 345793
rect 302394 345741 302406 345793
rect 302458 345741 302464 345793
rect 302144 345729 302464 345741
rect 302144 345677 302150 345729
rect 302202 345677 302214 345729
rect 302266 345677 302278 345729
rect 302330 345677 302342 345729
rect 302394 345677 302406 345729
rect 302458 345677 302464 345729
rect 302144 345655 302464 345677
rect 309144 345985 309464 346007
rect 309144 345933 309150 345985
rect 309202 345933 309214 345985
rect 309266 345933 309278 345985
rect 309330 345933 309342 345985
rect 309394 345933 309406 345985
rect 309458 345933 309464 345985
rect 309144 345921 309464 345933
rect 309144 345869 309150 345921
rect 309202 345869 309214 345921
rect 309266 345869 309278 345921
rect 309330 345869 309342 345921
rect 309394 345869 309406 345921
rect 309458 345869 309464 345921
rect 309144 345857 309464 345869
rect 309144 345805 309150 345857
rect 309202 345805 309214 345857
rect 309266 345805 309278 345857
rect 309330 345805 309342 345857
rect 309394 345805 309406 345857
rect 309458 345805 309464 345857
rect 309144 345793 309464 345805
rect 309144 345741 309150 345793
rect 309202 345741 309214 345793
rect 309266 345741 309278 345793
rect 309330 345741 309342 345793
rect 309394 345741 309406 345793
rect 309458 345741 309464 345793
rect 309144 345729 309464 345741
rect 309144 345677 309150 345729
rect 309202 345677 309214 345729
rect 309266 345677 309278 345729
rect 309330 345677 309342 345729
rect 309394 345677 309406 345729
rect 309458 345677 309464 345729
rect 309144 345655 309464 345677
rect 298652 345084 298704 345090
rect 298652 345026 298704 345032
rect 301688 345084 301740 345090
rect 301688 345026 301740 345032
rect 304724 345084 304776 345090
rect 307796 345083 307854 345089
rect 307796 345049 307808 345083
rect 307842 345080 307854 345083
rect 307938 345080 307944 345092
rect 307842 345052 307944 345080
rect 307842 345049 307854 345052
rect 307796 345043 307854 345049
rect 307938 345040 307944 345052
rect 307996 345040 308002 345092
rect 304724 345026 304776 345032
rect 296876 326086 297196 326092
rect 296876 326034 296882 326086
rect 296934 326034 296946 326086
rect 296998 326034 297010 326086
rect 297062 326034 297074 326086
rect 297126 326034 297138 326086
rect 297190 326034 297196 326086
rect 296876 326022 297196 326034
rect 296876 325970 296882 326022
rect 296934 325970 296946 326022
rect 296998 325970 297010 326022
rect 297062 325970 297074 326022
rect 297126 325970 297138 326022
rect 297190 325970 297196 326022
rect 296876 325958 297196 325970
rect 296876 325906 296882 325958
rect 296934 325906 296946 325958
rect 296998 325906 297010 325958
rect 297062 325906 297074 325958
rect 297126 325906 297138 325958
rect 297190 325906 297196 325958
rect 296876 325894 297196 325906
rect 296876 325842 296882 325894
rect 296934 325842 296946 325894
rect 296998 325842 297010 325894
rect 297062 325842 297074 325894
rect 297126 325842 297138 325894
rect 297190 325842 297196 325894
rect 296876 325830 297196 325842
rect 296876 325778 296882 325830
rect 296934 325778 296946 325830
rect 296998 325778 297010 325830
rect 297062 325778 297074 325830
rect 297126 325778 297138 325830
rect 297190 325778 297196 325830
rect 296876 325772 297196 325778
rect 303876 326086 304196 326092
rect 303876 326034 303882 326086
rect 303934 326034 303946 326086
rect 303998 326034 304010 326086
rect 304062 326034 304074 326086
rect 304126 326034 304138 326086
rect 304190 326034 304196 326086
rect 303876 326022 304196 326034
rect 303876 325970 303882 326022
rect 303934 325970 303946 326022
rect 303998 325970 304010 326022
rect 304062 325970 304074 326022
rect 304126 325970 304138 326022
rect 304190 325970 304196 326022
rect 303876 325958 304196 325970
rect 303876 325906 303882 325958
rect 303934 325906 303946 325958
rect 303998 325906 304010 325958
rect 304062 325906 304074 325958
rect 304126 325906 304138 325958
rect 304190 325906 304196 325958
rect 303876 325894 304196 325906
rect 303876 325842 303882 325894
rect 303934 325842 303946 325894
rect 303998 325842 304010 325894
rect 304062 325842 304074 325894
rect 304126 325842 304138 325894
rect 304190 325842 304196 325894
rect 303876 325830 304196 325842
rect 303876 325778 303882 325830
rect 303934 325778 303946 325830
rect 303998 325778 304010 325830
rect 304062 325778 304074 325830
rect 304126 325778 304138 325830
rect 304190 325778 304196 325830
rect 303876 325772 304196 325778
rect 310876 326086 311196 326092
rect 310876 326034 310882 326086
rect 310934 326034 310946 326086
rect 310998 326034 311010 326086
rect 311062 326034 311074 326086
rect 311126 326034 311138 326086
rect 311190 326034 311196 326086
rect 310876 326022 311196 326034
rect 310876 325970 310882 326022
rect 310934 325970 310946 326022
rect 310998 325970 311010 326022
rect 311062 325970 311074 326022
rect 311126 325970 311138 326022
rect 311190 325970 311196 326022
rect 310876 325958 311196 325970
rect 310876 325906 310882 325958
rect 310934 325906 310946 325958
rect 310998 325906 311010 325958
rect 311062 325906 311074 325958
rect 311126 325906 311138 325958
rect 311190 325906 311196 325958
rect 310876 325894 311196 325906
rect 310876 325842 310882 325894
rect 310934 325842 310946 325894
rect 310998 325842 311010 325894
rect 311062 325842 311074 325894
rect 311126 325842 311138 325894
rect 311190 325842 311196 325894
rect 310876 325830 311196 325842
rect 310876 325778 310882 325830
rect 310934 325778 310946 325830
rect 310998 325778 311010 325830
rect 311062 325778 311074 325830
rect 311126 325778 311138 325830
rect 311190 325778 311196 325830
rect 310876 325772 311196 325778
rect 292482 325252 292488 325304
rect 292540 325252 292546 325304
rect 292500 325224 292528 325252
rect 295168 325224 295196 325263
rect 292500 325196 295196 325224
rect 295150 324572 295156 324624
rect 295208 324612 295214 324624
rect 295208 324584 297956 324612
rect 295208 324572 295214 324584
rect 297928 324462 297956 324584
rect 301774 324028 301780 324080
rect 301832 324068 301838 324080
rect 301908 324071 301966 324077
rect 301908 324068 301920 324071
rect 301832 324040 301920 324068
rect 301832 324028 301838 324040
rect 301908 324037 301920 324040
rect 301954 324037 301966 324071
rect 301908 324031 301966 324037
rect 303876 323914 304196 323920
rect 303876 323862 303882 323914
rect 303934 323862 303946 323914
rect 303998 323862 304010 323914
rect 304062 323862 304074 323914
rect 304126 323862 304138 323914
rect 304190 323862 304196 323914
rect 303876 323850 304196 323862
rect 303876 323798 303882 323850
rect 303934 323798 303946 323850
rect 303998 323798 304010 323850
rect 304062 323798 304074 323850
rect 304126 323798 304138 323850
rect 304190 323798 304196 323850
rect 303876 323786 304196 323798
rect 303876 323734 303882 323786
rect 303934 323734 303946 323786
rect 303998 323734 304010 323786
rect 304062 323734 304074 323786
rect 304126 323734 304138 323786
rect 304190 323734 304196 323786
rect 303876 323722 304196 323734
rect 303876 323670 303882 323722
rect 303934 323670 303946 323722
rect 303998 323670 304010 323722
rect 304062 323670 304074 323722
rect 304126 323670 304138 323722
rect 304190 323670 304196 323722
rect 303876 323658 304196 323670
rect 303876 323606 303882 323658
rect 303934 323606 303946 323658
rect 303998 323606 304010 323658
rect 304062 323606 304074 323658
rect 304126 323606 304138 323658
rect 304190 323606 304196 323658
rect 303876 323600 304196 323606
rect 310876 323914 311196 323920
rect 310876 323862 310882 323914
rect 310934 323862 310946 323914
rect 310998 323862 311010 323914
rect 311062 323862 311074 323914
rect 311126 323862 311138 323914
rect 311190 323862 311196 323914
rect 310876 323850 311196 323862
rect 310876 323798 310882 323850
rect 310934 323798 310946 323850
rect 310998 323798 311010 323850
rect 311062 323798 311074 323850
rect 311126 323798 311138 323850
rect 311190 323798 311196 323850
rect 310876 323786 311196 323798
rect 310876 323734 310882 323786
rect 310934 323734 310946 323786
rect 310998 323734 311010 323786
rect 311062 323734 311074 323786
rect 311126 323734 311138 323786
rect 311190 323734 311196 323786
rect 310876 323722 311196 323734
rect 310876 323670 310882 323722
rect 310934 323670 310946 323722
rect 310998 323670 311010 323722
rect 311062 323670 311074 323722
rect 311126 323670 311138 323722
rect 311190 323670 311196 323722
rect 310876 323658 311196 323670
rect 310876 323606 310882 323658
rect 310934 323606 310946 323658
rect 310998 323606 311010 323658
rect 311062 323606 311074 323658
rect 311126 323606 311138 323658
rect 311190 323606 311196 323658
rect 310876 323600 311196 323606
rect 296876 305116 297196 305122
rect 296876 305064 296882 305116
rect 296934 305064 296946 305116
rect 296998 305064 297010 305116
rect 297062 305064 297074 305116
rect 297126 305064 297138 305116
rect 297190 305064 297196 305116
rect 296876 305052 297196 305064
rect 296876 305000 296882 305052
rect 296934 305000 296946 305052
rect 296998 305000 297010 305052
rect 297062 305000 297074 305052
rect 297126 305000 297138 305052
rect 297190 305000 297196 305052
rect 296876 304988 297196 305000
rect 296876 304936 296882 304988
rect 296934 304936 296946 304988
rect 296998 304936 297010 304988
rect 297062 304936 297074 304988
rect 297126 304936 297138 304988
rect 297190 304936 297196 304988
rect 296876 304924 297196 304936
rect 296876 304872 296882 304924
rect 296934 304872 296946 304924
rect 296998 304872 297010 304924
rect 297062 304872 297074 304924
rect 297126 304872 297138 304924
rect 297190 304872 297196 304924
rect 296876 304860 297196 304872
rect 296876 304808 296882 304860
rect 296934 304808 296946 304860
rect 296998 304808 297010 304860
rect 297062 304808 297074 304860
rect 297126 304808 297138 304860
rect 297190 304808 297196 304860
rect 296876 304802 297196 304808
rect 303876 305116 304196 305122
rect 303876 305064 303882 305116
rect 303934 305064 303946 305116
rect 303998 305064 304010 305116
rect 304062 305064 304074 305116
rect 304126 305064 304138 305116
rect 304190 305064 304196 305116
rect 303876 305052 304196 305064
rect 303876 305000 303882 305052
rect 303934 305000 303946 305052
rect 303998 305000 304010 305052
rect 304062 305000 304074 305052
rect 304126 305000 304138 305052
rect 304190 305000 304196 305052
rect 303876 304988 304196 305000
rect 303876 304936 303882 304988
rect 303934 304936 303946 304988
rect 303998 304936 304010 304988
rect 304062 304936 304074 304988
rect 304126 304936 304138 304988
rect 304190 304936 304196 304988
rect 303876 304924 304196 304936
rect 303876 304872 303882 304924
rect 303934 304872 303946 304924
rect 303998 304872 304010 304924
rect 304062 304872 304074 304924
rect 304126 304872 304138 304924
rect 304190 304872 304196 304924
rect 303876 304860 304196 304872
rect 303876 304808 303882 304860
rect 303934 304808 303946 304860
rect 303998 304808 304010 304860
rect 304062 304808 304074 304860
rect 304126 304808 304138 304860
rect 304190 304808 304196 304860
rect 303876 304802 304196 304808
rect 310876 305116 311196 305122
rect 310876 305064 310882 305116
rect 310934 305064 310946 305116
rect 310998 305064 311010 305116
rect 311062 305064 311074 305116
rect 311126 305064 311138 305116
rect 311190 305064 311196 305116
rect 310876 305052 311196 305064
rect 310876 305000 310882 305052
rect 310934 305000 310946 305052
rect 310998 305000 311010 305052
rect 311062 305000 311074 305052
rect 311126 305000 311138 305052
rect 311190 305000 311196 305052
rect 310876 304988 311196 305000
rect 310876 304936 310882 304988
rect 310934 304936 310946 304988
rect 310998 304936 311010 304988
rect 311062 304936 311074 304988
rect 311126 304936 311138 304988
rect 311190 304936 311196 304988
rect 310876 304924 311196 304936
rect 310876 304872 310882 304924
rect 310934 304872 310946 304924
rect 310998 304872 311010 304924
rect 311062 304872 311074 304924
rect 311126 304872 311138 304924
rect 311190 304872 311196 304924
rect 310876 304860 311196 304872
rect 310876 304808 310882 304860
rect 310934 304808 310946 304860
rect 310998 304808 311010 304860
rect 311062 304808 311074 304860
rect 311126 304808 311138 304860
rect 311190 304808 311196 304860
rect 310876 304802 311196 304808
rect 292482 304308 292488 304360
rect 292540 304308 292546 304360
rect 297456 304319 297508 304325
rect 292500 304280 292528 304308
rect 295260 304280 295288 304293
rect 292500 304252 295288 304280
rect 312354 304267 312360 304319
rect 312412 304267 312418 304319
rect 297456 304261 297508 304267
rect 295150 304172 295156 304224
rect 295208 304212 295214 304224
rect 297450 304212 297456 304224
rect 295208 304184 297456 304212
rect 295208 304172 295214 304184
rect 297450 304172 297456 304184
rect 297508 304212 297514 304224
rect 298094 304212 298100 304224
rect 297508 304184 298100 304212
rect 297508 304172 297514 304184
rect 298094 304172 298100 304184
rect 298152 304172 298158 304224
rect 312354 304104 312360 304156
rect 312412 304144 312418 304156
rect 313826 304144 313832 304156
rect 312412 304116 313832 304144
rect 312412 304104 312418 304116
rect 313826 304104 313832 304116
rect 313884 304104 313890 304156
rect 302144 304015 302464 304036
rect 302144 303963 302150 304015
rect 302202 303963 302214 304015
rect 302266 303963 302278 304015
rect 302330 303963 302342 304015
rect 302394 303963 302406 304015
rect 302458 303963 302464 304015
rect 302144 303951 302464 303963
rect 302144 303899 302150 303951
rect 302202 303899 302214 303951
rect 302266 303899 302278 303951
rect 302330 303899 302342 303951
rect 302394 303899 302406 303951
rect 302458 303899 302464 303951
rect 302144 303887 302464 303899
rect 302144 303835 302150 303887
rect 302202 303835 302214 303887
rect 302266 303835 302278 303887
rect 302330 303835 302342 303887
rect 302394 303835 302406 303887
rect 302458 303835 302464 303887
rect 302144 303823 302464 303835
rect 302144 303771 302150 303823
rect 302202 303771 302214 303823
rect 302266 303771 302278 303823
rect 302330 303771 302342 303823
rect 302394 303771 302406 303823
rect 302458 303771 302464 303823
rect 302144 303759 302464 303771
rect 302144 303707 302150 303759
rect 302202 303707 302214 303759
rect 302266 303707 302278 303759
rect 302330 303707 302342 303759
rect 302394 303707 302406 303759
rect 302458 303707 302464 303759
rect 302144 303686 302464 303707
rect 309144 304015 309464 304036
rect 309144 303963 309150 304015
rect 309202 303963 309214 304015
rect 309266 303963 309278 304015
rect 309330 303963 309342 304015
rect 309394 303963 309406 304015
rect 309458 303963 309464 304015
rect 309144 303951 309464 303963
rect 309144 303899 309150 303951
rect 309202 303899 309214 303951
rect 309266 303899 309278 303951
rect 309330 303899 309342 303951
rect 309394 303899 309406 303951
rect 309458 303899 309464 303951
rect 309144 303887 309464 303899
rect 309144 303835 309150 303887
rect 309202 303835 309214 303887
rect 309266 303835 309278 303887
rect 309330 303835 309342 303887
rect 309394 303835 309406 303887
rect 309458 303835 309464 303887
rect 309144 303823 309464 303835
rect 309144 303771 309150 303823
rect 309202 303771 309214 303823
rect 309266 303771 309278 303823
rect 309330 303771 309342 303823
rect 309394 303771 309406 303823
rect 309458 303771 309464 303823
rect 309144 303759 309464 303771
rect 309144 303707 309150 303759
rect 309202 303707 309214 303759
rect 309266 303707 309278 303759
rect 309330 303707 309342 303759
rect 309394 303707 309406 303759
rect 309458 303707 309464 303759
rect 309144 303686 309464 303707
rect 313642 303532 313648 303544
rect 309152 303504 313648 303532
rect 309152 303450 309180 303504
rect 313642 303492 313648 303504
rect 313700 303492 313706 303544
rect 314286 302880 314292 302932
rect 314344 302920 314350 302932
rect 515766 302920 515772 302932
rect 314344 302892 515772 302920
rect 314344 302880 314350 302892
rect 515766 302880 515772 302892
rect 515824 302880 515830 302932
rect 313642 302132 313648 302184
rect 313700 302172 313706 302184
rect 314470 302172 314476 302184
rect 313700 302144 314476 302172
rect 313700 302132 313706 302144
rect 314470 302132 314476 302144
rect 314528 302132 314534 302184
rect 376018 284316 376024 284368
rect 376076 284356 376082 284368
rect 514754 284356 514760 284368
rect 376076 284328 514760 284356
rect 376076 284316 376082 284328
rect 514754 284316 514760 284328
rect 514812 284316 514818 284368
rect 292482 283228 292488 283280
rect 292540 283268 292546 283280
rect 311466 283268 311572 283279
rect 312630 283268 312636 283280
rect 292540 283240 295288 283268
rect 311466 283251 312636 283268
rect 311544 283240 312636 283251
rect 292540 283228 292546 283240
rect 312630 283228 312636 283240
rect 312688 283268 312694 283280
rect 312814 283268 312820 283280
rect 312688 283240 312820 283268
rect 312688 283228 312694 283240
rect 312814 283228 312820 283240
rect 312872 283228 312878 283280
rect 302144 283000 302464 283006
rect 302144 282948 302150 283000
rect 302202 282948 302214 283000
rect 302266 282948 302278 283000
rect 302330 282948 302342 283000
rect 302394 282948 302406 283000
rect 302458 282948 302464 283000
rect 302144 282936 302464 282948
rect 302144 282884 302150 282936
rect 302202 282884 302214 282936
rect 302266 282884 302278 282936
rect 302330 282884 302342 282936
rect 302394 282884 302406 282936
rect 302458 282884 302464 282936
rect 302144 282872 302464 282884
rect 302144 282820 302150 282872
rect 302202 282820 302214 282872
rect 302266 282820 302278 282872
rect 302330 282820 302342 282872
rect 302394 282820 302406 282872
rect 302458 282820 302464 282872
rect 302144 282808 302464 282820
rect 302144 282756 302150 282808
rect 302202 282756 302214 282808
rect 302266 282756 302278 282808
rect 302330 282756 302342 282808
rect 302394 282756 302406 282808
rect 302458 282756 302464 282808
rect 302144 282744 302464 282756
rect 302144 282692 302150 282744
rect 302202 282692 302214 282744
rect 302266 282692 302278 282744
rect 302330 282692 302342 282744
rect 302394 282692 302406 282744
rect 302458 282692 302464 282744
rect 302144 282686 302464 282692
rect 309144 283001 309464 283008
rect 309144 282949 309150 283001
rect 309202 282949 309214 283001
rect 309266 282949 309278 283001
rect 309330 282949 309342 283001
rect 309394 282949 309406 283001
rect 309458 282949 309464 283001
rect 309144 282937 309464 282949
rect 309144 282885 309150 282937
rect 309202 282885 309214 282937
rect 309266 282885 309278 282937
rect 309330 282885 309342 282937
rect 309394 282885 309406 282937
rect 309458 282885 309464 282937
rect 309144 282873 309464 282885
rect 309144 282821 309150 282873
rect 309202 282821 309214 282873
rect 309266 282821 309278 282873
rect 309330 282821 309342 282873
rect 309394 282821 309406 282873
rect 309458 282821 309464 282873
rect 309144 282809 309464 282821
rect 309144 282757 309150 282809
rect 309202 282757 309214 282809
rect 309266 282757 309278 282809
rect 309330 282757 309342 282809
rect 309394 282757 309406 282809
rect 309458 282757 309464 282809
rect 309144 282745 309464 282757
rect 309144 282693 309150 282745
rect 309202 282693 309214 282745
rect 309266 282693 309278 282745
rect 309330 282693 309342 282745
rect 309394 282693 309406 282745
rect 309458 282693 309464 282745
rect 309144 282686 309464 282693
rect 303876 282239 304196 282250
rect 303876 282187 303882 282239
rect 303934 282187 303946 282239
rect 303998 282187 304010 282239
rect 304062 282187 304074 282239
rect 304126 282187 304138 282239
rect 304190 282187 304196 282239
rect 303876 282175 304196 282187
rect 303876 282123 303882 282175
rect 303934 282123 303946 282175
rect 303998 282123 304010 282175
rect 304062 282123 304074 282175
rect 304126 282123 304138 282175
rect 304190 282123 304196 282175
rect 303876 282111 304196 282123
rect 303876 282059 303882 282111
rect 303934 282059 303946 282111
rect 303998 282059 304010 282111
rect 304062 282059 304074 282111
rect 304126 282059 304138 282111
rect 304190 282059 304196 282111
rect 310876 282192 311196 282220
rect 310876 282140 310882 282192
rect 310934 282140 310946 282192
rect 310998 282140 311010 282192
rect 311062 282140 311074 282192
rect 311126 282140 311138 282192
rect 311190 282140 311196 282192
rect 310876 282128 311196 282140
rect 298974 282047 299032 282053
rect 298974 282013 298986 282047
rect 299020 282044 299032 282047
rect 299106 282044 299112 282056
rect 299020 282016 299112 282044
rect 299020 282013 299032 282016
rect 298974 282007 299032 282013
rect 299106 282004 299112 282016
rect 299164 282004 299170 282056
rect 302291 282047 302349 282053
rect 302291 282013 302303 282047
rect 302337 282044 302349 282047
rect 302418 282044 302424 282056
rect 302337 282016 302424 282044
rect 302337 282013 302349 282016
rect 302291 282007 302349 282013
rect 302418 282004 302424 282016
rect 302476 282004 302482 282056
rect 303876 282047 304196 282059
rect 308956 282087 309008 282093
rect 303876 281995 303882 282047
rect 303934 281995 303946 282047
rect 303998 281995 304010 282047
rect 304062 281995 304074 282047
rect 304126 281995 304138 282047
rect 304190 281995 304196 282047
rect 305608 282047 305666 282053
rect 305608 282013 305620 282047
rect 305654 282044 305666 282047
rect 305730 282044 305736 282056
rect 305654 282016 305736 282044
rect 305654 282013 305666 282016
rect 305608 282007 305666 282013
rect 305730 282004 305736 282016
rect 305788 282004 305794 282056
rect 308956 282029 309008 282035
rect 310876 282076 310882 282128
rect 310934 282076 310946 282128
rect 310998 282076 311010 282128
rect 311062 282076 311074 282128
rect 311126 282076 311138 282128
rect 311190 282076 311196 282128
rect 310876 282064 311196 282076
rect 310876 282012 310882 282064
rect 310934 282012 310946 282064
rect 310998 282012 311010 282064
rect 311062 282012 311074 282064
rect 311126 282012 311138 282064
rect 311190 282012 311196 282064
rect 312294 282056 312584 282075
rect 312294 282047 312544 282056
rect 303876 281983 304196 281995
rect 303876 281931 303882 281983
rect 303934 281931 303946 281983
rect 303998 281931 304010 281983
rect 304062 281931 304074 281983
rect 304126 281931 304138 281983
rect 304190 281931 304196 281983
rect 303876 281919 304196 281931
rect 303876 281867 303882 281919
rect 303934 281867 303946 281919
rect 303998 281867 304010 281919
rect 304062 281867 304074 281919
rect 304126 281867 304138 281919
rect 304190 281867 304196 281919
rect 303876 281855 304196 281867
rect 303876 281803 303882 281855
rect 303934 281803 303946 281855
rect 303998 281803 304010 281855
rect 304062 281803 304074 281855
rect 304126 281803 304138 281855
rect 304190 281803 304196 281855
rect 303876 281791 304196 281803
rect 303876 281739 303882 281791
rect 303934 281739 303946 281791
rect 303998 281739 304010 281791
rect 304062 281739 304074 281791
rect 304126 281739 304138 281791
rect 304190 281739 304196 281791
rect 303876 281727 304196 281739
rect 303876 281675 303882 281727
rect 303934 281675 303946 281727
rect 303998 281675 304010 281727
rect 304062 281675 304074 281727
rect 304126 281675 304138 281727
rect 304190 281675 304196 281727
rect 303876 281663 304196 281675
rect 303876 281611 303882 281663
rect 303934 281611 303946 281663
rect 303998 281611 304010 281663
rect 304062 281611 304074 281663
rect 304126 281611 304138 281663
rect 304190 281611 304196 281663
rect 303876 281600 304196 281611
rect 310876 282000 311196 282012
rect 312538 282004 312544 282047
rect 312596 282004 312602 282056
rect 310876 281948 310882 282000
rect 310934 281948 310946 282000
rect 310998 281948 311010 282000
rect 311062 281948 311074 282000
rect 311126 281948 311138 282000
rect 311190 281948 311196 282000
rect 310876 281936 311196 281948
rect 310876 281884 310882 281936
rect 310934 281884 310946 281936
rect 310998 281884 311010 281936
rect 311062 281884 311074 281936
rect 311126 281884 311138 281936
rect 311190 281884 311196 281936
rect 310876 281872 311196 281884
rect 310876 281820 310882 281872
rect 310934 281820 310946 281872
rect 310998 281820 311010 281872
rect 311062 281820 311074 281872
rect 311126 281820 311138 281872
rect 311190 281820 311196 281872
rect 310876 281808 311196 281820
rect 310876 281756 310882 281808
rect 310934 281756 310946 281808
rect 310998 281756 311010 281808
rect 311062 281756 311074 281808
rect 311126 281756 311138 281808
rect 311190 281756 311196 281808
rect 310876 281744 311196 281756
rect 310876 281692 310882 281744
rect 310934 281692 310946 281744
rect 310998 281692 311010 281744
rect 311062 281692 311074 281744
rect 311126 281692 311138 281744
rect 311190 281692 311196 281744
rect 310876 281680 311196 281692
rect 310876 281628 310882 281680
rect 310934 281628 310946 281680
rect 310998 281628 311010 281680
rect 311062 281628 311074 281680
rect 311126 281628 311138 281680
rect 311190 281628 311196 281680
rect 310876 281600 311196 281628
rect 298186 262692 298192 262744
rect 298244 262692 298250 262744
rect 299290 262692 299296 262744
rect 299348 262692 299354 262744
rect 305086 262692 305092 262744
rect 305144 262692 305150 262744
rect 308766 262692 308772 262744
rect 308824 262692 308830 262744
rect 292482 262420 292488 262472
rect 292540 262460 292546 262472
rect 292540 262432 295196 262460
rect 292540 262420 292546 262432
rect 295168 262263 295196 262432
rect 298204 262278 298232 262692
rect 299308 262469 299336 262692
rect 299305 262463 299363 262469
rect 299305 262429 299317 262463
rect 299351 262429 299363 262463
rect 299305 262423 299363 262429
rect 305104 262392 305132 262692
rect 305100 262364 305132 262392
rect 298204 262250 298239 262278
rect 305100 262250 305128 262364
rect 308784 262277 308812 262692
rect 298211 262249 298239 262250
rect 308614 262249 308812 262277
rect 312722 262256 312728 262268
rect 312018 262228 312728 262256
rect 312722 262216 312728 262228
rect 312780 262256 312786 262268
rect 312998 262256 313004 262268
rect 312780 262228 313004 262256
rect 312780 262216 312786 262228
rect 312998 262216 313004 262228
rect 313056 262216 313062 262268
rect 302144 262000 302464 262006
rect 302144 261948 302150 262000
rect 302202 261948 302214 262000
rect 302266 261948 302278 262000
rect 302330 261948 302342 262000
rect 302394 261948 302406 262000
rect 302458 261948 302464 262000
rect 302144 261936 302464 261948
rect 302144 261884 302150 261936
rect 302202 261884 302214 261936
rect 302266 261884 302278 261936
rect 302330 261884 302342 261936
rect 302394 261884 302406 261936
rect 302458 261884 302464 261936
rect 302144 261872 302464 261884
rect 302144 261820 302150 261872
rect 302202 261820 302214 261872
rect 302266 261820 302278 261872
rect 302330 261820 302342 261872
rect 302394 261820 302406 261872
rect 302458 261820 302464 261872
rect 302144 261808 302464 261820
rect 302144 261756 302150 261808
rect 302202 261756 302214 261808
rect 302266 261756 302278 261808
rect 302330 261756 302342 261808
rect 302394 261756 302406 261808
rect 302458 261756 302464 261808
rect 302144 261744 302464 261756
rect 302144 261692 302150 261744
rect 302202 261692 302214 261744
rect 302266 261692 302278 261744
rect 302330 261692 302342 261744
rect 302394 261692 302406 261744
rect 302458 261692 302464 261744
rect 302144 261686 302464 261692
rect 309144 262000 309464 262006
rect 309144 261948 309150 262000
rect 309202 261948 309214 262000
rect 309266 261948 309278 262000
rect 309330 261948 309342 262000
rect 309394 261948 309406 262000
rect 309458 261948 309464 262000
rect 309144 261936 309464 261948
rect 309144 261884 309150 261936
rect 309202 261884 309214 261936
rect 309266 261884 309278 261936
rect 309330 261884 309342 261936
rect 309394 261884 309406 261936
rect 309458 261884 309464 261936
rect 309144 261872 309464 261884
rect 309144 261820 309150 261872
rect 309202 261820 309214 261872
rect 309266 261820 309278 261872
rect 309330 261820 309342 261872
rect 309394 261820 309406 261872
rect 309458 261820 309464 261872
rect 309144 261808 309464 261820
rect 309144 261756 309150 261808
rect 309202 261756 309214 261808
rect 309266 261756 309278 261808
rect 309330 261756 309342 261808
rect 309394 261756 309406 261808
rect 309458 261756 309464 261808
rect 309144 261744 309464 261756
rect 309144 261692 309150 261744
rect 309202 261692 309214 261744
rect 309266 261692 309278 261744
rect 309330 261692 309342 261744
rect 309394 261692 309406 261744
rect 309458 261692 309464 261744
rect 309144 261686 309464 261692
rect 303876 261239 304196 261250
rect 303876 261187 303882 261239
rect 303934 261187 303946 261239
rect 303998 261187 304010 261239
rect 304062 261187 304074 261239
rect 304126 261187 304138 261239
rect 304190 261187 304196 261239
rect 303876 261175 304196 261187
rect 303876 261123 303882 261175
rect 303934 261123 303946 261175
rect 303998 261123 304010 261175
rect 304062 261123 304074 261175
rect 304126 261123 304138 261175
rect 304190 261123 304196 261175
rect 303876 261111 304196 261123
rect 303876 261059 303882 261111
rect 303934 261059 303946 261111
rect 303998 261059 304010 261111
rect 304062 261059 304074 261111
rect 304126 261059 304138 261111
rect 304190 261059 304196 261111
rect 303876 261047 304196 261059
rect 302472 261035 302530 261041
rect 302472 261001 302484 261035
rect 302518 261032 302530 261035
rect 302602 261032 302608 261044
rect 302518 261004 302608 261032
rect 302518 261001 302530 261004
rect 302472 260995 302530 261001
rect 302602 260992 302608 261004
rect 302660 260992 302666 261044
rect 303876 260995 303882 261047
rect 303934 260995 303946 261047
rect 303998 260995 304010 261047
rect 304062 260995 304074 261047
rect 304126 260995 304138 261047
rect 304190 260995 304196 261047
rect 303876 260983 304196 260995
rect 303876 260931 303882 260983
rect 303934 260931 303946 260983
rect 303998 260931 304010 260983
rect 304062 260931 304074 260983
rect 304126 260931 304138 260983
rect 304190 260931 304196 260983
rect 303876 260919 304196 260931
rect 303876 260867 303882 260919
rect 303934 260867 303946 260919
rect 303998 260867 304010 260919
rect 304062 260867 304074 260919
rect 304126 260867 304138 260919
rect 304190 260867 304196 260919
rect 303876 260855 304196 260867
rect 303876 260803 303882 260855
rect 303934 260803 303946 260855
rect 303998 260803 304010 260855
rect 304062 260803 304074 260855
rect 304126 260803 304138 260855
rect 304190 260803 304196 260855
rect 303876 260791 304196 260803
rect 303876 260739 303882 260791
rect 303934 260739 303946 260791
rect 303998 260739 304010 260791
rect 304062 260739 304074 260791
rect 304126 260739 304138 260791
rect 304190 260739 304196 260791
rect 303876 260727 304196 260739
rect 303876 260675 303882 260727
rect 303934 260675 303946 260727
rect 303998 260675 304010 260727
rect 304062 260675 304074 260727
rect 304126 260675 304138 260727
rect 304190 260675 304196 260727
rect 303876 260663 304196 260675
rect 303876 260611 303882 260663
rect 303934 260611 303946 260663
rect 303998 260611 304010 260663
rect 304062 260611 304074 260663
rect 304126 260611 304138 260663
rect 304190 260611 304196 260663
rect 303876 260600 304196 260611
rect 296876 242086 297196 242092
rect 296876 242034 296882 242086
rect 296934 242034 296946 242086
rect 296998 242034 297010 242086
rect 297062 242034 297074 242086
rect 297126 242034 297138 242086
rect 297190 242034 297196 242086
rect 296876 242022 297196 242034
rect 296876 241970 296882 242022
rect 296934 241970 296946 242022
rect 296998 241970 297010 242022
rect 297062 241970 297074 242022
rect 297126 241970 297138 242022
rect 297190 241970 297196 242022
rect 296876 241958 297196 241970
rect 296876 241906 296882 241958
rect 296934 241906 296946 241958
rect 296998 241906 297010 241958
rect 297062 241906 297074 241958
rect 297126 241906 297138 241958
rect 297190 241906 297196 241958
rect 296876 241894 297196 241906
rect 296876 241842 296882 241894
rect 296934 241842 296946 241894
rect 296998 241842 297010 241894
rect 297062 241842 297074 241894
rect 297126 241842 297138 241894
rect 297190 241842 297196 241894
rect 296876 241830 297196 241842
rect 296876 241778 296882 241830
rect 296934 241778 296946 241830
rect 296998 241778 297010 241830
rect 297062 241778 297074 241830
rect 297126 241778 297138 241830
rect 297190 241778 297196 241830
rect 296876 241772 297196 241778
rect 303876 242086 304196 242092
rect 303876 242034 303882 242086
rect 303934 242034 303946 242086
rect 303998 242034 304010 242086
rect 304062 242034 304074 242086
rect 304126 242034 304138 242086
rect 304190 242034 304196 242086
rect 303876 242022 304196 242034
rect 303876 241970 303882 242022
rect 303934 241970 303946 242022
rect 303998 241970 304010 242022
rect 304062 241970 304074 242022
rect 304126 241970 304138 242022
rect 304190 241970 304196 242022
rect 303876 241958 304196 241970
rect 303876 241906 303882 241958
rect 303934 241906 303946 241958
rect 303998 241906 304010 241958
rect 304062 241906 304074 241958
rect 304126 241906 304138 241958
rect 304190 241906 304196 241958
rect 303876 241894 304196 241906
rect 303876 241842 303882 241894
rect 303934 241842 303946 241894
rect 303998 241842 304010 241894
rect 304062 241842 304074 241894
rect 304126 241842 304138 241894
rect 304190 241842 304196 241894
rect 303876 241830 304196 241842
rect 303876 241778 303882 241830
rect 303934 241778 303946 241830
rect 303998 241778 304010 241830
rect 304062 241778 304074 241830
rect 304126 241778 304138 241830
rect 304190 241778 304196 241830
rect 303876 241772 304196 241778
rect 310876 242086 311196 242092
rect 310876 242034 310882 242086
rect 310934 242034 310946 242086
rect 310998 242034 311010 242086
rect 311062 242034 311074 242086
rect 311126 242034 311138 242086
rect 311190 242034 311196 242086
rect 310876 242022 311196 242034
rect 310876 241970 310882 242022
rect 310934 241970 310946 242022
rect 310998 241970 311010 242022
rect 311062 241970 311074 242022
rect 311126 241970 311138 242022
rect 311190 241970 311196 242022
rect 310876 241958 311196 241970
rect 310876 241906 310882 241958
rect 310934 241906 310946 241958
rect 310998 241906 311010 241958
rect 311062 241906 311074 241958
rect 311126 241906 311138 241958
rect 311190 241906 311196 241958
rect 310876 241894 311196 241906
rect 310876 241842 310882 241894
rect 310934 241842 310946 241894
rect 310998 241842 311010 241894
rect 311062 241842 311074 241894
rect 311126 241842 311138 241894
rect 311190 241842 311196 241894
rect 310876 241830 311196 241842
rect 310876 241778 310882 241830
rect 310934 241778 310946 241830
rect 310998 241778 311010 241830
rect 311062 241778 311074 241830
rect 311126 241778 311138 241830
rect 311190 241778 311196 241830
rect 310876 241772 311196 241778
rect 311066 241612 311072 241664
rect 311124 241652 311130 241664
rect 312446 241652 312452 241664
rect 311124 241624 312452 241652
rect 311124 241612 311130 241624
rect 312446 241612 312452 241624
rect 312504 241652 312510 241664
rect 314378 241652 314384 241664
rect 312504 241624 314384 241652
rect 312504 241612 312510 241624
rect 314378 241612 314384 241624
rect 314436 241612 314442 241664
rect 292482 241408 292488 241460
rect 292540 241448 292546 241460
rect 292540 241420 295196 241448
rect 292540 241408 292546 241420
rect 295168 241263 295196 241420
rect 296898 241237 296904 241289
rect 296956 241237 296962 241289
rect 300946 241237 300952 241289
rect 301004 241237 301010 241289
rect 295242 241136 295248 241188
rect 295300 241176 295306 241188
rect 296898 241176 296904 241188
rect 295300 241148 296904 241176
rect 295300 241136 295306 241148
rect 296898 241136 296904 241148
rect 296956 241136 296962 241188
rect 295144 241001 295464 241007
rect 295144 240949 295150 241001
rect 295202 240949 295214 241001
rect 295266 240949 295278 241001
rect 295330 240949 295342 241001
rect 295394 240949 295406 241001
rect 295458 240949 295464 241001
rect 295144 240937 295464 240949
rect 295144 240885 295150 240937
rect 295202 240885 295214 240937
rect 295266 240885 295278 240937
rect 295330 240885 295342 240937
rect 295394 240885 295406 240937
rect 295458 240885 295464 240937
rect 295144 240873 295464 240885
rect 295144 240821 295150 240873
rect 295202 240821 295214 240873
rect 295266 240821 295278 240873
rect 295330 240821 295342 240873
rect 295394 240821 295406 240873
rect 295458 240821 295464 240873
rect 295144 240809 295464 240821
rect 295144 240757 295150 240809
rect 295202 240757 295214 240809
rect 295266 240757 295278 240809
rect 295330 240757 295342 240809
rect 295394 240757 295406 240809
rect 295458 240757 295464 240809
rect 295144 240745 295464 240757
rect 295144 240693 295150 240745
rect 295202 240693 295214 240745
rect 295266 240693 295278 240745
rect 295330 240693 295342 240745
rect 295394 240693 295406 240745
rect 295458 240693 295464 240745
rect 295144 240687 295464 240693
rect 309144 240975 309464 241007
rect 309144 240923 309150 240975
rect 309202 240923 309214 240975
rect 309266 240923 309278 240975
rect 309330 240923 309342 240975
rect 309394 240923 309406 240975
rect 309458 240923 309464 240975
rect 309144 240911 309464 240923
rect 309144 240859 309150 240911
rect 309202 240859 309214 240911
rect 309266 240859 309278 240911
rect 309330 240859 309342 240911
rect 309394 240859 309406 240911
rect 309458 240859 309464 240911
rect 309144 240847 309464 240859
rect 309144 240795 309150 240847
rect 309202 240795 309214 240847
rect 309266 240795 309278 240847
rect 309330 240795 309342 240847
rect 309394 240795 309406 240847
rect 309458 240795 309464 240847
rect 309144 240783 309464 240795
rect 309144 240731 309150 240783
rect 309202 240731 309214 240783
rect 309266 240731 309278 240783
rect 309330 240731 309342 240783
rect 309394 240731 309406 240783
rect 309458 240731 309464 240783
rect 309144 240719 309464 240731
rect 309144 240667 309150 240719
rect 309202 240667 309214 240719
rect 309266 240667 309278 240719
rect 309330 240667 309342 240719
rect 309394 240667 309406 240719
rect 309458 240667 309464 240719
rect 309144 240635 309464 240667
rect 312538 240564 312544 240576
rect 307864 240536 312544 240564
rect 302142 240505 302148 240508
rect 302113 240499 302148 240505
rect 302113 240465 302125 240499
rect 302113 240459 302148 240465
rect 302142 240456 302148 240459
rect 302200 240456 302206 240508
rect 307864 240429 307892 240536
rect 312538 240524 312544 240536
rect 312596 240524 312602 240576
rect 308674 240505 308680 240508
rect 308643 240499 308680 240505
rect 308643 240465 308655 240499
rect 308643 240459 308680 240465
rect 308674 240456 308680 240459
rect 308732 240456 308738 240508
rect 298836 240085 298888 240091
rect 298836 240027 298888 240033
rect 305368 240085 305420 240091
rect 514754 240088 514760 240100
rect 311912 240060 514760 240088
rect 311912 240059 311940 240060
rect 514754 240048 514760 240060
rect 514812 240048 514818 240100
rect 305368 240027 305420 240033
rect 310876 239914 311196 239920
rect 310876 239862 310882 239914
rect 310934 239862 310946 239914
rect 310998 239862 311010 239914
rect 311062 239862 311074 239914
rect 311126 239862 311138 239914
rect 311190 239862 311196 239914
rect 310876 239850 311196 239862
rect 310876 239798 310882 239850
rect 310934 239798 310946 239850
rect 310998 239798 311010 239850
rect 311062 239798 311074 239850
rect 311126 239798 311138 239850
rect 311190 239798 311196 239850
rect 310876 239786 311196 239798
rect 310876 239734 310882 239786
rect 310934 239734 310946 239786
rect 310998 239734 311010 239786
rect 311062 239734 311074 239786
rect 311126 239734 311138 239786
rect 311190 239734 311196 239786
rect 310876 239722 311196 239734
rect 310876 239670 310882 239722
rect 310934 239670 310946 239722
rect 310998 239670 311010 239722
rect 311062 239670 311074 239722
rect 311126 239670 311138 239722
rect 311190 239670 311196 239722
rect 310876 239658 311196 239670
rect 310876 239606 310882 239658
rect 310934 239606 310946 239658
rect 310998 239606 311010 239658
rect 311062 239606 311074 239658
rect 311126 239606 311138 239658
rect 311190 239606 311196 239658
rect 310876 239600 311196 239606
rect 308674 238688 308680 238740
rect 308732 238728 308738 238740
rect 376018 238728 376024 238740
rect 308732 238700 376024 238728
rect 308732 238688 308738 238700
rect 376018 238688 376024 238700
rect 376076 238688 376082 238740
rect 298830 238620 298836 238672
rect 298888 238660 298894 238672
rect 316862 238660 316868 238672
rect 298888 238632 316868 238660
rect 298888 238620 298894 238632
rect 316862 238620 316868 238632
rect 316920 238620 316926 238672
rect 302142 238552 302148 238604
rect 302200 238592 302206 238604
rect 313918 238592 313924 238604
rect 302200 238564 313924 238592
rect 302200 238552 302206 238564
rect 313918 238552 313924 238564
rect 313976 238552 313982 238604
rect 305362 238484 305368 238536
rect 305420 238524 305426 238536
rect 314286 238524 314292 238536
rect 305420 238496 314292 238524
rect 305420 238484 305426 238496
rect 314286 238484 314292 238496
rect 314344 238484 314350 238536
rect 296876 221087 297196 221093
rect 296876 221035 296882 221087
rect 296934 221035 296946 221087
rect 296998 221035 297010 221087
rect 297062 221035 297074 221087
rect 297126 221035 297138 221087
rect 297190 221035 297196 221087
rect 296876 221023 297196 221035
rect 296876 220971 296882 221023
rect 296934 220971 296946 221023
rect 296998 220971 297010 221023
rect 297062 220971 297074 221023
rect 297126 220971 297138 221023
rect 297190 220971 297196 221023
rect 296876 220959 297196 220971
rect 296876 220907 296882 220959
rect 296934 220907 296946 220959
rect 296998 220907 297010 220959
rect 297062 220907 297074 220959
rect 297126 220907 297138 220959
rect 297190 220907 297196 220959
rect 296876 220895 297196 220907
rect 296876 220843 296882 220895
rect 296934 220843 296946 220895
rect 296998 220843 297010 220895
rect 297062 220843 297074 220895
rect 297126 220843 297138 220895
rect 297190 220843 297196 220895
rect 296876 220831 297196 220843
rect 296876 220779 296882 220831
rect 296934 220779 296946 220831
rect 296998 220779 297010 220831
rect 297062 220779 297074 220831
rect 297126 220779 297138 220831
rect 297190 220779 297196 220831
rect 296876 220773 297196 220779
rect 303876 221087 304196 221093
rect 303876 221035 303882 221087
rect 303934 221035 303946 221087
rect 303998 221035 304010 221087
rect 304062 221035 304074 221087
rect 304126 221035 304138 221087
rect 304190 221035 304196 221087
rect 303876 221023 304196 221035
rect 303876 220971 303882 221023
rect 303934 220971 303946 221023
rect 303998 220971 304010 221023
rect 304062 220971 304074 221023
rect 304126 220971 304138 221023
rect 304190 220971 304196 221023
rect 303876 220959 304196 220971
rect 303876 220907 303882 220959
rect 303934 220907 303946 220959
rect 303998 220907 304010 220959
rect 304062 220907 304074 220959
rect 304126 220907 304138 220959
rect 304190 220907 304196 220959
rect 303876 220895 304196 220907
rect 303876 220843 303882 220895
rect 303934 220843 303946 220895
rect 303998 220843 304010 220895
rect 304062 220843 304074 220895
rect 304126 220843 304138 220895
rect 304190 220843 304196 220895
rect 303876 220831 304196 220843
rect 303876 220779 303882 220831
rect 303934 220779 303946 220831
rect 303998 220779 304010 220831
rect 304062 220779 304074 220831
rect 304126 220779 304138 220831
rect 304190 220779 304196 220831
rect 303876 220773 304196 220779
rect 310876 221087 311196 221093
rect 310876 221035 310882 221087
rect 310934 221035 310946 221087
rect 310998 221035 311010 221087
rect 311062 221035 311074 221087
rect 311126 221035 311138 221087
rect 311190 221035 311196 221087
rect 310876 221023 311196 221035
rect 310876 220971 310882 221023
rect 310934 220971 310946 221023
rect 310998 220971 311010 221023
rect 311062 220971 311074 221023
rect 311126 220971 311138 221023
rect 311190 220971 311196 221023
rect 310876 220959 311196 220971
rect 310876 220907 310882 220959
rect 310934 220907 310946 220959
rect 310998 220907 311010 220959
rect 311062 220907 311074 220959
rect 311126 220907 311138 220959
rect 311190 220907 311196 220959
rect 310876 220895 311196 220907
rect 310876 220843 310882 220895
rect 310934 220843 310946 220895
rect 310998 220843 311010 220895
rect 311062 220843 311074 220895
rect 311126 220843 311138 220895
rect 311190 220843 311196 220895
rect 310876 220831 311196 220843
rect 310876 220779 310882 220831
rect 310934 220779 310946 220831
rect 310998 220779 311010 220831
rect 311062 220779 311074 220831
rect 311126 220779 311138 220831
rect 311190 220779 311196 220831
rect 310876 220773 311196 220779
rect 292482 220464 292488 220516
rect 292540 220464 292546 220516
rect 294966 220464 294972 220516
rect 295024 220504 295030 220516
rect 297341 220507 297399 220513
rect 297341 220504 297353 220507
rect 295024 220476 297353 220504
rect 295024 220464 295030 220476
rect 297341 220473 297353 220476
rect 297387 220473 297399 220507
rect 297341 220467 297399 220473
rect 292500 220436 292528 220464
rect 292500 220408 295196 220436
rect 295168 220265 295196 220408
rect 313918 220300 313924 220312
rect 313476 220278 313924 220300
rect 313398 220272 313924 220278
rect 313398 220250 313504 220272
rect 313918 220260 313924 220272
rect 313976 220300 313982 220312
rect 314378 220300 314384 220312
rect 313976 220272 314384 220300
rect 313976 220260 313982 220272
rect 314378 220260 314384 220272
rect 314436 220260 314442 220312
rect 295144 220002 295464 220008
rect 295144 219950 295150 220002
rect 295202 219950 295214 220002
rect 295266 219950 295278 220002
rect 295330 219950 295342 220002
rect 295394 219950 295406 220002
rect 295458 219950 295464 220002
rect 295144 219938 295464 219950
rect 295144 219886 295150 219938
rect 295202 219886 295214 219938
rect 295266 219886 295278 219938
rect 295330 219886 295342 219938
rect 295394 219886 295406 219938
rect 295458 219886 295464 219938
rect 295144 219874 295464 219886
rect 295144 219822 295150 219874
rect 295202 219822 295214 219874
rect 295266 219822 295278 219874
rect 295330 219822 295342 219874
rect 295394 219822 295406 219874
rect 295458 219822 295464 219874
rect 295144 219810 295464 219822
rect 295144 219758 295150 219810
rect 295202 219758 295214 219810
rect 295266 219758 295278 219810
rect 295330 219758 295342 219810
rect 295394 219758 295406 219810
rect 295458 219758 295464 219810
rect 295144 219746 295464 219758
rect 295144 219694 295150 219746
rect 295202 219694 295214 219746
rect 295266 219694 295278 219746
rect 295330 219694 295342 219746
rect 295394 219694 295406 219746
rect 295458 219694 295464 219746
rect 295144 219688 295464 219694
rect 302144 220001 302464 220008
rect 302144 219949 302150 220001
rect 302202 219949 302214 220001
rect 302266 219949 302278 220001
rect 302330 219949 302342 220001
rect 302394 219949 302406 220001
rect 302458 219949 302464 220001
rect 302144 219937 302464 219949
rect 302144 219885 302150 219937
rect 302202 219885 302214 219937
rect 302266 219885 302278 219937
rect 302330 219885 302342 219937
rect 302394 219885 302406 219937
rect 302458 219885 302464 219937
rect 302144 219873 302464 219885
rect 302144 219821 302150 219873
rect 302202 219821 302214 219873
rect 302266 219821 302278 219873
rect 302330 219821 302342 219873
rect 302394 219821 302406 219873
rect 302458 219821 302464 219873
rect 302144 219809 302464 219821
rect 302144 219757 302150 219809
rect 302202 219757 302214 219809
rect 302266 219757 302278 219809
rect 302330 219757 302342 219809
rect 302394 219757 302406 219809
rect 302458 219757 302464 219809
rect 302144 219745 302464 219757
rect 302144 219693 302150 219745
rect 302202 219693 302214 219745
rect 302266 219693 302278 219745
rect 302330 219693 302342 219745
rect 302394 219693 302406 219745
rect 302458 219693 302464 219745
rect 302144 219686 302464 219693
rect 309144 220001 309464 220008
rect 309144 219949 309150 220001
rect 309202 219949 309214 220001
rect 309266 219949 309278 220001
rect 309330 219949 309342 220001
rect 309394 219949 309406 220001
rect 309458 219949 309464 220001
rect 309144 219937 309464 219949
rect 309144 219885 309150 219937
rect 309202 219885 309214 219937
rect 309266 219885 309278 219937
rect 309330 219885 309342 219937
rect 309394 219885 309406 219937
rect 309458 219885 309464 219937
rect 309144 219873 309464 219885
rect 309144 219821 309150 219873
rect 309202 219821 309214 219873
rect 309266 219821 309278 219873
rect 309330 219821 309342 219873
rect 309394 219821 309406 219873
rect 309458 219821 309464 219873
rect 309144 219809 309464 219821
rect 309144 219757 309150 219809
rect 309202 219757 309214 219809
rect 309266 219757 309278 219809
rect 309330 219757 309342 219809
rect 309394 219757 309406 219809
rect 309458 219757 309464 219809
rect 309144 219745 309464 219757
rect 309144 219693 309150 219745
rect 309202 219693 309214 219745
rect 309266 219693 309278 219745
rect 309330 219693 309342 219745
rect 309394 219693 309406 219745
rect 309458 219693 309464 219745
rect 309144 219686 309464 219693
rect 311039 219461 311045 219513
rect 311097 219461 311103 219513
rect 303962 219396 304020 219407
rect 303962 219344 303965 219396
rect 304017 219344 304020 219396
rect 303962 219333 304020 219344
rect 299296 219085 299348 219091
rect 303007 219079 303065 219085
rect 303007 219045 303019 219079
rect 303053 219076 303065 219079
rect 303154 219076 303160 219088
rect 303053 219048 303160 219076
rect 303053 219045 303065 219048
rect 303007 219039 303065 219045
rect 303154 219036 303160 219048
rect 303212 219036 303218 219088
rect 306748 219085 306800 219091
rect 299296 219027 299348 219033
rect 306748 219027 306800 219033
rect 310428 219085 310480 219091
rect 310428 219027 310480 219033
rect 292482 206252 292488 206304
rect 292540 206292 292546 206304
rect 580166 206292 580172 206304
rect 292540 206264 580172 206292
rect 292540 206252 292546 206264
rect 580166 206252 580172 206264
rect 580224 206252 580230 206304
rect 295242 199316 295248 199368
rect 295300 199356 295306 199368
rect 296681 199359 296739 199365
rect 296681 199356 296693 199359
rect 295300 199328 296693 199356
rect 295300 199316 295306 199328
rect 296681 199325 296693 199328
rect 296727 199325 296739 199359
rect 296681 199319 296739 199325
rect 292482 199248 292488 199300
rect 292540 199288 292546 199300
rect 292540 199260 295196 199288
rect 292540 199248 292546 199260
rect 311066 198472 311072 198484
rect 310072 198444 311072 198472
rect 307050 198415 307156 198443
rect 310072 198429 310100 198444
rect 311066 198432 311072 198444
rect 311124 198472 311130 198484
rect 311250 198472 311256 198484
rect 311124 198444 311256 198472
rect 311124 198432 311130 198444
rect 311250 198432 311256 198444
rect 311308 198432 311314 198484
rect 307128 198404 307156 198415
rect 307662 198404 307668 198416
rect 307128 198376 307668 198404
rect 307662 198364 307668 198376
rect 307720 198364 307726 198416
rect 296876 179287 297196 179293
rect 296876 179235 296882 179287
rect 296934 179235 296946 179287
rect 296998 179235 297010 179287
rect 297062 179235 297074 179287
rect 297126 179235 297138 179287
rect 297190 179235 297196 179287
rect 296876 179223 297196 179235
rect 296876 179171 296882 179223
rect 296934 179171 296946 179223
rect 296998 179171 297010 179223
rect 297062 179171 297074 179223
rect 297126 179171 297138 179223
rect 297190 179171 297196 179223
rect 296876 179159 297196 179171
rect 296876 179107 296882 179159
rect 296934 179107 296946 179159
rect 296998 179107 297010 179159
rect 297062 179107 297074 179159
rect 297126 179107 297138 179159
rect 297190 179107 297196 179159
rect 296876 179095 297196 179107
rect 296876 179043 296882 179095
rect 296934 179043 296946 179095
rect 296998 179043 297010 179095
rect 297062 179043 297074 179095
rect 297126 179043 297138 179095
rect 297190 179043 297196 179095
rect 296876 179031 297196 179043
rect 296876 178979 296882 179031
rect 296934 178979 296946 179031
rect 296998 178979 297010 179031
rect 297062 178979 297074 179031
rect 297126 178979 297138 179031
rect 297190 178979 297196 179031
rect 296876 178973 297196 178979
rect 303876 179287 304196 179293
rect 303876 179235 303882 179287
rect 303934 179235 303946 179287
rect 303998 179235 304010 179287
rect 304062 179235 304074 179287
rect 304126 179235 304138 179287
rect 304190 179235 304196 179287
rect 303876 179223 304196 179235
rect 303876 179171 303882 179223
rect 303934 179171 303946 179223
rect 303998 179171 304010 179223
rect 304062 179171 304074 179223
rect 304126 179171 304138 179223
rect 304190 179171 304196 179223
rect 303876 179159 304196 179171
rect 303876 179107 303882 179159
rect 303934 179107 303946 179159
rect 303998 179107 304010 179159
rect 304062 179107 304074 179159
rect 304126 179107 304138 179159
rect 304190 179107 304196 179159
rect 303876 179095 304196 179107
rect 303876 179043 303882 179095
rect 303934 179043 303946 179095
rect 303998 179043 304010 179095
rect 304062 179043 304074 179095
rect 304126 179043 304138 179095
rect 304190 179043 304196 179095
rect 303876 179031 304196 179043
rect 303876 178979 303882 179031
rect 303934 178979 303946 179031
rect 303998 178979 304010 179031
rect 304062 178979 304074 179031
rect 304126 178979 304138 179031
rect 304190 178979 304196 179031
rect 303876 178973 304196 178979
rect 310876 179287 310964 179293
rect 310876 179235 310894 179287
rect 310946 179235 310964 179287
rect 310876 179223 310964 179235
rect 310876 179171 310894 179223
rect 310946 179171 310964 179223
rect 310876 179159 310964 179171
rect 310876 179107 310894 179159
rect 310946 179107 310964 179159
rect 310876 179095 310964 179107
rect 310876 179043 310894 179095
rect 310946 179043 310964 179095
rect 310876 179031 310964 179043
rect 310876 178979 310894 179031
rect 310946 178979 310964 179031
rect 310876 178973 310964 178979
rect 292482 178712 292488 178764
rect 292540 178752 292546 178764
rect 292540 178724 295196 178752
rect 292540 178712 292546 178724
rect 295168 178464 295196 178724
rect 297266 178438 297272 178490
rect 297324 178438 297330 178490
rect 295144 178201 295464 178207
rect 295144 178149 295150 178201
rect 295202 178149 295214 178201
rect 295266 178149 295278 178201
rect 295330 178149 295342 178201
rect 295394 178149 295406 178201
rect 295458 178149 295464 178201
rect 295144 178137 295464 178149
rect 295144 178085 295150 178137
rect 295202 178085 295214 178137
rect 295266 178085 295278 178137
rect 295330 178085 295342 178137
rect 295394 178085 295406 178137
rect 295458 178085 295464 178137
rect 295144 178073 295464 178085
rect 295144 178021 295150 178073
rect 295202 178021 295214 178073
rect 295266 178021 295278 178073
rect 295330 178021 295342 178073
rect 295394 178021 295406 178073
rect 295458 178021 295464 178073
rect 295144 178009 295464 178021
rect 295144 177957 295150 178009
rect 295202 177957 295214 178009
rect 295266 177957 295278 178009
rect 295330 177957 295342 178009
rect 295394 177957 295406 178009
rect 295458 177957 295464 178009
rect 295144 177945 295464 177957
rect 295144 177893 295150 177945
rect 295202 177893 295214 177945
rect 295266 177893 295278 177945
rect 295330 177893 295342 177945
rect 295394 177893 295406 177945
rect 295458 177893 295464 177945
rect 295144 177887 295464 177893
rect 302144 178185 302464 178207
rect 302144 178133 302150 178185
rect 302202 178133 302214 178185
rect 302266 178133 302278 178185
rect 302330 178133 302342 178185
rect 302394 178133 302406 178185
rect 302458 178133 302464 178185
rect 302144 178121 302464 178133
rect 302144 178069 302150 178121
rect 302202 178069 302214 178121
rect 302266 178069 302278 178121
rect 302330 178069 302342 178121
rect 302394 178069 302406 178121
rect 302458 178069 302464 178121
rect 302144 178057 302464 178069
rect 302144 178005 302150 178057
rect 302202 178005 302214 178057
rect 302266 178005 302278 178057
rect 302330 178005 302342 178057
rect 302394 178005 302406 178057
rect 302458 178005 302464 178057
rect 302144 177993 302464 178005
rect 302144 177941 302150 177993
rect 302202 177941 302214 177993
rect 302266 177941 302278 177993
rect 302330 177941 302342 177993
rect 302394 177941 302406 177993
rect 302458 177941 302464 177993
rect 302144 177929 302464 177941
rect 302144 177877 302150 177929
rect 302202 177877 302214 177929
rect 302266 177877 302278 177929
rect 302330 177877 302342 177929
rect 302394 177877 302406 177929
rect 302458 177877 302464 177929
rect 302144 177855 302464 177877
rect 309144 178185 309464 178207
rect 309144 178133 309150 178185
rect 309202 178133 309214 178185
rect 309266 178133 309278 178185
rect 309330 178133 309342 178185
rect 309394 178133 309406 178185
rect 309458 178133 309464 178185
rect 309144 178121 309464 178133
rect 309144 178069 309150 178121
rect 309202 178069 309214 178121
rect 309266 178069 309278 178121
rect 309330 178069 309342 178121
rect 309394 178069 309406 178121
rect 309458 178069 309464 178121
rect 309144 178057 309464 178069
rect 309144 178005 309150 178057
rect 309202 178005 309214 178057
rect 309266 178005 309278 178057
rect 309330 178005 309342 178057
rect 309394 178005 309406 178057
rect 309458 178005 309464 178057
rect 309144 177993 309464 178005
rect 309144 177941 309150 177993
rect 309202 177941 309214 177993
rect 309266 177941 309278 177993
rect 309330 177941 309342 177993
rect 309394 177941 309406 177993
rect 309458 177941 309464 177993
rect 309144 177929 309464 177941
rect 309144 177877 309150 177929
rect 309202 177877 309214 177929
rect 309266 177877 309278 177929
rect 309330 177877 309342 177929
rect 309394 177877 309406 177929
rect 309458 177877 309464 177929
rect 309144 177855 309464 177877
rect 311250 177664 311256 177676
rect 310072 177636 311256 177664
rect 310072 177629 310100 177636
rect 311250 177624 311256 177636
rect 311308 177664 311314 177676
rect 311526 177664 311532 177676
rect 311308 177636 311532 177664
rect 311308 177624 311314 177636
rect 311526 177624 311532 177636
rect 311584 177624 311590 177676
<< via1 >>
rect 296882 491604 296934 491656
rect 296946 491604 296998 491656
rect 297010 491604 297062 491656
rect 297074 491604 297126 491656
rect 297138 491604 297190 491656
rect 296882 491540 296934 491592
rect 296946 491540 296998 491592
rect 297010 491540 297062 491592
rect 297074 491540 297126 491592
rect 297138 491540 297190 491592
rect 296882 491476 296934 491528
rect 296946 491476 296998 491528
rect 297010 491476 297062 491528
rect 297074 491476 297126 491528
rect 297138 491476 297190 491528
rect 296882 491412 296934 491464
rect 296946 491412 296998 491464
rect 297010 491412 297062 491464
rect 297074 491412 297126 491464
rect 297138 491412 297190 491464
rect 296882 491348 296934 491400
rect 296946 491348 296998 491400
rect 297010 491348 297062 491400
rect 297074 491348 297126 491400
rect 297138 491348 297190 491400
rect 303882 491604 303934 491656
rect 303946 491604 303998 491656
rect 304010 491604 304062 491656
rect 304074 491604 304126 491656
rect 304138 491604 304190 491656
rect 303882 491540 303934 491592
rect 303946 491540 303998 491592
rect 304010 491540 304062 491592
rect 304074 491540 304126 491592
rect 304138 491540 304190 491592
rect 303882 491476 303934 491528
rect 303946 491476 303998 491528
rect 304010 491476 304062 491528
rect 304074 491476 304126 491528
rect 304138 491476 304190 491528
rect 303882 491412 303934 491464
rect 303946 491412 303998 491464
rect 304010 491412 304062 491464
rect 304074 491412 304126 491464
rect 304138 491412 304190 491464
rect 303882 491348 303934 491400
rect 303946 491348 303998 491400
rect 304010 491348 304062 491400
rect 304074 491348 304126 491400
rect 304138 491348 304190 491400
rect 310882 491604 310934 491656
rect 310946 491604 310998 491656
rect 311010 491604 311062 491656
rect 311074 491604 311126 491656
rect 311138 491604 311190 491656
rect 310882 491540 310934 491592
rect 310946 491540 310998 491592
rect 311010 491540 311062 491592
rect 311074 491540 311126 491592
rect 311138 491540 311190 491592
rect 310882 491476 310934 491528
rect 310946 491476 310998 491528
rect 311010 491476 311062 491528
rect 311074 491476 311126 491528
rect 311138 491476 311190 491528
rect 310882 491412 310934 491464
rect 310946 491412 310998 491464
rect 311010 491412 311062 491464
rect 311074 491412 311126 491464
rect 311138 491412 311190 491464
rect 310882 491348 310934 491400
rect 310946 491348 310998 491400
rect 311010 491348 311062 491400
rect 311074 491348 311126 491400
rect 311138 491348 311190 491400
rect 292488 490696 292540 490748
rect 296996 490807 297048 490859
rect 294880 490628 294932 490680
rect 296996 490628 297048 490680
rect 295150 490496 295202 490548
rect 295214 490496 295266 490548
rect 295278 490496 295330 490548
rect 295342 490496 295394 490548
rect 295406 490496 295458 490548
rect 295150 490432 295202 490484
rect 295214 490432 295266 490484
rect 295278 490432 295330 490484
rect 295342 490432 295394 490484
rect 295406 490432 295458 490484
rect 295150 490368 295202 490420
rect 295214 490368 295266 490420
rect 295278 490368 295330 490420
rect 295342 490368 295394 490420
rect 295406 490368 295458 490420
rect 295150 490304 295202 490356
rect 295214 490304 295266 490356
rect 295278 490304 295330 490356
rect 295342 490304 295394 490356
rect 295406 490304 295458 490356
rect 305092 490059 305144 490068
rect 305092 490025 305100 490059
rect 305100 490025 305144 490059
rect 305092 490016 305144 490025
rect 312084 490152 312136 490204
rect 298744 489744 298796 489796
rect 308128 489676 308180 489728
rect 301780 489603 301832 489655
rect 311532 489603 311584 489655
rect 303882 489432 303934 489484
rect 303946 489432 303998 489484
rect 304010 489432 304062 489484
rect 304074 489432 304126 489484
rect 304138 489432 304190 489484
rect 303882 489368 303934 489420
rect 303946 489368 303998 489420
rect 304010 489368 304062 489420
rect 304074 489368 304126 489420
rect 304138 489368 304190 489420
rect 303882 489304 303934 489356
rect 303946 489304 303998 489356
rect 304010 489304 304062 489356
rect 304074 489304 304126 489356
rect 304138 489304 304190 489356
rect 303882 489240 303934 489292
rect 303946 489240 303998 489292
rect 304010 489240 304062 489292
rect 304074 489240 304126 489292
rect 304138 489240 304190 489292
rect 303882 489176 303934 489228
rect 303946 489176 303998 489228
rect 304010 489176 304062 489228
rect 304074 489176 304126 489228
rect 304138 489176 304190 489228
rect 310882 489432 310934 489484
rect 310946 489432 310998 489484
rect 311010 489432 311062 489484
rect 311074 489432 311126 489484
rect 311138 489432 311190 489484
rect 310882 489368 310934 489420
rect 310946 489368 310998 489420
rect 311010 489368 311062 489420
rect 311074 489368 311126 489420
rect 311138 489368 311190 489420
rect 310882 489304 310934 489356
rect 310946 489304 310998 489356
rect 311010 489304 311062 489356
rect 311074 489304 311126 489356
rect 311138 489304 311190 489356
rect 310882 489240 310934 489292
rect 310946 489240 310998 489292
rect 311010 489240 311062 489292
rect 311074 489240 311126 489292
rect 311138 489240 311190 489292
rect 310882 489176 310934 489228
rect 310946 489176 310998 489228
rect 311010 489176 311062 489228
rect 311074 489176 311126 489228
rect 311138 489176 311190 489228
rect 296882 473064 296934 473116
rect 296946 473064 296998 473116
rect 297010 473064 297062 473116
rect 297074 473064 297126 473116
rect 297138 473064 297190 473116
rect 296882 473000 296934 473052
rect 296946 473000 296998 473052
rect 297010 473000 297062 473052
rect 297074 473000 297126 473052
rect 297138 473000 297190 473052
rect 296882 472936 296934 472988
rect 296946 472936 296998 472988
rect 297010 472936 297062 472988
rect 297074 472936 297126 472988
rect 297138 472936 297190 472988
rect 296882 472872 296934 472924
rect 296946 472872 296998 472924
rect 297010 472872 297062 472924
rect 297074 472872 297126 472924
rect 297138 472872 297190 472924
rect 296882 472808 296934 472860
rect 296946 472808 296998 472860
rect 297010 472808 297062 472860
rect 297074 472808 297126 472860
rect 297138 472808 297190 472860
rect 303882 473064 303934 473116
rect 303946 473064 303998 473116
rect 304010 473064 304062 473116
rect 304074 473064 304126 473116
rect 304138 473064 304190 473116
rect 303882 473000 303934 473052
rect 303946 473000 303998 473052
rect 304010 473000 304062 473052
rect 304074 473000 304126 473052
rect 304138 473000 304190 473052
rect 303882 472936 303934 472988
rect 303946 472936 303998 472988
rect 304010 472936 304062 472988
rect 304074 472936 304126 472988
rect 304138 472936 304190 472988
rect 303882 472872 303934 472924
rect 303946 472872 303998 472924
rect 304010 472872 304062 472924
rect 304074 472872 304126 472924
rect 304138 472872 304190 472924
rect 303882 472808 303934 472860
rect 303946 472808 303998 472860
rect 304010 472808 304062 472860
rect 304074 472808 304126 472860
rect 304138 472808 304190 472860
rect 310882 473064 310934 473116
rect 310946 473064 310998 473116
rect 311010 473064 311062 473116
rect 311074 473064 311126 473116
rect 311138 473064 311190 473116
rect 310882 473000 310934 473052
rect 310946 473000 310998 473052
rect 311010 473000 311062 473052
rect 311074 473000 311126 473052
rect 311138 473000 311190 473052
rect 310882 472936 310934 472988
rect 310946 472936 310998 472988
rect 311010 472936 311062 472988
rect 311074 472936 311126 472988
rect 311138 472936 311190 472988
rect 310882 472872 310934 472924
rect 310946 472872 310998 472924
rect 311010 472872 311062 472924
rect 311074 472872 311126 472924
rect 311138 472872 311190 472924
rect 310882 472808 310934 472860
rect 310946 472808 310998 472860
rect 311010 472808 311062 472860
rect 311074 472808 311126 472860
rect 311138 472808 311190 472860
rect 294880 472540 294932 472592
rect 295248 472540 295300 472592
rect 292488 472336 292540 472388
rect 309140 472267 309192 472319
rect 302150 471963 302202 472015
rect 302214 471963 302266 472015
rect 302278 471963 302330 472015
rect 302342 471963 302394 472015
rect 302406 471963 302458 472015
rect 302150 471899 302202 471951
rect 302214 471899 302266 471951
rect 302278 471899 302330 471951
rect 302342 471899 302394 471951
rect 302406 471899 302458 471951
rect 302150 471835 302202 471887
rect 302214 471835 302266 471887
rect 302278 471835 302330 471887
rect 302342 471835 302394 471887
rect 302406 471835 302458 471887
rect 302150 471771 302202 471823
rect 302214 471771 302266 471823
rect 302278 471771 302330 471823
rect 302342 471771 302394 471823
rect 302406 471771 302458 471823
rect 302150 471707 302202 471759
rect 302214 471707 302266 471759
rect 302278 471707 302330 471759
rect 302342 471707 302394 471759
rect 302406 471707 302458 471759
rect 309150 471963 309202 472015
rect 309214 471963 309266 472015
rect 309278 471963 309330 472015
rect 309342 471963 309394 472015
rect 309406 471963 309458 472015
rect 309150 471899 309202 471951
rect 309214 471899 309266 471951
rect 309278 471899 309330 471951
rect 309342 471899 309394 471951
rect 309406 471899 309458 471951
rect 309150 471835 309202 471887
rect 309214 471835 309266 471887
rect 309278 471835 309330 471887
rect 309342 471835 309394 471887
rect 309406 471835 309458 471887
rect 309150 471771 309202 471823
rect 309214 471771 309266 471823
rect 309278 471771 309330 471823
rect 309342 471771 309394 471823
rect 309406 471771 309458 471823
rect 309150 471707 309202 471759
rect 309214 471707 309266 471759
rect 309278 471707 309330 471759
rect 309342 471707 309394 471759
rect 309406 471707 309458 471759
rect 313740 471248 313792 471300
rect 299296 471044 299348 471096
rect 302884 471044 302936 471096
rect 306472 471044 306524 471096
rect 313648 471044 313700 471096
rect 313740 471044 313792 471096
rect 296882 452024 296934 452076
rect 296946 452024 296998 452076
rect 297010 452024 297062 452076
rect 297074 452024 297126 452076
rect 297138 452024 297190 452076
rect 296882 451960 296934 452012
rect 296946 451960 296998 452012
rect 297010 451960 297062 452012
rect 297074 451960 297126 452012
rect 297138 451960 297190 452012
rect 296882 451896 296934 451948
rect 296946 451896 296998 451948
rect 297010 451896 297062 451948
rect 297074 451896 297126 451948
rect 297138 451896 297190 451948
rect 296882 451832 296934 451884
rect 296946 451832 296998 451884
rect 297010 451832 297062 451884
rect 297074 451832 297126 451884
rect 297138 451832 297190 451884
rect 296882 451768 296934 451820
rect 296946 451768 296998 451820
rect 297010 451768 297062 451820
rect 297074 451768 297126 451820
rect 297138 451768 297190 451820
rect 296882 451704 296934 451756
rect 296946 451704 296998 451756
rect 297010 451704 297062 451756
rect 297074 451704 297126 451756
rect 297138 451704 297190 451756
rect 296882 451640 296934 451692
rect 296946 451640 296998 451692
rect 297010 451640 297062 451692
rect 297074 451640 297126 451692
rect 297138 451640 297190 451692
rect 296882 451576 296934 451628
rect 296946 451576 296998 451628
rect 297010 451576 297062 451628
rect 297074 451576 297126 451628
rect 297138 451576 297190 451628
rect 296882 451512 296934 451564
rect 296946 451512 296998 451564
rect 297010 451512 297062 451564
rect 297074 451512 297126 451564
rect 297138 451512 297190 451564
rect 296882 451448 296934 451500
rect 296946 451448 296998 451500
rect 297010 451448 297062 451500
rect 297074 451448 297126 451500
rect 297138 451448 297190 451500
rect 296882 451384 296934 451436
rect 296946 451384 296998 451436
rect 297010 451384 297062 451436
rect 297074 451384 297126 451436
rect 297138 451384 297190 451436
rect 292488 451324 292540 451376
rect 296882 451320 296934 451372
rect 296946 451320 296998 451372
rect 297010 451320 297062 451372
rect 297074 451320 297126 451372
rect 297138 451320 297190 451372
rect 296882 451256 296934 451308
rect 296946 451256 296998 451308
rect 297010 451256 297062 451308
rect 297074 451256 297126 451308
rect 297138 451256 297190 451308
rect 295248 451120 295300 451172
rect 303882 452024 303934 452076
rect 303946 452024 303998 452076
rect 304010 452024 304062 452076
rect 304074 452024 304126 452076
rect 304138 452024 304190 452076
rect 303882 451960 303934 452012
rect 303946 451960 303998 452012
rect 304010 451960 304062 452012
rect 304074 451960 304126 452012
rect 304138 451960 304190 452012
rect 303882 451896 303934 451948
rect 303946 451896 303998 451948
rect 304010 451896 304062 451948
rect 304074 451896 304126 451948
rect 304138 451896 304190 451948
rect 303882 451832 303934 451884
rect 303946 451832 303998 451884
rect 304010 451832 304062 451884
rect 304074 451832 304126 451884
rect 304138 451832 304190 451884
rect 303882 451768 303934 451820
rect 303946 451768 303998 451820
rect 304010 451768 304062 451820
rect 304074 451768 304126 451820
rect 304138 451768 304190 451820
rect 303882 451704 303934 451756
rect 303946 451704 303998 451756
rect 304010 451704 304062 451756
rect 304074 451704 304126 451756
rect 304138 451704 304190 451756
rect 303882 451640 303934 451692
rect 303946 451640 303998 451692
rect 304010 451640 304062 451692
rect 304074 451640 304126 451692
rect 304138 451640 304190 451692
rect 303882 451576 303934 451628
rect 303946 451576 303998 451628
rect 304010 451576 304062 451628
rect 304074 451576 304126 451628
rect 304138 451576 304190 451628
rect 303882 451512 303934 451564
rect 303946 451512 303998 451564
rect 304010 451512 304062 451564
rect 304074 451512 304126 451564
rect 304138 451512 304190 451564
rect 303882 451448 303934 451500
rect 303946 451448 303998 451500
rect 304010 451448 304062 451500
rect 304074 451448 304126 451500
rect 304138 451448 304190 451500
rect 303882 451384 303934 451436
rect 303946 451384 303998 451436
rect 304010 451384 304062 451436
rect 304074 451384 304126 451436
rect 304138 451384 304190 451436
rect 303882 451320 303934 451372
rect 303946 451320 303998 451372
rect 304010 451320 304062 451372
rect 304074 451320 304126 451372
rect 304138 451320 304190 451372
rect 303882 451256 303934 451308
rect 303946 451256 303998 451308
rect 304010 451256 304062 451308
rect 304074 451256 304126 451308
rect 304138 451256 304190 451308
rect 310897 452024 310949 452076
rect 310961 452024 311013 452076
rect 311025 452024 311077 452076
rect 310897 451960 310949 452012
rect 310961 451960 311013 452012
rect 311025 451960 311077 452012
rect 310897 451896 310949 451948
rect 310961 451896 311013 451948
rect 311025 451896 311077 451948
rect 310897 451832 310949 451884
rect 310961 451832 311013 451884
rect 311025 451832 311077 451884
rect 310897 451768 310949 451820
rect 310961 451768 311013 451820
rect 311025 451768 311077 451820
rect 310897 451704 310949 451756
rect 310961 451704 311013 451756
rect 311025 451704 311077 451756
rect 310897 451640 310949 451692
rect 310961 451640 311013 451692
rect 311025 451640 311077 451692
rect 310897 451576 310949 451628
rect 310961 451576 311013 451628
rect 311025 451576 311077 451628
rect 310897 451512 310949 451564
rect 310961 451512 311013 451564
rect 311025 451512 311077 451564
rect 310897 451448 310949 451500
rect 310961 451448 311013 451500
rect 311025 451448 311077 451500
rect 310897 451384 310949 451436
rect 310961 451384 311013 451436
rect 311025 451384 311077 451436
rect 310897 451320 310949 451372
rect 310961 451320 311013 451372
rect 311025 451320 311077 451372
rect 310897 451256 310949 451308
rect 310961 451256 311013 451308
rect 311025 451256 311077 451308
rect 313004 450508 313056 450560
rect 300860 450372 300912 450424
rect 306196 450440 306248 450492
rect 310884 450139 310936 450191
rect 310948 450139 311000 450191
rect 311012 450139 311064 450191
rect 311076 450139 311128 450191
rect 310884 450075 310936 450127
rect 310948 450075 311000 450127
rect 311012 450075 311064 450127
rect 311076 450075 311128 450127
rect 310884 450011 310936 450063
rect 310948 450011 311000 450063
rect 311012 450011 311064 450063
rect 311076 450011 311128 450063
rect 310884 449947 310936 449999
rect 310948 449947 311000 449999
rect 311012 449947 311064 449999
rect 311076 449947 311128 449999
rect 310884 449883 310936 449935
rect 310948 449883 311000 449935
rect 311012 449883 311064 449935
rect 311076 449883 311128 449935
rect 310884 449819 310936 449871
rect 310948 449819 311000 449871
rect 311012 449819 311064 449871
rect 311076 449819 311128 449871
rect 310884 449755 310936 449807
rect 310948 449755 311000 449807
rect 311012 449755 311064 449807
rect 311076 449755 311128 449807
rect 310884 449691 310936 449743
rect 310948 449691 311000 449743
rect 311012 449691 311064 449743
rect 311076 449691 311128 449743
rect 310884 449627 310936 449679
rect 310948 449627 311000 449679
rect 311012 449627 311064 449679
rect 311076 449627 311128 449679
rect 292488 430244 292540 430296
rect 295892 430237 295944 430289
rect 312452 430244 312504 430296
rect 312820 430244 312872 430296
rect 309177 429948 309229 430000
rect 309241 429948 309293 430000
rect 309305 429948 309357 430000
rect 309369 429948 309421 430000
rect 309177 429884 309229 429936
rect 309241 429884 309293 429936
rect 309305 429884 309357 429936
rect 309369 429884 309421 429936
rect 309177 429820 309229 429872
rect 309241 429820 309293 429872
rect 309305 429820 309357 429872
rect 309369 429820 309421 429872
rect 309177 429756 309229 429808
rect 309241 429756 309293 429808
rect 309305 429756 309357 429808
rect 309369 429756 309421 429808
rect 309177 429692 309229 429744
rect 309241 429692 309293 429744
rect 309305 429692 309357 429744
rect 309369 429692 309421 429744
rect 301688 429403 301740 429455
rect 301688 429156 301740 429208
rect 299020 429032 299072 429084
rect 305920 429020 305972 429072
rect 313004 429032 313056 429084
rect 302516 428995 302568 429004
rect 302516 428961 302522 428995
rect 302522 428961 302568 428995
rect 302516 428952 302568 428961
rect 526996 421336 527048 421388
rect 529204 421336 529256 421388
rect 296882 410034 296934 410086
rect 296946 410034 296998 410086
rect 297010 410034 297062 410086
rect 297074 410034 297126 410086
rect 297138 410034 297190 410086
rect 296882 409970 296934 410022
rect 296946 409970 296998 410022
rect 297010 409970 297062 410022
rect 297074 409970 297126 410022
rect 297138 409970 297190 410022
rect 296882 409906 296934 409958
rect 296946 409906 296998 409958
rect 297010 409906 297062 409958
rect 297074 409906 297126 409958
rect 297138 409906 297190 409958
rect 296882 409842 296934 409894
rect 296946 409842 296998 409894
rect 297010 409842 297062 409894
rect 297074 409842 297126 409894
rect 297138 409842 297190 409894
rect 296882 409778 296934 409830
rect 296946 409778 296998 409830
rect 297010 409778 297062 409830
rect 297074 409778 297126 409830
rect 297138 409778 297190 409830
rect 303882 410034 303934 410086
rect 303946 410034 303998 410086
rect 304010 410034 304062 410086
rect 304074 410034 304126 410086
rect 304138 410034 304190 410086
rect 303882 409970 303934 410022
rect 303946 409970 303998 410022
rect 304010 409970 304062 410022
rect 304074 409970 304126 410022
rect 304138 409970 304190 410022
rect 303882 409906 303934 409958
rect 303946 409906 303998 409958
rect 304010 409906 304062 409958
rect 304074 409906 304126 409958
rect 304138 409906 304190 409958
rect 303882 409842 303934 409894
rect 303946 409842 303998 409894
rect 304010 409842 304062 409894
rect 304074 409842 304126 409894
rect 304138 409842 304190 409894
rect 303882 409778 303934 409830
rect 303946 409778 303998 409830
rect 304010 409778 304062 409830
rect 304074 409778 304126 409830
rect 304138 409778 304190 409830
rect 310882 410034 310934 410086
rect 310946 410034 310998 410086
rect 311010 410034 311062 410086
rect 311074 410034 311126 410086
rect 311138 410034 311190 410086
rect 310882 409970 310934 410022
rect 310946 409970 310998 410022
rect 311010 409970 311062 410022
rect 311074 409970 311126 410022
rect 311138 409970 311190 410022
rect 310882 409906 310934 409958
rect 310946 409906 310998 409958
rect 311010 409906 311062 409958
rect 311074 409906 311126 409958
rect 311138 409906 311190 409958
rect 310882 409842 310934 409894
rect 310946 409842 310998 409894
rect 311010 409842 311062 409894
rect 311074 409842 311126 409894
rect 311138 409842 311190 409894
rect 310882 409778 310934 409830
rect 310946 409778 310998 409830
rect 311010 409778 311062 409830
rect 311074 409778 311126 409830
rect 311138 409778 311190 409830
rect 295248 409504 295300 409556
rect 292488 409232 292540 409284
rect 302150 408948 302202 409000
rect 302214 408948 302266 409000
rect 302278 408948 302330 409000
rect 302342 408948 302394 409000
rect 302406 408948 302458 409000
rect 302150 408884 302202 408936
rect 302214 408884 302266 408936
rect 302278 408884 302330 408936
rect 302342 408884 302394 408936
rect 302406 408884 302458 408936
rect 302150 408820 302202 408872
rect 302214 408820 302266 408872
rect 302278 408820 302330 408872
rect 302342 408820 302394 408872
rect 302406 408820 302458 408872
rect 302150 408756 302202 408808
rect 302214 408756 302266 408808
rect 302278 408756 302330 408808
rect 302342 408756 302394 408808
rect 302406 408756 302458 408808
rect 302150 408692 302202 408744
rect 302214 408692 302266 408744
rect 302278 408692 302330 408744
rect 302342 408692 302394 408744
rect 302406 408692 302458 408744
rect 313280 408416 313332 408468
rect 314568 408416 314620 408468
rect 312176 408008 312228 408060
rect 310882 407862 310934 407914
rect 310946 407862 310998 407914
rect 311010 407862 311062 407914
rect 311074 407862 311126 407914
rect 311138 407862 311190 407914
rect 310882 407798 310934 407850
rect 310946 407798 310998 407850
rect 311010 407798 311062 407850
rect 311074 407798 311126 407850
rect 311138 407798 311190 407850
rect 310882 407734 310934 407786
rect 310946 407734 310998 407786
rect 311010 407734 311062 407786
rect 311074 407734 311126 407786
rect 311138 407734 311190 407786
rect 310882 407670 310934 407722
rect 310946 407670 310998 407722
rect 311010 407670 311062 407722
rect 311074 407670 311126 407722
rect 311138 407670 311190 407722
rect 310882 407606 310934 407658
rect 310946 407606 310998 407658
rect 311010 407606 311062 407658
rect 311074 407606 311126 407658
rect 311138 407606 311190 407658
rect 316868 404336 316920 404388
rect 514760 404336 514812 404388
rect 296882 389035 296934 389087
rect 296946 389035 296998 389087
rect 297010 389035 297062 389087
rect 297074 389035 297126 389087
rect 297138 389035 297190 389087
rect 296882 388971 296934 389023
rect 296946 388971 296998 389023
rect 297010 388971 297062 389023
rect 297074 388971 297126 389023
rect 297138 388971 297190 389023
rect 296882 388907 296934 388959
rect 296946 388907 296998 388959
rect 297010 388907 297062 388959
rect 297074 388907 297126 388959
rect 297138 388907 297190 388959
rect 296882 388843 296934 388895
rect 296946 388843 296998 388895
rect 297010 388843 297062 388895
rect 297074 388843 297126 388895
rect 297138 388843 297190 388895
rect 296882 388779 296934 388831
rect 296946 388779 296998 388831
rect 297010 388779 297062 388831
rect 297074 388779 297126 388831
rect 297138 388779 297190 388831
rect 303882 389035 303934 389087
rect 303946 389035 303998 389087
rect 304010 389035 304062 389087
rect 304074 389035 304126 389087
rect 304138 389035 304190 389087
rect 303882 388971 303934 389023
rect 303946 388971 303998 389023
rect 304010 388971 304062 389023
rect 304074 388971 304126 389023
rect 304138 388971 304190 389023
rect 303882 388907 303934 388959
rect 303946 388907 303998 388959
rect 304010 388907 304062 388959
rect 304074 388907 304126 388959
rect 304138 388907 304190 388959
rect 303882 388843 303934 388895
rect 303946 388843 303998 388895
rect 304010 388843 304062 388895
rect 304074 388843 304126 388895
rect 304138 388843 304190 388895
rect 303882 388779 303934 388831
rect 303946 388779 303998 388831
rect 304010 388779 304062 388831
rect 304074 388779 304126 388831
rect 304138 388779 304190 388831
rect 310882 389035 310934 389087
rect 310946 389035 310998 389087
rect 311010 389035 311062 389087
rect 311074 389035 311126 389087
rect 311138 389035 311190 389087
rect 310882 388971 310934 389023
rect 310946 388971 310998 389023
rect 311010 388971 311062 389023
rect 311074 388971 311126 389023
rect 311138 388971 311190 389023
rect 310882 388907 310934 388959
rect 310946 388907 310998 388959
rect 311010 388907 311062 388959
rect 311074 388907 311126 388959
rect 311138 388907 311190 388959
rect 310882 388843 310934 388895
rect 310946 388843 310998 388895
rect 311010 388843 311062 388895
rect 311074 388843 311126 388895
rect 311138 388843 311190 388895
rect 310882 388779 310934 388831
rect 310946 388779 310998 388831
rect 311010 388779 311062 388831
rect 311074 388779 311126 388831
rect 311138 388779 311190 388831
rect 295064 388492 295116 388544
rect 292488 388424 292540 388476
rect 301596 388238 301648 388290
rect 295150 387952 295202 388004
rect 295214 387952 295266 388004
rect 295278 387952 295330 388004
rect 295342 387952 295394 388004
rect 295406 387952 295458 388004
rect 295150 387888 295202 387940
rect 295214 387888 295266 387940
rect 295278 387888 295330 387940
rect 295342 387888 295394 387940
rect 295406 387888 295458 387940
rect 295150 387824 295202 387876
rect 295214 387824 295266 387876
rect 295278 387824 295330 387876
rect 295342 387824 295394 387876
rect 295406 387824 295458 387876
rect 295150 387760 295202 387812
rect 295214 387760 295266 387812
rect 295278 387760 295330 387812
rect 295342 387760 295394 387812
rect 295406 387760 295458 387812
rect 295150 387696 295202 387748
rect 295214 387696 295266 387748
rect 295278 387696 295330 387748
rect 295342 387696 295394 387748
rect 295406 387696 295458 387748
rect 302150 387947 302202 387999
rect 302214 387947 302266 387999
rect 302278 387947 302330 387999
rect 302342 387947 302394 387999
rect 302406 387947 302458 387999
rect 302150 387883 302202 387935
rect 302214 387883 302266 387935
rect 302278 387883 302330 387935
rect 302342 387883 302394 387935
rect 302406 387883 302458 387935
rect 302150 387819 302202 387871
rect 302214 387819 302266 387871
rect 302278 387819 302330 387871
rect 302342 387819 302394 387871
rect 302406 387819 302458 387871
rect 302150 387755 302202 387807
rect 302214 387755 302266 387807
rect 302278 387755 302330 387807
rect 302342 387755 302394 387807
rect 302406 387755 302458 387807
rect 302150 387691 302202 387743
rect 302214 387691 302266 387743
rect 302278 387691 302330 387743
rect 302342 387691 302394 387743
rect 302406 387691 302458 387743
rect 309150 387947 309202 387999
rect 309214 387947 309266 387999
rect 309278 387947 309330 387999
rect 309342 387947 309394 387999
rect 309406 387947 309458 387999
rect 309150 387883 309202 387935
rect 309214 387883 309266 387935
rect 309278 387883 309330 387935
rect 309342 387883 309394 387935
rect 309406 387883 309458 387935
rect 309150 387819 309202 387871
rect 309214 387819 309266 387871
rect 309278 387819 309330 387871
rect 309342 387819 309394 387871
rect 309406 387819 309458 387871
rect 309150 387755 309202 387807
rect 309214 387755 309266 387807
rect 309278 387755 309330 387807
rect 309342 387755 309394 387807
rect 309406 387755 309458 387807
rect 309150 387691 309202 387743
rect 309214 387691 309266 387743
rect 309278 387691 309330 387743
rect 309342 387691 309394 387743
rect 309406 387691 309458 387743
rect 311046 387461 311098 387513
rect 303966 387344 304018 387396
rect 299296 387033 299348 387085
rect 303160 386996 303212 387048
rect 306748 387033 306800 387085
rect 310428 387033 310480 387085
rect 295064 374688 295116 374740
rect 295064 374484 295116 374536
rect 294972 370744 295024 370796
rect 295248 370744 295300 370796
rect 292488 367412 292540 367464
rect 296720 367238 296772 367290
rect 299756 367238 299808 367290
rect 295064 367140 295116 367192
rect 296720 367140 296772 367192
rect 307668 366392 307720 366444
rect 307944 366324 307996 366376
rect 298652 366032 298704 366084
rect 301688 366032 301740 366084
rect 304724 366032 304776 366084
rect 313924 364352 313976 364404
rect 514760 364352 514812 364404
rect 310520 347148 310572 347200
rect 311440 347148 311492 347200
rect 296882 347035 296934 347087
rect 296946 347035 296998 347087
rect 297010 347035 297062 347087
rect 297074 347035 297126 347087
rect 297138 347035 297190 347087
rect 296882 346971 296934 347023
rect 296946 346971 296998 347023
rect 297010 346971 297062 347023
rect 297074 346971 297126 347023
rect 297138 346971 297190 347023
rect 296882 346907 296934 346959
rect 296946 346907 296998 346959
rect 297010 346907 297062 346959
rect 297074 346907 297126 346959
rect 297138 346907 297190 346959
rect 296882 346843 296934 346895
rect 296946 346843 296998 346895
rect 297010 346843 297062 346895
rect 297074 346843 297126 346895
rect 297138 346843 297190 346895
rect 296882 346779 296934 346831
rect 296946 346779 296998 346831
rect 297010 346779 297062 346831
rect 297074 346779 297126 346831
rect 297138 346779 297190 346831
rect 303882 347035 303934 347087
rect 303946 347035 303998 347087
rect 304010 347035 304062 347087
rect 304074 347035 304126 347087
rect 304138 347035 304190 347087
rect 303882 346971 303934 347023
rect 303946 346971 303998 347023
rect 304010 346971 304062 347023
rect 304074 346971 304126 347023
rect 304138 346971 304190 347023
rect 303882 346907 303934 346959
rect 303946 346907 303998 346959
rect 304010 346907 304062 346959
rect 304074 346907 304126 346959
rect 304138 346907 304190 346959
rect 303882 346843 303934 346895
rect 303946 346843 303998 346895
rect 304010 346843 304062 346895
rect 304074 346843 304126 346895
rect 304138 346843 304190 346895
rect 303882 346779 303934 346831
rect 303946 346779 303998 346831
rect 304010 346779 304062 346831
rect 304074 346779 304126 346831
rect 304138 346779 304190 346831
rect 295156 346468 295208 346520
rect 292488 346332 292540 346384
rect 302150 345933 302202 345985
rect 302214 345933 302266 345985
rect 302278 345933 302330 345985
rect 302342 345933 302394 345985
rect 302406 345933 302458 345985
rect 302150 345869 302202 345921
rect 302214 345869 302266 345921
rect 302278 345869 302330 345921
rect 302342 345869 302394 345921
rect 302406 345869 302458 345921
rect 302150 345805 302202 345857
rect 302214 345805 302266 345857
rect 302278 345805 302330 345857
rect 302342 345805 302394 345857
rect 302406 345805 302458 345857
rect 302150 345741 302202 345793
rect 302214 345741 302266 345793
rect 302278 345741 302330 345793
rect 302342 345741 302394 345793
rect 302406 345741 302458 345793
rect 302150 345677 302202 345729
rect 302214 345677 302266 345729
rect 302278 345677 302330 345729
rect 302342 345677 302394 345729
rect 302406 345677 302458 345729
rect 309150 345933 309202 345985
rect 309214 345933 309266 345985
rect 309278 345933 309330 345985
rect 309342 345933 309394 345985
rect 309406 345933 309458 345985
rect 309150 345869 309202 345921
rect 309214 345869 309266 345921
rect 309278 345869 309330 345921
rect 309342 345869 309394 345921
rect 309406 345869 309458 345921
rect 309150 345805 309202 345857
rect 309214 345805 309266 345857
rect 309278 345805 309330 345857
rect 309342 345805 309394 345857
rect 309406 345805 309458 345857
rect 309150 345741 309202 345793
rect 309214 345741 309266 345793
rect 309278 345741 309330 345793
rect 309342 345741 309394 345793
rect 309406 345741 309458 345793
rect 309150 345677 309202 345729
rect 309214 345677 309266 345729
rect 309278 345677 309330 345729
rect 309342 345677 309394 345729
rect 309406 345677 309458 345729
rect 298652 345032 298704 345084
rect 301688 345032 301740 345084
rect 304724 345032 304776 345084
rect 307944 345040 307996 345092
rect 296882 326034 296934 326086
rect 296946 326034 296998 326086
rect 297010 326034 297062 326086
rect 297074 326034 297126 326086
rect 297138 326034 297190 326086
rect 296882 325970 296934 326022
rect 296946 325970 296998 326022
rect 297010 325970 297062 326022
rect 297074 325970 297126 326022
rect 297138 325970 297190 326022
rect 296882 325906 296934 325958
rect 296946 325906 296998 325958
rect 297010 325906 297062 325958
rect 297074 325906 297126 325958
rect 297138 325906 297190 325958
rect 296882 325842 296934 325894
rect 296946 325842 296998 325894
rect 297010 325842 297062 325894
rect 297074 325842 297126 325894
rect 297138 325842 297190 325894
rect 296882 325778 296934 325830
rect 296946 325778 296998 325830
rect 297010 325778 297062 325830
rect 297074 325778 297126 325830
rect 297138 325778 297190 325830
rect 303882 326034 303934 326086
rect 303946 326034 303998 326086
rect 304010 326034 304062 326086
rect 304074 326034 304126 326086
rect 304138 326034 304190 326086
rect 303882 325970 303934 326022
rect 303946 325970 303998 326022
rect 304010 325970 304062 326022
rect 304074 325970 304126 326022
rect 304138 325970 304190 326022
rect 303882 325906 303934 325958
rect 303946 325906 303998 325958
rect 304010 325906 304062 325958
rect 304074 325906 304126 325958
rect 304138 325906 304190 325958
rect 303882 325842 303934 325894
rect 303946 325842 303998 325894
rect 304010 325842 304062 325894
rect 304074 325842 304126 325894
rect 304138 325842 304190 325894
rect 303882 325778 303934 325830
rect 303946 325778 303998 325830
rect 304010 325778 304062 325830
rect 304074 325778 304126 325830
rect 304138 325778 304190 325830
rect 310882 326034 310934 326086
rect 310946 326034 310998 326086
rect 311010 326034 311062 326086
rect 311074 326034 311126 326086
rect 311138 326034 311190 326086
rect 310882 325970 310934 326022
rect 310946 325970 310998 326022
rect 311010 325970 311062 326022
rect 311074 325970 311126 326022
rect 311138 325970 311190 326022
rect 310882 325906 310934 325958
rect 310946 325906 310998 325958
rect 311010 325906 311062 325958
rect 311074 325906 311126 325958
rect 311138 325906 311190 325958
rect 310882 325842 310934 325894
rect 310946 325842 310998 325894
rect 311010 325842 311062 325894
rect 311074 325842 311126 325894
rect 311138 325842 311190 325894
rect 310882 325778 310934 325830
rect 310946 325778 310998 325830
rect 311010 325778 311062 325830
rect 311074 325778 311126 325830
rect 311138 325778 311190 325830
rect 292488 325252 292540 325304
rect 295156 324572 295208 324624
rect 301780 324028 301832 324080
rect 303882 323862 303934 323914
rect 303946 323862 303998 323914
rect 304010 323862 304062 323914
rect 304074 323862 304126 323914
rect 304138 323862 304190 323914
rect 303882 323798 303934 323850
rect 303946 323798 303998 323850
rect 304010 323798 304062 323850
rect 304074 323798 304126 323850
rect 304138 323798 304190 323850
rect 303882 323734 303934 323786
rect 303946 323734 303998 323786
rect 304010 323734 304062 323786
rect 304074 323734 304126 323786
rect 304138 323734 304190 323786
rect 303882 323670 303934 323722
rect 303946 323670 303998 323722
rect 304010 323670 304062 323722
rect 304074 323670 304126 323722
rect 304138 323670 304190 323722
rect 303882 323606 303934 323658
rect 303946 323606 303998 323658
rect 304010 323606 304062 323658
rect 304074 323606 304126 323658
rect 304138 323606 304190 323658
rect 310882 323862 310934 323914
rect 310946 323862 310998 323914
rect 311010 323862 311062 323914
rect 311074 323862 311126 323914
rect 311138 323862 311190 323914
rect 310882 323798 310934 323850
rect 310946 323798 310998 323850
rect 311010 323798 311062 323850
rect 311074 323798 311126 323850
rect 311138 323798 311190 323850
rect 310882 323734 310934 323786
rect 310946 323734 310998 323786
rect 311010 323734 311062 323786
rect 311074 323734 311126 323786
rect 311138 323734 311190 323786
rect 310882 323670 310934 323722
rect 310946 323670 310998 323722
rect 311010 323670 311062 323722
rect 311074 323670 311126 323722
rect 311138 323670 311190 323722
rect 310882 323606 310934 323658
rect 310946 323606 310998 323658
rect 311010 323606 311062 323658
rect 311074 323606 311126 323658
rect 311138 323606 311190 323658
rect 296882 305064 296934 305116
rect 296946 305064 296998 305116
rect 297010 305064 297062 305116
rect 297074 305064 297126 305116
rect 297138 305064 297190 305116
rect 296882 305000 296934 305052
rect 296946 305000 296998 305052
rect 297010 305000 297062 305052
rect 297074 305000 297126 305052
rect 297138 305000 297190 305052
rect 296882 304936 296934 304988
rect 296946 304936 296998 304988
rect 297010 304936 297062 304988
rect 297074 304936 297126 304988
rect 297138 304936 297190 304988
rect 296882 304872 296934 304924
rect 296946 304872 296998 304924
rect 297010 304872 297062 304924
rect 297074 304872 297126 304924
rect 297138 304872 297190 304924
rect 296882 304808 296934 304860
rect 296946 304808 296998 304860
rect 297010 304808 297062 304860
rect 297074 304808 297126 304860
rect 297138 304808 297190 304860
rect 303882 305064 303934 305116
rect 303946 305064 303998 305116
rect 304010 305064 304062 305116
rect 304074 305064 304126 305116
rect 304138 305064 304190 305116
rect 303882 305000 303934 305052
rect 303946 305000 303998 305052
rect 304010 305000 304062 305052
rect 304074 305000 304126 305052
rect 304138 305000 304190 305052
rect 303882 304936 303934 304988
rect 303946 304936 303998 304988
rect 304010 304936 304062 304988
rect 304074 304936 304126 304988
rect 304138 304936 304190 304988
rect 303882 304872 303934 304924
rect 303946 304872 303998 304924
rect 304010 304872 304062 304924
rect 304074 304872 304126 304924
rect 304138 304872 304190 304924
rect 303882 304808 303934 304860
rect 303946 304808 303998 304860
rect 304010 304808 304062 304860
rect 304074 304808 304126 304860
rect 304138 304808 304190 304860
rect 310882 305064 310934 305116
rect 310946 305064 310998 305116
rect 311010 305064 311062 305116
rect 311074 305064 311126 305116
rect 311138 305064 311190 305116
rect 310882 305000 310934 305052
rect 310946 305000 310998 305052
rect 311010 305000 311062 305052
rect 311074 305000 311126 305052
rect 311138 305000 311190 305052
rect 310882 304936 310934 304988
rect 310946 304936 310998 304988
rect 311010 304936 311062 304988
rect 311074 304936 311126 304988
rect 311138 304936 311190 304988
rect 310882 304872 310934 304924
rect 310946 304872 310998 304924
rect 311010 304872 311062 304924
rect 311074 304872 311126 304924
rect 311138 304872 311190 304924
rect 310882 304808 310934 304860
rect 310946 304808 310998 304860
rect 311010 304808 311062 304860
rect 311074 304808 311126 304860
rect 311138 304808 311190 304860
rect 292488 304308 292540 304360
rect 297456 304267 297508 304319
rect 312360 304267 312412 304319
rect 295156 304172 295208 304224
rect 297456 304172 297508 304224
rect 298100 304172 298152 304224
rect 312360 304104 312412 304156
rect 313832 304104 313884 304156
rect 302150 303963 302202 304015
rect 302214 303963 302266 304015
rect 302278 303963 302330 304015
rect 302342 303963 302394 304015
rect 302406 303963 302458 304015
rect 302150 303899 302202 303951
rect 302214 303899 302266 303951
rect 302278 303899 302330 303951
rect 302342 303899 302394 303951
rect 302406 303899 302458 303951
rect 302150 303835 302202 303887
rect 302214 303835 302266 303887
rect 302278 303835 302330 303887
rect 302342 303835 302394 303887
rect 302406 303835 302458 303887
rect 302150 303771 302202 303823
rect 302214 303771 302266 303823
rect 302278 303771 302330 303823
rect 302342 303771 302394 303823
rect 302406 303771 302458 303823
rect 302150 303707 302202 303759
rect 302214 303707 302266 303759
rect 302278 303707 302330 303759
rect 302342 303707 302394 303759
rect 302406 303707 302458 303759
rect 309150 303963 309202 304015
rect 309214 303963 309266 304015
rect 309278 303963 309330 304015
rect 309342 303963 309394 304015
rect 309406 303963 309458 304015
rect 309150 303899 309202 303951
rect 309214 303899 309266 303951
rect 309278 303899 309330 303951
rect 309342 303899 309394 303951
rect 309406 303899 309458 303951
rect 309150 303835 309202 303887
rect 309214 303835 309266 303887
rect 309278 303835 309330 303887
rect 309342 303835 309394 303887
rect 309406 303835 309458 303887
rect 309150 303771 309202 303823
rect 309214 303771 309266 303823
rect 309278 303771 309330 303823
rect 309342 303771 309394 303823
rect 309406 303771 309458 303823
rect 309150 303707 309202 303759
rect 309214 303707 309266 303759
rect 309278 303707 309330 303759
rect 309342 303707 309394 303759
rect 309406 303707 309458 303759
rect 313648 303492 313700 303544
rect 314292 302880 314344 302932
rect 515772 302880 515824 302932
rect 313648 302132 313700 302184
rect 314476 302132 314528 302184
rect 376024 284316 376076 284368
rect 514760 284316 514812 284368
rect 292488 283228 292540 283280
rect 312636 283228 312688 283280
rect 312820 283228 312872 283280
rect 302150 282948 302202 283000
rect 302214 282948 302266 283000
rect 302278 282948 302330 283000
rect 302342 282948 302394 283000
rect 302406 282948 302458 283000
rect 302150 282884 302202 282936
rect 302214 282884 302266 282936
rect 302278 282884 302330 282936
rect 302342 282884 302394 282936
rect 302406 282884 302458 282936
rect 302150 282820 302202 282872
rect 302214 282820 302266 282872
rect 302278 282820 302330 282872
rect 302342 282820 302394 282872
rect 302406 282820 302458 282872
rect 302150 282756 302202 282808
rect 302214 282756 302266 282808
rect 302278 282756 302330 282808
rect 302342 282756 302394 282808
rect 302406 282756 302458 282808
rect 302150 282692 302202 282744
rect 302214 282692 302266 282744
rect 302278 282692 302330 282744
rect 302342 282692 302394 282744
rect 302406 282692 302458 282744
rect 309150 282949 309202 283001
rect 309214 282949 309266 283001
rect 309278 282949 309330 283001
rect 309342 282949 309394 283001
rect 309406 282949 309458 283001
rect 309150 282885 309202 282937
rect 309214 282885 309266 282937
rect 309278 282885 309330 282937
rect 309342 282885 309394 282937
rect 309406 282885 309458 282937
rect 309150 282821 309202 282873
rect 309214 282821 309266 282873
rect 309278 282821 309330 282873
rect 309342 282821 309394 282873
rect 309406 282821 309458 282873
rect 309150 282757 309202 282809
rect 309214 282757 309266 282809
rect 309278 282757 309330 282809
rect 309342 282757 309394 282809
rect 309406 282757 309458 282809
rect 309150 282693 309202 282745
rect 309214 282693 309266 282745
rect 309278 282693 309330 282745
rect 309342 282693 309394 282745
rect 309406 282693 309458 282745
rect 303882 282187 303934 282239
rect 303946 282187 303998 282239
rect 304010 282187 304062 282239
rect 304074 282187 304126 282239
rect 304138 282187 304190 282239
rect 303882 282123 303934 282175
rect 303946 282123 303998 282175
rect 304010 282123 304062 282175
rect 304074 282123 304126 282175
rect 304138 282123 304190 282175
rect 303882 282059 303934 282111
rect 303946 282059 303998 282111
rect 304010 282059 304062 282111
rect 304074 282059 304126 282111
rect 304138 282059 304190 282111
rect 310882 282140 310934 282192
rect 310946 282140 310998 282192
rect 311010 282140 311062 282192
rect 311074 282140 311126 282192
rect 311138 282140 311190 282192
rect 299112 282004 299164 282056
rect 302424 282004 302476 282056
rect 303882 281995 303934 282047
rect 303946 281995 303998 282047
rect 304010 281995 304062 282047
rect 304074 281995 304126 282047
rect 304138 281995 304190 282047
rect 305736 282004 305788 282056
rect 308956 282035 309008 282087
rect 310882 282076 310934 282128
rect 310946 282076 310998 282128
rect 311010 282076 311062 282128
rect 311074 282076 311126 282128
rect 311138 282076 311190 282128
rect 310882 282012 310934 282064
rect 310946 282012 310998 282064
rect 311010 282012 311062 282064
rect 311074 282012 311126 282064
rect 311138 282012 311190 282064
rect 303882 281931 303934 281983
rect 303946 281931 303998 281983
rect 304010 281931 304062 281983
rect 304074 281931 304126 281983
rect 304138 281931 304190 281983
rect 303882 281867 303934 281919
rect 303946 281867 303998 281919
rect 304010 281867 304062 281919
rect 304074 281867 304126 281919
rect 304138 281867 304190 281919
rect 303882 281803 303934 281855
rect 303946 281803 303998 281855
rect 304010 281803 304062 281855
rect 304074 281803 304126 281855
rect 304138 281803 304190 281855
rect 303882 281739 303934 281791
rect 303946 281739 303998 281791
rect 304010 281739 304062 281791
rect 304074 281739 304126 281791
rect 304138 281739 304190 281791
rect 303882 281675 303934 281727
rect 303946 281675 303998 281727
rect 304010 281675 304062 281727
rect 304074 281675 304126 281727
rect 304138 281675 304190 281727
rect 303882 281611 303934 281663
rect 303946 281611 303998 281663
rect 304010 281611 304062 281663
rect 304074 281611 304126 281663
rect 304138 281611 304190 281663
rect 312544 282004 312596 282056
rect 310882 281948 310934 282000
rect 310946 281948 310998 282000
rect 311010 281948 311062 282000
rect 311074 281948 311126 282000
rect 311138 281948 311190 282000
rect 310882 281884 310934 281936
rect 310946 281884 310998 281936
rect 311010 281884 311062 281936
rect 311074 281884 311126 281936
rect 311138 281884 311190 281936
rect 310882 281820 310934 281872
rect 310946 281820 310998 281872
rect 311010 281820 311062 281872
rect 311074 281820 311126 281872
rect 311138 281820 311190 281872
rect 310882 281756 310934 281808
rect 310946 281756 310998 281808
rect 311010 281756 311062 281808
rect 311074 281756 311126 281808
rect 311138 281756 311190 281808
rect 310882 281692 310934 281744
rect 310946 281692 310998 281744
rect 311010 281692 311062 281744
rect 311074 281692 311126 281744
rect 311138 281692 311190 281744
rect 310882 281628 310934 281680
rect 310946 281628 310998 281680
rect 311010 281628 311062 281680
rect 311074 281628 311126 281680
rect 311138 281628 311190 281680
rect 298192 262692 298244 262744
rect 299296 262692 299348 262744
rect 305092 262692 305144 262744
rect 308772 262692 308824 262744
rect 292488 262420 292540 262472
rect 312728 262216 312780 262268
rect 313004 262216 313056 262268
rect 302150 261948 302202 262000
rect 302214 261948 302266 262000
rect 302278 261948 302330 262000
rect 302342 261948 302394 262000
rect 302406 261948 302458 262000
rect 302150 261884 302202 261936
rect 302214 261884 302266 261936
rect 302278 261884 302330 261936
rect 302342 261884 302394 261936
rect 302406 261884 302458 261936
rect 302150 261820 302202 261872
rect 302214 261820 302266 261872
rect 302278 261820 302330 261872
rect 302342 261820 302394 261872
rect 302406 261820 302458 261872
rect 302150 261756 302202 261808
rect 302214 261756 302266 261808
rect 302278 261756 302330 261808
rect 302342 261756 302394 261808
rect 302406 261756 302458 261808
rect 302150 261692 302202 261744
rect 302214 261692 302266 261744
rect 302278 261692 302330 261744
rect 302342 261692 302394 261744
rect 302406 261692 302458 261744
rect 309150 261948 309202 262000
rect 309214 261948 309266 262000
rect 309278 261948 309330 262000
rect 309342 261948 309394 262000
rect 309406 261948 309458 262000
rect 309150 261884 309202 261936
rect 309214 261884 309266 261936
rect 309278 261884 309330 261936
rect 309342 261884 309394 261936
rect 309406 261884 309458 261936
rect 309150 261820 309202 261872
rect 309214 261820 309266 261872
rect 309278 261820 309330 261872
rect 309342 261820 309394 261872
rect 309406 261820 309458 261872
rect 309150 261756 309202 261808
rect 309214 261756 309266 261808
rect 309278 261756 309330 261808
rect 309342 261756 309394 261808
rect 309406 261756 309458 261808
rect 309150 261692 309202 261744
rect 309214 261692 309266 261744
rect 309278 261692 309330 261744
rect 309342 261692 309394 261744
rect 309406 261692 309458 261744
rect 303882 261187 303934 261239
rect 303946 261187 303998 261239
rect 304010 261187 304062 261239
rect 304074 261187 304126 261239
rect 304138 261187 304190 261239
rect 303882 261123 303934 261175
rect 303946 261123 303998 261175
rect 304010 261123 304062 261175
rect 304074 261123 304126 261175
rect 304138 261123 304190 261175
rect 303882 261059 303934 261111
rect 303946 261059 303998 261111
rect 304010 261059 304062 261111
rect 304074 261059 304126 261111
rect 304138 261059 304190 261111
rect 302608 260992 302660 261044
rect 303882 260995 303934 261047
rect 303946 260995 303998 261047
rect 304010 260995 304062 261047
rect 304074 260995 304126 261047
rect 304138 260995 304190 261047
rect 303882 260931 303934 260983
rect 303946 260931 303998 260983
rect 304010 260931 304062 260983
rect 304074 260931 304126 260983
rect 304138 260931 304190 260983
rect 303882 260867 303934 260919
rect 303946 260867 303998 260919
rect 304010 260867 304062 260919
rect 304074 260867 304126 260919
rect 304138 260867 304190 260919
rect 303882 260803 303934 260855
rect 303946 260803 303998 260855
rect 304010 260803 304062 260855
rect 304074 260803 304126 260855
rect 304138 260803 304190 260855
rect 303882 260739 303934 260791
rect 303946 260739 303998 260791
rect 304010 260739 304062 260791
rect 304074 260739 304126 260791
rect 304138 260739 304190 260791
rect 303882 260675 303934 260727
rect 303946 260675 303998 260727
rect 304010 260675 304062 260727
rect 304074 260675 304126 260727
rect 304138 260675 304190 260727
rect 303882 260611 303934 260663
rect 303946 260611 303998 260663
rect 304010 260611 304062 260663
rect 304074 260611 304126 260663
rect 304138 260611 304190 260663
rect 296882 242034 296934 242086
rect 296946 242034 296998 242086
rect 297010 242034 297062 242086
rect 297074 242034 297126 242086
rect 297138 242034 297190 242086
rect 296882 241970 296934 242022
rect 296946 241970 296998 242022
rect 297010 241970 297062 242022
rect 297074 241970 297126 242022
rect 297138 241970 297190 242022
rect 296882 241906 296934 241958
rect 296946 241906 296998 241958
rect 297010 241906 297062 241958
rect 297074 241906 297126 241958
rect 297138 241906 297190 241958
rect 296882 241842 296934 241894
rect 296946 241842 296998 241894
rect 297010 241842 297062 241894
rect 297074 241842 297126 241894
rect 297138 241842 297190 241894
rect 296882 241778 296934 241830
rect 296946 241778 296998 241830
rect 297010 241778 297062 241830
rect 297074 241778 297126 241830
rect 297138 241778 297190 241830
rect 303882 242034 303934 242086
rect 303946 242034 303998 242086
rect 304010 242034 304062 242086
rect 304074 242034 304126 242086
rect 304138 242034 304190 242086
rect 303882 241970 303934 242022
rect 303946 241970 303998 242022
rect 304010 241970 304062 242022
rect 304074 241970 304126 242022
rect 304138 241970 304190 242022
rect 303882 241906 303934 241958
rect 303946 241906 303998 241958
rect 304010 241906 304062 241958
rect 304074 241906 304126 241958
rect 304138 241906 304190 241958
rect 303882 241842 303934 241894
rect 303946 241842 303998 241894
rect 304010 241842 304062 241894
rect 304074 241842 304126 241894
rect 304138 241842 304190 241894
rect 303882 241778 303934 241830
rect 303946 241778 303998 241830
rect 304010 241778 304062 241830
rect 304074 241778 304126 241830
rect 304138 241778 304190 241830
rect 310882 242034 310934 242086
rect 310946 242034 310998 242086
rect 311010 242034 311062 242086
rect 311074 242034 311126 242086
rect 311138 242034 311190 242086
rect 310882 241970 310934 242022
rect 310946 241970 310998 242022
rect 311010 241970 311062 242022
rect 311074 241970 311126 242022
rect 311138 241970 311190 242022
rect 310882 241906 310934 241958
rect 310946 241906 310998 241958
rect 311010 241906 311062 241958
rect 311074 241906 311126 241958
rect 311138 241906 311190 241958
rect 310882 241842 310934 241894
rect 310946 241842 310998 241894
rect 311010 241842 311062 241894
rect 311074 241842 311126 241894
rect 311138 241842 311190 241894
rect 310882 241778 310934 241830
rect 310946 241778 310998 241830
rect 311010 241778 311062 241830
rect 311074 241778 311126 241830
rect 311138 241778 311190 241830
rect 311072 241612 311124 241664
rect 312452 241612 312504 241664
rect 314384 241612 314436 241664
rect 292488 241408 292540 241460
rect 296904 241237 296956 241289
rect 300952 241237 301004 241289
rect 295248 241136 295300 241188
rect 296904 241136 296956 241188
rect 295150 240949 295202 241001
rect 295214 240949 295266 241001
rect 295278 240949 295330 241001
rect 295342 240949 295394 241001
rect 295406 240949 295458 241001
rect 295150 240885 295202 240937
rect 295214 240885 295266 240937
rect 295278 240885 295330 240937
rect 295342 240885 295394 240937
rect 295406 240885 295458 240937
rect 295150 240821 295202 240873
rect 295214 240821 295266 240873
rect 295278 240821 295330 240873
rect 295342 240821 295394 240873
rect 295406 240821 295458 240873
rect 295150 240757 295202 240809
rect 295214 240757 295266 240809
rect 295278 240757 295330 240809
rect 295342 240757 295394 240809
rect 295406 240757 295458 240809
rect 295150 240693 295202 240745
rect 295214 240693 295266 240745
rect 295278 240693 295330 240745
rect 295342 240693 295394 240745
rect 295406 240693 295458 240745
rect 309150 240923 309202 240975
rect 309214 240923 309266 240975
rect 309278 240923 309330 240975
rect 309342 240923 309394 240975
rect 309406 240923 309458 240975
rect 309150 240859 309202 240911
rect 309214 240859 309266 240911
rect 309278 240859 309330 240911
rect 309342 240859 309394 240911
rect 309406 240859 309458 240911
rect 309150 240795 309202 240847
rect 309214 240795 309266 240847
rect 309278 240795 309330 240847
rect 309342 240795 309394 240847
rect 309406 240795 309458 240847
rect 309150 240731 309202 240783
rect 309214 240731 309266 240783
rect 309278 240731 309330 240783
rect 309342 240731 309394 240783
rect 309406 240731 309458 240783
rect 309150 240667 309202 240719
rect 309214 240667 309266 240719
rect 309278 240667 309330 240719
rect 309342 240667 309394 240719
rect 309406 240667 309458 240719
rect 302148 240499 302200 240508
rect 302148 240465 302159 240499
rect 302159 240465 302200 240499
rect 302148 240456 302200 240465
rect 312544 240524 312596 240576
rect 308680 240499 308732 240508
rect 308680 240465 308689 240499
rect 308689 240465 308732 240499
rect 308680 240456 308732 240465
rect 298836 240033 298888 240085
rect 305368 240033 305420 240085
rect 514760 240048 514812 240100
rect 310882 239862 310934 239914
rect 310946 239862 310998 239914
rect 311010 239862 311062 239914
rect 311074 239862 311126 239914
rect 311138 239862 311190 239914
rect 310882 239798 310934 239850
rect 310946 239798 310998 239850
rect 311010 239798 311062 239850
rect 311074 239798 311126 239850
rect 311138 239798 311190 239850
rect 310882 239734 310934 239786
rect 310946 239734 310998 239786
rect 311010 239734 311062 239786
rect 311074 239734 311126 239786
rect 311138 239734 311190 239786
rect 310882 239670 310934 239722
rect 310946 239670 310998 239722
rect 311010 239670 311062 239722
rect 311074 239670 311126 239722
rect 311138 239670 311190 239722
rect 310882 239606 310934 239658
rect 310946 239606 310998 239658
rect 311010 239606 311062 239658
rect 311074 239606 311126 239658
rect 311138 239606 311190 239658
rect 308680 238688 308732 238740
rect 376024 238688 376076 238740
rect 298836 238620 298888 238672
rect 316868 238620 316920 238672
rect 302148 238552 302200 238604
rect 313924 238552 313976 238604
rect 305368 238484 305420 238536
rect 314292 238484 314344 238536
rect 296882 221035 296934 221087
rect 296946 221035 296998 221087
rect 297010 221035 297062 221087
rect 297074 221035 297126 221087
rect 297138 221035 297190 221087
rect 296882 220971 296934 221023
rect 296946 220971 296998 221023
rect 297010 220971 297062 221023
rect 297074 220971 297126 221023
rect 297138 220971 297190 221023
rect 296882 220907 296934 220959
rect 296946 220907 296998 220959
rect 297010 220907 297062 220959
rect 297074 220907 297126 220959
rect 297138 220907 297190 220959
rect 296882 220843 296934 220895
rect 296946 220843 296998 220895
rect 297010 220843 297062 220895
rect 297074 220843 297126 220895
rect 297138 220843 297190 220895
rect 296882 220779 296934 220831
rect 296946 220779 296998 220831
rect 297010 220779 297062 220831
rect 297074 220779 297126 220831
rect 297138 220779 297190 220831
rect 303882 221035 303934 221087
rect 303946 221035 303998 221087
rect 304010 221035 304062 221087
rect 304074 221035 304126 221087
rect 304138 221035 304190 221087
rect 303882 220971 303934 221023
rect 303946 220971 303998 221023
rect 304010 220971 304062 221023
rect 304074 220971 304126 221023
rect 304138 220971 304190 221023
rect 303882 220907 303934 220959
rect 303946 220907 303998 220959
rect 304010 220907 304062 220959
rect 304074 220907 304126 220959
rect 304138 220907 304190 220959
rect 303882 220843 303934 220895
rect 303946 220843 303998 220895
rect 304010 220843 304062 220895
rect 304074 220843 304126 220895
rect 304138 220843 304190 220895
rect 303882 220779 303934 220831
rect 303946 220779 303998 220831
rect 304010 220779 304062 220831
rect 304074 220779 304126 220831
rect 304138 220779 304190 220831
rect 310882 221035 310934 221087
rect 310946 221035 310998 221087
rect 311010 221035 311062 221087
rect 311074 221035 311126 221087
rect 311138 221035 311190 221087
rect 310882 220971 310934 221023
rect 310946 220971 310998 221023
rect 311010 220971 311062 221023
rect 311074 220971 311126 221023
rect 311138 220971 311190 221023
rect 310882 220907 310934 220959
rect 310946 220907 310998 220959
rect 311010 220907 311062 220959
rect 311074 220907 311126 220959
rect 311138 220907 311190 220959
rect 310882 220843 310934 220895
rect 310946 220843 310998 220895
rect 311010 220843 311062 220895
rect 311074 220843 311126 220895
rect 311138 220843 311190 220895
rect 310882 220779 310934 220831
rect 310946 220779 310998 220831
rect 311010 220779 311062 220831
rect 311074 220779 311126 220831
rect 311138 220779 311190 220831
rect 292488 220464 292540 220516
rect 294972 220464 295024 220516
rect 313924 220260 313976 220312
rect 314384 220260 314436 220312
rect 295150 219950 295202 220002
rect 295214 219950 295266 220002
rect 295278 219950 295330 220002
rect 295342 219950 295394 220002
rect 295406 219950 295458 220002
rect 295150 219886 295202 219938
rect 295214 219886 295266 219938
rect 295278 219886 295330 219938
rect 295342 219886 295394 219938
rect 295406 219886 295458 219938
rect 295150 219822 295202 219874
rect 295214 219822 295266 219874
rect 295278 219822 295330 219874
rect 295342 219822 295394 219874
rect 295406 219822 295458 219874
rect 295150 219758 295202 219810
rect 295214 219758 295266 219810
rect 295278 219758 295330 219810
rect 295342 219758 295394 219810
rect 295406 219758 295458 219810
rect 295150 219694 295202 219746
rect 295214 219694 295266 219746
rect 295278 219694 295330 219746
rect 295342 219694 295394 219746
rect 295406 219694 295458 219746
rect 302150 219949 302202 220001
rect 302214 219949 302266 220001
rect 302278 219949 302330 220001
rect 302342 219949 302394 220001
rect 302406 219949 302458 220001
rect 302150 219885 302202 219937
rect 302214 219885 302266 219937
rect 302278 219885 302330 219937
rect 302342 219885 302394 219937
rect 302406 219885 302458 219937
rect 302150 219821 302202 219873
rect 302214 219821 302266 219873
rect 302278 219821 302330 219873
rect 302342 219821 302394 219873
rect 302406 219821 302458 219873
rect 302150 219757 302202 219809
rect 302214 219757 302266 219809
rect 302278 219757 302330 219809
rect 302342 219757 302394 219809
rect 302406 219757 302458 219809
rect 302150 219693 302202 219745
rect 302214 219693 302266 219745
rect 302278 219693 302330 219745
rect 302342 219693 302394 219745
rect 302406 219693 302458 219745
rect 309150 219949 309202 220001
rect 309214 219949 309266 220001
rect 309278 219949 309330 220001
rect 309342 219949 309394 220001
rect 309406 219949 309458 220001
rect 309150 219885 309202 219937
rect 309214 219885 309266 219937
rect 309278 219885 309330 219937
rect 309342 219885 309394 219937
rect 309406 219885 309458 219937
rect 309150 219821 309202 219873
rect 309214 219821 309266 219873
rect 309278 219821 309330 219873
rect 309342 219821 309394 219873
rect 309406 219821 309458 219873
rect 309150 219757 309202 219809
rect 309214 219757 309266 219809
rect 309278 219757 309330 219809
rect 309342 219757 309394 219809
rect 309406 219757 309458 219809
rect 309150 219693 309202 219745
rect 309214 219693 309266 219745
rect 309278 219693 309330 219745
rect 309342 219693 309394 219745
rect 309406 219693 309458 219745
rect 311045 219461 311097 219513
rect 303965 219344 304017 219396
rect 299296 219033 299348 219085
rect 303160 219036 303212 219088
rect 306748 219033 306800 219085
rect 310428 219033 310480 219085
rect 292488 206252 292540 206304
rect 580172 206252 580224 206304
rect 295248 199316 295300 199368
rect 292488 199248 292540 199300
rect 311072 198432 311124 198484
rect 311256 198432 311308 198484
rect 307668 198364 307720 198416
rect 296882 179235 296934 179287
rect 296946 179235 296998 179287
rect 297010 179235 297062 179287
rect 297074 179235 297126 179287
rect 297138 179235 297190 179287
rect 296882 179171 296934 179223
rect 296946 179171 296998 179223
rect 297010 179171 297062 179223
rect 297074 179171 297126 179223
rect 297138 179171 297190 179223
rect 296882 179107 296934 179159
rect 296946 179107 296998 179159
rect 297010 179107 297062 179159
rect 297074 179107 297126 179159
rect 297138 179107 297190 179159
rect 296882 179043 296934 179095
rect 296946 179043 296998 179095
rect 297010 179043 297062 179095
rect 297074 179043 297126 179095
rect 297138 179043 297190 179095
rect 296882 178979 296934 179031
rect 296946 178979 296998 179031
rect 297010 178979 297062 179031
rect 297074 178979 297126 179031
rect 297138 178979 297190 179031
rect 303882 179235 303934 179287
rect 303946 179235 303998 179287
rect 304010 179235 304062 179287
rect 304074 179235 304126 179287
rect 304138 179235 304190 179287
rect 303882 179171 303934 179223
rect 303946 179171 303998 179223
rect 304010 179171 304062 179223
rect 304074 179171 304126 179223
rect 304138 179171 304190 179223
rect 303882 179107 303934 179159
rect 303946 179107 303998 179159
rect 304010 179107 304062 179159
rect 304074 179107 304126 179159
rect 304138 179107 304190 179159
rect 303882 179043 303934 179095
rect 303946 179043 303998 179095
rect 304010 179043 304062 179095
rect 304074 179043 304126 179095
rect 304138 179043 304190 179095
rect 303882 178979 303934 179031
rect 303946 178979 303998 179031
rect 304010 178979 304062 179031
rect 304074 178979 304126 179031
rect 304138 178979 304190 179031
rect 310894 179235 310946 179287
rect 310894 179171 310946 179223
rect 310894 179107 310946 179159
rect 310894 179043 310946 179095
rect 310894 178979 310946 179031
rect 292488 178712 292540 178764
rect 297272 178438 297324 178490
rect 295150 178149 295202 178201
rect 295214 178149 295266 178201
rect 295278 178149 295330 178201
rect 295342 178149 295394 178201
rect 295406 178149 295458 178201
rect 295150 178085 295202 178137
rect 295214 178085 295266 178137
rect 295278 178085 295330 178137
rect 295342 178085 295394 178137
rect 295406 178085 295458 178137
rect 295150 178021 295202 178073
rect 295214 178021 295266 178073
rect 295278 178021 295330 178073
rect 295342 178021 295394 178073
rect 295406 178021 295458 178073
rect 295150 177957 295202 178009
rect 295214 177957 295266 178009
rect 295278 177957 295330 178009
rect 295342 177957 295394 178009
rect 295406 177957 295458 178009
rect 295150 177893 295202 177945
rect 295214 177893 295266 177945
rect 295278 177893 295330 177945
rect 295342 177893 295394 177945
rect 295406 177893 295458 177945
rect 302150 178133 302202 178185
rect 302214 178133 302266 178185
rect 302278 178133 302330 178185
rect 302342 178133 302394 178185
rect 302406 178133 302458 178185
rect 302150 178069 302202 178121
rect 302214 178069 302266 178121
rect 302278 178069 302330 178121
rect 302342 178069 302394 178121
rect 302406 178069 302458 178121
rect 302150 178005 302202 178057
rect 302214 178005 302266 178057
rect 302278 178005 302330 178057
rect 302342 178005 302394 178057
rect 302406 178005 302458 178057
rect 302150 177941 302202 177993
rect 302214 177941 302266 177993
rect 302278 177941 302330 177993
rect 302342 177941 302394 177993
rect 302406 177941 302458 177993
rect 302150 177877 302202 177929
rect 302214 177877 302266 177929
rect 302278 177877 302330 177929
rect 302342 177877 302394 177929
rect 302406 177877 302458 177929
rect 309150 178133 309202 178185
rect 309214 178133 309266 178185
rect 309278 178133 309330 178185
rect 309342 178133 309394 178185
rect 309406 178133 309458 178185
rect 309150 178069 309202 178121
rect 309214 178069 309266 178121
rect 309278 178069 309330 178121
rect 309342 178069 309394 178121
rect 309406 178069 309458 178121
rect 309150 178005 309202 178057
rect 309214 178005 309266 178057
rect 309278 178005 309330 178057
rect 309342 178005 309394 178057
rect 309406 178005 309458 178057
rect 309150 177941 309202 177993
rect 309214 177941 309266 177993
rect 309278 177941 309330 177993
rect 309342 177941 309394 177993
rect 309406 177941 309458 177993
rect 309150 177877 309202 177929
rect 309214 177877 309266 177929
rect 309278 177877 309330 177929
rect 309342 177877 309394 177929
rect 309406 177877 309458 177929
rect 311256 177624 311308 177676
rect 311532 177624 311584 177676
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 304446 492824 304502 492833
rect 304446 492759 304502 492768
rect 311990 492824 312046 492833
rect 311990 492759 312046 492768
rect 295062 491872 295118 491881
rect 295062 491807 295118 491816
rect 292488 490748 292540 490754
rect 292488 490690 292540 490696
rect 292500 472394 292528 490690
rect 294880 490680 294932 490686
rect 294880 490622 294932 490628
rect 293866 474056 293922 474065
rect 293866 473991 293922 474000
rect 292488 472388 292540 472394
rect 292488 472330 292540 472336
rect 292500 451382 292528 472330
rect 292488 451376 292540 451382
rect 292488 451318 292540 451324
rect 292500 430302 292528 451318
rect 293880 449177 293908 473991
rect 294892 472598 294920 490622
rect 295076 474065 295104 491807
rect 296882 491656 297190 491662
rect 296934 491650 296946 491656
rect 296998 491650 297010 491656
rect 297062 491650 297074 491656
rect 297126 491650 297138 491656
rect 296944 491604 296946 491650
rect 297126 491604 297128 491650
rect 296882 491594 296888 491604
rect 296944 491594 296968 491604
rect 297024 491594 297048 491604
rect 297104 491594 297128 491604
rect 297184 491594 297190 491604
rect 296882 491592 297190 491594
rect 296934 491570 296946 491592
rect 296998 491570 297010 491592
rect 297062 491570 297074 491592
rect 297126 491570 297138 491592
rect 296944 491540 296946 491570
rect 297126 491540 297128 491570
rect 296882 491528 296888 491540
rect 296944 491528 296968 491540
rect 297024 491528 297048 491540
rect 297104 491528 297128 491540
rect 297184 491528 297190 491540
rect 296944 491514 296946 491528
rect 297126 491514 297128 491528
rect 296934 491490 296946 491514
rect 296998 491490 297010 491514
rect 297062 491490 297074 491514
rect 297126 491490 297138 491514
rect 296944 491476 296946 491490
rect 297126 491476 297128 491490
rect 296882 491464 296888 491476
rect 296944 491464 296968 491476
rect 297024 491464 297048 491476
rect 297104 491464 297128 491476
rect 297184 491464 297190 491476
rect 296944 491434 296946 491464
rect 297126 491434 297128 491464
rect 296934 491412 296946 491434
rect 296998 491412 297010 491434
rect 297062 491412 297074 491434
rect 297126 491412 297138 491434
rect 296882 491410 297190 491412
rect 296882 491400 296888 491410
rect 296944 491400 296968 491410
rect 297024 491400 297048 491410
rect 297104 491400 297128 491410
rect 297184 491400 297190 491410
rect 296944 491354 296946 491400
rect 297126 491354 297128 491400
rect 296934 491348 296946 491354
rect 296998 491348 297010 491354
rect 297062 491348 297074 491354
rect 297126 491348 297138 491354
rect 296882 491342 297190 491348
rect 303882 491656 304190 491662
rect 303934 491650 303946 491656
rect 303998 491650 304010 491656
rect 304062 491650 304074 491656
rect 304126 491650 304138 491656
rect 303944 491604 303946 491650
rect 304126 491604 304128 491650
rect 303882 491594 303888 491604
rect 303944 491594 303968 491604
rect 304024 491594 304048 491604
rect 304104 491594 304128 491604
rect 304184 491594 304190 491604
rect 303882 491592 304190 491594
rect 303934 491570 303946 491592
rect 303998 491570 304010 491592
rect 304062 491570 304074 491592
rect 304126 491570 304138 491592
rect 303944 491540 303946 491570
rect 304126 491540 304128 491570
rect 303882 491528 303888 491540
rect 303944 491528 303968 491540
rect 304024 491528 304048 491540
rect 304104 491528 304128 491540
rect 304184 491528 304190 491540
rect 303944 491514 303946 491528
rect 304126 491514 304128 491528
rect 303934 491490 303946 491514
rect 303998 491490 304010 491514
rect 304062 491490 304074 491514
rect 304126 491490 304138 491514
rect 303944 491476 303946 491490
rect 304126 491476 304128 491490
rect 303882 491464 303888 491476
rect 303944 491464 303968 491476
rect 304024 491464 304048 491476
rect 304104 491464 304128 491476
rect 304184 491464 304190 491476
rect 304460 491473 304488 492759
rect 310882 491656 311190 491662
rect 310934 491650 310946 491656
rect 310998 491650 311010 491656
rect 311062 491650 311074 491656
rect 311126 491650 311138 491656
rect 310944 491604 310946 491650
rect 311126 491604 311128 491650
rect 310882 491594 310888 491604
rect 310944 491594 310968 491604
rect 311024 491594 311048 491604
rect 311104 491594 311128 491604
rect 311184 491594 311190 491604
rect 310882 491592 311190 491594
rect 310934 491570 310946 491592
rect 310998 491570 311010 491592
rect 311062 491570 311074 491592
rect 311126 491570 311138 491592
rect 310944 491540 310946 491570
rect 311126 491540 311128 491570
rect 310882 491528 310888 491540
rect 310944 491528 310968 491540
rect 311024 491528 311048 491540
rect 311104 491528 311128 491540
rect 311184 491528 311190 491540
rect 310944 491514 310946 491528
rect 311126 491514 311128 491528
rect 310934 491490 310946 491514
rect 310998 491490 311010 491514
rect 311062 491490 311074 491514
rect 311126 491490 311138 491514
rect 310944 491476 310946 491490
rect 311126 491476 311128 491490
rect 303944 491434 303946 491464
rect 304126 491434 304128 491464
rect 303934 491412 303946 491434
rect 303998 491412 304010 491434
rect 304062 491412 304074 491434
rect 304126 491412 304138 491434
rect 303882 491410 304190 491412
rect 303882 491400 303888 491410
rect 303944 491400 303968 491410
rect 304024 491400 304048 491410
rect 304104 491400 304128 491410
rect 304184 491400 304190 491410
rect 303944 491354 303946 491400
rect 304126 491354 304128 491400
rect 304446 491464 304502 491473
rect 304446 491399 304502 491408
rect 310882 491464 310888 491476
rect 310944 491464 310968 491476
rect 311024 491464 311048 491476
rect 311104 491464 311128 491476
rect 311184 491464 311190 491476
rect 310944 491434 310946 491464
rect 311126 491434 311128 491464
rect 310934 491412 310946 491434
rect 310998 491412 311010 491434
rect 311062 491412 311074 491434
rect 311126 491412 311138 491434
rect 310882 491410 311190 491412
rect 310882 491400 310888 491410
rect 310944 491400 310968 491410
rect 311024 491400 311048 491410
rect 311104 491400 311128 491410
rect 311184 491400 311190 491410
rect 303934 491348 303946 491354
rect 303998 491348 304010 491354
rect 304062 491348 304074 491354
rect 304126 491348 304138 491354
rect 303882 491342 304190 491348
rect 310944 491354 310946 491400
rect 311126 491354 311128 491400
rect 310934 491348 310946 491354
rect 310998 491348 311010 491354
rect 311062 491348 311074 491354
rect 311126 491348 311138 491354
rect 310882 491342 311190 491348
rect 300858 491192 300914 491201
rect 300858 491127 300914 491136
rect 296996 490859 297048 490865
rect 296996 490801 297048 490807
rect 297008 490686 297036 490801
rect 300872 490770 300900 491127
rect 304221 491056 304277 491065
rect 304221 490991 304277 491000
rect 300872 490742 301094 490770
rect 304235 490756 304263 490991
rect 296996 490680 297048 490686
rect 296996 490622 297048 490628
rect 295150 490548 295458 490554
rect 295202 490534 295214 490548
rect 295266 490534 295278 490548
rect 295330 490534 295342 490548
rect 295394 490534 295406 490548
rect 295212 490496 295214 490534
rect 295394 490496 295396 490534
rect 295150 490484 295156 490496
rect 295212 490484 295236 490496
rect 295292 490484 295316 490496
rect 295372 490484 295396 490496
rect 295452 490484 295458 490496
rect 295212 490478 295214 490484
rect 295394 490478 295396 490484
rect 295202 490454 295214 490478
rect 295266 490454 295278 490478
rect 295330 490454 295342 490478
rect 295394 490454 295406 490478
rect 295212 490432 295214 490454
rect 295394 490432 295396 490454
rect 295150 490420 295156 490432
rect 295212 490420 295236 490432
rect 295292 490420 295316 490432
rect 295372 490420 295396 490432
rect 295452 490420 295458 490432
rect 295212 490398 295214 490420
rect 295394 490398 295396 490420
rect 295202 490374 295214 490398
rect 295266 490374 295278 490398
rect 295330 490374 295342 490398
rect 295394 490374 295406 490398
rect 295212 490368 295214 490374
rect 295394 490368 295396 490374
rect 295150 490356 295156 490368
rect 295212 490356 295236 490368
rect 295292 490356 295316 490368
rect 295372 490356 295396 490368
rect 295452 490356 295458 490368
rect 295212 490318 295214 490356
rect 295394 490318 295396 490356
rect 295202 490304 295214 490318
rect 295266 490304 295278 490318
rect 295330 490304 295342 490318
rect 295394 490304 295406 490318
rect 295150 490298 295458 490304
rect 305092 490068 305144 490074
rect 305092 490010 305144 490016
rect 298744 489796 298796 489802
rect 298744 489738 298796 489744
rect 298756 486441 298784 489738
rect 301780 489655 301832 489661
rect 301780 489597 301832 489603
rect 301792 486577 301820 489597
rect 303882 489484 304190 489490
rect 303934 489478 303946 489484
rect 303998 489478 304010 489484
rect 304062 489478 304074 489484
rect 304126 489478 304138 489484
rect 303944 489432 303946 489478
rect 304126 489432 304128 489478
rect 303882 489422 303888 489432
rect 303944 489422 303968 489432
rect 304024 489422 304048 489432
rect 304104 489422 304128 489432
rect 304184 489422 304190 489432
rect 303882 489420 304190 489422
rect 303934 489398 303946 489420
rect 303998 489398 304010 489420
rect 304062 489398 304074 489420
rect 304126 489398 304138 489420
rect 303944 489368 303946 489398
rect 304126 489368 304128 489398
rect 303882 489356 303888 489368
rect 303944 489356 303968 489368
rect 304024 489356 304048 489368
rect 304104 489356 304128 489368
rect 304184 489356 304190 489368
rect 303944 489342 303946 489356
rect 304126 489342 304128 489356
rect 303934 489318 303946 489342
rect 303998 489318 304010 489342
rect 304062 489318 304074 489342
rect 304126 489318 304138 489342
rect 303944 489304 303946 489318
rect 304126 489304 304128 489318
rect 303882 489292 303888 489304
rect 303944 489292 303968 489304
rect 304024 489292 304048 489304
rect 304104 489292 304128 489304
rect 304184 489292 304190 489304
rect 303944 489262 303946 489292
rect 304126 489262 304128 489292
rect 303934 489240 303946 489262
rect 303998 489240 304010 489262
rect 304062 489240 304074 489262
rect 304126 489240 304138 489262
rect 303882 489238 304190 489240
rect 303882 489228 303888 489238
rect 303944 489228 303968 489238
rect 304024 489228 304048 489238
rect 304104 489228 304128 489238
rect 304184 489228 304190 489238
rect 303944 489182 303946 489228
rect 304126 489182 304128 489228
rect 303934 489176 303946 489182
rect 303998 489176 304010 489182
rect 304062 489176 304074 489182
rect 304126 489176 304138 489182
rect 303882 489170 304190 489176
rect 305104 486713 305132 490010
rect 310549 489914 310577 490076
rect 310532 489886 310577 489914
rect 308128 489728 308180 489734
rect 308128 489670 308180 489676
rect 305090 486704 305146 486713
rect 305090 486639 305146 486648
rect 301778 486568 301834 486577
rect 301778 486503 301834 486512
rect 298742 486432 298798 486441
rect 298742 486367 298798 486376
rect 305550 474736 305606 474745
rect 305550 474671 305606 474680
rect 295062 474056 295118 474065
rect 295062 473991 295118 474000
rect 301410 474056 301466 474065
rect 301410 473991 301466 474000
rect 296882 473116 297190 473122
rect 296934 473110 296946 473116
rect 296998 473110 297010 473116
rect 297062 473110 297074 473116
rect 297126 473110 297138 473116
rect 296944 473064 296946 473110
rect 297126 473064 297128 473110
rect 296882 473054 296888 473064
rect 296944 473054 296968 473064
rect 297024 473054 297048 473064
rect 297104 473054 297128 473064
rect 297184 473054 297190 473064
rect 296882 473052 297190 473054
rect 296934 473030 296946 473052
rect 296998 473030 297010 473052
rect 297062 473030 297074 473052
rect 297126 473030 297138 473052
rect 296944 473000 296946 473030
rect 297126 473000 297128 473030
rect 296882 472988 296888 473000
rect 296944 472988 296968 473000
rect 297024 472988 297048 473000
rect 297104 472988 297128 473000
rect 297184 472988 297190 473000
rect 296944 472974 296946 472988
rect 297126 472974 297128 472988
rect 301424 472977 301452 473991
rect 303882 473116 304190 473122
rect 303934 473110 303946 473116
rect 303998 473110 304010 473116
rect 304062 473110 304074 473116
rect 304126 473110 304138 473116
rect 303944 473064 303946 473110
rect 304126 473064 304128 473110
rect 303882 473054 303888 473064
rect 303944 473054 303968 473064
rect 304024 473054 304048 473064
rect 304104 473054 304128 473064
rect 304184 473054 304190 473064
rect 303882 473052 304190 473054
rect 303934 473030 303946 473052
rect 303998 473030 304010 473052
rect 304062 473030 304074 473052
rect 304126 473030 304138 473052
rect 303944 473000 303946 473030
rect 304126 473000 304128 473030
rect 303882 472988 303888 473000
rect 303944 472988 303968 473000
rect 304024 472988 304048 473000
rect 304104 472988 304128 473000
rect 304184 472988 304190 473000
rect 296934 472950 296946 472974
rect 296998 472950 297010 472974
rect 297062 472950 297074 472974
rect 297126 472950 297138 472974
rect 296944 472936 296946 472950
rect 297126 472936 297128 472950
rect 296882 472924 296888 472936
rect 296944 472924 296968 472936
rect 297024 472924 297048 472936
rect 297104 472924 297128 472936
rect 297184 472924 297190 472936
rect 296944 472894 296946 472924
rect 297126 472894 297128 472924
rect 301410 472968 301466 472977
rect 301410 472903 301466 472912
rect 303944 472974 303946 472988
rect 304126 472974 304128 472988
rect 305564 472977 305592 474671
rect 308140 474065 308168 489670
rect 308126 474056 308182 474065
rect 308126 473991 308182 474000
rect 310532 473385 310560 489886
rect 311530 489696 311586 489705
rect 311530 489631 311532 489640
rect 311584 489631 311586 489640
rect 311532 489597 311584 489603
rect 310882 489484 311190 489490
rect 310934 489478 310946 489484
rect 310998 489478 311010 489484
rect 311062 489478 311074 489484
rect 311126 489478 311138 489484
rect 310944 489432 310946 489478
rect 311126 489432 311128 489478
rect 310882 489422 310888 489432
rect 310944 489422 310968 489432
rect 311024 489422 311048 489432
rect 311104 489422 311128 489432
rect 311184 489422 311190 489432
rect 310882 489420 311190 489422
rect 310934 489398 310946 489420
rect 310998 489398 311010 489420
rect 311062 489398 311074 489420
rect 311126 489398 311138 489420
rect 310944 489368 310946 489398
rect 311126 489368 311128 489398
rect 310882 489356 310888 489368
rect 310944 489356 310968 489368
rect 311024 489356 311048 489368
rect 311104 489356 311128 489368
rect 311184 489356 311190 489368
rect 310944 489342 310946 489356
rect 311126 489342 311128 489356
rect 310934 489318 310946 489342
rect 310998 489318 311010 489342
rect 311062 489318 311074 489342
rect 311126 489318 311138 489342
rect 310944 489304 310946 489318
rect 311126 489304 311128 489318
rect 310882 489292 310888 489304
rect 310944 489292 310968 489304
rect 311024 489292 311048 489304
rect 311104 489292 311128 489304
rect 311184 489292 311190 489304
rect 310944 489262 310946 489292
rect 311126 489262 311128 489292
rect 310934 489240 310946 489262
rect 310998 489240 311010 489262
rect 311062 489240 311074 489262
rect 311126 489240 311138 489262
rect 310882 489238 311190 489240
rect 310882 489228 310888 489238
rect 310944 489228 310968 489238
rect 311024 489228 311048 489238
rect 311104 489228 311128 489238
rect 311184 489228 311190 489238
rect 310944 489182 310946 489228
rect 311126 489182 311128 489228
rect 310934 489176 310946 489182
rect 310998 489176 311010 489182
rect 311062 489176 311074 489182
rect 311126 489176 311138 489182
rect 310882 489170 311190 489176
rect 312004 474745 312032 492759
rect 312084 490204 312136 490210
rect 312084 490146 312136 490152
rect 312096 489914 312124 490146
rect 312096 489886 312216 489914
rect 311990 474736 312046 474745
rect 311990 474671 312046 474680
rect 312188 473521 312216 489886
rect 319442 489696 319498 489705
rect 319442 489631 319498 489640
rect 318338 486704 318394 486713
rect 318338 486639 318394 486648
rect 313646 474736 313702 474745
rect 313646 474671 313702 474680
rect 312174 473512 312230 473521
rect 312174 473447 312230 473456
rect 310518 473376 310574 473385
rect 310518 473311 310574 473320
rect 310882 473116 311190 473122
rect 310934 473110 310946 473116
rect 310998 473110 311010 473116
rect 311062 473110 311074 473116
rect 311126 473110 311138 473116
rect 310944 473064 310946 473110
rect 311126 473064 311128 473110
rect 310882 473054 310888 473064
rect 310944 473054 310968 473064
rect 311024 473054 311048 473064
rect 311104 473054 311128 473064
rect 311184 473054 311190 473064
rect 310882 473052 311190 473054
rect 310934 473030 310946 473052
rect 310998 473030 311010 473052
rect 311062 473030 311074 473052
rect 311126 473030 311138 473052
rect 310944 473000 310946 473030
rect 311126 473000 311128 473030
rect 310882 472988 310888 473000
rect 310944 472988 310968 473000
rect 311024 472988 311048 473000
rect 311104 472988 311128 473000
rect 311184 472988 311190 473000
rect 303934 472950 303946 472974
rect 303998 472950 304010 472974
rect 304062 472950 304074 472974
rect 304126 472950 304138 472974
rect 303944 472936 303946 472950
rect 304126 472936 304128 472950
rect 303882 472924 303888 472936
rect 303944 472924 303968 472936
rect 304024 472924 304048 472936
rect 304104 472924 304128 472936
rect 304184 472924 304190 472936
rect 296934 472872 296946 472894
rect 296998 472872 297010 472894
rect 297062 472872 297074 472894
rect 297126 472872 297138 472894
rect 296882 472870 297190 472872
rect 296882 472860 296888 472870
rect 296944 472860 296968 472870
rect 297024 472860 297048 472870
rect 297104 472860 297128 472870
rect 297184 472860 297190 472870
rect 296944 472814 296946 472860
rect 297126 472814 297128 472860
rect 296934 472808 296946 472814
rect 296998 472808 297010 472814
rect 297062 472808 297074 472814
rect 297126 472808 297138 472814
rect 296882 472802 297190 472808
rect 303944 472894 303946 472924
rect 304126 472894 304128 472924
rect 305550 472968 305606 472977
rect 305550 472903 305606 472912
rect 310944 472974 310946 472988
rect 311126 472974 311128 472988
rect 310934 472950 310946 472974
rect 310998 472950 311010 472974
rect 311062 472950 311074 472974
rect 311126 472950 311138 472974
rect 310944 472936 310946 472950
rect 311126 472936 311128 472950
rect 310882 472924 310888 472936
rect 310944 472924 310968 472936
rect 311024 472924 311048 472936
rect 311104 472924 311128 472936
rect 311184 472924 311190 472936
rect 303934 472872 303946 472894
rect 303998 472872 304010 472894
rect 304062 472872 304074 472894
rect 304126 472872 304138 472894
rect 303882 472870 304190 472872
rect 303882 472860 303888 472870
rect 303944 472860 303968 472870
rect 304024 472860 304048 472870
rect 304104 472860 304128 472870
rect 304184 472860 304190 472870
rect 303944 472814 303946 472860
rect 304126 472814 304128 472860
rect 303934 472808 303946 472814
rect 303998 472808 304010 472814
rect 304062 472808 304074 472814
rect 304126 472808 304138 472814
rect 303882 472802 304190 472808
rect 310944 472894 310946 472924
rect 311126 472894 311128 472924
rect 310934 472872 310946 472894
rect 310998 472872 311010 472894
rect 311062 472872 311074 472894
rect 311126 472872 311138 472894
rect 310882 472870 311190 472872
rect 310882 472860 310888 472870
rect 310944 472860 310968 472870
rect 311024 472860 311048 472870
rect 311104 472860 311128 472870
rect 311184 472860 311190 472870
rect 310944 472814 310946 472860
rect 311126 472814 311128 472860
rect 310934 472808 310946 472814
rect 310998 472808 311010 472814
rect 311062 472808 311074 472814
rect 311126 472808 311138 472814
rect 310882 472802 311190 472808
rect 301594 472696 301650 472705
rect 301594 472631 301650 472640
rect 309138 472696 309194 472705
rect 309138 472631 309194 472640
rect 312358 472696 312414 472705
rect 312358 472631 312414 472640
rect 294880 472592 294932 472598
rect 294880 472534 294932 472540
rect 295248 472592 295300 472598
rect 295248 472534 295300 472540
rect 295260 451178 295288 472534
rect 301608 472274 301636 472631
rect 305508 472560 305564 472569
rect 305508 472495 305564 472504
rect 301608 472246 301951 472274
rect 305522 472260 305550 472495
rect 309152 472325 309180 472631
rect 309140 472319 309192 472325
rect 309140 472261 309192 472267
rect 312372 472274 312400 472631
rect 312372 472246 312706 472274
rect 302150 472015 302458 472021
rect 302202 472009 302214 472015
rect 302266 472009 302278 472015
rect 302330 472009 302342 472015
rect 302394 472009 302406 472015
rect 302212 471963 302214 472009
rect 302394 471963 302396 472009
rect 302150 471953 302156 471963
rect 302212 471953 302236 471963
rect 302292 471953 302316 471963
rect 302372 471953 302396 471963
rect 302452 471953 302458 471963
rect 302150 471951 302458 471953
rect 302202 471929 302214 471951
rect 302266 471929 302278 471951
rect 302330 471929 302342 471951
rect 302394 471929 302406 471951
rect 302212 471899 302214 471929
rect 302394 471899 302396 471929
rect 302150 471887 302156 471899
rect 302212 471887 302236 471899
rect 302292 471887 302316 471899
rect 302372 471887 302396 471899
rect 302452 471887 302458 471899
rect 302212 471873 302214 471887
rect 302394 471873 302396 471887
rect 302202 471849 302214 471873
rect 302266 471849 302278 471873
rect 302330 471849 302342 471873
rect 302394 471849 302406 471873
rect 302212 471835 302214 471849
rect 302394 471835 302396 471849
rect 302150 471823 302156 471835
rect 302212 471823 302236 471835
rect 302292 471823 302316 471835
rect 302372 471823 302396 471835
rect 302452 471823 302458 471835
rect 302212 471793 302214 471823
rect 302394 471793 302396 471823
rect 302202 471771 302214 471793
rect 302266 471771 302278 471793
rect 302330 471771 302342 471793
rect 302394 471771 302406 471793
rect 302150 471769 302458 471771
rect 302150 471759 302156 471769
rect 302212 471759 302236 471769
rect 302292 471759 302316 471769
rect 302372 471759 302396 471769
rect 302452 471759 302458 471769
rect 302212 471713 302214 471759
rect 302394 471713 302396 471759
rect 302202 471707 302214 471713
rect 302266 471707 302278 471713
rect 302330 471707 302342 471713
rect 302394 471707 302406 471713
rect 302150 471701 302458 471707
rect 309150 472015 309458 472021
rect 309202 472009 309214 472015
rect 309266 472009 309278 472015
rect 309330 472009 309342 472015
rect 309394 472009 309406 472015
rect 309212 471963 309214 472009
rect 309394 471963 309396 472009
rect 309150 471953 309156 471963
rect 309212 471953 309236 471963
rect 309292 471953 309316 471963
rect 309372 471953 309396 471963
rect 309452 471953 309458 471963
rect 309150 471951 309458 471953
rect 309202 471929 309214 471951
rect 309266 471929 309278 471951
rect 309330 471929 309342 471951
rect 309394 471929 309406 471951
rect 309212 471899 309214 471929
rect 309394 471899 309396 471929
rect 309150 471887 309156 471899
rect 309212 471887 309236 471899
rect 309292 471887 309316 471899
rect 309372 471887 309396 471899
rect 309452 471887 309458 471899
rect 309212 471873 309214 471887
rect 309394 471873 309396 471887
rect 309202 471849 309214 471873
rect 309266 471849 309278 471873
rect 309330 471849 309342 471873
rect 309394 471849 309406 471873
rect 309212 471835 309214 471849
rect 309394 471835 309396 471849
rect 309150 471823 309156 471835
rect 309212 471823 309236 471835
rect 309292 471823 309316 471835
rect 309372 471823 309396 471835
rect 309452 471823 309458 471835
rect 309212 471793 309214 471823
rect 309394 471793 309396 471823
rect 309202 471771 309214 471793
rect 309266 471771 309278 471793
rect 309330 471771 309342 471793
rect 309394 471771 309406 471793
rect 309150 471769 309458 471771
rect 309150 471759 309156 471769
rect 309212 471759 309236 471769
rect 309292 471759 309316 471769
rect 309372 471759 309396 471769
rect 309452 471759 309458 471769
rect 309212 471713 309214 471759
rect 309394 471713 309396 471759
rect 309202 471707 309214 471713
rect 309266 471707 309278 471713
rect 309330 471707 309342 471713
rect 309394 471707 309406 471713
rect 309150 471701 309458 471707
rect 313660 471458 313688 474671
rect 318246 474056 318302 474065
rect 318246 473991 318302 474000
rect 313738 473512 313794 473521
rect 313738 473447 313794 473456
rect 313568 471430 313688 471458
rect 299296 471096 299348 471102
rect 299296 471038 299348 471044
rect 302884 471096 302936 471102
rect 302884 471038 302936 471044
rect 306472 471096 306524 471102
rect 306472 471038 306524 471044
rect 299308 468625 299336 471038
rect 299294 468616 299350 468625
rect 299294 468551 299350 468560
rect 302896 468489 302924 471038
rect 302882 468480 302938 468489
rect 302882 468415 302938 468424
rect 306484 467945 306512 471038
rect 310058 470656 310114 470665
rect 310058 470591 310114 470600
rect 313568 470594 313596 471430
rect 313752 471306 313780 473447
rect 313830 473376 313886 473385
rect 313830 473311 313886 473320
rect 313740 471300 313792 471306
rect 313740 471242 313792 471248
rect 313648 471096 313700 471102
rect 313646 471064 313648 471073
rect 313740 471096 313792 471102
rect 313700 471064 313702 471073
rect 313740 471038 313792 471044
rect 313646 470999 313702 471008
rect 310072 468761 310100 470591
rect 313568 470566 313688 470594
rect 310058 468752 310114 468761
rect 310058 468687 310114 468696
rect 306470 467936 306526 467945
rect 306470 467871 306526 467880
rect 313002 455424 313058 455433
rect 313002 455359 313058 455368
rect 312542 453928 312598 453937
rect 312542 453863 312598 453872
rect 312556 452713 312584 453863
rect 308310 452704 308366 452713
rect 308310 452639 308366 452648
rect 312542 452704 312598 452713
rect 312542 452639 312598 452648
rect 296882 452076 297190 452082
rect 296934 452054 296946 452076
rect 296998 452054 297010 452076
rect 297062 452054 297074 452076
rect 297126 452054 297138 452076
rect 296944 452024 296946 452054
rect 297126 452024 297128 452054
rect 296882 452012 296888 452024
rect 296944 452012 296968 452024
rect 297024 452012 297048 452024
rect 297104 452012 297128 452024
rect 297184 452012 297190 452024
rect 296944 451998 296946 452012
rect 297126 451998 297128 452012
rect 296934 451974 296946 451998
rect 296998 451974 297010 451998
rect 297062 451974 297074 451998
rect 297126 451974 297138 451998
rect 296944 451960 296946 451974
rect 297126 451960 297128 451974
rect 296882 451948 296888 451960
rect 296944 451948 296968 451960
rect 297024 451948 297048 451960
rect 297104 451948 297128 451960
rect 297184 451948 297190 451960
rect 296944 451918 296946 451948
rect 297126 451918 297128 451948
rect 296934 451896 296946 451918
rect 296998 451896 297010 451918
rect 297062 451896 297074 451918
rect 297126 451896 297138 451918
rect 296882 451894 297190 451896
rect 296882 451884 296888 451894
rect 296944 451884 296968 451894
rect 297024 451884 297048 451894
rect 297104 451884 297128 451894
rect 297184 451884 297190 451894
rect 296944 451838 296946 451884
rect 297126 451838 297128 451884
rect 296934 451832 296946 451838
rect 296998 451832 297010 451838
rect 297062 451832 297074 451838
rect 297126 451832 297138 451838
rect 296882 451820 297190 451832
rect 296934 451814 296946 451820
rect 296998 451814 297010 451820
rect 297062 451814 297074 451820
rect 297126 451814 297138 451820
rect 296944 451768 296946 451814
rect 297126 451768 297128 451814
rect 296882 451758 296888 451768
rect 296944 451758 296968 451768
rect 297024 451758 297048 451768
rect 297104 451758 297128 451768
rect 297184 451758 297190 451768
rect 296882 451756 297190 451758
rect 296934 451734 296946 451756
rect 296998 451734 297010 451756
rect 297062 451734 297074 451756
rect 297126 451734 297138 451756
rect 296944 451704 296946 451734
rect 297126 451704 297128 451734
rect 296882 451692 296888 451704
rect 296944 451692 296968 451704
rect 297024 451692 297048 451704
rect 297104 451692 297128 451704
rect 297184 451692 297190 451704
rect 296944 451678 296946 451692
rect 297126 451678 297128 451692
rect 296934 451654 296946 451678
rect 296998 451654 297010 451678
rect 297062 451654 297074 451678
rect 297126 451654 297138 451678
rect 296944 451640 296946 451654
rect 297126 451640 297128 451654
rect 296882 451628 296888 451640
rect 296944 451628 296968 451640
rect 297024 451628 297048 451640
rect 297104 451628 297128 451640
rect 297184 451628 297190 451640
rect 296944 451598 296946 451628
rect 297126 451598 297128 451628
rect 296934 451576 296946 451598
rect 296998 451576 297010 451598
rect 297062 451576 297074 451598
rect 297126 451576 297138 451598
rect 296882 451574 297190 451576
rect 296882 451564 296888 451574
rect 296944 451564 296968 451574
rect 297024 451564 297048 451574
rect 297104 451564 297128 451574
rect 297184 451564 297190 451574
rect 296944 451518 296946 451564
rect 297126 451518 297128 451564
rect 296934 451512 296946 451518
rect 296998 451512 297010 451518
rect 297062 451512 297074 451518
rect 297126 451512 297138 451518
rect 296882 451500 297190 451512
rect 296934 451494 296946 451500
rect 296998 451494 297010 451500
rect 297062 451494 297074 451500
rect 297126 451494 297138 451500
rect 296944 451448 296946 451494
rect 297126 451448 297128 451494
rect 296882 451438 296888 451448
rect 296944 451438 296968 451448
rect 297024 451438 297048 451448
rect 297104 451438 297128 451448
rect 297184 451438 297190 451448
rect 296882 451436 297190 451438
rect 296934 451414 296946 451436
rect 296998 451414 297010 451436
rect 297062 451414 297074 451436
rect 297126 451414 297138 451436
rect 296944 451384 296946 451414
rect 297126 451384 297128 451414
rect 296882 451372 296888 451384
rect 296944 451372 296968 451384
rect 297024 451372 297048 451384
rect 297104 451372 297128 451384
rect 297184 451372 297190 451384
rect 296944 451358 296946 451372
rect 297126 451358 297128 451372
rect 296934 451334 296946 451358
rect 296998 451334 297010 451358
rect 297062 451334 297074 451358
rect 297126 451334 297138 451358
rect 296944 451320 296946 451334
rect 297126 451320 297128 451334
rect 296882 451308 296888 451320
rect 296944 451308 296968 451320
rect 297024 451308 297048 451320
rect 297104 451308 297128 451320
rect 297184 451308 297190 451320
rect 296944 451278 296946 451308
rect 297126 451278 297128 451308
rect 296934 451256 296946 451278
rect 296998 451256 297010 451278
rect 297062 451256 297074 451278
rect 297126 451256 297138 451278
rect 296882 451250 297190 451256
rect 303882 452076 304190 452082
rect 303934 452054 303946 452076
rect 303998 452054 304010 452076
rect 304062 452054 304074 452076
rect 304126 452054 304138 452076
rect 303944 452024 303946 452054
rect 304126 452024 304128 452054
rect 303882 452012 303888 452024
rect 303944 452012 303968 452024
rect 304024 452012 304048 452024
rect 304104 452012 304128 452024
rect 304184 452012 304190 452024
rect 303944 451998 303946 452012
rect 304126 451998 304128 452012
rect 303934 451974 303946 451998
rect 303998 451974 304010 451998
rect 304062 451974 304074 451998
rect 304126 451974 304138 451998
rect 303944 451960 303946 451974
rect 304126 451960 304128 451974
rect 303882 451948 303888 451960
rect 303944 451948 303968 451960
rect 304024 451948 304048 451960
rect 304104 451948 304128 451960
rect 304184 451948 304190 451960
rect 303944 451918 303946 451948
rect 304126 451918 304128 451948
rect 303934 451896 303946 451918
rect 303998 451896 304010 451918
rect 304062 451896 304074 451918
rect 304126 451896 304138 451918
rect 303882 451894 304190 451896
rect 303882 451884 303888 451894
rect 303944 451884 303968 451894
rect 304024 451884 304048 451894
rect 304104 451884 304128 451894
rect 304184 451884 304190 451894
rect 303944 451838 303946 451884
rect 304126 451838 304128 451884
rect 303934 451832 303946 451838
rect 303998 451832 304010 451838
rect 304062 451832 304074 451838
rect 304126 451832 304138 451838
rect 303882 451820 304190 451832
rect 303934 451814 303946 451820
rect 303998 451814 304010 451820
rect 304062 451814 304074 451820
rect 304126 451814 304138 451820
rect 303944 451768 303946 451814
rect 304126 451768 304128 451814
rect 303882 451758 303888 451768
rect 303944 451758 303968 451768
rect 304024 451758 304048 451768
rect 304104 451758 304128 451768
rect 304184 451758 304190 451768
rect 308324 451761 308352 452639
rect 310897 452076 311077 452082
rect 310949 452054 310961 452076
rect 311013 452054 311025 452076
rect 310897 452012 310919 452024
rect 310975 452012 310999 452024
rect 311055 452012 311077 452024
rect 310949 451974 310961 451998
rect 311013 451974 311025 451998
rect 310897 451948 310919 451960
rect 310975 451948 310999 451960
rect 311055 451948 311077 451960
rect 310949 451896 310961 451918
rect 311013 451896 311025 451918
rect 310897 451894 311077 451896
rect 310897 451884 310919 451894
rect 310975 451884 310999 451894
rect 311055 451884 311077 451894
rect 310949 451832 310961 451838
rect 311013 451832 311025 451838
rect 310897 451820 311077 451832
rect 310949 451814 310961 451820
rect 311013 451814 311025 451820
rect 303882 451756 304190 451758
rect 303934 451734 303946 451756
rect 303998 451734 304010 451756
rect 304062 451734 304074 451756
rect 304126 451734 304138 451756
rect 303944 451704 303946 451734
rect 304126 451704 304128 451734
rect 303882 451692 303888 451704
rect 303944 451692 303968 451704
rect 304024 451692 304048 451704
rect 304104 451692 304128 451704
rect 304184 451692 304190 451704
rect 303944 451678 303946 451692
rect 304126 451678 304128 451692
rect 308310 451752 308366 451761
rect 308310 451687 308366 451696
rect 310897 451758 310919 451768
rect 310975 451758 310999 451768
rect 311055 451758 311077 451768
rect 310897 451756 311077 451758
rect 310949 451734 310961 451756
rect 311013 451734 311025 451756
rect 310897 451692 310919 451704
rect 310975 451692 310999 451704
rect 311055 451692 311077 451704
rect 303934 451654 303946 451678
rect 303998 451654 304010 451678
rect 304062 451654 304074 451678
rect 304126 451654 304138 451678
rect 303944 451640 303946 451654
rect 304126 451640 304128 451654
rect 303882 451628 303888 451640
rect 303944 451628 303968 451640
rect 304024 451628 304048 451640
rect 304104 451628 304128 451640
rect 304184 451628 304190 451640
rect 303944 451598 303946 451628
rect 304126 451598 304128 451628
rect 303934 451576 303946 451598
rect 303998 451576 304010 451598
rect 304062 451576 304074 451598
rect 304126 451576 304138 451598
rect 303882 451574 304190 451576
rect 303882 451564 303888 451574
rect 303944 451564 303968 451574
rect 304024 451564 304048 451574
rect 304104 451564 304128 451574
rect 304184 451564 304190 451574
rect 303944 451518 303946 451564
rect 304126 451518 304128 451564
rect 303934 451512 303946 451518
rect 303998 451512 304010 451518
rect 304062 451512 304074 451518
rect 304126 451512 304138 451518
rect 303882 451500 304190 451512
rect 303934 451494 303946 451500
rect 303998 451494 304010 451500
rect 304062 451494 304074 451500
rect 304126 451494 304138 451500
rect 303944 451448 303946 451494
rect 304126 451448 304128 451494
rect 310949 451654 310961 451678
rect 311013 451654 311025 451678
rect 310897 451628 310919 451640
rect 310975 451628 310999 451640
rect 311055 451628 311077 451640
rect 310949 451576 310961 451598
rect 311013 451576 311025 451598
rect 310897 451574 311077 451576
rect 310897 451564 310919 451574
rect 310975 451564 310999 451574
rect 311055 451564 311077 451574
rect 310949 451512 310961 451518
rect 311013 451512 311025 451518
rect 310897 451500 311077 451512
rect 310949 451494 310961 451500
rect 311013 451494 311025 451500
rect 303882 451438 303888 451448
rect 303944 451438 303968 451448
rect 304024 451438 304048 451448
rect 304104 451438 304128 451448
rect 304184 451438 304190 451448
rect 303882 451436 304190 451438
rect 303934 451414 303946 451436
rect 303998 451414 304010 451436
rect 304062 451414 304074 451436
rect 304126 451414 304138 451436
rect 308015 451424 308024 451480
rect 308080 451424 308089 451480
rect 310897 451438 310919 451448
rect 310975 451438 310999 451448
rect 311055 451438 311077 451448
rect 310897 451436 311077 451438
rect 303944 451384 303946 451414
rect 304126 451384 304128 451414
rect 303882 451372 303888 451384
rect 303944 451372 303968 451384
rect 304024 451372 304048 451384
rect 304104 451372 304128 451384
rect 304184 451372 304190 451384
rect 303944 451358 303946 451372
rect 304126 451358 304128 451372
rect 303934 451334 303946 451358
rect 303998 451334 304010 451358
rect 304062 451334 304074 451358
rect 304126 451334 304138 451358
rect 303944 451320 303946 451334
rect 304126 451320 304128 451334
rect 303882 451308 303888 451320
rect 303944 451308 303968 451320
rect 304024 451308 304048 451320
rect 304104 451308 304128 451320
rect 304184 451308 304190 451320
rect 303944 451278 303946 451308
rect 304126 451278 304128 451308
rect 303934 451256 303946 451278
rect 303998 451256 304010 451278
rect 304062 451256 304074 451278
rect 304126 451256 304138 451278
rect 303882 451250 304190 451256
rect 310949 451414 310961 451436
rect 311013 451414 311025 451436
rect 310897 451372 310919 451384
rect 310975 451372 310999 451384
rect 311055 451372 311077 451384
rect 310949 451334 310961 451358
rect 311013 451334 311025 451358
rect 310897 451308 310919 451320
rect 310975 451308 310999 451320
rect 311055 451308 311077 451320
rect 310949 451256 310961 451278
rect 311013 451256 311025 451278
rect 310897 451250 311077 451256
rect 295248 451172 295300 451178
rect 295248 451114 295300 451120
rect 293866 449168 293922 449177
rect 293866 449103 293922 449112
rect 292488 430296 292540 430302
rect 292488 430238 292540 430244
rect 295260 430250 295288 451114
rect 298940 448089 298968 450636
rect 300860 450424 300912 450430
rect 300860 450366 300912 450372
rect 300872 449177 300900 450366
rect 300858 449168 300914 449177
rect 300858 449103 300914 449112
rect 298926 448080 298982 448089
rect 298926 448015 298982 448024
rect 300872 430817 300900 449103
rect 302252 448225 302280 450636
rect 302238 448216 302294 448225
rect 302238 448151 302294 448160
rect 305564 447953 305592 450636
rect 306196 450492 306248 450498
rect 306196 450434 306248 450440
rect 306208 449177 306236 450434
rect 306194 449168 306250 449177
rect 306194 449103 306250 449112
rect 305550 447944 305606 447953
rect 305550 447879 305606 447888
rect 306208 447134 306236 449103
rect 308876 447817 308904 450636
rect 312165 450608 312174 450664
rect 312230 450608 312239 450664
rect 310884 450191 311128 450197
rect 310936 450177 310948 450191
rect 311000 450177 311012 450191
rect 311064 450177 311076 450191
rect 310884 450127 310898 450139
rect 310954 450127 310978 450139
rect 311034 450127 311058 450139
rect 311114 450127 311128 450139
rect 310936 450097 310948 450121
rect 311000 450097 311012 450121
rect 311064 450097 311076 450121
rect 310884 450063 310898 450075
rect 310954 450063 310978 450075
rect 311034 450063 311058 450075
rect 311114 450063 311128 450075
rect 310936 450017 310948 450041
rect 311000 450017 311012 450041
rect 311064 450017 311076 450041
rect 310884 449999 310898 450011
rect 310954 449999 310978 450011
rect 311034 449999 311058 450011
rect 311114 449999 311128 450011
rect 310936 449947 310948 449961
rect 311000 449947 311012 449961
rect 311064 449947 311076 449961
rect 310884 449937 311128 449947
rect 310884 449935 310898 449937
rect 310954 449935 310978 449937
rect 311034 449935 311058 449937
rect 311114 449935 311128 449937
rect 310884 449881 310898 449883
rect 310954 449881 310978 449883
rect 311034 449881 311058 449883
rect 311114 449881 311128 449883
rect 310884 449871 311128 449881
rect 310936 449857 310948 449871
rect 311000 449857 311012 449871
rect 311064 449857 311076 449871
rect 310884 449807 310898 449819
rect 310954 449807 310978 449819
rect 311034 449807 311058 449819
rect 311114 449807 311128 449819
rect 310936 449777 310948 449801
rect 311000 449777 311012 449801
rect 311064 449777 311076 449801
rect 310884 449743 310898 449755
rect 310954 449743 310978 449755
rect 311034 449743 311058 449755
rect 311114 449743 311128 449755
rect 310936 449697 310948 449721
rect 311000 449697 311012 449721
rect 311064 449697 311076 449721
rect 310884 449679 310898 449691
rect 310954 449679 310978 449691
rect 311034 449679 311058 449691
rect 311114 449679 311128 449691
rect 310936 449627 310948 449641
rect 311000 449627 311012 449641
rect 311064 449627 311076 449641
rect 310884 449621 311128 449627
rect 308862 447808 308918 447817
rect 308862 447743 308918 447752
rect 306208 447106 306328 447134
rect 306300 432177 306328 447106
rect 312556 433265 312584 452639
rect 313016 450566 313044 455359
rect 313660 451274 313688 470566
rect 313752 453937 313780 471038
rect 313844 455433 313872 473311
rect 318062 471064 318118 471073
rect 318062 470999 318118 471008
rect 313922 467936 313978 467945
rect 313922 467871 313978 467880
rect 313830 455424 313886 455433
rect 313830 455359 313886 455368
rect 313738 453928 313794 453937
rect 313738 453863 313794 453872
rect 313476 451246 313688 451274
rect 313004 450560 313056 450566
rect 313004 450502 313056 450508
rect 312634 448080 312690 448089
rect 312634 448015 312690 448024
rect 308494 433256 308550 433265
rect 308494 433191 308550 433200
rect 312542 433256 312598 433265
rect 312542 433191 312598 433200
rect 305182 432168 305238 432177
rect 305182 432103 305238 432112
rect 306286 432168 306342 432177
rect 306286 432103 306342 432112
rect 305196 430817 305224 432103
rect 308508 430817 308536 433191
rect 312648 431225 312676 448015
rect 312634 431216 312690 431225
rect 312634 431151 312690 431160
rect 300858 430808 300914 430817
rect 300858 430743 300914 430752
rect 305182 430808 305238 430817
rect 305182 430743 305238 430752
rect 308494 430808 308550 430817
rect 308494 430743 308550 430752
rect 301502 430400 301558 430409
rect 301502 430335 301558 430344
rect 305091 430400 305147 430409
rect 305091 430335 305147 430344
rect 308402 430400 308458 430409
rect 313016 430386 313044 450502
rect 313476 449177 313504 451246
rect 313462 449168 313518 449177
rect 313462 449103 313518 449112
rect 313370 433256 313426 433265
rect 313370 433191 313426 433200
rect 313278 432168 313334 432177
rect 313278 432103 313334 432112
rect 308458 430358 308562 430386
rect 312832 430358 313044 430386
rect 308402 430335 308458 430344
rect 295892 430289 295944 430295
rect 292500 409290 292528 430238
rect 295260 430237 295892 430250
rect 295260 430231 295944 430237
rect 295260 430222 295932 430231
rect 295154 410272 295210 410281
rect 295154 410207 295210 410216
rect 292488 409284 292540 409290
rect 292488 409226 292540 409232
rect 292500 388482 292528 409226
rect 295168 402974 295196 410207
rect 295260 409562 295288 430222
rect 301516 430114 301544 430335
rect 312832 430302 312860 430358
rect 312452 430296 312504 430302
rect 312452 430238 312504 430244
rect 312820 430296 312872 430302
rect 312820 430238 312872 430244
rect 301516 430100 301674 430114
rect 301516 430086 301688 430100
rect 301660 429461 301688 430086
rect 309151 430000 309447 430006
rect 309151 429994 309177 430000
rect 309229 429994 309241 430000
rect 309229 429948 309231 429994
rect 309293 429948 309305 430000
rect 309357 429994 309369 430000
rect 309421 429994 309447 430000
rect 309367 429948 309369 429994
rect 309207 429938 309231 429948
rect 309287 429938 309311 429948
rect 309367 429938 309391 429948
rect 309151 429936 309447 429938
rect 309151 429914 309177 429936
rect 309229 429914 309241 429936
rect 309229 429884 309231 429914
rect 309293 429884 309305 429936
rect 309357 429914 309369 429936
rect 309421 429914 309447 429936
rect 309367 429884 309369 429914
rect 309207 429872 309231 429884
rect 309287 429872 309311 429884
rect 309367 429872 309391 429884
rect 309229 429858 309231 429872
rect 309151 429834 309177 429858
rect 309229 429834 309241 429858
rect 309229 429820 309231 429834
rect 309293 429820 309305 429872
rect 309367 429858 309369 429872
rect 309357 429834 309369 429858
rect 309421 429834 309447 429858
rect 309367 429820 309369 429834
rect 309207 429808 309231 429820
rect 309287 429808 309311 429820
rect 309367 429808 309391 429820
rect 309229 429778 309231 429808
rect 309151 429756 309177 429778
rect 309229 429756 309241 429778
rect 309293 429756 309305 429808
rect 309367 429778 309369 429808
rect 309357 429756 309369 429778
rect 309421 429756 309447 429778
rect 309151 429754 309447 429756
rect 309207 429744 309231 429754
rect 309287 429744 309311 429754
rect 309367 429744 309391 429754
rect 309229 429698 309231 429744
rect 309151 429692 309177 429698
rect 309229 429692 309241 429698
rect 309293 429692 309305 429744
rect 309367 429698 309369 429744
rect 309357 429692 309369 429698
rect 309421 429692 309447 429698
rect 309151 429686 309447 429692
rect 301660 429455 301740 429461
rect 301660 429406 301688 429455
rect 301688 429397 301740 429403
rect 301688 429208 301740 429214
rect 301688 429150 301740 429156
rect 299020 429084 299072 429090
rect 299020 429026 299072 429032
rect 299032 417081 299060 429026
rect 301700 427961 301728 429150
rect 305920 429072 305972 429078
rect 305920 429014 305972 429020
rect 302516 429004 302568 429010
rect 302516 428946 302568 428952
rect 300858 427952 300914 427961
rect 300858 427887 300914 427896
rect 301686 427952 301742 427961
rect 301686 427887 301742 427896
rect 300872 422294 300900 427887
rect 302528 427417 302556 428946
rect 302514 427408 302570 427417
rect 302514 427343 302570 427352
rect 305932 427281 305960 429014
rect 309414 428496 309470 428505
rect 309414 428431 309470 428440
rect 305918 427272 305974 427281
rect 305918 427207 305974 427216
rect 309428 427145 309456 428431
rect 309414 427136 309470 427145
rect 309414 427071 309470 427080
rect 309046 423600 309102 423609
rect 309046 423535 309102 423544
rect 300872 422266 301084 422294
rect 299018 417072 299074 417081
rect 299018 417007 299074 417016
rect 301056 410281 301084 422266
rect 305182 411360 305238 411369
rect 305182 411295 305238 411304
rect 301042 410272 301098 410281
rect 301042 410207 301098 410216
rect 296882 410086 297190 410092
rect 296934 410080 296946 410086
rect 296998 410080 297010 410086
rect 297062 410080 297074 410086
rect 297126 410080 297138 410086
rect 296944 410034 296946 410080
rect 297126 410034 297128 410080
rect 296882 410024 296888 410034
rect 296944 410024 296968 410034
rect 297024 410024 297048 410034
rect 297104 410024 297128 410034
rect 297184 410024 297190 410034
rect 296882 410022 297190 410024
rect 296934 410000 296946 410022
rect 296998 410000 297010 410022
rect 297062 410000 297074 410022
rect 297126 410000 297138 410022
rect 296944 409970 296946 410000
rect 297126 409970 297128 410000
rect 296882 409958 296888 409970
rect 296944 409958 296968 409970
rect 297024 409958 297048 409970
rect 297104 409958 297128 409970
rect 297184 409958 297190 409970
rect 296944 409944 296946 409958
rect 297126 409944 297128 409958
rect 296934 409920 296946 409944
rect 296998 409920 297010 409944
rect 297062 409920 297074 409944
rect 297126 409920 297138 409944
rect 296944 409906 296946 409920
rect 297126 409906 297128 409920
rect 296882 409894 296888 409906
rect 296944 409894 296968 409906
rect 297024 409894 297048 409906
rect 297104 409894 297128 409906
rect 297184 409894 297190 409906
rect 296944 409864 296946 409894
rect 297126 409864 297128 409894
rect 301056 409873 301084 410207
rect 303882 410086 304190 410092
rect 303934 410080 303946 410086
rect 303998 410080 304010 410086
rect 304062 410080 304074 410086
rect 304126 410080 304138 410086
rect 303944 410034 303946 410080
rect 304126 410034 304128 410080
rect 303882 410024 303888 410034
rect 303944 410024 303968 410034
rect 304024 410024 304048 410034
rect 304104 410024 304128 410034
rect 304184 410024 304190 410034
rect 303882 410022 304190 410024
rect 303934 410000 303946 410022
rect 303998 410000 304010 410022
rect 304062 410000 304074 410022
rect 304126 410000 304138 410022
rect 303944 409970 303946 410000
rect 304126 409970 304128 410000
rect 303882 409958 303888 409970
rect 303944 409958 303968 409970
rect 304024 409958 304048 409970
rect 304104 409958 304128 409970
rect 304184 409958 304190 409970
rect 303944 409944 303946 409958
rect 304126 409944 304128 409958
rect 303934 409920 303946 409944
rect 303998 409920 304010 409944
rect 304062 409920 304074 409944
rect 304126 409920 304138 409944
rect 303944 409906 303946 409920
rect 304126 409906 304128 409920
rect 303882 409894 303888 409906
rect 303944 409894 303968 409906
rect 304024 409894 304048 409906
rect 304104 409894 304128 409906
rect 304184 409894 304190 409906
rect 296934 409842 296946 409864
rect 296998 409842 297010 409864
rect 297062 409842 297074 409864
rect 297126 409842 297138 409864
rect 296882 409840 297190 409842
rect 296882 409830 296888 409840
rect 296944 409830 296968 409840
rect 297024 409830 297048 409840
rect 297104 409830 297128 409840
rect 297184 409830 297190 409840
rect 296944 409784 296946 409830
rect 297126 409784 297128 409830
rect 301042 409864 301098 409873
rect 301042 409799 301098 409808
rect 303944 409864 303946 409894
rect 304126 409864 304128 409894
rect 305196 409873 305224 411295
rect 309060 410281 309088 423535
rect 312464 411505 312492 430238
rect 313004 429084 313056 429090
rect 313002 429040 313004 429049
rect 313056 429040 313058 429049
rect 313002 428975 313058 428984
rect 313292 412634 313320 432103
rect 313384 423609 313412 433191
rect 313370 423600 313426 423609
rect 313370 423535 313426 423544
rect 313200 412606 313320 412634
rect 312450 411496 312506 411505
rect 312450 411431 312506 411440
rect 313200 411369 313228 412606
rect 313278 411496 313334 411505
rect 313278 411431 313334 411440
rect 312266 411360 312322 411369
rect 312266 411295 312322 411304
rect 313186 411360 313242 411369
rect 313186 411295 313242 411304
rect 309046 410272 309102 410281
rect 309046 410207 309102 410216
rect 312082 410272 312138 410281
rect 312082 410207 312138 410216
rect 310882 410086 311190 410092
rect 310934 410080 310946 410086
rect 310998 410080 311010 410086
rect 311062 410080 311074 410086
rect 311126 410080 311138 410086
rect 310944 410034 310946 410080
rect 311126 410034 311128 410080
rect 310882 410024 310888 410034
rect 310944 410024 310968 410034
rect 311024 410024 311048 410034
rect 311104 410024 311128 410034
rect 311184 410024 311190 410034
rect 310882 410022 311190 410024
rect 310934 410000 310946 410022
rect 310998 410000 311010 410022
rect 311062 410000 311074 410022
rect 311126 410000 311138 410022
rect 310944 409970 310946 410000
rect 311126 409970 311128 410000
rect 310882 409958 310888 409970
rect 310944 409958 310968 409970
rect 311024 409958 311048 409970
rect 311104 409958 311128 409970
rect 311184 409958 311190 409970
rect 310944 409944 310946 409958
rect 311126 409944 311128 409958
rect 310934 409920 310946 409944
rect 310998 409920 311010 409944
rect 311062 409920 311074 409944
rect 311126 409920 311138 409944
rect 310944 409906 310946 409920
rect 311126 409906 311128 409920
rect 310882 409894 310888 409906
rect 310944 409894 310968 409906
rect 311024 409894 311048 409906
rect 311104 409894 311128 409906
rect 311184 409894 311190 409906
rect 303934 409842 303946 409864
rect 303998 409842 304010 409864
rect 304062 409842 304074 409864
rect 304126 409842 304138 409864
rect 303882 409840 304190 409842
rect 303882 409830 303888 409840
rect 303944 409830 303968 409840
rect 304024 409830 304048 409840
rect 304104 409830 304128 409840
rect 304184 409830 304190 409840
rect 296934 409778 296946 409784
rect 296998 409778 297010 409784
rect 297062 409778 297074 409784
rect 297126 409778 297138 409784
rect 296882 409772 297190 409778
rect 303944 409784 303946 409830
rect 304126 409784 304128 409830
rect 305182 409864 305238 409873
rect 305182 409799 305238 409808
rect 310944 409864 310946 409894
rect 311126 409864 311128 409894
rect 310934 409842 310946 409864
rect 310998 409842 311010 409864
rect 311062 409842 311074 409864
rect 311126 409842 311138 409864
rect 310882 409840 311190 409842
rect 310882 409830 310888 409840
rect 310944 409830 310968 409840
rect 311024 409830 311048 409840
rect 311104 409830 311128 409840
rect 311184 409830 311190 409840
rect 303934 409778 303946 409784
rect 303998 409778 304010 409784
rect 304062 409778 304074 409784
rect 304126 409778 304138 409784
rect 303882 409772 304190 409778
rect 310944 409784 310946 409830
rect 311126 409784 311128 409830
rect 310934 409778 310946 409784
rect 310998 409778 311010 409784
rect 311062 409778 311074 409784
rect 311126 409778 311138 409784
rect 310882 409772 311190 409778
rect 301226 409592 301282 409601
rect 295248 409556 295300 409562
rect 301226 409527 301282 409536
rect 304549 409592 304605 409601
rect 304549 409527 304605 409536
rect 307814 409592 307870 409601
rect 307814 409527 307870 409536
rect 295248 409498 295300 409504
rect 294984 402946 295196 402974
rect 294984 390697 295012 402946
rect 295260 393314 295288 409498
rect 301240 409306 301268 409527
rect 301240 409278 301312 409306
rect 304563 409292 304591 409527
rect 307828 409292 307856 409527
rect 302150 409000 302458 409006
rect 302202 408994 302214 409000
rect 302266 408994 302278 409000
rect 302330 408994 302342 409000
rect 302394 408994 302406 409000
rect 302212 408948 302214 408994
rect 302394 408948 302396 408994
rect 302150 408938 302156 408948
rect 302212 408938 302236 408948
rect 302292 408938 302316 408948
rect 302372 408938 302396 408948
rect 302452 408938 302458 408948
rect 302150 408936 302458 408938
rect 302202 408914 302214 408936
rect 302266 408914 302278 408936
rect 302330 408914 302342 408936
rect 302394 408914 302406 408936
rect 302212 408884 302214 408914
rect 302394 408884 302396 408914
rect 302150 408872 302156 408884
rect 302212 408872 302236 408884
rect 302292 408872 302316 408884
rect 302372 408872 302396 408884
rect 302452 408872 302458 408884
rect 302212 408858 302214 408872
rect 302394 408858 302396 408872
rect 302202 408834 302214 408858
rect 302266 408834 302278 408858
rect 302330 408834 302342 408858
rect 302394 408834 302406 408858
rect 302212 408820 302214 408834
rect 302394 408820 302396 408834
rect 302150 408808 302156 408820
rect 302212 408808 302236 408820
rect 302292 408808 302316 408820
rect 302372 408808 302396 408820
rect 302452 408808 302458 408820
rect 302212 408778 302214 408808
rect 302394 408778 302396 408808
rect 302202 408756 302214 408778
rect 302266 408756 302278 408778
rect 302330 408756 302342 408778
rect 302394 408756 302406 408778
rect 302150 408754 302458 408756
rect 302150 408744 302156 408754
rect 302212 408744 302236 408754
rect 302292 408744 302316 408754
rect 302372 408744 302396 408754
rect 302452 408744 302458 408754
rect 302212 408698 302214 408744
rect 302394 408698 302396 408744
rect 302202 408692 302214 408698
rect 302266 408692 302278 408698
rect 302330 408692 302342 408698
rect 302394 408692 302406 408698
rect 302150 408686 302458 408692
rect 298848 407017 298876 408612
rect 301976 408598 302174 408626
rect 305394 408598 305592 408626
rect 298834 407008 298890 407017
rect 298834 406943 298890 406952
rect 295076 393286 295288 393314
rect 294970 390688 295026 390697
rect 294970 390623 295026 390632
rect 292488 388476 292540 388482
rect 292488 388418 292540 388424
rect 292500 367470 292528 388418
rect 294984 370802 295012 390623
rect 295076 388550 295104 393286
rect 301594 390688 301650 390697
rect 301594 390623 301650 390632
rect 296882 389087 297190 389093
rect 296934 389081 296946 389087
rect 296998 389081 297010 389087
rect 297062 389081 297074 389087
rect 297126 389081 297138 389087
rect 296944 389035 296946 389081
rect 297126 389035 297128 389081
rect 296882 389025 296888 389035
rect 296944 389025 296968 389035
rect 297024 389025 297048 389035
rect 297104 389025 297128 389035
rect 297184 389025 297190 389035
rect 296882 389023 297190 389025
rect 296934 389001 296946 389023
rect 296998 389001 297010 389023
rect 297062 389001 297074 389023
rect 297126 389001 297138 389023
rect 296944 388971 296946 389001
rect 297126 388971 297128 389001
rect 296882 388959 296888 388971
rect 296944 388959 296968 388971
rect 297024 388959 297048 388971
rect 297104 388959 297128 388971
rect 297184 388959 297190 388971
rect 296944 388945 296946 388959
rect 297126 388945 297128 388959
rect 296934 388921 296946 388945
rect 296998 388921 297010 388945
rect 297062 388921 297074 388945
rect 297126 388921 297138 388945
rect 301608 388929 301636 390623
rect 301976 389881 302004 408598
rect 305564 391241 305592 408598
rect 308692 406337 308720 408612
rect 310882 407914 311190 407920
rect 310934 407908 310946 407914
rect 310998 407908 311010 407914
rect 311062 407908 311074 407914
rect 311126 407908 311138 407914
rect 310944 407862 310946 407908
rect 311126 407862 311128 407908
rect 310882 407852 310888 407862
rect 310944 407852 310968 407862
rect 311024 407852 311048 407862
rect 311104 407852 311128 407862
rect 311184 407852 311190 407862
rect 310882 407850 311190 407852
rect 310934 407828 310946 407850
rect 310998 407828 311010 407850
rect 311062 407828 311074 407850
rect 311126 407828 311138 407850
rect 310944 407798 310946 407828
rect 311126 407798 311128 407828
rect 310882 407786 310888 407798
rect 310944 407786 310968 407798
rect 311024 407786 311048 407798
rect 311104 407786 311128 407798
rect 311184 407786 311190 407798
rect 310944 407772 310946 407786
rect 311126 407772 311128 407786
rect 310934 407748 310946 407772
rect 310998 407748 311010 407772
rect 311062 407748 311074 407772
rect 311126 407748 311138 407772
rect 310944 407734 310946 407748
rect 311126 407734 311128 407748
rect 310882 407722 310888 407734
rect 310944 407722 310968 407734
rect 311024 407722 311048 407734
rect 311104 407722 311128 407734
rect 311184 407722 311190 407734
rect 310944 407692 310946 407722
rect 311126 407692 311128 407722
rect 310934 407670 310946 407692
rect 310998 407670 311010 407692
rect 311062 407670 311074 407692
rect 311126 407670 311138 407692
rect 310882 407668 311190 407670
rect 310882 407658 310888 407668
rect 310944 407658 310968 407668
rect 311024 407658 311048 407668
rect 311104 407658 311128 407668
rect 311184 407658 311190 407668
rect 310944 407612 310946 407658
rect 311126 407612 311128 407658
rect 310934 407606 310946 407612
rect 310998 407606 311010 407612
rect 311062 407606 311074 407612
rect 311126 407606 311138 407612
rect 310882 407600 311190 407606
rect 308678 406328 308734 406337
rect 308678 406263 308734 406272
rect 305918 391504 305974 391513
rect 305918 391439 305974 391448
rect 305550 391232 305606 391241
rect 305550 391167 305606 391176
rect 301962 389872 302018 389881
rect 301962 389807 302018 389816
rect 303882 389087 304190 389093
rect 303934 389081 303946 389087
rect 303998 389081 304010 389087
rect 304062 389081 304074 389087
rect 304126 389081 304138 389087
rect 303944 389035 303946 389081
rect 304126 389035 304128 389081
rect 303882 389025 303888 389035
rect 303944 389025 303968 389035
rect 304024 389025 304048 389035
rect 304104 389025 304128 389035
rect 304184 389025 304190 389035
rect 303882 389023 304190 389025
rect 303934 389001 303946 389023
rect 303998 389001 304010 389023
rect 304062 389001 304074 389023
rect 304126 389001 304138 389023
rect 303944 388971 303946 389001
rect 304126 388971 304128 389001
rect 303882 388959 303888 388971
rect 303944 388959 303968 388971
rect 304024 388959 304048 388971
rect 304104 388959 304128 388971
rect 304184 388959 304190 388971
rect 303944 388945 303946 388959
rect 304126 388945 304128 388959
rect 296944 388907 296946 388921
rect 297126 388907 297128 388921
rect 296882 388895 296888 388907
rect 296944 388895 296968 388907
rect 297024 388895 297048 388907
rect 297104 388895 297128 388907
rect 297184 388895 297190 388907
rect 296944 388865 296946 388895
rect 297126 388865 297128 388895
rect 296934 388843 296946 388865
rect 296998 388843 297010 388865
rect 297062 388843 297074 388865
rect 297126 388843 297138 388865
rect 301594 388920 301650 388929
rect 301594 388855 301650 388864
rect 303934 388921 303946 388945
rect 303998 388921 304010 388945
rect 304062 388921 304074 388945
rect 304126 388921 304138 388945
rect 305932 388929 305960 391439
rect 312096 390697 312124 410207
rect 312176 408060 312228 408066
rect 312176 408002 312228 408008
rect 312188 407969 312216 408002
rect 312174 407960 312230 407969
rect 312174 407895 312230 407904
rect 312280 391513 312308 411295
rect 313292 408474 313320 411431
rect 313280 408468 313332 408474
rect 313280 408410 313332 408416
rect 312266 391504 312322 391513
rect 312266 391439 312322 391448
rect 312280 390697 312308 391439
rect 309506 390688 309562 390697
rect 309506 390623 309562 390632
rect 312082 390688 312138 390697
rect 312082 390623 312138 390632
rect 312266 390688 312322 390697
rect 312266 390623 312322 390632
rect 309520 388929 309548 390623
rect 313936 390017 313964 467871
rect 315302 450664 315358 450673
rect 315302 450599 315358 450608
rect 314290 448216 314346 448225
rect 314290 448151 314346 448160
rect 313922 390008 313978 390017
rect 313922 389943 313978 389952
rect 310882 389087 311190 389093
rect 310934 389081 310946 389087
rect 310998 389081 311010 389087
rect 311062 389081 311074 389087
rect 311126 389081 311138 389087
rect 310944 389035 310946 389081
rect 311126 389035 311128 389081
rect 310882 389025 310888 389035
rect 310944 389025 310968 389035
rect 311024 389025 311048 389035
rect 311104 389025 311128 389035
rect 311184 389025 311190 389035
rect 310882 389023 311190 389025
rect 310934 389001 310946 389023
rect 310998 389001 311010 389023
rect 311062 389001 311074 389023
rect 311126 389001 311138 389023
rect 310944 388971 310946 389001
rect 311126 388971 311128 389001
rect 310882 388959 310888 388971
rect 310944 388959 310968 388971
rect 311024 388959 311048 388971
rect 311104 388959 311128 388971
rect 311184 388959 311190 388971
rect 310944 388945 310946 388959
rect 311126 388945 311128 388959
rect 303944 388907 303946 388921
rect 304126 388907 304128 388921
rect 303882 388895 303888 388907
rect 303944 388895 303968 388907
rect 304024 388895 304048 388907
rect 304104 388895 304128 388907
rect 304184 388895 304190 388907
rect 303944 388865 303946 388895
rect 304126 388865 304128 388895
rect 296882 388841 297190 388843
rect 296882 388831 296888 388841
rect 296944 388831 296968 388841
rect 297024 388831 297048 388841
rect 297104 388831 297128 388841
rect 297184 388831 297190 388841
rect 296944 388785 296946 388831
rect 297126 388785 297128 388831
rect 296934 388779 296946 388785
rect 296998 388779 297010 388785
rect 297062 388779 297074 388785
rect 297126 388779 297138 388785
rect 296882 388773 297190 388779
rect 303934 388843 303946 388865
rect 303998 388843 304010 388865
rect 304062 388843 304074 388865
rect 304126 388843 304138 388865
rect 305918 388920 305974 388929
rect 305918 388855 305974 388864
rect 309506 388920 309562 388929
rect 309506 388855 309562 388864
rect 310934 388921 310946 388945
rect 310998 388921 311010 388945
rect 311062 388921 311074 388945
rect 311126 388921 311138 388945
rect 310944 388907 310946 388921
rect 311126 388907 311128 388921
rect 310882 388895 310888 388907
rect 310944 388895 310968 388907
rect 311024 388895 311048 388907
rect 311104 388895 311128 388907
rect 311184 388895 311190 388907
rect 310944 388865 310946 388895
rect 311126 388865 311128 388895
rect 303882 388841 304190 388843
rect 303882 388831 303888 388841
rect 303944 388831 303968 388841
rect 304024 388831 304048 388841
rect 304104 388831 304128 388841
rect 304184 388831 304190 388841
rect 303944 388785 303946 388831
rect 304126 388785 304128 388831
rect 303934 388779 303946 388785
rect 303998 388779 304010 388785
rect 304062 388779 304074 388785
rect 304126 388779 304138 388785
rect 303882 388773 304190 388779
rect 310934 388843 310946 388865
rect 310998 388843 311010 388865
rect 311062 388843 311074 388865
rect 311126 388843 311138 388865
rect 310882 388841 311190 388843
rect 310882 388831 310888 388841
rect 310944 388831 310968 388841
rect 311024 388831 311048 388841
rect 311104 388831 311128 388841
rect 311184 388831 311190 388841
rect 310944 388785 310946 388831
rect 311126 388785 311128 388831
rect 310934 388779 310946 388785
rect 310998 388779 311010 388785
rect 311062 388779 311074 388785
rect 311126 388779 311138 388785
rect 310882 388773 311190 388779
rect 301594 388648 301650 388657
rect 301594 388583 301650 388592
rect 309506 388648 309562 388657
rect 309506 388583 309562 388592
rect 295064 388544 295116 388550
rect 295064 388486 295116 388492
rect 295076 374746 295104 388486
rect 301608 388296 301636 388583
rect 305890 388512 305946 388521
rect 305890 388447 305946 388456
rect 301596 388290 301648 388296
rect 301596 388232 301648 388238
rect 305904 388212 305932 388447
rect 309520 388090 309548 388583
rect 314304 388385 314332 448151
rect 314474 427408 314530 427417
rect 314474 427343 314530 427352
rect 314382 390688 314438 390697
rect 314382 390623 314438 390632
rect 314290 388376 314346 388385
rect 314290 388311 314346 388320
rect 309520 388062 309640 388090
rect 295150 388004 295458 388010
rect 295202 387998 295214 388004
rect 295266 387998 295278 388004
rect 295330 387998 295342 388004
rect 295394 387998 295406 388004
rect 295212 387952 295214 387998
rect 295394 387952 295396 387998
rect 295150 387942 295156 387952
rect 295212 387942 295236 387952
rect 295292 387942 295316 387952
rect 295372 387942 295396 387952
rect 295452 387942 295458 387952
rect 295150 387940 295458 387942
rect 295202 387918 295214 387940
rect 295266 387918 295278 387940
rect 295330 387918 295342 387940
rect 295394 387918 295406 387940
rect 295212 387888 295214 387918
rect 295394 387888 295396 387918
rect 295150 387876 295156 387888
rect 295212 387876 295236 387888
rect 295292 387876 295316 387888
rect 295372 387876 295396 387888
rect 295452 387876 295458 387888
rect 295212 387862 295214 387876
rect 295394 387862 295396 387876
rect 295202 387838 295214 387862
rect 295266 387838 295278 387862
rect 295330 387838 295342 387862
rect 295394 387838 295406 387862
rect 295212 387824 295214 387838
rect 295394 387824 295396 387838
rect 295150 387812 295156 387824
rect 295212 387812 295236 387824
rect 295292 387812 295316 387824
rect 295372 387812 295396 387824
rect 295452 387812 295458 387824
rect 295212 387782 295214 387812
rect 295394 387782 295396 387812
rect 295202 387760 295214 387782
rect 295266 387760 295278 387782
rect 295330 387760 295342 387782
rect 295394 387760 295406 387782
rect 295150 387758 295458 387760
rect 295150 387748 295156 387758
rect 295212 387748 295236 387758
rect 295292 387748 295316 387758
rect 295372 387748 295396 387758
rect 295452 387748 295458 387758
rect 295212 387702 295214 387748
rect 295394 387702 295396 387748
rect 295202 387696 295214 387702
rect 295266 387696 295278 387702
rect 295330 387696 295342 387702
rect 295394 387696 295406 387702
rect 295150 387690 295458 387696
rect 302150 387999 302458 388005
rect 302202 387993 302214 387999
rect 302266 387993 302278 387999
rect 302330 387993 302342 387999
rect 302394 387993 302406 387999
rect 302212 387947 302214 387993
rect 302394 387947 302396 387993
rect 302150 387937 302156 387947
rect 302212 387937 302236 387947
rect 302292 387937 302316 387947
rect 302372 387937 302396 387947
rect 302452 387937 302458 387947
rect 302150 387935 302458 387937
rect 302202 387913 302214 387935
rect 302266 387913 302278 387935
rect 302330 387913 302342 387935
rect 302394 387913 302406 387935
rect 302212 387883 302214 387913
rect 302394 387883 302396 387913
rect 302150 387871 302156 387883
rect 302212 387871 302236 387883
rect 302292 387871 302316 387883
rect 302372 387871 302396 387883
rect 302452 387871 302458 387883
rect 302212 387857 302214 387871
rect 302394 387857 302396 387871
rect 302202 387833 302214 387857
rect 302266 387833 302278 387857
rect 302330 387833 302342 387857
rect 302394 387833 302406 387857
rect 302212 387819 302214 387833
rect 302394 387819 302396 387833
rect 302150 387807 302156 387819
rect 302212 387807 302236 387819
rect 302292 387807 302316 387819
rect 302372 387807 302396 387819
rect 302452 387807 302458 387819
rect 302212 387777 302214 387807
rect 302394 387777 302396 387807
rect 302202 387755 302214 387777
rect 302266 387755 302278 387777
rect 302330 387755 302342 387777
rect 302394 387755 302406 387777
rect 302150 387753 302458 387755
rect 302150 387743 302156 387753
rect 302212 387743 302236 387753
rect 302292 387743 302316 387753
rect 302372 387743 302396 387753
rect 302452 387743 302458 387753
rect 302212 387697 302214 387743
rect 302394 387697 302396 387743
rect 302202 387691 302214 387697
rect 302266 387691 302278 387697
rect 302330 387691 302342 387697
rect 302394 387691 302406 387697
rect 302150 387685 302458 387691
rect 309150 387999 309458 388005
rect 309202 387993 309214 387999
rect 309266 387993 309278 387999
rect 309330 387993 309342 387999
rect 309394 387993 309406 387999
rect 309212 387947 309214 387993
rect 309394 387947 309396 387993
rect 309150 387937 309156 387947
rect 309212 387937 309236 387947
rect 309292 387937 309316 387947
rect 309372 387937 309396 387947
rect 309452 387937 309458 387947
rect 309150 387935 309458 387937
rect 309202 387913 309214 387935
rect 309266 387913 309278 387935
rect 309330 387913 309342 387935
rect 309394 387913 309406 387935
rect 309212 387883 309214 387913
rect 309394 387883 309396 387913
rect 309150 387871 309156 387883
rect 309212 387871 309236 387883
rect 309292 387871 309316 387883
rect 309372 387871 309396 387883
rect 309452 387871 309458 387883
rect 309212 387857 309214 387871
rect 309394 387857 309396 387871
rect 309202 387833 309214 387857
rect 309266 387833 309278 387857
rect 309330 387833 309342 387857
rect 309394 387833 309406 387857
rect 309212 387819 309214 387833
rect 309394 387819 309396 387833
rect 309150 387807 309156 387819
rect 309212 387807 309236 387819
rect 309292 387807 309316 387819
rect 309372 387807 309396 387819
rect 309452 387807 309458 387819
rect 309212 387777 309214 387807
rect 309394 387777 309396 387807
rect 309202 387755 309214 387777
rect 309266 387755 309278 387777
rect 309330 387755 309342 387777
rect 309394 387755 309406 387777
rect 309150 387753 309458 387755
rect 309150 387743 309156 387753
rect 309212 387743 309236 387753
rect 309292 387743 309316 387753
rect 309372 387743 309396 387753
rect 309452 387743 309458 387753
rect 309212 387697 309214 387743
rect 309394 387697 309396 387743
rect 309202 387691 309214 387697
rect 309266 387691 309278 387697
rect 309330 387691 309342 387697
rect 309394 387691 309406 387697
rect 309150 387685 309458 387691
rect 303964 387398 304020 387407
rect 303964 387333 304020 387342
rect 299296 387085 299348 387091
rect 306748 387085 306800 387091
rect 299296 387027 299348 387033
rect 303160 387048 303212 387054
rect 299308 384985 299336 387027
rect 306748 387027 306800 387033
rect 303160 386990 303212 386996
rect 299294 384976 299350 384985
rect 299294 384911 299350 384920
rect 295064 374740 295116 374746
rect 295064 374682 295116 374688
rect 295064 374536 295116 374542
rect 295064 374478 295116 374484
rect 294972 370796 295024 370802
rect 294972 370738 295024 370744
rect 292488 367464 292540 367470
rect 292488 367406 292540 367412
rect 292500 346390 292528 367406
rect 295076 367198 295104 374478
rect 303172 374241 303200 386990
rect 306760 384305 306788 387027
rect 309612 386345 309640 388062
rect 311044 387515 311100 387524
rect 311044 387450 311100 387459
rect 313328 387410 313356 387532
rect 313292 387382 313356 387410
rect 310428 387085 310480 387091
rect 310428 387027 310480 387033
rect 310058 386472 310114 386481
rect 310058 386407 310114 386416
rect 307666 386336 307722 386345
rect 307666 386271 307722 386280
rect 309598 386336 309654 386345
rect 309598 386271 309654 386280
rect 306746 384296 306802 384305
rect 306746 384231 306802 384240
rect 307680 376754 307708 386271
rect 307588 376726 307708 376754
rect 303158 374232 303214 374241
rect 303158 374167 303214 374176
rect 295248 370796 295300 370802
rect 295248 370738 295300 370744
rect 295260 368529 295288 370738
rect 304538 368928 304594 368937
rect 304538 368863 304594 368872
rect 295246 368520 295302 368529
rect 295246 368455 295302 368464
rect 295064 367192 295116 367198
rect 295064 367134 295116 367140
rect 295076 360194 295104 367134
rect 295076 360166 295196 360194
rect 295168 346526 295196 360166
rect 295260 347857 295288 368455
rect 304552 367985 304580 368863
rect 307588 367985 307616 376726
rect 310072 367985 310100 386407
rect 310440 384849 310468 387027
rect 313292 386481 313320 387382
rect 313278 386472 313334 386481
rect 313278 386407 313334 386416
rect 310426 384840 310482 384849
rect 310426 384775 310482 384784
rect 312542 384840 312598 384849
rect 312542 384775 312598 384784
rect 310978 368928 311034 368937
rect 310978 368863 311034 368872
rect 304538 367976 304594 367985
rect 304538 367911 304594 367920
rect 307574 367976 307630 367985
rect 307574 367911 307630 367920
rect 310058 367976 310114 367985
rect 310058 367911 310114 367920
rect 303909 367568 303965 367577
rect 303909 367503 303965 367512
rect 307574 367568 307630 367577
rect 310058 367568 310114 367577
rect 307574 367503 307630 367512
rect 309888 367526 310058 367554
rect 299754 367296 299810 367305
rect 296720 367290 296772 367296
rect 296720 367232 296772 367238
rect 303923 367268 303951 367503
rect 299754 367238 299756 367240
rect 299808 367238 299810 367240
rect 296732 367198 296760 367232
rect 299754 367231 299810 367238
rect 296720 367192 296772 367198
rect 296720 367134 296772 367140
rect 307588 367094 307616 367503
rect 309888 367094 309916 367526
rect 310058 367503 310114 367512
rect 307588 367066 307708 367094
rect 309888 367066 310055 367094
rect 307680 366450 307708 367066
rect 307668 366444 307720 366450
rect 307668 366386 307720 366392
rect 298652 366084 298704 366090
rect 298652 366026 298704 366032
rect 301688 366084 301740 366090
rect 301688 366026 301740 366032
rect 304724 366084 304776 366090
rect 304724 366026 304776 366032
rect 298664 364177 298692 366026
rect 301700 364313 301728 366026
rect 301686 364304 301742 364313
rect 301686 364239 301742 364248
rect 298650 364168 298706 364177
rect 298650 364103 298706 364112
rect 304736 348401 304764 366026
rect 304722 348392 304778 348401
rect 304722 348327 304778 348336
rect 295246 347848 295302 347857
rect 295246 347783 295302 347792
rect 300858 347848 300914 347857
rect 300858 347783 300914 347792
rect 304446 347848 304502 347857
rect 304446 347783 304502 347792
rect 295156 346520 295208 346526
rect 295156 346462 295208 346468
rect 292488 346384 292540 346390
rect 292488 346326 292540 346332
rect 292500 325310 292528 346326
rect 292488 325304 292540 325310
rect 292488 325246 292540 325252
rect 292500 304366 292528 325246
rect 295168 324630 295196 346462
rect 295260 327185 295288 347783
rect 296882 347087 297190 347093
rect 296934 347081 296946 347087
rect 296998 347081 297010 347087
rect 297062 347081 297074 347087
rect 297126 347081 297138 347087
rect 296944 347035 296946 347081
rect 297126 347035 297128 347081
rect 296882 347025 296888 347035
rect 296944 347025 296968 347035
rect 297024 347025 297048 347035
rect 297104 347025 297128 347035
rect 297184 347025 297190 347035
rect 296882 347023 297190 347025
rect 296934 347001 296946 347023
rect 296998 347001 297010 347023
rect 297062 347001 297074 347023
rect 297126 347001 297138 347023
rect 296944 346971 296946 347001
rect 297126 346971 297128 347001
rect 296882 346959 296888 346971
rect 296944 346959 296968 346971
rect 297024 346959 297048 346971
rect 297104 346959 297128 346971
rect 297184 346959 297190 346971
rect 296944 346945 296946 346959
rect 297126 346945 297128 346959
rect 296934 346921 296946 346945
rect 296998 346921 297010 346945
rect 297062 346921 297074 346945
rect 297126 346921 297138 346945
rect 296944 346907 296946 346921
rect 297126 346907 297128 346921
rect 296882 346895 296888 346907
rect 296944 346895 296968 346907
rect 297024 346895 297048 346907
rect 297104 346895 297128 346907
rect 297184 346895 297190 346907
rect 300872 346905 300900 347783
rect 303882 347087 304190 347093
rect 303934 347081 303946 347087
rect 303998 347081 304010 347087
rect 304062 347081 304074 347087
rect 304126 347081 304138 347087
rect 303944 347035 303946 347081
rect 304126 347035 304128 347081
rect 303882 347025 303888 347035
rect 303944 347025 303968 347035
rect 304024 347025 304048 347035
rect 304104 347025 304128 347035
rect 304184 347025 304190 347035
rect 303882 347023 304190 347025
rect 303934 347001 303946 347023
rect 303998 347001 304010 347023
rect 304062 347001 304074 347023
rect 304126 347001 304138 347023
rect 303944 346971 303946 347001
rect 304126 346971 304128 347001
rect 303882 346959 303888 346971
rect 303944 346959 303968 346971
rect 304024 346959 304048 346971
rect 304104 346959 304128 346971
rect 304184 346959 304190 346971
rect 303944 346945 303946 346959
rect 304126 346945 304128 346959
rect 303934 346921 303946 346945
rect 303998 346921 304010 346945
rect 304062 346921 304074 346945
rect 304126 346921 304138 346945
rect 303944 346907 303946 346921
rect 304126 346907 304128 346921
rect 296944 346865 296946 346895
rect 297126 346865 297128 346895
rect 296934 346843 296946 346865
rect 296998 346843 297010 346865
rect 297062 346843 297074 346865
rect 297126 346843 297138 346865
rect 296882 346841 297190 346843
rect 296882 346831 296888 346841
rect 296944 346831 296968 346841
rect 297024 346831 297048 346841
rect 297104 346831 297128 346841
rect 297184 346831 297190 346841
rect 300858 346896 300914 346905
rect 300858 346831 300914 346840
rect 303882 346895 303888 346907
rect 303944 346895 303968 346907
rect 304024 346895 304048 346907
rect 304104 346895 304128 346907
rect 304184 346895 304190 346907
rect 304460 346905 304488 347783
rect 307680 347313 307708 366386
rect 307944 366376 307996 366382
rect 307944 366318 307996 366324
rect 310027 366330 310055 367066
rect 307956 363089 307984 366318
rect 310027 366302 310100 366330
rect 310072 365786 310100 366302
rect 310072 365758 310560 365786
rect 307942 363080 307998 363089
rect 307942 363015 307998 363024
rect 307666 347304 307722 347313
rect 307666 347239 307722 347248
rect 307680 346905 307708 347239
rect 310532 347206 310560 365758
rect 310992 347857 311020 368863
rect 310978 347848 311034 347857
rect 310978 347783 311034 347792
rect 310520 347200 310572 347206
rect 310520 347142 310572 347148
rect 310532 346905 310560 347142
rect 303944 346865 303946 346895
rect 304126 346865 304128 346895
rect 303934 346843 303946 346865
rect 303998 346843 304010 346865
rect 304062 346843 304074 346865
rect 304126 346843 304138 346865
rect 303882 346841 304190 346843
rect 303882 346831 303888 346841
rect 303944 346831 303968 346841
rect 304024 346831 304048 346841
rect 304104 346831 304128 346841
rect 304184 346831 304190 346841
rect 304446 346896 304502 346905
rect 304446 346831 304502 346840
rect 307666 346896 307722 346905
rect 307666 346831 307722 346840
rect 310518 346896 310574 346905
rect 310518 346831 310574 346840
rect 296944 346785 296946 346831
rect 297126 346785 297128 346831
rect 296934 346779 296946 346785
rect 296998 346779 297010 346785
rect 297062 346779 297074 346785
rect 297126 346779 297138 346785
rect 296882 346773 297190 346779
rect 303944 346785 303946 346831
rect 304126 346785 304128 346831
rect 303934 346779 303946 346785
rect 303998 346779 304010 346785
rect 304062 346779 304074 346785
rect 304126 346779 304138 346785
rect 303882 346773 304190 346779
rect 300858 346624 300914 346633
rect 300858 346559 300914 346568
rect 303894 346624 303950 346633
rect 303894 346559 303950 346568
rect 306746 346624 306802 346633
rect 306746 346559 306802 346568
rect 309874 346624 309930 346633
rect 309874 346559 309930 346568
rect 300872 346174 300900 346559
rect 303908 346202 303936 346559
rect 306760 346202 306788 346559
rect 309888 346202 309916 346559
rect 303908 346174 303942 346202
rect 306760 346174 306880 346202
rect 309888 346174 310046 346202
rect 306852 346066 306880 346174
rect 306852 346038 306994 346066
rect 302150 345985 302458 345991
rect 302202 345979 302214 345985
rect 302266 345979 302278 345985
rect 302330 345979 302342 345985
rect 302394 345979 302406 345985
rect 302212 345933 302214 345979
rect 302394 345933 302396 345979
rect 302150 345923 302156 345933
rect 302212 345923 302236 345933
rect 302292 345923 302316 345933
rect 302372 345923 302396 345933
rect 302452 345923 302458 345933
rect 302150 345921 302458 345923
rect 302202 345899 302214 345921
rect 302266 345899 302278 345921
rect 302330 345899 302342 345921
rect 302394 345899 302406 345921
rect 302212 345869 302214 345899
rect 302394 345869 302396 345899
rect 302150 345857 302156 345869
rect 302212 345857 302236 345869
rect 302292 345857 302316 345869
rect 302372 345857 302396 345869
rect 302452 345857 302458 345869
rect 302212 345843 302214 345857
rect 302394 345843 302396 345857
rect 302202 345819 302214 345843
rect 302266 345819 302278 345843
rect 302330 345819 302342 345843
rect 302394 345819 302406 345843
rect 302212 345805 302214 345819
rect 302394 345805 302396 345819
rect 302150 345793 302156 345805
rect 302212 345793 302236 345805
rect 302292 345793 302316 345805
rect 302372 345793 302396 345805
rect 302452 345793 302458 345805
rect 302212 345763 302214 345793
rect 302394 345763 302396 345793
rect 302202 345741 302214 345763
rect 302266 345741 302278 345763
rect 302330 345741 302342 345763
rect 302394 345741 302406 345763
rect 302150 345739 302458 345741
rect 302150 345729 302156 345739
rect 302212 345729 302236 345739
rect 302292 345729 302316 345739
rect 302372 345729 302396 345739
rect 302452 345729 302458 345739
rect 302212 345683 302214 345729
rect 302394 345683 302396 345729
rect 302202 345677 302214 345683
rect 302266 345677 302278 345683
rect 302330 345677 302342 345683
rect 302394 345677 302406 345683
rect 302150 345671 302458 345677
rect 309150 345985 309458 345991
rect 309202 345979 309214 345985
rect 309266 345979 309278 345985
rect 309330 345979 309342 345985
rect 309394 345979 309406 345985
rect 309212 345933 309214 345979
rect 309394 345933 309396 345979
rect 309150 345923 309156 345933
rect 309212 345923 309236 345933
rect 309292 345923 309316 345933
rect 309372 345923 309396 345933
rect 309452 345923 309458 345933
rect 309150 345921 309458 345923
rect 309202 345899 309214 345921
rect 309266 345899 309278 345921
rect 309330 345899 309342 345921
rect 309394 345899 309406 345921
rect 309212 345869 309214 345899
rect 309394 345869 309396 345899
rect 309150 345857 309156 345869
rect 309212 345857 309236 345869
rect 309292 345857 309316 345869
rect 309372 345857 309396 345869
rect 309452 345857 309458 345869
rect 309212 345843 309214 345857
rect 309394 345843 309396 345857
rect 309202 345819 309214 345843
rect 309266 345819 309278 345843
rect 309330 345819 309342 345843
rect 309394 345819 309406 345843
rect 309212 345805 309214 345819
rect 309394 345805 309396 345819
rect 309150 345793 309156 345805
rect 309212 345793 309236 345805
rect 309292 345793 309316 345805
rect 309372 345793 309396 345805
rect 309452 345793 309458 345805
rect 309212 345763 309214 345793
rect 309394 345763 309396 345793
rect 309202 345741 309214 345763
rect 309266 345741 309278 345763
rect 309330 345741 309342 345763
rect 309394 345741 309406 345763
rect 309150 345739 309458 345741
rect 309150 345729 309156 345739
rect 309212 345729 309236 345739
rect 309292 345729 309316 345739
rect 309372 345729 309396 345739
rect 309452 345729 309458 345739
rect 309212 345683 309214 345729
rect 309394 345683 309396 345729
rect 309202 345677 309214 345683
rect 309266 345677 309278 345683
rect 309330 345677 309342 345683
rect 309394 345677 309406 345683
rect 309150 345671 309458 345677
rect 307944 345092 307996 345098
rect 298652 345084 298704 345090
rect 298652 345026 298704 345032
rect 301688 345084 301740 345090
rect 301688 345026 301740 345032
rect 304724 345084 304776 345090
rect 307944 345034 307996 345040
rect 304724 345026 304776 345032
rect 298664 343505 298692 345026
rect 301700 343641 301728 345026
rect 301686 343632 301742 343641
rect 301686 343567 301742 343576
rect 298650 343496 298706 343505
rect 298650 343431 298706 343440
rect 304736 331537 304764 345026
rect 307956 342281 307984 345034
rect 307942 342272 307998 342281
rect 307942 342207 307998 342216
rect 307666 340232 307722 340241
rect 307666 340167 307722 340176
rect 304722 331528 304778 331537
rect 304722 331463 304778 331472
rect 304906 327720 304962 327729
rect 304906 327655 304962 327664
rect 295246 327176 295302 327185
rect 295246 327111 295302 327120
rect 300858 327176 300914 327185
rect 300858 327111 300914 327120
rect 295156 324624 295208 324630
rect 295156 324566 295208 324572
rect 292488 304360 292540 304366
rect 292488 304302 292540 304308
rect 292500 283286 292528 304302
rect 295168 304230 295196 324566
rect 295260 306513 295288 327111
rect 296882 326086 297190 326092
rect 296934 326080 296946 326086
rect 296998 326080 297010 326086
rect 297062 326080 297074 326086
rect 297126 326080 297138 326086
rect 296944 326034 296946 326080
rect 297126 326034 297128 326080
rect 296882 326024 296888 326034
rect 296944 326024 296968 326034
rect 297024 326024 297048 326034
rect 297104 326024 297128 326034
rect 297184 326024 297190 326034
rect 296882 326022 297190 326024
rect 296934 326000 296946 326022
rect 296998 326000 297010 326022
rect 297062 326000 297074 326022
rect 297126 326000 297138 326022
rect 296944 325970 296946 326000
rect 297126 325970 297128 326000
rect 296882 325958 296888 325970
rect 296944 325958 296968 325970
rect 297024 325958 297048 325970
rect 297104 325958 297128 325970
rect 297184 325958 297190 325970
rect 300872 325961 300900 327111
rect 303882 326086 304190 326092
rect 303934 326080 303946 326086
rect 303998 326080 304010 326086
rect 304062 326080 304074 326086
rect 304126 326080 304138 326086
rect 303944 326034 303946 326080
rect 304126 326034 304128 326080
rect 303882 326024 303888 326034
rect 303944 326024 303968 326034
rect 304024 326024 304048 326034
rect 304104 326024 304128 326034
rect 304184 326024 304190 326034
rect 303882 326022 304190 326024
rect 303934 326000 303946 326022
rect 303998 326000 304010 326022
rect 304062 326000 304074 326022
rect 304126 326000 304138 326022
rect 303944 325970 303946 326000
rect 304126 325970 304128 326000
rect 296944 325944 296946 325958
rect 297126 325944 297128 325958
rect 296934 325920 296946 325944
rect 296998 325920 297010 325944
rect 297062 325920 297074 325944
rect 297126 325920 297138 325944
rect 296944 325906 296946 325920
rect 297126 325906 297128 325920
rect 296882 325894 296888 325906
rect 296944 325894 296968 325906
rect 297024 325894 297048 325906
rect 297104 325894 297128 325906
rect 297184 325894 297190 325906
rect 296944 325864 296946 325894
rect 297126 325864 297128 325894
rect 300858 325952 300914 325961
rect 300858 325887 300914 325896
rect 303882 325958 303888 325970
rect 303944 325958 303968 325970
rect 304024 325958 304048 325970
rect 304104 325958 304128 325970
rect 304184 325958 304190 325970
rect 304920 325961 304948 327655
rect 307680 326233 307708 340167
rect 310992 328409 311020 347783
rect 311440 347200 311492 347206
rect 311440 347142 311492 347148
rect 311070 346760 311126 346769
rect 311070 346695 311126 346704
rect 311084 340241 311112 346695
rect 311452 345014 311480 347142
rect 311452 344986 311572 345014
rect 311070 340232 311126 340241
rect 311070 340167 311126 340176
rect 310978 328400 311034 328409
rect 310978 328335 311034 328344
rect 310992 327729 311020 328335
rect 310978 327720 311034 327729
rect 310978 327655 311034 327664
rect 307666 326224 307722 326233
rect 307666 326159 307722 326168
rect 307680 325961 307708 326159
rect 310882 326086 311190 326092
rect 310934 326080 310946 326086
rect 310998 326080 311010 326086
rect 311062 326080 311074 326086
rect 311126 326080 311138 326086
rect 310944 326034 310946 326080
rect 311126 326034 311128 326080
rect 310882 326024 310888 326034
rect 310944 326024 310968 326034
rect 311024 326024 311048 326034
rect 311104 326024 311128 326034
rect 311184 326024 311190 326034
rect 310882 326022 311190 326024
rect 310934 326000 310946 326022
rect 310998 326000 311010 326022
rect 311062 326000 311074 326022
rect 311126 326000 311138 326022
rect 310944 325970 310946 326000
rect 311126 325970 311128 326000
rect 303944 325944 303946 325958
rect 304126 325944 304128 325958
rect 303934 325920 303946 325944
rect 303998 325920 304010 325944
rect 304062 325920 304074 325944
rect 304126 325920 304138 325944
rect 303944 325906 303946 325920
rect 304126 325906 304128 325920
rect 303882 325894 303888 325906
rect 303944 325894 303968 325906
rect 304024 325894 304048 325906
rect 304104 325894 304128 325906
rect 304184 325894 304190 325906
rect 296934 325842 296946 325864
rect 296998 325842 297010 325864
rect 297062 325842 297074 325864
rect 297126 325842 297138 325864
rect 296882 325840 297190 325842
rect 296882 325830 296888 325840
rect 296944 325830 296968 325840
rect 297024 325830 297048 325840
rect 297104 325830 297128 325840
rect 297184 325830 297190 325840
rect 296944 325784 296946 325830
rect 297126 325784 297128 325830
rect 296934 325778 296946 325784
rect 296998 325778 297010 325784
rect 297062 325778 297074 325784
rect 297126 325778 297138 325784
rect 296882 325772 297190 325778
rect 303944 325864 303946 325894
rect 304126 325864 304128 325894
rect 304906 325952 304962 325961
rect 304906 325887 304962 325896
rect 307666 325952 307722 325961
rect 307666 325887 307722 325896
rect 310882 325958 310888 325970
rect 310944 325958 310968 325970
rect 311024 325958 311048 325970
rect 311104 325958 311128 325970
rect 311184 325958 311190 325970
rect 310944 325944 310946 325958
rect 311126 325944 311128 325958
rect 310934 325920 310946 325944
rect 310998 325920 311010 325944
rect 311062 325920 311074 325944
rect 311126 325920 311138 325944
rect 310944 325906 310946 325920
rect 311126 325906 311128 325920
rect 310882 325894 310888 325906
rect 310944 325894 310968 325906
rect 311024 325894 311048 325906
rect 311104 325894 311128 325906
rect 311184 325894 311190 325906
rect 303934 325842 303946 325864
rect 303998 325842 304010 325864
rect 304062 325842 304074 325864
rect 304126 325842 304138 325864
rect 303882 325840 304190 325842
rect 303882 325830 303888 325840
rect 303944 325830 303968 325840
rect 304024 325830 304048 325840
rect 304104 325830 304128 325840
rect 304184 325830 304190 325840
rect 303944 325784 303946 325830
rect 304126 325784 304128 325830
rect 303934 325778 303946 325784
rect 303998 325778 304010 325784
rect 304062 325778 304074 325784
rect 304126 325778 304138 325784
rect 303882 325772 304190 325778
rect 310944 325864 310946 325894
rect 311126 325864 311128 325894
rect 310934 325842 310946 325864
rect 310998 325842 311010 325864
rect 311062 325842 311074 325864
rect 311126 325842 311138 325864
rect 310882 325840 311190 325842
rect 310882 325830 310888 325840
rect 310944 325830 310968 325840
rect 311024 325830 311048 325840
rect 311104 325830 311128 325840
rect 311184 325830 311190 325840
rect 310944 325784 310946 325830
rect 311126 325784 311128 325830
rect 310934 325778 310946 325784
rect 310998 325778 311010 325784
rect 311062 325778 311074 325784
rect 311126 325778 311138 325784
rect 310882 325772 311190 325778
rect 300950 325680 301006 325689
rect 300950 325615 301006 325624
rect 304262 325680 304318 325689
rect 304262 325615 304318 325624
rect 307390 325680 307446 325689
rect 307390 325615 307446 325624
rect 300964 325258 300992 325615
rect 300964 325230 301104 325258
rect 304276 325244 304304 325615
rect 307404 325244 307432 325615
rect 310559 324306 310587 324428
rect 311544 324306 311572 344986
rect 311898 328400 311954 328409
rect 311898 328335 311954 328344
rect 310559 324278 310652 324306
rect 310624 324170 310652 324278
rect 311268 324278 311572 324306
rect 311268 324170 311296 324278
rect 298756 321473 298784 324156
rect 301780 324080 301832 324086
rect 301780 324022 301832 324028
rect 298742 321464 298798 321473
rect 298742 321399 298798 321408
rect 301792 321337 301820 324022
rect 303882 323914 304190 323920
rect 303934 323908 303946 323914
rect 303998 323908 304010 323914
rect 304062 323908 304074 323914
rect 304126 323908 304138 323914
rect 303944 323862 303946 323908
rect 304126 323862 304128 323908
rect 303882 323852 303888 323862
rect 303944 323852 303968 323862
rect 304024 323852 304048 323862
rect 304104 323852 304128 323862
rect 304184 323852 304190 323862
rect 303882 323850 304190 323852
rect 303934 323828 303946 323850
rect 303998 323828 304010 323850
rect 304062 323828 304074 323850
rect 304126 323828 304138 323850
rect 303944 323798 303946 323828
rect 304126 323798 304128 323828
rect 303882 323786 303888 323798
rect 303944 323786 303968 323798
rect 304024 323786 304048 323798
rect 304104 323786 304128 323798
rect 304184 323786 304190 323798
rect 303944 323772 303946 323786
rect 304126 323772 304128 323786
rect 303934 323748 303946 323772
rect 303998 323748 304010 323772
rect 304062 323748 304074 323772
rect 304126 323748 304138 323772
rect 303944 323734 303946 323748
rect 304126 323734 304128 323748
rect 303882 323722 303888 323734
rect 303944 323722 303968 323734
rect 304024 323722 304048 323734
rect 304104 323722 304128 323734
rect 304184 323722 304190 323734
rect 303944 323692 303946 323722
rect 304126 323692 304128 323722
rect 303934 323670 303946 323692
rect 303998 323670 304010 323692
rect 304062 323670 304074 323692
rect 304126 323670 304138 323692
rect 303882 323668 304190 323670
rect 303882 323658 303888 323668
rect 303944 323658 303968 323668
rect 304024 323658 304048 323668
rect 304104 323658 304128 323668
rect 304184 323658 304190 323668
rect 303944 323612 303946 323658
rect 304126 323612 304128 323658
rect 303934 323606 303946 323612
rect 303998 323606 304010 323612
rect 304062 323606 304074 323612
rect 304126 323606 304138 323612
rect 303882 323600 304190 323606
rect 305104 322833 305132 324156
rect 305090 322824 305146 322833
rect 305090 322759 305146 322768
rect 301778 321328 301834 321337
rect 301778 321263 301834 321272
rect 308232 308417 308260 324156
rect 310624 324142 311296 324170
rect 308218 308408 308274 308417
rect 308218 308343 308274 308352
rect 306194 307456 306250 307465
rect 306194 307391 306250 307400
rect 295246 306504 295302 306513
rect 295246 306439 295302 306448
rect 301686 306504 301742 306513
rect 301686 306439 301742 306448
rect 295156 304224 295208 304230
rect 295156 304166 295208 304172
rect 295260 294545 295288 306439
rect 296882 305116 297190 305122
rect 296934 305110 296946 305116
rect 296998 305110 297010 305116
rect 297062 305110 297074 305116
rect 297126 305110 297138 305116
rect 296944 305064 296946 305110
rect 297126 305064 297128 305110
rect 296882 305054 296888 305064
rect 296944 305054 296968 305064
rect 297024 305054 297048 305064
rect 297104 305054 297128 305064
rect 297184 305054 297190 305064
rect 296882 305052 297190 305054
rect 296934 305030 296946 305052
rect 296998 305030 297010 305052
rect 297062 305030 297074 305052
rect 297126 305030 297138 305052
rect 296944 305000 296946 305030
rect 297126 305000 297128 305030
rect 301700 305017 301728 306439
rect 303882 305116 304190 305122
rect 303934 305110 303946 305116
rect 303998 305110 304010 305116
rect 304062 305110 304074 305116
rect 304126 305110 304138 305116
rect 303944 305064 303946 305110
rect 304126 305064 304128 305110
rect 303882 305054 303888 305064
rect 303944 305054 303968 305064
rect 304024 305054 304048 305064
rect 304104 305054 304128 305064
rect 304184 305054 304190 305064
rect 303882 305052 304190 305054
rect 303934 305030 303946 305052
rect 303998 305030 304010 305052
rect 304062 305030 304074 305052
rect 304126 305030 304138 305052
rect 296882 304988 296888 305000
rect 296944 304988 296968 305000
rect 297024 304988 297048 305000
rect 297104 304988 297128 305000
rect 297184 304988 297190 305000
rect 296944 304974 296946 304988
rect 297126 304974 297128 304988
rect 296934 304950 296946 304974
rect 296998 304950 297010 304974
rect 297062 304950 297074 304974
rect 297126 304950 297138 304974
rect 296944 304936 296946 304950
rect 297126 304936 297128 304950
rect 301686 305008 301742 305017
rect 301686 304943 301742 304952
rect 303944 305000 303946 305030
rect 304126 305000 304128 305030
rect 306208 305017 306236 307391
rect 310624 305017 310652 324142
rect 310882 323914 311190 323920
rect 310934 323908 310946 323914
rect 310998 323908 311010 323914
rect 311062 323908 311074 323914
rect 311126 323908 311138 323914
rect 310944 323862 310946 323908
rect 311126 323862 311128 323908
rect 310882 323852 310888 323862
rect 310944 323852 310968 323862
rect 311024 323852 311048 323862
rect 311104 323852 311128 323862
rect 311184 323852 311190 323862
rect 310882 323850 311190 323852
rect 310934 323828 310946 323850
rect 310998 323828 311010 323850
rect 311062 323828 311074 323850
rect 311126 323828 311138 323850
rect 310944 323798 310946 323828
rect 311126 323798 311128 323828
rect 310882 323786 310888 323798
rect 310944 323786 310968 323798
rect 311024 323786 311048 323798
rect 311104 323786 311128 323798
rect 311184 323786 311190 323798
rect 310944 323772 310946 323786
rect 311126 323772 311128 323786
rect 310934 323748 310946 323772
rect 310998 323748 311010 323772
rect 311062 323748 311074 323772
rect 311126 323748 311138 323772
rect 310944 323734 310946 323748
rect 311126 323734 311128 323748
rect 310882 323722 310888 323734
rect 310944 323722 310968 323734
rect 311024 323722 311048 323734
rect 311104 323722 311128 323734
rect 311184 323722 311190 323734
rect 310944 323692 310946 323722
rect 311126 323692 311128 323722
rect 310934 323670 310946 323692
rect 310998 323670 311010 323692
rect 311062 323670 311074 323692
rect 311126 323670 311138 323692
rect 310882 323668 311190 323670
rect 310882 323658 310888 323668
rect 310944 323658 310968 323668
rect 311024 323658 311048 323668
rect 311104 323658 311128 323668
rect 311184 323658 311190 323668
rect 310944 323612 310946 323658
rect 311126 323612 311128 323658
rect 310934 323606 310946 323612
rect 310998 323606 311010 323612
rect 311062 323606 311074 323612
rect 311126 323606 311138 323612
rect 310882 323600 311190 323606
rect 311912 307465 311940 328335
rect 311990 326224 312046 326233
rect 311990 326159 312046 326168
rect 311898 307456 311954 307465
rect 311898 307391 311954 307400
rect 312004 306513 312032 326159
rect 312556 307057 312584 384775
rect 314396 368937 314424 390623
rect 314488 388521 314516 427343
rect 314568 408468 314620 408474
rect 314568 408410 314620 408416
rect 314474 388512 314530 388521
rect 314474 388447 314530 388456
rect 314580 386481 314608 408410
rect 314566 386472 314622 386481
rect 314566 386407 314622 386416
rect 314382 368928 314438 368937
rect 314382 368863 314438 368872
rect 314014 366072 314070 366081
rect 314014 366007 314070 366016
rect 313924 364404 313976 364410
rect 313924 364346 313976 364352
rect 312910 363080 312966 363089
rect 312910 363015 312966 363024
rect 312634 342272 312690 342281
rect 312634 342207 312690 342216
rect 312648 325009 312676 342207
rect 312634 325000 312690 325009
rect 312634 324935 312690 324944
rect 312924 307193 312952 363015
rect 313738 307456 313794 307465
rect 313738 307391 313794 307400
rect 312910 307184 312966 307193
rect 312910 307119 312966 307128
rect 312542 307048 312598 307057
rect 312542 306983 312598 306992
rect 311990 306504 312046 306513
rect 311990 306439 312046 306448
rect 313646 306504 313702 306513
rect 313646 306439 313702 306448
rect 310882 305116 311190 305122
rect 310934 305110 310946 305116
rect 310998 305110 311010 305116
rect 311062 305110 311074 305116
rect 311126 305110 311138 305116
rect 310944 305064 310946 305110
rect 311126 305064 311128 305110
rect 310882 305054 310888 305064
rect 310944 305054 310968 305064
rect 311024 305054 311048 305064
rect 311104 305054 311128 305064
rect 311184 305054 311190 305064
rect 310882 305052 311190 305054
rect 310934 305030 310946 305052
rect 310998 305030 311010 305052
rect 311062 305030 311074 305052
rect 311126 305030 311138 305052
rect 303882 304988 303888 305000
rect 303944 304988 303968 305000
rect 304024 304988 304048 305000
rect 304104 304988 304128 305000
rect 304184 304988 304190 305000
rect 303944 304974 303946 304988
rect 304126 304974 304128 304988
rect 303934 304950 303946 304974
rect 303998 304950 304010 304974
rect 304062 304950 304074 304974
rect 304126 304950 304138 304974
rect 296882 304924 296888 304936
rect 296944 304924 296968 304936
rect 297024 304924 297048 304936
rect 297104 304924 297128 304936
rect 297184 304924 297190 304936
rect 296944 304894 296946 304924
rect 297126 304894 297128 304924
rect 296934 304872 296946 304894
rect 296998 304872 297010 304894
rect 297062 304872 297074 304894
rect 297126 304872 297138 304894
rect 296882 304870 297190 304872
rect 296882 304860 296888 304870
rect 296944 304860 296968 304870
rect 297024 304860 297048 304870
rect 297104 304860 297128 304870
rect 297184 304860 297190 304870
rect 296944 304814 296946 304860
rect 297126 304814 297128 304860
rect 296934 304808 296946 304814
rect 296998 304808 297010 304814
rect 297062 304808 297074 304814
rect 297126 304808 297138 304814
rect 296882 304802 297190 304808
rect 303944 304936 303946 304950
rect 304126 304936 304128 304950
rect 306194 305008 306250 305017
rect 306194 304943 306250 304952
rect 310610 305008 310666 305017
rect 310610 304943 310666 304952
rect 310944 305000 310946 305030
rect 311126 305000 311128 305030
rect 310882 304988 310888 305000
rect 310944 304988 310968 305000
rect 311024 304988 311048 305000
rect 311104 304988 311128 305000
rect 311184 304988 311190 305000
rect 310944 304974 310946 304988
rect 311126 304974 311128 304988
rect 310934 304950 310946 304974
rect 310998 304950 311010 304974
rect 311062 304950 311074 304974
rect 311126 304950 311138 304974
rect 303882 304924 303888 304936
rect 303944 304924 303968 304936
rect 304024 304924 304048 304936
rect 304104 304924 304128 304936
rect 304184 304924 304190 304936
rect 303944 304894 303946 304924
rect 304126 304894 304128 304924
rect 303934 304872 303946 304894
rect 303998 304872 304010 304894
rect 304062 304872 304074 304894
rect 304126 304872 304138 304894
rect 303882 304870 304190 304872
rect 303882 304860 303888 304870
rect 303944 304860 303968 304870
rect 304024 304860 304048 304870
rect 304104 304860 304128 304870
rect 304184 304860 304190 304870
rect 303944 304814 303946 304860
rect 304126 304814 304128 304860
rect 303934 304808 303946 304814
rect 303998 304808 304010 304814
rect 304062 304808 304074 304814
rect 304126 304808 304138 304814
rect 303882 304802 304190 304808
rect 310944 304936 310946 304950
rect 311126 304936 311128 304950
rect 310882 304924 310888 304936
rect 310944 304924 310968 304936
rect 311024 304924 311048 304936
rect 311104 304924 311128 304936
rect 311184 304924 311190 304936
rect 310944 304894 310946 304924
rect 311126 304894 311128 304924
rect 310934 304872 310946 304894
rect 310998 304872 311010 304894
rect 311062 304872 311074 304894
rect 311126 304872 311138 304894
rect 310882 304870 311190 304872
rect 310882 304860 310888 304870
rect 310944 304860 310968 304870
rect 311024 304860 311048 304870
rect 311104 304860 311128 304870
rect 311184 304860 311190 304870
rect 310944 304814 310946 304860
rect 311126 304814 311128 304860
rect 310934 304808 310946 304814
rect 310998 304808 311010 304814
rect 311062 304808 311074 304814
rect 311126 304808 311138 304814
rect 310882 304802 311190 304808
rect 301956 304600 302012 304609
rect 301956 304535 302012 304544
rect 305550 304600 305606 304609
rect 305550 304535 305606 304544
rect 312358 304600 312414 304609
rect 312358 304535 312414 304544
rect 297456 304319 297508 304325
rect 301970 304300 301998 304535
rect 305564 304300 305592 304535
rect 312372 304325 312400 304535
rect 312360 304319 312412 304325
rect 297456 304261 297508 304267
rect 312360 304261 312412 304267
rect 297468 304230 297496 304261
rect 297456 304224 297508 304230
rect 297456 304166 297508 304172
rect 298100 304224 298152 304230
rect 298100 304166 298152 304172
rect 298112 303906 298140 304166
rect 312372 304162 312400 304261
rect 312360 304156 312412 304162
rect 312360 304098 312412 304104
rect 302150 304015 302458 304021
rect 302202 304009 302214 304015
rect 302266 304009 302278 304015
rect 302330 304009 302342 304015
rect 302394 304009 302406 304015
rect 302212 303963 302214 304009
rect 302394 303963 302396 304009
rect 302150 303953 302156 303963
rect 302212 303953 302236 303963
rect 302292 303953 302316 303963
rect 302372 303953 302396 303963
rect 302452 303953 302458 303963
rect 302150 303951 302458 303953
rect 302202 303929 302214 303951
rect 302266 303929 302278 303951
rect 302330 303929 302342 303951
rect 302394 303929 302406 303951
rect 298112 303892 298399 303906
rect 302212 303899 302214 303929
rect 302394 303899 302396 303929
rect 298112 303878 298413 303892
rect 298385 303362 298413 303878
rect 302150 303887 302156 303899
rect 302212 303887 302236 303899
rect 302292 303887 302316 303899
rect 302372 303887 302396 303899
rect 302452 303887 302458 303899
rect 302212 303873 302214 303887
rect 302394 303873 302396 303887
rect 302202 303849 302214 303873
rect 302266 303849 302278 303873
rect 302330 303849 302342 303873
rect 302394 303849 302406 303873
rect 302212 303835 302214 303849
rect 302394 303835 302396 303849
rect 302150 303823 302156 303835
rect 302212 303823 302236 303835
rect 302292 303823 302316 303835
rect 302372 303823 302396 303835
rect 302452 303823 302458 303835
rect 302212 303793 302214 303823
rect 302394 303793 302396 303823
rect 302202 303771 302214 303793
rect 302266 303771 302278 303793
rect 302330 303771 302342 303793
rect 302394 303771 302406 303793
rect 302150 303769 302458 303771
rect 302150 303759 302156 303769
rect 302212 303759 302236 303769
rect 302292 303759 302316 303769
rect 302372 303759 302396 303769
rect 302452 303759 302458 303769
rect 302212 303713 302214 303759
rect 302394 303713 302396 303759
rect 302202 303707 302214 303713
rect 302266 303707 302278 303713
rect 302330 303707 302342 303713
rect 302394 303707 302406 303713
rect 302150 303701 302458 303707
rect 309150 304015 309458 304021
rect 309202 304009 309214 304015
rect 309266 304009 309278 304015
rect 309330 304009 309342 304015
rect 309394 304009 309406 304015
rect 309212 303963 309214 304009
rect 309394 303963 309396 304009
rect 309150 303953 309156 303963
rect 309212 303953 309236 303963
rect 309292 303953 309316 303963
rect 309372 303953 309396 303963
rect 309452 303953 309458 303963
rect 309150 303951 309458 303953
rect 309202 303929 309214 303951
rect 309266 303929 309278 303951
rect 309330 303929 309342 303951
rect 309394 303929 309406 303951
rect 309212 303899 309214 303929
rect 309394 303899 309396 303929
rect 309150 303887 309156 303899
rect 309212 303887 309236 303899
rect 309292 303887 309316 303899
rect 309372 303887 309396 303899
rect 309452 303887 309458 303899
rect 309212 303873 309214 303887
rect 309394 303873 309396 303887
rect 309202 303849 309214 303873
rect 309266 303849 309278 303873
rect 309330 303849 309342 303873
rect 309394 303849 309406 303873
rect 309212 303835 309214 303849
rect 309394 303835 309396 303849
rect 309150 303823 309156 303835
rect 309212 303823 309236 303835
rect 309292 303823 309316 303835
rect 309372 303823 309396 303835
rect 309452 303823 309458 303835
rect 309212 303793 309214 303823
rect 309394 303793 309396 303823
rect 309202 303771 309214 303793
rect 309266 303771 309278 303793
rect 309330 303771 309342 303793
rect 309394 303771 309406 303793
rect 309150 303769 309458 303771
rect 309150 303759 309156 303769
rect 309212 303759 309236 303769
rect 309292 303759 309316 303769
rect 309372 303759 309396 303769
rect 309452 303759 309458 303769
rect 309212 303713 309214 303759
rect 309394 303713 309396 303759
rect 309202 303707 309214 303713
rect 309266 303707 309278 303713
rect 309330 303707 309342 303713
rect 309394 303707 309406 303713
rect 309150 303701 309458 303707
rect 298385 303334 298416 303362
rect 298388 296714 298416 303334
rect 299216 302025 299244 303620
rect 299202 302016 299258 302025
rect 299202 301951 299258 301960
rect 302804 301889 302832 303620
rect 306392 302161 306420 303620
rect 306378 302152 306434 302161
rect 306378 302087 306434 302096
rect 302790 301880 302846 301889
rect 302790 301815 302846 301824
rect 298112 296686 298416 296714
rect 295246 294536 295302 294545
rect 295246 294471 295302 294480
rect 295246 284472 295302 284481
rect 295168 284430 295246 284458
rect 292488 283280 292540 283286
rect 292488 283222 292540 283228
rect 292500 262478 292528 283222
rect 295168 277394 295196 284430
rect 295246 284407 295302 284416
rect 298112 284345 298140 296686
rect 299478 294536 299534 294545
rect 299478 294471 299534 294480
rect 299492 284481 299520 294471
rect 309980 288833 310008 303620
rect 313384 303606 313582 303634
rect 313384 303521 313412 303606
rect 313660 303550 313688 306439
rect 313648 303544 313700 303550
rect 313370 303512 313426 303521
rect 313648 303486 313700 303492
rect 313370 303447 313426 303456
rect 313660 302190 313688 303486
rect 313648 302184 313700 302190
rect 313648 302126 313700 302132
rect 309966 288824 310022 288833
rect 309966 288759 310022 288768
rect 313752 288425 313780 307391
rect 313832 304156 313884 304162
rect 313832 304098 313884 304104
rect 311898 288416 311954 288425
rect 311898 288351 311954 288360
rect 313738 288416 313794 288425
rect 313738 288351 313794 288360
rect 311912 287054 311940 288351
rect 311912 287026 312400 287054
rect 308126 285968 308182 285977
rect 308126 285903 308182 285912
rect 304814 285832 304870 285841
rect 304814 285767 304870 285776
rect 299478 284472 299534 284481
rect 299478 284407 299534 284416
rect 295246 284336 295302 284345
rect 295246 284271 295302 284280
rect 298098 284336 298154 284345
rect 298098 284271 298154 284280
rect 295260 277545 295288 284271
rect 299492 283801 299520 284407
rect 304828 283801 304856 285767
rect 308140 283801 308168 285903
rect 312372 285841 312400 287026
rect 312726 285968 312782 285977
rect 312726 285903 312782 285912
rect 312358 285832 312414 285841
rect 312358 285767 312414 285776
rect 299478 283792 299534 283801
rect 299478 283727 299534 283736
rect 304814 283792 304870 283801
rect 304814 283727 304870 283736
rect 308126 283792 308182 283801
rect 308126 283727 308182 283736
rect 299754 283384 299810 283393
rect 298133 283328 298142 283384
rect 298198 283328 298207 283384
rect 299705 283342 299754 283370
rect 304767 283328 304776 283384
rect 304832 283328 304841 283384
rect 308084 283328 308093 283384
rect 308149 283328 308158 283384
rect 299754 283319 299810 283328
rect 302150 283000 302458 283006
rect 302202 282994 302214 283000
rect 302266 282994 302278 283000
rect 302330 282994 302342 283000
rect 302394 282994 302406 283000
rect 302212 282948 302214 282994
rect 302394 282948 302396 282994
rect 302150 282938 302156 282948
rect 302212 282938 302236 282948
rect 302292 282938 302316 282948
rect 302372 282938 302396 282948
rect 302452 282938 302458 282948
rect 302150 282936 302458 282938
rect 302202 282914 302214 282936
rect 302266 282914 302278 282936
rect 302330 282914 302342 282936
rect 302394 282914 302406 282936
rect 302212 282884 302214 282914
rect 302394 282884 302396 282914
rect 302150 282872 302156 282884
rect 302212 282872 302236 282884
rect 302292 282872 302316 282884
rect 302372 282872 302396 282884
rect 302452 282872 302458 282884
rect 302212 282858 302214 282872
rect 302394 282858 302396 282872
rect 302202 282834 302214 282858
rect 302266 282834 302278 282858
rect 302330 282834 302342 282858
rect 302394 282834 302406 282858
rect 302212 282820 302214 282834
rect 302394 282820 302396 282834
rect 302150 282808 302156 282820
rect 302212 282808 302236 282820
rect 302292 282808 302316 282820
rect 302372 282808 302396 282820
rect 302452 282808 302458 282820
rect 302212 282778 302214 282808
rect 302394 282778 302396 282808
rect 302202 282756 302214 282778
rect 302266 282756 302278 282778
rect 302330 282756 302342 282778
rect 302394 282756 302406 282778
rect 302150 282754 302458 282756
rect 302150 282744 302156 282754
rect 302212 282744 302236 282754
rect 302292 282744 302316 282754
rect 302372 282744 302396 282754
rect 302452 282744 302458 282754
rect 302212 282698 302214 282744
rect 302394 282698 302396 282744
rect 302202 282692 302214 282698
rect 302266 282692 302278 282698
rect 302330 282692 302342 282698
rect 302394 282692 302406 282698
rect 302150 282686 302458 282692
rect 309150 283001 309458 283007
rect 309202 282995 309214 283001
rect 309266 282995 309278 283001
rect 309330 282995 309342 283001
rect 309394 282995 309406 283001
rect 309212 282949 309214 282995
rect 309394 282949 309396 282995
rect 309150 282939 309156 282949
rect 309212 282939 309236 282949
rect 309292 282939 309316 282949
rect 309372 282939 309396 282949
rect 309452 282939 309458 282949
rect 309150 282937 309458 282939
rect 309202 282915 309214 282937
rect 309266 282915 309278 282937
rect 309330 282915 309342 282937
rect 309394 282915 309406 282937
rect 309212 282885 309214 282915
rect 309394 282885 309396 282915
rect 309150 282873 309156 282885
rect 309212 282873 309236 282885
rect 309292 282873 309316 282885
rect 309372 282873 309396 282885
rect 309452 282873 309458 282885
rect 309212 282859 309214 282873
rect 309394 282859 309396 282873
rect 309202 282835 309214 282859
rect 309266 282835 309278 282859
rect 309330 282835 309342 282859
rect 309394 282835 309406 282859
rect 309212 282821 309214 282835
rect 309394 282821 309396 282835
rect 309150 282809 309156 282821
rect 309212 282809 309236 282821
rect 309292 282809 309316 282821
rect 309372 282809 309396 282821
rect 309452 282809 309458 282821
rect 309212 282779 309214 282809
rect 309394 282779 309396 282809
rect 309202 282757 309214 282779
rect 309266 282757 309278 282779
rect 309330 282757 309342 282779
rect 309394 282757 309406 282779
rect 309150 282755 309458 282757
rect 309150 282745 309156 282755
rect 309212 282745 309236 282755
rect 309292 282745 309316 282755
rect 309372 282745 309396 282755
rect 309452 282745 309458 282755
rect 309212 282699 309214 282745
rect 309394 282699 309396 282745
rect 309202 282693 309214 282699
rect 309266 282693 309278 282699
rect 309330 282693 309342 282699
rect 309394 282693 309406 282699
rect 309150 282687 309458 282693
rect 303882 282239 304190 282245
rect 303934 282233 303946 282239
rect 303998 282233 304010 282239
rect 304062 282233 304074 282239
rect 304126 282233 304138 282239
rect 303944 282187 303946 282233
rect 304126 282187 304128 282233
rect 303882 282177 303888 282187
rect 303944 282177 303968 282187
rect 304024 282177 304048 282187
rect 304104 282177 304128 282187
rect 304184 282177 304190 282187
rect 303882 282175 304190 282177
rect 303934 282153 303946 282175
rect 303998 282153 304010 282175
rect 304062 282153 304074 282175
rect 304126 282153 304138 282175
rect 303944 282123 303946 282153
rect 304126 282123 304128 282153
rect 303882 282111 303888 282123
rect 303944 282111 303968 282123
rect 304024 282111 304048 282123
rect 304104 282111 304128 282123
rect 304184 282111 304190 282123
rect 303944 282097 303946 282111
rect 304126 282097 304128 282111
rect 303934 282073 303946 282097
rect 303998 282073 304010 282097
rect 304062 282073 304074 282097
rect 304126 282073 304138 282097
rect 310882 282192 311190 282198
rect 310934 282178 310946 282192
rect 310998 282178 311010 282192
rect 311062 282178 311074 282192
rect 311126 282178 311138 282192
rect 310944 282140 310946 282178
rect 311126 282140 311128 282178
rect 310882 282128 310888 282140
rect 310944 282128 310968 282140
rect 311024 282128 311048 282140
rect 311104 282128 311128 282140
rect 311184 282128 311190 282140
rect 310944 282122 310946 282128
rect 311126 282122 311128 282128
rect 310934 282098 310946 282122
rect 310998 282098 311010 282122
rect 311062 282098 311074 282122
rect 311126 282098 311138 282122
rect 299112 282056 299164 282062
rect 299112 281998 299164 282004
rect 302424 282056 302476 282062
rect 302424 281998 302476 282004
rect 303944 282059 303946 282073
rect 304126 282059 304128 282073
rect 308956 282087 309008 282093
rect 303882 282047 303888 282059
rect 303944 282047 303968 282059
rect 304024 282047 304048 282059
rect 304104 282047 304128 282059
rect 304184 282047 304190 282059
rect 303944 282017 303946 282047
rect 304126 282017 304128 282047
rect 299124 281353 299152 281998
rect 299110 281344 299166 281353
rect 299110 281279 299166 281288
rect 302436 279993 302464 281998
rect 303934 281995 303946 282017
rect 303998 281995 304010 282017
rect 304062 281995 304074 282017
rect 304126 281995 304138 282017
rect 305736 282056 305788 282062
rect 308956 282029 309008 282035
rect 310944 282076 310946 282098
rect 311126 282076 311128 282098
rect 310882 282064 310888 282076
rect 310944 282064 310968 282076
rect 311024 282064 311048 282076
rect 311104 282064 311128 282076
rect 311184 282064 311190 282076
rect 310944 282042 310946 282064
rect 311126 282042 311128 282064
rect 305736 281998 305788 282004
rect 303882 281993 304190 281995
rect 303882 281983 303888 281993
rect 303944 281983 303968 281993
rect 304024 281983 304048 281993
rect 304104 281983 304128 281993
rect 304184 281983 304190 281993
rect 303944 281937 303946 281983
rect 304126 281937 304128 281983
rect 303934 281931 303946 281937
rect 303998 281931 304010 281937
rect 304062 281931 304074 281937
rect 304126 281931 304138 281937
rect 303882 281919 304190 281931
rect 303934 281913 303946 281919
rect 303998 281913 304010 281919
rect 304062 281913 304074 281919
rect 304126 281913 304138 281919
rect 303944 281867 303946 281913
rect 304126 281867 304128 281913
rect 303882 281857 303888 281867
rect 303944 281857 303968 281867
rect 304024 281857 304048 281867
rect 304104 281857 304128 281867
rect 304184 281857 304190 281867
rect 303882 281855 304190 281857
rect 303934 281833 303946 281855
rect 303998 281833 304010 281855
rect 304062 281833 304074 281855
rect 304126 281833 304138 281855
rect 303944 281803 303946 281833
rect 304126 281803 304128 281833
rect 303882 281791 303888 281803
rect 303944 281791 303968 281803
rect 304024 281791 304048 281803
rect 304104 281791 304128 281803
rect 304184 281791 304190 281803
rect 303944 281777 303946 281791
rect 304126 281777 304128 281791
rect 303934 281753 303946 281777
rect 303998 281753 304010 281777
rect 304062 281753 304074 281777
rect 304126 281753 304138 281777
rect 303944 281739 303946 281753
rect 304126 281739 304128 281753
rect 303882 281727 303888 281739
rect 303944 281727 303968 281739
rect 304024 281727 304048 281739
rect 304104 281727 304128 281739
rect 304184 281727 304190 281739
rect 303944 281697 303946 281727
rect 304126 281697 304128 281727
rect 303934 281675 303946 281697
rect 303998 281675 304010 281697
rect 304062 281675 304074 281697
rect 304126 281675 304138 281697
rect 303882 281673 304190 281675
rect 303882 281663 303888 281673
rect 303944 281663 303968 281673
rect 304024 281663 304048 281673
rect 304104 281663 304128 281673
rect 304184 281663 304190 281673
rect 303944 281617 303946 281663
rect 304126 281617 304128 281663
rect 303934 281611 303946 281617
rect 303998 281611 304010 281617
rect 304062 281611 304074 281617
rect 304126 281611 304138 281617
rect 303882 281605 304190 281611
rect 305748 281489 305776 281998
rect 305734 281480 305790 281489
rect 305734 281415 305790 281424
rect 308968 280129 308996 282029
rect 310934 282018 310946 282042
rect 310998 282018 311010 282042
rect 311062 282018 311074 282042
rect 311126 282018 311138 282042
rect 310944 282012 310946 282018
rect 311126 282012 311128 282018
rect 310882 282000 310888 282012
rect 310944 282000 310968 282012
rect 311024 282000 311048 282012
rect 311104 282000 311128 282012
rect 311184 282000 311190 282012
rect 310944 281962 310946 282000
rect 311126 281962 311128 282000
rect 310934 281948 310946 281962
rect 310998 281948 311010 281962
rect 311062 281948 311074 281962
rect 311126 281948 311138 281962
rect 310882 281938 311190 281948
rect 310882 281936 310888 281938
rect 310944 281936 310968 281938
rect 311024 281936 311048 281938
rect 311104 281936 311128 281938
rect 311184 281936 311190 281938
rect 310944 281884 310946 281936
rect 311126 281884 311128 281936
rect 310882 281882 310888 281884
rect 310944 281882 310968 281884
rect 311024 281882 311048 281884
rect 311104 281882 311128 281884
rect 311184 281882 311190 281884
rect 310882 281872 311190 281882
rect 310934 281858 310946 281872
rect 310998 281858 311010 281872
rect 311062 281858 311074 281872
rect 311126 281858 311138 281872
rect 310944 281820 310946 281858
rect 311126 281820 311128 281858
rect 310882 281808 310888 281820
rect 310944 281808 310968 281820
rect 311024 281808 311048 281820
rect 311104 281808 311128 281820
rect 311184 281808 311190 281820
rect 310944 281802 310946 281808
rect 311126 281802 311128 281808
rect 310934 281778 310946 281802
rect 310998 281778 311010 281802
rect 311062 281778 311074 281802
rect 311126 281778 311138 281802
rect 310944 281756 310946 281778
rect 311126 281756 311128 281778
rect 310882 281744 310888 281756
rect 310944 281744 310968 281756
rect 311024 281744 311048 281756
rect 311104 281744 311128 281756
rect 311184 281744 311190 281756
rect 310944 281722 310946 281744
rect 311126 281722 311128 281744
rect 310934 281698 310946 281722
rect 310998 281698 311010 281722
rect 311062 281698 311074 281722
rect 311126 281698 311138 281722
rect 310944 281692 310946 281698
rect 311126 281692 311128 281698
rect 310882 281680 310888 281692
rect 310944 281680 310968 281692
rect 311024 281680 311048 281692
rect 311104 281680 311128 281692
rect 311184 281680 311190 281692
rect 310944 281642 310946 281680
rect 311126 281642 311128 281680
rect 310934 281628 310946 281642
rect 310998 281628 311010 281642
rect 311062 281628 311074 281642
rect 311126 281628 311138 281642
rect 310882 281622 311190 281628
rect 308954 280120 309010 280129
rect 308954 280055 309010 280064
rect 302422 279984 302478 279993
rect 302422 279919 302478 279928
rect 295246 277536 295302 277545
rect 295246 277471 295302 277480
rect 298190 277536 298246 277545
rect 298190 277471 298246 277480
rect 295168 277366 295288 277394
rect 295260 265033 295288 277366
rect 295246 265024 295302 265033
rect 295246 264959 295302 264968
rect 295154 262848 295210 262857
rect 295154 262783 295210 262792
rect 292488 262472 292540 262478
rect 292488 262414 292540 262420
rect 292500 241466 292528 262414
rect 292488 241460 292540 241466
rect 292488 241402 292540 241408
rect 292500 220522 292528 241402
rect 295168 241210 295196 262783
rect 295260 243545 295288 264959
rect 298204 262857 298232 277471
rect 308770 265160 308826 265169
rect 308770 265095 308826 265104
rect 299478 265024 299534 265033
rect 299478 264959 299534 264968
rect 305090 265024 305146 265033
rect 305090 264959 305146 264968
rect 298190 262848 298246 262857
rect 298190 262783 298246 262792
rect 298204 262750 298232 262783
rect 298192 262744 298244 262750
rect 298192 262686 298244 262692
rect 299296 262744 299348 262750
rect 299492 262732 299520 264959
rect 305104 262750 305132 264959
rect 308784 262750 308812 265095
rect 312372 265033 312400 285767
rect 312634 285696 312690 285705
rect 312634 285631 312690 285640
rect 312648 283286 312676 285631
rect 312636 283280 312688 283286
rect 312636 283222 312688 283228
rect 312544 282056 312596 282062
rect 312542 282024 312544 282033
rect 312596 282024 312598 282033
rect 312542 281959 312598 281968
rect 312740 277394 312768 285903
rect 313844 285705 313872 304098
rect 313830 285696 313886 285705
rect 313830 285631 313886 285640
rect 312820 283280 312872 283286
rect 312820 283222 312872 283228
rect 312556 277366 312768 277394
rect 312832 277394 312860 283222
rect 312832 277366 313044 277394
rect 312556 265033 312584 277366
rect 312358 265024 312414 265033
rect 312358 264959 312414 264968
rect 312542 265024 312598 265033
rect 312542 264959 312598 264968
rect 312372 263650 312400 264959
rect 312372 263622 312952 263650
rect 299348 262704 299520 262732
rect 305092 262744 305144 262750
rect 299296 262686 299348 262692
rect 305092 262686 305144 262692
rect 308772 262744 308824 262750
rect 308772 262686 308824 262692
rect 312728 262268 312780 262274
rect 312728 262210 312780 262216
rect 302150 262000 302458 262006
rect 302202 261994 302214 262000
rect 302266 261994 302278 262000
rect 302330 261994 302342 262000
rect 302394 261994 302406 262000
rect 302212 261948 302214 261994
rect 302394 261948 302396 261994
rect 302150 261938 302156 261948
rect 302212 261938 302236 261948
rect 302292 261938 302316 261948
rect 302372 261938 302396 261948
rect 302452 261938 302458 261948
rect 302150 261936 302458 261938
rect 302202 261914 302214 261936
rect 302266 261914 302278 261936
rect 302330 261914 302342 261936
rect 302394 261914 302406 261936
rect 302212 261884 302214 261914
rect 302394 261884 302396 261914
rect 302150 261872 302156 261884
rect 302212 261872 302236 261884
rect 302292 261872 302316 261884
rect 302372 261872 302396 261884
rect 302452 261872 302458 261884
rect 302212 261858 302214 261872
rect 302394 261858 302396 261872
rect 302202 261834 302214 261858
rect 302266 261834 302278 261858
rect 302330 261834 302342 261858
rect 302394 261834 302406 261858
rect 302212 261820 302214 261834
rect 302394 261820 302396 261834
rect 302150 261808 302156 261820
rect 302212 261808 302236 261820
rect 302292 261808 302316 261820
rect 302372 261808 302396 261820
rect 302452 261808 302458 261820
rect 302212 261778 302214 261808
rect 302394 261778 302396 261808
rect 302202 261756 302214 261778
rect 302266 261756 302278 261778
rect 302330 261756 302342 261778
rect 302394 261756 302406 261778
rect 302150 261754 302458 261756
rect 302150 261744 302156 261754
rect 302212 261744 302236 261754
rect 302292 261744 302316 261754
rect 302372 261744 302396 261754
rect 302452 261744 302458 261754
rect 302212 261698 302214 261744
rect 302394 261698 302396 261744
rect 302202 261692 302214 261698
rect 302266 261692 302278 261698
rect 302330 261692 302342 261698
rect 302394 261692 302406 261698
rect 302150 261686 302458 261692
rect 309150 262000 309458 262006
rect 309202 261994 309214 262000
rect 309266 261994 309278 262000
rect 309330 261994 309342 262000
rect 309394 261994 309406 262000
rect 309212 261948 309214 261994
rect 309394 261948 309396 261994
rect 309150 261938 309156 261948
rect 309212 261938 309236 261948
rect 309292 261938 309316 261948
rect 309372 261938 309396 261948
rect 309452 261938 309458 261948
rect 309150 261936 309458 261938
rect 309202 261914 309214 261936
rect 309266 261914 309278 261936
rect 309330 261914 309342 261936
rect 309394 261914 309406 261936
rect 309212 261884 309214 261914
rect 309394 261884 309396 261914
rect 309150 261872 309156 261884
rect 309212 261872 309236 261884
rect 309292 261872 309316 261884
rect 309372 261872 309396 261884
rect 309452 261872 309458 261884
rect 309212 261858 309214 261872
rect 309394 261858 309396 261872
rect 309202 261834 309214 261858
rect 309266 261834 309278 261858
rect 309330 261834 309342 261858
rect 309394 261834 309406 261858
rect 309212 261820 309214 261834
rect 309394 261820 309396 261834
rect 309150 261808 309156 261820
rect 309212 261808 309236 261820
rect 309292 261808 309316 261820
rect 309372 261808 309396 261820
rect 309452 261808 309458 261820
rect 309212 261778 309214 261808
rect 309394 261778 309396 261808
rect 309202 261756 309214 261778
rect 309266 261756 309278 261778
rect 309330 261756 309342 261778
rect 309394 261756 309406 261778
rect 309150 261754 309458 261756
rect 309150 261744 309156 261754
rect 309212 261744 309236 261754
rect 309292 261744 309316 261754
rect 309372 261744 309396 261754
rect 309452 261744 309458 261754
rect 312740 261746 312768 262210
rect 309212 261698 309214 261744
rect 309394 261698 309396 261744
rect 309202 261692 309214 261698
rect 309266 261692 309278 261698
rect 309330 261692 309342 261698
rect 309394 261692 309406 261698
rect 309150 261686 309458 261692
rect 312648 261718 312768 261746
rect 299032 259321 299060 261596
rect 303882 261239 304190 261245
rect 303934 261233 303946 261239
rect 303998 261233 304010 261239
rect 304062 261233 304074 261239
rect 304126 261233 304138 261239
rect 303944 261187 303946 261233
rect 304126 261187 304128 261233
rect 303882 261177 303888 261187
rect 303944 261177 303968 261187
rect 304024 261177 304048 261187
rect 304104 261177 304128 261187
rect 304184 261177 304190 261187
rect 303882 261175 304190 261177
rect 303934 261153 303946 261175
rect 303998 261153 304010 261175
rect 304062 261153 304074 261175
rect 304126 261153 304138 261175
rect 303944 261123 303946 261153
rect 304126 261123 304128 261153
rect 303882 261111 303888 261123
rect 303944 261111 303968 261123
rect 304024 261111 304048 261123
rect 304104 261111 304128 261123
rect 304184 261111 304190 261123
rect 303944 261097 303946 261111
rect 304126 261097 304128 261111
rect 303934 261073 303946 261097
rect 303998 261073 304010 261097
rect 304062 261073 304074 261097
rect 304126 261073 304138 261097
rect 303944 261059 303946 261073
rect 304126 261059 304128 261073
rect 302608 261044 302660 261050
rect 302608 260986 302660 260992
rect 303882 261047 303888 261059
rect 303944 261047 303968 261059
rect 304024 261047 304048 261059
rect 304104 261047 304128 261059
rect 304184 261047 304190 261059
rect 303944 261017 303946 261047
rect 304126 261017 304128 261047
rect 303934 260995 303946 261017
rect 303998 260995 304010 261017
rect 304062 260995 304074 261017
rect 304126 260995 304138 261017
rect 303882 260993 304190 260995
rect 299018 259312 299074 259321
rect 299018 259247 299074 259256
rect 302620 259185 302648 260986
rect 303882 260983 303888 260993
rect 303944 260983 303968 260993
rect 304024 260983 304048 260993
rect 304104 260983 304128 260993
rect 304184 260983 304190 260993
rect 303944 260937 303946 260983
rect 304126 260937 304128 260983
rect 303934 260931 303946 260937
rect 303998 260931 304010 260937
rect 304062 260931 304074 260937
rect 304126 260931 304138 260937
rect 303882 260919 304190 260931
rect 303934 260913 303946 260919
rect 303998 260913 304010 260919
rect 304062 260913 304074 260919
rect 304126 260913 304138 260919
rect 303944 260867 303946 260913
rect 304126 260867 304128 260913
rect 303882 260857 303888 260867
rect 303944 260857 303968 260867
rect 304024 260857 304048 260867
rect 304104 260857 304128 260867
rect 304184 260857 304190 260867
rect 303882 260855 304190 260857
rect 303934 260833 303946 260855
rect 303998 260833 304010 260855
rect 304062 260833 304074 260855
rect 304126 260833 304138 260855
rect 303944 260803 303946 260833
rect 304126 260803 304128 260833
rect 303882 260791 303888 260803
rect 303944 260791 303968 260803
rect 304024 260791 304048 260803
rect 304104 260791 304128 260803
rect 304184 260791 304190 260803
rect 303944 260777 303946 260791
rect 304126 260777 304128 260791
rect 303934 260753 303946 260777
rect 303998 260753 304010 260777
rect 304062 260753 304074 260777
rect 304126 260753 304138 260777
rect 303944 260739 303946 260753
rect 304126 260739 304128 260753
rect 303882 260727 303888 260739
rect 303944 260727 303968 260739
rect 304024 260727 304048 260739
rect 304104 260727 304128 260739
rect 304184 260727 304190 260739
rect 303944 260697 303946 260727
rect 304126 260697 304128 260727
rect 303934 260675 303946 260697
rect 303998 260675 304010 260697
rect 304062 260675 304074 260697
rect 304126 260675 304138 260697
rect 303882 260673 304190 260675
rect 303882 260663 303888 260673
rect 303944 260663 303968 260673
rect 304024 260663 304048 260673
rect 304104 260663 304128 260673
rect 304184 260663 304190 260673
rect 303944 260617 303946 260663
rect 304126 260617 304128 260663
rect 303934 260611 303946 260617
rect 303998 260611 304010 260617
rect 304062 260611 304074 260617
rect 304126 260611 304138 260617
rect 303882 260605 304190 260611
rect 305932 260545 305960 261596
rect 309506 260672 309562 260681
rect 309506 260607 309562 260616
rect 305918 260536 305974 260545
rect 305918 260471 305974 260480
rect 309520 259457 309548 260607
rect 309506 259448 309562 259457
rect 309506 259383 309562 259392
rect 302606 259176 302662 259185
rect 302606 259111 302662 259120
rect 312648 258074 312676 261718
rect 312818 261624 312874 261633
rect 312818 261559 312874 261568
rect 312648 258046 312768 258074
rect 312740 248414 312768 258046
rect 312464 248386 312768 248414
rect 295246 243536 295302 243545
rect 295246 243471 295302 243480
rect 300858 243536 300914 243545
rect 300858 243471 300914 243480
rect 296882 242086 297190 242092
rect 296934 242080 296946 242086
rect 296998 242080 297010 242086
rect 297062 242080 297074 242086
rect 297126 242080 297138 242086
rect 296944 242034 296946 242080
rect 297126 242034 297128 242080
rect 296882 242024 296888 242034
rect 296944 242024 296968 242034
rect 297024 242024 297048 242034
rect 297104 242024 297128 242034
rect 297184 242024 297190 242034
rect 296882 242022 297190 242024
rect 296934 242000 296946 242022
rect 296998 242000 297010 242022
rect 297062 242000 297074 242022
rect 297126 242000 297138 242022
rect 296944 241970 296946 242000
rect 297126 241970 297128 242000
rect 296882 241958 296888 241970
rect 296944 241958 296968 241970
rect 297024 241958 297048 241970
rect 297104 241958 297128 241970
rect 297184 241958 297190 241970
rect 296944 241944 296946 241958
rect 297126 241944 297128 241958
rect 296934 241920 296946 241944
rect 296998 241920 297010 241944
rect 297062 241920 297074 241944
rect 297126 241920 297138 241944
rect 296944 241906 296946 241920
rect 297126 241906 297128 241920
rect 300872 241913 300900 243471
rect 304630 243400 304686 243409
rect 304630 243335 304686 243344
rect 312082 243400 312138 243409
rect 312082 243335 312138 243344
rect 303882 242086 304190 242092
rect 303934 242080 303946 242086
rect 303998 242080 304010 242086
rect 304062 242080 304074 242086
rect 304126 242080 304138 242086
rect 303944 242034 303946 242080
rect 304126 242034 304128 242080
rect 303882 242024 303888 242034
rect 303944 242024 303968 242034
rect 304024 242024 304048 242034
rect 304104 242024 304128 242034
rect 304184 242024 304190 242034
rect 303882 242022 304190 242024
rect 303934 242000 303946 242022
rect 303998 242000 304010 242022
rect 304062 242000 304074 242022
rect 304126 242000 304138 242022
rect 303944 241970 303946 242000
rect 304126 241970 304128 242000
rect 303882 241958 303888 241970
rect 303944 241958 303968 241970
rect 304024 241958 304048 241970
rect 304104 241958 304128 241970
rect 304184 241958 304190 241970
rect 303944 241944 303946 241958
rect 304126 241944 304128 241958
rect 303934 241920 303946 241944
rect 303998 241920 304010 241944
rect 304062 241920 304074 241944
rect 304126 241920 304138 241944
rect 296882 241894 296888 241906
rect 296944 241894 296968 241906
rect 297024 241894 297048 241906
rect 297104 241894 297128 241906
rect 297184 241894 297190 241906
rect 296944 241864 296946 241894
rect 297126 241864 297128 241894
rect 296934 241842 296946 241864
rect 296998 241842 297010 241864
rect 297062 241842 297074 241864
rect 297126 241842 297138 241864
rect 296882 241840 297190 241842
rect 296882 241830 296888 241840
rect 296944 241830 296968 241840
rect 297024 241830 297048 241840
rect 297104 241830 297128 241840
rect 297184 241830 297190 241840
rect 300858 241904 300914 241913
rect 300858 241839 300914 241848
rect 303944 241906 303946 241920
rect 304126 241906 304128 241920
rect 304644 241913 304672 243335
rect 310882 242086 311190 242092
rect 310934 242080 310946 242086
rect 310998 242080 311010 242086
rect 311062 242080 311074 242086
rect 311126 242080 311138 242086
rect 310944 242034 310946 242080
rect 311126 242034 311128 242080
rect 310882 242024 310888 242034
rect 310944 242024 310968 242034
rect 311024 242024 311048 242034
rect 311104 242024 311128 242034
rect 311184 242024 311190 242034
rect 310882 242022 311190 242024
rect 310934 242000 310946 242022
rect 310998 242000 311010 242022
rect 311062 242000 311074 242022
rect 311126 242000 311138 242022
rect 310944 241970 310946 242000
rect 311126 241970 311128 242000
rect 310882 241958 310888 241970
rect 310944 241958 310968 241970
rect 311024 241958 311048 241970
rect 311104 241958 311128 241970
rect 311184 241958 311190 241970
rect 310944 241944 310946 241958
rect 311126 241944 311128 241958
rect 310934 241920 310946 241944
rect 310998 241920 311010 241944
rect 311062 241920 311074 241944
rect 311126 241920 311138 241944
rect 303882 241894 303888 241906
rect 303944 241894 303968 241906
rect 304024 241894 304048 241906
rect 304104 241894 304128 241906
rect 304184 241894 304190 241906
rect 303944 241864 303946 241894
rect 304126 241864 304128 241894
rect 303934 241842 303946 241864
rect 303998 241842 304010 241864
rect 304062 241842 304074 241864
rect 304126 241842 304138 241864
rect 303882 241840 304190 241842
rect 296944 241784 296946 241830
rect 297126 241784 297128 241830
rect 296934 241778 296946 241784
rect 296998 241778 297010 241784
rect 297062 241778 297074 241784
rect 297126 241778 297138 241784
rect 296882 241772 297190 241778
rect 303882 241830 303888 241840
rect 303944 241830 303968 241840
rect 304024 241830 304048 241840
rect 304104 241830 304128 241840
rect 304184 241830 304190 241840
rect 304630 241904 304686 241913
rect 304630 241839 304686 241848
rect 310944 241906 310946 241920
rect 311126 241906 311128 241920
rect 310882 241894 310888 241906
rect 310944 241894 310968 241906
rect 311024 241894 311048 241906
rect 311104 241894 311128 241906
rect 311184 241894 311190 241906
rect 310944 241864 310946 241894
rect 311126 241864 311128 241894
rect 310934 241842 310946 241864
rect 310998 241842 311010 241864
rect 311062 241842 311074 241864
rect 311126 241842 311138 241864
rect 310882 241840 311190 241842
rect 303944 241784 303946 241830
rect 304126 241784 304128 241830
rect 303934 241778 303946 241784
rect 303998 241778 304010 241784
rect 304062 241778 304074 241784
rect 304126 241778 304138 241784
rect 303882 241772 304190 241778
rect 310882 241830 310888 241840
rect 310944 241830 310968 241840
rect 311024 241830 311048 241840
rect 311104 241830 311128 241840
rect 311184 241830 311190 241840
rect 310944 241784 310946 241830
rect 311126 241784 311128 241830
rect 310934 241778 310946 241784
rect 310998 241778 311010 241784
rect 311062 241778 311074 241784
rect 311126 241778 311138 241784
rect 310882 241772 311190 241778
rect 311072 241664 311124 241670
rect 300950 241632 301006 241641
rect 311072 241606 311124 241612
rect 300950 241567 301006 241576
rect 300964 241295 300992 241567
rect 304548 241496 304604 241505
rect 311084 241482 311112 241606
rect 311084 241454 311120 241482
rect 304548 241431 304604 241440
rect 296904 241289 296956 241295
rect 296904 241231 296956 241237
rect 300952 241289 301004 241295
rect 300952 241231 301004 241237
rect 295076 241194 295288 241210
rect 296916 241194 296944 241231
rect 295076 241188 295300 241194
rect 295076 241182 295248 241188
rect 295076 229094 295104 241182
rect 295248 241130 295300 241136
rect 296904 241188 296956 241194
rect 296904 241130 296956 241136
rect 295150 241001 295458 241007
rect 295202 240995 295214 241001
rect 295266 240995 295278 241001
rect 295330 240995 295342 241001
rect 295394 240995 295406 241001
rect 295212 240949 295214 240995
rect 295394 240949 295396 240995
rect 295150 240939 295156 240949
rect 295212 240939 295236 240949
rect 295292 240939 295316 240949
rect 295372 240939 295396 240949
rect 295452 240939 295458 240949
rect 295150 240937 295458 240939
rect 295202 240915 295214 240937
rect 295266 240915 295278 240937
rect 295330 240915 295342 240937
rect 295394 240915 295406 240937
rect 295212 240885 295214 240915
rect 295394 240885 295396 240915
rect 300964 240938 300992 241231
rect 304562 241196 304590 241431
rect 311092 241196 311120 241454
rect 309150 240975 309458 240981
rect 309202 240969 309214 240975
rect 309266 240969 309278 240975
rect 309330 240969 309342 240975
rect 309394 240969 309406 240975
rect 300964 240924 301311 240938
rect 300964 240910 301325 240924
rect 295150 240873 295156 240885
rect 295212 240873 295236 240885
rect 295292 240873 295316 240885
rect 295372 240873 295396 240885
rect 295452 240873 295458 240885
rect 295212 240859 295214 240873
rect 295394 240859 295396 240873
rect 295202 240835 295214 240859
rect 295266 240835 295278 240859
rect 295330 240835 295342 240859
rect 295394 240835 295406 240859
rect 295212 240821 295214 240835
rect 295394 240821 295396 240835
rect 295150 240809 295156 240821
rect 295212 240809 295236 240821
rect 295292 240809 295316 240821
rect 295372 240809 295396 240821
rect 295452 240809 295458 240821
rect 295212 240779 295214 240809
rect 295394 240779 295396 240809
rect 295202 240757 295214 240779
rect 295266 240757 295278 240779
rect 295330 240757 295342 240779
rect 295394 240757 295406 240779
rect 295150 240755 295458 240757
rect 295150 240745 295156 240755
rect 295212 240745 295236 240755
rect 295292 240745 295316 240755
rect 295372 240745 295396 240755
rect 295452 240745 295458 240755
rect 295212 240699 295214 240745
rect 295394 240699 295396 240745
rect 295202 240693 295214 240699
rect 295266 240693 295278 240699
rect 295330 240693 295342 240699
rect 295394 240693 295406 240699
rect 295150 240687 295458 240693
rect 301297 240258 301325 240910
rect 309212 240923 309214 240969
rect 309394 240923 309396 240969
rect 309150 240913 309156 240923
rect 309212 240913 309236 240923
rect 309292 240913 309316 240923
rect 309372 240913 309396 240923
rect 309452 240913 309458 240923
rect 309150 240911 309458 240913
rect 309202 240889 309214 240911
rect 309266 240889 309278 240911
rect 309330 240889 309342 240911
rect 309394 240889 309406 240911
rect 309212 240859 309214 240889
rect 309394 240859 309396 240889
rect 309150 240847 309156 240859
rect 309212 240847 309236 240859
rect 309292 240847 309316 240859
rect 309372 240847 309396 240859
rect 309452 240847 309458 240859
rect 309212 240833 309214 240847
rect 309394 240833 309396 240847
rect 309202 240809 309214 240833
rect 309266 240809 309278 240833
rect 309330 240809 309342 240833
rect 309394 240809 309406 240833
rect 309212 240795 309214 240809
rect 309394 240795 309396 240809
rect 309150 240783 309156 240795
rect 309212 240783 309236 240795
rect 309292 240783 309316 240795
rect 309372 240783 309396 240795
rect 309452 240783 309458 240795
rect 309212 240753 309214 240783
rect 309394 240753 309396 240783
rect 309202 240731 309214 240753
rect 309266 240731 309278 240753
rect 309330 240731 309342 240753
rect 309394 240731 309406 240753
rect 309150 240729 309458 240731
rect 309150 240719 309156 240729
rect 309212 240719 309236 240729
rect 309292 240719 309316 240729
rect 309372 240719 309396 240729
rect 309452 240719 309458 240729
rect 309212 240673 309214 240719
rect 309394 240673 309396 240719
rect 309202 240667 309214 240673
rect 309266 240667 309278 240673
rect 309330 240667 309342 240673
rect 309394 240667 309406 240673
rect 309150 240661 309458 240667
rect 302148 240508 302200 240514
rect 302148 240450 302200 240456
rect 308680 240508 308732 240514
rect 308680 240450 308732 240456
rect 301297 240230 301360 240258
rect 298836 240085 298888 240091
rect 298836 240027 298888 240033
rect 298848 238678 298876 240027
rect 298836 238672 298888 238678
rect 298836 238614 298888 238620
rect 294984 229066 295104 229094
rect 294878 222456 294934 222465
rect 294878 222391 294934 222400
rect 292488 220516 292540 220522
rect 292488 220458 292540 220464
rect 292500 206310 292528 220458
rect 292488 206304 292540 206310
rect 292488 206246 292540 206252
rect 292500 199306 292528 206246
rect 294892 202201 294920 222391
rect 294984 220522 295012 229066
rect 295062 221232 295118 221241
rect 295062 221167 295118 221176
rect 294972 220516 295024 220522
rect 294972 220458 295024 220464
rect 294984 202881 295012 220458
rect 294970 202872 295026 202881
rect 294970 202807 295026 202816
rect 294878 202192 294934 202201
rect 294878 202127 294934 202136
rect 295076 201521 295104 221167
rect 296882 221087 297190 221093
rect 296934 221081 296946 221087
rect 296998 221081 297010 221087
rect 297062 221081 297074 221087
rect 297126 221081 297138 221087
rect 296944 221035 296946 221081
rect 297126 221035 297128 221081
rect 296882 221025 296888 221035
rect 296944 221025 296968 221035
rect 297024 221025 297048 221035
rect 297104 221025 297128 221035
rect 297184 221025 297190 221035
rect 296882 221023 297190 221025
rect 296934 221001 296946 221023
rect 296998 221001 297010 221023
rect 297062 221001 297074 221023
rect 297126 221001 297138 221023
rect 296944 220971 296946 221001
rect 297126 220971 297128 221001
rect 296882 220959 296888 220971
rect 296944 220959 296968 220971
rect 297024 220959 297048 220971
rect 297104 220959 297128 220971
rect 297184 220959 297190 220971
rect 301332 220969 301360 240230
rect 302160 238610 302188 240450
rect 305368 240085 305420 240091
rect 305368 240027 305420 240033
rect 302148 238604 302200 238610
rect 302148 238546 302200 238552
rect 305380 238542 305408 240027
rect 308692 238746 308720 240450
rect 310882 239914 311190 239920
rect 310934 239908 310946 239914
rect 310998 239908 311010 239914
rect 311062 239908 311074 239914
rect 311126 239908 311138 239914
rect 310944 239862 310946 239908
rect 311126 239862 311128 239908
rect 310882 239852 310888 239862
rect 310944 239852 310968 239862
rect 311024 239852 311048 239862
rect 311104 239852 311128 239862
rect 311184 239852 311190 239862
rect 310882 239850 311190 239852
rect 310934 239828 310946 239850
rect 310998 239828 311010 239850
rect 311062 239828 311074 239850
rect 311126 239828 311138 239850
rect 310944 239798 310946 239828
rect 311126 239798 311128 239828
rect 310882 239786 310888 239798
rect 310944 239786 310968 239798
rect 311024 239786 311048 239798
rect 311104 239786 311128 239798
rect 311184 239786 311190 239798
rect 310944 239772 310946 239786
rect 311126 239772 311128 239786
rect 310934 239748 310946 239772
rect 310998 239748 311010 239772
rect 311062 239748 311074 239772
rect 311126 239748 311138 239772
rect 310944 239734 310946 239748
rect 311126 239734 311128 239748
rect 310882 239722 310888 239734
rect 310944 239722 310968 239734
rect 311024 239722 311048 239734
rect 311104 239722 311128 239734
rect 311184 239722 311190 239734
rect 310944 239692 310946 239722
rect 311126 239692 311128 239722
rect 310934 239670 310946 239692
rect 310998 239670 311010 239692
rect 311062 239670 311074 239692
rect 311126 239670 311138 239692
rect 310882 239668 311190 239670
rect 310882 239658 310888 239668
rect 310944 239658 310968 239668
rect 311024 239658 311048 239668
rect 311104 239658 311128 239668
rect 311184 239658 311190 239668
rect 310944 239612 310946 239658
rect 311126 239612 311128 239658
rect 310934 239606 310946 239612
rect 310998 239606 311010 239612
rect 311062 239606 311074 239612
rect 311126 239606 311138 239612
rect 310882 239600 311190 239606
rect 308680 238740 308732 238746
rect 308680 238682 308732 238688
rect 305368 238536 305420 238542
rect 305368 238478 305420 238484
rect 309874 222728 309930 222737
rect 309874 222663 309930 222672
rect 305734 222456 305790 222465
rect 305734 222391 305790 222400
rect 303882 221087 304190 221093
rect 303934 221081 303946 221087
rect 303998 221081 304010 221087
rect 304062 221081 304074 221087
rect 304126 221081 304138 221087
rect 303944 221035 303946 221081
rect 304126 221035 304128 221081
rect 303882 221025 303888 221035
rect 303944 221025 303968 221035
rect 304024 221025 304048 221035
rect 304104 221025 304128 221035
rect 304184 221025 304190 221035
rect 303882 221023 304190 221025
rect 303934 221001 303946 221023
rect 303998 221001 304010 221023
rect 304062 221001 304074 221023
rect 304126 221001 304138 221023
rect 303944 220971 303946 221001
rect 304126 220971 304128 221001
rect 296944 220945 296946 220959
rect 297126 220945 297128 220959
rect 296934 220921 296946 220945
rect 296998 220921 297010 220945
rect 297062 220921 297074 220945
rect 297126 220921 297138 220945
rect 296944 220907 296946 220921
rect 297126 220907 297128 220921
rect 296882 220895 296888 220907
rect 296944 220895 296968 220907
rect 297024 220895 297048 220907
rect 297104 220895 297128 220907
rect 297184 220895 297190 220907
rect 301318 220960 301374 220969
rect 301318 220895 301374 220904
rect 303882 220959 303888 220971
rect 303944 220959 303968 220971
rect 304024 220959 304048 220971
rect 304104 220959 304128 220971
rect 304184 220959 304190 220971
rect 305748 220969 305776 222391
rect 309888 220969 309916 222663
rect 312096 222329 312124 243335
rect 312464 241670 312492 248386
rect 312924 243409 312952 263622
rect 313016 262274 313044 277366
rect 313278 265024 313334 265033
rect 313278 264959 313334 264968
rect 313004 262268 313056 262274
rect 313004 262210 313056 262216
rect 312910 243400 312966 243409
rect 312910 243335 312966 243344
rect 313292 242978 313320 264959
rect 312556 242950 313320 242978
rect 312452 241664 312504 241670
rect 312452 241606 312504 241612
rect 312556 240582 312584 242950
rect 312544 240576 312596 240582
rect 312544 240518 312596 240524
rect 312556 222737 312584 240518
rect 313936 238610 313964 364346
rect 314028 259185 314056 366007
rect 314106 345128 314162 345137
rect 314106 345063 314162 345072
rect 314014 259176 314070 259185
rect 314014 259111 314070 259120
rect 314120 251569 314148 345063
rect 314198 323096 314254 323105
rect 314198 323031 314254 323040
rect 314106 251560 314162 251569
rect 314106 251495 314162 251504
rect 314212 250209 314240 323031
rect 314292 302932 314344 302938
rect 314292 302874 314344 302880
rect 314198 250200 314254 250209
rect 314198 250135 314254 250144
rect 313924 238604 313976 238610
rect 313924 238546 313976 238552
rect 314304 238542 314332 302874
rect 314476 302184 314528 302190
rect 314476 302126 314528 302132
rect 314488 285977 314516 302126
rect 314474 285968 314530 285977
rect 314474 285903 314530 285912
rect 315316 258369 315344 450599
rect 315486 429040 315542 429049
rect 315486 428975 315542 428984
rect 315394 403472 315450 403481
rect 315394 403407 315450 403416
rect 315302 258360 315358 258369
rect 315302 258295 315358 258304
rect 314384 241664 314436 241670
rect 314384 241606 314436 241612
rect 314292 238536 314344 238542
rect 314292 238478 314344 238484
rect 312542 222728 312598 222737
rect 312542 222663 312598 222672
rect 312082 222320 312138 222329
rect 312082 222255 312138 222264
rect 310882 221087 311190 221093
rect 310934 221081 310946 221087
rect 310998 221081 311010 221087
rect 311062 221081 311074 221087
rect 311126 221081 311138 221087
rect 310944 221035 310946 221081
rect 311126 221035 311128 221081
rect 310882 221025 310888 221035
rect 310944 221025 310968 221035
rect 311024 221025 311048 221035
rect 311104 221025 311128 221035
rect 311184 221025 311190 221035
rect 310882 221023 311190 221025
rect 310934 221001 310946 221023
rect 310998 221001 311010 221023
rect 311062 221001 311074 221023
rect 311126 221001 311138 221023
rect 310944 220971 310946 221001
rect 311126 220971 311128 221001
rect 303944 220945 303946 220959
rect 304126 220945 304128 220959
rect 303934 220921 303946 220945
rect 303998 220921 304010 220945
rect 304062 220921 304074 220945
rect 304126 220921 304138 220945
rect 303944 220907 303946 220921
rect 304126 220907 304128 220921
rect 303882 220895 303888 220907
rect 303944 220895 303968 220907
rect 304024 220895 304048 220907
rect 304104 220895 304128 220907
rect 304184 220895 304190 220907
rect 305734 220960 305790 220969
rect 305734 220895 305790 220904
rect 309874 220960 309930 220969
rect 309874 220895 309930 220904
rect 310882 220959 310888 220971
rect 310944 220959 310968 220971
rect 311024 220959 311048 220971
rect 311104 220959 311128 220971
rect 311184 220959 311190 220971
rect 310944 220945 310946 220959
rect 311126 220945 311128 220959
rect 310934 220921 310946 220945
rect 310998 220921 311010 220945
rect 311062 220921 311074 220945
rect 311126 220921 311138 220945
rect 310944 220907 310946 220921
rect 311126 220907 311128 220921
rect 310882 220895 310888 220907
rect 310944 220895 310968 220907
rect 311024 220895 311048 220907
rect 311104 220895 311128 220907
rect 311184 220895 311190 220907
rect 296944 220865 296946 220895
rect 297126 220865 297128 220895
rect 296934 220843 296946 220865
rect 296998 220843 297010 220865
rect 297062 220843 297074 220865
rect 297126 220843 297138 220865
rect 296882 220841 297190 220843
rect 296882 220831 296888 220841
rect 296944 220831 296968 220841
rect 297024 220831 297048 220841
rect 297104 220831 297128 220841
rect 297184 220831 297190 220841
rect 296944 220785 296946 220831
rect 297126 220785 297128 220831
rect 296934 220779 296946 220785
rect 296998 220779 297010 220785
rect 297062 220779 297074 220785
rect 297126 220779 297138 220785
rect 296882 220773 297190 220779
rect 303944 220865 303946 220895
rect 304126 220865 304128 220895
rect 303934 220843 303946 220865
rect 303998 220843 304010 220865
rect 304062 220843 304074 220865
rect 304126 220843 304138 220865
rect 303882 220841 304190 220843
rect 303882 220831 303888 220841
rect 303944 220831 303968 220841
rect 304024 220831 304048 220841
rect 304104 220831 304128 220841
rect 304184 220831 304190 220841
rect 303944 220785 303946 220831
rect 304126 220785 304128 220831
rect 303934 220779 303946 220785
rect 303998 220779 304010 220785
rect 304062 220779 304074 220785
rect 304126 220779 304138 220785
rect 303882 220773 304190 220779
rect 310944 220865 310946 220895
rect 311126 220865 311128 220895
rect 310934 220843 310946 220865
rect 310998 220843 311010 220865
rect 311062 220843 311074 220865
rect 311126 220843 311138 220865
rect 310882 220841 311190 220843
rect 310882 220831 310888 220841
rect 310944 220831 310968 220841
rect 311024 220831 311048 220841
rect 311104 220831 311128 220841
rect 311184 220831 311190 220841
rect 310944 220785 310946 220831
rect 311126 220785 311128 220831
rect 310934 220779 310946 220785
rect 310998 220779 311010 220785
rect 311062 220779 311074 220785
rect 311126 220779 311138 220785
rect 310882 220773 311190 220779
rect 301870 220688 301926 220697
rect 301870 220623 301926 220632
rect 305734 220688 305790 220697
rect 305734 220623 305790 220632
rect 309690 220688 309746 220697
rect 309690 220623 309746 220632
rect 301884 220266 301912 220623
rect 305748 220266 305776 220623
rect 309704 220538 309732 220623
rect 309615 220510 309732 220538
rect 301884 220238 302174 220266
rect 305748 220238 305917 220266
rect 309615 220252 309643 220510
rect 314396 220318 314424 241606
rect 313924 220312 313976 220318
rect 313924 220254 313976 220260
rect 314384 220312 314436 220318
rect 314384 220254 314436 220260
rect 295150 220002 295458 220008
rect 295202 219996 295214 220002
rect 295266 219996 295278 220002
rect 295330 219996 295342 220002
rect 295394 219996 295406 220002
rect 295212 219950 295214 219996
rect 295394 219950 295396 219996
rect 295150 219940 295156 219950
rect 295212 219940 295236 219950
rect 295292 219940 295316 219950
rect 295372 219940 295396 219950
rect 295452 219940 295458 219950
rect 295150 219938 295458 219940
rect 295202 219916 295214 219938
rect 295266 219916 295278 219938
rect 295330 219916 295342 219938
rect 295394 219916 295406 219938
rect 295212 219886 295214 219916
rect 295394 219886 295396 219916
rect 295150 219874 295156 219886
rect 295212 219874 295236 219886
rect 295292 219874 295316 219886
rect 295372 219874 295396 219886
rect 295452 219874 295458 219886
rect 295212 219860 295214 219874
rect 295394 219860 295396 219874
rect 295202 219836 295214 219860
rect 295266 219836 295278 219860
rect 295330 219836 295342 219860
rect 295394 219836 295406 219860
rect 295212 219822 295214 219836
rect 295394 219822 295396 219836
rect 295150 219810 295156 219822
rect 295212 219810 295236 219822
rect 295292 219810 295316 219822
rect 295372 219810 295396 219822
rect 295452 219810 295458 219822
rect 295212 219780 295214 219810
rect 295394 219780 295396 219810
rect 295202 219758 295214 219780
rect 295266 219758 295278 219780
rect 295330 219758 295342 219780
rect 295394 219758 295406 219780
rect 295150 219756 295458 219758
rect 295150 219746 295156 219756
rect 295212 219746 295236 219756
rect 295292 219746 295316 219756
rect 295372 219746 295396 219756
rect 295452 219746 295458 219756
rect 295212 219700 295214 219746
rect 295394 219700 295396 219746
rect 295202 219694 295214 219700
rect 295266 219694 295278 219700
rect 295330 219694 295342 219700
rect 295394 219694 295406 219700
rect 295150 219688 295458 219694
rect 302150 220001 302458 220007
rect 302202 219995 302214 220001
rect 302266 219995 302278 220001
rect 302330 219995 302342 220001
rect 302394 219995 302406 220001
rect 302212 219949 302214 219995
rect 302394 219949 302396 219995
rect 302150 219939 302156 219949
rect 302212 219939 302236 219949
rect 302292 219939 302316 219949
rect 302372 219939 302396 219949
rect 302452 219939 302458 219949
rect 302150 219937 302458 219939
rect 302202 219915 302214 219937
rect 302266 219915 302278 219937
rect 302330 219915 302342 219937
rect 302394 219915 302406 219937
rect 302212 219885 302214 219915
rect 302394 219885 302396 219915
rect 302150 219873 302156 219885
rect 302212 219873 302236 219885
rect 302292 219873 302316 219885
rect 302372 219873 302396 219885
rect 302452 219873 302458 219885
rect 302212 219859 302214 219873
rect 302394 219859 302396 219873
rect 302202 219835 302214 219859
rect 302266 219835 302278 219859
rect 302330 219835 302342 219859
rect 302394 219835 302406 219859
rect 302212 219821 302214 219835
rect 302394 219821 302396 219835
rect 302150 219809 302156 219821
rect 302212 219809 302236 219821
rect 302292 219809 302316 219821
rect 302372 219809 302396 219821
rect 302452 219809 302458 219821
rect 302212 219779 302214 219809
rect 302394 219779 302396 219809
rect 302202 219757 302214 219779
rect 302266 219757 302278 219779
rect 302330 219757 302342 219779
rect 302394 219757 302406 219779
rect 302150 219755 302458 219757
rect 302150 219745 302156 219755
rect 302212 219745 302236 219755
rect 302292 219745 302316 219755
rect 302372 219745 302396 219755
rect 302452 219745 302458 219755
rect 302212 219699 302214 219745
rect 302394 219699 302396 219745
rect 302202 219693 302214 219699
rect 302266 219693 302278 219699
rect 302330 219693 302342 219699
rect 302394 219693 302406 219699
rect 302150 219687 302458 219693
rect 309150 220001 309458 220007
rect 309202 219995 309214 220001
rect 309266 219995 309278 220001
rect 309330 219995 309342 220001
rect 309394 219995 309406 220001
rect 309212 219949 309214 219995
rect 309394 219949 309396 219995
rect 309150 219939 309156 219949
rect 309212 219939 309236 219949
rect 309292 219939 309316 219949
rect 309372 219939 309396 219949
rect 309452 219939 309458 219949
rect 309150 219937 309458 219939
rect 309202 219915 309214 219937
rect 309266 219915 309278 219937
rect 309330 219915 309342 219937
rect 309394 219915 309406 219937
rect 309212 219885 309214 219915
rect 309394 219885 309396 219915
rect 309150 219873 309156 219885
rect 309212 219873 309236 219885
rect 309292 219873 309316 219885
rect 309372 219873 309396 219885
rect 309452 219873 309458 219885
rect 309212 219859 309214 219873
rect 309394 219859 309396 219873
rect 309202 219835 309214 219859
rect 309266 219835 309278 219859
rect 309330 219835 309342 219859
rect 309394 219835 309406 219859
rect 309212 219821 309214 219835
rect 309394 219821 309396 219835
rect 309150 219809 309156 219821
rect 309212 219809 309236 219821
rect 309292 219809 309316 219821
rect 309372 219809 309396 219821
rect 309452 219809 309458 219821
rect 309212 219779 309214 219809
rect 309394 219779 309396 219809
rect 309202 219757 309214 219779
rect 309266 219757 309278 219779
rect 309330 219757 309342 219779
rect 309394 219757 309406 219779
rect 309150 219755 309458 219757
rect 309150 219745 309156 219755
rect 309212 219745 309236 219755
rect 309292 219745 309316 219755
rect 309372 219745 309396 219755
rect 309452 219745 309458 219755
rect 309212 219699 309214 219745
rect 309394 219699 309396 219745
rect 309202 219693 309214 219699
rect 309266 219693 309278 219699
rect 309330 219693 309342 219699
rect 309394 219693 309406 219699
rect 309150 219687 309458 219693
rect 303963 219398 304019 219407
rect 303963 219333 304019 219342
rect 299296 219085 299348 219091
rect 299296 219027 299348 219033
rect 303160 219088 303212 219094
rect 303160 219030 303212 219036
rect 306748 219085 306800 219091
rect 299308 217841 299336 219027
rect 299294 217832 299350 217841
rect 299294 217767 299350 217776
rect 303172 217569 303200 219030
rect 306748 219027 306800 219033
rect 303158 217560 303214 217569
rect 303158 217495 303214 217504
rect 306760 217433 306788 219027
rect 309612 217977 309640 220252
rect 311043 219515 311099 219524
rect 311043 219450 311099 219459
rect 310428 219085 310480 219091
rect 310428 219027 310480 219033
rect 307666 217968 307722 217977
rect 307666 217903 307722 217912
rect 309598 217968 309654 217977
rect 309598 217903 309654 217912
rect 306746 217424 306802 217433
rect 306746 217359 306802 217368
rect 295246 202872 295302 202881
rect 295246 202807 295302 202816
rect 295062 201512 295118 201521
rect 295062 201447 295118 201456
rect 292488 199300 292540 199306
rect 292488 199242 292540 199248
rect 292500 178770 292528 199242
rect 295076 181393 295104 201447
rect 295260 199374 295288 202807
rect 303618 202192 303674 202201
rect 303618 202127 303674 202136
rect 303632 201521 303660 202127
rect 300858 201512 300914 201521
rect 300858 201447 300914 201456
rect 303618 201512 303674 201521
rect 303618 201447 303674 201456
rect 300872 199889 300900 201447
rect 303632 199889 303660 201447
rect 307680 200297 307708 217903
rect 310440 217841 310468 219027
rect 310426 217832 310482 217841
rect 310426 217767 310482 217776
rect 313936 216753 313964 220254
rect 315408 217977 315436 403407
rect 315500 257009 315528 428975
rect 317050 408912 317106 408921
rect 317050 408847 317106 408856
rect 315578 407960 315634 407969
rect 315578 407895 315634 407904
rect 315486 257000 315542 257009
rect 315486 256935 315542 256944
rect 315592 255649 315620 407895
rect 315762 407552 315818 407561
rect 315762 407487 315818 407496
rect 315670 406192 315726 406201
rect 315670 406127 315726 406136
rect 315684 259321 315712 406127
rect 315776 281353 315804 407487
rect 316868 404388 316920 404394
rect 316868 404330 316920 404336
rect 316774 402112 316830 402121
rect 316774 402047 316830 402056
rect 316682 400752 316738 400761
rect 316682 400687 316738 400696
rect 315762 281344 315818 281353
rect 315762 281279 315818 281288
rect 315762 261624 315818 261633
rect 315762 261559 315818 261568
rect 315670 259312 315726 259321
rect 315670 259247 315726 259256
rect 315578 255640 315634 255649
rect 315578 255575 315634 255584
rect 315776 246129 315804 261559
rect 315762 246120 315818 246129
rect 315762 246055 315818 246064
rect 315394 217968 315450 217977
rect 315394 217903 315450 217912
rect 310426 216744 310482 216753
rect 310426 216679 310482 216688
rect 313922 216744 313978 216753
rect 313922 216679 313978 216688
rect 307666 200288 307722 200297
rect 307666 200223 307722 200232
rect 310440 200114 310468 216679
rect 311162 201512 311218 201521
rect 311162 201447 311218 201456
rect 310440 200086 311112 200114
rect 300858 199880 300914 199889
rect 300858 199815 300914 199824
rect 303618 199880 303674 199889
rect 303618 199815 303674 199824
rect 300858 199608 300914 199617
rect 300858 199543 300914 199552
rect 303710 199608 303766 199617
rect 303710 199543 303766 199552
rect 307574 199608 307630 199617
rect 307630 199566 307708 199594
rect 307574 199543 307630 199552
rect 295248 199368 295300 199374
rect 300872 199322 300900 199543
rect 295248 199310 295300 199316
rect 295062 181384 295118 181393
rect 295062 181319 295118 181328
rect 295260 180849 295288 199310
rect 300871 199294 300900 199322
rect 300871 199172 300899 199294
rect 303724 199186 303752 199543
rect 303724 199158 303937 199186
rect 298664 195809 298692 198628
rect 301700 197169 301728 198628
rect 304736 197305 304764 198628
rect 307680 198422 307708 199566
rect 307668 198416 307720 198422
rect 307668 198358 307720 198364
rect 304722 197296 304778 197305
rect 304722 197231 304778 197240
rect 301686 197160 301742 197169
rect 301686 197095 301742 197104
rect 298650 195800 298706 195809
rect 298650 195735 298706 195744
rect 304446 181384 304502 181393
rect 304446 181319 304502 181328
rect 300858 181112 300914 181121
rect 300858 181047 300914 181056
rect 297270 180976 297326 180985
rect 297270 180911 297326 180920
rect 295246 180840 295302 180849
rect 295246 180775 295302 180784
rect 296882 179287 297190 179293
rect 296934 179281 296946 179287
rect 296998 179281 297010 179287
rect 297062 179281 297074 179287
rect 297126 179281 297138 179287
rect 296944 179235 296946 179281
rect 297126 179235 297128 179281
rect 296882 179225 296888 179235
rect 296944 179225 296968 179235
rect 297024 179225 297048 179235
rect 297104 179225 297128 179235
rect 297184 179225 297190 179235
rect 296882 179223 297190 179225
rect 296934 179201 296946 179223
rect 296998 179201 297010 179223
rect 297062 179201 297074 179223
rect 297126 179201 297138 179223
rect 296944 179171 296946 179201
rect 297126 179171 297128 179201
rect 296882 179159 296888 179171
rect 296944 179159 296968 179171
rect 297024 179159 297048 179171
rect 297104 179159 297128 179171
rect 297184 179159 297190 179171
rect 296944 179145 296946 179159
rect 297126 179145 297128 179159
rect 296934 179121 296946 179145
rect 296998 179121 297010 179145
rect 297062 179121 297074 179145
rect 297126 179121 297138 179145
rect 296944 179107 296946 179121
rect 297126 179107 297128 179121
rect 296882 179095 296888 179107
rect 296944 179095 296968 179107
rect 297024 179095 297048 179107
rect 297104 179095 297128 179107
rect 297184 179095 297190 179107
rect 296944 179065 296946 179095
rect 297126 179065 297128 179095
rect 297284 179081 297312 180911
rect 300872 179081 300900 181047
rect 303882 179287 304190 179293
rect 303934 179281 303946 179287
rect 303998 179281 304010 179287
rect 304062 179281 304074 179287
rect 304126 179281 304138 179287
rect 303944 179235 303946 179281
rect 304126 179235 304128 179281
rect 303882 179225 303888 179235
rect 303944 179225 303968 179235
rect 304024 179225 304048 179235
rect 304104 179225 304128 179235
rect 304184 179225 304190 179235
rect 303882 179223 304190 179225
rect 303934 179201 303946 179223
rect 303998 179201 304010 179223
rect 304062 179201 304074 179223
rect 304126 179201 304138 179223
rect 303944 179171 303946 179201
rect 304126 179171 304128 179201
rect 303882 179159 303888 179171
rect 303944 179159 303968 179171
rect 304024 179159 304048 179171
rect 304104 179159 304128 179171
rect 304184 179159 304190 179171
rect 303944 179145 303946 179159
rect 304126 179145 304128 179159
rect 303934 179121 303946 179145
rect 303998 179121 304010 179145
rect 304062 179121 304074 179145
rect 304126 179121 304138 179145
rect 303944 179107 303946 179121
rect 304126 179107 304128 179121
rect 303882 179095 303888 179107
rect 303944 179095 303968 179107
rect 304024 179095 304048 179107
rect 304104 179095 304128 179107
rect 304184 179095 304190 179107
rect 296934 179043 296946 179065
rect 296998 179043 297010 179065
rect 297062 179043 297074 179065
rect 297126 179043 297138 179065
rect 296882 179041 297190 179043
rect 296882 179031 296888 179041
rect 296944 179031 296968 179041
rect 297024 179031 297048 179041
rect 297104 179031 297128 179041
rect 297184 179031 297190 179041
rect 296944 178985 296946 179031
rect 297126 178985 297128 179031
rect 297270 179072 297326 179081
rect 297270 179007 297326 179016
rect 300858 179072 300914 179081
rect 300858 179007 300914 179016
rect 303944 179065 303946 179095
rect 304126 179065 304128 179095
rect 304460 179081 304488 181319
rect 307680 179489 307708 198358
rect 307772 195945 307800 198628
rect 311084 198490 311112 200086
rect 311072 198484 311124 198490
rect 311072 198426 311124 198432
rect 307758 195936 307814 195945
rect 307758 195871 307814 195880
rect 311176 181393 311204 201447
rect 311256 198484 311308 198490
rect 311256 198426 311308 198432
rect 311162 181384 311218 181393
rect 311162 181319 311218 181328
rect 311162 180976 311218 180985
rect 311162 180911 311218 180920
rect 307666 179480 307722 179489
rect 307666 179415 307722 179424
rect 310892 179287 310948 179293
rect 310892 179281 310894 179287
rect 310946 179281 310948 179287
rect 310892 179223 310948 179225
rect 310892 179201 310894 179223
rect 310946 179201 310948 179223
rect 310892 179121 310894 179145
rect 310946 179121 310948 179145
rect 303934 179043 303946 179065
rect 303998 179043 304010 179065
rect 304062 179043 304074 179065
rect 304126 179043 304138 179065
rect 303882 179041 304190 179043
rect 303882 179031 303888 179041
rect 303944 179031 303968 179041
rect 304024 179031 304048 179041
rect 304104 179031 304128 179041
rect 304184 179031 304190 179041
rect 296934 178979 296946 178985
rect 296998 178979 297010 178985
rect 297062 178979 297074 178985
rect 297126 178979 297138 178985
rect 296882 178973 297190 178979
rect 303944 178985 303946 179031
rect 304126 178985 304128 179031
rect 304446 179072 304502 179081
rect 304446 179007 304502 179016
rect 310892 179043 310894 179065
rect 310946 179043 310948 179065
rect 310892 179041 310948 179043
rect 303934 178979 303946 178985
rect 303998 178979 304010 178985
rect 304062 178979 304074 178985
rect 304126 178979 304138 178985
rect 303882 178973 304190 178979
rect 310892 178979 310894 178985
rect 310946 178979 310948 178985
rect 310892 178973 310948 178979
rect 297270 178800 297326 178809
rect 292488 178764 292540 178770
rect 297270 178735 297326 178744
rect 300857 178800 300913 178809
rect 300857 178735 300913 178744
rect 303909 178800 303965 178809
rect 307114 178800 307170 178809
rect 303909 178735 303965 178744
rect 306975 178758 307114 178786
rect 292488 178706 292540 178712
rect 297284 178496 297312 178735
rect 300871 178500 300899 178735
rect 303923 178500 303951 178735
rect 306975 178500 307003 178758
rect 307114 178735 307170 178744
rect 297272 178490 297324 178496
rect 297272 178432 297324 178438
rect 295150 178201 295458 178207
rect 295202 178195 295214 178201
rect 295266 178195 295278 178201
rect 295330 178195 295342 178201
rect 295394 178195 295406 178201
rect 295212 178149 295214 178195
rect 295394 178149 295396 178195
rect 295150 178139 295156 178149
rect 295212 178139 295236 178149
rect 295292 178139 295316 178149
rect 295372 178139 295396 178149
rect 295452 178139 295458 178149
rect 295150 178137 295458 178139
rect 295202 178115 295214 178137
rect 295266 178115 295278 178137
rect 295330 178115 295342 178137
rect 295394 178115 295406 178137
rect 295212 178085 295214 178115
rect 295394 178085 295396 178115
rect 295150 178073 295156 178085
rect 295212 178073 295236 178085
rect 295292 178073 295316 178085
rect 295372 178073 295396 178085
rect 295452 178073 295458 178085
rect 295212 178059 295214 178073
rect 295394 178059 295396 178073
rect 295202 178035 295214 178059
rect 295266 178035 295278 178059
rect 295330 178035 295342 178059
rect 295394 178035 295406 178059
rect 295212 178021 295214 178035
rect 295394 178021 295396 178035
rect 295150 178009 295156 178021
rect 295212 178009 295236 178021
rect 295292 178009 295316 178021
rect 295372 178009 295396 178021
rect 295452 178009 295458 178021
rect 295212 177979 295214 178009
rect 295394 177979 295396 178009
rect 295202 177957 295214 177979
rect 295266 177957 295278 177979
rect 295330 177957 295342 177979
rect 295394 177957 295406 177979
rect 295150 177955 295458 177957
rect 295150 177945 295156 177955
rect 295212 177945 295236 177955
rect 295292 177945 295316 177955
rect 295372 177945 295396 177955
rect 295452 177945 295458 177955
rect 295212 177899 295214 177945
rect 295394 177899 295396 177945
rect 295202 177893 295214 177899
rect 295266 177893 295278 177899
rect 295330 177893 295342 177899
rect 295394 177893 295406 177899
rect 295150 177887 295458 177893
rect 302150 178185 302458 178191
rect 302202 178179 302214 178185
rect 302266 178179 302278 178185
rect 302330 178179 302342 178185
rect 302394 178179 302406 178185
rect 302212 178133 302214 178179
rect 302394 178133 302396 178179
rect 302150 178123 302156 178133
rect 302212 178123 302236 178133
rect 302292 178123 302316 178133
rect 302372 178123 302396 178133
rect 302452 178123 302458 178133
rect 302150 178121 302458 178123
rect 302202 178099 302214 178121
rect 302266 178099 302278 178121
rect 302330 178099 302342 178121
rect 302394 178099 302406 178121
rect 302212 178069 302214 178099
rect 302394 178069 302396 178099
rect 302150 178057 302156 178069
rect 302212 178057 302236 178069
rect 302292 178057 302316 178069
rect 302372 178057 302396 178069
rect 302452 178057 302458 178069
rect 302212 178043 302214 178057
rect 302394 178043 302396 178057
rect 302202 178019 302214 178043
rect 302266 178019 302278 178043
rect 302330 178019 302342 178043
rect 302394 178019 302406 178043
rect 302212 178005 302214 178019
rect 302394 178005 302396 178019
rect 302150 177993 302156 178005
rect 302212 177993 302236 178005
rect 302292 177993 302316 178005
rect 302372 177993 302396 178005
rect 302452 177993 302458 178005
rect 302212 177963 302214 177993
rect 302394 177963 302396 177993
rect 302202 177941 302214 177963
rect 302266 177941 302278 177963
rect 302330 177941 302342 177963
rect 302394 177941 302406 177963
rect 302150 177939 302458 177941
rect 302150 177929 302156 177939
rect 302212 177929 302236 177939
rect 302292 177929 302316 177939
rect 302372 177929 302396 177939
rect 302452 177929 302458 177939
rect 302212 177883 302214 177929
rect 302394 177883 302396 177929
rect 302202 177877 302214 177883
rect 302266 177877 302278 177883
rect 302330 177877 302342 177883
rect 302394 177877 302406 177883
rect 302150 177871 302458 177877
rect 309150 178185 309458 178191
rect 309202 178179 309214 178185
rect 309266 178179 309278 178185
rect 309330 178179 309342 178185
rect 309394 178179 309406 178185
rect 309212 178133 309214 178179
rect 309394 178133 309396 178179
rect 309150 178123 309156 178133
rect 309212 178123 309236 178133
rect 309292 178123 309316 178133
rect 309372 178123 309396 178133
rect 309452 178123 309458 178133
rect 309150 178121 309458 178123
rect 309202 178099 309214 178121
rect 309266 178099 309278 178121
rect 309330 178099 309342 178121
rect 309394 178099 309406 178121
rect 309212 178069 309214 178099
rect 309394 178069 309396 178099
rect 309150 178057 309156 178069
rect 309212 178057 309236 178069
rect 309292 178057 309316 178069
rect 309372 178057 309396 178069
rect 309452 178057 309458 178069
rect 309212 178043 309214 178057
rect 309394 178043 309396 178057
rect 309202 178019 309214 178043
rect 309266 178019 309278 178043
rect 309330 178019 309342 178043
rect 309394 178019 309406 178043
rect 309212 178005 309214 178019
rect 309394 178005 309396 178019
rect 309150 177993 309156 178005
rect 309212 177993 309236 178005
rect 309292 177993 309316 178005
rect 309372 177993 309396 178005
rect 309452 177993 309458 178005
rect 309212 177963 309214 177993
rect 309394 177963 309396 177993
rect 309202 177941 309214 177963
rect 309266 177941 309278 177963
rect 309330 177941 309342 177963
rect 309394 177941 309406 177963
rect 309150 177939 309458 177941
rect 309150 177929 309156 177939
rect 309212 177929 309236 177939
rect 309292 177929 309316 177939
rect 309372 177929 309396 177939
rect 309452 177929 309458 177939
rect 309212 177883 309214 177929
rect 309394 177883 309396 177929
rect 309202 177877 309214 177883
rect 309266 177877 309278 177883
rect 309330 177877 309342 177883
rect 309394 177877 309406 177883
rect 309150 177871 309458 177877
rect 298664 175137 298692 177820
rect 301700 176497 301728 177820
rect 301686 176488 301742 176497
rect 301686 176423 301742 176432
rect 304736 175273 304764 177820
rect 307772 176633 307800 177820
rect 307758 176624 307814 176633
rect 307758 176559 307814 176568
rect 304722 175264 304778 175273
rect 304722 175199 304778 175208
rect 298650 175128 298706 175137
rect 298650 175063 298706 175072
rect 311176 6633 311204 180911
rect 311268 177682 311296 198426
rect 311256 177676 311308 177682
rect 311256 177618 311308 177624
rect 311532 177676 311584 177682
rect 311532 177618 311584 177624
rect 311544 177313 311572 177618
rect 311530 177304 311586 177313
rect 311530 177239 311586 177248
rect 316696 175137 316724 400687
rect 316788 195809 316816 402047
rect 316880 238678 316908 404330
rect 316958 361992 317014 362001
rect 316958 361927 317014 361936
rect 316868 238672 316920 238678
rect 316868 238614 316920 238620
rect 316972 197169 317000 361927
rect 317064 302025 317092 408847
rect 317142 303512 317198 303521
rect 317142 303447 317198 303456
rect 317050 302016 317106 302025
rect 317050 301951 317106 301960
rect 317050 283384 317106 283393
rect 317050 283319 317106 283328
rect 317064 217841 317092 283319
rect 317156 248849 317184 303447
rect 318076 259729 318104 470999
rect 318154 360632 318210 360641
rect 318154 360567 318210 360576
rect 318062 259720 318118 259729
rect 318062 259655 318118 259664
rect 317142 248840 317198 248849
rect 317142 248775 317198 248784
rect 317050 217832 317106 217841
rect 317050 217767 317106 217776
rect 316958 197160 317014 197169
rect 316958 197095 317014 197104
rect 316774 195800 316830 195809
rect 316774 195735 316830 195744
rect 318168 176497 318196 360567
rect 318260 301073 318288 473991
rect 318352 344321 318380 486639
rect 318338 344312 318394 344321
rect 318338 344247 318394 344256
rect 318430 326088 318486 326097
rect 318430 326023 318486 326032
rect 318338 323368 318394 323377
rect 318338 323303 318394 323312
rect 318246 301064 318302 301073
rect 318246 300999 318302 301008
rect 318352 217433 318380 323303
rect 318444 260545 318472 326023
rect 319456 261089 319484 489631
rect 369122 486568 369178 486577
rect 369122 486503 369178 486512
rect 366362 486432 366418 486441
rect 366362 486367 366418 486376
rect 319534 468752 319590 468761
rect 319534 468687 319590 468696
rect 319548 304201 319576 468687
rect 324962 447944 325018 447953
rect 324962 447879 325018 447888
rect 319718 406328 319774 406337
rect 319718 406263 319774 406272
rect 319732 304337 319760 406263
rect 324976 342961 325004 447879
rect 366376 421161 366404 486367
rect 366454 468616 366510 468625
rect 366454 468551 366510 468560
rect 366362 421152 366418 421161
rect 366362 421087 366418 421096
rect 366468 419801 366496 468551
rect 366454 419792 366510 419801
rect 366454 419727 366510 419736
rect 366454 412992 366510 413001
rect 366454 412927 366510 412936
rect 366362 411632 366418 411641
rect 366362 411567 366418 411576
rect 339406 407960 339462 407969
rect 339406 407895 339462 407904
rect 338762 407824 338818 407833
rect 338762 407759 338818 407768
rect 338776 384985 338804 407759
rect 339420 407017 339448 407895
rect 339406 407008 339462 407017
rect 339406 406943 339462 406952
rect 338762 384976 338818 384985
rect 338762 384911 338818 384920
rect 326342 367432 326398 367441
rect 326342 367367 326398 367376
rect 324962 342952 325018 342961
rect 324962 342887 325018 342896
rect 319718 304328 319774 304337
rect 319718 304263 319774 304272
rect 319534 304192 319590 304201
rect 319534 304127 319590 304136
rect 326356 279993 326384 367367
rect 347042 363352 347098 363361
rect 347042 363287 347098 363296
rect 329102 320648 329158 320657
rect 329102 320583 329158 320592
rect 326342 279984 326398 279993
rect 326342 279919 326398 279928
rect 319442 261080 319498 261089
rect 319442 261015 319498 261024
rect 318430 260536 318486 260545
rect 318430 260471 318486 260480
rect 318338 217424 318394 217433
rect 318338 217359 318394 217368
rect 318154 176488 318210 176497
rect 318154 176423 318210 176432
rect 329116 175273 329144 320583
rect 347056 217569 347084 363287
rect 366376 343505 366404 411567
rect 366468 364177 366496 412927
rect 369136 381041 369164 486503
rect 370502 468480 370558 468489
rect 370502 468415 370558 468424
rect 369122 381032 369178 381041
rect 369122 380967 369178 380976
rect 370516 379681 370544 468415
rect 464342 447808 464398 447817
rect 464342 447743 464398 447752
rect 373262 427272 373318 427281
rect 373262 427207 373318 427216
rect 370502 379672 370558 379681
rect 370502 379607 370558 379616
rect 370502 368792 370558 368801
rect 370502 368727 370558 368736
rect 366454 364168 366510 364177
rect 366454 364103 366510 364112
rect 366362 343496 366418 343505
rect 366362 343431 366418 343440
rect 370516 301889 370544 368727
rect 373276 336977 373304 427207
rect 377402 427136 377458 427145
rect 377402 427071 377458 427080
rect 373354 391232 373410 391241
rect 373354 391167 373410 391176
rect 373262 336968 373318 336977
rect 373262 336903 373318 336912
rect 373368 335617 373396 391167
rect 373354 335608 373410 335617
rect 373354 335543 373410 335552
rect 373262 327448 373318 327457
rect 373262 327383 373318 327392
rect 371882 322008 371938 322017
rect 371882 321943 371938 321952
rect 370502 301880 370558 301889
rect 370502 301815 370558 301824
rect 347042 217560 347098 217569
rect 347042 217495 347098 217504
rect 371896 197305 371924 321943
rect 373276 281489 373304 327383
rect 377416 296993 377444 427071
rect 384302 386744 384358 386753
rect 384302 386679 384358 386688
rect 381542 365800 381598 365809
rect 381542 365735 381598 365744
rect 377494 348392 377550 348401
rect 377494 348327 377550 348336
rect 377508 332897 377536 348327
rect 377494 332888 377550 332897
rect 377494 332823 377550 332832
rect 377402 296984 377458 296993
rect 377402 296919 377458 296928
rect 376024 284368 376076 284374
rect 376024 284310 376076 284316
rect 373262 281480 373318 281489
rect 373262 281415 373318 281424
rect 376036 238746 376064 284310
rect 381556 252929 381584 365735
rect 382922 282160 382978 282169
rect 382922 282095 382978 282104
rect 381542 252920 381598 252929
rect 381542 252855 381598 252864
rect 382936 247489 382964 282095
rect 384316 254289 384344 386679
rect 433982 384296 434038 384305
rect 433982 384231 434038 384240
rect 433996 334257 434024 384231
rect 433982 334248 434038 334257
rect 433982 334183 434038 334192
rect 384394 308408 384450 308417
rect 384394 308343 384450 308352
rect 384408 290193 384436 308343
rect 464356 298353 464384 447743
rect 515402 431216 515458 431225
rect 515402 431151 515458 431160
rect 515416 418305 515444 431151
rect 517426 423872 517482 423881
rect 517426 423807 517482 423816
rect 521658 423872 521714 423881
rect 521658 423807 521714 423816
rect 515402 418296 515458 418305
rect 515402 418231 515458 418240
rect 515494 415576 515550 415585
rect 515494 415511 515550 415520
rect 514942 414216 514998 414225
rect 514942 414151 514998 414160
rect 514956 407833 514984 414151
rect 515402 410136 515458 410145
rect 515402 410071 515458 410080
rect 514942 407824 514998 407833
rect 514942 407759 514998 407768
rect 514758 404696 514814 404705
rect 514758 404631 514814 404640
rect 514772 404394 514800 404631
rect 514760 404388 514812 404394
rect 514760 404330 514812 404336
rect 514758 364712 514814 364721
rect 514758 364647 514814 364656
rect 514772 364410 514800 364647
rect 514760 364404 514812 364410
rect 514760 364346 514812 364352
rect 514758 344312 514814 344321
rect 514758 344247 514814 344256
rect 514772 341057 514800 344247
rect 514850 342952 514906 342961
rect 514850 342887 514906 342896
rect 514758 341048 514814 341057
rect 514758 340983 514814 340992
rect 514864 338337 514892 342887
rect 514850 338328 514906 338337
rect 514850 338263 514906 338272
rect 515416 321473 515444 410071
rect 515508 407969 515536 415511
rect 515494 407960 515550 407969
rect 515494 407895 515550 407904
rect 517440 399537 517468 423807
rect 521672 421954 521700 423807
rect 524326 423736 524382 423745
rect 524326 423671 524382 423680
rect 528558 423736 528614 423745
rect 528558 423671 528614 423680
rect 524340 421954 524368 423671
rect 521672 421926 521732 421954
rect 524216 421926 524368 421954
rect 518636 421382 519248 421410
rect 526700 421394 527036 421410
rect 526700 421388 527048 421394
rect 526700 421382 526996 421388
rect 518636 400194 518664 421382
rect 526996 421330 527048 421336
rect 528572 400217 528600 423671
rect 529204 421388 529256 421394
rect 529204 421330 529256 421336
rect 529216 404977 529244 421330
rect 529938 410952 529994 410961
rect 529938 410887 529994 410896
rect 529202 404968 529258 404977
rect 529202 404903 529258 404912
rect 529216 402974 529244 404903
rect 529216 402946 529428 402974
rect 524326 400208 524382 400217
rect 518636 400166 518940 400194
rect 517426 399528 517482 399537
rect 517426 399463 517482 399472
rect 515494 390008 515550 390017
rect 515494 389943 515550 389952
rect 515508 339697 515536 389943
rect 515678 389872 515734 389881
rect 515678 389807 515734 389816
rect 515586 388512 515642 388521
rect 515586 388447 515642 388456
rect 515600 376961 515628 388447
rect 515586 376952 515642 376961
rect 515586 376887 515642 376896
rect 515692 375601 515720 389807
rect 515770 388376 515826 388385
rect 515770 388311 515826 388320
rect 515784 378321 515812 388311
rect 517426 383888 517482 383897
rect 517426 383823 517482 383832
rect 515770 378312 515826 378321
rect 515770 378247 515826 378256
rect 515678 375592 515734 375601
rect 515678 375527 515734 375536
rect 515770 372872 515826 372881
rect 515770 372807 515826 372816
rect 515678 371512 515734 371521
rect 515678 371447 515734 371456
rect 515586 370152 515642 370161
rect 515586 370087 515642 370096
rect 515494 339688 515550 339697
rect 515494 339623 515550 339632
rect 515494 325000 515550 325009
rect 515494 324935 515550 324944
rect 515402 321464 515458 321473
rect 515402 321399 515458 321408
rect 515402 307184 515458 307193
rect 515402 307119 515458 307128
rect 514758 304192 514814 304201
rect 514758 304127 514814 304136
rect 514772 299713 514800 304127
rect 514758 299704 514814 299713
rect 514758 299639 514814 299648
rect 464342 298344 464398 298353
rect 464342 298279 464398 298288
rect 515416 292913 515444 307119
rect 515402 292904 515458 292913
rect 515402 292839 515458 292848
rect 515508 291553 515536 324935
rect 515600 321337 515628 370087
rect 515692 343641 515720 371447
rect 515784 364313 515812 372807
rect 515770 364304 515826 364313
rect 515770 364239 515826 364248
rect 517440 359417 517468 383823
rect 518912 381970 518940 400166
rect 524326 400143 524382 400152
rect 528558 400208 528614 400217
rect 528558 400143 528614 400152
rect 521658 399528 521714 399537
rect 521658 399463 521714 399472
rect 521672 383897 521700 399463
rect 524340 383897 524368 400143
rect 521658 383888 521714 383897
rect 521658 383823 521714 383832
rect 524326 383888 524382 383897
rect 524326 383823 524382 383832
rect 529202 383888 529258 383897
rect 529202 383823 529258 383832
rect 521672 381970 521700 383823
rect 524340 381970 524368 383823
rect 527086 383752 527142 383761
rect 527086 383687 527142 383696
rect 528558 383752 528614 383761
rect 528558 383687 528614 383696
rect 527100 381970 527128 383687
rect 518912 381942 519248 381970
rect 521672 381942 521732 381970
rect 524216 381942 524368 381970
rect 526700 381942 527128 381970
rect 518912 381426 518940 381942
rect 518636 381398 518940 381426
rect 518636 360074 518664 381398
rect 518636 360046 518940 360074
rect 517426 359408 517482 359417
rect 517426 359343 517482 359352
rect 517426 343904 517482 343913
rect 517426 343839 517482 343848
rect 515678 343632 515734 343641
rect 515678 343567 515734 343576
rect 515862 330168 515918 330177
rect 515862 330103 515918 330112
rect 515678 328808 515734 328817
rect 515678 328743 515734 328752
rect 515586 321328 515642 321337
rect 515586 321263 515642 321272
rect 515586 307048 515642 307057
rect 515586 306983 515642 306992
rect 515600 294273 515628 306983
rect 515692 302841 515720 328743
rect 515770 324728 515826 324737
rect 515770 324663 515826 324672
rect 515784 302938 515812 324663
rect 515876 322833 515904 330103
rect 515862 322824 515918 322833
rect 515862 322759 515918 322768
rect 517440 319433 517468 343839
rect 518912 341986 518940 360046
rect 521658 359408 521714 359417
rect 521658 359343 521714 359352
rect 521672 343913 521700 359343
rect 521658 343904 521714 343913
rect 521658 343839 521714 343848
rect 524326 343904 524382 343913
rect 524326 343839 524382 343848
rect 527270 343904 527326 343913
rect 527270 343839 527326 343848
rect 521672 341986 521700 343839
rect 524340 341986 524368 343839
rect 527086 343768 527142 343777
rect 527086 343703 527142 343712
rect 527100 341986 527128 343703
rect 518636 341958 519248 341986
rect 521672 341958 521732 341986
rect 524216 341958 524368 341986
rect 526700 341958 527128 341986
rect 517426 319424 517482 319433
rect 517426 319359 517482 319368
rect 518636 318794 518664 341958
rect 522302 319424 522358 319433
rect 522302 319359 522358 319368
rect 518636 318766 518940 318794
rect 515862 304328 515918 304337
rect 515862 304263 515918 304272
rect 515772 302932 515824 302938
rect 515772 302874 515824 302880
rect 515678 302832 515734 302841
rect 515678 302767 515734 302776
rect 515876 295633 515904 304263
rect 518912 301866 518940 318766
rect 522316 306374 522344 319359
rect 522132 306346 522344 306374
rect 522132 302297 522160 306346
rect 527086 303784 527142 303793
rect 527086 303719 527142 303728
rect 524326 303648 524382 303657
rect 524326 303583 524382 303592
rect 522118 302288 522174 302297
rect 522118 302223 522174 302232
rect 522132 301866 522160 302223
rect 524340 301866 524368 303583
rect 527100 301866 527128 303719
rect 527284 303657 527312 343839
rect 528572 343777 528600 383687
rect 529216 351937 529244 383823
rect 529400 383761 529428 402946
rect 529386 383752 529442 383761
rect 529386 383687 529442 383696
rect 529952 370977 529980 410887
rect 529938 370968 529994 370977
rect 529938 370903 529994 370912
rect 529202 351928 529258 351937
rect 529202 351863 529258 351872
rect 529216 343913 529244 351863
rect 529202 343904 529258 343913
rect 529202 343839 529258 343848
rect 528558 343768 528614 343777
rect 528558 343703 528614 343712
rect 528572 303793 528600 343703
rect 529952 330993 529980 370903
rect 529938 330984 529994 330993
rect 529938 330919 529994 330928
rect 528558 303784 528614 303793
rect 528558 303719 528614 303728
rect 527270 303648 527326 303657
rect 527270 303583 527326 303592
rect 518636 301838 519248 301866
rect 521732 301838 522160 301866
rect 524216 301838 524368 301866
rect 526700 301838 527128 301866
rect 515862 295624 515918 295633
rect 515862 295559 515918 295568
rect 515586 294264 515642 294273
rect 515586 294199 515642 294208
rect 515494 291544 515550 291553
rect 515494 291479 515550 291488
rect 384394 290184 384450 290193
rect 384394 290119 384450 290128
rect 515678 287464 515734 287473
rect 515678 287399 515734 287408
rect 515586 286104 515642 286113
rect 515586 286039 515642 286048
rect 514758 284744 514814 284753
rect 514758 284679 514814 284688
rect 514772 284374 514800 284679
rect 514760 284368 514812 284374
rect 514760 284310 514812 284316
rect 515494 282024 515550 282033
rect 515494 281959 515550 281968
rect 515402 280664 515458 280673
rect 515402 280599 515458 280608
rect 384302 254280 384358 254289
rect 384302 254215 384358 254224
rect 382922 247480 382978 247489
rect 382922 247415 382978 247424
rect 514758 244760 514814 244769
rect 514758 244695 514814 244704
rect 402242 240680 402298 240689
rect 402242 240615 402298 240624
rect 376024 238740 376076 238746
rect 376024 238682 376076 238688
rect 371882 197296 371938 197305
rect 371882 197231 371938 197240
rect 371882 181384 371938 181393
rect 371882 181319 371938 181328
rect 342902 181112 342958 181121
rect 342902 181047 342958 181056
rect 329102 175264 329158 175273
rect 329102 175199 329158 175208
rect 316682 175128 316738 175137
rect 316682 175063 316738 175072
rect 342916 46345 342944 181047
rect 371896 86193 371924 181319
rect 402256 176905 402284 240615
rect 514772 240106 514800 244695
rect 514760 240100 514812 240106
rect 514760 240042 514812 240048
rect 402242 176896 402298 176905
rect 402242 176831 402298 176840
rect 515416 176633 515444 280599
rect 515508 195945 515536 281959
rect 515600 259457 515628 286039
rect 515692 280129 515720 287399
rect 515678 280120 515734 280129
rect 515678 280055 515734 280064
rect 518636 278905 518664 301838
rect 518622 278896 518678 278905
rect 518622 278831 518678 278840
rect 519542 278896 519598 278905
rect 519542 278831 519598 278840
rect 519556 267734 519584 278831
rect 519556 267706 519676 267734
rect 519648 263673 519676 267706
rect 527086 264888 527142 264897
rect 527086 264823 527142 264832
rect 524326 264616 524382 264625
rect 524326 264551 524382 264560
rect 522118 264480 522174 264489
rect 522118 264415 522174 264424
rect 519634 263664 519690 263673
rect 519634 263599 519690 263608
rect 519648 261882 519676 263599
rect 522132 261882 522160 264415
rect 524340 261882 524368 264551
rect 527100 261882 527128 264823
rect 527284 264625 527312 303583
rect 528572 264897 528600 303719
rect 528650 302288 528706 302297
rect 528650 302223 528706 302232
rect 528558 264888 528614 264897
rect 528558 264823 528614 264832
rect 527270 264616 527326 264625
rect 527270 264551 527326 264560
rect 528664 264489 528692 302223
rect 529952 291009 529980 330919
rect 580170 302288 580226 302297
rect 580170 302223 580226 302232
rect 580184 298761 580212 302223
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 529938 291000 529994 291009
rect 529938 290935 529994 290944
rect 528650 264480 528706 264489
rect 528650 264415 528706 264424
rect 527822 263664 527878 263673
rect 527822 263599 527878 263608
rect 519248 261854 519676 261882
rect 521732 261854 522160 261882
rect 524216 261854 524368 261882
rect 526700 261854 527128 261882
rect 515586 259448 515642 259457
rect 515586 259383 515642 259392
rect 527836 245585 527864 263599
rect 529952 251025 529980 290935
rect 529938 251016 529994 251025
rect 529938 250951 529994 250960
rect 530582 251016 530638 251025
rect 530582 250951 530638 250960
rect 527822 245576 527878 245585
rect 527822 245511 527878 245520
rect 515678 243400 515734 243409
rect 515678 243335 515734 243344
rect 515586 242040 515642 242049
rect 515586 241975 515642 241984
rect 515600 197713 515628 241975
rect 515692 218657 515720 243335
rect 515678 218648 515734 218657
rect 515678 218583 515734 218592
rect 515586 197704 515642 197713
rect 515586 197639 515642 197648
rect 515494 195936 515550 195945
rect 515494 195871 515550 195880
rect 515402 176624 515458 176633
rect 515402 176559 515458 176568
rect 371882 86184 371938 86193
rect 371882 86119 371938 86128
rect 342902 46336 342958 46345
rect 342902 46271 342958 46280
rect 530596 19825 530624 250951
rect 580172 206304 580224 206310
rect 580172 206246 580224 206252
rect 580184 205737 580212 206246
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580262 179480 580318 179489
rect 580262 179415 580318 179424
rect 580276 126041 580304 179415
rect 580354 177304 580410 177313
rect 580354 177239 580410 177248
rect 580368 165889 580396 177239
rect 580354 165880 580410 165889
rect 580354 165815 580410 165824
rect 580262 126032 580318 126041
rect 580262 125967 580318 125976
rect 530582 19816 530638 19825
rect 530582 19751 530638 19760
rect 311162 6624 311218 6633
rect 311162 6559 311218 6568
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
<< via2 >>
rect 304446 492768 304502 492824
rect 311990 492768 312046 492824
rect 295062 491816 295118 491872
rect 293866 474000 293922 474056
rect 296888 491604 296934 491650
rect 296934 491604 296944 491650
rect 296968 491604 296998 491650
rect 296998 491604 297010 491650
rect 297010 491604 297024 491650
rect 297048 491604 297062 491650
rect 297062 491604 297074 491650
rect 297074 491604 297104 491650
rect 297128 491604 297138 491650
rect 297138 491604 297184 491650
rect 296888 491594 296944 491604
rect 296968 491594 297024 491604
rect 297048 491594 297104 491604
rect 297128 491594 297184 491604
rect 296888 491540 296934 491570
rect 296934 491540 296944 491570
rect 296968 491540 296998 491570
rect 296998 491540 297010 491570
rect 297010 491540 297024 491570
rect 297048 491540 297062 491570
rect 297062 491540 297074 491570
rect 297074 491540 297104 491570
rect 297128 491540 297138 491570
rect 297138 491540 297184 491570
rect 296888 491528 296944 491540
rect 296968 491528 297024 491540
rect 297048 491528 297104 491540
rect 297128 491528 297184 491540
rect 296888 491514 296934 491528
rect 296934 491514 296944 491528
rect 296968 491514 296998 491528
rect 296998 491514 297010 491528
rect 297010 491514 297024 491528
rect 297048 491514 297062 491528
rect 297062 491514 297074 491528
rect 297074 491514 297104 491528
rect 297128 491514 297138 491528
rect 297138 491514 297184 491528
rect 296888 491476 296934 491490
rect 296934 491476 296944 491490
rect 296968 491476 296998 491490
rect 296998 491476 297010 491490
rect 297010 491476 297024 491490
rect 297048 491476 297062 491490
rect 297062 491476 297074 491490
rect 297074 491476 297104 491490
rect 297128 491476 297138 491490
rect 297138 491476 297184 491490
rect 296888 491464 296944 491476
rect 296968 491464 297024 491476
rect 297048 491464 297104 491476
rect 297128 491464 297184 491476
rect 296888 491434 296934 491464
rect 296934 491434 296944 491464
rect 296968 491434 296998 491464
rect 296998 491434 297010 491464
rect 297010 491434 297024 491464
rect 297048 491434 297062 491464
rect 297062 491434 297074 491464
rect 297074 491434 297104 491464
rect 297128 491434 297138 491464
rect 297138 491434 297184 491464
rect 296888 491400 296944 491410
rect 296968 491400 297024 491410
rect 297048 491400 297104 491410
rect 297128 491400 297184 491410
rect 296888 491354 296934 491400
rect 296934 491354 296944 491400
rect 296968 491354 296998 491400
rect 296998 491354 297010 491400
rect 297010 491354 297024 491400
rect 297048 491354 297062 491400
rect 297062 491354 297074 491400
rect 297074 491354 297104 491400
rect 297128 491354 297138 491400
rect 297138 491354 297184 491400
rect 303888 491604 303934 491650
rect 303934 491604 303944 491650
rect 303968 491604 303998 491650
rect 303998 491604 304010 491650
rect 304010 491604 304024 491650
rect 304048 491604 304062 491650
rect 304062 491604 304074 491650
rect 304074 491604 304104 491650
rect 304128 491604 304138 491650
rect 304138 491604 304184 491650
rect 303888 491594 303944 491604
rect 303968 491594 304024 491604
rect 304048 491594 304104 491604
rect 304128 491594 304184 491604
rect 303888 491540 303934 491570
rect 303934 491540 303944 491570
rect 303968 491540 303998 491570
rect 303998 491540 304010 491570
rect 304010 491540 304024 491570
rect 304048 491540 304062 491570
rect 304062 491540 304074 491570
rect 304074 491540 304104 491570
rect 304128 491540 304138 491570
rect 304138 491540 304184 491570
rect 303888 491528 303944 491540
rect 303968 491528 304024 491540
rect 304048 491528 304104 491540
rect 304128 491528 304184 491540
rect 303888 491514 303934 491528
rect 303934 491514 303944 491528
rect 303968 491514 303998 491528
rect 303998 491514 304010 491528
rect 304010 491514 304024 491528
rect 304048 491514 304062 491528
rect 304062 491514 304074 491528
rect 304074 491514 304104 491528
rect 304128 491514 304138 491528
rect 304138 491514 304184 491528
rect 303888 491476 303934 491490
rect 303934 491476 303944 491490
rect 303968 491476 303998 491490
rect 303998 491476 304010 491490
rect 304010 491476 304024 491490
rect 304048 491476 304062 491490
rect 304062 491476 304074 491490
rect 304074 491476 304104 491490
rect 304128 491476 304138 491490
rect 304138 491476 304184 491490
rect 303888 491464 303944 491476
rect 303968 491464 304024 491476
rect 304048 491464 304104 491476
rect 304128 491464 304184 491476
rect 310888 491604 310934 491650
rect 310934 491604 310944 491650
rect 310968 491604 310998 491650
rect 310998 491604 311010 491650
rect 311010 491604 311024 491650
rect 311048 491604 311062 491650
rect 311062 491604 311074 491650
rect 311074 491604 311104 491650
rect 311128 491604 311138 491650
rect 311138 491604 311184 491650
rect 310888 491594 310944 491604
rect 310968 491594 311024 491604
rect 311048 491594 311104 491604
rect 311128 491594 311184 491604
rect 310888 491540 310934 491570
rect 310934 491540 310944 491570
rect 310968 491540 310998 491570
rect 310998 491540 311010 491570
rect 311010 491540 311024 491570
rect 311048 491540 311062 491570
rect 311062 491540 311074 491570
rect 311074 491540 311104 491570
rect 311128 491540 311138 491570
rect 311138 491540 311184 491570
rect 310888 491528 310944 491540
rect 310968 491528 311024 491540
rect 311048 491528 311104 491540
rect 311128 491528 311184 491540
rect 310888 491514 310934 491528
rect 310934 491514 310944 491528
rect 310968 491514 310998 491528
rect 310998 491514 311010 491528
rect 311010 491514 311024 491528
rect 311048 491514 311062 491528
rect 311062 491514 311074 491528
rect 311074 491514 311104 491528
rect 311128 491514 311138 491528
rect 311138 491514 311184 491528
rect 310888 491476 310934 491490
rect 310934 491476 310944 491490
rect 310968 491476 310998 491490
rect 310998 491476 311010 491490
rect 311010 491476 311024 491490
rect 311048 491476 311062 491490
rect 311062 491476 311074 491490
rect 311074 491476 311104 491490
rect 311128 491476 311138 491490
rect 311138 491476 311184 491490
rect 303888 491434 303934 491464
rect 303934 491434 303944 491464
rect 303968 491434 303998 491464
rect 303998 491434 304010 491464
rect 304010 491434 304024 491464
rect 304048 491434 304062 491464
rect 304062 491434 304074 491464
rect 304074 491434 304104 491464
rect 304128 491434 304138 491464
rect 304138 491434 304184 491464
rect 303888 491400 303944 491410
rect 303968 491400 304024 491410
rect 304048 491400 304104 491410
rect 304128 491400 304184 491410
rect 303888 491354 303934 491400
rect 303934 491354 303944 491400
rect 303968 491354 303998 491400
rect 303998 491354 304010 491400
rect 304010 491354 304024 491400
rect 304048 491354 304062 491400
rect 304062 491354 304074 491400
rect 304074 491354 304104 491400
rect 304128 491354 304138 491400
rect 304138 491354 304184 491400
rect 304446 491408 304502 491464
rect 310888 491464 310944 491476
rect 310968 491464 311024 491476
rect 311048 491464 311104 491476
rect 311128 491464 311184 491476
rect 310888 491434 310934 491464
rect 310934 491434 310944 491464
rect 310968 491434 310998 491464
rect 310998 491434 311010 491464
rect 311010 491434 311024 491464
rect 311048 491434 311062 491464
rect 311062 491434 311074 491464
rect 311074 491434 311104 491464
rect 311128 491434 311138 491464
rect 311138 491434 311184 491464
rect 310888 491400 310944 491410
rect 310968 491400 311024 491410
rect 311048 491400 311104 491410
rect 311128 491400 311184 491410
rect 310888 491354 310934 491400
rect 310934 491354 310944 491400
rect 310968 491354 310998 491400
rect 310998 491354 311010 491400
rect 311010 491354 311024 491400
rect 311048 491354 311062 491400
rect 311062 491354 311074 491400
rect 311074 491354 311104 491400
rect 311128 491354 311138 491400
rect 311138 491354 311184 491400
rect 300858 491136 300914 491192
rect 304221 491000 304277 491056
rect 295156 490496 295202 490534
rect 295202 490496 295212 490534
rect 295236 490496 295266 490534
rect 295266 490496 295278 490534
rect 295278 490496 295292 490534
rect 295316 490496 295330 490534
rect 295330 490496 295342 490534
rect 295342 490496 295372 490534
rect 295396 490496 295406 490534
rect 295406 490496 295452 490534
rect 295156 490484 295212 490496
rect 295236 490484 295292 490496
rect 295316 490484 295372 490496
rect 295396 490484 295452 490496
rect 295156 490478 295202 490484
rect 295202 490478 295212 490484
rect 295236 490478 295266 490484
rect 295266 490478 295278 490484
rect 295278 490478 295292 490484
rect 295316 490478 295330 490484
rect 295330 490478 295342 490484
rect 295342 490478 295372 490484
rect 295396 490478 295406 490484
rect 295406 490478 295452 490484
rect 295156 490432 295202 490454
rect 295202 490432 295212 490454
rect 295236 490432 295266 490454
rect 295266 490432 295278 490454
rect 295278 490432 295292 490454
rect 295316 490432 295330 490454
rect 295330 490432 295342 490454
rect 295342 490432 295372 490454
rect 295396 490432 295406 490454
rect 295406 490432 295452 490454
rect 295156 490420 295212 490432
rect 295236 490420 295292 490432
rect 295316 490420 295372 490432
rect 295396 490420 295452 490432
rect 295156 490398 295202 490420
rect 295202 490398 295212 490420
rect 295236 490398 295266 490420
rect 295266 490398 295278 490420
rect 295278 490398 295292 490420
rect 295316 490398 295330 490420
rect 295330 490398 295342 490420
rect 295342 490398 295372 490420
rect 295396 490398 295406 490420
rect 295406 490398 295452 490420
rect 295156 490368 295202 490374
rect 295202 490368 295212 490374
rect 295236 490368 295266 490374
rect 295266 490368 295278 490374
rect 295278 490368 295292 490374
rect 295316 490368 295330 490374
rect 295330 490368 295342 490374
rect 295342 490368 295372 490374
rect 295396 490368 295406 490374
rect 295406 490368 295452 490374
rect 295156 490356 295212 490368
rect 295236 490356 295292 490368
rect 295316 490356 295372 490368
rect 295396 490356 295452 490368
rect 295156 490318 295202 490356
rect 295202 490318 295212 490356
rect 295236 490318 295266 490356
rect 295266 490318 295278 490356
rect 295278 490318 295292 490356
rect 295316 490318 295330 490356
rect 295330 490318 295342 490356
rect 295342 490318 295372 490356
rect 295396 490318 295406 490356
rect 295406 490318 295452 490356
rect 303888 489432 303934 489478
rect 303934 489432 303944 489478
rect 303968 489432 303998 489478
rect 303998 489432 304010 489478
rect 304010 489432 304024 489478
rect 304048 489432 304062 489478
rect 304062 489432 304074 489478
rect 304074 489432 304104 489478
rect 304128 489432 304138 489478
rect 304138 489432 304184 489478
rect 303888 489422 303944 489432
rect 303968 489422 304024 489432
rect 304048 489422 304104 489432
rect 304128 489422 304184 489432
rect 303888 489368 303934 489398
rect 303934 489368 303944 489398
rect 303968 489368 303998 489398
rect 303998 489368 304010 489398
rect 304010 489368 304024 489398
rect 304048 489368 304062 489398
rect 304062 489368 304074 489398
rect 304074 489368 304104 489398
rect 304128 489368 304138 489398
rect 304138 489368 304184 489398
rect 303888 489356 303944 489368
rect 303968 489356 304024 489368
rect 304048 489356 304104 489368
rect 304128 489356 304184 489368
rect 303888 489342 303934 489356
rect 303934 489342 303944 489356
rect 303968 489342 303998 489356
rect 303998 489342 304010 489356
rect 304010 489342 304024 489356
rect 304048 489342 304062 489356
rect 304062 489342 304074 489356
rect 304074 489342 304104 489356
rect 304128 489342 304138 489356
rect 304138 489342 304184 489356
rect 303888 489304 303934 489318
rect 303934 489304 303944 489318
rect 303968 489304 303998 489318
rect 303998 489304 304010 489318
rect 304010 489304 304024 489318
rect 304048 489304 304062 489318
rect 304062 489304 304074 489318
rect 304074 489304 304104 489318
rect 304128 489304 304138 489318
rect 304138 489304 304184 489318
rect 303888 489292 303944 489304
rect 303968 489292 304024 489304
rect 304048 489292 304104 489304
rect 304128 489292 304184 489304
rect 303888 489262 303934 489292
rect 303934 489262 303944 489292
rect 303968 489262 303998 489292
rect 303998 489262 304010 489292
rect 304010 489262 304024 489292
rect 304048 489262 304062 489292
rect 304062 489262 304074 489292
rect 304074 489262 304104 489292
rect 304128 489262 304138 489292
rect 304138 489262 304184 489292
rect 303888 489228 303944 489238
rect 303968 489228 304024 489238
rect 304048 489228 304104 489238
rect 304128 489228 304184 489238
rect 303888 489182 303934 489228
rect 303934 489182 303944 489228
rect 303968 489182 303998 489228
rect 303998 489182 304010 489228
rect 304010 489182 304024 489228
rect 304048 489182 304062 489228
rect 304062 489182 304074 489228
rect 304074 489182 304104 489228
rect 304128 489182 304138 489228
rect 304138 489182 304184 489228
rect 305090 486648 305146 486704
rect 301778 486512 301834 486568
rect 298742 486376 298798 486432
rect 305550 474680 305606 474736
rect 295062 474000 295118 474056
rect 301410 474000 301466 474056
rect 296888 473064 296934 473110
rect 296934 473064 296944 473110
rect 296968 473064 296998 473110
rect 296998 473064 297010 473110
rect 297010 473064 297024 473110
rect 297048 473064 297062 473110
rect 297062 473064 297074 473110
rect 297074 473064 297104 473110
rect 297128 473064 297138 473110
rect 297138 473064 297184 473110
rect 296888 473054 296944 473064
rect 296968 473054 297024 473064
rect 297048 473054 297104 473064
rect 297128 473054 297184 473064
rect 296888 473000 296934 473030
rect 296934 473000 296944 473030
rect 296968 473000 296998 473030
rect 296998 473000 297010 473030
rect 297010 473000 297024 473030
rect 297048 473000 297062 473030
rect 297062 473000 297074 473030
rect 297074 473000 297104 473030
rect 297128 473000 297138 473030
rect 297138 473000 297184 473030
rect 296888 472988 296944 473000
rect 296968 472988 297024 473000
rect 297048 472988 297104 473000
rect 297128 472988 297184 473000
rect 296888 472974 296934 472988
rect 296934 472974 296944 472988
rect 296968 472974 296998 472988
rect 296998 472974 297010 472988
rect 297010 472974 297024 472988
rect 297048 472974 297062 472988
rect 297062 472974 297074 472988
rect 297074 472974 297104 472988
rect 297128 472974 297138 472988
rect 297138 472974 297184 472988
rect 303888 473064 303934 473110
rect 303934 473064 303944 473110
rect 303968 473064 303998 473110
rect 303998 473064 304010 473110
rect 304010 473064 304024 473110
rect 304048 473064 304062 473110
rect 304062 473064 304074 473110
rect 304074 473064 304104 473110
rect 304128 473064 304138 473110
rect 304138 473064 304184 473110
rect 303888 473054 303944 473064
rect 303968 473054 304024 473064
rect 304048 473054 304104 473064
rect 304128 473054 304184 473064
rect 303888 473000 303934 473030
rect 303934 473000 303944 473030
rect 303968 473000 303998 473030
rect 303998 473000 304010 473030
rect 304010 473000 304024 473030
rect 304048 473000 304062 473030
rect 304062 473000 304074 473030
rect 304074 473000 304104 473030
rect 304128 473000 304138 473030
rect 304138 473000 304184 473030
rect 303888 472988 303944 473000
rect 303968 472988 304024 473000
rect 304048 472988 304104 473000
rect 304128 472988 304184 473000
rect 296888 472936 296934 472950
rect 296934 472936 296944 472950
rect 296968 472936 296998 472950
rect 296998 472936 297010 472950
rect 297010 472936 297024 472950
rect 297048 472936 297062 472950
rect 297062 472936 297074 472950
rect 297074 472936 297104 472950
rect 297128 472936 297138 472950
rect 297138 472936 297184 472950
rect 296888 472924 296944 472936
rect 296968 472924 297024 472936
rect 297048 472924 297104 472936
rect 297128 472924 297184 472936
rect 296888 472894 296934 472924
rect 296934 472894 296944 472924
rect 296968 472894 296998 472924
rect 296998 472894 297010 472924
rect 297010 472894 297024 472924
rect 297048 472894 297062 472924
rect 297062 472894 297074 472924
rect 297074 472894 297104 472924
rect 297128 472894 297138 472924
rect 297138 472894 297184 472924
rect 301410 472912 301466 472968
rect 303888 472974 303934 472988
rect 303934 472974 303944 472988
rect 303968 472974 303998 472988
rect 303998 472974 304010 472988
rect 304010 472974 304024 472988
rect 304048 472974 304062 472988
rect 304062 472974 304074 472988
rect 304074 472974 304104 472988
rect 304128 472974 304138 472988
rect 304138 472974 304184 472988
rect 308126 474000 308182 474056
rect 311530 489655 311586 489696
rect 311530 489640 311532 489655
rect 311532 489640 311584 489655
rect 311584 489640 311586 489655
rect 310888 489432 310934 489478
rect 310934 489432 310944 489478
rect 310968 489432 310998 489478
rect 310998 489432 311010 489478
rect 311010 489432 311024 489478
rect 311048 489432 311062 489478
rect 311062 489432 311074 489478
rect 311074 489432 311104 489478
rect 311128 489432 311138 489478
rect 311138 489432 311184 489478
rect 310888 489422 310944 489432
rect 310968 489422 311024 489432
rect 311048 489422 311104 489432
rect 311128 489422 311184 489432
rect 310888 489368 310934 489398
rect 310934 489368 310944 489398
rect 310968 489368 310998 489398
rect 310998 489368 311010 489398
rect 311010 489368 311024 489398
rect 311048 489368 311062 489398
rect 311062 489368 311074 489398
rect 311074 489368 311104 489398
rect 311128 489368 311138 489398
rect 311138 489368 311184 489398
rect 310888 489356 310944 489368
rect 310968 489356 311024 489368
rect 311048 489356 311104 489368
rect 311128 489356 311184 489368
rect 310888 489342 310934 489356
rect 310934 489342 310944 489356
rect 310968 489342 310998 489356
rect 310998 489342 311010 489356
rect 311010 489342 311024 489356
rect 311048 489342 311062 489356
rect 311062 489342 311074 489356
rect 311074 489342 311104 489356
rect 311128 489342 311138 489356
rect 311138 489342 311184 489356
rect 310888 489304 310934 489318
rect 310934 489304 310944 489318
rect 310968 489304 310998 489318
rect 310998 489304 311010 489318
rect 311010 489304 311024 489318
rect 311048 489304 311062 489318
rect 311062 489304 311074 489318
rect 311074 489304 311104 489318
rect 311128 489304 311138 489318
rect 311138 489304 311184 489318
rect 310888 489292 310944 489304
rect 310968 489292 311024 489304
rect 311048 489292 311104 489304
rect 311128 489292 311184 489304
rect 310888 489262 310934 489292
rect 310934 489262 310944 489292
rect 310968 489262 310998 489292
rect 310998 489262 311010 489292
rect 311010 489262 311024 489292
rect 311048 489262 311062 489292
rect 311062 489262 311074 489292
rect 311074 489262 311104 489292
rect 311128 489262 311138 489292
rect 311138 489262 311184 489292
rect 310888 489228 310944 489238
rect 310968 489228 311024 489238
rect 311048 489228 311104 489238
rect 311128 489228 311184 489238
rect 310888 489182 310934 489228
rect 310934 489182 310944 489228
rect 310968 489182 310998 489228
rect 310998 489182 311010 489228
rect 311010 489182 311024 489228
rect 311048 489182 311062 489228
rect 311062 489182 311074 489228
rect 311074 489182 311104 489228
rect 311128 489182 311138 489228
rect 311138 489182 311184 489228
rect 311990 474680 312046 474736
rect 319442 489640 319498 489696
rect 318338 486648 318394 486704
rect 313646 474680 313702 474736
rect 312174 473456 312230 473512
rect 310518 473320 310574 473376
rect 310888 473064 310934 473110
rect 310934 473064 310944 473110
rect 310968 473064 310998 473110
rect 310998 473064 311010 473110
rect 311010 473064 311024 473110
rect 311048 473064 311062 473110
rect 311062 473064 311074 473110
rect 311074 473064 311104 473110
rect 311128 473064 311138 473110
rect 311138 473064 311184 473110
rect 310888 473054 310944 473064
rect 310968 473054 311024 473064
rect 311048 473054 311104 473064
rect 311128 473054 311184 473064
rect 310888 473000 310934 473030
rect 310934 473000 310944 473030
rect 310968 473000 310998 473030
rect 310998 473000 311010 473030
rect 311010 473000 311024 473030
rect 311048 473000 311062 473030
rect 311062 473000 311074 473030
rect 311074 473000 311104 473030
rect 311128 473000 311138 473030
rect 311138 473000 311184 473030
rect 310888 472988 310944 473000
rect 310968 472988 311024 473000
rect 311048 472988 311104 473000
rect 311128 472988 311184 473000
rect 303888 472936 303934 472950
rect 303934 472936 303944 472950
rect 303968 472936 303998 472950
rect 303998 472936 304010 472950
rect 304010 472936 304024 472950
rect 304048 472936 304062 472950
rect 304062 472936 304074 472950
rect 304074 472936 304104 472950
rect 304128 472936 304138 472950
rect 304138 472936 304184 472950
rect 303888 472924 303944 472936
rect 303968 472924 304024 472936
rect 304048 472924 304104 472936
rect 304128 472924 304184 472936
rect 296888 472860 296944 472870
rect 296968 472860 297024 472870
rect 297048 472860 297104 472870
rect 297128 472860 297184 472870
rect 296888 472814 296934 472860
rect 296934 472814 296944 472860
rect 296968 472814 296998 472860
rect 296998 472814 297010 472860
rect 297010 472814 297024 472860
rect 297048 472814 297062 472860
rect 297062 472814 297074 472860
rect 297074 472814 297104 472860
rect 297128 472814 297138 472860
rect 297138 472814 297184 472860
rect 303888 472894 303934 472924
rect 303934 472894 303944 472924
rect 303968 472894 303998 472924
rect 303998 472894 304010 472924
rect 304010 472894 304024 472924
rect 304048 472894 304062 472924
rect 304062 472894 304074 472924
rect 304074 472894 304104 472924
rect 304128 472894 304138 472924
rect 304138 472894 304184 472924
rect 305550 472912 305606 472968
rect 310888 472974 310934 472988
rect 310934 472974 310944 472988
rect 310968 472974 310998 472988
rect 310998 472974 311010 472988
rect 311010 472974 311024 472988
rect 311048 472974 311062 472988
rect 311062 472974 311074 472988
rect 311074 472974 311104 472988
rect 311128 472974 311138 472988
rect 311138 472974 311184 472988
rect 310888 472936 310934 472950
rect 310934 472936 310944 472950
rect 310968 472936 310998 472950
rect 310998 472936 311010 472950
rect 311010 472936 311024 472950
rect 311048 472936 311062 472950
rect 311062 472936 311074 472950
rect 311074 472936 311104 472950
rect 311128 472936 311138 472950
rect 311138 472936 311184 472950
rect 310888 472924 310944 472936
rect 310968 472924 311024 472936
rect 311048 472924 311104 472936
rect 311128 472924 311184 472936
rect 303888 472860 303944 472870
rect 303968 472860 304024 472870
rect 304048 472860 304104 472870
rect 304128 472860 304184 472870
rect 303888 472814 303934 472860
rect 303934 472814 303944 472860
rect 303968 472814 303998 472860
rect 303998 472814 304010 472860
rect 304010 472814 304024 472860
rect 304048 472814 304062 472860
rect 304062 472814 304074 472860
rect 304074 472814 304104 472860
rect 304128 472814 304138 472860
rect 304138 472814 304184 472860
rect 310888 472894 310934 472924
rect 310934 472894 310944 472924
rect 310968 472894 310998 472924
rect 310998 472894 311010 472924
rect 311010 472894 311024 472924
rect 311048 472894 311062 472924
rect 311062 472894 311074 472924
rect 311074 472894 311104 472924
rect 311128 472894 311138 472924
rect 311138 472894 311184 472924
rect 310888 472860 310944 472870
rect 310968 472860 311024 472870
rect 311048 472860 311104 472870
rect 311128 472860 311184 472870
rect 310888 472814 310934 472860
rect 310934 472814 310944 472860
rect 310968 472814 310998 472860
rect 310998 472814 311010 472860
rect 311010 472814 311024 472860
rect 311048 472814 311062 472860
rect 311062 472814 311074 472860
rect 311074 472814 311104 472860
rect 311128 472814 311138 472860
rect 311138 472814 311184 472860
rect 301594 472640 301650 472696
rect 309138 472640 309194 472696
rect 312358 472640 312414 472696
rect 305508 472504 305564 472560
rect 302156 471963 302202 472009
rect 302202 471963 302212 472009
rect 302236 471963 302266 472009
rect 302266 471963 302278 472009
rect 302278 471963 302292 472009
rect 302316 471963 302330 472009
rect 302330 471963 302342 472009
rect 302342 471963 302372 472009
rect 302396 471963 302406 472009
rect 302406 471963 302452 472009
rect 302156 471953 302212 471963
rect 302236 471953 302292 471963
rect 302316 471953 302372 471963
rect 302396 471953 302452 471963
rect 302156 471899 302202 471929
rect 302202 471899 302212 471929
rect 302236 471899 302266 471929
rect 302266 471899 302278 471929
rect 302278 471899 302292 471929
rect 302316 471899 302330 471929
rect 302330 471899 302342 471929
rect 302342 471899 302372 471929
rect 302396 471899 302406 471929
rect 302406 471899 302452 471929
rect 302156 471887 302212 471899
rect 302236 471887 302292 471899
rect 302316 471887 302372 471899
rect 302396 471887 302452 471899
rect 302156 471873 302202 471887
rect 302202 471873 302212 471887
rect 302236 471873 302266 471887
rect 302266 471873 302278 471887
rect 302278 471873 302292 471887
rect 302316 471873 302330 471887
rect 302330 471873 302342 471887
rect 302342 471873 302372 471887
rect 302396 471873 302406 471887
rect 302406 471873 302452 471887
rect 302156 471835 302202 471849
rect 302202 471835 302212 471849
rect 302236 471835 302266 471849
rect 302266 471835 302278 471849
rect 302278 471835 302292 471849
rect 302316 471835 302330 471849
rect 302330 471835 302342 471849
rect 302342 471835 302372 471849
rect 302396 471835 302406 471849
rect 302406 471835 302452 471849
rect 302156 471823 302212 471835
rect 302236 471823 302292 471835
rect 302316 471823 302372 471835
rect 302396 471823 302452 471835
rect 302156 471793 302202 471823
rect 302202 471793 302212 471823
rect 302236 471793 302266 471823
rect 302266 471793 302278 471823
rect 302278 471793 302292 471823
rect 302316 471793 302330 471823
rect 302330 471793 302342 471823
rect 302342 471793 302372 471823
rect 302396 471793 302406 471823
rect 302406 471793 302452 471823
rect 302156 471759 302212 471769
rect 302236 471759 302292 471769
rect 302316 471759 302372 471769
rect 302396 471759 302452 471769
rect 302156 471713 302202 471759
rect 302202 471713 302212 471759
rect 302236 471713 302266 471759
rect 302266 471713 302278 471759
rect 302278 471713 302292 471759
rect 302316 471713 302330 471759
rect 302330 471713 302342 471759
rect 302342 471713 302372 471759
rect 302396 471713 302406 471759
rect 302406 471713 302452 471759
rect 309156 471963 309202 472009
rect 309202 471963 309212 472009
rect 309236 471963 309266 472009
rect 309266 471963 309278 472009
rect 309278 471963 309292 472009
rect 309316 471963 309330 472009
rect 309330 471963 309342 472009
rect 309342 471963 309372 472009
rect 309396 471963 309406 472009
rect 309406 471963 309452 472009
rect 309156 471953 309212 471963
rect 309236 471953 309292 471963
rect 309316 471953 309372 471963
rect 309396 471953 309452 471963
rect 309156 471899 309202 471929
rect 309202 471899 309212 471929
rect 309236 471899 309266 471929
rect 309266 471899 309278 471929
rect 309278 471899 309292 471929
rect 309316 471899 309330 471929
rect 309330 471899 309342 471929
rect 309342 471899 309372 471929
rect 309396 471899 309406 471929
rect 309406 471899 309452 471929
rect 309156 471887 309212 471899
rect 309236 471887 309292 471899
rect 309316 471887 309372 471899
rect 309396 471887 309452 471899
rect 309156 471873 309202 471887
rect 309202 471873 309212 471887
rect 309236 471873 309266 471887
rect 309266 471873 309278 471887
rect 309278 471873 309292 471887
rect 309316 471873 309330 471887
rect 309330 471873 309342 471887
rect 309342 471873 309372 471887
rect 309396 471873 309406 471887
rect 309406 471873 309452 471887
rect 309156 471835 309202 471849
rect 309202 471835 309212 471849
rect 309236 471835 309266 471849
rect 309266 471835 309278 471849
rect 309278 471835 309292 471849
rect 309316 471835 309330 471849
rect 309330 471835 309342 471849
rect 309342 471835 309372 471849
rect 309396 471835 309406 471849
rect 309406 471835 309452 471849
rect 309156 471823 309212 471835
rect 309236 471823 309292 471835
rect 309316 471823 309372 471835
rect 309396 471823 309452 471835
rect 309156 471793 309202 471823
rect 309202 471793 309212 471823
rect 309236 471793 309266 471823
rect 309266 471793 309278 471823
rect 309278 471793 309292 471823
rect 309316 471793 309330 471823
rect 309330 471793 309342 471823
rect 309342 471793 309372 471823
rect 309396 471793 309406 471823
rect 309406 471793 309452 471823
rect 309156 471759 309212 471769
rect 309236 471759 309292 471769
rect 309316 471759 309372 471769
rect 309396 471759 309452 471769
rect 309156 471713 309202 471759
rect 309202 471713 309212 471759
rect 309236 471713 309266 471759
rect 309266 471713 309278 471759
rect 309278 471713 309292 471759
rect 309316 471713 309330 471759
rect 309330 471713 309342 471759
rect 309342 471713 309372 471759
rect 309396 471713 309406 471759
rect 309406 471713 309452 471759
rect 318246 474000 318302 474056
rect 313738 473456 313794 473512
rect 299294 468560 299350 468616
rect 302882 468424 302938 468480
rect 310058 470600 310114 470656
rect 313830 473320 313886 473376
rect 313646 471044 313648 471064
rect 313648 471044 313700 471064
rect 313700 471044 313702 471064
rect 313646 471008 313702 471044
rect 310058 468696 310114 468752
rect 306470 467880 306526 467936
rect 313002 455368 313058 455424
rect 312542 453872 312598 453928
rect 308310 452648 308366 452704
rect 312542 452648 312598 452704
rect 296888 452024 296934 452054
rect 296934 452024 296944 452054
rect 296968 452024 296998 452054
rect 296998 452024 297010 452054
rect 297010 452024 297024 452054
rect 297048 452024 297062 452054
rect 297062 452024 297074 452054
rect 297074 452024 297104 452054
rect 297128 452024 297138 452054
rect 297138 452024 297184 452054
rect 296888 452012 296944 452024
rect 296968 452012 297024 452024
rect 297048 452012 297104 452024
rect 297128 452012 297184 452024
rect 296888 451998 296934 452012
rect 296934 451998 296944 452012
rect 296968 451998 296998 452012
rect 296998 451998 297010 452012
rect 297010 451998 297024 452012
rect 297048 451998 297062 452012
rect 297062 451998 297074 452012
rect 297074 451998 297104 452012
rect 297128 451998 297138 452012
rect 297138 451998 297184 452012
rect 296888 451960 296934 451974
rect 296934 451960 296944 451974
rect 296968 451960 296998 451974
rect 296998 451960 297010 451974
rect 297010 451960 297024 451974
rect 297048 451960 297062 451974
rect 297062 451960 297074 451974
rect 297074 451960 297104 451974
rect 297128 451960 297138 451974
rect 297138 451960 297184 451974
rect 296888 451948 296944 451960
rect 296968 451948 297024 451960
rect 297048 451948 297104 451960
rect 297128 451948 297184 451960
rect 296888 451918 296934 451948
rect 296934 451918 296944 451948
rect 296968 451918 296998 451948
rect 296998 451918 297010 451948
rect 297010 451918 297024 451948
rect 297048 451918 297062 451948
rect 297062 451918 297074 451948
rect 297074 451918 297104 451948
rect 297128 451918 297138 451948
rect 297138 451918 297184 451948
rect 296888 451884 296944 451894
rect 296968 451884 297024 451894
rect 297048 451884 297104 451894
rect 297128 451884 297184 451894
rect 296888 451838 296934 451884
rect 296934 451838 296944 451884
rect 296968 451838 296998 451884
rect 296998 451838 297010 451884
rect 297010 451838 297024 451884
rect 297048 451838 297062 451884
rect 297062 451838 297074 451884
rect 297074 451838 297104 451884
rect 297128 451838 297138 451884
rect 297138 451838 297184 451884
rect 296888 451768 296934 451814
rect 296934 451768 296944 451814
rect 296968 451768 296998 451814
rect 296998 451768 297010 451814
rect 297010 451768 297024 451814
rect 297048 451768 297062 451814
rect 297062 451768 297074 451814
rect 297074 451768 297104 451814
rect 297128 451768 297138 451814
rect 297138 451768 297184 451814
rect 296888 451758 296944 451768
rect 296968 451758 297024 451768
rect 297048 451758 297104 451768
rect 297128 451758 297184 451768
rect 296888 451704 296934 451734
rect 296934 451704 296944 451734
rect 296968 451704 296998 451734
rect 296998 451704 297010 451734
rect 297010 451704 297024 451734
rect 297048 451704 297062 451734
rect 297062 451704 297074 451734
rect 297074 451704 297104 451734
rect 297128 451704 297138 451734
rect 297138 451704 297184 451734
rect 296888 451692 296944 451704
rect 296968 451692 297024 451704
rect 297048 451692 297104 451704
rect 297128 451692 297184 451704
rect 296888 451678 296934 451692
rect 296934 451678 296944 451692
rect 296968 451678 296998 451692
rect 296998 451678 297010 451692
rect 297010 451678 297024 451692
rect 297048 451678 297062 451692
rect 297062 451678 297074 451692
rect 297074 451678 297104 451692
rect 297128 451678 297138 451692
rect 297138 451678 297184 451692
rect 296888 451640 296934 451654
rect 296934 451640 296944 451654
rect 296968 451640 296998 451654
rect 296998 451640 297010 451654
rect 297010 451640 297024 451654
rect 297048 451640 297062 451654
rect 297062 451640 297074 451654
rect 297074 451640 297104 451654
rect 297128 451640 297138 451654
rect 297138 451640 297184 451654
rect 296888 451628 296944 451640
rect 296968 451628 297024 451640
rect 297048 451628 297104 451640
rect 297128 451628 297184 451640
rect 296888 451598 296934 451628
rect 296934 451598 296944 451628
rect 296968 451598 296998 451628
rect 296998 451598 297010 451628
rect 297010 451598 297024 451628
rect 297048 451598 297062 451628
rect 297062 451598 297074 451628
rect 297074 451598 297104 451628
rect 297128 451598 297138 451628
rect 297138 451598 297184 451628
rect 296888 451564 296944 451574
rect 296968 451564 297024 451574
rect 297048 451564 297104 451574
rect 297128 451564 297184 451574
rect 296888 451518 296934 451564
rect 296934 451518 296944 451564
rect 296968 451518 296998 451564
rect 296998 451518 297010 451564
rect 297010 451518 297024 451564
rect 297048 451518 297062 451564
rect 297062 451518 297074 451564
rect 297074 451518 297104 451564
rect 297128 451518 297138 451564
rect 297138 451518 297184 451564
rect 296888 451448 296934 451494
rect 296934 451448 296944 451494
rect 296968 451448 296998 451494
rect 296998 451448 297010 451494
rect 297010 451448 297024 451494
rect 297048 451448 297062 451494
rect 297062 451448 297074 451494
rect 297074 451448 297104 451494
rect 297128 451448 297138 451494
rect 297138 451448 297184 451494
rect 296888 451438 296944 451448
rect 296968 451438 297024 451448
rect 297048 451438 297104 451448
rect 297128 451438 297184 451448
rect 296888 451384 296934 451414
rect 296934 451384 296944 451414
rect 296968 451384 296998 451414
rect 296998 451384 297010 451414
rect 297010 451384 297024 451414
rect 297048 451384 297062 451414
rect 297062 451384 297074 451414
rect 297074 451384 297104 451414
rect 297128 451384 297138 451414
rect 297138 451384 297184 451414
rect 296888 451372 296944 451384
rect 296968 451372 297024 451384
rect 297048 451372 297104 451384
rect 297128 451372 297184 451384
rect 296888 451358 296934 451372
rect 296934 451358 296944 451372
rect 296968 451358 296998 451372
rect 296998 451358 297010 451372
rect 297010 451358 297024 451372
rect 297048 451358 297062 451372
rect 297062 451358 297074 451372
rect 297074 451358 297104 451372
rect 297128 451358 297138 451372
rect 297138 451358 297184 451372
rect 296888 451320 296934 451334
rect 296934 451320 296944 451334
rect 296968 451320 296998 451334
rect 296998 451320 297010 451334
rect 297010 451320 297024 451334
rect 297048 451320 297062 451334
rect 297062 451320 297074 451334
rect 297074 451320 297104 451334
rect 297128 451320 297138 451334
rect 297138 451320 297184 451334
rect 296888 451308 296944 451320
rect 296968 451308 297024 451320
rect 297048 451308 297104 451320
rect 297128 451308 297184 451320
rect 296888 451278 296934 451308
rect 296934 451278 296944 451308
rect 296968 451278 296998 451308
rect 296998 451278 297010 451308
rect 297010 451278 297024 451308
rect 297048 451278 297062 451308
rect 297062 451278 297074 451308
rect 297074 451278 297104 451308
rect 297128 451278 297138 451308
rect 297138 451278 297184 451308
rect 303888 452024 303934 452054
rect 303934 452024 303944 452054
rect 303968 452024 303998 452054
rect 303998 452024 304010 452054
rect 304010 452024 304024 452054
rect 304048 452024 304062 452054
rect 304062 452024 304074 452054
rect 304074 452024 304104 452054
rect 304128 452024 304138 452054
rect 304138 452024 304184 452054
rect 303888 452012 303944 452024
rect 303968 452012 304024 452024
rect 304048 452012 304104 452024
rect 304128 452012 304184 452024
rect 303888 451998 303934 452012
rect 303934 451998 303944 452012
rect 303968 451998 303998 452012
rect 303998 451998 304010 452012
rect 304010 451998 304024 452012
rect 304048 451998 304062 452012
rect 304062 451998 304074 452012
rect 304074 451998 304104 452012
rect 304128 451998 304138 452012
rect 304138 451998 304184 452012
rect 303888 451960 303934 451974
rect 303934 451960 303944 451974
rect 303968 451960 303998 451974
rect 303998 451960 304010 451974
rect 304010 451960 304024 451974
rect 304048 451960 304062 451974
rect 304062 451960 304074 451974
rect 304074 451960 304104 451974
rect 304128 451960 304138 451974
rect 304138 451960 304184 451974
rect 303888 451948 303944 451960
rect 303968 451948 304024 451960
rect 304048 451948 304104 451960
rect 304128 451948 304184 451960
rect 303888 451918 303934 451948
rect 303934 451918 303944 451948
rect 303968 451918 303998 451948
rect 303998 451918 304010 451948
rect 304010 451918 304024 451948
rect 304048 451918 304062 451948
rect 304062 451918 304074 451948
rect 304074 451918 304104 451948
rect 304128 451918 304138 451948
rect 304138 451918 304184 451948
rect 303888 451884 303944 451894
rect 303968 451884 304024 451894
rect 304048 451884 304104 451894
rect 304128 451884 304184 451894
rect 303888 451838 303934 451884
rect 303934 451838 303944 451884
rect 303968 451838 303998 451884
rect 303998 451838 304010 451884
rect 304010 451838 304024 451884
rect 304048 451838 304062 451884
rect 304062 451838 304074 451884
rect 304074 451838 304104 451884
rect 304128 451838 304138 451884
rect 304138 451838 304184 451884
rect 303888 451768 303934 451814
rect 303934 451768 303944 451814
rect 303968 451768 303998 451814
rect 303998 451768 304010 451814
rect 304010 451768 304024 451814
rect 304048 451768 304062 451814
rect 304062 451768 304074 451814
rect 304074 451768 304104 451814
rect 304128 451768 304138 451814
rect 304138 451768 304184 451814
rect 303888 451758 303944 451768
rect 303968 451758 304024 451768
rect 304048 451758 304104 451768
rect 304128 451758 304184 451768
rect 310919 452024 310949 452054
rect 310949 452024 310961 452054
rect 310961 452024 310975 452054
rect 310999 452024 311013 452054
rect 311013 452024 311025 452054
rect 311025 452024 311055 452054
rect 310919 452012 310975 452024
rect 310999 452012 311055 452024
rect 310919 451998 310949 452012
rect 310949 451998 310961 452012
rect 310961 451998 310975 452012
rect 310999 451998 311013 452012
rect 311013 451998 311025 452012
rect 311025 451998 311055 452012
rect 310919 451960 310949 451974
rect 310949 451960 310961 451974
rect 310961 451960 310975 451974
rect 310999 451960 311013 451974
rect 311013 451960 311025 451974
rect 311025 451960 311055 451974
rect 310919 451948 310975 451960
rect 310999 451948 311055 451960
rect 310919 451918 310949 451948
rect 310949 451918 310961 451948
rect 310961 451918 310975 451948
rect 310999 451918 311013 451948
rect 311013 451918 311025 451948
rect 311025 451918 311055 451948
rect 310919 451884 310975 451894
rect 310999 451884 311055 451894
rect 310919 451838 310949 451884
rect 310949 451838 310961 451884
rect 310961 451838 310975 451884
rect 310999 451838 311013 451884
rect 311013 451838 311025 451884
rect 311025 451838 311055 451884
rect 310919 451768 310949 451814
rect 310949 451768 310961 451814
rect 310961 451768 310975 451814
rect 310999 451768 311013 451814
rect 311013 451768 311025 451814
rect 311025 451768 311055 451814
rect 303888 451704 303934 451734
rect 303934 451704 303944 451734
rect 303968 451704 303998 451734
rect 303998 451704 304010 451734
rect 304010 451704 304024 451734
rect 304048 451704 304062 451734
rect 304062 451704 304074 451734
rect 304074 451704 304104 451734
rect 304128 451704 304138 451734
rect 304138 451704 304184 451734
rect 303888 451692 303944 451704
rect 303968 451692 304024 451704
rect 304048 451692 304104 451704
rect 304128 451692 304184 451704
rect 303888 451678 303934 451692
rect 303934 451678 303944 451692
rect 303968 451678 303998 451692
rect 303998 451678 304010 451692
rect 304010 451678 304024 451692
rect 304048 451678 304062 451692
rect 304062 451678 304074 451692
rect 304074 451678 304104 451692
rect 304128 451678 304138 451692
rect 304138 451678 304184 451692
rect 308310 451696 308366 451752
rect 310919 451758 310975 451768
rect 310999 451758 311055 451768
rect 310919 451704 310949 451734
rect 310949 451704 310961 451734
rect 310961 451704 310975 451734
rect 310999 451704 311013 451734
rect 311013 451704 311025 451734
rect 311025 451704 311055 451734
rect 310919 451692 310975 451704
rect 310999 451692 311055 451704
rect 303888 451640 303934 451654
rect 303934 451640 303944 451654
rect 303968 451640 303998 451654
rect 303998 451640 304010 451654
rect 304010 451640 304024 451654
rect 304048 451640 304062 451654
rect 304062 451640 304074 451654
rect 304074 451640 304104 451654
rect 304128 451640 304138 451654
rect 304138 451640 304184 451654
rect 303888 451628 303944 451640
rect 303968 451628 304024 451640
rect 304048 451628 304104 451640
rect 304128 451628 304184 451640
rect 303888 451598 303934 451628
rect 303934 451598 303944 451628
rect 303968 451598 303998 451628
rect 303998 451598 304010 451628
rect 304010 451598 304024 451628
rect 304048 451598 304062 451628
rect 304062 451598 304074 451628
rect 304074 451598 304104 451628
rect 304128 451598 304138 451628
rect 304138 451598 304184 451628
rect 303888 451564 303944 451574
rect 303968 451564 304024 451574
rect 304048 451564 304104 451574
rect 304128 451564 304184 451574
rect 303888 451518 303934 451564
rect 303934 451518 303944 451564
rect 303968 451518 303998 451564
rect 303998 451518 304010 451564
rect 304010 451518 304024 451564
rect 304048 451518 304062 451564
rect 304062 451518 304074 451564
rect 304074 451518 304104 451564
rect 304128 451518 304138 451564
rect 304138 451518 304184 451564
rect 303888 451448 303934 451494
rect 303934 451448 303944 451494
rect 303968 451448 303998 451494
rect 303998 451448 304010 451494
rect 304010 451448 304024 451494
rect 304048 451448 304062 451494
rect 304062 451448 304074 451494
rect 304074 451448 304104 451494
rect 304128 451448 304138 451494
rect 304138 451448 304184 451494
rect 310919 451678 310949 451692
rect 310949 451678 310961 451692
rect 310961 451678 310975 451692
rect 310999 451678 311013 451692
rect 311013 451678 311025 451692
rect 311025 451678 311055 451692
rect 310919 451640 310949 451654
rect 310949 451640 310961 451654
rect 310961 451640 310975 451654
rect 310999 451640 311013 451654
rect 311013 451640 311025 451654
rect 311025 451640 311055 451654
rect 310919 451628 310975 451640
rect 310999 451628 311055 451640
rect 310919 451598 310949 451628
rect 310949 451598 310961 451628
rect 310961 451598 310975 451628
rect 310999 451598 311013 451628
rect 311013 451598 311025 451628
rect 311025 451598 311055 451628
rect 310919 451564 310975 451574
rect 310999 451564 311055 451574
rect 310919 451518 310949 451564
rect 310949 451518 310961 451564
rect 310961 451518 310975 451564
rect 310999 451518 311013 451564
rect 311013 451518 311025 451564
rect 311025 451518 311055 451564
rect 303888 451438 303944 451448
rect 303968 451438 304024 451448
rect 304048 451438 304104 451448
rect 304128 451438 304184 451448
rect 308024 451424 308080 451480
rect 310919 451448 310949 451494
rect 310949 451448 310961 451494
rect 310961 451448 310975 451494
rect 310999 451448 311013 451494
rect 311013 451448 311025 451494
rect 311025 451448 311055 451494
rect 310919 451438 310975 451448
rect 310999 451438 311055 451448
rect 303888 451384 303934 451414
rect 303934 451384 303944 451414
rect 303968 451384 303998 451414
rect 303998 451384 304010 451414
rect 304010 451384 304024 451414
rect 304048 451384 304062 451414
rect 304062 451384 304074 451414
rect 304074 451384 304104 451414
rect 304128 451384 304138 451414
rect 304138 451384 304184 451414
rect 303888 451372 303944 451384
rect 303968 451372 304024 451384
rect 304048 451372 304104 451384
rect 304128 451372 304184 451384
rect 303888 451358 303934 451372
rect 303934 451358 303944 451372
rect 303968 451358 303998 451372
rect 303998 451358 304010 451372
rect 304010 451358 304024 451372
rect 304048 451358 304062 451372
rect 304062 451358 304074 451372
rect 304074 451358 304104 451372
rect 304128 451358 304138 451372
rect 304138 451358 304184 451372
rect 303888 451320 303934 451334
rect 303934 451320 303944 451334
rect 303968 451320 303998 451334
rect 303998 451320 304010 451334
rect 304010 451320 304024 451334
rect 304048 451320 304062 451334
rect 304062 451320 304074 451334
rect 304074 451320 304104 451334
rect 304128 451320 304138 451334
rect 304138 451320 304184 451334
rect 303888 451308 303944 451320
rect 303968 451308 304024 451320
rect 304048 451308 304104 451320
rect 304128 451308 304184 451320
rect 303888 451278 303934 451308
rect 303934 451278 303944 451308
rect 303968 451278 303998 451308
rect 303998 451278 304010 451308
rect 304010 451278 304024 451308
rect 304048 451278 304062 451308
rect 304062 451278 304074 451308
rect 304074 451278 304104 451308
rect 304128 451278 304138 451308
rect 304138 451278 304184 451308
rect 310919 451384 310949 451414
rect 310949 451384 310961 451414
rect 310961 451384 310975 451414
rect 310999 451384 311013 451414
rect 311013 451384 311025 451414
rect 311025 451384 311055 451414
rect 310919 451372 310975 451384
rect 310999 451372 311055 451384
rect 310919 451358 310949 451372
rect 310949 451358 310961 451372
rect 310961 451358 310975 451372
rect 310999 451358 311013 451372
rect 311013 451358 311025 451372
rect 311025 451358 311055 451372
rect 310919 451320 310949 451334
rect 310949 451320 310961 451334
rect 310961 451320 310975 451334
rect 310999 451320 311013 451334
rect 311013 451320 311025 451334
rect 311025 451320 311055 451334
rect 310919 451308 310975 451320
rect 310999 451308 311055 451320
rect 310919 451278 310949 451308
rect 310949 451278 310961 451308
rect 310961 451278 310975 451308
rect 310999 451278 311013 451308
rect 311013 451278 311025 451308
rect 311025 451278 311055 451308
rect 293866 449112 293922 449168
rect 300858 449112 300914 449168
rect 298926 448024 298982 448080
rect 302238 448160 302294 448216
rect 306194 449112 306250 449168
rect 305550 447888 305606 447944
rect 312174 450608 312230 450664
rect 310898 450139 310936 450177
rect 310936 450139 310948 450177
rect 310948 450139 310954 450177
rect 310978 450139 311000 450177
rect 311000 450139 311012 450177
rect 311012 450139 311034 450177
rect 311058 450139 311064 450177
rect 311064 450139 311076 450177
rect 311076 450139 311114 450177
rect 310898 450127 310954 450139
rect 310978 450127 311034 450139
rect 311058 450127 311114 450139
rect 310898 450121 310936 450127
rect 310936 450121 310948 450127
rect 310948 450121 310954 450127
rect 310978 450121 311000 450127
rect 311000 450121 311012 450127
rect 311012 450121 311034 450127
rect 311058 450121 311064 450127
rect 311064 450121 311076 450127
rect 311076 450121 311114 450127
rect 310898 450075 310936 450097
rect 310936 450075 310948 450097
rect 310948 450075 310954 450097
rect 310978 450075 311000 450097
rect 311000 450075 311012 450097
rect 311012 450075 311034 450097
rect 311058 450075 311064 450097
rect 311064 450075 311076 450097
rect 311076 450075 311114 450097
rect 310898 450063 310954 450075
rect 310978 450063 311034 450075
rect 311058 450063 311114 450075
rect 310898 450041 310936 450063
rect 310936 450041 310948 450063
rect 310948 450041 310954 450063
rect 310978 450041 311000 450063
rect 311000 450041 311012 450063
rect 311012 450041 311034 450063
rect 311058 450041 311064 450063
rect 311064 450041 311076 450063
rect 311076 450041 311114 450063
rect 310898 450011 310936 450017
rect 310936 450011 310948 450017
rect 310948 450011 310954 450017
rect 310978 450011 311000 450017
rect 311000 450011 311012 450017
rect 311012 450011 311034 450017
rect 311058 450011 311064 450017
rect 311064 450011 311076 450017
rect 311076 450011 311114 450017
rect 310898 449999 310954 450011
rect 310978 449999 311034 450011
rect 311058 449999 311114 450011
rect 310898 449961 310936 449999
rect 310936 449961 310948 449999
rect 310948 449961 310954 449999
rect 310978 449961 311000 449999
rect 311000 449961 311012 449999
rect 311012 449961 311034 449999
rect 311058 449961 311064 449999
rect 311064 449961 311076 449999
rect 311076 449961 311114 449999
rect 310898 449935 310954 449937
rect 310978 449935 311034 449937
rect 311058 449935 311114 449937
rect 310898 449883 310936 449935
rect 310936 449883 310948 449935
rect 310948 449883 310954 449935
rect 310978 449883 311000 449935
rect 311000 449883 311012 449935
rect 311012 449883 311034 449935
rect 311058 449883 311064 449935
rect 311064 449883 311076 449935
rect 311076 449883 311114 449935
rect 310898 449881 310954 449883
rect 310978 449881 311034 449883
rect 311058 449881 311114 449883
rect 310898 449819 310936 449857
rect 310936 449819 310948 449857
rect 310948 449819 310954 449857
rect 310978 449819 311000 449857
rect 311000 449819 311012 449857
rect 311012 449819 311034 449857
rect 311058 449819 311064 449857
rect 311064 449819 311076 449857
rect 311076 449819 311114 449857
rect 310898 449807 310954 449819
rect 310978 449807 311034 449819
rect 311058 449807 311114 449819
rect 310898 449801 310936 449807
rect 310936 449801 310948 449807
rect 310948 449801 310954 449807
rect 310978 449801 311000 449807
rect 311000 449801 311012 449807
rect 311012 449801 311034 449807
rect 311058 449801 311064 449807
rect 311064 449801 311076 449807
rect 311076 449801 311114 449807
rect 310898 449755 310936 449777
rect 310936 449755 310948 449777
rect 310948 449755 310954 449777
rect 310978 449755 311000 449777
rect 311000 449755 311012 449777
rect 311012 449755 311034 449777
rect 311058 449755 311064 449777
rect 311064 449755 311076 449777
rect 311076 449755 311114 449777
rect 310898 449743 310954 449755
rect 310978 449743 311034 449755
rect 311058 449743 311114 449755
rect 310898 449721 310936 449743
rect 310936 449721 310948 449743
rect 310948 449721 310954 449743
rect 310978 449721 311000 449743
rect 311000 449721 311012 449743
rect 311012 449721 311034 449743
rect 311058 449721 311064 449743
rect 311064 449721 311076 449743
rect 311076 449721 311114 449743
rect 310898 449691 310936 449697
rect 310936 449691 310948 449697
rect 310948 449691 310954 449697
rect 310978 449691 311000 449697
rect 311000 449691 311012 449697
rect 311012 449691 311034 449697
rect 311058 449691 311064 449697
rect 311064 449691 311076 449697
rect 311076 449691 311114 449697
rect 310898 449679 310954 449691
rect 310978 449679 311034 449691
rect 311058 449679 311114 449691
rect 310898 449641 310936 449679
rect 310936 449641 310948 449679
rect 310948 449641 310954 449679
rect 310978 449641 311000 449679
rect 311000 449641 311012 449679
rect 311012 449641 311034 449679
rect 311058 449641 311064 449679
rect 311064 449641 311076 449679
rect 311076 449641 311114 449679
rect 308862 447752 308918 447808
rect 318062 471008 318118 471064
rect 313922 467880 313978 467936
rect 313830 455368 313886 455424
rect 313738 453872 313794 453928
rect 312634 448024 312690 448080
rect 308494 433200 308550 433256
rect 312542 433200 312598 433256
rect 305182 432112 305238 432168
rect 306286 432112 306342 432168
rect 312634 431160 312690 431216
rect 300858 430752 300914 430808
rect 305182 430752 305238 430808
rect 308494 430752 308550 430808
rect 301502 430344 301558 430400
rect 305091 430344 305147 430400
rect 308402 430344 308458 430400
rect 313462 449112 313518 449168
rect 313370 433200 313426 433256
rect 313278 432112 313334 432168
rect 295154 410216 295210 410272
rect 309151 429948 309177 429994
rect 309177 429948 309207 429994
rect 309231 429948 309241 429994
rect 309241 429948 309287 429994
rect 309311 429948 309357 429994
rect 309357 429948 309367 429994
rect 309391 429948 309421 429994
rect 309421 429948 309447 429994
rect 309151 429938 309207 429948
rect 309231 429938 309287 429948
rect 309311 429938 309367 429948
rect 309391 429938 309447 429948
rect 309151 429884 309177 429914
rect 309177 429884 309207 429914
rect 309231 429884 309241 429914
rect 309241 429884 309287 429914
rect 309311 429884 309357 429914
rect 309357 429884 309367 429914
rect 309391 429884 309421 429914
rect 309421 429884 309447 429914
rect 309151 429872 309207 429884
rect 309231 429872 309287 429884
rect 309311 429872 309367 429884
rect 309391 429872 309447 429884
rect 309151 429858 309177 429872
rect 309177 429858 309207 429872
rect 309231 429858 309241 429872
rect 309241 429858 309287 429872
rect 309151 429820 309177 429834
rect 309177 429820 309207 429834
rect 309231 429820 309241 429834
rect 309241 429820 309287 429834
rect 309311 429858 309357 429872
rect 309357 429858 309367 429872
rect 309391 429858 309421 429872
rect 309421 429858 309447 429872
rect 309311 429820 309357 429834
rect 309357 429820 309367 429834
rect 309391 429820 309421 429834
rect 309421 429820 309447 429834
rect 309151 429808 309207 429820
rect 309231 429808 309287 429820
rect 309311 429808 309367 429820
rect 309391 429808 309447 429820
rect 309151 429778 309177 429808
rect 309177 429778 309207 429808
rect 309231 429778 309241 429808
rect 309241 429778 309287 429808
rect 309311 429778 309357 429808
rect 309357 429778 309367 429808
rect 309391 429778 309421 429808
rect 309421 429778 309447 429808
rect 309151 429744 309207 429754
rect 309231 429744 309287 429754
rect 309311 429744 309367 429754
rect 309391 429744 309447 429754
rect 309151 429698 309177 429744
rect 309177 429698 309207 429744
rect 309231 429698 309241 429744
rect 309241 429698 309287 429744
rect 309311 429698 309357 429744
rect 309357 429698 309367 429744
rect 309391 429698 309421 429744
rect 309421 429698 309447 429744
rect 300858 427896 300914 427952
rect 301686 427896 301742 427952
rect 302514 427352 302570 427408
rect 309414 428440 309470 428496
rect 305918 427216 305974 427272
rect 309414 427080 309470 427136
rect 309046 423544 309102 423600
rect 299018 417016 299074 417072
rect 305182 411304 305238 411360
rect 301042 410216 301098 410272
rect 296888 410034 296934 410080
rect 296934 410034 296944 410080
rect 296968 410034 296998 410080
rect 296998 410034 297010 410080
rect 297010 410034 297024 410080
rect 297048 410034 297062 410080
rect 297062 410034 297074 410080
rect 297074 410034 297104 410080
rect 297128 410034 297138 410080
rect 297138 410034 297184 410080
rect 296888 410024 296944 410034
rect 296968 410024 297024 410034
rect 297048 410024 297104 410034
rect 297128 410024 297184 410034
rect 296888 409970 296934 410000
rect 296934 409970 296944 410000
rect 296968 409970 296998 410000
rect 296998 409970 297010 410000
rect 297010 409970 297024 410000
rect 297048 409970 297062 410000
rect 297062 409970 297074 410000
rect 297074 409970 297104 410000
rect 297128 409970 297138 410000
rect 297138 409970 297184 410000
rect 296888 409958 296944 409970
rect 296968 409958 297024 409970
rect 297048 409958 297104 409970
rect 297128 409958 297184 409970
rect 296888 409944 296934 409958
rect 296934 409944 296944 409958
rect 296968 409944 296998 409958
rect 296998 409944 297010 409958
rect 297010 409944 297024 409958
rect 297048 409944 297062 409958
rect 297062 409944 297074 409958
rect 297074 409944 297104 409958
rect 297128 409944 297138 409958
rect 297138 409944 297184 409958
rect 296888 409906 296934 409920
rect 296934 409906 296944 409920
rect 296968 409906 296998 409920
rect 296998 409906 297010 409920
rect 297010 409906 297024 409920
rect 297048 409906 297062 409920
rect 297062 409906 297074 409920
rect 297074 409906 297104 409920
rect 297128 409906 297138 409920
rect 297138 409906 297184 409920
rect 296888 409894 296944 409906
rect 296968 409894 297024 409906
rect 297048 409894 297104 409906
rect 297128 409894 297184 409906
rect 296888 409864 296934 409894
rect 296934 409864 296944 409894
rect 296968 409864 296998 409894
rect 296998 409864 297010 409894
rect 297010 409864 297024 409894
rect 297048 409864 297062 409894
rect 297062 409864 297074 409894
rect 297074 409864 297104 409894
rect 297128 409864 297138 409894
rect 297138 409864 297184 409894
rect 303888 410034 303934 410080
rect 303934 410034 303944 410080
rect 303968 410034 303998 410080
rect 303998 410034 304010 410080
rect 304010 410034 304024 410080
rect 304048 410034 304062 410080
rect 304062 410034 304074 410080
rect 304074 410034 304104 410080
rect 304128 410034 304138 410080
rect 304138 410034 304184 410080
rect 303888 410024 303944 410034
rect 303968 410024 304024 410034
rect 304048 410024 304104 410034
rect 304128 410024 304184 410034
rect 303888 409970 303934 410000
rect 303934 409970 303944 410000
rect 303968 409970 303998 410000
rect 303998 409970 304010 410000
rect 304010 409970 304024 410000
rect 304048 409970 304062 410000
rect 304062 409970 304074 410000
rect 304074 409970 304104 410000
rect 304128 409970 304138 410000
rect 304138 409970 304184 410000
rect 303888 409958 303944 409970
rect 303968 409958 304024 409970
rect 304048 409958 304104 409970
rect 304128 409958 304184 409970
rect 303888 409944 303934 409958
rect 303934 409944 303944 409958
rect 303968 409944 303998 409958
rect 303998 409944 304010 409958
rect 304010 409944 304024 409958
rect 304048 409944 304062 409958
rect 304062 409944 304074 409958
rect 304074 409944 304104 409958
rect 304128 409944 304138 409958
rect 304138 409944 304184 409958
rect 303888 409906 303934 409920
rect 303934 409906 303944 409920
rect 303968 409906 303998 409920
rect 303998 409906 304010 409920
rect 304010 409906 304024 409920
rect 304048 409906 304062 409920
rect 304062 409906 304074 409920
rect 304074 409906 304104 409920
rect 304128 409906 304138 409920
rect 304138 409906 304184 409920
rect 303888 409894 303944 409906
rect 303968 409894 304024 409906
rect 304048 409894 304104 409906
rect 304128 409894 304184 409906
rect 296888 409830 296944 409840
rect 296968 409830 297024 409840
rect 297048 409830 297104 409840
rect 297128 409830 297184 409840
rect 296888 409784 296934 409830
rect 296934 409784 296944 409830
rect 296968 409784 296998 409830
rect 296998 409784 297010 409830
rect 297010 409784 297024 409830
rect 297048 409784 297062 409830
rect 297062 409784 297074 409830
rect 297074 409784 297104 409830
rect 297128 409784 297138 409830
rect 297138 409784 297184 409830
rect 301042 409808 301098 409864
rect 303888 409864 303934 409894
rect 303934 409864 303944 409894
rect 303968 409864 303998 409894
rect 303998 409864 304010 409894
rect 304010 409864 304024 409894
rect 304048 409864 304062 409894
rect 304062 409864 304074 409894
rect 304074 409864 304104 409894
rect 304128 409864 304138 409894
rect 304138 409864 304184 409894
rect 313002 429032 313004 429040
rect 313004 429032 313056 429040
rect 313056 429032 313058 429040
rect 313002 428984 313058 429032
rect 313370 423544 313426 423600
rect 312450 411440 312506 411496
rect 313278 411440 313334 411496
rect 312266 411304 312322 411360
rect 313186 411304 313242 411360
rect 309046 410216 309102 410272
rect 312082 410216 312138 410272
rect 310888 410034 310934 410080
rect 310934 410034 310944 410080
rect 310968 410034 310998 410080
rect 310998 410034 311010 410080
rect 311010 410034 311024 410080
rect 311048 410034 311062 410080
rect 311062 410034 311074 410080
rect 311074 410034 311104 410080
rect 311128 410034 311138 410080
rect 311138 410034 311184 410080
rect 310888 410024 310944 410034
rect 310968 410024 311024 410034
rect 311048 410024 311104 410034
rect 311128 410024 311184 410034
rect 310888 409970 310934 410000
rect 310934 409970 310944 410000
rect 310968 409970 310998 410000
rect 310998 409970 311010 410000
rect 311010 409970 311024 410000
rect 311048 409970 311062 410000
rect 311062 409970 311074 410000
rect 311074 409970 311104 410000
rect 311128 409970 311138 410000
rect 311138 409970 311184 410000
rect 310888 409958 310944 409970
rect 310968 409958 311024 409970
rect 311048 409958 311104 409970
rect 311128 409958 311184 409970
rect 310888 409944 310934 409958
rect 310934 409944 310944 409958
rect 310968 409944 310998 409958
rect 310998 409944 311010 409958
rect 311010 409944 311024 409958
rect 311048 409944 311062 409958
rect 311062 409944 311074 409958
rect 311074 409944 311104 409958
rect 311128 409944 311138 409958
rect 311138 409944 311184 409958
rect 310888 409906 310934 409920
rect 310934 409906 310944 409920
rect 310968 409906 310998 409920
rect 310998 409906 311010 409920
rect 311010 409906 311024 409920
rect 311048 409906 311062 409920
rect 311062 409906 311074 409920
rect 311074 409906 311104 409920
rect 311128 409906 311138 409920
rect 311138 409906 311184 409920
rect 310888 409894 310944 409906
rect 310968 409894 311024 409906
rect 311048 409894 311104 409906
rect 311128 409894 311184 409906
rect 303888 409830 303944 409840
rect 303968 409830 304024 409840
rect 304048 409830 304104 409840
rect 304128 409830 304184 409840
rect 303888 409784 303934 409830
rect 303934 409784 303944 409830
rect 303968 409784 303998 409830
rect 303998 409784 304010 409830
rect 304010 409784 304024 409830
rect 304048 409784 304062 409830
rect 304062 409784 304074 409830
rect 304074 409784 304104 409830
rect 304128 409784 304138 409830
rect 304138 409784 304184 409830
rect 305182 409808 305238 409864
rect 310888 409864 310934 409894
rect 310934 409864 310944 409894
rect 310968 409864 310998 409894
rect 310998 409864 311010 409894
rect 311010 409864 311024 409894
rect 311048 409864 311062 409894
rect 311062 409864 311074 409894
rect 311074 409864 311104 409894
rect 311128 409864 311138 409894
rect 311138 409864 311184 409894
rect 310888 409830 310944 409840
rect 310968 409830 311024 409840
rect 311048 409830 311104 409840
rect 311128 409830 311184 409840
rect 310888 409784 310934 409830
rect 310934 409784 310944 409830
rect 310968 409784 310998 409830
rect 310998 409784 311010 409830
rect 311010 409784 311024 409830
rect 311048 409784 311062 409830
rect 311062 409784 311074 409830
rect 311074 409784 311104 409830
rect 311128 409784 311138 409830
rect 311138 409784 311184 409830
rect 301226 409536 301282 409592
rect 304549 409536 304605 409592
rect 307814 409536 307870 409592
rect 302156 408948 302202 408994
rect 302202 408948 302212 408994
rect 302236 408948 302266 408994
rect 302266 408948 302278 408994
rect 302278 408948 302292 408994
rect 302316 408948 302330 408994
rect 302330 408948 302342 408994
rect 302342 408948 302372 408994
rect 302396 408948 302406 408994
rect 302406 408948 302452 408994
rect 302156 408938 302212 408948
rect 302236 408938 302292 408948
rect 302316 408938 302372 408948
rect 302396 408938 302452 408948
rect 302156 408884 302202 408914
rect 302202 408884 302212 408914
rect 302236 408884 302266 408914
rect 302266 408884 302278 408914
rect 302278 408884 302292 408914
rect 302316 408884 302330 408914
rect 302330 408884 302342 408914
rect 302342 408884 302372 408914
rect 302396 408884 302406 408914
rect 302406 408884 302452 408914
rect 302156 408872 302212 408884
rect 302236 408872 302292 408884
rect 302316 408872 302372 408884
rect 302396 408872 302452 408884
rect 302156 408858 302202 408872
rect 302202 408858 302212 408872
rect 302236 408858 302266 408872
rect 302266 408858 302278 408872
rect 302278 408858 302292 408872
rect 302316 408858 302330 408872
rect 302330 408858 302342 408872
rect 302342 408858 302372 408872
rect 302396 408858 302406 408872
rect 302406 408858 302452 408872
rect 302156 408820 302202 408834
rect 302202 408820 302212 408834
rect 302236 408820 302266 408834
rect 302266 408820 302278 408834
rect 302278 408820 302292 408834
rect 302316 408820 302330 408834
rect 302330 408820 302342 408834
rect 302342 408820 302372 408834
rect 302396 408820 302406 408834
rect 302406 408820 302452 408834
rect 302156 408808 302212 408820
rect 302236 408808 302292 408820
rect 302316 408808 302372 408820
rect 302396 408808 302452 408820
rect 302156 408778 302202 408808
rect 302202 408778 302212 408808
rect 302236 408778 302266 408808
rect 302266 408778 302278 408808
rect 302278 408778 302292 408808
rect 302316 408778 302330 408808
rect 302330 408778 302342 408808
rect 302342 408778 302372 408808
rect 302396 408778 302406 408808
rect 302406 408778 302452 408808
rect 302156 408744 302212 408754
rect 302236 408744 302292 408754
rect 302316 408744 302372 408754
rect 302396 408744 302452 408754
rect 302156 408698 302202 408744
rect 302202 408698 302212 408744
rect 302236 408698 302266 408744
rect 302266 408698 302278 408744
rect 302278 408698 302292 408744
rect 302316 408698 302330 408744
rect 302330 408698 302342 408744
rect 302342 408698 302372 408744
rect 302396 408698 302406 408744
rect 302406 408698 302452 408744
rect 298834 406952 298890 407008
rect 294970 390632 295026 390688
rect 301594 390632 301650 390688
rect 296888 389035 296934 389081
rect 296934 389035 296944 389081
rect 296968 389035 296998 389081
rect 296998 389035 297010 389081
rect 297010 389035 297024 389081
rect 297048 389035 297062 389081
rect 297062 389035 297074 389081
rect 297074 389035 297104 389081
rect 297128 389035 297138 389081
rect 297138 389035 297184 389081
rect 296888 389025 296944 389035
rect 296968 389025 297024 389035
rect 297048 389025 297104 389035
rect 297128 389025 297184 389035
rect 296888 388971 296934 389001
rect 296934 388971 296944 389001
rect 296968 388971 296998 389001
rect 296998 388971 297010 389001
rect 297010 388971 297024 389001
rect 297048 388971 297062 389001
rect 297062 388971 297074 389001
rect 297074 388971 297104 389001
rect 297128 388971 297138 389001
rect 297138 388971 297184 389001
rect 296888 388959 296944 388971
rect 296968 388959 297024 388971
rect 297048 388959 297104 388971
rect 297128 388959 297184 388971
rect 296888 388945 296934 388959
rect 296934 388945 296944 388959
rect 296968 388945 296998 388959
rect 296998 388945 297010 388959
rect 297010 388945 297024 388959
rect 297048 388945 297062 388959
rect 297062 388945 297074 388959
rect 297074 388945 297104 388959
rect 297128 388945 297138 388959
rect 297138 388945 297184 388959
rect 310888 407862 310934 407908
rect 310934 407862 310944 407908
rect 310968 407862 310998 407908
rect 310998 407862 311010 407908
rect 311010 407862 311024 407908
rect 311048 407862 311062 407908
rect 311062 407862 311074 407908
rect 311074 407862 311104 407908
rect 311128 407862 311138 407908
rect 311138 407862 311184 407908
rect 310888 407852 310944 407862
rect 310968 407852 311024 407862
rect 311048 407852 311104 407862
rect 311128 407852 311184 407862
rect 310888 407798 310934 407828
rect 310934 407798 310944 407828
rect 310968 407798 310998 407828
rect 310998 407798 311010 407828
rect 311010 407798 311024 407828
rect 311048 407798 311062 407828
rect 311062 407798 311074 407828
rect 311074 407798 311104 407828
rect 311128 407798 311138 407828
rect 311138 407798 311184 407828
rect 310888 407786 310944 407798
rect 310968 407786 311024 407798
rect 311048 407786 311104 407798
rect 311128 407786 311184 407798
rect 310888 407772 310934 407786
rect 310934 407772 310944 407786
rect 310968 407772 310998 407786
rect 310998 407772 311010 407786
rect 311010 407772 311024 407786
rect 311048 407772 311062 407786
rect 311062 407772 311074 407786
rect 311074 407772 311104 407786
rect 311128 407772 311138 407786
rect 311138 407772 311184 407786
rect 310888 407734 310934 407748
rect 310934 407734 310944 407748
rect 310968 407734 310998 407748
rect 310998 407734 311010 407748
rect 311010 407734 311024 407748
rect 311048 407734 311062 407748
rect 311062 407734 311074 407748
rect 311074 407734 311104 407748
rect 311128 407734 311138 407748
rect 311138 407734 311184 407748
rect 310888 407722 310944 407734
rect 310968 407722 311024 407734
rect 311048 407722 311104 407734
rect 311128 407722 311184 407734
rect 310888 407692 310934 407722
rect 310934 407692 310944 407722
rect 310968 407692 310998 407722
rect 310998 407692 311010 407722
rect 311010 407692 311024 407722
rect 311048 407692 311062 407722
rect 311062 407692 311074 407722
rect 311074 407692 311104 407722
rect 311128 407692 311138 407722
rect 311138 407692 311184 407722
rect 310888 407658 310944 407668
rect 310968 407658 311024 407668
rect 311048 407658 311104 407668
rect 311128 407658 311184 407668
rect 310888 407612 310934 407658
rect 310934 407612 310944 407658
rect 310968 407612 310998 407658
rect 310998 407612 311010 407658
rect 311010 407612 311024 407658
rect 311048 407612 311062 407658
rect 311062 407612 311074 407658
rect 311074 407612 311104 407658
rect 311128 407612 311138 407658
rect 311138 407612 311184 407658
rect 308678 406272 308734 406328
rect 305918 391448 305974 391504
rect 305550 391176 305606 391232
rect 301962 389816 302018 389872
rect 303888 389035 303934 389081
rect 303934 389035 303944 389081
rect 303968 389035 303998 389081
rect 303998 389035 304010 389081
rect 304010 389035 304024 389081
rect 304048 389035 304062 389081
rect 304062 389035 304074 389081
rect 304074 389035 304104 389081
rect 304128 389035 304138 389081
rect 304138 389035 304184 389081
rect 303888 389025 303944 389035
rect 303968 389025 304024 389035
rect 304048 389025 304104 389035
rect 304128 389025 304184 389035
rect 303888 388971 303934 389001
rect 303934 388971 303944 389001
rect 303968 388971 303998 389001
rect 303998 388971 304010 389001
rect 304010 388971 304024 389001
rect 304048 388971 304062 389001
rect 304062 388971 304074 389001
rect 304074 388971 304104 389001
rect 304128 388971 304138 389001
rect 304138 388971 304184 389001
rect 303888 388959 303944 388971
rect 303968 388959 304024 388971
rect 304048 388959 304104 388971
rect 304128 388959 304184 388971
rect 303888 388945 303934 388959
rect 303934 388945 303944 388959
rect 303968 388945 303998 388959
rect 303998 388945 304010 388959
rect 304010 388945 304024 388959
rect 304048 388945 304062 388959
rect 304062 388945 304074 388959
rect 304074 388945 304104 388959
rect 304128 388945 304138 388959
rect 304138 388945 304184 388959
rect 296888 388907 296934 388921
rect 296934 388907 296944 388921
rect 296968 388907 296998 388921
rect 296998 388907 297010 388921
rect 297010 388907 297024 388921
rect 297048 388907 297062 388921
rect 297062 388907 297074 388921
rect 297074 388907 297104 388921
rect 297128 388907 297138 388921
rect 297138 388907 297184 388921
rect 296888 388895 296944 388907
rect 296968 388895 297024 388907
rect 297048 388895 297104 388907
rect 297128 388895 297184 388907
rect 296888 388865 296934 388895
rect 296934 388865 296944 388895
rect 296968 388865 296998 388895
rect 296998 388865 297010 388895
rect 297010 388865 297024 388895
rect 297048 388865 297062 388895
rect 297062 388865 297074 388895
rect 297074 388865 297104 388895
rect 297128 388865 297138 388895
rect 297138 388865 297184 388895
rect 301594 388864 301650 388920
rect 312174 407904 312230 407960
rect 312266 391448 312322 391504
rect 309506 390632 309562 390688
rect 312082 390632 312138 390688
rect 312266 390632 312322 390688
rect 315302 450608 315358 450664
rect 314290 448160 314346 448216
rect 313922 389952 313978 390008
rect 310888 389035 310934 389081
rect 310934 389035 310944 389081
rect 310968 389035 310998 389081
rect 310998 389035 311010 389081
rect 311010 389035 311024 389081
rect 311048 389035 311062 389081
rect 311062 389035 311074 389081
rect 311074 389035 311104 389081
rect 311128 389035 311138 389081
rect 311138 389035 311184 389081
rect 310888 389025 310944 389035
rect 310968 389025 311024 389035
rect 311048 389025 311104 389035
rect 311128 389025 311184 389035
rect 310888 388971 310934 389001
rect 310934 388971 310944 389001
rect 310968 388971 310998 389001
rect 310998 388971 311010 389001
rect 311010 388971 311024 389001
rect 311048 388971 311062 389001
rect 311062 388971 311074 389001
rect 311074 388971 311104 389001
rect 311128 388971 311138 389001
rect 311138 388971 311184 389001
rect 310888 388959 310944 388971
rect 310968 388959 311024 388971
rect 311048 388959 311104 388971
rect 311128 388959 311184 388971
rect 310888 388945 310934 388959
rect 310934 388945 310944 388959
rect 310968 388945 310998 388959
rect 310998 388945 311010 388959
rect 311010 388945 311024 388959
rect 311048 388945 311062 388959
rect 311062 388945 311074 388959
rect 311074 388945 311104 388959
rect 311128 388945 311138 388959
rect 311138 388945 311184 388959
rect 303888 388907 303934 388921
rect 303934 388907 303944 388921
rect 303968 388907 303998 388921
rect 303998 388907 304010 388921
rect 304010 388907 304024 388921
rect 304048 388907 304062 388921
rect 304062 388907 304074 388921
rect 304074 388907 304104 388921
rect 304128 388907 304138 388921
rect 304138 388907 304184 388921
rect 303888 388895 303944 388907
rect 303968 388895 304024 388907
rect 304048 388895 304104 388907
rect 304128 388895 304184 388907
rect 303888 388865 303934 388895
rect 303934 388865 303944 388895
rect 303968 388865 303998 388895
rect 303998 388865 304010 388895
rect 304010 388865 304024 388895
rect 304048 388865 304062 388895
rect 304062 388865 304074 388895
rect 304074 388865 304104 388895
rect 304128 388865 304138 388895
rect 304138 388865 304184 388895
rect 296888 388831 296944 388841
rect 296968 388831 297024 388841
rect 297048 388831 297104 388841
rect 297128 388831 297184 388841
rect 296888 388785 296934 388831
rect 296934 388785 296944 388831
rect 296968 388785 296998 388831
rect 296998 388785 297010 388831
rect 297010 388785 297024 388831
rect 297048 388785 297062 388831
rect 297062 388785 297074 388831
rect 297074 388785 297104 388831
rect 297128 388785 297138 388831
rect 297138 388785 297184 388831
rect 305918 388864 305974 388920
rect 309506 388864 309562 388920
rect 310888 388907 310934 388921
rect 310934 388907 310944 388921
rect 310968 388907 310998 388921
rect 310998 388907 311010 388921
rect 311010 388907 311024 388921
rect 311048 388907 311062 388921
rect 311062 388907 311074 388921
rect 311074 388907 311104 388921
rect 311128 388907 311138 388921
rect 311138 388907 311184 388921
rect 310888 388895 310944 388907
rect 310968 388895 311024 388907
rect 311048 388895 311104 388907
rect 311128 388895 311184 388907
rect 310888 388865 310934 388895
rect 310934 388865 310944 388895
rect 310968 388865 310998 388895
rect 310998 388865 311010 388895
rect 311010 388865 311024 388895
rect 311048 388865 311062 388895
rect 311062 388865 311074 388895
rect 311074 388865 311104 388895
rect 311128 388865 311138 388895
rect 311138 388865 311184 388895
rect 303888 388831 303944 388841
rect 303968 388831 304024 388841
rect 304048 388831 304104 388841
rect 304128 388831 304184 388841
rect 303888 388785 303934 388831
rect 303934 388785 303944 388831
rect 303968 388785 303998 388831
rect 303998 388785 304010 388831
rect 304010 388785 304024 388831
rect 304048 388785 304062 388831
rect 304062 388785 304074 388831
rect 304074 388785 304104 388831
rect 304128 388785 304138 388831
rect 304138 388785 304184 388831
rect 310888 388831 310944 388841
rect 310968 388831 311024 388841
rect 311048 388831 311104 388841
rect 311128 388831 311184 388841
rect 310888 388785 310934 388831
rect 310934 388785 310944 388831
rect 310968 388785 310998 388831
rect 310998 388785 311010 388831
rect 311010 388785 311024 388831
rect 311048 388785 311062 388831
rect 311062 388785 311074 388831
rect 311074 388785 311104 388831
rect 311128 388785 311138 388831
rect 311138 388785 311184 388831
rect 301594 388592 301650 388648
rect 309506 388592 309562 388648
rect 305890 388456 305946 388512
rect 314474 427352 314530 427408
rect 314382 390632 314438 390688
rect 314290 388320 314346 388376
rect 295156 387952 295202 387998
rect 295202 387952 295212 387998
rect 295236 387952 295266 387998
rect 295266 387952 295278 387998
rect 295278 387952 295292 387998
rect 295316 387952 295330 387998
rect 295330 387952 295342 387998
rect 295342 387952 295372 387998
rect 295396 387952 295406 387998
rect 295406 387952 295452 387998
rect 295156 387942 295212 387952
rect 295236 387942 295292 387952
rect 295316 387942 295372 387952
rect 295396 387942 295452 387952
rect 295156 387888 295202 387918
rect 295202 387888 295212 387918
rect 295236 387888 295266 387918
rect 295266 387888 295278 387918
rect 295278 387888 295292 387918
rect 295316 387888 295330 387918
rect 295330 387888 295342 387918
rect 295342 387888 295372 387918
rect 295396 387888 295406 387918
rect 295406 387888 295452 387918
rect 295156 387876 295212 387888
rect 295236 387876 295292 387888
rect 295316 387876 295372 387888
rect 295396 387876 295452 387888
rect 295156 387862 295202 387876
rect 295202 387862 295212 387876
rect 295236 387862 295266 387876
rect 295266 387862 295278 387876
rect 295278 387862 295292 387876
rect 295316 387862 295330 387876
rect 295330 387862 295342 387876
rect 295342 387862 295372 387876
rect 295396 387862 295406 387876
rect 295406 387862 295452 387876
rect 295156 387824 295202 387838
rect 295202 387824 295212 387838
rect 295236 387824 295266 387838
rect 295266 387824 295278 387838
rect 295278 387824 295292 387838
rect 295316 387824 295330 387838
rect 295330 387824 295342 387838
rect 295342 387824 295372 387838
rect 295396 387824 295406 387838
rect 295406 387824 295452 387838
rect 295156 387812 295212 387824
rect 295236 387812 295292 387824
rect 295316 387812 295372 387824
rect 295396 387812 295452 387824
rect 295156 387782 295202 387812
rect 295202 387782 295212 387812
rect 295236 387782 295266 387812
rect 295266 387782 295278 387812
rect 295278 387782 295292 387812
rect 295316 387782 295330 387812
rect 295330 387782 295342 387812
rect 295342 387782 295372 387812
rect 295396 387782 295406 387812
rect 295406 387782 295452 387812
rect 295156 387748 295212 387758
rect 295236 387748 295292 387758
rect 295316 387748 295372 387758
rect 295396 387748 295452 387758
rect 295156 387702 295202 387748
rect 295202 387702 295212 387748
rect 295236 387702 295266 387748
rect 295266 387702 295278 387748
rect 295278 387702 295292 387748
rect 295316 387702 295330 387748
rect 295330 387702 295342 387748
rect 295342 387702 295372 387748
rect 295396 387702 295406 387748
rect 295406 387702 295452 387748
rect 302156 387947 302202 387993
rect 302202 387947 302212 387993
rect 302236 387947 302266 387993
rect 302266 387947 302278 387993
rect 302278 387947 302292 387993
rect 302316 387947 302330 387993
rect 302330 387947 302342 387993
rect 302342 387947 302372 387993
rect 302396 387947 302406 387993
rect 302406 387947 302452 387993
rect 302156 387937 302212 387947
rect 302236 387937 302292 387947
rect 302316 387937 302372 387947
rect 302396 387937 302452 387947
rect 302156 387883 302202 387913
rect 302202 387883 302212 387913
rect 302236 387883 302266 387913
rect 302266 387883 302278 387913
rect 302278 387883 302292 387913
rect 302316 387883 302330 387913
rect 302330 387883 302342 387913
rect 302342 387883 302372 387913
rect 302396 387883 302406 387913
rect 302406 387883 302452 387913
rect 302156 387871 302212 387883
rect 302236 387871 302292 387883
rect 302316 387871 302372 387883
rect 302396 387871 302452 387883
rect 302156 387857 302202 387871
rect 302202 387857 302212 387871
rect 302236 387857 302266 387871
rect 302266 387857 302278 387871
rect 302278 387857 302292 387871
rect 302316 387857 302330 387871
rect 302330 387857 302342 387871
rect 302342 387857 302372 387871
rect 302396 387857 302406 387871
rect 302406 387857 302452 387871
rect 302156 387819 302202 387833
rect 302202 387819 302212 387833
rect 302236 387819 302266 387833
rect 302266 387819 302278 387833
rect 302278 387819 302292 387833
rect 302316 387819 302330 387833
rect 302330 387819 302342 387833
rect 302342 387819 302372 387833
rect 302396 387819 302406 387833
rect 302406 387819 302452 387833
rect 302156 387807 302212 387819
rect 302236 387807 302292 387819
rect 302316 387807 302372 387819
rect 302396 387807 302452 387819
rect 302156 387777 302202 387807
rect 302202 387777 302212 387807
rect 302236 387777 302266 387807
rect 302266 387777 302278 387807
rect 302278 387777 302292 387807
rect 302316 387777 302330 387807
rect 302330 387777 302342 387807
rect 302342 387777 302372 387807
rect 302396 387777 302406 387807
rect 302406 387777 302452 387807
rect 302156 387743 302212 387753
rect 302236 387743 302292 387753
rect 302316 387743 302372 387753
rect 302396 387743 302452 387753
rect 302156 387697 302202 387743
rect 302202 387697 302212 387743
rect 302236 387697 302266 387743
rect 302266 387697 302278 387743
rect 302278 387697 302292 387743
rect 302316 387697 302330 387743
rect 302330 387697 302342 387743
rect 302342 387697 302372 387743
rect 302396 387697 302406 387743
rect 302406 387697 302452 387743
rect 309156 387947 309202 387993
rect 309202 387947 309212 387993
rect 309236 387947 309266 387993
rect 309266 387947 309278 387993
rect 309278 387947 309292 387993
rect 309316 387947 309330 387993
rect 309330 387947 309342 387993
rect 309342 387947 309372 387993
rect 309396 387947 309406 387993
rect 309406 387947 309452 387993
rect 309156 387937 309212 387947
rect 309236 387937 309292 387947
rect 309316 387937 309372 387947
rect 309396 387937 309452 387947
rect 309156 387883 309202 387913
rect 309202 387883 309212 387913
rect 309236 387883 309266 387913
rect 309266 387883 309278 387913
rect 309278 387883 309292 387913
rect 309316 387883 309330 387913
rect 309330 387883 309342 387913
rect 309342 387883 309372 387913
rect 309396 387883 309406 387913
rect 309406 387883 309452 387913
rect 309156 387871 309212 387883
rect 309236 387871 309292 387883
rect 309316 387871 309372 387883
rect 309396 387871 309452 387883
rect 309156 387857 309202 387871
rect 309202 387857 309212 387871
rect 309236 387857 309266 387871
rect 309266 387857 309278 387871
rect 309278 387857 309292 387871
rect 309316 387857 309330 387871
rect 309330 387857 309342 387871
rect 309342 387857 309372 387871
rect 309396 387857 309406 387871
rect 309406 387857 309452 387871
rect 309156 387819 309202 387833
rect 309202 387819 309212 387833
rect 309236 387819 309266 387833
rect 309266 387819 309278 387833
rect 309278 387819 309292 387833
rect 309316 387819 309330 387833
rect 309330 387819 309342 387833
rect 309342 387819 309372 387833
rect 309396 387819 309406 387833
rect 309406 387819 309452 387833
rect 309156 387807 309212 387819
rect 309236 387807 309292 387819
rect 309316 387807 309372 387819
rect 309396 387807 309452 387819
rect 309156 387777 309202 387807
rect 309202 387777 309212 387807
rect 309236 387777 309266 387807
rect 309266 387777 309278 387807
rect 309278 387777 309292 387807
rect 309316 387777 309330 387807
rect 309330 387777 309342 387807
rect 309342 387777 309372 387807
rect 309396 387777 309406 387807
rect 309406 387777 309452 387807
rect 309156 387743 309212 387753
rect 309236 387743 309292 387753
rect 309316 387743 309372 387753
rect 309396 387743 309452 387753
rect 309156 387697 309202 387743
rect 309202 387697 309212 387743
rect 309236 387697 309266 387743
rect 309266 387697 309278 387743
rect 309278 387697 309292 387743
rect 309316 387697 309330 387743
rect 309330 387697 309342 387743
rect 309342 387697 309372 387743
rect 309396 387697 309406 387743
rect 309406 387697 309452 387743
rect 303964 387396 304020 387398
rect 303964 387344 303966 387396
rect 303966 387344 304018 387396
rect 304018 387344 304020 387396
rect 303964 387342 304020 387344
rect 299294 384920 299350 384976
rect 311044 387513 311100 387515
rect 311044 387461 311046 387513
rect 311046 387461 311098 387513
rect 311098 387461 311100 387513
rect 311044 387459 311100 387461
rect 310058 386416 310114 386472
rect 307666 386280 307722 386336
rect 309598 386280 309654 386336
rect 306746 384240 306802 384296
rect 303158 374176 303214 374232
rect 304538 368872 304594 368928
rect 295246 368464 295302 368520
rect 313278 386416 313334 386472
rect 310426 384784 310482 384840
rect 312542 384784 312598 384840
rect 310978 368872 311034 368928
rect 304538 367920 304594 367976
rect 307574 367920 307630 367976
rect 310058 367920 310114 367976
rect 303909 367512 303965 367568
rect 307574 367512 307630 367568
rect 299754 367290 299810 367296
rect 299754 367240 299756 367290
rect 299756 367240 299808 367290
rect 299808 367240 299810 367290
rect 310058 367512 310114 367568
rect 301686 364248 301742 364304
rect 298650 364112 298706 364168
rect 304722 348336 304778 348392
rect 295246 347792 295302 347848
rect 300858 347792 300914 347848
rect 304446 347792 304502 347848
rect 296888 347035 296934 347081
rect 296934 347035 296944 347081
rect 296968 347035 296998 347081
rect 296998 347035 297010 347081
rect 297010 347035 297024 347081
rect 297048 347035 297062 347081
rect 297062 347035 297074 347081
rect 297074 347035 297104 347081
rect 297128 347035 297138 347081
rect 297138 347035 297184 347081
rect 296888 347025 296944 347035
rect 296968 347025 297024 347035
rect 297048 347025 297104 347035
rect 297128 347025 297184 347035
rect 296888 346971 296934 347001
rect 296934 346971 296944 347001
rect 296968 346971 296998 347001
rect 296998 346971 297010 347001
rect 297010 346971 297024 347001
rect 297048 346971 297062 347001
rect 297062 346971 297074 347001
rect 297074 346971 297104 347001
rect 297128 346971 297138 347001
rect 297138 346971 297184 347001
rect 296888 346959 296944 346971
rect 296968 346959 297024 346971
rect 297048 346959 297104 346971
rect 297128 346959 297184 346971
rect 296888 346945 296934 346959
rect 296934 346945 296944 346959
rect 296968 346945 296998 346959
rect 296998 346945 297010 346959
rect 297010 346945 297024 346959
rect 297048 346945 297062 346959
rect 297062 346945 297074 346959
rect 297074 346945 297104 346959
rect 297128 346945 297138 346959
rect 297138 346945 297184 346959
rect 296888 346907 296934 346921
rect 296934 346907 296944 346921
rect 296968 346907 296998 346921
rect 296998 346907 297010 346921
rect 297010 346907 297024 346921
rect 297048 346907 297062 346921
rect 297062 346907 297074 346921
rect 297074 346907 297104 346921
rect 297128 346907 297138 346921
rect 297138 346907 297184 346921
rect 296888 346895 296944 346907
rect 296968 346895 297024 346907
rect 297048 346895 297104 346907
rect 297128 346895 297184 346907
rect 303888 347035 303934 347081
rect 303934 347035 303944 347081
rect 303968 347035 303998 347081
rect 303998 347035 304010 347081
rect 304010 347035 304024 347081
rect 304048 347035 304062 347081
rect 304062 347035 304074 347081
rect 304074 347035 304104 347081
rect 304128 347035 304138 347081
rect 304138 347035 304184 347081
rect 303888 347025 303944 347035
rect 303968 347025 304024 347035
rect 304048 347025 304104 347035
rect 304128 347025 304184 347035
rect 303888 346971 303934 347001
rect 303934 346971 303944 347001
rect 303968 346971 303998 347001
rect 303998 346971 304010 347001
rect 304010 346971 304024 347001
rect 304048 346971 304062 347001
rect 304062 346971 304074 347001
rect 304074 346971 304104 347001
rect 304128 346971 304138 347001
rect 304138 346971 304184 347001
rect 303888 346959 303944 346971
rect 303968 346959 304024 346971
rect 304048 346959 304104 346971
rect 304128 346959 304184 346971
rect 303888 346945 303934 346959
rect 303934 346945 303944 346959
rect 303968 346945 303998 346959
rect 303998 346945 304010 346959
rect 304010 346945 304024 346959
rect 304048 346945 304062 346959
rect 304062 346945 304074 346959
rect 304074 346945 304104 346959
rect 304128 346945 304138 346959
rect 304138 346945 304184 346959
rect 303888 346907 303934 346921
rect 303934 346907 303944 346921
rect 303968 346907 303998 346921
rect 303998 346907 304010 346921
rect 304010 346907 304024 346921
rect 304048 346907 304062 346921
rect 304062 346907 304074 346921
rect 304074 346907 304104 346921
rect 304128 346907 304138 346921
rect 304138 346907 304184 346921
rect 296888 346865 296934 346895
rect 296934 346865 296944 346895
rect 296968 346865 296998 346895
rect 296998 346865 297010 346895
rect 297010 346865 297024 346895
rect 297048 346865 297062 346895
rect 297062 346865 297074 346895
rect 297074 346865 297104 346895
rect 297128 346865 297138 346895
rect 297138 346865 297184 346895
rect 296888 346831 296944 346841
rect 296968 346831 297024 346841
rect 297048 346831 297104 346841
rect 297128 346831 297184 346841
rect 300858 346840 300914 346896
rect 303888 346895 303944 346907
rect 303968 346895 304024 346907
rect 304048 346895 304104 346907
rect 304128 346895 304184 346907
rect 307942 363024 307998 363080
rect 307666 347248 307722 347304
rect 310978 347792 311034 347848
rect 303888 346865 303934 346895
rect 303934 346865 303944 346895
rect 303968 346865 303998 346895
rect 303998 346865 304010 346895
rect 304010 346865 304024 346895
rect 304048 346865 304062 346895
rect 304062 346865 304074 346895
rect 304074 346865 304104 346895
rect 304128 346865 304138 346895
rect 304138 346865 304184 346895
rect 303888 346831 303944 346841
rect 303968 346831 304024 346841
rect 304048 346831 304104 346841
rect 304128 346831 304184 346841
rect 304446 346840 304502 346896
rect 307666 346840 307722 346896
rect 310518 346840 310574 346896
rect 296888 346785 296934 346831
rect 296934 346785 296944 346831
rect 296968 346785 296998 346831
rect 296998 346785 297010 346831
rect 297010 346785 297024 346831
rect 297048 346785 297062 346831
rect 297062 346785 297074 346831
rect 297074 346785 297104 346831
rect 297128 346785 297138 346831
rect 297138 346785 297184 346831
rect 303888 346785 303934 346831
rect 303934 346785 303944 346831
rect 303968 346785 303998 346831
rect 303998 346785 304010 346831
rect 304010 346785 304024 346831
rect 304048 346785 304062 346831
rect 304062 346785 304074 346831
rect 304074 346785 304104 346831
rect 304128 346785 304138 346831
rect 304138 346785 304184 346831
rect 300858 346568 300914 346624
rect 303894 346568 303950 346624
rect 306746 346568 306802 346624
rect 309874 346568 309930 346624
rect 302156 345933 302202 345979
rect 302202 345933 302212 345979
rect 302236 345933 302266 345979
rect 302266 345933 302278 345979
rect 302278 345933 302292 345979
rect 302316 345933 302330 345979
rect 302330 345933 302342 345979
rect 302342 345933 302372 345979
rect 302396 345933 302406 345979
rect 302406 345933 302452 345979
rect 302156 345923 302212 345933
rect 302236 345923 302292 345933
rect 302316 345923 302372 345933
rect 302396 345923 302452 345933
rect 302156 345869 302202 345899
rect 302202 345869 302212 345899
rect 302236 345869 302266 345899
rect 302266 345869 302278 345899
rect 302278 345869 302292 345899
rect 302316 345869 302330 345899
rect 302330 345869 302342 345899
rect 302342 345869 302372 345899
rect 302396 345869 302406 345899
rect 302406 345869 302452 345899
rect 302156 345857 302212 345869
rect 302236 345857 302292 345869
rect 302316 345857 302372 345869
rect 302396 345857 302452 345869
rect 302156 345843 302202 345857
rect 302202 345843 302212 345857
rect 302236 345843 302266 345857
rect 302266 345843 302278 345857
rect 302278 345843 302292 345857
rect 302316 345843 302330 345857
rect 302330 345843 302342 345857
rect 302342 345843 302372 345857
rect 302396 345843 302406 345857
rect 302406 345843 302452 345857
rect 302156 345805 302202 345819
rect 302202 345805 302212 345819
rect 302236 345805 302266 345819
rect 302266 345805 302278 345819
rect 302278 345805 302292 345819
rect 302316 345805 302330 345819
rect 302330 345805 302342 345819
rect 302342 345805 302372 345819
rect 302396 345805 302406 345819
rect 302406 345805 302452 345819
rect 302156 345793 302212 345805
rect 302236 345793 302292 345805
rect 302316 345793 302372 345805
rect 302396 345793 302452 345805
rect 302156 345763 302202 345793
rect 302202 345763 302212 345793
rect 302236 345763 302266 345793
rect 302266 345763 302278 345793
rect 302278 345763 302292 345793
rect 302316 345763 302330 345793
rect 302330 345763 302342 345793
rect 302342 345763 302372 345793
rect 302396 345763 302406 345793
rect 302406 345763 302452 345793
rect 302156 345729 302212 345739
rect 302236 345729 302292 345739
rect 302316 345729 302372 345739
rect 302396 345729 302452 345739
rect 302156 345683 302202 345729
rect 302202 345683 302212 345729
rect 302236 345683 302266 345729
rect 302266 345683 302278 345729
rect 302278 345683 302292 345729
rect 302316 345683 302330 345729
rect 302330 345683 302342 345729
rect 302342 345683 302372 345729
rect 302396 345683 302406 345729
rect 302406 345683 302452 345729
rect 309156 345933 309202 345979
rect 309202 345933 309212 345979
rect 309236 345933 309266 345979
rect 309266 345933 309278 345979
rect 309278 345933 309292 345979
rect 309316 345933 309330 345979
rect 309330 345933 309342 345979
rect 309342 345933 309372 345979
rect 309396 345933 309406 345979
rect 309406 345933 309452 345979
rect 309156 345923 309212 345933
rect 309236 345923 309292 345933
rect 309316 345923 309372 345933
rect 309396 345923 309452 345933
rect 309156 345869 309202 345899
rect 309202 345869 309212 345899
rect 309236 345869 309266 345899
rect 309266 345869 309278 345899
rect 309278 345869 309292 345899
rect 309316 345869 309330 345899
rect 309330 345869 309342 345899
rect 309342 345869 309372 345899
rect 309396 345869 309406 345899
rect 309406 345869 309452 345899
rect 309156 345857 309212 345869
rect 309236 345857 309292 345869
rect 309316 345857 309372 345869
rect 309396 345857 309452 345869
rect 309156 345843 309202 345857
rect 309202 345843 309212 345857
rect 309236 345843 309266 345857
rect 309266 345843 309278 345857
rect 309278 345843 309292 345857
rect 309316 345843 309330 345857
rect 309330 345843 309342 345857
rect 309342 345843 309372 345857
rect 309396 345843 309406 345857
rect 309406 345843 309452 345857
rect 309156 345805 309202 345819
rect 309202 345805 309212 345819
rect 309236 345805 309266 345819
rect 309266 345805 309278 345819
rect 309278 345805 309292 345819
rect 309316 345805 309330 345819
rect 309330 345805 309342 345819
rect 309342 345805 309372 345819
rect 309396 345805 309406 345819
rect 309406 345805 309452 345819
rect 309156 345793 309212 345805
rect 309236 345793 309292 345805
rect 309316 345793 309372 345805
rect 309396 345793 309452 345805
rect 309156 345763 309202 345793
rect 309202 345763 309212 345793
rect 309236 345763 309266 345793
rect 309266 345763 309278 345793
rect 309278 345763 309292 345793
rect 309316 345763 309330 345793
rect 309330 345763 309342 345793
rect 309342 345763 309372 345793
rect 309396 345763 309406 345793
rect 309406 345763 309452 345793
rect 309156 345729 309212 345739
rect 309236 345729 309292 345739
rect 309316 345729 309372 345739
rect 309396 345729 309452 345739
rect 309156 345683 309202 345729
rect 309202 345683 309212 345729
rect 309236 345683 309266 345729
rect 309266 345683 309278 345729
rect 309278 345683 309292 345729
rect 309316 345683 309330 345729
rect 309330 345683 309342 345729
rect 309342 345683 309372 345729
rect 309396 345683 309406 345729
rect 309406 345683 309452 345729
rect 301686 343576 301742 343632
rect 298650 343440 298706 343496
rect 307942 342216 307998 342272
rect 307666 340176 307722 340232
rect 304722 331472 304778 331528
rect 304906 327664 304962 327720
rect 295246 327120 295302 327176
rect 300858 327120 300914 327176
rect 296888 326034 296934 326080
rect 296934 326034 296944 326080
rect 296968 326034 296998 326080
rect 296998 326034 297010 326080
rect 297010 326034 297024 326080
rect 297048 326034 297062 326080
rect 297062 326034 297074 326080
rect 297074 326034 297104 326080
rect 297128 326034 297138 326080
rect 297138 326034 297184 326080
rect 296888 326024 296944 326034
rect 296968 326024 297024 326034
rect 297048 326024 297104 326034
rect 297128 326024 297184 326034
rect 296888 325970 296934 326000
rect 296934 325970 296944 326000
rect 296968 325970 296998 326000
rect 296998 325970 297010 326000
rect 297010 325970 297024 326000
rect 297048 325970 297062 326000
rect 297062 325970 297074 326000
rect 297074 325970 297104 326000
rect 297128 325970 297138 326000
rect 297138 325970 297184 326000
rect 296888 325958 296944 325970
rect 296968 325958 297024 325970
rect 297048 325958 297104 325970
rect 297128 325958 297184 325970
rect 303888 326034 303934 326080
rect 303934 326034 303944 326080
rect 303968 326034 303998 326080
rect 303998 326034 304010 326080
rect 304010 326034 304024 326080
rect 304048 326034 304062 326080
rect 304062 326034 304074 326080
rect 304074 326034 304104 326080
rect 304128 326034 304138 326080
rect 304138 326034 304184 326080
rect 303888 326024 303944 326034
rect 303968 326024 304024 326034
rect 304048 326024 304104 326034
rect 304128 326024 304184 326034
rect 303888 325970 303934 326000
rect 303934 325970 303944 326000
rect 303968 325970 303998 326000
rect 303998 325970 304010 326000
rect 304010 325970 304024 326000
rect 304048 325970 304062 326000
rect 304062 325970 304074 326000
rect 304074 325970 304104 326000
rect 304128 325970 304138 326000
rect 304138 325970 304184 326000
rect 296888 325944 296934 325958
rect 296934 325944 296944 325958
rect 296968 325944 296998 325958
rect 296998 325944 297010 325958
rect 297010 325944 297024 325958
rect 297048 325944 297062 325958
rect 297062 325944 297074 325958
rect 297074 325944 297104 325958
rect 297128 325944 297138 325958
rect 297138 325944 297184 325958
rect 296888 325906 296934 325920
rect 296934 325906 296944 325920
rect 296968 325906 296998 325920
rect 296998 325906 297010 325920
rect 297010 325906 297024 325920
rect 297048 325906 297062 325920
rect 297062 325906 297074 325920
rect 297074 325906 297104 325920
rect 297128 325906 297138 325920
rect 297138 325906 297184 325920
rect 296888 325894 296944 325906
rect 296968 325894 297024 325906
rect 297048 325894 297104 325906
rect 297128 325894 297184 325906
rect 296888 325864 296934 325894
rect 296934 325864 296944 325894
rect 296968 325864 296998 325894
rect 296998 325864 297010 325894
rect 297010 325864 297024 325894
rect 297048 325864 297062 325894
rect 297062 325864 297074 325894
rect 297074 325864 297104 325894
rect 297128 325864 297138 325894
rect 297138 325864 297184 325894
rect 300858 325896 300914 325952
rect 303888 325958 303944 325970
rect 303968 325958 304024 325970
rect 304048 325958 304104 325970
rect 304128 325958 304184 325970
rect 311070 346704 311126 346760
rect 311070 340176 311126 340232
rect 310978 328344 311034 328400
rect 310978 327664 311034 327720
rect 307666 326168 307722 326224
rect 310888 326034 310934 326080
rect 310934 326034 310944 326080
rect 310968 326034 310998 326080
rect 310998 326034 311010 326080
rect 311010 326034 311024 326080
rect 311048 326034 311062 326080
rect 311062 326034 311074 326080
rect 311074 326034 311104 326080
rect 311128 326034 311138 326080
rect 311138 326034 311184 326080
rect 310888 326024 310944 326034
rect 310968 326024 311024 326034
rect 311048 326024 311104 326034
rect 311128 326024 311184 326034
rect 310888 325970 310934 326000
rect 310934 325970 310944 326000
rect 310968 325970 310998 326000
rect 310998 325970 311010 326000
rect 311010 325970 311024 326000
rect 311048 325970 311062 326000
rect 311062 325970 311074 326000
rect 311074 325970 311104 326000
rect 311128 325970 311138 326000
rect 311138 325970 311184 326000
rect 303888 325944 303934 325958
rect 303934 325944 303944 325958
rect 303968 325944 303998 325958
rect 303998 325944 304010 325958
rect 304010 325944 304024 325958
rect 304048 325944 304062 325958
rect 304062 325944 304074 325958
rect 304074 325944 304104 325958
rect 304128 325944 304138 325958
rect 304138 325944 304184 325958
rect 303888 325906 303934 325920
rect 303934 325906 303944 325920
rect 303968 325906 303998 325920
rect 303998 325906 304010 325920
rect 304010 325906 304024 325920
rect 304048 325906 304062 325920
rect 304062 325906 304074 325920
rect 304074 325906 304104 325920
rect 304128 325906 304138 325920
rect 304138 325906 304184 325920
rect 303888 325894 303944 325906
rect 303968 325894 304024 325906
rect 304048 325894 304104 325906
rect 304128 325894 304184 325906
rect 296888 325830 296944 325840
rect 296968 325830 297024 325840
rect 297048 325830 297104 325840
rect 297128 325830 297184 325840
rect 296888 325784 296934 325830
rect 296934 325784 296944 325830
rect 296968 325784 296998 325830
rect 296998 325784 297010 325830
rect 297010 325784 297024 325830
rect 297048 325784 297062 325830
rect 297062 325784 297074 325830
rect 297074 325784 297104 325830
rect 297128 325784 297138 325830
rect 297138 325784 297184 325830
rect 303888 325864 303934 325894
rect 303934 325864 303944 325894
rect 303968 325864 303998 325894
rect 303998 325864 304010 325894
rect 304010 325864 304024 325894
rect 304048 325864 304062 325894
rect 304062 325864 304074 325894
rect 304074 325864 304104 325894
rect 304128 325864 304138 325894
rect 304138 325864 304184 325894
rect 304906 325896 304962 325952
rect 307666 325896 307722 325952
rect 310888 325958 310944 325970
rect 310968 325958 311024 325970
rect 311048 325958 311104 325970
rect 311128 325958 311184 325970
rect 310888 325944 310934 325958
rect 310934 325944 310944 325958
rect 310968 325944 310998 325958
rect 310998 325944 311010 325958
rect 311010 325944 311024 325958
rect 311048 325944 311062 325958
rect 311062 325944 311074 325958
rect 311074 325944 311104 325958
rect 311128 325944 311138 325958
rect 311138 325944 311184 325958
rect 310888 325906 310934 325920
rect 310934 325906 310944 325920
rect 310968 325906 310998 325920
rect 310998 325906 311010 325920
rect 311010 325906 311024 325920
rect 311048 325906 311062 325920
rect 311062 325906 311074 325920
rect 311074 325906 311104 325920
rect 311128 325906 311138 325920
rect 311138 325906 311184 325920
rect 310888 325894 310944 325906
rect 310968 325894 311024 325906
rect 311048 325894 311104 325906
rect 311128 325894 311184 325906
rect 303888 325830 303944 325840
rect 303968 325830 304024 325840
rect 304048 325830 304104 325840
rect 304128 325830 304184 325840
rect 303888 325784 303934 325830
rect 303934 325784 303944 325830
rect 303968 325784 303998 325830
rect 303998 325784 304010 325830
rect 304010 325784 304024 325830
rect 304048 325784 304062 325830
rect 304062 325784 304074 325830
rect 304074 325784 304104 325830
rect 304128 325784 304138 325830
rect 304138 325784 304184 325830
rect 310888 325864 310934 325894
rect 310934 325864 310944 325894
rect 310968 325864 310998 325894
rect 310998 325864 311010 325894
rect 311010 325864 311024 325894
rect 311048 325864 311062 325894
rect 311062 325864 311074 325894
rect 311074 325864 311104 325894
rect 311128 325864 311138 325894
rect 311138 325864 311184 325894
rect 310888 325830 310944 325840
rect 310968 325830 311024 325840
rect 311048 325830 311104 325840
rect 311128 325830 311184 325840
rect 310888 325784 310934 325830
rect 310934 325784 310944 325830
rect 310968 325784 310998 325830
rect 310998 325784 311010 325830
rect 311010 325784 311024 325830
rect 311048 325784 311062 325830
rect 311062 325784 311074 325830
rect 311074 325784 311104 325830
rect 311128 325784 311138 325830
rect 311138 325784 311184 325830
rect 300950 325624 301006 325680
rect 304262 325624 304318 325680
rect 307390 325624 307446 325680
rect 311898 328344 311954 328400
rect 298742 321408 298798 321464
rect 303888 323862 303934 323908
rect 303934 323862 303944 323908
rect 303968 323862 303998 323908
rect 303998 323862 304010 323908
rect 304010 323862 304024 323908
rect 304048 323862 304062 323908
rect 304062 323862 304074 323908
rect 304074 323862 304104 323908
rect 304128 323862 304138 323908
rect 304138 323862 304184 323908
rect 303888 323852 303944 323862
rect 303968 323852 304024 323862
rect 304048 323852 304104 323862
rect 304128 323852 304184 323862
rect 303888 323798 303934 323828
rect 303934 323798 303944 323828
rect 303968 323798 303998 323828
rect 303998 323798 304010 323828
rect 304010 323798 304024 323828
rect 304048 323798 304062 323828
rect 304062 323798 304074 323828
rect 304074 323798 304104 323828
rect 304128 323798 304138 323828
rect 304138 323798 304184 323828
rect 303888 323786 303944 323798
rect 303968 323786 304024 323798
rect 304048 323786 304104 323798
rect 304128 323786 304184 323798
rect 303888 323772 303934 323786
rect 303934 323772 303944 323786
rect 303968 323772 303998 323786
rect 303998 323772 304010 323786
rect 304010 323772 304024 323786
rect 304048 323772 304062 323786
rect 304062 323772 304074 323786
rect 304074 323772 304104 323786
rect 304128 323772 304138 323786
rect 304138 323772 304184 323786
rect 303888 323734 303934 323748
rect 303934 323734 303944 323748
rect 303968 323734 303998 323748
rect 303998 323734 304010 323748
rect 304010 323734 304024 323748
rect 304048 323734 304062 323748
rect 304062 323734 304074 323748
rect 304074 323734 304104 323748
rect 304128 323734 304138 323748
rect 304138 323734 304184 323748
rect 303888 323722 303944 323734
rect 303968 323722 304024 323734
rect 304048 323722 304104 323734
rect 304128 323722 304184 323734
rect 303888 323692 303934 323722
rect 303934 323692 303944 323722
rect 303968 323692 303998 323722
rect 303998 323692 304010 323722
rect 304010 323692 304024 323722
rect 304048 323692 304062 323722
rect 304062 323692 304074 323722
rect 304074 323692 304104 323722
rect 304128 323692 304138 323722
rect 304138 323692 304184 323722
rect 303888 323658 303944 323668
rect 303968 323658 304024 323668
rect 304048 323658 304104 323668
rect 304128 323658 304184 323668
rect 303888 323612 303934 323658
rect 303934 323612 303944 323658
rect 303968 323612 303998 323658
rect 303998 323612 304010 323658
rect 304010 323612 304024 323658
rect 304048 323612 304062 323658
rect 304062 323612 304074 323658
rect 304074 323612 304104 323658
rect 304128 323612 304138 323658
rect 304138 323612 304184 323658
rect 305090 322768 305146 322824
rect 301778 321272 301834 321328
rect 308218 308352 308274 308408
rect 306194 307400 306250 307456
rect 295246 306448 295302 306504
rect 301686 306448 301742 306504
rect 296888 305064 296934 305110
rect 296934 305064 296944 305110
rect 296968 305064 296998 305110
rect 296998 305064 297010 305110
rect 297010 305064 297024 305110
rect 297048 305064 297062 305110
rect 297062 305064 297074 305110
rect 297074 305064 297104 305110
rect 297128 305064 297138 305110
rect 297138 305064 297184 305110
rect 296888 305054 296944 305064
rect 296968 305054 297024 305064
rect 297048 305054 297104 305064
rect 297128 305054 297184 305064
rect 296888 305000 296934 305030
rect 296934 305000 296944 305030
rect 296968 305000 296998 305030
rect 296998 305000 297010 305030
rect 297010 305000 297024 305030
rect 297048 305000 297062 305030
rect 297062 305000 297074 305030
rect 297074 305000 297104 305030
rect 297128 305000 297138 305030
rect 297138 305000 297184 305030
rect 303888 305064 303934 305110
rect 303934 305064 303944 305110
rect 303968 305064 303998 305110
rect 303998 305064 304010 305110
rect 304010 305064 304024 305110
rect 304048 305064 304062 305110
rect 304062 305064 304074 305110
rect 304074 305064 304104 305110
rect 304128 305064 304138 305110
rect 304138 305064 304184 305110
rect 303888 305054 303944 305064
rect 303968 305054 304024 305064
rect 304048 305054 304104 305064
rect 304128 305054 304184 305064
rect 296888 304988 296944 305000
rect 296968 304988 297024 305000
rect 297048 304988 297104 305000
rect 297128 304988 297184 305000
rect 296888 304974 296934 304988
rect 296934 304974 296944 304988
rect 296968 304974 296998 304988
rect 296998 304974 297010 304988
rect 297010 304974 297024 304988
rect 297048 304974 297062 304988
rect 297062 304974 297074 304988
rect 297074 304974 297104 304988
rect 297128 304974 297138 304988
rect 297138 304974 297184 304988
rect 296888 304936 296934 304950
rect 296934 304936 296944 304950
rect 296968 304936 296998 304950
rect 296998 304936 297010 304950
rect 297010 304936 297024 304950
rect 297048 304936 297062 304950
rect 297062 304936 297074 304950
rect 297074 304936 297104 304950
rect 297128 304936 297138 304950
rect 297138 304936 297184 304950
rect 301686 304952 301742 305008
rect 303888 305000 303934 305030
rect 303934 305000 303944 305030
rect 303968 305000 303998 305030
rect 303998 305000 304010 305030
rect 304010 305000 304024 305030
rect 304048 305000 304062 305030
rect 304062 305000 304074 305030
rect 304074 305000 304104 305030
rect 304128 305000 304138 305030
rect 304138 305000 304184 305030
rect 310888 323862 310934 323908
rect 310934 323862 310944 323908
rect 310968 323862 310998 323908
rect 310998 323862 311010 323908
rect 311010 323862 311024 323908
rect 311048 323862 311062 323908
rect 311062 323862 311074 323908
rect 311074 323862 311104 323908
rect 311128 323862 311138 323908
rect 311138 323862 311184 323908
rect 310888 323852 310944 323862
rect 310968 323852 311024 323862
rect 311048 323852 311104 323862
rect 311128 323852 311184 323862
rect 310888 323798 310934 323828
rect 310934 323798 310944 323828
rect 310968 323798 310998 323828
rect 310998 323798 311010 323828
rect 311010 323798 311024 323828
rect 311048 323798 311062 323828
rect 311062 323798 311074 323828
rect 311074 323798 311104 323828
rect 311128 323798 311138 323828
rect 311138 323798 311184 323828
rect 310888 323786 310944 323798
rect 310968 323786 311024 323798
rect 311048 323786 311104 323798
rect 311128 323786 311184 323798
rect 310888 323772 310934 323786
rect 310934 323772 310944 323786
rect 310968 323772 310998 323786
rect 310998 323772 311010 323786
rect 311010 323772 311024 323786
rect 311048 323772 311062 323786
rect 311062 323772 311074 323786
rect 311074 323772 311104 323786
rect 311128 323772 311138 323786
rect 311138 323772 311184 323786
rect 310888 323734 310934 323748
rect 310934 323734 310944 323748
rect 310968 323734 310998 323748
rect 310998 323734 311010 323748
rect 311010 323734 311024 323748
rect 311048 323734 311062 323748
rect 311062 323734 311074 323748
rect 311074 323734 311104 323748
rect 311128 323734 311138 323748
rect 311138 323734 311184 323748
rect 310888 323722 310944 323734
rect 310968 323722 311024 323734
rect 311048 323722 311104 323734
rect 311128 323722 311184 323734
rect 310888 323692 310934 323722
rect 310934 323692 310944 323722
rect 310968 323692 310998 323722
rect 310998 323692 311010 323722
rect 311010 323692 311024 323722
rect 311048 323692 311062 323722
rect 311062 323692 311074 323722
rect 311074 323692 311104 323722
rect 311128 323692 311138 323722
rect 311138 323692 311184 323722
rect 310888 323658 310944 323668
rect 310968 323658 311024 323668
rect 311048 323658 311104 323668
rect 311128 323658 311184 323668
rect 310888 323612 310934 323658
rect 310934 323612 310944 323658
rect 310968 323612 310998 323658
rect 310998 323612 311010 323658
rect 311010 323612 311024 323658
rect 311048 323612 311062 323658
rect 311062 323612 311074 323658
rect 311074 323612 311104 323658
rect 311128 323612 311138 323658
rect 311138 323612 311184 323658
rect 311990 326168 312046 326224
rect 311898 307400 311954 307456
rect 314474 388456 314530 388512
rect 314566 386416 314622 386472
rect 314382 368872 314438 368928
rect 314014 366016 314070 366072
rect 312910 363024 312966 363080
rect 312634 342216 312690 342272
rect 312634 324944 312690 325000
rect 313738 307400 313794 307456
rect 312910 307128 312966 307184
rect 312542 306992 312598 307048
rect 311990 306448 312046 306504
rect 313646 306448 313702 306504
rect 310888 305064 310934 305110
rect 310934 305064 310944 305110
rect 310968 305064 310998 305110
rect 310998 305064 311010 305110
rect 311010 305064 311024 305110
rect 311048 305064 311062 305110
rect 311062 305064 311074 305110
rect 311074 305064 311104 305110
rect 311128 305064 311138 305110
rect 311138 305064 311184 305110
rect 310888 305054 310944 305064
rect 310968 305054 311024 305064
rect 311048 305054 311104 305064
rect 311128 305054 311184 305064
rect 303888 304988 303944 305000
rect 303968 304988 304024 305000
rect 304048 304988 304104 305000
rect 304128 304988 304184 305000
rect 303888 304974 303934 304988
rect 303934 304974 303944 304988
rect 303968 304974 303998 304988
rect 303998 304974 304010 304988
rect 304010 304974 304024 304988
rect 304048 304974 304062 304988
rect 304062 304974 304074 304988
rect 304074 304974 304104 304988
rect 304128 304974 304138 304988
rect 304138 304974 304184 304988
rect 296888 304924 296944 304936
rect 296968 304924 297024 304936
rect 297048 304924 297104 304936
rect 297128 304924 297184 304936
rect 296888 304894 296934 304924
rect 296934 304894 296944 304924
rect 296968 304894 296998 304924
rect 296998 304894 297010 304924
rect 297010 304894 297024 304924
rect 297048 304894 297062 304924
rect 297062 304894 297074 304924
rect 297074 304894 297104 304924
rect 297128 304894 297138 304924
rect 297138 304894 297184 304924
rect 296888 304860 296944 304870
rect 296968 304860 297024 304870
rect 297048 304860 297104 304870
rect 297128 304860 297184 304870
rect 296888 304814 296934 304860
rect 296934 304814 296944 304860
rect 296968 304814 296998 304860
rect 296998 304814 297010 304860
rect 297010 304814 297024 304860
rect 297048 304814 297062 304860
rect 297062 304814 297074 304860
rect 297074 304814 297104 304860
rect 297128 304814 297138 304860
rect 297138 304814 297184 304860
rect 303888 304936 303934 304950
rect 303934 304936 303944 304950
rect 303968 304936 303998 304950
rect 303998 304936 304010 304950
rect 304010 304936 304024 304950
rect 304048 304936 304062 304950
rect 304062 304936 304074 304950
rect 304074 304936 304104 304950
rect 304128 304936 304138 304950
rect 304138 304936 304184 304950
rect 306194 304952 306250 305008
rect 310610 304952 310666 305008
rect 310888 305000 310934 305030
rect 310934 305000 310944 305030
rect 310968 305000 310998 305030
rect 310998 305000 311010 305030
rect 311010 305000 311024 305030
rect 311048 305000 311062 305030
rect 311062 305000 311074 305030
rect 311074 305000 311104 305030
rect 311128 305000 311138 305030
rect 311138 305000 311184 305030
rect 310888 304988 310944 305000
rect 310968 304988 311024 305000
rect 311048 304988 311104 305000
rect 311128 304988 311184 305000
rect 310888 304974 310934 304988
rect 310934 304974 310944 304988
rect 310968 304974 310998 304988
rect 310998 304974 311010 304988
rect 311010 304974 311024 304988
rect 311048 304974 311062 304988
rect 311062 304974 311074 304988
rect 311074 304974 311104 304988
rect 311128 304974 311138 304988
rect 311138 304974 311184 304988
rect 303888 304924 303944 304936
rect 303968 304924 304024 304936
rect 304048 304924 304104 304936
rect 304128 304924 304184 304936
rect 303888 304894 303934 304924
rect 303934 304894 303944 304924
rect 303968 304894 303998 304924
rect 303998 304894 304010 304924
rect 304010 304894 304024 304924
rect 304048 304894 304062 304924
rect 304062 304894 304074 304924
rect 304074 304894 304104 304924
rect 304128 304894 304138 304924
rect 304138 304894 304184 304924
rect 303888 304860 303944 304870
rect 303968 304860 304024 304870
rect 304048 304860 304104 304870
rect 304128 304860 304184 304870
rect 303888 304814 303934 304860
rect 303934 304814 303944 304860
rect 303968 304814 303998 304860
rect 303998 304814 304010 304860
rect 304010 304814 304024 304860
rect 304048 304814 304062 304860
rect 304062 304814 304074 304860
rect 304074 304814 304104 304860
rect 304128 304814 304138 304860
rect 304138 304814 304184 304860
rect 310888 304936 310934 304950
rect 310934 304936 310944 304950
rect 310968 304936 310998 304950
rect 310998 304936 311010 304950
rect 311010 304936 311024 304950
rect 311048 304936 311062 304950
rect 311062 304936 311074 304950
rect 311074 304936 311104 304950
rect 311128 304936 311138 304950
rect 311138 304936 311184 304950
rect 310888 304924 310944 304936
rect 310968 304924 311024 304936
rect 311048 304924 311104 304936
rect 311128 304924 311184 304936
rect 310888 304894 310934 304924
rect 310934 304894 310944 304924
rect 310968 304894 310998 304924
rect 310998 304894 311010 304924
rect 311010 304894 311024 304924
rect 311048 304894 311062 304924
rect 311062 304894 311074 304924
rect 311074 304894 311104 304924
rect 311128 304894 311138 304924
rect 311138 304894 311184 304924
rect 310888 304860 310944 304870
rect 310968 304860 311024 304870
rect 311048 304860 311104 304870
rect 311128 304860 311184 304870
rect 310888 304814 310934 304860
rect 310934 304814 310944 304860
rect 310968 304814 310998 304860
rect 310998 304814 311010 304860
rect 311010 304814 311024 304860
rect 311048 304814 311062 304860
rect 311062 304814 311074 304860
rect 311074 304814 311104 304860
rect 311128 304814 311138 304860
rect 311138 304814 311184 304860
rect 301956 304544 302012 304600
rect 305550 304544 305606 304600
rect 312358 304544 312414 304600
rect 302156 303963 302202 304009
rect 302202 303963 302212 304009
rect 302236 303963 302266 304009
rect 302266 303963 302278 304009
rect 302278 303963 302292 304009
rect 302316 303963 302330 304009
rect 302330 303963 302342 304009
rect 302342 303963 302372 304009
rect 302396 303963 302406 304009
rect 302406 303963 302452 304009
rect 302156 303953 302212 303963
rect 302236 303953 302292 303963
rect 302316 303953 302372 303963
rect 302396 303953 302452 303963
rect 302156 303899 302202 303929
rect 302202 303899 302212 303929
rect 302236 303899 302266 303929
rect 302266 303899 302278 303929
rect 302278 303899 302292 303929
rect 302316 303899 302330 303929
rect 302330 303899 302342 303929
rect 302342 303899 302372 303929
rect 302396 303899 302406 303929
rect 302406 303899 302452 303929
rect 302156 303887 302212 303899
rect 302236 303887 302292 303899
rect 302316 303887 302372 303899
rect 302396 303887 302452 303899
rect 302156 303873 302202 303887
rect 302202 303873 302212 303887
rect 302236 303873 302266 303887
rect 302266 303873 302278 303887
rect 302278 303873 302292 303887
rect 302316 303873 302330 303887
rect 302330 303873 302342 303887
rect 302342 303873 302372 303887
rect 302396 303873 302406 303887
rect 302406 303873 302452 303887
rect 302156 303835 302202 303849
rect 302202 303835 302212 303849
rect 302236 303835 302266 303849
rect 302266 303835 302278 303849
rect 302278 303835 302292 303849
rect 302316 303835 302330 303849
rect 302330 303835 302342 303849
rect 302342 303835 302372 303849
rect 302396 303835 302406 303849
rect 302406 303835 302452 303849
rect 302156 303823 302212 303835
rect 302236 303823 302292 303835
rect 302316 303823 302372 303835
rect 302396 303823 302452 303835
rect 302156 303793 302202 303823
rect 302202 303793 302212 303823
rect 302236 303793 302266 303823
rect 302266 303793 302278 303823
rect 302278 303793 302292 303823
rect 302316 303793 302330 303823
rect 302330 303793 302342 303823
rect 302342 303793 302372 303823
rect 302396 303793 302406 303823
rect 302406 303793 302452 303823
rect 302156 303759 302212 303769
rect 302236 303759 302292 303769
rect 302316 303759 302372 303769
rect 302396 303759 302452 303769
rect 302156 303713 302202 303759
rect 302202 303713 302212 303759
rect 302236 303713 302266 303759
rect 302266 303713 302278 303759
rect 302278 303713 302292 303759
rect 302316 303713 302330 303759
rect 302330 303713 302342 303759
rect 302342 303713 302372 303759
rect 302396 303713 302406 303759
rect 302406 303713 302452 303759
rect 309156 303963 309202 304009
rect 309202 303963 309212 304009
rect 309236 303963 309266 304009
rect 309266 303963 309278 304009
rect 309278 303963 309292 304009
rect 309316 303963 309330 304009
rect 309330 303963 309342 304009
rect 309342 303963 309372 304009
rect 309396 303963 309406 304009
rect 309406 303963 309452 304009
rect 309156 303953 309212 303963
rect 309236 303953 309292 303963
rect 309316 303953 309372 303963
rect 309396 303953 309452 303963
rect 309156 303899 309202 303929
rect 309202 303899 309212 303929
rect 309236 303899 309266 303929
rect 309266 303899 309278 303929
rect 309278 303899 309292 303929
rect 309316 303899 309330 303929
rect 309330 303899 309342 303929
rect 309342 303899 309372 303929
rect 309396 303899 309406 303929
rect 309406 303899 309452 303929
rect 309156 303887 309212 303899
rect 309236 303887 309292 303899
rect 309316 303887 309372 303899
rect 309396 303887 309452 303899
rect 309156 303873 309202 303887
rect 309202 303873 309212 303887
rect 309236 303873 309266 303887
rect 309266 303873 309278 303887
rect 309278 303873 309292 303887
rect 309316 303873 309330 303887
rect 309330 303873 309342 303887
rect 309342 303873 309372 303887
rect 309396 303873 309406 303887
rect 309406 303873 309452 303887
rect 309156 303835 309202 303849
rect 309202 303835 309212 303849
rect 309236 303835 309266 303849
rect 309266 303835 309278 303849
rect 309278 303835 309292 303849
rect 309316 303835 309330 303849
rect 309330 303835 309342 303849
rect 309342 303835 309372 303849
rect 309396 303835 309406 303849
rect 309406 303835 309452 303849
rect 309156 303823 309212 303835
rect 309236 303823 309292 303835
rect 309316 303823 309372 303835
rect 309396 303823 309452 303835
rect 309156 303793 309202 303823
rect 309202 303793 309212 303823
rect 309236 303793 309266 303823
rect 309266 303793 309278 303823
rect 309278 303793 309292 303823
rect 309316 303793 309330 303823
rect 309330 303793 309342 303823
rect 309342 303793 309372 303823
rect 309396 303793 309406 303823
rect 309406 303793 309452 303823
rect 309156 303759 309212 303769
rect 309236 303759 309292 303769
rect 309316 303759 309372 303769
rect 309396 303759 309452 303769
rect 309156 303713 309202 303759
rect 309202 303713 309212 303759
rect 309236 303713 309266 303759
rect 309266 303713 309278 303759
rect 309278 303713 309292 303759
rect 309316 303713 309330 303759
rect 309330 303713 309342 303759
rect 309342 303713 309372 303759
rect 309396 303713 309406 303759
rect 309406 303713 309452 303759
rect 299202 301960 299258 302016
rect 306378 302096 306434 302152
rect 302790 301824 302846 301880
rect 295246 294480 295302 294536
rect 295246 284416 295302 284472
rect 299478 294480 299534 294536
rect 313370 303456 313426 303512
rect 309966 288768 310022 288824
rect 311898 288360 311954 288416
rect 313738 288360 313794 288416
rect 308126 285912 308182 285968
rect 304814 285776 304870 285832
rect 299478 284416 299534 284472
rect 295246 284280 295302 284336
rect 298098 284280 298154 284336
rect 312726 285912 312782 285968
rect 312358 285776 312414 285832
rect 299478 283736 299534 283792
rect 304814 283736 304870 283792
rect 308126 283736 308182 283792
rect 298142 283328 298198 283384
rect 299754 283328 299810 283384
rect 304776 283328 304832 283384
rect 308093 283328 308149 283384
rect 302156 282948 302202 282994
rect 302202 282948 302212 282994
rect 302236 282948 302266 282994
rect 302266 282948 302278 282994
rect 302278 282948 302292 282994
rect 302316 282948 302330 282994
rect 302330 282948 302342 282994
rect 302342 282948 302372 282994
rect 302396 282948 302406 282994
rect 302406 282948 302452 282994
rect 302156 282938 302212 282948
rect 302236 282938 302292 282948
rect 302316 282938 302372 282948
rect 302396 282938 302452 282948
rect 302156 282884 302202 282914
rect 302202 282884 302212 282914
rect 302236 282884 302266 282914
rect 302266 282884 302278 282914
rect 302278 282884 302292 282914
rect 302316 282884 302330 282914
rect 302330 282884 302342 282914
rect 302342 282884 302372 282914
rect 302396 282884 302406 282914
rect 302406 282884 302452 282914
rect 302156 282872 302212 282884
rect 302236 282872 302292 282884
rect 302316 282872 302372 282884
rect 302396 282872 302452 282884
rect 302156 282858 302202 282872
rect 302202 282858 302212 282872
rect 302236 282858 302266 282872
rect 302266 282858 302278 282872
rect 302278 282858 302292 282872
rect 302316 282858 302330 282872
rect 302330 282858 302342 282872
rect 302342 282858 302372 282872
rect 302396 282858 302406 282872
rect 302406 282858 302452 282872
rect 302156 282820 302202 282834
rect 302202 282820 302212 282834
rect 302236 282820 302266 282834
rect 302266 282820 302278 282834
rect 302278 282820 302292 282834
rect 302316 282820 302330 282834
rect 302330 282820 302342 282834
rect 302342 282820 302372 282834
rect 302396 282820 302406 282834
rect 302406 282820 302452 282834
rect 302156 282808 302212 282820
rect 302236 282808 302292 282820
rect 302316 282808 302372 282820
rect 302396 282808 302452 282820
rect 302156 282778 302202 282808
rect 302202 282778 302212 282808
rect 302236 282778 302266 282808
rect 302266 282778 302278 282808
rect 302278 282778 302292 282808
rect 302316 282778 302330 282808
rect 302330 282778 302342 282808
rect 302342 282778 302372 282808
rect 302396 282778 302406 282808
rect 302406 282778 302452 282808
rect 302156 282744 302212 282754
rect 302236 282744 302292 282754
rect 302316 282744 302372 282754
rect 302396 282744 302452 282754
rect 302156 282698 302202 282744
rect 302202 282698 302212 282744
rect 302236 282698 302266 282744
rect 302266 282698 302278 282744
rect 302278 282698 302292 282744
rect 302316 282698 302330 282744
rect 302330 282698 302342 282744
rect 302342 282698 302372 282744
rect 302396 282698 302406 282744
rect 302406 282698 302452 282744
rect 309156 282949 309202 282995
rect 309202 282949 309212 282995
rect 309236 282949 309266 282995
rect 309266 282949 309278 282995
rect 309278 282949 309292 282995
rect 309316 282949 309330 282995
rect 309330 282949 309342 282995
rect 309342 282949 309372 282995
rect 309396 282949 309406 282995
rect 309406 282949 309452 282995
rect 309156 282939 309212 282949
rect 309236 282939 309292 282949
rect 309316 282939 309372 282949
rect 309396 282939 309452 282949
rect 309156 282885 309202 282915
rect 309202 282885 309212 282915
rect 309236 282885 309266 282915
rect 309266 282885 309278 282915
rect 309278 282885 309292 282915
rect 309316 282885 309330 282915
rect 309330 282885 309342 282915
rect 309342 282885 309372 282915
rect 309396 282885 309406 282915
rect 309406 282885 309452 282915
rect 309156 282873 309212 282885
rect 309236 282873 309292 282885
rect 309316 282873 309372 282885
rect 309396 282873 309452 282885
rect 309156 282859 309202 282873
rect 309202 282859 309212 282873
rect 309236 282859 309266 282873
rect 309266 282859 309278 282873
rect 309278 282859 309292 282873
rect 309316 282859 309330 282873
rect 309330 282859 309342 282873
rect 309342 282859 309372 282873
rect 309396 282859 309406 282873
rect 309406 282859 309452 282873
rect 309156 282821 309202 282835
rect 309202 282821 309212 282835
rect 309236 282821 309266 282835
rect 309266 282821 309278 282835
rect 309278 282821 309292 282835
rect 309316 282821 309330 282835
rect 309330 282821 309342 282835
rect 309342 282821 309372 282835
rect 309396 282821 309406 282835
rect 309406 282821 309452 282835
rect 309156 282809 309212 282821
rect 309236 282809 309292 282821
rect 309316 282809 309372 282821
rect 309396 282809 309452 282821
rect 309156 282779 309202 282809
rect 309202 282779 309212 282809
rect 309236 282779 309266 282809
rect 309266 282779 309278 282809
rect 309278 282779 309292 282809
rect 309316 282779 309330 282809
rect 309330 282779 309342 282809
rect 309342 282779 309372 282809
rect 309396 282779 309406 282809
rect 309406 282779 309452 282809
rect 309156 282745 309212 282755
rect 309236 282745 309292 282755
rect 309316 282745 309372 282755
rect 309396 282745 309452 282755
rect 309156 282699 309202 282745
rect 309202 282699 309212 282745
rect 309236 282699 309266 282745
rect 309266 282699 309278 282745
rect 309278 282699 309292 282745
rect 309316 282699 309330 282745
rect 309330 282699 309342 282745
rect 309342 282699 309372 282745
rect 309396 282699 309406 282745
rect 309406 282699 309452 282745
rect 303888 282187 303934 282233
rect 303934 282187 303944 282233
rect 303968 282187 303998 282233
rect 303998 282187 304010 282233
rect 304010 282187 304024 282233
rect 304048 282187 304062 282233
rect 304062 282187 304074 282233
rect 304074 282187 304104 282233
rect 304128 282187 304138 282233
rect 304138 282187 304184 282233
rect 303888 282177 303944 282187
rect 303968 282177 304024 282187
rect 304048 282177 304104 282187
rect 304128 282177 304184 282187
rect 303888 282123 303934 282153
rect 303934 282123 303944 282153
rect 303968 282123 303998 282153
rect 303998 282123 304010 282153
rect 304010 282123 304024 282153
rect 304048 282123 304062 282153
rect 304062 282123 304074 282153
rect 304074 282123 304104 282153
rect 304128 282123 304138 282153
rect 304138 282123 304184 282153
rect 303888 282111 303944 282123
rect 303968 282111 304024 282123
rect 304048 282111 304104 282123
rect 304128 282111 304184 282123
rect 303888 282097 303934 282111
rect 303934 282097 303944 282111
rect 303968 282097 303998 282111
rect 303998 282097 304010 282111
rect 304010 282097 304024 282111
rect 304048 282097 304062 282111
rect 304062 282097 304074 282111
rect 304074 282097 304104 282111
rect 304128 282097 304138 282111
rect 304138 282097 304184 282111
rect 310888 282140 310934 282178
rect 310934 282140 310944 282178
rect 310968 282140 310998 282178
rect 310998 282140 311010 282178
rect 311010 282140 311024 282178
rect 311048 282140 311062 282178
rect 311062 282140 311074 282178
rect 311074 282140 311104 282178
rect 311128 282140 311138 282178
rect 311138 282140 311184 282178
rect 310888 282128 310944 282140
rect 310968 282128 311024 282140
rect 311048 282128 311104 282140
rect 311128 282128 311184 282140
rect 310888 282122 310934 282128
rect 310934 282122 310944 282128
rect 310968 282122 310998 282128
rect 310998 282122 311010 282128
rect 311010 282122 311024 282128
rect 311048 282122 311062 282128
rect 311062 282122 311074 282128
rect 311074 282122 311104 282128
rect 311128 282122 311138 282128
rect 311138 282122 311184 282128
rect 303888 282059 303934 282073
rect 303934 282059 303944 282073
rect 303968 282059 303998 282073
rect 303998 282059 304010 282073
rect 304010 282059 304024 282073
rect 304048 282059 304062 282073
rect 304062 282059 304074 282073
rect 304074 282059 304104 282073
rect 304128 282059 304138 282073
rect 304138 282059 304184 282073
rect 303888 282047 303944 282059
rect 303968 282047 304024 282059
rect 304048 282047 304104 282059
rect 304128 282047 304184 282059
rect 303888 282017 303934 282047
rect 303934 282017 303944 282047
rect 303968 282017 303998 282047
rect 303998 282017 304010 282047
rect 304010 282017 304024 282047
rect 304048 282017 304062 282047
rect 304062 282017 304074 282047
rect 304074 282017 304104 282047
rect 304128 282017 304138 282047
rect 304138 282017 304184 282047
rect 299110 281288 299166 281344
rect 310888 282076 310934 282098
rect 310934 282076 310944 282098
rect 310968 282076 310998 282098
rect 310998 282076 311010 282098
rect 311010 282076 311024 282098
rect 311048 282076 311062 282098
rect 311062 282076 311074 282098
rect 311074 282076 311104 282098
rect 311128 282076 311138 282098
rect 311138 282076 311184 282098
rect 310888 282064 310944 282076
rect 310968 282064 311024 282076
rect 311048 282064 311104 282076
rect 311128 282064 311184 282076
rect 310888 282042 310934 282064
rect 310934 282042 310944 282064
rect 310968 282042 310998 282064
rect 310998 282042 311010 282064
rect 311010 282042 311024 282064
rect 311048 282042 311062 282064
rect 311062 282042 311074 282064
rect 311074 282042 311104 282064
rect 311128 282042 311138 282064
rect 311138 282042 311184 282064
rect 303888 281983 303944 281993
rect 303968 281983 304024 281993
rect 304048 281983 304104 281993
rect 304128 281983 304184 281993
rect 303888 281937 303934 281983
rect 303934 281937 303944 281983
rect 303968 281937 303998 281983
rect 303998 281937 304010 281983
rect 304010 281937 304024 281983
rect 304048 281937 304062 281983
rect 304062 281937 304074 281983
rect 304074 281937 304104 281983
rect 304128 281937 304138 281983
rect 304138 281937 304184 281983
rect 303888 281867 303934 281913
rect 303934 281867 303944 281913
rect 303968 281867 303998 281913
rect 303998 281867 304010 281913
rect 304010 281867 304024 281913
rect 304048 281867 304062 281913
rect 304062 281867 304074 281913
rect 304074 281867 304104 281913
rect 304128 281867 304138 281913
rect 304138 281867 304184 281913
rect 303888 281857 303944 281867
rect 303968 281857 304024 281867
rect 304048 281857 304104 281867
rect 304128 281857 304184 281867
rect 303888 281803 303934 281833
rect 303934 281803 303944 281833
rect 303968 281803 303998 281833
rect 303998 281803 304010 281833
rect 304010 281803 304024 281833
rect 304048 281803 304062 281833
rect 304062 281803 304074 281833
rect 304074 281803 304104 281833
rect 304128 281803 304138 281833
rect 304138 281803 304184 281833
rect 303888 281791 303944 281803
rect 303968 281791 304024 281803
rect 304048 281791 304104 281803
rect 304128 281791 304184 281803
rect 303888 281777 303934 281791
rect 303934 281777 303944 281791
rect 303968 281777 303998 281791
rect 303998 281777 304010 281791
rect 304010 281777 304024 281791
rect 304048 281777 304062 281791
rect 304062 281777 304074 281791
rect 304074 281777 304104 281791
rect 304128 281777 304138 281791
rect 304138 281777 304184 281791
rect 303888 281739 303934 281753
rect 303934 281739 303944 281753
rect 303968 281739 303998 281753
rect 303998 281739 304010 281753
rect 304010 281739 304024 281753
rect 304048 281739 304062 281753
rect 304062 281739 304074 281753
rect 304074 281739 304104 281753
rect 304128 281739 304138 281753
rect 304138 281739 304184 281753
rect 303888 281727 303944 281739
rect 303968 281727 304024 281739
rect 304048 281727 304104 281739
rect 304128 281727 304184 281739
rect 303888 281697 303934 281727
rect 303934 281697 303944 281727
rect 303968 281697 303998 281727
rect 303998 281697 304010 281727
rect 304010 281697 304024 281727
rect 304048 281697 304062 281727
rect 304062 281697 304074 281727
rect 304074 281697 304104 281727
rect 304128 281697 304138 281727
rect 304138 281697 304184 281727
rect 303888 281663 303944 281673
rect 303968 281663 304024 281673
rect 304048 281663 304104 281673
rect 304128 281663 304184 281673
rect 303888 281617 303934 281663
rect 303934 281617 303944 281663
rect 303968 281617 303998 281663
rect 303998 281617 304010 281663
rect 304010 281617 304024 281663
rect 304048 281617 304062 281663
rect 304062 281617 304074 281663
rect 304074 281617 304104 281663
rect 304128 281617 304138 281663
rect 304138 281617 304184 281663
rect 305734 281424 305790 281480
rect 310888 282012 310934 282018
rect 310934 282012 310944 282018
rect 310968 282012 310998 282018
rect 310998 282012 311010 282018
rect 311010 282012 311024 282018
rect 311048 282012 311062 282018
rect 311062 282012 311074 282018
rect 311074 282012 311104 282018
rect 311128 282012 311138 282018
rect 311138 282012 311184 282018
rect 310888 282000 310944 282012
rect 310968 282000 311024 282012
rect 311048 282000 311104 282012
rect 311128 282000 311184 282012
rect 310888 281962 310934 282000
rect 310934 281962 310944 282000
rect 310968 281962 310998 282000
rect 310998 281962 311010 282000
rect 311010 281962 311024 282000
rect 311048 281962 311062 282000
rect 311062 281962 311074 282000
rect 311074 281962 311104 282000
rect 311128 281962 311138 282000
rect 311138 281962 311184 282000
rect 310888 281936 310944 281938
rect 310968 281936 311024 281938
rect 311048 281936 311104 281938
rect 311128 281936 311184 281938
rect 310888 281884 310934 281936
rect 310934 281884 310944 281936
rect 310968 281884 310998 281936
rect 310998 281884 311010 281936
rect 311010 281884 311024 281936
rect 311048 281884 311062 281936
rect 311062 281884 311074 281936
rect 311074 281884 311104 281936
rect 311128 281884 311138 281936
rect 311138 281884 311184 281936
rect 310888 281882 310944 281884
rect 310968 281882 311024 281884
rect 311048 281882 311104 281884
rect 311128 281882 311184 281884
rect 310888 281820 310934 281858
rect 310934 281820 310944 281858
rect 310968 281820 310998 281858
rect 310998 281820 311010 281858
rect 311010 281820 311024 281858
rect 311048 281820 311062 281858
rect 311062 281820 311074 281858
rect 311074 281820 311104 281858
rect 311128 281820 311138 281858
rect 311138 281820 311184 281858
rect 310888 281808 310944 281820
rect 310968 281808 311024 281820
rect 311048 281808 311104 281820
rect 311128 281808 311184 281820
rect 310888 281802 310934 281808
rect 310934 281802 310944 281808
rect 310968 281802 310998 281808
rect 310998 281802 311010 281808
rect 311010 281802 311024 281808
rect 311048 281802 311062 281808
rect 311062 281802 311074 281808
rect 311074 281802 311104 281808
rect 311128 281802 311138 281808
rect 311138 281802 311184 281808
rect 310888 281756 310934 281778
rect 310934 281756 310944 281778
rect 310968 281756 310998 281778
rect 310998 281756 311010 281778
rect 311010 281756 311024 281778
rect 311048 281756 311062 281778
rect 311062 281756 311074 281778
rect 311074 281756 311104 281778
rect 311128 281756 311138 281778
rect 311138 281756 311184 281778
rect 310888 281744 310944 281756
rect 310968 281744 311024 281756
rect 311048 281744 311104 281756
rect 311128 281744 311184 281756
rect 310888 281722 310934 281744
rect 310934 281722 310944 281744
rect 310968 281722 310998 281744
rect 310998 281722 311010 281744
rect 311010 281722 311024 281744
rect 311048 281722 311062 281744
rect 311062 281722 311074 281744
rect 311074 281722 311104 281744
rect 311128 281722 311138 281744
rect 311138 281722 311184 281744
rect 310888 281692 310934 281698
rect 310934 281692 310944 281698
rect 310968 281692 310998 281698
rect 310998 281692 311010 281698
rect 311010 281692 311024 281698
rect 311048 281692 311062 281698
rect 311062 281692 311074 281698
rect 311074 281692 311104 281698
rect 311128 281692 311138 281698
rect 311138 281692 311184 281698
rect 310888 281680 310944 281692
rect 310968 281680 311024 281692
rect 311048 281680 311104 281692
rect 311128 281680 311184 281692
rect 310888 281642 310934 281680
rect 310934 281642 310944 281680
rect 310968 281642 310998 281680
rect 310998 281642 311010 281680
rect 311010 281642 311024 281680
rect 311048 281642 311062 281680
rect 311062 281642 311074 281680
rect 311074 281642 311104 281680
rect 311128 281642 311138 281680
rect 311138 281642 311184 281680
rect 308954 280064 309010 280120
rect 302422 279928 302478 279984
rect 295246 277480 295302 277536
rect 298190 277480 298246 277536
rect 295246 264968 295302 265024
rect 295154 262792 295210 262848
rect 308770 265104 308826 265160
rect 299478 264968 299534 265024
rect 305090 264968 305146 265024
rect 298190 262792 298246 262848
rect 312634 285640 312690 285696
rect 312542 282004 312544 282024
rect 312544 282004 312596 282024
rect 312596 282004 312598 282024
rect 312542 281968 312598 282004
rect 313830 285640 313886 285696
rect 312358 264968 312414 265024
rect 312542 264968 312598 265024
rect 302156 261948 302202 261994
rect 302202 261948 302212 261994
rect 302236 261948 302266 261994
rect 302266 261948 302278 261994
rect 302278 261948 302292 261994
rect 302316 261948 302330 261994
rect 302330 261948 302342 261994
rect 302342 261948 302372 261994
rect 302396 261948 302406 261994
rect 302406 261948 302452 261994
rect 302156 261938 302212 261948
rect 302236 261938 302292 261948
rect 302316 261938 302372 261948
rect 302396 261938 302452 261948
rect 302156 261884 302202 261914
rect 302202 261884 302212 261914
rect 302236 261884 302266 261914
rect 302266 261884 302278 261914
rect 302278 261884 302292 261914
rect 302316 261884 302330 261914
rect 302330 261884 302342 261914
rect 302342 261884 302372 261914
rect 302396 261884 302406 261914
rect 302406 261884 302452 261914
rect 302156 261872 302212 261884
rect 302236 261872 302292 261884
rect 302316 261872 302372 261884
rect 302396 261872 302452 261884
rect 302156 261858 302202 261872
rect 302202 261858 302212 261872
rect 302236 261858 302266 261872
rect 302266 261858 302278 261872
rect 302278 261858 302292 261872
rect 302316 261858 302330 261872
rect 302330 261858 302342 261872
rect 302342 261858 302372 261872
rect 302396 261858 302406 261872
rect 302406 261858 302452 261872
rect 302156 261820 302202 261834
rect 302202 261820 302212 261834
rect 302236 261820 302266 261834
rect 302266 261820 302278 261834
rect 302278 261820 302292 261834
rect 302316 261820 302330 261834
rect 302330 261820 302342 261834
rect 302342 261820 302372 261834
rect 302396 261820 302406 261834
rect 302406 261820 302452 261834
rect 302156 261808 302212 261820
rect 302236 261808 302292 261820
rect 302316 261808 302372 261820
rect 302396 261808 302452 261820
rect 302156 261778 302202 261808
rect 302202 261778 302212 261808
rect 302236 261778 302266 261808
rect 302266 261778 302278 261808
rect 302278 261778 302292 261808
rect 302316 261778 302330 261808
rect 302330 261778 302342 261808
rect 302342 261778 302372 261808
rect 302396 261778 302406 261808
rect 302406 261778 302452 261808
rect 302156 261744 302212 261754
rect 302236 261744 302292 261754
rect 302316 261744 302372 261754
rect 302396 261744 302452 261754
rect 302156 261698 302202 261744
rect 302202 261698 302212 261744
rect 302236 261698 302266 261744
rect 302266 261698 302278 261744
rect 302278 261698 302292 261744
rect 302316 261698 302330 261744
rect 302330 261698 302342 261744
rect 302342 261698 302372 261744
rect 302396 261698 302406 261744
rect 302406 261698 302452 261744
rect 309156 261948 309202 261994
rect 309202 261948 309212 261994
rect 309236 261948 309266 261994
rect 309266 261948 309278 261994
rect 309278 261948 309292 261994
rect 309316 261948 309330 261994
rect 309330 261948 309342 261994
rect 309342 261948 309372 261994
rect 309396 261948 309406 261994
rect 309406 261948 309452 261994
rect 309156 261938 309212 261948
rect 309236 261938 309292 261948
rect 309316 261938 309372 261948
rect 309396 261938 309452 261948
rect 309156 261884 309202 261914
rect 309202 261884 309212 261914
rect 309236 261884 309266 261914
rect 309266 261884 309278 261914
rect 309278 261884 309292 261914
rect 309316 261884 309330 261914
rect 309330 261884 309342 261914
rect 309342 261884 309372 261914
rect 309396 261884 309406 261914
rect 309406 261884 309452 261914
rect 309156 261872 309212 261884
rect 309236 261872 309292 261884
rect 309316 261872 309372 261884
rect 309396 261872 309452 261884
rect 309156 261858 309202 261872
rect 309202 261858 309212 261872
rect 309236 261858 309266 261872
rect 309266 261858 309278 261872
rect 309278 261858 309292 261872
rect 309316 261858 309330 261872
rect 309330 261858 309342 261872
rect 309342 261858 309372 261872
rect 309396 261858 309406 261872
rect 309406 261858 309452 261872
rect 309156 261820 309202 261834
rect 309202 261820 309212 261834
rect 309236 261820 309266 261834
rect 309266 261820 309278 261834
rect 309278 261820 309292 261834
rect 309316 261820 309330 261834
rect 309330 261820 309342 261834
rect 309342 261820 309372 261834
rect 309396 261820 309406 261834
rect 309406 261820 309452 261834
rect 309156 261808 309212 261820
rect 309236 261808 309292 261820
rect 309316 261808 309372 261820
rect 309396 261808 309452 261820
rect 309156 261778 309202 261808
rect 309202 261778 309212 261808
rect 309236 261778 309266 261808
rect 309266 261778 309278 261808
rect 309278 261778 309292 261808
rect 309316 261778 309330 261808
rect 309330 261778 309342 261808
rect 309342 261778 309372 261808
rect 309396 261778 309406 261808
rect 309406 261778 309452 261808
rect 309156 261744 309212 261754
rect 309236 261744 309292 261754
rect 309316 261744 309372 261754
rect 309396 261744 309452 261754
rect 309156 261698 309202 261744
rect 309202 261698 309212 261744
rect 309236 261698 309266 261744
rect 309266 261698 309278 261744
rect 309278 261698 309292 261744
rect 309316 261698 309330 261744
rect 309330 261698 309342 261744
rect 309342 261698 309372 261744
rect 309396 261698 309406 261744
rect 309406 261698 309452 261744
rect 303888 261187 303934 261233
rect 303934 261187 303944 261233
rect 303968 261187 303998 261233
rect 303998 261187 304010 261233
rect 304010 261187 304024 261233
rect 304048 261187 304062 261233
rect 304062 261187 304074 261233
rect 304074 261187 304104 261233
rect 304128 261187 304138 261233
rect 304138 261187 304184 261233
rect 303888 261177 303944 261187
rect 303968 261177 304024 261187
rect 304048 261177 304104 261187
rect 304128 261177 304184 261187
rect 303888 261123 303934 261153
rect 303934 261123 303944 261153
rect 303968 261123 303998 261153
rect 303998 261123 304010 261153
rect 304010 261123 304024 261153
rect 304048 261123 304062 261153
rect 304062 261123 304074 261153
rect 304074 261123 304104 261153
rect 304128 261123 304138 261153
rect 304138 261123 304184 261153
rect 303888 261111 303944 261123
rect 303968 261111 304024 261123
rect 304048 261111 304104 261123
rect 304128 261111 304184 261123
rect 303888 261097 303934 261111
rect 303934 261097 303944 261111
rect 303968 261097 303998 261111
rect 303998 261097 304010 261111
rect 304010 261097 304024 261111
rect 304048 261097 304062 261111
rect 304062 261097 304074 261111
rect 304074 261097 304104 261111
rect 304128 261097 304138 261111
rect 304138 261097 304184 261111
rect 303888 261059 303934 261073
rect 303934 261059 303944 261073
rect 303968 261059 303998 261073
rect 303998 261059 304010 261073
rect 304010 261059 304024 261073
rect 304048 261059 304062 261073
rect 304062 261059 304074 261073
rect 304074 261059 304104 261073
rect 304128 261059 304138 261073
rect 304138 261059 304184 261073
rect 303888 261047 303944 261059
rect 303968 261047 304024 261059
rect 304048 261047 304104 261059
rect 304128 261047 304184 261059
rect 303888 261017 303934 261047
rect 303934 261017 303944 261047
rect 303968 261017 303998 261047
rect 303998 261017 304010 261047
rect 304010 261017 304024 261047
rect 304048 261017 304062 261047
rect 304062 261017 304074 261047
rect 304074 261017 304104 261047
rect 304128 261017 304138 261047
rect 304138 261017 304184 261047
rect 299018 259256 299074 259312
rect 303888 260983 303944 260993
rect 303968 260983 304024 260993
rect 304048 260983 304104 260993
rect 304128 260983 304184 260993
rect 303888 260937 303934 260983
rect 303934 260937 303944 260983
rect 303968 260937 303998 260983
rect 303998 260937 304010 260983
rect 304010 260937 304024 260983
rect 304048 260937 304062 260983
rect 304062 260937 304074 260983
rect 304074 260937 304104 260983
rect 304128 260937 304138 260983
rect 304138 260937 304184 260983
rect 303888 260867 303934 260913
rect 303934 260867 303944 260913
rect 303968 260867 303998 260913
rect 303998 260867 304010 260913
rect 304010 260867 304024 260913
rect 304048 260867 304062 260913
rect 304062 260867 304074 260913
rect 304074 260867 304104 260913
rect 304128 260867 304138 260913
rect 304138 260867 304184 260913
rect 303888 260857 303944 260867
rect 303968 260857 304024 260867
rect 304048 260857 304104 260867
rect 304128 260857 304184 260867
rect 303888 260803 303934 260833
rect 303934 260803 303944 260833
rect 303968 260803 303998 260833
rect 303998 260803 304010 260833
rect 304010 260803 304024 260833
rect 304048 260803 304062 260833
rect 304062 260803 304074 260833
rect 304074 260803 304104 260833
rect 304128 260803 304138 260833
rect 304138 260803 304184 260833
rect 303888 260791 303944 260803
rect 303968 260791 304024 260803
rect 304048 260791 304104 260803
rect 304128 260791 304184 260803
rect 303888 260777 303934 260791
rect 303934 260777 303944 260791
rect 303968 260777 303998 260791
rect 303998 260777 304010 260791
rect 304010 260777 304024 260791
rect 304048 260777 304062 260791
rect 304062 260777 304074 260791
rect 304074 260777 304104 260791
rect 304128 260777 304138 260791
rect 304138 260777 304184 260791
rect 303888 260739 303934 260753
rect 303934 260739 303944 260753
rect 303968 260739 303998 260753
rect 303998 260739 304010 260753
rect 304010 260739 304024 260753
rect 304048 260739 304062 260753
rect 304062 260739 304074 260753
rect 304074 260739 304104 260753
rect 304128 260739 304138 260753
rect 304138 260739 304184 260753
rect 303888 260727 303944 260739
rect 303968 260727 304024 260739
rect 304048 260727 304104 260739
rect 304128 260727 304184 260739
rect 303888 260697 303934 260727
rect 303934 260697 303944 260727
rect 303968 260697 303998 260727
rect 303998 260697 304010 260727
rect 304010 260697 304024 260727
rect 304048 260697 304062 260727
rect 304062 260697 304074 260727
rect 304074 260697 304104 260727
rect 304128 260697 304138 260727
rect 304138 260697 304184 260727
rect 303888 260663 303944 260673
rect 303968 260663 304024 260673
rect 304048 260663 304104 260673
rect 304128 260663 304184 260673
rect 303888 260617 303934 260663
rect 303934 260617 303944 260663
rect 303968 260617 303998 260663
rect 303998 260617 304010 260663
rect 304010 260617 304024 260663
rect 304048 260617 304062 260663
rect 304062 260617 304074 260663
rect 304074 260617 304104 260663
rect 304128 260617 304138 260663
rect 304138 260617 304184 260663
rect 309506 260616 309562 260672
rect 305918 260480 305974 260536
rect 309506 259392 309562 259448
rect 302606 259120 302662 259176
rect 312818 261568 312874 261624
rect 295246 243480 295302 243536
rect 300858 243480 300914 243536
rect 296888 242034 296934 242080
rect 296934 242034 296944 242080
rect 296968 242034 296998 242080
rect 296998 242034 297010 242080
rect 297010 242034 297024 242080
rect 297048 242034 297062 242080
rect 297062 242034 297074 242080
rect 297074 242034 297104 242080
rect 297128 242034 297138 242080
rect 297138 242034 297184 242080
rect 296888 242024 296944 242034
rect 296968 242024 297024 242034
rect 297048 242024 297104 242034
rect 297128 242024 297184 242034
rect 296888 241970 296934 242000
rect 296934 241970 296944 242000
rect 296968 241970 296998 242000
rect 296998 241970 297010 242000
rect 297010 241970 297024 242000
rect 297048 241970 297062 242000
rect 297062 241970 297074 242000
rect 297074 241970 297104 242000
rect 297128 241970 297138 242000
rect 297138 241970 297184 242000
rect 296888 241958 296944 241970
rect 296968 241958 297024 241970
rect 297048 241958 297104 241970
rect 297128 241958 297184 241970
rect 296888 241944 296934 241958
rect 296934 241944 296944 241958
rect 296968 241944 296998 241958
rect 296998 241944 297010 241958
rect 297010 241944 297024 241958
rect 297048 241944 297062 241958
rect 297062 241944 297074 241958
rect 297074 241944 297104 241958
rect 297128 241944 297138 241958
rect 297138 241944 297184 241958
rect 296888 241906 296934 241920
rect 296934 241906 296944 241920
rect 296968 241906 296998 241920
rect 296998 241906 297010 241920
rect 297010 241906 297024 241920
rect 297048 241906 297062 241920
rect 297062 241906 297074 241920
rect 297074 241906 297104 241920
rect 297128 241906 297138 241920
rect 297138 241906 297184 241920
rect 304630 243344 304686 243400
rect 312082 243344 312138 243400
rect 303888 242034 303934 242080
rect 303934 242034 303944 242080
rect 303968 242034 303998 242080
rect 303998 242034 304010 242080
rect 304010 242034 304024 242080
rect 304048 242034 304062 242080
rect 304062 242034 304074 242080
rect 304074 242034 304104 242080
rect 304128 242034 304138 242080
rect 304138 242034 304184 242080
rect 303888 242024 303944 242034
rect 303968 242024 304024 242034
rect 304048 242024 304104 242034
rect 304128 242024 304184 242034
rect 303888 241970 303934 242000
rect 303934 241970 303944 242000
rect 303968 241970 303998 242000
rect 303998 241970 304010 242000
rect 304010 241970 304024 242000
rect 304048 241970 304062 242000
rect 304062 241970 304074 242000
rect 304074 241970 304104 242000
rect 304128 241970 304138 242000
rect 304138 241970 304184 242000
rect 303888 241958 303944 241970
rect 303968 241958 304024 241970
rect 304048 241958 304104 241970
rect 304128 241958 304184 241970
rect 303888 241944 303934 241958
rect 303934 241944 303944 241958
rect 303968 241944 303998 241958
rect 303998 241944 304010 241958
rect 304010 241944 304024 241958
rect 304048 241944 304062 241958
rect 304062 241944 304074 241958
rect 304074 241944 304104 241958
rect 304128 241944 304138 241958
rect 304138 241944 304184 241958
rect 296888 241894 296944 241906
rect 296968 241894 297024 241906
rect 297048 241894 297104 241906
rect 297128 241894 297184 241906
rect 296888 241864 296934 241894
rect 296934 241864 296944 241894
rect 296968 241864 296998 241894
rect 296998 241864 297010 241894
rect 297010 241864 297024 241894
rect 297048 241864 297062 241894
rect 297062 241864 297074 241894
rect 297074 241864 297104 241894
rect 297128 241864 297138 241894
rect 297138 241864 297184 241894
rect 296888 241830 296944 241840
rect 296968 241830 297024 241840
rect 297048 241830 297104 241840
rect 297128 241830 297184 241840
rect 300858 241848 300914 241904
rect 303888 241906 303934 241920
rect 303934 241906 303944 241920
rect 303968 241906 303998 241920
rect 303998 241906 304010 241920
rect 304010 241906 304024 241920
rect 304048 241906 304062 241920
rect 304062 241906 304074 241920
rect 304074 241906 304104 241920
rect 304128 241906 304138 241920
rect 304138 241906 304184 241920
rect 310888 242034 310934 242080
rect 310934 242034 310944 242080
rect 310968 242034 310998 242080
rect 310998 242034 311010 242080
rect 311010 242034 311024 242080
rect 311048 242034 311062 242080
rect 311062 242034 311074 242080
rect 311074 242034 311104 242080
rect 311128 242034 311138 242080
rect 311138 242034 311184 242080
rect 310888 242024 310944 242034
rect 310968 242024 311024 242034
rect 311048 242024 311104 242034
rect 311128 242024 311184 242034
rect 310888 241970 310934 242000
rect 310934 241970 310944 242000
rect 310968 241970 310998 242000
rect 310998 241970 311010 242000
rect 311010 241970 311024 242000
rect 311048 241970 311062 242000
rect 311062 241970 311074 242000
rect 311074 241970 311104 242000
rect 311128 241970 311138 242000
rect 311138 241970 311184 242000
rect 310888 241958 310944 241970
rect 310968 241958 311024 241970
rect 311048 241958 311104 241970
rect 311128 241958 311184 241970
rect 310888 241944 310934 241958
rect 310934 241944 310944 241958
rect 310968 241944 310998 241958
rect 310998 241944 311010 241958
rect 311010 241944 311024 241958
rect 311048 241944 311062 241958
rect 311062 241944 311074 241958
rect 311074 241944 311104 241958
rect 311128 241944 311138 241958
rect 311138 241944 311184 241958
rect 303888 241894 303944 241906
rect 303968 241894 304024 241906
rect 304048 241894 304104 241906
rect 304128 241894 304184 241906
rect 303888 241864 303934 241894
rect 303934 241864 303944 241894
rect 303968 241864 303998 241894
rect 303998 241864 304010 241894
rect 304010 241864 304024 241894
rect 304048 241864 304062 241894
rect 304062 241864 304074 241894
rect 304074 241864 304104 241894
rect 304128 241864 304138 241894
rect 304138 241864 304184 241894
rect 296888 241784 296934 241830
rect 296934 241784 296944 241830
rect 296968 241784 296998 241830
rect 296998 241784 297010 241830
rect 297010 241784 297024 241830
rect 297048 241784 297062 241830
rect 297062 241784 297074 241830
rect 297074 241784 297104 241830
rect 297128 241784 297138 241830
rect 297138 241784 297184 241830
rect 303888 241830 303944 241840
rect 303968 241830 304024 241840
rect 304048 241830 304104 241840
rect 304128 241830 304184 241840
rect 304630 241848 304686 241904
rect 310888 241906 310934 241920
rect 310934 241906 310944 241920
rect 310968 241906 310998 241920
rect 310998 241906 311010 241920
rect 311010 241906 311024 241920
rect 311048 241906 311062 241920
rect 311062 241906 311074 241920
rect 311074 241906 311104 241920
rect 311128 241906 311138 241920
rect 311138 241906 311184 241920
rect 310888 241894 310944 241906
rect 310968 241894 311024 241906
rect 311048 241894 311104 241906
rect 311128 241894 311184 241906
rect 310888 241864 310934 241894
rect 310934 241864 310944 241894
rect 310968 241864 310998 241894
rect 310998 241864 311010 241894
rect 311010 241864 311024 241894
rect 311048 241864 311062 241894
rect 311062 241864 311074 241894
rect 311074 241864 311104 241894
rect 311128 241864 311138 241894
rect 311138 241864 311184 241894
rect 303888 241784 303934 241830
rect 303934 241784 303944 241830
rect 303968 241784 303998 241830
rect 303998 241784 304010 241830
rect 304010 241784 304024 241830
rect 304048 241784 304062 241830
rect 304062 241784 304074 241830
rect 304074 241784 304104 241830
rect 304128 241784 304138 241830
rect 304138 241784 304184 241830
rect 310888 241830 310944 241840
rect 310968 241830 311024 241840
rect 311048 241830 311104 241840
rect 311128 241830 311184 241840
rect 310888 241784 310934 241830
rect 310934 241784 310944 241830
rect 310968 241784 310998 241830
rect 310998 241784 311010 241830
rect 311010 241784 311024 241830
rect 311048 241784 311062 241830
rect 311062 241784 311074 241830
rect 311074 241784 311104 241830
rect 311128 241784 311138 241830
rect 311138 241784 311184 241830
rect 300950 241576 301006 241632
rect 304548 241440 304604 241496
rect 295156 240949 295202 240995
rect 295202 240949 295212 240995
rect 295236 240949 295266 240995
rect 295266 240949 295278 240995
rect 295278 240949 295292 240995
rect 295316 240949 295330 240995
rect 295330 240949 295342 240995
rect 295342 240949 295372 240995
rect 295396 240949 295406 240995
rect 295406 240949 295452 240995
rect 295156 240939 295212 240949
rect 295236 240939 295292 240949
rect 295316 240939 295372 240949
rect 295396 240939 295452 240949
rect 295156 240885 295202 240915
rect 295202 240885 295212 240915
rect 295236 240885 295266 240915
rect 295266 240885 295278 240915
rect 295278 240885 295292 240915
rect 295316 240885 295330 240915
rect 295330 240885 295342 240915
rect 295342 240885 295372 240915
rect 295396 240885 295406 240915
rect 295406 240885 295452 240915
rect 295156 240873 295212 240885
rect 295236 240873 295292 240885
rect 295316 240873 295372 240885
rect 295396 240873 295452 240885
rect 295156 240859 295202 240873
rect 295202 240859 295212 240873
rect 295236 240859 295266 240873
rect 295266 240859 295278 240873
rect 295278 240859 295292 240873
rect 295316 240859 295330 240873
rect 295330 240859 295342 240873
rect 295342 240859 295372 240873
rect 295396 240859 295406 240873
rect 295406 240859 295452 240873
rect 295156 240821 295202 240835
rect 295202 240821 295212 240835
rect 295236 240821 295266 240835
rect 295266 240821 295278 240835
rect 295278 240821 295292 240835
rect 295316 240821 295330 240835
rect 295330 240821 295342 240835
rect 295342 240821 295372 240835
rect 295396 240821 295406 240835
rect 295406 240821 295452 240835
rect 295156 240809 295212 240821
rect 295236 240809 295292 240821
rect 295316 240809 295372 240821
rect 295396 240809 295452 240821
rect 295156 240779 295202 240809
rect 295202 240779 295212 240809
rect 295236 240779 295266 240809
rect 295266 240779 295278 240809
rect 295278 240779 295292 240809
rect 295316 240779 295330 240809
rect 295330 240779 295342 240809
rect 295342 240779 295372 240809
rect 295396 240779 295406 240809
rect 295406 240779 295452 240809
rect 295156 240745 295212 240755
rect 295236 240745 295292 240755
rect 295316 240745 295372 240755
rect 295396 240745 295452 240755
rect 295156 240699 295202 240745
rect 295202 240699 295212 240745
rect 295236 240699 295266 240745
rect 295266 240699 295278 240745
rect 295278 240699 295292 240745
rect 295316 240699 295330 240745
rect 295330 240699 295342 240745
rect 295342 240699 295372 240745
rect 295396 240699 295406 240745
rect 295406 240699 295452 240745
rect 309156 240923 309202 240969
rect 309202 240923 309212 240969
rect 309236 240923 309266 240969
rect 309266 240923 309278 240969
rect 309278 240923 309292 240969
rect 309316 240923 309330 240969
rect 309330 240923 309342 240969
rect 309342 240923 309372 240969
rect 309396 240923 309406 240969
rect 309406 240923 309452 240969
rect 309156 240913 309212 240923
rect 309236 240913 309292 240923
rect 309316 240913 309372 240923
rect 309396 240913 309452 240923
rect 309156 240859 309202 240889
rect 309202 240859 309212 240889
rect 309236 240859 309266 240889
rect 309266 240859 309278 240889
rect 309278 240859 309292 240889
rect 309316 240859 309330 240889
rect 309330 240859 309342 240889
rect 309342 240859 309372 240889
rect 309396 240859 309406 240889
rect 309406 240859 309452 240889
rect 309156 240847 309212 240859
rect 309236 240847 309292 240859
rect 309316 240847 309372 240859
rect 309396 240847 309452 240859
rect 309156 240833 309202 240847
rect 309202 240833 309212 240847
rect 309236 240833 309266 240847
rect 309266 240833 309278 240847
rect 309278 240833 309292 240847
rect 309316 240833 309330 240847
rect 309330 240833 309342 240847
rect 309342 240833 309372 240847
rect 309396 240833 309406 240847
rect 309406 240833 309452 240847
rect 309156 240795 309202 240809
rect 309202 240795 309212 240809
rect 309236 240795 309266 240809
rect 309266 240795 309278 240809
rect 309278 240795 309292 240809
rect 309316 240795 309330 240809
rect 309330 240795 309342 240809
rect 309342 240795 309372 240809
rect 309396 240795 309406 240809
rect 309406 240795 309452 240809
rect 309156 240783 309212 240795
rect 309236 240783 309292 240795
rect 309316 240783 309372 240795
rect 309396 240783 309452 240795
rect 309156 240753 309202 240783
rect 309202 240753 309212 240783
rect 309236 240753 309266 240783
rect 309266 240753 309278 240783
rect 309278 240753 309292 240783
rect 309316 240753 309330 240783
rect 309330 240753 309342 240783
rect 309342 240753 309372 240783
rect 309396 240753 309406 240783
rect 309406 240753 309452 240783
rect 309156 240719 309212 240729
rect 309236 240719 309292 240729
rect 309316 240719 309372 240729
rect 309396 240719 309452 240729
rect 309156 240673 309202 240719
rect 309202 240673 309212 240719
rect 309236 240673 309266 240719
rect 309266 240673 309278 240719
rect 309278 240673 309292 240719
rect 309316 240673 309330 240719
rect 309330 240673 309342 240719
rect 309342 240673 309372 240719
rect 309396 240673 309406 240719
rect 309406 240673 309452 240719
rect 294878 222400 294934 222456
rect 295062 221176 295118 221232
rect 294970 202816 295026 202872
rect 294878 202136 294934 202192
rect 296888 221035 296934 221081
rect 296934 221035 296944 221081
rect 296968 221035 296998 221081
rect 296998 221035 297010 221081
rect 297010 221035 297024 221081
rect 297048 221035 297062 221081
rect 297062 221035 297074 221081
rect 297074 221035 297104 221081
rect 297128 221035 297138 221081
rect 297138 221035 297184 221081
rect 296888 221025 296944 221035
rect 296968 221025 297024 221035
rect 297048 221025 297104 221035
rect 297128 221025 297184 221035
rect 296888 220971 296934 221001
rect 296934 220971 296944 221001
rect 296968 220971 296998 221001
rect 296998 220971 297010 221001
rect 297010 220971 297024 221001
rect 297048 220971 297062 221001
rect 297062 220971 297074 221001
rect 297074 220971 297104 221001
rect 297128 220971 297138 221001
rect 297138 220971 297184 221001
rect 296888 220959 296944 220971
rect 296968 220959 297024 220971
rect 297048 220959 297104 220971
rect 297128 220959 297184 220971
rect 310888 239862 310934 239908
rect 310934 239862 310944 239908
rect 310968 239862 310998 239908
rect 310998 239862 311010 239908
rect 311010 239862 311024 239908
rect 311048 239862 311062 239908
rect 311062 239862 311074 239908
rect 311074 239862 311104 239908
rect 311128 239862 311138 239908
rect 311138 239862 311184 239908
rect 310888 239852 310944 239862
rect 310968 239852 311024 239862
rect 311048 239852 311104 239862
rect 311128 239852 311184 239862
rect 310888 239798 310934 239828
rect 310934 239798 310944 239828
rect 310968 239798 310998 239828
rect 310998 239798 311010 239828
rect 311010 239798 311024 239828
rect 311048 239798 311062 239828
rect 311062 239798 311074 239828
rect 311074 239798 311104 239828
rect 311128 239798 311138 239828
rect 311138 239798 311184 239828
rect 310888 239786 310944 239798
rect 310968 239786 311024 239798
rect 311048 239786 311104 239798
rect 311128 239786 311184 239798
rect 310888 239772 310934 239786
rect 310934 239772 310944 239786
rect 310968 239772 310998 239786
rect 310998 239772 311010 239786
rect 311010 239772 311024 239786
rect 311048 239772 311062 239786
rect 311062 239772 311074 239786
rect 311074 239772 311104 239786
rect 311128 239772 311138 239786
rect 311138 239772 311184 239786
rect 310888 239734 310934 239748
rect 310934 239734 310944 239748
rect 310968 239734 310998 239748
rect 310998 239734 311010 239748
rect 311010 239734 311024 239748
rect 311048 239734 311062 239748
rect 311062 239734 311074 239748
rect 311074 239734 311104 239748
rect 311128 239734 311138 239748
rect 311138 239734 311184 239748
rect 310888 239722 310944 239734
rect 310968 239722 311024 239734
rect 311048 239722 311104 239734
rect 311128 239722 311184 239734
rect 310888 239692 310934 239722
rect 310934 239692 310944 239722
rect 310968 239692 310998 239722
rect 310998 239692 311010 239722
rect 311010 239692 311024 239722
rect 311048 239692 311062 239722
rect 311062 239692 311074 239722
rect 311074 239692 311104 239722
rect 311128 239692 311138 239722
rect 311138 239692 311184 239722
rect 310888 239658 310944 239668
rect 310968 239658 311024 239668
rect 311048 239658 311104 239668
rect 311128 239658 311184 239668
rect 310888 239612 310934 239658
rect 310934 239612 310944 239658
rect 310968 239612 310998 239658
rect 310998 239612 311010 239658
rect 311010 239612 311024 239658
rect 311048 239612 311062 239658
rect 311062 239612 311074 239658
rect 311074 239612 311104 239658
rect 311128 239612 311138 239658
rect 311138 239612 311184 239658
rect 309874 222672 309930 222728
rect 305734 222400 305790 222456
rect 303888 221035 303934 221081
rect 303934 221035 303944 221081
rect 303968 221035 303998 221081
rect 303998 221035 304010 221081
rect 304010 221035 304024 221081
rect 304048 221035 304062 221081
rect 304062 221035 304074 221081
rect 304074 221035 304104 221081
rect 304128 221035 304138 221081
rect 304138 221035 304184 221081
rect 303888 221025 303944 221035
rect 303968 221025 304024 221035
rect 304048 221025 304104 221035
rect 304128 221025 304184 221035
rect 303888 220971 303934 221001
rect 303934 220971 303944 221001
rect 303968 220971 303998 221001
rect 303998 220971 304010 221001
rect 304010 220971 304024 221001
rect 304048 220971 304062 221001
rect 304062 220971 304074 221001
rect 304074 220971 304104 221001
rect 304128 220971 304138 221001
rect 304138 220971 304184 221001
rect 296888 220945 296934 220959
rect 296934 220945 296944 220959
rect 296968 220945 296998 220959
rect 296998 220945 297010 220959
rect 297010 220945 297024 220959
rect 297048 220945 297062 220959
rect 297062 220945 297074 220959
rect 297074 220945 297104 220959
rect 297128 220945 297138 220959
rect 297138 220945 297184 220959
rect 296888 220907 296934 220921
rect 296934 220907 296944 220921
rect 296968 220907 296998 220921
rect 296998 220907 297010 220921
rect 297010 220907 297024 220921
rect 297048 220907 297062 220921
rect 297062 220907 297074 220921
rect 297074 220907 297104 220921
rect 297128 220907 297138 220921
rect 297138 220907 297184 220921
rect 296888 220895 296944 220907
rect 296968 220895 297024 220907
rect 297048 220895 297104 220907
rect 297128 220895 297184 220907
rect 301318 220904 301374 220960
rect 303888 220959 303944 220971
rect 303968 220959 304024 220971
rect 304048 220959 304104 220971
rect 304128 220959 304184 220971
rect 313278 264968 313334 265024
rect 312910 243344 312966 243400
rect 314106 345072 314162 345128
rect 314014 259120 314070 259176
rect 314198 323040 314254 323096
rect 314106 251504 314162 251560
rect 314198 250144 314254 250200
rect 314474 285912 314530 285968
rect 315486 428984 315542 429040
rect 315394 403416 315450 403472
rect 315302 258304 315358 258360
rect 312542 222672 312598 222728
rect 312082 222264 312138 222320
rect 310888 221035 310934 221081
rect 310934 221035 310944 221081
rect 310968 221035 310998 221081
rect 310998 221035 311010 221081
rect 311010 221035 311024 221081
rect 311048 221035 311062 221081
rect 311062 221035 311074 221081
rect 311074 221035 311104 221081
rect 311128 221035 311138 221081
rect 311138 221035 311184 221081
rect 310888 221025 310944 221035
rect 310968 221025 311024 221035
rect 311048 221025 311104 221035
rect 311128 221025 311184 221035
rect 310888 220971 310934 221001
rect 310934 220971 310944 221001
rect 310968 220971 310998 221001
rect 310998 220971 311010 221001
rect 311010 220971 311024 221001
rect 311048 220971 311062 221001
rect 311062 220971 311074 221001
rect 311074 220971 311104 221001
rect 311128 220971 311138 221001
rect 311138 220971 311184 221001
rect 303888 220945 303934 220959
rect 303934 220945 303944 220959
rect 303968 220945 303998 220959
rect 303998 220945 304010 220959
rect 304010 220945 304024 220959
rect 304048 220945 304062 220959
rect 304062 220945 304074 220959
rect 304074 220945 304104 220959
rect 304128 220945 304138 220959
rect 304138 220945 304184 220959
rect 303888 220907 303934 220921
rect 303934 220907 303944 220921
rect 303968 220907 303998 220921
rect 303998 220907 304010 220921
rect 304010 220907 304024 220921
rect 304048 220907 304062 220921
rect 304062 220907 304074 220921
rect 304074 220907 304104 220921
rect 304128 220907 304138 220921
rect 304138 220907 304184 220921
rect 303888 220895 303944 220907
rect 303968 220895 304024 220907
rect 304048 220895 304104 220907
rect 304128 220895 304184 220907
rect 305734 220904 305790 220960
rect 309874 220904 309930 220960
rect 310888 220959 310944 220971
rect 310968 220959 311024 220971
rect 311048 220959 311104 220971
rect 311128 220959 311184 220971
rect 310888 220945 310934 220959
rect 310934 220945 310944 220959
rect 310968 220945 310998 220959
rect 310998 220945 311010 220959
rect 311010 220945 311024 220959
rect 311048 220945 311062 220959
rect 311062 220945 311074 220959
rect 311074 220945 311104 220959
rect 311128 220945 311138 220959
rect 311138 220945 311184 220959
rect 310888 220907 310934 220921
rect 310934 220907 310944 220921
rect 310968 220907 310998 220921
rect 310998 220907 311010 220921
rect 311010 220907 311024 220921
rect 311048 220907 311062 220921
rect 311062 220907 311074 220921
rect 311074 220907 311104 220921
rect 311128 220907 311138 220921
rect 311138 220907 311184 220921
rect 310888 220895 310944 220907
rect 310968 220895 311024 220907
rect 311048 220895 311104 220907
rect 311128 220895 311184 220907
rect 296888 220865 296934 220895
rect 296934 220865 296944 220895
rect 296968 220865 296998 220895
rect 296998 220865 297010 220895
rect 297010 220865 297024 220895
rect 297048 220865 297062 220895
rect 297062 220865 297074 220895
rect 297074 220865 297104 220895
rect 297128 220865 297138 220895
rect 297138 220865 297184 220895
rect 296888 220831 296944 220841
rect 296968 220831 297024 220841
rect 297048 220831 297104 220841
rect 297128 220831 297184 220841
rect 296888 220785 296934 220831
rect 296934 220785 296944 220831
rect 296968 220785 296998 220831
rect 296998 220785 297010 220831
rect 297010 220785 297024 220831
rect 297048 220785 297062 220831
rect 297062 220785 297074 220831
rect 297074 220785 297104 220831
rect 297128 220785 297138 220831
rect 297138 220785 297184 220831
rect 303888 220865 303934 220895
rect 303934 220865 303944 220895
rect 303968 220865 303998 220895
rect 303998 220865 304010 220895
rect 304010 220865 304024 220895
rect 304048 220865 304062 220895
rect 304062 220865 304074 220895
rect 304074 220865 304104 220895
rect 304128 220865 304138 220895
rect 304138 220865 304184 220895
rect 303888 220831 303944 220841
rect 303968 220831 304024 220841
rect 304048 220831 304104 220841
rect 304128 220831 304184 220841
rect 303888 220785 303934 220831
rect 303934 220785 303944 220831
rect 303968 220785 303998 220831
rect 303998 220785 304010 220831
rect 304010 220785 304024 220831
rect 304048 220785 304062 220831
rect 304062 220785 304074 220831
rect 304074 220785 304104 220831
rect 304128 220785 304138 220831
rect 304138 220785 304184 220831
rect 310888 220865 310934 220895
rect 310934 220865 310944 220895
rect 310968 220865 310998 220895
rect 310998 220865 311010 220895
rect 311010 220865 311024 220895
rect 311048 220865 311062 220895
rect 311062 220865 311074 220895
rect 311074 220865 311104 220895
rect 311128 220865 311138 220895
rect 311138 220865 311184 220895
rect 310888 220831 310944 220841
rect 310968 220831 311024 220841
rect 311048 220831 311104 220841
rect 311128 220831 311184 220841
rect 310888 220785 310934 220831
rect 310934 220785 310944 220831
rect 310968 220785 310998 220831
rect 310998 220785 311010 220831
rect 311010 220785 311024 220831
rect 311048 220785 311062 220831
rect 311062 220785 311074 220831
rect 311074 220785 311104 220831
rect 311128 220785 311138 220831
rect 311138 220785 311184 220831
rect 301870 220632 301926 220688
rect 305734 220632 305790 220688
rect 309690 220632 309746 220688
rect 295156 219950 295202 219996
rect 295202 219950 295212 219996
rect 295236 219950 295266 219996
rect 295266 219950 295278 219996
rect 295278 219950 295292 219996
rect 295316 219950 295330 219996
rect 295330 219950 295342 219996
rect 295342 219950 295372 219996
rect 295396 219950 295406 219996
rect 295406 219950 295452 219996
rect 295156 219940 295212 219950
rect 295236 219940 295292 219950
rect 295316 219940 295372 219950
rect 295396 219940 295452 219950
rect 295156 219886 295202 219916
rect 295202 219886 295212 219916
rect 295236 219886 295266 219916
rect 295266 219886 295278 219916
rect 295278 219886 295292 219916
rect 295316 219886 295330 219916
rect 295330 219886 295342 219916
rect 295342 219886 295372 219916
rect 295396 219886 295406 219916
rect 295406 219886 295452 219916
rect 295156 219874 295212 219886
rect 295236 219874 295292 219886
rect 295316 219874 295372 219886
rect 295396 219874 295452 219886
rect 295156 219860 295202 219874
rect 295202 219860 295212 219874
rect 295236 219860 295266 219874
rect 295266 219860 295278 219874
rect 295278 219860 295292 219874
rect 295316 219860 295330 219874
rect 295330 219860 295342 219874
rect 295342 219860 295372 219874
rect 295396 219860 295406 219874
rect 295406 219860 295452 219874
rect 295156 219822 295202 219836
rect 295202 219822 295212 219836
rect 295236 219822 295266 219836
rect 295266 219822 295278 219836
rect 295278 219822 295292 219836
rect 295316 219822 295330 219836
rect 295330 219822 295342 219836
rect 295342 219822 295372 219836
rect 295396 219822 295406 219836
rect 295406 219822 295452 219836
rect 295156 219810 295212 219822
rect 295236 219810 295292 219822
rect 295316 219810 295372 219822
rect 295396 219810 295452 219822
rect 295156 219780 295202 219810
rect 295202 219780 295212 219810
rect 295236 219780 295266 219810
rect 295266 219780 295278 219810
rect 295278 219780 295292 219810
rect 295316 219780 295330 219810
rect 295330 219780 295342 219810
rect 295342 219780 295372 219810
rect 295396 219780 295406 219810
rect 295406 219780 295452 219810
rect 295156 219746 295212 219756
rect 295236 219746 295292 219756
rect 295316 219746 295372 219756
rect 295396 219746 295452 219756
rect 295156 219700 295202 219746
rect 295202 219700 295212 219746
rect 295236 219700 295266 219746
rect 295266 219700 295278 219746
rect 295278 219700 295292 219746
rect 295316 219700 295330 219746
rect 295330 219700 295342 219746
rect 295342 219700 295372 219746
rect 295396 219700 295406 219746
rect 295406 219700 295452 219746
rect 302156 219949 302202 219995
rect 302202 219949 302212 219995
rect 302236 219949 302266 219995
rect 302266 219949 302278 219995
rect 302278 219949 302292 219995
rect 302316 219949 302330 219995
rect 302330 219949 302342 219995
rect 302342 219949 302372 219995
rect 302396 219949 302406 219995
rect 302406 219949 302452 219995
rect 302156 219939 302212 219949
rect 302236 219939 302292 219949
rect 302316 219939 302372 219949
rect 302396 219939 302452 219949
rect 302156 219885 302202 219915
rect 302202 219885 302212 219915
rect 302236 219885 302266 219915
rect 302266 219885 302278 219915
rect 302278 219885 302292 219915
rect 302316 219885 302330 219915
rect 302330 219885 302342 219915
rect 302342 219885 302372 219915
rect 302396 219885 302406 219915
rect 302406 219885 302452 219915
rect 302156 219873 302212 219885
rect 302236 219873 302292 219885
rect 302316 219873 302372 219885
rect 302396 219873 302452 219885
rect 302156 219859 302202 219873
rect 302202 219859 302212 219873
rect 302236 219859 302266 219873
rect 302266 219859 302278 219873
rect 302278 219859 302292 219873
rect 302316 219859 302330 219873
rect 302330 219859 302342 219873
rect 302342 219859 302372 219873
rect 302396 219859 302406 219873
rect 302406 219859 302452 219873
rect 302156 219821 302202 219835
rect 302202 219821 302212 219835
rect 302236 219821 302266 219835
rect 302266 219821 302278 219835
rect 302278 219821 302292 219835
rect 302316 219821 302330 219835
rect 302330 219821 302342 219835
rect 302342 219821 302372 219835
rect 302396 219821 302406 219835
rect 302406 219821 302452 219835
rect 302156 219809 302212 219821
rect 302236 219809 302292 219821
rect 302316 219809 302372 219821
rect 302396 219809 302452 219821
rect 302156 219779 302202 219809
rect 302202 219779 302212 219809
rect 302236 219779 302266 219809
rect 302266 219779 302278 219809
rect 302278 219779 302292 219809
rect 302316 219779 302330 219809
rect 302330 219779 302342 219809
rect 302342 219779 302372 219809
rect 302396 219779 302406 219809
rect 302406 219779 302452 219809
rect 302156 219745 302212 219755
rect 302236 219745 302292 219755
rect 302316 219745 302372 219755
rect 302396 219745 302452 219755
rect 302156 219699 302202 219745
rect 302202 219699 302212 219745
rect 302236 219699 302266 219745
rect 302266 219699 302278 219745
rect 302278 219699 302292 219745
rect 302316 219699 302330 219745
rect 302330 219699 302342 219745
rect 302342 219699 302372 219745
rect 302396 219699 302406 219745
rect 302406 219699 302452 219745
rect 309156 219949 309202 219995
rect 309202 219949 309212 219995
rect 309236 219949 309266 219995
rect 309266 219949 309278 219995
rect 309278 219949 309292 219995
rect 309316 219949 309330 219995
rect 309330 219949 309342 219995
rect 309342 219949 309372 219995
rect 309396 219949 309406 219995
rect 309406 219949 309452 219995
rect 309156 219939 309212 219949
rect 309236 219939 309292 219949
rect 309316 219939 309372 219949
rect 309396 219939 309452 219949
rect 309156 219885 309202 219915
rect 309202 219885 309212 219915
rect 309236 219885 309266 219915
rect 309266 219885 309278 219915
rect 309278 219885 309292 219915
rect 309316 219885 309330 219915
rect 309330 219885 309342 219915
rect 309342 219885 309372 219915
rect 309396 219885 309406 219915
rect 309406 219885 309452 219915
rect 309156 219873 309212 219885
rect 309236 219873 309292 219885
rect 309316 219873 309372 219885
rect 309396 219873 309452 219885
rect 309156 219859 309202 219873
rect 309202 219859 309212 219873
rect 309236 219859 309266 219873
rect 309266 219859 309278 219873
rect 309278 219859 309292 219873
rect 309316 219859 309330 219873
rect 309330 219859 309342 219873
rect 309342 219859 309372 219873
rect 309396 219859 309406 219873
rect 309406 219859 309452 219873
rect 309156 219821 309202 219835
rect 309202 219821 309212 219835
rect 309236 219821 309266 219835
rect 309266 219821 309278 219835
rect 309278 219821 309292 219835
rect 309316 219821 309330 219835
rect 309330 219821 309342 219835
rect 309342 219821 309372 219835
rect 309396 219821 309406 219835
rect 309406 219821 309452 219835
rect 309156 219809 309212 219821
rect 309236 219809 309292 219821
rect 309316 219809 309372 219821
rect 309396 219809 309452 219821
rect 309156 219779 309202 219809
rect 309202 219779 309212 219809
rect 309236 219779 309266 219809
rect 309266 219779 309278 219809
rect 309278 219779 309292 219809
rect 309316 219779 309330 219809
rect 309330 219779 309342 219809
rect 309342 219779 309372 219809
rect 309396 219779 309406 219809
rect 309406 219779 309452 219809
rect 309156 219745 309212 219755
rect 309236 219745 309292 219755
rect 309316 219745 309372 219755
rect 309396 219745 309452 219755
rect 309156 219699 309202 219745
rect 309202 219699 309212 219745
rect 309236 219699 309266 219745
rect 309266 219699 309278 219745
rect 309278 219699 309292 219745
rect 309316 219699 309330 219745
rect 309330 219699 309342 219745
rect 309342 219699 309372 219745
rect 309396 219699 309406 219745
rect 309406 219699 309452 219745
rect 303963 219396 304019 219398
rect 303963 219344 303965 219396
rect 303965 219344 304017 219396
rect 304017 219344 304019 219396
rect 303963 219342 304019 219344
rect 299294 217776 299350 217832
rect 303158 217504 303214 217560
rect 311043 219513 311099 219515
rect 311043 219461 311045 219513
rect 311045 219461 311097 219513
rect 311097 219461 311099 219513
rect 311043 219459 311099 219461
rect 307666 217912 307722 217968
rect 309598 217912 309654 217968
rect 306746 217368 306802 217424
rect 295246 202816 295302 202872
rect 295062 201456 295118 201512
rect 303618 202136 303674 202192
rect 300858 201456 300914 201512
rect 303618 201456 303674 201512
rect 310426 217776 310482 217832
rect 317050 408856 317106 408912
rect 315578 407904 315634 407960
rect 315486 256944 315542 257000
rect 315762 407496 315818 407552
rect 315670 406136 315726 406192
rect 316774 402056 316830 402112
rect 316682 400696 316738 400752
rect 315762 281288 315818 281344
rect 315762 261568 315818 261624
rect 315670 259256 315726 259312
rect 315578 255584 315634 255640
rect 315762 246064 315818 246120
rect 315394 217912 315450 217968
rect 310426 216688 310482 216744
rect 313922 216688 313978 216744
rect 307666 200232 307722 200288
rect 311162 201456 311218 201512
rect 300858 199824 300914 199880
rect 303618 199824 303674 199880
rect 300858 199552 300914 199608
rect 303710 199552 303766 199608
rect 307574 199552 307630 199608
rect 295062 181328 295118 181384
rect 304722 197240 304778 197296
rect 301686 197104 301742 197160
rect 298650 195744 298706 195800
rect 304446 181328 304502 181384
rect 300858 181056 300914 181112
rect 297270 180920 297326 180976
rect 295246 180784 295302 180840
rect 296888 179235 296934 179281
rect 296934 179235 296944 179281
rect 296968 179235 296998 179281
rect 296998 179235 297010 179281
rect 297010 179235 297024 179281
rect 297048 179235 297062 179281
rect 297062 179235 297074 179281
rect 297074 179235 297104 179281
rect 297128 179235 297138 179281
rect 297138 179235 297184 179281
rect 296888 179225 296944 179235
rect 296968 179225 297024 179235
rect 297048 179225 297104 179235
rect 297128 179225 297184 179235
rect 296888 179171 296934 179201
rect 296934 179171 296944 179201
rect 296968 179171 296998 179201
rect 296998 179171 297010 179201
rect 297010 179171 297024 179201
rect 297048 179171 297062 179201
rect 297062 179171 297074 179201
rect 297074 179171 297104 179201
rect 297128 179171 297138 179201
rect 297138 179171 297184 179201
rect 296888 179159 296944 179171
rect 296968 179159 297024 179171
rect 297048 179159 297104 179171
rect 297128 179159 297184 179171
rect 296888 179145 296934 179159
rect 296934 179145 296944 179159
rect 296968 179145 296998 179159
rect 296998 179145 297010 179159
rect 297010 179145 297024 179159
rect 297048 179145 297062 179159
rect 297062 179145 297074 179159
rect 297074 179145 297104 179159
rect 297128 179145 297138 179159
rect 297138 179145 297184 179159
rect 296888 179107 296934 179121
rect 296934 179107 296944 179121
rect 296968 179107 296998 179121
rect 296998 179107 297010 179121
rect 297010 179107 297024 179121
rect 297048 179107 297062 179121
rect 297062 179107 297074 179121
rect 297074 179107 297104 179121
rect 297128 179107 297138 179121
rect 297138 179107 297184 179121
rect 296888 179095 296944 179107
rect 296968 179095 297024 179107
rect 297048 179095 297104 179107
rect 297128 179095 297184 179107
rect 296888 179065 296934 179095
rect 296934 179065 296944 179095
rect 296968 179065 296998 179095
rect 296998 179065 297010 179095
rect 297010 179065 297024 179095
rect 297048 179065 297062 179095
rect 297062 179065 297074 179095
rect 297074 179065 297104 179095
rect 297128 179065 297138 179095
rect 297138 179065 297184 179095
rect 303888 179235 303934 179281
rect 303934 179235 303944 179281
rect 303968 179235 303998 179281
rect 303998 179235 304010 179281
rect 304010 179235 304024 179281
rect 304048 179235 304062 179281
rect 304062 179235 304074 179281
rect 304074 179235 304104 179281
rect 304128 179235 304138 179281
rect 304138 179235 304184 179281
rect 303888 179225 303944 179235
rect 303968 179225 304024 179235
rect 304048 179225 304104 179235
rect 304128 179225 304184 179235
rect 303888 179171 303934 179201
rect 303934 179171 303944 179201
rect 303968 179171 303998 179201
rect 303998 179171 304010 179201
rect 304010 179171 304024 179201
rect 304048 179171 304062 179201
rect 304062 179171 304074 179201
rect 304074 179171 304104 179201
rect 304128 179171 304138 179201
rect 304138 179171 304184 179201
rect 303888 179159 303944 179171
rect 303968 179159 304024 179171
rect 304048 179159 304104 179171
rect 304128 179159 304184 179171
rect 303888 179145 303934 179159
rect 303934 179145 303944 179159
rect 303968 179145 303998 179159
rect 303998 179145 304010 179159
rect 304010 179145 304024 179159
rect 304048 179145 304062 179159
rect 304062 179145 304074 179159
rect 304074 179145 304104 179159
rect 304128 179145 304138 179159
rect 304138 179145 304184 179159
rect 303888 179107 303934 179121
rect 303934 179107 303944 179121
rect 303968 179107 303998 179121
rect 303998 179107 304010 179121
rect 304010 179107 304024 179121
rect 304048 179107 304062 179121
rect 304062 179107 304074 179121
rect 304074 179107 304104 179121
rect 304128 179107 304138 179121
rect 304138 179107 304184 179121
rect 303888 179095 303944 179107
rect 303968 179095 304024 179107
rect 304048 179095 304104 179107
rect 304128 179095 304184 179107
rect 296888 179031 296944 179041
rect 296968 179031 297024 179041
rect 297048 179031 297104 179041
rect 297128 179031 297184 179041
rect 296888 178985 296934 179031
rect 296934 178985 296944 179031
rect 296968 178985 296998 179031
rect 296998 178985 297010 179031
rect 297010 178985 297024 179031
rect 297048 178985 297062 179031
rect 297062 178985 297074 179031
rect 297074 178985 297104 179031
rect 297128 178985 297138 179031
rect 297138 178985 297184 179031
rect 297270 179016 297326 179072
rect 300858 179016 300914 179072
rect 303888 179065 303934 179095
rect 303934 179065 303944 179095
rect 303968 179065 303998 179095
rect 303998 179065 304010 179095
rect 304010 179065 304024 179095
rect 304048 179065 304062 179095
rect 304062 179065 304074 179095
rect 304074 179065 304104 179095
rect 304128 179065 304138 179095
rect 304138 179065 304184 179095
rect 307758 195880 307814 195936
rect 311162 181328 311218 181384
rect 311162 180920 311218 180976
rect 307666 179424 307722 179480
rect 310892 179235 310894 179281
rect 310894 179235 310946 179281
rect 310946 179235 310948 179281
rect 310892 179225 310948 179235
rect 310892 179171 310894 179201
rect 310894 179171 310946 179201
rect 310946 179171 310948 179201
rect 310892 179159 310948 179171
rect 310892 179145 310894 179159
rect 310894 179145 310946 179159
rect 310946 179145 310948 179159
rect 310892 179107 310894 179121
rect 310894 179107 310946 179121
rect 310946 179107 310948 179121
rect 310892 179095 310948 179107
rect 303888 179031 303944 179041
rect 303968 179031 304024 179041
rect 304048 179031 304104 179041
rect 304128 179031 304184 179041
rect 303888 178985 303934 179031
rect 303934 178985 303944 179031
rect 303968 178985 303998 179031
rect 303998 178985 304010 179031
rect 304010 178985 304024 179031
rect 304048 178985 304062 179031
rect 304062 178985 304074 179031
rect 304074 178985 304104 179031
rect 304128 178985 304138 179031
rect 304138 178985 304184 179031
rect 304446 179016 304502 179072
rect 310892 179065 310894 179095
rect 310894 179065 310946 179095
rect 310946 179065 310948 179095
rect 310892 179031 310948 179041
rect 310892 178985 310894 179031
rect 310894 178985 310946 179031
rect 310946 178985 310948 179031
rect 297270 178744 297326 178800
rect 300857 178744 300913 178800
rect 303909 178744 303965 178800
rect 307114 178744 307170 178800
rect 295156 178149 295202 178195
rect 295202 178149 295212 178195
rect 295236 178149 295266 178195
rect 295266 178149 295278 178195
rect 295278 178149 295292 178195
rect 295316 178149 295330 178195
rect 295330 178149 295342 178195
rect 295342 178149 295372 178195
rect 295396 178149 295406 178195
rect 295406 178149 295452 178195
rect 295156 178139 295212 178149
rect 295236 178139 295292 178149
rect 295316 178139 295372 178149
rect 295396 178139 295452 178149
rect 295156 178085 295202 178115
rect 295202 178085 295212 178115
rect 295236 178085 295266 178115
rect 295266 178085 295278 178115
rect 295278 178085 295292 178115
rect 295316 178085 295330 178115
rect 295330 178085 295342 178115
rect 295342 178085 295372 178115
rect 295396 178085 295406 178115
rect 295406 178085 295452 178115
rect 295156 178073 295212 178085
rect 295236 178073 295292 178085
rect 295316 178073 295372 178085
rect 295396 178073 295452 178085
rect 295156 178059 295202 178073
rect 295202 178059 295212 178073
rect 295236 178059 295266 178073
rect 295266 178059 295278 178073
rect 295278 178059 295292 178073
rect 295316 178059 295330 178073
rect 295330 178059 295342 178073
rect 295342 178059 295372 178073
rect 295396 178059 295406 178073
rect 295406 178059 295452 178073
rect 295156 178021 295202 178035
rect 295202 178021 295212 178035
rect 295236 178021 295266 178035
rect 295266 178021 295278 178035
rect 295278 178021 295292 178035
rect 295316 178021 295330 178035
rect 295330 178021 295342 178035
rect 295342 178021 295372 178035
rect 295396 178021 295406 178035
rect 295406 178021 295452 178035
rect 295156 178009 295212 178021
rect 295236 178009 295292 178021
rect 295316 178009 295372 178021
rect 295396 178009 295452 178021
rect 295156 177979 295202 178009
rect 295202 177979 295212 178009
rect 295236 177979 295266 178009
rect 295266 177979 295278 178009
rect 295278 177979 295292 178009
rect 295316 177979 295330 178009
rect 295330 177979 295342 178009
rect 295342 177979 295372 178009
rect 295396 177979 295406 178009
rect 295406 177979 295452 178009
rect 295156 177945 295212 177955
rect 295236 177945 295292 177955
rect 295316 177945 295372 177955
rect 295396 177945 295452 177955
rect 295156 177899 295202 177945
rect 295202 177899 295212 177945
rect 295236 177899 295266 177945
rect 295266 177899 295278 177945
rect 295278 177899 295292 177945
rect 295316 177899 295330 177945
rect 295330 177899 295342 177945
rect 295342 177899 295372 177945
rect 295396 177899 295406 177945
rect 295406 177899 295452 177945
rect 302156 178133 302202 178179
rect 302202 178133 302212 178179
rect 302236 178133 302266 178179
rect 302266 178133 302278 178179
rect 302278 178133 302292 178179
rect 302316 178133 302330 178179
rect 302330 178133 302342 178179
rect 302342 178133 302372 178179
rect 302396 178133 302406 178179
rect 302406 178133 302452 178179
rect 302156 178123 302212 178133
rect 302236 178123 302292 178133
rect 302316 178123 302372 178133
rect 302396 178123 302452 178133
rect 302156 178069 302202 178099
rect 302202 178069 302212 178099
rect 302236 178069 302266 178099
rect 302266 178069 302278 178099
rect 302278 178069 302292 178099
rect 302316 178069 302330 178099
rect 302330 178069 302342 178099
rect 302342 178069 302372 178099
rect 302396 178069 302406 178099
rect 302406 178069 302452 178099
rect 302156 178057 302212 178069
rect 302236 178057 302292 178069
rect 302316 178057 302372 178069
rect 302396 178057 302452 178069
rect 302156 178043 302202 178057
rect 302202 178043 302212 178057
rect 302236 178043 302266 178057
rect 302266 178043 302278 178057
rect 302278 178043 302292 178057
rect 302316 178043 302330 178057
rect 302330 178043 302342 178057
rect 302342 178043 302372 178057
rect 302396 178043 302406 178057
rect 302406 178043 302452 178057
rect 302156 178005 302202 178019
rect 302202 178005 302212 178019
rect 302236 178005 302266 178019
rect 302266 178005 302278 178019
rect 302278 178005 302292 178019
rect 302316 178005 302330 178019
rect 302330 178005 302342 178019
rect 302342 178005 302372 178019
rect 302396 178005 302406 178019
rect 302406 178005 302452 178019
rect 302156 177993 302212 178005
rect 302236 177993 302292 178005
rect 302316 177993 302372 178005
rect 302396 177993 302452 178005
rect 302156 177963 302202 177993
rect 302202 177963 302212 177993
rect 302236 177963 302266 177993
rect 302266 177963 302278 177993
rect 302278 177963 302292 177993
rect 302316 177963 302330 177993
rect 302330 177963 302342 177993
rect 302342 177963 302372 177993
rect 302396 177963 302406 177993
rect 302406 177963 302452 177993
rect 302156 177929 302212 177939
rect 302236 177929 302292 177939
rect 302316 177929 302372 177939
rect 302396 177929 302452 177939
rect 302156 177883 302202 177929
rect 302202 177883 302212 177929
rect 302236 177883 302266 177929
rect 302266 177883 302278 177929
rect 302278 177883 302292 177929
rect 302316 177883 302330 177929
rect 302330 177883 302342 177929
rect 302342 177883 302372 177929
rect 302396 177883 302406 177929
rect 302406 177883 302452 177929
rect 309156 178133 309202 178179
rect 309202 178133 309212 178179
rect 309236 178133 309266 178179
rect 309266 178133 309278 178179
rect 309278 178133 309292 178179
rect 309316 178133 309330 178179
rect 309330 178133 309342 178179
rect 309342 178133 309372 178179
rect 309396 178133 309406 178179
rect 309406 178133 309452 178179
rect 309156 178123 309212 178133
rect 309236 178123 309292 178133
rect 309316 178123 309372 178133
rect 309396 178123 309452 178133
rect 309156 178069 309202 178099
rect 309202 178069 309212 178099
rect 309236 178069 309266 178099
rect 309266 178069 309278 178099
rect 309278 178069 309292 178099
rect 309316 178069 309330 178099
rect 309330 178069 309342 178099
rect 309342 178069 309372 178099
rect 309396 178069 309406 178099
rect 309406 178069 309452 178099
rect 309156 178057 309212 178069
rect 309236 178057 309292 178069
rect 309316 178057 309372 178069
rect 309396 178057 309452 178069
rect 309156 178043 309202 178057
rect 309202 178043 309212 178057
rect 309236 178043 309266 178057
rect 309266 178043 309278 178057
rect 309278 178043 309292 178057
rect 309316 178043 309330 178057
rect 309330 178043 309342 178057
rect 309342 178043 309372 178057
rect 309396 178043 309406 178057
rect 309406 178043 309452 178057
rect 309156 178005 309202 178019
rect 309202 178005 309212 178019
rect 309236 178005 309266 178019
rect 309266 178005 309278 178019
rect 309278 178005 309292 178019
rect 309316 178005 309330 178019
rect 309330 178005 309342 178019
rect 309342 178005 309372 178019
rect 309396 178005 309406 178019
rect 309406 178005 309452 178019
rect 309156 177993 309212 178005
rect 309236 177993 309292 178005
rect 309316 177993 309372 178005
rect 309396 177993 309452 178005
rect 309156 177963 309202 177993
rect 309202 177963 309212 177993
rect 309236 177963 309266 177993
rect 309266 177963 309278 177993
rect 309278 177963 309292 177993
rect 309316 177963 309330 177993
rect 309330 177963 309342 177993
rect 309342 177963 309372 177993
rect 309396 177963 309406 177993
rect 309406 177963 309452 177993
rect 309156 177929 309212 177939
rect 309236 177929 309292 177939
rect 309316 177929 309372 177939
rect 309396 177929 309452 177939
rect 309156 177883 309202 177929
rect 309202 177883 309212 177929
rect 309236 177883 309266 177929
rect 309266 177883 309278 177929
rect 309278 177883 309292 177929
rect 309316 177883 309330 177929
rect 309330 177883 309342 177929
rect 309342 177883 309372 177929
rect 309396 177883 309406 177929
rect 309406 177883 309452 177929
rect 301686 176432 301742 176488
rect 307758 176568 307814 176624
rect 304722 175208 304778 175264
rect 298650 175072 298706 175128
rect 311530 177248 311586 177304
rect 316958 361936 317014 361992
rect 317142 303456 317198 303512
rect 317050 301960 317106 302016
rect 317050 283328 317106 283384
rect 318154 360576 318210 360632
rect 318062 259664 318118 259720
rect 317142 248784 317198 248840
rect 317050 217776 317106 217832
rect 316958 197104 317014 197160
rect 316774 195744 316830 195800
rect 318338 344256 318394 344312
rect 318430 326032 318486 326088
rect 318338 323312 318394 323368
rect 318246 301008 318302 301064
rect 369122 486512 369178 486568
rect 366362 486376 366418 486432
rect 319534 468696 319590 468752
rect 324962 447888 325018 447944
rect 319718 406272 319774 406328
rect 366454 468560 366510 468616
rect 366362 421096 366418 421152
rect 366454 419736 366510 419792
rect 366454 412936 366510 412992
rect 366362 411576 366418 411632
rect 339406 407904 339462 407960
rect 338762 407768 338818 407824
rect 339406 406952 339462 407008
rect 338762 384920 338818 384976
rect 326342 367376 326398 367432
rect 324962 342896 325018 342952
rect 319718 304272 319774 304328
rect 319534 304136 319590 304192
rect 347042 363296 347098 363352
rect 329102 320592 329158 320648
rect 326342 279928 326398 279984
rect 319442 261024 319498 261080
rect 318430 260480 318486 260536
rect 318338 217368 318394 217424
rect 318154 176432 318210 176488
rect 370502 468424 370558 468480
rect 369122 380976 369178 381032
rect 464342 447752 464398 447808
rect 373262 427216 373318 427272
rect 370502 379616 370558 379672
rect 370502 368736 370558 368792
rect 366454 364112 366510 364168
rect 366362 343440 366418 343496
rect 377402 427080 377458 427136
rect 373354 391176 373410 391232
rect 373262 336912 373318 336968
rect 373354 335552 373410 335608
rect 373262 327392 373318 327448
rect 371882 321952 371938 322008
rect 370502 301824 370558 301880
rect 347042 217504 347098 217560
rect 384302 386688 384358 386744
rect 381542 365744 381598 365800
rect 377494 348336 377550 348392
rect 377494 332832 377550 332888
rect 377402 296928 377458 296984
rect 373262 281424 373318 281480
rect 382922 282104 382978 282160
rect 381542 252864 381598 252920
rect 433982 384240 434038 384296
rect 433982 334192 434038 334248
rect 384394 308352 384450 308408
rect 515402 431160 515458 431216
rect 517426 423816 517482 423872
rect 521658 423816 521714 423872
rect 515402 418240 515458 418296
rect 515494 415520 515550 415576
rect 514942 414160 514998 414216
rect 515402 410080 515458 410136
rect 514942 407768 514998 407824
rect 514758 404640 514814 404696
rect 514758 364656 514814 364712
rect 514758 344256 514814 344312
rect 514850 342896 514906 342952
rect 514758 340992 514814 341048
rect 514850 338272 514906 338328
rect 515494 407904 515550 407960
rect 524326 423680 524382 423736
rect 528558 423680 528614 423736
rect 529938 410896 529994 410952
rect 529202 404912 529258 404968
rect 517426 399472 517482 399528
rect 515494 389952 515550 390008
rect 515678 389816 515734 389872
rect 515586 388456 515642 388512
rect 515586 376896 515642 376952
rect 515770 388320 515826 388376
rect 517426 383832 517482 383888
rect 515770 378256 515826 378312
rect 515678 375536 515734 375592
rect 515770 372816 515826 372872
rect 515678 371456 515734 371512
rect 515586 370096 515642 370152
rect 515494 339632 515550 339688
rect 515494 324944 515550 325000
rect 515402 321408 515458 321464
rect 515402 307128 515458 307184
rect 514758 304136 514814 304192
rect 514758 299648 514814 299704
rect 464342 298288 464398 298344
rect 515402 292848 515458 292904
rect 515770 364248 515826 364304
rect 524326 400152 524382 400208
rect 528558 400152 528614 400208
rect 521658 399472 521714 399528
rect 521658 383832 521714 383888
rect 524326 383832 524382 383888
rect 529202 383832 529258 383888
rect 527086 383696 527142 383752
rect 528558 383696 528614 383752
rect 517426 359352 517482 359408
rect 517426 343848 517482 343904
rect 515678 343576 515734 343632
rect 515862 330112 515918 330168
rect 515678 328752 515734 328808
rect 515586 321272 515642 321328
rect 515586 306992 515642 307048
rect 515770 324672 515826 324728
rect 515862 322768 515918 322824
rect 521658 359352 521714 359408
rect 521658 343848 521714 343904
rect 524326 343848 524382 343904
rect 527270 343848 527326 343904
rect 527086 343712 527142 343768
rect 517426 319368 517482 319424
rect 522302 319368 522358 319424
rect 515862 304272 515918 304328
rect 515678 302776 515734 302832
rect 527086 303728 527142 303784
rect 524326 303592 524382 303648
rect 522118 302232 522174 302288
rect 529386 383696 529442 383752
rect 529938 370912 529994 370968
rect 529202 351872 529258 351928
rect 529202 343848 529258 343904
rect 528558 343712 528614 343768
rect 529938 330928 529994 330984
rect 528558 303728 528614 303784
rect 527270 303592 527326 303648
rect 515862 295568 515918 295624
rect 515586 294208 515642 294264
rect 515494 291488 515550 291544
rect 384394 290128 384450 290184
rect 515678 287408 515734 287464
rect 515586 286048 515642 286104
rect 514758 284688 514814 284744
rect 515494 281968 515550 282024
rect 515402 280608 515458 280664
rect 384302 254224 384358 254280
rect 382922 247424 382978 247480
rect 514758 244704 514814 244760
rect 402242 240624 402298 240680
rect 371882 197240 371938 197296
rect 371882 181328 371938 181384
rect 342902 181056 342958 181112
rect 329102 175208 329158 175264
rect 316682 175072 316738 175128
rect 402242 176840 402298 176896
rect 515678 280064 515734 280120
rect 518622 278840 518678 278896
rect 519542 278840 519598 278896
rect 527086 264832 527142 264888
rect 524326 264560 524382 264616
rect 522118 264424 522174 264480
rect 519634 263608 519690 263664
rect 528650 302232 528706 302288
rect 528558 264832 528614 264888
rect 527270 264560 527326 264616
rect 580170 302232 580226 302288
rect 580170 298696 580226 298752
rect 529938 290944 529994 291000
rect 528650 264424 528706 264480
rect 527822 263608 527878 263664
rect 515586 259392 515642 259448
rect 529938 250960 529994 251016
rect 530582 250960 530638 251016
rect 527822 245520 527878 245576
rect 515678 243344 515734 243400
rect 515586 241984 515642 242040
rect 515678 218592 515734 218648
rect 515586 197648 515642 197704
rect 515494 195880 515550 195936
rect 515402 176568 515458 176624
rect 371882 86128 371938 86184
rect 342902 46280 342958 46336
rect 580170 205672 580226 205728
rect 580262 179424 580318 179480
rect 580354 177248 580410 177304
rect 580354 165824 580410 165880
rect 580262 125976 580318 126032
rect 530582 19760 530638 19816
rect 311162 6568 311218 6624
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect 304441 492826 304507 492829
rect 311985 492826 312051 492829
rect 304441 492824 312051 492826
rect 304441 492768 304446 492824
rect 304502 492768 311990 492824
rect 312046 492768 312051 492824
rect 304441 492766 312051 492768
rect 304441 492763 304507 492766
rect 311985 492763 312051 492766
rect 295057 491874 295123 491877
rect 295057 491872 300778 491874
rect 295057 491816 295062 491872
rect 295118 491816 300778 491872
rect 295057 491814 300778 491816
rect 295057 491811 295123 491814
rect 296878 491654 297194 491655
rect 296878 491590 296884 491654
rect 296948 491590 296964 491654
rect 297028 491590 297044 491654
rect 297108 491590 297124 491654
rect 297188 491590 297194 491654
rect 296878 491574 297194 491590
rect 296878 491510 296884 491574
rect 296948 491510 296964 491574
rect 297028 491510 297044 491574
rect 297108 491510 297124 491574
rect 297188 491510 297194 491574
rect 296878 491494 297194 491510
rect 296878 491430 296884 491494
rect 296948 491430 296964 491494
rect 297028 491430 297044 491494
rect 297108 491430 297124 491494
rect 297188 491430 297194 491494
rect 296878 491414 297194 491430
rect 296878 491350 296884 491414
rect 296948 491350 296964 491414
rect 297028 491350 297044 491414
rect 297108 491350 297124 491414
rect 297188 491350 297194 491414
rect 296878 491349 297194 491350
rect 300718 491194 300778 491814
rect 303878 491654 304194 491655
rect 303878 491590 303884 491654
rect 303948 491590 303964 491654
rect 304028 491590 304044 491654
rect 304108 491590 304124 491654
rect 304188 491590 304194 491654
rect 303878 491574 304194 491590
rect 303878 491510 303884 491574
rect 303948 491510 303964 491574
rect 304028 491510 304044 491574
rect 304108 491510 304124 491574
rect 304188 491510 304194 491574
rect 303878 491494 304194 491510
rect 303878 491430 303884 491494
rect 303948 491430 303964 491494
rect 304028 491430 304044 491494
rect 304108 491430 304124 491494
rect 304188 491430 304194 491494
rect 310878 491654 311194 491655
rect 310878 491590 310884 491654
rect 310948 491590 310964 491654
rect 311028 491590 311044 491654
rect 311108 491590 311124 491654
rect 311188 491590 311194 491654
rect 310878 491574 311194 491590
rect 310878 491510 310884 491574
rect 310948 491510 310964 491574
rect 311028 491510 311044 491574
rect 311108 491510 311124 491574
rect 311188 491510 311194 491574
rect 310878 491494 311194 491510
rect 304441 491466 304507 491469
rect 303878 491414 304194 491430
rect 303878 491350 303884 491414
rect 303948 491350 303964 491414
rect 304028 491350 304044 491414
rect 304108 491350 304124 491414
rect 304188 491350 304194 491414
rect 303878 491349 304194 491350
rect 304398 491464 304507 491466
rect 304398 491408 304446 491464
rect 304502 491408 304507 491464
rect 304398 491403 304507 491408
rect 310878 491430 310884 491494
rect 310948 491430 310964 491494
rect 311028 491430 311044 491494
rect 311108 491430 311124 491494
rect 311188 491430 311194 491494
rect 310878 491414 311194 491430
rect 300853 491194 300919 491197
rect 300718 491192 300919 491194
rect 300718 491136 300858 491192
rect 300914 491136 300919 491192
rect 300718 491134 300919 491136
rect 300853 491131 300919 491134
rect 304216 491058 304282 491061
rect 304398 491058 304458 491403
rect 310878 491350 310884 491414
rect 310948 491350 310964 491414
rect 311028 491350 311044 491414
rect 311108 491350 311124 491414
rect 311188 491350 311194 491414
rect 310878 491349 311194 491350
rect 304216 491056 304458 491058
rect 304216 491000 304221 491056
rect 304277 491000 304458 491056
rect 304216 490998 304458 491000
rect 304216 490995 304282 490998
rect 295146 490538 295462 490539
rect 295146 490474 295152 490538
rect 295216 490474 295232 490538
rect 295296 490474 295312 490538
rect 295376 490474 295392 490538
rect 295456 490474 295462 490538
rect 295146 490458 295462 490474
rect 295146 490394 295152 490458
rect 295216 490394 295232 490458
rect 295296 490394 295312 490458
rect 295376 490394 295392 490458
rect 295456 490394 295462 490458
rect 295146 490378 295462 490394
rect 295146 490314 295152 490378
rect 295216 490314 295232 490378
rect 295296 490314 295312 490378
rect 295376 490314 295392 490378
rect 295456 490314 295462 490378
rect 295146 490313 295462 490314
rect 311525 489698 311591 489701
rect 319437 489698 319503 489701
rect 311525 489696 319503 489698
rect 311525 489640 311530 489696
rect 311586 489640 319442 489696
rect 319498 489640 319503 489696
rect 311525 489638 319503 489640
rect 311525 489635 311591 489638
rect 319437 489635 319503 489638
rect 303878 489482 304194 489483
rect 303878 489418 303884 489482
rect 303948 489418 303964 489482
rect 304028 489418 304044 489482
rect 304108 489418 304124 489482
rect 304188 489418 304194 489482
rect 303878 489402 304194 489418
rect 303878 489338 303884 489402
rect 303948 489338 303964 489402
rect 304028 489338 304044 489402
rect 304108 489338 304124 489402
rect 304188 489338 304194 489402
rect 303878 489322 304194 489338
rect 303878 489258 303884 489322
rect 303948 489258 303964 489322
rect 304028 489258 304044 489322
rect 304108 489258 304124 489322
rect 304188 489258 304194 489322
rect 303878 489242 304194 489258
rect 303878 489178 303884 489242
rect 303948 489178 303964 489242
rect 304028 489178 304044 489242
rect 304108 489178 304124 489242
rect 304188 489178 304194 489242
rect 303878 489177 304194 489178
rect 310878 489482 311194 489483
rect 310878 489418 310884 489482
rect 310948 489418 310964 489482
rect 311028 489418 311044 489482
rect 311108 489418 311124 489482
rect 311188 489418 311194 489482
rect 310878 489402 311194 489418
rect 310878 489338 310884 489402
rect 310948 489338 310964 489402
rect 311028 489338 311044 489402
rect 311108 489338 311124 489402
rect 311188 489338 311194 489402
rect 310878 489322 311194 489338
rect 310878 489258 310884 489322
rect 310948 489258 310964 489322
rect 311028 489258 311044 489322
rect 311108 489258 311124 489322
rect 311188 489258 311194 489322
rect 310878 489242 311194 489258
rect 310878 489178 310884 489242
rect 310948 489178 310964 489242
rect 311028 489178 311044 489242
rect 311108 489178 311124 489242
rect 311188 489178 311194 489242
rect 310878 489177 311194 489178
rect -960 488596 480 488836
rect 305085 486706 305151 486709
rect 318333 486706 318399 486709
rect 305085 486704 318399 486706
rect 305085 486648 305090 486704
rect 305146 486648 318338 486704
rect 318394 486648 318399 486704
rect 305085 486646 318399 486648
rect 305085 486643 305151 486646
rect 318333 486643 318399 486646
rect 301773 486570 301839 486573
rect 369117 486570 369183 486573
rect 301773 486568 369183 486570
rect 301773 486512 301778 486568
rect 301834 486512 369122 486568
rect 369178 486512 369183 486568
rect 301773 486510 369183 486512
rect 301773 486507 301839 486510
rect 369117 486507 369183 486510
rect 298737 486434 298803 486437
rect 366357 486434 366423 486437
rect 298737 486432 366423 486434
rect 298737 486376 298742 486432
rect 298798 486376 366362 486432
rect 366418 486376 366423 486432
rect 298737 486374 366423 486376
rect 298737 486371 298803 486374
rect 366357 486371 366423 486374
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 305545 474738 305611 474741
rect 311985 474738 312051 474741
rect 313641 474738 313707 474741
rect 305545 474736 313707 474738
rect 305545 474680 305550 474736
rect 305606 474680 311990 474736
rect 312046 474680 313646 474736
rect 313702 474680 313707 474736
rect 305545 474678 313707 474680
rect 305545 474675 305611 474678
rect 311985 474675 312051 474678
rect 313641 474675 313707 474678
rect 293861 474058 293927 474061
rect 295057 474058 295123 474061
rect 301405 474058 301471 474061
rect 293861 474056 301471 474058
rect 293861 474000 293866 474056
rect 293922 474000 295062 474056
rect 295118 474000 301410 474056
rect 301466 474000 301471 474056
rect 293861 473998 301471 474000
rect 293861 473995 293927 473998
rect 295057 473995 295123 473998
rect 301405 473995 301471 473998
rect 308121 474058 308187 474061
rect 318241 474058 318307 474061
rect 308121 474056 318307 474058
rect 308121 474000 308126 474056
rect 308182 474000 318246 474056
rect 318302 474000 318307 474056
rect 308121 473998 318307 474000
rect 308121 473995 308187 473998
rect 318241 473995 318307 473998
rect 312169 473514 312235 473517
rect 313733 473514 313799 473517
rect 309182 473512 313799 473514
rect 309182 473456 312174 473512
rect 312230 473456 313738 473512
rect 313794 473456 313799 473512
rect 309182 473454 313799 473456
rect 296878 473114 297194 473115
rect 296878 473050 296884 473114
rect 296948 473050 296964 473114
rect 297028 473050 297044 473114
rect 297108 473050 297124 473114
rect 297188 473050 297194 473114
rect 296878 473034 297194 473050
rect 296878 472970 296884 473034
rect 296948 472970 296964 473034
rect 297028 472970 297044 473034
rect 297108 472970 297124 473034
rect 297188 472970 297194 473034
rect 303878 473114 304194 473115
rect 303878 473050 303884 473114
rect 303948 473050 303964 473114
rect 304028 473050 304044 473114
rect 304108 473050 304124 473114
rect 304188 473050 304194 473114
rect 303878 473034 304194 473050
rect 296878 472954 297194 472970
rect 296878 472890 296884 472954
rect 296948 472890 296964 472954
rect 297028 472890 297044 472954
rect 297108 472890 297124 472954
rect 297188 472890 297194 472954
rect 301405 472970 301471 472973
rect 303878 472970 303884 473034
rect 303948 472970 303964 473034
rect 304028 472970 304044 473034
rect 304108 472970 304124 473034
rect 304188 472970 304194 473034
rect 305545 472970 305611 472973
rect 301405 472968 301514 472970
rect 301405 472912 301410 472968
rect 301466 472912 301514 472968
rect 301405 472907 301514 472912
rect 296878 472874 297194 472890
rect 296878 472810 296884 472874
rect 296948 472810 296964 472874
rect 297028 472810 297044 472874
rect 297108 472810 297124 472874
rect 297188 472810 297194 472874
rect 296878 472809 297194 472810
rect 301454 472698 301514 472907
rect 303878 472954 304194 472970
rect 303878 472890 303884 472954
rect 303948 472890 303964 472954
rect 304028 472890 304044 472954
rect 304108 472890 304124 472954
rect 304188 472890 304194 472954
rect 303878 472874 304194 472890
rect 303878 472810 303884 472874
rect 303948 472810 303964 472874
rect 304028 472810 304044 472874
rect 304108 472810 304124 472874
rect 304188 472810 304194 472874
rect 303878 472809 304194 472810
rect 305502 472968 305611 472970
rect 305502 472912 305550 472968
rect 305606 472912 305611 472968
rect 305502 472907 305611 472912
rect 301589 472698 301655 472701
rect 301454 472696 301655 472698
rect 301454 472640 301594 472696
rect 301650 472640 301655 472696
rect 301454 472638 301655 472640
rect 301589 472635 301655 472638
rect 305502 472565 305562 472907
rect 309182 472701 309242 473454
rect 312169 473451 312235 473454
rect 313733 473451 313799 473454
rect 310513 473378 310579 473381
rect 313825 473378 313891 473381
rect 310513 473376 313891 473378
rect 310513 473320 310518 473376
rect 310574 473320 313830 473376
rect 313886 473320 313891 473376
rect 310513 473318 313891 473320
rect 310513 473315 310579 473318
rect 310878 473114 311194 473115
rect 310878 473050 310884 473114
rect 310948 473050 310964 473114
rect 311028 473050 311044 473114
rect 311108 473050 311124 473114
rect 311188 473050 311194 473114
rect 310878 473034 311194 473050
rect 310878 472970 310884 473034
rect 310948 472970 310964 473034
rect 311028 472970 311044 473034
rect 311108 472970 311124 473034
rect 311188 472970 311194 473034
rect 310878 472954 311194 472970
rect 310878 472890 310884 472954
rect 310948 472890 310964 472954
rect 311028 472890 311044 472954
rect 311108 472890 311124 472954
rect 311188 472890 311194 472954
rect 310878 472874 311194 472890
rect 310878 472810 310884 472874
rect 310948 472810 310964 472874
rect 311028 472810 311044 472874
rect 311108 472810 311124 472874
rect 311188 472810 311194 472874
rect 310878 472809 311194 472810
rect 309133 472696 309242 472701
rect 309133 472640 309138 472696
rect 309194 472640 309242 472696
rect 309133 472638 309242 472640
rect 312310 472701 312370 473318
rect 313825 473315 313891 473318
rect 312310 472696 312419 472701
rect 312310 472640 312358 472696
rect 312414 472640 312419 472696
rect 312310 472638 312419 472640
rect 309133 472635 309199 472638
rect 312353 472635 312419 472638
rect 305502 472560 305569 472565
rect 305502 472504 305508 472560
rect 305564 472504 305569 472560
rect 305502 472502 305569 472504
rect 305503 472499 305569 472502
rect 302146 472013 302462 472014
rect 302146 471949 302152 472013
rect 302216 471949 302232 472013
rect 302296 471949 302312 472013
rect 302376 471949 302392 472013
rect 302456 471949 302462 472013
rect 302146 471933 302462 471949
rect 302146 471869 302152 471933
rect 302216 471869 302232 471933
rect 302296 471869 302312 471933
rect 302376 471869 302392 471933
rect 302456 471869 302462 471933
rect 302146 471853 302462 471869
rect 302146 471789 302152 471853
rect 302216 471789 302232 471853
rect 302296 471789 302312 471853
rect 302376 471789 302392 471853
rect 302456 471789 302462 471853
rect 302146 471773 302462 471789
rect 302146 471709 302152 471773
rect 302216 471709 302232 471773
rect 302296 471709 302312 471773
rect 302376 471709 302392 471773
rect 302456 471709 302462 471773
rect 302146 471708 302462 471709
rect 309146 472013 309462 472014
rect 309146 471949 309152 472013
rect 309216 471949 309232 472013
rect 309296 471949 309312 472013
rect 309376 471949 309392 472013
rect 309456 471949 309462 472013
rect 309146 471933 309462 471949
rect 309146 471869 309152 471933
rect 309216 471869 309232 471933
rect 309296 471869 309312 471933
rect 309376 471869 309392 471933
rect 309456 471869 309462 471933
rect 309146 471853 309462 471869
rect 309146 471789 309152 471853
rect 309216 471789 309232 471853
rect 309296 471789 309312 471853
rect 309376 471789 309392 471853
rect 309456 471789 309462 471853
rect 309146 471773 309462 471789
rect 309146 471709 309152 471773
rect 309216 471709 309232 471773
rect 309296 471709 309312 471773
rect 309376 471709 309392 471773
rect 309456 471709 309462 471773
rect 309146 471708 309462 471709
rect 583520 471324 584960 471564
rect 313641 471066 313707 471069
rect 318057 471066 318123 471069
rect 313641 471064 318123 471066
rect 313641 471008 313646 471064
rect 313702 471008 318062 471064
rect 318118 471008 318123 471064
rect 313641 471006 318123 471008
rect 313641 471003 313707 471006
rect 318057 471003 318123 471006
rect 310053 470658 310119 470661
rect 309948 470656 310119 470658
rect 309948 470600 310058 470656
rect 310114 470600 310119 470656
rect 309948 470598 310119 470600
rect 310053 470595 310119 470598
rect 310053 468754 310119 468757
rect 319529 468754 319595 468757
rect 310053 468752 319595 468754
rect 310053 468696 310058 468752
rect 310114 468696 319534 468752
rect 319590 468696 319595 468752
rect 310053 468694 319595 468696
rect 310053 468691 310119 468694
rect 319529 468691 319595 468694
rect 299289 468618 299355 468621
rect 366449 468618 366515 468621
rect 299289 468616 366515 468618
rect 299289 468560 299294 468616
rect 299350 468560 366454 468616
rect 366510 468560 366515 468616
rect 299289 468558 366515 468560
rect 299289 468555 299355 468558
rect 366449 468555 366515 468558
rect 302877 468482 302943 468485
rect 370497 468482 370563 468485
rect 302877 468480 370563 468482
rect 302877 468424 302882 468480
rect 302938 468424 370502 468480
rect 370558 468424 370563 468480
rect 302877 468422 370563 468424
rect 302877 468419 302943 468422
rect 370497 468419 370563 468422
rect 306465 467938 306531 467941
rect 313917 467938 313983 467941
rect 306465 467936 313983 467938
rect 306465 467880 306470 467936
rect 306526 467880 313922 467936
rect 313978 467880 313983 467936
rect 306465 467878 313983 467880
rect 306465 467875 306531 467878
rect 313917 467875 313983 467878
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect 312997 455426 313063 455429
rect 313825 455426 313891 455429
rect 312997 455424 313891 455426
rect 312997 455368 313002 455424
rect 313058 455368 313830 455424
rect 313886 455368 313891 455424
rect 312997 455366 313891 455368
rect 312997 455363 313063 455366
rect 313825 455363 313891 455366
rect 312537 453930 312603 453933
rect 313733 453930 313799 453933
rect 312537 453928 313799 453930
rect 312537 453872 312542 453928
rect 312598 453872 313738 453928
rect 313794 453872 313799 453928
rect 312537 453870 313799 453872
rect 312537 453867 312603 453870
rect 313733 453867 313799 453870
rect 308305 452706 308371 452709
rect 312537 452706 312603 452709
rect 308305 452704 312603 452706
rect 308305 452648 308310 452704
rect 308366 452648 312542 452704
rect 312598 452648 312603 452704
rect 308305 452646 312603 452648
rect 308305 452643 308371 452646
rect 312537 452643 312603 452646
rect 296878 452058 297194 452059
rect 296878 451994 296884 452058
rect 296948 451994 296964 452058
rect 297028 451994 297044 452058
rect 297108 451994 297124 452058
rect 297188 451994 297194 452058
rect 296878 451978 297194 451994
rect 296878 451914 296884 451978
rect 296948 451914 296964 451978
rect 297028 451914 297044 451978
rect 297108 451914 297124 451978
rect 297188 451914 297194 451978
rect 296878 451898 297194 451914
rect 296878 451834 296884 451898
rect 296948 451834 296964 451898
rect 297028 451834 297044 451898
rect 297108 451834 297124 451898
rect 297188 451834 297194 451898
rect 296878 451818 297194 451834
rect 296878 451754 296884 451818
rect 296948 451754 296964 451818
rect 297028 451754 297044 451818
rect 297108 451754 297124 451818
rect 297188 451754 297194 451818
rect 296878 451738 297194 451754
rect 296878 451674 296884 451738
rect 296948 451674 296964 451738
rect 297028 451674 297044 451738
rect 297108 451674 297124 451738
rect 297188 451674 297194 451738
rect 296878 451658 297194 451674
rect 296878 451594 296884 451658
rect 296948 451594 296964 451658
rect 297028 451594 297044 451658
rect 297108 451594 297124 451658
rect 297188 451594 297194 451658
rect 296878 451578 297194 451594
rect 296878 451514 296884 451578
rect 296948 451514 296964 451578
rect 297028 451514 297044 451578
rect 297108 451514 297124 451578
rect 297188 451514 297194 451578
rect 296878 451498 297194 451514
rect 296878 451434 296884 451498
rect 296948 451434 296964 451498
rect 297028 451434 297044 451498
rect 297108 451434 297124 451498
rect 297188 451434 297194 451498
rect 296878 451418 297194 451434
rect 296878 451354 296884 451418
rect 296948 451354 296964 451418
rect 297028 451354 297044 451418
rect 297108 451354 297124 451418
rect 297188 451354 297194 451418
rect 296878 451338 297194 451354
rect 296878 451274 296884 451338
rect 296948 451274 296964 451338
rect 297028 451274 297044 451338
rect 297108 451274 297124 451338
rect 297188 451274 297194 451338
rect 296878 451273 297194 451274
rect 303878 452058 304194 452059
rect 303878 451994 303884 452058
rect 303948 451994 303964 452058
rect 304028 451994 304044 452058
rect 304108 451994 304124 452058
rect 304188 451994 304194 452058
rect 303878 451978 304194 451994
rect 303878 451914 303884 451978
rect 303948 451914 303964 451978
rect 304028 451914 304044 451978
rect 304108 451914 304124 451978
rect 304188 451914 304194 451978
rect 303878 451898 304194 451914
rect 303878 451834 303884 451898
rect 303948 451834 303964 451898
rect 304028 451834 304044 451898
rect 304108 451834 304124 451898
rect 304188 451834 304194 451898
rect 303878 451818 304194 451834
rect 303878 451754 303884 451818
rect 303948 451754 303964 451818
rect 304028 451754 304044 451818
rect 304108 451754 304124 451818
rect 304188 451754 304194 451818
rect 310909 452058 311065 452059
rect 310909 451994 310915 452058
rect 310979 451994 310995 452058
rect 311059 451994 311065 452058
rect 310909 451978 311065 451994
rect 310909 451914 310915 451978
rect 310979 451914 310995 451978
rect 311059 451914 311065 451978
rect 310909 451898 311065 451914
rect 310909 451834 310915 451898
rect 310979 451834 310995 451898
rect 311059 451834 311065 451898
rect 310909 451818 311065 451834
rect 303878 451738 304194 451754
rect 303878 451674 303884 451738
rect 303948 451674 303964 451738
rect 304028 451674 304044 451738
rect 304108 451674 304124 451738
rect 304188 451674 304194 451738
rect 308305 451752 308371 451757
rect 308305 451696 308310 451752
rect 308366 451696 308371 451752
rect 308305 451691 308371 451696
rect 310909 451754 310915 451818
rect 310979 451754 310995 451818
rect 311059 451754 311065 451818
rect 310909 451738 311065 451754
rect 303878 451658 304194 451674
rect 303878 451594 303884 451658
rect 303948 451594 303964 451658
rect 304028 451594 304044 451658
rect 304108 451594 304124 451658
rect 304188 451594 304194 451658
rect 303878 451578 304194 451594
rect 303878 451514 303884 451578
rect 303948 451514 303964 451578
rect 304028 451514 304044 451578
rect 304108 451514 304124 451578
rect 304188 451514 304194 451578
rect 303878 451498 304194 451514
rect 303878 451434 303884 451498
rect 303948 451434 303964 451498
rect 304028 451434 304044 451498
rect 304108 451434 304124 451498
rect 304188 451434 304194 451498
rect 303878 451418 304194 451434
rect 308019 451482 308085 451485
rect 308308 451482 308368 451691
rect 308019 451480 308368 451482
rect 308019 451424 308024 451480
rect 308080 451424 308368 451480
rect 308019 451422 308368 451424
rect 310909 451674 310915 451738
rect 310979 451674 310995 451738
rect 311059 451674 311065 451738
rect 310909 451658 311065 451674
rect 310909 451594 310915 451658
rect 310979 451594 310995 451658
rect 311059 451594 311065 451658
rect 310909 451578 311065 451594
rect 310909 451514 310915 451578
rect 310979 451514 310995 451578
rect 311059 451514 311065 451578
rect 310909 451498 311065 451514
rect 310909 451434 310915 451498
rect 310979 451434 310995 451498
rect 311059 451434 311065 451498
rect 308019 451419 308085 451422
rect 303878 451354 303884 451418
rect 303948 451354 303964 451418
rect 304028 451354 304044 451418
rect 304108 451354 304124 451418
rect 304188 451354 304194 451418
rect 303878 451338 304194 451354
rect 303878 451274 303884 451338
rect 303948 451274 303964 451338
rect 304028 451274 304044 451338
rect 304108 451274 304124 451338
rect 304188 451274 304194 451338
rect 303878 451273 304194 451274
rect 310909 451418 311065 451434
rect 310909 451354 310915 451418
rect 310979 451354 310995 451418
rect 311059 451354 311065 451418
rect 310909 451338 311065 451354
rect 310909 451274 310915 451338
rect 310979 451274 310995 451338
rect 311059 451274 311065 451338
rect 310909 451273 311065 451274
rect 312169 450666 312235 450669
rect 315297 450666 315363 450669
rect 312169 450664 315363 450666
rect 312169 450608 312174 450664
rect 312230 450608 315302 450664
rect 315358 450608 315363 450664
rect 312169 450606 315363 450608
rect 312169 450603 312235 450606
rect 315297 450603 315363 450606
rect 310888 450181 311124 450182
rect 310888 450117 310894 450181
rect 310958 450117 310974 450181
rect 311038 450117 311054 450181
rect 311118 450117 311124 450181
rect 310888 450101 311124 450117
rect 310888 450037 310894 450101
rect 310958 450037 310974 450101
rect 311038 450037 311054 450101
rect 311118 450037 311124 450101
rect 310888 450021 311124 450037
rect 310888 449957 310894 450021
rect 310958 449957 310974 450021
rect 311038 449957 311054 450021
rect 311118 449957 311124 450021
rect 310888 449941 311124 449957
rect 310888 449877 310894 449941
rect 310958 449877 310974 449941
rect 311038 449877 311054 449941
rect 311118 449877 311124 449941
rect 310888 449861 311124 449877
rect 310888 449797 310894 449861
rect 310958 449797 310974 449861
rect 311038 449797 311054 449861
rect 311118 449797 311124 449861
rect 310888 449781 311124 449797
rect 310888 449717 310894 449781
rect 310958 449717 310974 449781
rect 311038 449717 311054 449781
rect 311118 449717 311124 449781
rect 310888 449701 311124 449717
rect -960 449428 480 449668
rect 310888 449637 310894 449701
rect 310958 449637 310974 449701
rect 311038 449637 311054 449701
rect 311118 449637 311124 449701
rect 310888 449636 311124 449637
rect 293861 449170 293927 449173
rect 300853 449170 300919 449173
rect 293861 449168 300919 449170
rect 293861 449112 293866 449168
rect 293922 449112 300858 449168
rect 300914 449112 300919 449168
rect 293861 449110 300919 449112
rect 293861 449107 293927 449110
rect 300853 449107 300919 449110
rect 306189 449170 306255 449173
rect 313457 449170 313523 449173
rect 306189 449168 313523 449170
rect 306189 449112 306194 449168
rect 306250 449112 313462 449168
rect 313518 449112 313523 449168
rect 306189 449110 313523 449112
rect 306189 449107 306255 449110
rect 313457 449107 313523 449110
rect 302233 448218 302299 448221
rect 314285 448218 314351 448221
rect 302233 448216 314351 448218
rect 302233 448160 302238 448216
rect 302294 448160 314290 448216
rect 314346 448160 314351 448216
rect 302233 448158 314351 448160
rect 302233 448155 302299 448158
rect 314285 448155 314351 448158
rect 298921 448082 298987 448085
rect 312629 448082 312695 448085
rect 298921 448080 312695 448082
rect 298921 448024 298926 448080
rect 298982 448024 312634 448080
rect 312690 448024 312695 448080
rect 298921 448022 312695 448024
rect 298921 448019 298987 448022
rect 312629 448019 312695 448022
rect 305545 447946 305611 447949
rect 324957 447946 325023 447949
rect 305545 447944 325023 447946
rect 305545 447888 305550 447944
rect 305606 447888 324962 447944
rect 325018 447888 325023 447944
rect 305545 447886 325023 447888
rect 305545 447883 305611 447886
rect 324957 447883 325023 447886
rect 308857 447810 308923 447813
rect 464337 447810 464403 447813
rect 308857 447808 464403 447810
rect 308857 447752 308862 447808
rect 308918 447752 464342 447808
rect 464398 447752 464403 447808
rect 308857 447750 464403 447752
rect 308857 447747 308923 447750
rect 464337 447747 464403 447750
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 308489 433258 308555 433261
rect 312537 433258 312603 433261
rect 313365 433258 313431 433261
rect 308489 433256 313431 433258
rect 308489 433200 308494 433256
rect 308550 433200 312542 433256
rect 312598 433200 313370 433256
rect 313426 433200 313431 433256
rect 308489 433198 313431 433200
rect 308489 433195 308555 433198
rect 312537 433195 312603 433198
rect 313365 433195 313431 433198
rect 305177 432170 305243 432173
rect 306281 432170 306347 432173
rect 313273 432170 313339 432173
rect 305177 432168 313339 432170
rect 305177 432112 305182 432168
rect 305238 432112 306286 432168
rect 306342 432112 313278 432168
rect 313334 432112 313339 432168
rect 305177 432110 313339 432112
rect 305177 432107 305243 432110
rect 306281 432107 306347 432110
rect 313273 432107 313339 432110
rect 583520 431476 584960 431716
rect 312629 431218 312695 431221
rect 515397 431218 515463 431221
rect 312629 431216 515463 431218
rect 312629 431160 312634 431216
rect 312690 431160 515402 431216
rect 515458 431160 515463 431216
rect 312629 431158 515463 431160
rect 312629 431155 312695 431158
rect 515397 431155 515463 431158
rect 300853 430810 300919 430813
rect 305177 430810 305243 430813
rect 308489 430810 308555 430813
rect 300853 430808 301514 430810
rect 300853 430752 300858 430808
rect 300914 430752 301514 430808
rect 300853 430750 301514 430752
rect 300853 430747 300919 430750
rect 301454 430405 301514 430750
rect 305134 430808 305243 430810
rect 305134 430752 305182 430808
rect 305238 430752 305243 430808
rect 305134 430747 305243 430752
rect 308446 430808 308555 430810
rect 308446 430752 308494 430808
rect 308550 430752 308555 430808
rect 308446 430747 308555 430752
rect 305134 430405 305194 430747
rect 308446 430405 308506 430747
rect 301454 430400 301563 430405
rect 301454 430344 301502 430400
rect 301558 430344 301563 430400
rect 301454 430342 301563 430344
rect 301497 430339 301563 430342
rect 305086 430400 305194 430405
rect 305086 430344 305091 430400
rect 305147 430344 305194 430400
rect 305086 430342 305194 430344
rect 308397 430400 308506 430405
rect 308397 430344 308402 430400
rect 308458 430344 308506 430400
rect 308397 430342 308506 430344
rect 305086 430339 305152 430342
rect 308397 430339 308463 430342
rect 309146 429998 309452 429999
rect 309146 429994 309187 429998
rect 309251 429994 309267 429998
rect 309331 429994 309347 429998
rect 309411 429994 309452 429998
rect 309146 429938 309151 429994
rect 309447 429938 309452 429994
rect 309146 429934 309187 429938
rect 309251 429934 309267 429938
rect 309331 429934 309347 429938
rect 309411 429934 309452 429938
rect 309146 429918 309452 429934
rect 309146 429914 309187 429918
rect 309251 429914 309267 429918
rect 309331 429914 309347 429918
rect 309411 429914 309452 429918
rect 309146 429858 309151 429914
rect 309447 429858 309452 429914
rect 309146 429854 309187 429858
rect 309251 429854 309267 429858
rect 309331 429854 309347 429858
rect 309411 429854 309452 429858
rect 309146 429838 309452 429854
rect 309146 429834 309187 429838
rect 309251 429834 309267 429838
rect 309331 429834 309347 429838
rect 309411 429834 309452 429838
rect 309146 429778 309151 429834
rect 309447 429778 309452 429834
rect 309146 429774 309187 429778
rect 309251 429774 309267 429778
rect 309331 429774 309347 429778
rect 309411 429774 309452 429778
rect 309146 429758 309452 429774
rect 309146 429754 309187 429758
rect 309251 429754 309267 429758
rect 309331 429754 309347 429758
rect 309411 429754 309452 429758
rect 309146 429698 309151 429754
rect 309447 429698 309452 429754
rect 309146 429694 309187 429698
rect 309251 429694 309267 429698
rect 309331 429694 309347 429698
rect 309411 429694 309452 429698
rect 309146 429693 309452 429694
rect 312997 429042 313063 429045
rect 315481 429042 315547 429045
rect 312997 429040 315547 429042
rect 312997 428984 313002 429040
rect 313058 428984 315486 429040
rect 315542 428984 315547 429040
rect 312997 428982 315547 428984
rect 312997 428979 313063 428982
rect 315481 428979 315547 428982
rect 309366 428501 309426 428604
rect 309366 428496 309475 428501
rect 309366 428440 309414 428496
rect 309470 428440 309475 428496
rect 309366 428438 309475 428440
rect 309409 428435 309475 428438
rect 300853 427954 300919 427957
rect 301681 427954 301747 427957
rect 300853 427952 301747 427954
rect 300853 427896 300858 427952
rect 300914 427896 301686 427952
rect 301742 427896 301747 427952
rect 300853 427894 301747 427896
rect 300853 427891 300919 427894
rect 301681 427891 301747 427894
rect 302509 427410 302575 427413
rect 314469 427410 314535 427413
rect 302509 427408 314535 427410
rect 302509 427352 302514 427408
rect 302570 427352 314474 427408
rect 314530 427352 314535 427408
rect 302509 427350 314535 427352
rect 302509 427347 302575 427350
rect 314469 427347 314535 427350
rect 305913 427274 305979 427277
rect 373257 427274 373323 427277
rect 305913 427272 373323 427274
rect 305913 427216 305918 427272
rect 305974 427216 373262 427272
rect 373318 427216 373323 427272
rect 305913 427214 373323 427216
rect 305913 427211 305979 427214
rect 373257 427211 373323 427214
rect 309409 427138 309475 427141
rect 377397 427138 377463 427141
rect 309409 427136 377463 427138
rect 309409 427080 309414 427136
rect 309470 427080 377402 427136
rect 377458 427080 377463 427136
rect 309409 427078 377463 427080
rect 309409 427075 309475 427078
rect 377397 427075 377463 427078
rect 517421 423874 517487 423877
rect 521653 423874 521719 423877
rect 517421 423872 521719 423874
rect 517421 423816 517426 423872
rect 517482 423816 521658 423872
rect 521714 423816 521719 423872
rect 517421 423814 521719 423816
rect 517421 423811 517487 423814
rect 521653 423811 521719 423814
rect 524321 423738 524387 423741
rect 528553 423738 528619 423741
rect 524321 423736 528619 423738
rect -960 423452 480 423692
rect 524321 423680 524326 423736
rect 524382 423680 528558 423736
rect 528614 423680 528619 423736
rect 524321 423678 528619 423680
rect 524321 423675 524387 423678
rect 528553 423675 528619 423678
rect 309041 423602 309107 423605
rect 313365 423602 313431 423605
rect 309041 423600 313431 423602
rect 309041 423544 309046 423600
rect 309102 423544 313370 423600
rect 313426 423544 313431 423600
rect 309041 423542 313431 423544
rect 309041 423539 309107 423542
rect 313365 423539 313431 423542
rect 366357 421154 366423 421157
rect 366357 421152 509250 421154
rect 366357 421096 366362 421152
rect 366418 421096 509250 421152
rect 366357 421094 509250 421096
rect 366357 421091 366423 421094
rect 509190 421018 509250 421094
rect 509190 420958 518052 421018
rect 366449 419794 366515 419797
rect 366449 419792 509250 419794
rect 366449 419736 366454 419792
rect 366510 419736 509250 419792
rect 366449 419734 509250 419736
rect 366449 419731 366515 419734
rect 509190 419658 509250 419734
rect 509190 419598 518052 419658
rect 515397 418298 515463 418301
rect 515397 418296 518052 418298
rect 515397 418240 515402 418296
rect 515458 418240 518052 418296
rect 515397 418238 518052 418240
rect 515397 418235 515463 418238
rect 583520 418148 584960 418388
rect 299013 417074 299079 417077
rect 299013 417072 509250 417074
rect 299013 417016 299018 417072
rect 299074 417016 509250 417072
rect 299013 417014 509250 417016
rect 299013 417011 299079 417014
rect 509190 416938 509250 417014
rect 509190 416878 518052 416938
rect 515489 415578 515555 415581
rect 515489 415576 518052 415578
rect 515489 415520 515494 415576
rect 515550 415520 518052 415576
rect 515489 415518 518052 415520
rect 515489 415515 515555 415518
rect 514937 414218 515003 414221
rect 514937 414216 518052 414218
rect 514937 414160 514942 414216
rect 514998 414160 518052 414216
rect 514937 414158 518052 414160
rect 514937 414155 515003 414158
rect 366449 412994 366515 412997
rect 366449 412992 509250 412994
rect 366449 412936 366454 412992
rect 366510 412936 509250 412992
rect 366449 412934 509250 412936
rect 366449 412931 366515 412934
rect 509190 412858 509250 412934
rect 509190 412798 518052 412858
rect 366357 411634 366423 411637
rect 366357 411632 509250 411634
rect 366357 411576 366362 411632
rect 366418 411576 509250 411632
rect 366357 411574 509250 411576
rect 366357 411571 366423 411574
rect 312445 411498 312511 411501
rect 313273 411498 313339 411501
rect 312445 411496 313339 411498
rect 312445 411440 312450 411496
rect 312506 411440 313278 411496
rect 313334 411440 313339 411496
rect 312445 411438 313339 411440
rect 509190 411498 509250 411574
rect 509190 411438 518052 411498
rect 312445 411435 312511 411438
rect 313273 411435 313339 411438
rect 305177 411362 305243 411365
rect 312261 411362 312327 411365
rect 313181 411362 313247 411365
rect 305177 411360 313247 411362
rect 305177 411304 305182 411360
rect 305238 411304 312266 411360
rect 312322 411304 313186 411360
rect 313242 411304 313247 411360
rect 305177 411302 313247 411304
rect 305177 411299 305243 411302
rect 312261 411299 312327 411302
rect 313181 411299 313247 411302
rect 529933 410954 529999 410957
rect 527804 410952 529999 410954
rect 527804 410896 529938 410952
rect 529994 410896 529999 410952
rect 527804 410894 529999 410896
rect 529933 410891 529999 410894
rect -960 410396 480 410636
rect 295149 410274 295215 410277
rect 301037 410274 301103 410277
rect 309041 410274 309107 410277
rect 312077 410274 312143 410277
rect 295149 410272 301103 410274
rect 295149 410216 295154 410272
rect 295210 410216 301042 410272
rect 301098 410216 301103 410272
rect 295149 410214 301103 410216
rect 295149 410211 295215 410214
rect 301037 410211 301103 410214
rect 308446 410272 312143 410274
rect 308446 410216 309046 410272
rect 309102 410216 312082 410272
rect 312138 410216 312143 410272
rect 308446 410214 312143 410216
rect 296878 410084 297194 410085
rect 296878 410020 296884 410084
rect 296948 410020 296964 410084
rect 297028 410020 297044 410084
rect 297108 410020 297124 410084
rect 297188 410020 297194 410084
rect 296878 410004 297194 410020
rect 296878 409940 296884 410004
rect 296948 409940 296964 410004
rect 297028 409940 297044 410004
rect 297108 409940 297124 410004
rect 297188 409940 297194 410004
rect 296878 409924 297194 409940
rect 296878 409860 296884 409924
rect 296948 409860 296964 409924
rect 297028 409860 297044 409924
rect 297108 409860 297124 409924
rect 297188 409860 297194 409924
rect 303878 410084 304194 410085
rect 303878 410020 303884 410084
rect 303948 410020 303964 410084
rect 304028 410020 304044 410084
rect 304108 410020 304124 410084
rect 304188 410020 304194 410084
rect 303878 410004 304194 410020
rect 303878 409940 303884 410004
rect 303948 409940 303964 410004
rect 304028 409940 304044 410004
rect 304108 409940 304124 410004
rect 304188 409940 304194 410004
rect 303878 409924 304194 409940
rect 296878 409844 297194 409860
rect 296878 409780 296884 409844
rect 296948 409780 296964 409844
rect 297028 409780 297044 409844
rect 297108 409780 297124 409844
rect 297188 409780 297194 409844
rect 301037 409864 301103 409869
rect 301037 409808 301042 409864
rect 301098 409808 301103 409864
rect 301037 409803 301103 409808
rect 303878 409860 303884 409924
rect 303948 409860 303964 409924
rect 304028 409860 304044 409924
rect 304108 409860 304124 409924
rect 304188 409860 304194 409924
rect 305177 409866 305243 409869
rect 303878 409844 304194 409860
rect 296878 409779 297194 409780
rect 301040 409594 301100 409803
rect 303878 409780 303884 409844
rect 303948 409780 303964 409844
rect 304028 409780 304044 409844
rect 304108 409780 304124 409844
rect 304188 409780 304194 409844
rect 303878 409779 304194 409780
rect 305134 409864 305243 409866
rect 305134 409808 305182 409864
rect 305238 409808 305243 409864
rect 305134 409803 305243 409808
rect 301221 409594 301287 409597
rect 301040 409592 301287 409594
rect 301040 409536 301226 409592
rect 301282 409536 301287 409592
rect 301040 409534 301287 409536
rect 301221 409531 301287 409534
rect 304544 409594 304610 409597
rect 305134 409594 305194 409803
rect 304544 409592 305194 409594
rect 304544 409536 304549 409592
rect 304605 409536 305194 409592
rect 304544 409534 305194 409536
rect 307809 409594 307875 409597
rect 308446 409594 308506 410214
rect 309041 410211 309107 410214
rect 312077 410211 312143 410214
rect 515397 410138 515463 410141
rect 515397 410136 518052 410138
rect 310878 410084 311194 410085
rect 310878 410020 310884 410084
rect 310948 410020 310964 410084
rect 311028 410020 311044 410084
rect 311108 410020 311124 410084
rect 311188 410020 311194 410084
rect 515397 410080 515402 410136
rect 515458 410080 518052 410136
rect 515397 410078 518052 410080
rect 515397 410075 515463 410078
rect 310878 410004 311194 410020
rect 310878 409940 310884 410004
rect 310948 409940 310964 410004
rect 311028 409940 311044 410004
rect 311108 409940 311124 410004
rect 311188 409940 311194 410004
rect 310878 409924 311194 409940
rect 310878 409860 310884 409924
rect 310948 409860 310964 409924
rect 311028 409860 311044 409924
rect 311108 409860 311124 409924
rect 311188 409860 311194 409924
rect 310878 409844 311194 409860
rect 310878 409780 310884 409844
rect 310948 409780 310964 409844
rect 311028 409780 311044 409844
rect 311108 409780 311124 409844
rect 311188 409780 311194 409844
rect 310878 409779 311194 409780
rect 307809 409592 308506 409594
rect 307809 409536 307814 409592
rect 307870 409536 308506 409592
rect 307809 409534 308506 409536
rect 304544 409531 304610 409534
rect 307809 409531 307875 409534
rect 302146 408998 302462 408999
rect 302146 408934 302152 408998
rect 302216 408934 302232 408998
rect 302296 408934 302312 408998
rect 302376 408934 302392 408998
rect 302456 408934 302462 408998
rect 302146 408918 302462 408934
rect 302146 408854 302152 408918
rect 302216 408854 302232 408918
rect 302296 408854 302312 408918
rect 302376 408854 302392 408918
rect 302456 408854 302462 408918
rect 302146 408838 302462 408854
rect 317045 408914 317111 408917
rect 317045 408912 509250 408914
rect 317045 408856 317050 408912
rect 317106 408856 509250 408912
rect 317045 408854 509250 408856
rect 317045 408851 317111 408854
rect 302146 408774 302152 408838
rect 302216 408774 302232 408838
rect 302296 408774 302312 408838
rect 302376 408774 302392 408838
rect 302456 408774 302462 408838
rect 302146 408758 302462 408774
rect 302146 408694 302152 408758
rect 302216 408694 302232 408758
rect 302296 408694 302312 408758
rect 302376 408694 302392 408758
rect 302456 408694 302462 408758
rect 509190 408778 509250 408854
rect 509190 408718 518052 408778
rect 302146 408693 302462 408694
rect 312169 407962 312235 407965
rect 315573 407962 315639 407965
rect 312169 407960 315639 407962
rect 310878 407912 311194 407913
rect 310878 407848 310884 407912
rect 310948 407848 310964 407912
rect 311028 407848 311044 407912
rect 311108 407848 311124 407912
rect 311188 407848 311194 407912
rect 312169 407904 312174 407960
rect 312230 407904 315578 407960
rect 315634 407904 315639 407960
rect 312169 407902 315639 407904
rect 312169 407899 312235 407902
rect 315573 407899 315639 407902
rect 339401 407962 339467 407965
rect 515489 407962 515555 407965
rect 339401 407960 515555 407962
rect 339401 407904 339406 407960
rect 339462 407904 515494 407960
rect 515550 407904 515555 407960
rect 339401 407902 515555 407904
rect 339401 407899 339467 407902
rect 515489 407899 515555 407902
rect 310878 407832 311194 407848
rect 310878 407768 310884 407832
rect 310948 407768 310964 407832
rect 311028 407768 311044 407832
rect 311108 407768 311124 407832
rect 311188 407768 311194 407832
rect 310878 407752 311194 407768
rect 338757 407826 338823 407829
rect 514937 407826 515003 407829
rect 338757 407824 515003 407826
rect 338757 407768 338762 407824
rect 338818 407768 514942 407824
rect 514998 407768 515003 407824
rect 338757 407766 515003 407768
rect 338757 407763 338823 407766
rect 514937 407763 515003 407766
rect 310878 407688 310884 407752
rect 310948 407688 310964 407752
rect 311028 407688 311044 407752
rect 311108 407688 311124 407752
rect 311188 407688 311194 407752
rect 310878 407672 311194 407688
rect 310878 407608 310884 407672
rect 310948 407608 310964 407672
rect 311028 407608 311044 407672
rect 311108 407608 311124 407672
rect 311188 407608 311194 407672
rect 310878 407607 311194 407608
rect 315757 407554 315823 407557
rect 315757 407552 509250 407554
rect 315757 407496 315762 407552
rect 315818 407496 509250 407552
rect 315757 407494 509250 407496
rect 315757 407491 315823 407494
rect 509190 407418 509250 407494
rect 509190 407358 518052 407418
rect 298829 407010 298895 407013
rect 339401 407010 339467 407013
rect 298829 407008 339467 407010
rect 298829 406952 298834 407008
rect 298890 406952 339406 407008
rect 339462 406952 339467 407008
rect 298829 406950 339467 406952
rect 298829 406947 298895 406950
rect 339401 406947 339467 406950
rect 308673 406330 308739 406333
rect 319713 406330 319779 406333
rect 308673 406328 319779 406330
rect 308673 406272 308678 406328
rect 308734 406272 319718 406328
rect 319774 406272 319779 406328
rect 308673 406270 319779 406272
rect 308673 406267 308739 406270
rect 319713 406267 319779 406270
rect 315665 406194 315731 406197
rect 315665 406192 509250 406194
rect 315665 406136 315670 406192
rect 315726 406136 509250 406192
rect 315665 406134 509250 406136
rect 315665 406131 315731 406134
rect 509190 406058 509250 406134
rect 509190 405998 518052 406058
rect 529197 404970 529263 404973
rect 583520 404970 584960 405060
rect 529197 404968 584960 404970
rect 529197 404912 529202 404968
rect 529258 404912 584960 404968
rect 529197 404910 584960 404912
rect 529197 404907 529263 404910
rect 583520 404820 584960 404910
rect 514753 404698 514819 404701
rect 514753 404696 518052 404698
rect 514753 404640 514758 404696
rect 514814 404640 518052 404696
rect 514753 404638 518052 404640
rect 514753 404635 514819 404638
rect 315389 403474 315455 403477
rect 315389 403472 509250 403474
rect 315389 403416 315394 403472
rect 315450 403416 509250 403472
rect 315389 403414 509250 403416
rect 315389 403411 315455 403414
rect 509190 403338 509250 403414
rect 509190 403278 518052 403338
rect 316769 402114 316835 402117
rect 316769 402112 509250 402114
rect 316769 402056 316774 402112
rect 316830 402056 509250 402112
rect 316769 402054 509250 402056
rect 316769 402051 316835 402054
rect 509190 401978 509250 402054
rect 509190 401918 518052 401978
rect 316677 400754 316743 400757
rect 316677 400752 509250 400754
rect 316677 400696 316682 400752
rect 316738 400696 509250 400752
rect 316677 400694 509250 400696
rect 316677 400691 316743 400694
rect 509190 400618 509250 400694
rect 509190 400558 518052 400618
rect 524321 400210 524387 400213
rect 528553 400210 528619 400213
rect 524321 400208 528619 400210
rect 524321 400152 524326 400208
rect 524382 400152 528558 400208
rect 528614 400152 528619 400208
rect 524321 400150 528619 400152
rect 524321 400147 524387 400150
rect 528553 400147 528619 400150
rect 517421 399530 517487 399533
rect 521653 399530 521719 399533
rect 517421 399528 521719 399530
rect 517421 399472 517426 399528
rect 517482 399472 521658 399528
rect 521714 399472 521719 399528
rect 517421 399470 521719 399472
rect 517421 399467 517487 399470
rect 521653 399467 521719 399470
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect 305913 391506 305979 391509
rect 312261 391506 312327 391509
rect 305913 391504 312327 391506
rect 305913 391448 305918 391504
rect 305974 391448 312266 391504
rect 312322 391448 312327 391504
rect 305913 391446 312327 391448
rect 305913 391443 305979 391446
rect 312261 391443 312327 391446
rect 305545 391234 305611 391237
rect 373349 391234 373415 391237
rect 305545 391232 373415 391234
rect 305545 391176 305550 391232
rect 305606 391176 373354 391232
rect 373410 391176 373415 391232
rect 305545 391174 373415 391176
rect 305545 391171 305611 391174
rect 373349 391171 373415 391174
rect 294965 390690 295031 390693
rect 301589 390690 301655 390693
rect 294965 390688 301655 390690
rect 294965 390632 294970 390688
rect 295026 390632 301594 390688
rect 301650 390632 301655 390688
rect 294965 390630 301655 390632
rect 294965 390627 295031 390630
rect 301589 390627 301655 390630
rect 309501 390690 309567 390693
rect 312077 390690 312143 390693
rect 309501 390688 312143 390690
rect 309501 390632 309506 390688
rect 309562 390632 312082 390688
rect 312138 390632 312143 390688
rect 309501 390630 312143 390632
rect 309501 390627 309567 390630
rect 312077 390627 312143 390630
rect 312261 390690 312327 390693
rect 314377 390690 314443 390693
rect 312261 390688 314443 390690
rect 312261 390632 312266 390688
rect 312322 390632 314382 390688
rect 314438 390632 314443 390688
rect 312261 390630 314443 390632
rect 312261 390627 312327 390630
rect 314377 390627 314443 390630
rect 313917 390010 313983 390013
rect 515489 390010 515555 390013
rect 313917 390008 515555 390010
rect 313917 389952 313922 390008
rect 313978 389952 515494 390008
rect 515550 389952 515555 390008
rect 313917 389950 515555 389952
rect 313917 389947 313983 389950
rect 515489 389947 515555 389950
rect 301957 389874 302023 389877
rect 515673 389874 515739 389877
rect 301957 389872 515739 389874
rect 301957 389816 301962 389872
rect 302018 389816 515678 389872
rect 515734 389816 515739 389872
rect 301957 389814 515739 389816
rect 301957 389811 302023 389814
rect 515673 389811 515739 389814
rect 296878 389085 297194 389086
rect 296878 389021 296884 389085
rect 296948 389021 296964 389085
rect 297028 389021 297044 389085
rect 297108 389021 297124 389085
rect 297188 389021 297194 389085
rect 296878 389005 297194 389021
rect 296878 388941 296884 389005
rect 296948 388941 296964 389005
rect 297028 388941 297044 389005
rect 297108 388941 297124 389005
rect 297188 388941 297194 389005
rect 296878 388925 297194 388941
rect 303878 389085 304194 389086
rect 303878 389021 303884 389085
rect 303948 389021 303964 389085
rect 304028 389021 304044 389085
rect 304108 389021 304124 389085
rect 304188 389021 304194 389085
rect 303878 389005 304194 389021
rect 303878 388941 303884 389005
rect 303948 388941 303964 389005
rect 304028 388941 304044 389005
rect 304108 388941 304124 389005
rect 304188 388941 304194 389005
rect 303878 388925 304194 388941
rect 310878 389085 311194 389086
rect 310878 389021 310884 389085
rect 310948 389021 310964 389085
rect 311028 389021 311044 389085
rect 311108 389021 311124 389085
rect 311188 389021 311194 389085
rect 310878 389005 311194 389021
rect 310878 388941 310884 389005
rect 310948 388941 310964 389005
rect 311028 388941 311044 389005
rect 311108 388941 311124 389005
rect 311188 388941 311194 389005
rect 310878 388925 311194 388941
rect 296878 388861 296884 388925
rect 296948 388861 296964 388925
rect 297028 388861 297044 388925
rect 297108 388861 297124 388925
rect 297188 388861 297194 388925
rect 296878 388845 297194 388861
rect 301589 388922 301655 388925
rect 301589 388920 301698 388922
rect 301589 388864 301594 388920
rect 301650 388864 301698 388920
rect 301589 388859 301698 388864
rect 296878 388781 296884 388845
rect 296948 388781 296964 388845
rect 297028 388781 297044 388845
rect 297108 388781 297124 388845
rect 297188 388781 297194 388845
rect 296878 388780 297194 388781
rect 301638 388653 301698 388859
rect 303878 388861 303884 388925
rect 303948 388861 303964 388925
rect 304028 388861 304044 388925
rect 304108 388861 304124 388925
rect 304188 388861 304194 388925
rect 305913 388922 305979 388925
rect 303878 388845 304194 388861
rect 303878 388781 303884 388845
rect 303948 388781 303964 388845
rect 304028 388781 304044 388845
rect 304108 388781 304124 388845
rect 304188 388781 304194 388845
rect 303878 388780 304194 388781
rect 305870 388920 305979 388922
rect 305870 388864 305918 388920
rect 305974 388864 305979 388920
rect 305870 388859 305979 388864
rect 309501 388922 309567 388925
rect 309501 388920 309610 388922
rect 309501 388864 309506 388920
rect 309562 388864 309610 388920
rect 309501 388859 309610 388864
rect 301589 388648 301698 388653
rect 301589 388592 301594 388648
rect 301650 388592 301698 388648
rect 301589 388590 301698 388592
rect 301589 388587 301655 388590
rect 305870 388517 305930 388859
rect 309550 388653 309610 388859
rect 310878 388861 310884 388925
rect 310948 388861 310964 388925
rect 311028 388861 311044 388925
rect 311108 388861 311124 388925
rect 311188 388861 311194 388925
rect 310878 388845 311194 388861
rect 310878 388781 310884 388845
rect 310948 388781 310964 388845
rect 311028 388781 311044 388845
rect 311108 388781 311124 388845
rect 311188 388781 311194 388845
rect 310878 388780 311194 388781
rect 309501 388648 309610 388653
rect 309501 388592 309506 388648
rect 309562 388592 309610 388648
rect 309501 388590 309610 388592
rect 309501 388587 309567 388590
rect 305870 388512 305951 388517
rect 305870 388456 305890 388512
rect 305946 388456 305951 388512
rect 305870 388454 305951 388456
rect 305885 388451 305951 388454
rect 314469 388514 314535 388517
rect 515581 388514 515647 388517
rect 314469 388512 515647 388514
rect 314469 388456 314474 388512
rect 314530 388456 515586 388512
rect 515642 388456 515647 388512
rect 314469 388454 515647 388456
rect 314469 388451 314535 388454
rect 515581 388451 515647 388454
rect 314285 388378 314351 388381
rect 515765 388378 515831 388381
rect 314285 388376 515831 388378
rect 314285 388320 314290 388376
rect 314346 388320 515770 388376
rect 515826 388320 515831 388376
rect 314285 388318 515831 388320
rect 314285 388315 314351 388318
rect 515765 388315 515831 388318
rect 295146 388002 295462 388003
rect 295146 387938 295152 388002
rect 295216 387938 295232 388002
rect 295296 387938 295312 388002
rect 295376 387938 295392 388002
rect 295456 387938 295462 388002
rect 295146 387922 295462 387938
rect 295146 387858 295152 387922
rect 295216 387858 295232 387922
rect 295296 387858 295312 387922
rect 295376 387858 295392 387922
rect 295456 387858 295462 387922
rect 295146 387842 295462 387858
rect 295146 387778 295152 387842
rect 295216 387778 295232 387842
rect 295296 387778 295312 387842
rect 295376 387778 295392 387842
rect 295456 387778 295462 387842
rect 295146 387762 295462 387778
rect 295146 387698 295152 387762
rect 295216 387698 295232 387762
rect 295296 387698 295312 387762
rect 295376 387698 295392 387762
rect 295456 387698 295462 387762
rect 295146 387697 295462 387698
rect 302146 387997 302462 387998
rect 302146 387933 302152 387997
rect 302216 387933 302232 387997
rect 302296 387933 302312 387997
rect 302376 387933 302392 387997
rect 302456 387933 302462 387997
rect 302146 387917 302462 387933
rect 302146 387853 302152 387917
rect 302216 387853 302232 387917
rect 302296 387853 302312 387917
rect 302376 387853 302392 387917
rect 302456 387853 302462 387917
rect 302146 387837 302462 387853
rect 302146 387773 302152 387837
rect 302216 387773 302232 387837
rect 302296 387773 302312 387837
rect 302376 387773 302392 387837
rect 302456 387773 302462 387837
rect 302146 387757 302462 387773
rect 302146 387693 302152 387757
rect 302216 387693 302232 387757
rect 302296 387693 302312 387757
rect 302376 387693 302392 387757
rect 302456 387693 302462 387757
rect 302146 387692 302462 387693
rect 309146 387997 309462 387998
rect 309146 387933 309152 387997
rect 309216 387933 309232 387997
rect 309296 387933 309312 387997
rect 309376 387933 309392 387997
rect 309456 387933 309462 387997
rect 309146 387917 309462 387933
rect 309146 387853 309152 387917
rect 309216 387853 309232 387917
rect 309296 387853 309312 387917
rect 309376 387853 309392 387917
rect 309456 387853 309462 387917
rect 309146 387837 309462 387853
rect 309146 387773 309152 387837
rect 309216 387773 309232 387837
rect 309296 387773 309312 387837
rect 309376 387773 309392 387837
rect 309456 387773 309462 387837
rect 309146 387757 309462 387773
rect 309146 387693 309152 387757
rect 309216 387693 309232 387757
rect 309296 387693 309312 387757
rect 309376 387693 309392 387757
rect 309456 387693 309462 387757
rect 309146 387692 309462 387693
rect 310999 387519 311145 387520
rect 310999 387455 311040 387519
rect 311104 387455 311145 387519
rect 310999 387454 311145 387455
rect 303919 387402 304065 387403
rect 303919 387338 303960 387402
rect 304024 387338 304065 387402
rect 303919 387337 304065 387338
rect 384297 386746 384363 386749
rect 314180 386744 384363 386746
rect 314180 386688 384302 386744
rect 384358 386688 384363 386744
rect 314180 386686 384363 386688
rect 384297 386683 384363 386686
rect 310053 386474 310119 386477
rect 313273 386474 313339 386477
rect 314561 386474 314627 386477
rect 310053 386472 314627 386474
rect 310053 386416 310058 386472
rect 310114 386416 313278 386472
rect 313334 386416 314566 386472
rect 314622 386416 314627 386472
rect 310053 386414 314627 386416
rect 310053 386411 310119 386414
rect 313273 386411 313339 386414
rect 314561 386411 314627 386414
rect 307661 386338 307727 386341
rect 309593 386338 309659 386341
rect 307661 386336 309659 386338
rect 307661 386280 307666 386336
rect 307722 386280 309598 386336
rect 309654 386280 309659 386336
rect 307661 386278 309659 386280
rect 307661 386275 307727 386278
rect 309593 386275 309659 386278
rect 299289 384978 299355 384981
rect 338757 384978 338823 384981
rect 299289 384976 338823 384978
rect 299289 384920 299294 384976
rect 299350 384920 338762 384976
rect 338818 384920 338823 384976
rect 299289 384918 338823 384920
rect 299289 384915 299355 384918
rect 338757 384915 338823 384918
rect 310421 384842 310487 384845
rect 312537 384842 312603 384845
rect 310421 384840 312603 384842
rect 310421 384784 310426 384840
rect 310482 384784 312542 384840
rect 312598 384784 312603 384840
rect 310421 384782 312603 384784
rect 310421 384779 310487 384782
rect 312537 384779 312603 384782
rect -960 384284 480 384524
rect 306741 384298 306807 384301
rect 433977 384298 434043 384301
rect 306741 384296 434043 384298
rect 306741 384240 306746 384296
rect 306802 384240 433982 384296
rect 434038 384240 434043 384296
rect 306741 384238 434043 384240
rect 306741 384235 306807 384238
rect 433977 384235 434043 384238
rect 517421 383890 517487 383893
rect 521653 383890 521719 383893
rect 517421 383888 521719 383890
rect 517421 383832 517426 383888
rect 517482 383832 521658 383888
rect 521714 383832 521719 383888
rect 517421 383830 521719 383832
rect 517421 383827 517487 383830
rect 521653 383827 521719 383830
rect 524321 383890 524387 383893
rect 529197 383890 529263 383893
rect 524321 383888 529263 383890
rect 524321 383832 524326 383888
rect 524382 383832 529202 383888
rect 529258 383832 529263 383888
rect 524321 383830 529263 383832
rect 524321 383827 524387 383830
rect 529197 383827 529263 383830
rect 527081 383754 527147 383757
rect 528553 383754 528619 383757
rect 529381 383754 529447 383757
rect 527081 383752 529447 383754
rect 527081 383696 527086 383752
rect 527142 383696 528558 383752
rect 528614 383696 529386 383752
rect 529442 383696 529447 383752
rect 527081 383694 529447 383696
rect 527081 383691 527147 383694
rect 528553 383691 528619 383694
rect 529381 383691 529447 383694
rect 369117 381034 369183 381037
rect 369117 381032 518052 381034
rect 369117 380976 369122 381032
rect 369178 380976 518052 381032
rect 369117 380974 518052 380976
rect 369117 380971 369183 380974
rect 370497 379674 370563 379677
rect 370497 379672 518052 379674
rect 370497 379616 370502 379672
rect 370558 379616 518052 379672
rect 370497 379614 518052 379616
rect 370497 379611 370563 379614
rect 515765 378314 515831 378317
rect 515765 378312 518052 378314
rect 515765 378256 515770 378312
rect 515826 378256 518052 378312
rect 583520 378300 584960 378540
rect 515765 378254 518052 378256
rect 515765 378251 515831 378254
rect 515581 376954 515647 376957
rect 515581 376952 518052 376954
rect 515581 376896 515586 376952
rect 515642 376896 518052 376952
rect 515581 376894 518052 376896
rect 515581 376891 515647 376894
rect 515673 375594 515739 375597
rect 515673 375592 518052 375594
rect 515673 375536 515678 375592
rect 515734 375536 518052 375592
rect 515673 375534 518052 375536
rect 515673 375531 515739 375534
rect 303153 374234 303219 374237
rect 303153 374232 518052 374234
rect 303153 374176 303158 374232
rect 303214 374176 518052 374232
rect 303153 374174 518052 374176
rect 303153 374171 303219 374174
rect 515765 372874 515831 372877
rect 515765 372872 518052 372874
rect 515765 372816 515770 372872
rect 515826 372816 518052 372872
rect 515765 372814 518052 372816
rect 515765 372811 515831 372814
rect 515673 371514 515739 371517
rect 515673 371512 518052 371514
rect -960 371228 480 371468
rect 515673 371456 515678 371512
rect 515734 371456 518052 371512
rect 515673 371454 518052 371456
rect 515673 371451 515739 371454
rect 529933 370970 529999 370973
rect 527804 370968 529999 370970
rect 527804 370912 529938 370968
rect 529994 370912 529999 370968
rect 527804 370910 529999 370912
rect 529933 370907 529999 370910
rect 515581 370154 515647 370157
rect 515581 370152 518052 370154
rect 515581 370096 515586 370152
rect 515642 370096 518052 370152
rect 515581 370094 518052 370096
rect 515581 370091 515647 370094
rect 304533 368930 304599 368933
rect 310973 368930 311039 368933
rect 314377 368930 314443 368933
rect 304533 368928 314443 368930
rect 304533 368872 304538 368928
rect 304594 368872 310978 368928
rect 311034 368872 314382 368928
rect 314438 368872 314443 368928
rect 304533 368870 314443 368872
rect 304533 368867 304599 368870
rect 310973 368867 311039 368870
rect 314377 368867 314443 368870
rect 370497 368794 370563 368797
rect 370497 368792 518052 368794
rect 370497 368736 370502 368792
rect 370558 368736 518052 368792
rect 370497 368734 518052 368736
rect 370497 368731 370563 368734
rect 295241 368522 295307 368525
rect 295241 368520 299490 368522
rect 295241 368464 295246 368520
rect 295302 368464 299490 368520
rect 295241 368462 299490 368464
rect 295241 368459 295307 368462
rect 299430 367298 299490 368462
rect 304533 367978 304599 367981
rect 307569 367978 307635 367981
rect 304398 367976 304599 367978
rect 304398 367920 304538 367976
rect 304594 367920 304599 367976
rect 304398 367918 304599 367920
rect 303904 367570 303970 367573
rect 304398 367570 304458 367918
rect 304533 367915 304599 367918
rect 307526 367976 307635 367978
rect 307526 367920 307574 367976
rect 307630 367920 307635 367976
rect 307526 367915 307635 367920
rect 310053 367978 310119 367981
rect 310053 367976 310162 367978
rect 310053 367920 310058 367976
rect 310114 367920 310162 367976
rect 310053 367915 310162 367920
rect 303904 367568 304458 367570
rect 303904 367512 303909 367568
rect 303965 367512 304458 367568
rect 303904 367510 304458 367512
rect 307526 367573 307586 367915
rect 310102 367573 310162 367915
rect 307526 367568 307635 367573
rect 307526 367512 307574 367568
rect 307630 367512 307635 367568
rect 307526 367510 307635 367512
rect 303904 367507 303970 367510
rect 307569 367507 307635 367510
rect 310053 367568 310162 367573
rect 310053 367512 310058 367568
rect 310114 367512 310162 367568
rect 310053 367510 310162 367512
rect 310053 367507 310119 367510
rect 326337 367434 326403 367437
rect 326337 367432 518052 367434
rect 326337 367376 326342 367432
rect 326398 367376 518052 367432
rect 326337 367374 518052 367376
rect 326337 367371 326403 367374
rect 299749 367298 299815 367301
rect 299430 367296 299815 367298
rect 299430 367240 299754 367296
rect 299810 367240 299815 367296
rect 299430 367238 299815 367240
rect 299749 367235 299815 367238
rect 314009 366074 314075 366077
rect 314009 366072 518052 366074
rect 314009 366016 314014 366072
rect 314070 366016 518052 366072
rect 314009 366014 518052 366016
rect 314009 366011 314075 366014
rect 381537 365802 381603 365805
rect 310868 365800 381603 365802
rect 310868 365744 381542 365800
rect 381598 365744 381603 365800
rect 310868 365742 381603 365744
rect 381537 365739 381603 365742
rect 583520 364972 584960 365212
rect 514753 364714 514819 364717
rect 514753 364712 518052 364714
rect 514753 364656 514758 364712
rect 514814 364656 518052 364712
rect 514753 364654 518052 364656
rect 514753 364651 514819 364654
rect 301681 364306 301747 364309
rect 515765 364306 515831 364309
rect 301681 364304 515831 364306
rect 301681 364248 301686 364304
rect 301742 364248 515770 364304
rect 515826 364248 515831 364304
rect 301681 364246 515831 364248
rect 301681 364243 301747 364246
rect 515765 364243 515831 364246
rect 298645 364170 298711 364173
rect 366449 364170 366515 364173
rect 298645 364168 366515 364170
rect 298645 364112 298650 364168
rect 298706 364112 366454 364168
rect 366510 364112 366515 364168
rect 298645 364110 366515 364112
rect 298645 364107 298711 364110
rect 366449 364107 366515 364110
rect 347037 363354 347103 363357
rect 347037 363352 518052 363354
rect 347037 363296 347042 363352
rect 347098 363296 518052 363352
rect 347037 363294 518052 363296
rect 347037 363291 347103 363294
rect 307937 363082 308003 363085
rect 312905 363082 312971 363085
rect 307937 363080 312971 363082
rect 307937 363024 307942 363080
rect 307998 363024 312910 363080
rect 312966 363024 312971 363080
rect 307937 363022 312971 363024
rect 307937 363019 308003 363022
rect 312905 363019 312971 363022
rect 316953 361994 317019 361997
rect 316953 361992 518052 361994
rect 316953 361936 316958 361992
rect 317014 361936 518052 361992
rect 316953 361934 518052 361936
rect 316953 361931 317019 361934
rect 318149 360634 318215 360637
rect 318149 360632 518052 360634
rect 318149 360576 318154 360632
rect 318210 360576 518052 360632
rect 318149 360574 518052 360576
rect 318149 360571 318215 360574
rect 517421 359410 517487 359413
rect 521653 359410 521719 359413
rect 517421 359408 521719 359410
rect 517421 359352 517426 359408
rect 517482 359352 521658 359408
rect 521714 359352 521719 359408
rect 517421 359350 521719 359352
rect 517421 359347 517487 359350
rect 521653 359347 521719 359350
rect -960 358308 480 358548
rect 529197 351930 529263 351933
rect 583520 351930 584960 352020
rect 529197 351928 584960 351930
rect 529197 351872 529202 351928
rect 529258 351872 584960 351928
rect 529197 351870 584960 351872
rect 529197 351867 529263 351870
rect 583520 351780 584960 351870
rect 304717 348394 304783 348397
rect 377489 348394 377555 348397
rect 304717 348392 377555 348394
rect 304717 348336 304722 348392
rect 304778 348336 377494 348392
rect 377550 348336 377555 348392
rect 304717 348334 377555 348336
rect 304717 348331 304783 348334
rect 377489 348331 377555 348334
rect 295241 347850 295307 347853
rect 300853 347850 300919 347853
rect 295241 347848 300919 347850
rect 295241 347792 295246 347848
rect 295302 347792 300858 347848
rect 300914 347792 300919 347848
rect 295241 347790 300919 347792
rect 295241 347787 295307 347790
rect 300853 347787 300919 347790
rect 304441 347850 304507 347853
rect 310973 347850 311039 347853
rect 304441 347848 311039 347850
rect 304441 347792 304446 347848
rect 304502 347792 310978 347848
rect 311034 347792 311039 347848
rect 304441 347790 311039 347792
rect 304441 347787 304507 347790
rect 310973 347787 311039 347790
rect 307661 347306 307727 347309
rect 307661 347304 311082 347306
rect 307661 347248 307666 347304
rect 307722 347248 311082 347304
rect 307661 347246 311082 347248
rect 307661 347243 307727 347246
rect 296878 347085 297194 347086
rect 296878 347021 296884 347085
rect 296948 347021 296964 347085
rect 297028 347021 297044 347085
rect 297108 347021 297124 347085
rect 297188 347021 297194 347085
rect 296878 347005 297194 347021
rect 296878 346941 296884 347005
rect 296948 346941 296964 347005
rect 297028 346941 297044 347005
rect 297108 346941 297124 347005
rect 297188 346941 297194 347005
rect 296878 346925 297194 346941
rect 296878 346861 296884 346925
rect 296948 346861 296964 346925
rect 297028 346861 297044 346925
rect 297108 346861 297124 346925
rect 297188 346861 297194 346925
rect 303878 347085 304194 347086
rect 303878 347021 303884 347085
rect 303948 347021 303964 347085
rect 304028 347021 304044 347085
rect 304108 347021 304124 347085
rect 304188 347021 304194 347085
rect 303878 347005 304194 347021
rect 303878 346941 303884 347005
rect 303948 346941 303964 347005
rect 304028 346941 304044 347005
rect 304108 346941 304124 347005
rect 304188 346941 304194 347005
rect 303878 346925 304194 346941
rect 296878 346845 297194 346861
rect 296878 346781 296884 346845
rect 296948 346781 296964 346845
rect 297028 346781 297044 346845
rect 297108 346781 297124 346845
rect 297188 346781 297194 346845
rect 300853 346898 300919 346901
rect 300853 346896 300962 346898
rect 300853 346840 300858 346896
rect 300914 346840 300962 346896
rect 300853 346835 300962 346840
rect 296878 346780 297194 346781
rect 300902 346629 300962 346835
rect 303878 346861 303884 346925
rect 303948 346861 303964 346925
rect 304028 346861 304044 346925
rect 304108 346861 304124 346925
rect 304188 346861 304194 346925
rect 304441 346898 304507 346901
rect 307661 346898 307727 346901
rect 310513 346898 310579 346901
rect 303878 346845 304194 346861
rect 303878 346781 303884 346845
rect 303948 346781 303964 346845
rect 304028 346781 304044 346845
rect 304108 346781 304124 346845
rect 304188 346781 304194 346845
rect 303878 346780 304194 346781
rect 304398 346896 304507 346898
rect 304398 346840 304446 346896
rect 304502 346840 304507 346896
rect 304398 346835 304507 346840
rect 306790 346896 307727 346898
rect 306790 346840 307666 346896
rect 307722 346840 307727 346896
rect 306790 346838 307727 346840
rect 300853 346624 300962 346629
rect 300853 346568 300858 346624
rect 300914 346568 300962 346624
rect 300853 346566 300962 346568
rect 303889 346626 303955 346629
rect 304398 346626 304458 346835
rect 306790 346629 306850 346838
rect 307661 346835 307727 346838
rect 310470 346896 310579 346898
rect 310470 346840 310518 346896
rect 310574 346840 310579 346896
rect 310470 346835 310579 346840
rect 303889 346624 304458 346626
rect 303889 346568 303894 346624
rect 303950 346568 304458 346624
rect 303889 346566 304458 346568
rect 306741 346624 306850 346629
rect 306741 346568 306746 346624
rect 306802 346568 306850 346624
rect 306741 346566 306850 346568
rect 309869 346626 309935 346629
rect 310470 346626 310530 346835
rect 311022 346765 311082 347246
rect 311022 346760 311131 346765
rect 311022 346704 311070 346760
rect 311126 346704 311131 346760
rect 311022 346702 311131 346704
rect 311065 346699 311131 346702
rect 309869 346624 310530 346626
rect 309869 346568 309874 346624
rect 309930 346568 310530 346624
rect 309869 346566 310530 346568
rect 300853 346563 300919 346566
rect 303889 346563 303955 346566
rect 306741 346563 306807 346566
rect 309869 346563 309935 346566
rect 302146 345983 302462 345984
rect 302146 345919 302152 345983
rect 302216 345919 302232 345983
rect 302296 345919 302312 345983
rect 302376 345919 302392 345983
rect 302456 345919 302462 345983
rect 302146 345903 302462 345919
rect 302146 345839 302152 345903
rect 302216 345839 302232 345903
rect 302296 345839 302312 345903
rect 302376 345839 302392 345903
rect 302456 345839 302462 345903
rect 302146 345823 302462 345839
rect 302146 345759 302152 345823
rect 302216 345759 302232 345823
rect 302296 345759 302312 345823
rect 302376 345759 302392 345823
rect 302456 345759 302462 345823
rect 302146 345743 302462 345759
rect 302146 345679 302152 345743
rect 302216 345679 302232 345743
rect 302296 345679 302312 345743
rect 302376 345679 302392 345743
rect 302456 345679 302462 345743
rect 302146 345678 302462 345679
rect 309146 345983 309462 345984
rect 309146 345919 309152 345983
rect 309216 345919 309232 345983
rect 309296 345919 309312 345983
rect 309376 345919 309392 345983
rect 309456 345919 309462 345983
rect 309146 345903 309462 345919
rect 309146 345839 309152 345903
rect 309216 345839 309232 345903
rect 309296 345839 309312 345903
rect 309376 345839 309392 345903
rect 309456 345839 309462 345903
rect 309146 345823 309462 345839
rect 309146 345759 309152 345823
rect 309216 345759 309232 345823
rect 309296 345759 309312 345823
rect 309376 345759 309392 345823
rect 309456 345759 309462 345823
rect 309146 345743 309462 345759
rect 309146 345679 309152 345743
rect 309216 345679 309232 345743
rect 309296 345679 309312 345743
rect 309376 345679 309392 345743
rect 309456 345679 309462 345743
rect 309146 345678 309462 345679
rect -960 345252 480 345492
rect 314101 345130 314167 345133
rect 310868 345128 314167 345130
rect 310868 345072 314106 345128
rect 314162 345072 314167 345128
rect 310868 345070 314167 345072
rect 314101 345067 314167 345070
rect 318333 344314 318399 344317
rect 514753 344314 514819 344317
rect 318333 344312 514819 344314
rect 318333 344256 318338 344312
rect 318394 344256 514758 344312
rect 514814 344256 514819 344312
rect 318333 344254 514819 344256
rect 318333 344251 318399 344254
rect 514753 344251 514819 344254
rect 517421 343906 517487 343909
rect 521653 343906 521719 343909
rect 517421 343904 521719 343906
rect 517421 343848 517426 343904
rect 517482 343848 521658 343904
rect 521714 343848 521719 343904
rect 517421 343846 521719 343848
rect 517421 343843 517487 343846
rect 521653 343843 521719 343846
rect 524321 343906 524387 343909
rect 527265 343906 527331 343909
rect 529197 343906 529263 343909
rect 524321 343904 529263 343906
rect 524321 343848 524326 343904
rect 524382 343848 527270 343904
rect 527326 343848 529202 343904
rect 529258 343848 529263 343904
rect 524321 343846 529263 343848
rect 524321 343843 524387 343846
rect 527265 343843 527331 343846
rect 529197 343843 529263 343846
rect 527081 343770 527147 343773
rect 528553 343770 528619 343773
rect 527081 343768 528619 343770
rect 527081 343712 527086 343768
rect 527142 343712 528558 343768
rect 528614 343712 528619 343768
rect 527081 343710 528619 343712
rect 527081 343707 527147 343710
rect 528553 343707 528619 343710
rect 301681 343634 301747 343637
rect 515673 343634 515739 343637
rect 301681 343632 515739 343634
rect 301681 343576 301686 343632
rect 301742 343576 515678 343632
rect 515734 343576 515739 343632
rect 301681 343574 515739 343576
rect 301681 343571 301747 343574
rect 515673 343571 515739 343574
rect 298645 343498 298711 343501
rect 366357 343498 366423 343501
rect 298645 343496 366423 343498
rect 298645 343440 298650 343496
rect 298706 343440 366362 343496
rect 366418 343440 366423 343496
rect 298645 343438 366423 343440
rect 298645 343435 298711 343438
rect 366357 343435 366423 343438
rect 324957 342954 325023 342957
rect 514845 342954 514911 342957
rect 324957 342952 514911 342954
rect 324957 342896 324962 342952
rect 325018 342896 514850 342952
rect 514906 342896 514911 342952
rect 324957 342894 514911 342896
rect 324957 342891 325023 342894
rect 514845 342891 514911 342894
rect 307937 342274 308003 342277
rect 312629 342274 312695 342277
rect 307937 342272 312695 342274
rect 307937 342216 307942 342272
rect 307998 342216 312634 342272
rect 312690 342216 312695 342272
rect 307937 342214 312695 342216
rect 307937 342211 308003 342214
rect 312629 342211 312695 342214
rect 514753 341050 514819 341053
rect 514753 341048 518052 341050
rect 514753 340992 514758 341048
rect 514814 340992 518052 341048
rect 514753 340990 518052 340992
rect 514753 340987 514819 340990
rect 307661 340234 307727 340237
rect 311065 340234 311131 340237
rect 307661 340232 311131 340234
rect 307661 340176 307666 340232
rect 307722 340176 311070 340232
rect 311126 340176 311131 340232
rect 307661 340174 311131 340176
rect 307661 340171 307727 340174
rect 311065 340171 311131 340174
rect 515489 339690 515555 339693
rect 515489 339688 518052 339690
rect 515489 339632 515494 339688
rect 515550 339632 518052 339688
rect 515489 339630 518052 339632
rect 515489 339627 515555 339630
rect 583520 338452 584960 338692
rect 514845 338330 514911 338333
rect 514845 338328 518052 338330
rect 514845 338272 514850 338328
rect 514906 338272 518052 338328
rect 514845 338270 518052 338272
rect 514845 338267 514911 338270
rect 373257 336970 373323 336973
rect 373257 336968 518052 336970
rect 373257 336912 373262 336968
rect 373318 336912 518052 336968
rect 373257 336910 518052 336912
rect 373257 336907 373323 336910
rect 373349 335610 373415 335613
rect 373349 335608 518052 335610
rect 373349 335552 373354 335608
rect 373410 335552 518052 335608
rect 373349 335550 518052 335552
rect 373349 335547 373415 335550
rect 433977 334250 434043 334253
rect 433977 334248 518052 334250
rect 433977 334192 433982 334248
rect 434038 334192 518052 334248
rect 433977 334190 518052 334192
rect 433977 334187 434043 334190
rect 377489 332890 377555 332893
rect 377489 332888 518052 332890
rect 377489 332832 377494 332888
rect 377550 332832 518052 332888
rect 377489 332830 518052 332832
rect 377489 332827 377555 332830
rect -960 332196 480 332436
rect 304717 331530 304783 331533
rect 304717 331528 518052 331530
rect 304717 331472 304722 331528
rect 304778 331472 518052 331528
rect 304717 331470 518052 331472
rect 304717 331467 304783 331470
rect 529933 330986 529999 330989
rect 527804 330984 529999 330986
rect 527804 330928 529938 330984
rect 529994 330928 529999 330984
rect 527804 330926 529999 330928
rect 529933 330923 529999 330926
rect 515857 330170 515923 330173
rect 515857 330168 518052 330170
rect 515857 330112 515862 330168
rect 515918 330112 518052 330168
rect 515857 330110 518052 330112
rect 515857 330107 515923 330110
rect 515673 328810 515739 328813
rect 515673 328808 518052 328810
rect 515673 328752 515678 328808
rect 515734 328752 518052 328808
rect 515673 328750 518052 328752
rect 515673 328747 515739 328750
rect 310973 328402 311039 328405
rect 311893 328402 311959 328405
rect 310973 328400 311959 328402
rect 310973 328344 310978 328400
rect 311034 328344 311898 328400
rect 311954 328344 311959 328400
rect 310973 328342 311959 328344
rect 310973 328339 311039 328342
rect 311893 328339 311959 328342
rect 304901 327722 304967 327725
rect 310973 327722 311039 327725
rect 304901 327720 311039 327722
rect 304901 327664 304906 327720
rect 304962 327664 310978 327720
rect 311034 327664 311039 327720
rect 304901 327662 311039 327664
rect 304901 327659 304967 327662
rect 310973 327659 311039 327662
rect 373257 327450 373323 327453
rect 373257 327448 518052 327450
rect 373257 327392 373262 327448
rect 373318 327392 518052 327448
rect 373257 327390 518052 327392
rect 373257 327387 373323 327390
rect 295241 327178 295307 327181
rect 300853 327178 300919 327181
rect 295241 327176 300919 327178
rect 295241 327120 295246 327176
rect 295302 327120 300858 327176
rect 300914 327120 300919 327176
rect 295241 327118 300919 327120
rect 295241 327115 295307 327118
rect 300853 327115 300919 327118
rect 307661 326226 307727 326229
rect 311985 326226 312051 326229
rect 307661 326224 312051 326226
rect 307661 326168 307666 326224
rect 307722 326168 311990 326224
rect 312046 326168 312051 326224
rect 307661 326166 312051 326168
rect 307661 326163 307727 326166
rect 311985 326163 312051 326166
rect 318425 326090 318491 326093
rect 318425 326088 518052 326090
rect 296878 326084 297194 326085
rect 296878 326020 296884 326084
rect 296948 326020 296964 326084
rect 297028 326020 297044 326084
rect 297108 326020 297124 326084
rect 297188 326020 297194 326084
rect 296878 326004 297194 326020
rect 296878 325940 296884 326004
rect 296948 325940 296964 326004
rect 297028 325940 297044 326004
rect 297108 325940 297124 326004
rect 297188 325940 297194 326004
rect 303878 326084 304194 326085
rect 303878 326020 303884 326084
rect 303948 326020 303964 326084
rect 304028 326020 304044 326084
rect 304108 326020 304124 326084
rect 304188 326020 304194 326084
rect 303878 326004 304194 326020
rect 296878 325924 297194 325940
rect 296878 325860 296884 325924
rect 296948 325860 296964 325924
rect 297028 325860 297044 325924
rect 297108 325860 297124 325924
rect 297188 325860 297194 325924
rect 300853 325954 300919 325957
rect 300853 325952 300962 325954
rect 300853 325896 300858 325952
rect 300914 325896 300962 325952
rect 300853 325891 300962 325896
rect 296878 325844 297194 325860
rect 296878 325780 296884 325844
rect 296948 325780 296964 325844
rect 297028 325780 297044 325844
rect 297108 325780 297124 325844
rect 297188 325780 297194 325844
rect 296878 325779 297194 325780
rect 300902 325685 300962 325891
rect 303878 325940 303884 326004
rect 303948 325940 303964 326004
rect 304028 325940 304044 326004
rect 304108 325940 304124 326004
rect 304188 325940 304194 326004
rect 310878 326084 311194 326085
rect 310878 326020 310884 326084
rect 310948 326020 310964 326084
rect 311028 326020 311044 326084
rect 311108 326020 311124 326084
rect 311188 326020 311194 326084
rect 318425 326032 318430 326088
rect 318486 326032 518052 326088
rect 318425 326030 518052 326032
rect 318425 326027 318491 326030
rect 310878 326004 311194 326020
rect 304901 325954 304967 325957
rect 307661 325954 307727 325957
rect 303878 325924 304194 325940
rect 303878 325860 303884 325924
rect 303948 325860 303964 325924
rect 304028 325860 304044 325924
rect 304108 325860 304124 325924
rect 304188 325860 304194 325924
rect 303878 325844 304194 325860
rect 303878 325780 303884 325844
rect 303948 325780 303964 325844
rect 304028 325780 304044 325844
rect 304108 325780 304124 325844
rect 304188 325780 304194 325844
rect 303878 325779 304194 325780
rect 304398 325952 304967 325954
rect 304398 325896 304906 325952
rect 304962 325896 304967 325952
rect 304398 325894 304967 325896
rect 300902 325680 301011 325685
rect 300902 325624 300950 325680
rect 301006 325624 301011 325680
rect 300902 325622 301011 325624
rect 300945 325619 301011 325622
rect 304257 325682 304323 325685
rect 304398 325682 304458 325894
rect 304901 325891 304967 325894
rect 307526 325952 307727 325954
rect 307526 325896 307666 325952
rect 307722 325896 307727 325952
rect 307526 325894 307727 325896
rect 304257 325680 304458 325682
rect 304257 325624 304262 325680
rect 304318 325624 304458 325680
rect 304257 325622 304458 325624
rect 307385 325682 307451 325685
rect 307526 325682 307586 325894
rect 307661 325891 307727 325894
rect 310878 325940 310884 326004
rect 310948 325940 310964 326004
rect 311028 325940 311044 326004
rect 311108 325940 311124 326004
rect 311188 325940 311194 326004
rect 310878 325924 311194 325940
rect 310878 325860 310884 325924
rect 310948 325860 310964 325924
rect 311028 325860 311044 325924
rect 311108 325860 311124 325924
rect 311188 325860 311194 325924
rect 310878 325844 311194 325860
rect 310878 325780 310884 325844
rect 310948 325780 310964 325844
rect 311028 325780 311044 325844
rect 311108 325780 311124 325844
rect 311188 325780 311194 325844
rect 310878 325779 311194 325780
rect 307385 325680 307586 325682
rect 307385 325624 307390 325680
rect 307446 325624 307586 325680
rect 307385 325622 307586 325624
rect 304257 325619 304323 325622
rect 307385 325619 307451 325622
rect 583520 325124 584960 325364
rect 312629 325002 312695 325005
rect 515489 325002 515555 325005
rect 312629 325000 515555 325002
rect 312629 324944 312634 325000
rect 312690 324944 515494 325000
rect 515550 324944 515555 325000
rect 312629 324942 515555 324944
rect 312629 324939 312695 324942
rect 515489 324939 515555 324942
rect 515765 324730 515831 324733
rect 515765 324728 518052 324730
rect 515765 324672 515770 324728
rect 515826 324672 518052 324728
rect 515765 324670 518052 324672
rect 515765 324667 515831 324670
rect 303878 323912 304194 323913
rect 303878 323848 303884 323912
rect 303948 323848 303964 323912
rect 304028 323848 304044 323912
rect 304108 323848 304124 323912
rect 304188 323848 304194 323912
rect 303878 323832 304194 323848
rect 303878 323768 303884 323832
rect 303948 323768 303964 323832
rect 304028 323768 304044 323832
rect 304108 323768 304124 323832
rect 304188 323768 304194 323832
rect 303878 323752 304194 323768
rect 303878 323688 303884 323752
rect 303948 323688 303964 323752
rect 304028 323688 304044 323752
rect 304108 323688 304124 323752
rect 304188 323688 304194 323752
rect 303878 323672 304194 323688
rect 303878 323608 303884 323672
rect 303948 323608 303964 323672
rect 304028 323608 304044 323672
rect 304108 323608 304124 323672
rect 304188 323608 304194 323672
rect 303878 323607 304194 323608
rect 310878 323912 311194 323913
rect 310878 323848 310884 323912
rect 310948 323848 310964 323912
rect 311028 323848 311044 323912
rect 311108 323848 311124 323912
rect 311188 323848 311194 323912
rect 310878 323832 311194 323848
rect 310878 323768 310884 323832
rect 310948 323768 310964 323832
rect 311028 323768 311044 323832
rect 311108 323768 311124 323832
rect 311188 323768 311194 323832
rect 310878 323752 311194 323768
rect 310878 323688 310884 323752
rect 310948 323688 310964 323752
rect 311028 323688 311044 323752
rect 311108 323688 311124 323752
rect 311188 323688 311194 323752
rect 310878 323672 311194 323688
rect 310878 323608 310884 323672
rect 310948 323608 310964 323672
rect 311028 323608 311044 323672
rect 311108 323608 311124 323672
rect 311188 323608 311194 323672
rect 310878 323607 311194 323608
rect 311390 323098 311450 323612
rect 318333 323370 318399 323373
rect 318333 323368 518052 323370
rect 318333 323312 318338 323368
rect 318394 323312 518052 323368
rect 318333 323310 518052 323312
rect 318333 323307 318399 323310
rect 314193 323098 314259 323101
rect 311390 323096 314259 323098
rect 311390 323040 314198 323096
rect 314254 323040 314259 323096
rect 311390 323038 314259 323040
rect 314193 323035 314259 323038
rect 305085 322826 305151 322829
rect 515857 322826 515923 322829
rect 305085 322824 515923 322826
rect 305085 322768 305090 322824
rect 305146 322768 515862 322824
rect 515918 322768 515923 322824
rect 305085 322766 515923 322768
rect 305085 322763 305151 322766
rect 515857 322763 515923 322766
rect 371877 322010 371943 322013
rect 371877 322008 518052 322010
rect 371877 321952 371882 322008
rect 371938 321952 518052 322008
rect 371877 321950 518052 321952
rect 371877 321947 371943 321950
rect 298737 321466 298803 321469
rect 515397 321466 515463 321469
rect 298737 321464 515463 321466
rect 298737 321408 298742 321464
rect 298798 321408 515402 321464
rect 515458 321408 515463 321464
rect 298737 321406 515463 321408
rect 298737 321403 298803 321406
rect 515397 321403 515463 321406
rect 301773 321330 301839 321333
rect 515581 321330 515647 321333
rect 301773 321328 515647 321330
rect 301773 321272 301778 321328
rect 301834 321272 515586 321328
rect 515642 321272 515647 321328
rect 301773 321270 515647 321272
rect 301773 321267 301839 321270
rect 515581 321267 515647 321270
rect 329097 320650 329163 320653
rect 329097 320648 518052 320650
rect 329097 320592 329102 320648
rect 329158 320592 518052 320648
rect 329097 320590 518052 320592
rect 329097 320587 329163 320590
rect 517421 319426 517487 319429
rect 522297 319426 522363 319429
rect 517421 319424 522363 319426
rect -960 319140 480 319380
rect 517421 319368 517426 319424
rect 517482 319368 522302 319424
rect 522358 319368 522363 319424
rect 517421 319366 522363 319368
rect 517421 319363 517487 319366
rect 522297 319363 522363 319366
rect 583520 311932 584960 312172
rect 308213 308410 308279 308413
rect 384389 308410 384455 308413
rect 308213 308408 384455 308410
rect 308213 308352 308218 308408
rect 308274 308352 384394 308408
rect 384450 308352 384455 308408
rect 308213 308350 384455 308352
rect 308213 308347 308279 308350
rect 384389 308347 384455 308350
rect 306189 307458 306255 307461
rect 311893 307458 311959 307461
rect 313733 307458 313799 307461
rect 306189 307456 313799 307458
rect 306189 307400 306194 307456
rect 306250 307400 311898 307456
rect 311954 307400 313738 307456
rect 313794 307400 313799 307456
rect 306189 307398 313799 307400
rect 306189 307395 306255 307398
rect 311893 307395 311959 307398
rect 313733 307395 313799 307398
rect 312905 307186 312971 307189
rect 515397 307186 515463 307189
rect 312905 307184 515463 307186
rect 312905 307128 312910 307184
rect 312966 307128 515402 307184
rect 515458 307128 515463 307184
rect 312905 307126 515463 307128
rect 312905 307123 312971 307126
rect 515397 307123 515463 307126
rect 312537 307050 312603 307053
rect 515581 307050 515647 307053
rect 312537 307048 515647 307050
rect 312537 306992 312542 307048
rect 312598 306992 515586 307048
rect 515642 306992 515647 307048
rect 312537 306990 515647 306992
rect 312537 306987 312603 306990
rect 515581 306987 515647 306990
rect 295241 306506 295307 306509
rect 301681 306506 301747 306509
rect 295241 306504 301747 306506
rect 295241 306448 295246 306504
rect 295302 306448 301686 306504
rect 301742 306448 301747 306504
rect 295241 306446 301747 306448
rect 295241 306443 295307 306446
rect 301681 306443 301747 306446
rect 311985 306506 312051 306509
rect 313641 306506 313707 306509
rect 311985 306504 313707 306506
rect 311985 306448 311990 306504
rect 312046 306448 313646 306504
rect 313702 306448 313707 306504
rect 311985 306446 313707 306448
rect 311985 306443 312051 306446
rect 313641 306443 313707 306446
rect -960 306084 480 306324
rect 296878 305114 297194 305115
rect 296878 305050 296884 305114
rect 296948 305050 296964 305114
rect 297028 305050 297044 305114
rect 297108 305050 297124 305114
rect 297188 305050 297194 305114
rect 296878 305034 297194 305050
rect 296878 304970 296884 305034
rect 296948 304970 296964 305034
rect 297028 304970 297044 305034
rect 297108 304970 297124 305034
rect 297188 304970 297194 305034
rect 303878 305114 304194 305115
rect 303878 305050 303884 305114
rect 303948 305050 303964 305114
rect 304028 305050 304044 305114
rect 304108 305050 304124 305114
rect 304188 305050 304194 305114
rect 303878 305034 304194 305050
rect 296878 304954 297194 304970
rect 296878 304890 296884 304954
rect 296948 304890 296964 304954
rect 297028 304890 297044 304954
rect 297108 304890 297124 304954
rect 297188 304890 297194 304954
rect 301681 305008 301747 305013
rect 301681 304952 301686 305008
rect 301742 304952 301747 305008
rect 301681 304947 301747 304952
rect 303878 304970 303884 305034
rect 303948 304970 303964 305034
rect 304028 304970 304044 305034
rect 304108 304970 304124 305034
rect 304188 304970 304194 305034
rect 310878 305114 311194 305115
rect 310878 305050 310884 305114
rect 310948 305050 310964 305114
rect 311028 305050 311044 305114
rect 311108 305050 311124 305114
rect 311188 305050 311194 305114
rect 310878 305034 311194 305050
rect 306189 305010 306255 305013
rect 303878 304954 304194 304970
rect 296878 304874 297194 304890
rect 296878 304810 296884 304874
rect 296948 304810 296964 304874
rect 297028 304810 297044 304874
rect 297108 304810 297124 304874
rect 297188 304810 297194 304874
rect 296878 304809 297194 304810
rect 301684 304602 301744 304947
rect 303878 304890 303884 304954
rect 303948 304890 303964 304954
rect 304028 304890 304044 304954
rect 304108 304890 304124 304954
rect 304188 304890 304194 304954
rect 303878 304874 304194 304890
rect 303878 304810 303884 304874
rect 303948 304810 303964 304874
rect 304028 304810 304044 304874
rect 304108 304810 304124 304874
rect 304188 304810 304194 304874
rect 303878 304809 304194 304810
rect 306054 305008 306255 305010
rect 306054 304952 306194 305008
rect 306250 304952 306255 305008
rect 306054 304950 306255 304952
rect 301951 304602 302017 304605
rect 301684 304600 302017 304602
rect 301684 304544 301956 304600
rect 302012 304544 302017 304600
rect 301684 304542 302017 304544
rect 301951 304539 302017 304542
rect 305545 304602 305611 304605
rect 306054 304602 306114 304950
rect 306189 304947 306255 304950
rect 310605 305008 310671 305013
rect 310605 304952 310610 305008
rect 310666 304952 310671 305008
rect 310605 304947 310671 304952
rect 310878 304970 310884 305034
rect 310948 304970 310964 305034
rect 311028 304970 311044 305034
rect 311108 304970 311124 305034
rect 311188 304970 311194 305034
rect 310878 304954 311194 304970
rect 310608 304738 310668 304947
rect 310878 304890 310884 304954
rect 310948 304890 310964 304954
rect 311028 304890 311044 304954
rect 311108 304890 311124 304954
rect 311188 304890 311194 304954
rect 310878 304874 311194 304890
rect 310878 304810 310884 304874
rect 310948 304810 310964 304874
rect 311028 304810 311044 304874
rect 311108 304810 311124 304874
rect 311188 304810 311194 304874
rect 310878 304809 311194 304810
rect 310608 304678 312416 304738
rect 312356 304605 312416 304678
rect 305545 304600 306114 304602
rect 305545 304544 305550 304600
rect 305606 304544 306114 304600
rect 305545 304542 306114 304544
rect 312353 304600 312419 304605
rect 312353 304544 312358 304600
rect 312414 304544 312419 304600
rect 305545 304539 305611 304542
rect 312353 304539 312419 304544
rect 319713 304330 319779 304333
rect 515857 304330 515923 304333
rect 319713 304328 515923 304330
rect 319713 304272 319718 304328
rect 319774 304272 515862 304328
rect 515918 304272 515923 304328
rect 319713 304270 515923 304272
rect 319713 304267 319779 304270
rect 515857 304267 515923 304270
rect 319529 304194 319595 304197
rect 514753 304194 514819 304197
rect 319529 304192 514819 304194
rect 319529 304136 319534 304192
rect 319590 304136 514758 304192
rect 514814 304136 514819 304192
rect 319529 304134 514819 304136
rect 319529 304131 319595 304134
rect 514753 304131 514819 304134
rect 302146 304013 302462 304014
rect 302146 303949 302152 304013
rect 302216 303949 302232 304013
rect 302296 303949 302312 304013
rect 302376 303949 302392 304013
rect 302456 303949 302462 304013
rect 302146 303933 302462 303949
rect 302146 303869 302152 303933
rect 302216 303869 302232 303933
rect 302296 303869 302312 303933
rect 302376 303869 302392 303933
rect 302456 303869 302462 303933
rect 302146 303853 302462 303869
rect 302146 303789 302152 303853
rect 302216 303789 302232 303853
rect 302296 303789 302312 303853
rect 302376 303789 302392 303853
rect 302456 303789 302462 303853
rect 302146 303773 302462 303789
rect 302146 303709 302152 303773
rect 302216 303709 302232 303773
rect 302296 303709 302312 303773
rect 302376 303709 302392 303773
rect 302456 303709 302462 303773
rect 302146 303708 302462 303709
rect 309146 304013 309462 304014
rect 309146 303949 309152 304013
rect 309216 303949 309232 304013
rect 309296 303949 309312 304013
rect 309376 303949 309392 304013
rect 309456 303949 309462 304013
rect 309146 303933 309462 303949
rect 309146 303869 309152 303933
rect 309216 303869 309232 303933
rect 309296 303869 309312 303933
rect 309376 303869 309392 303933
rect 309456 303869 309462 303933
rect 309146 303853 309462 303869
rect 309146 303789 309152 303853
rect 309216 303789 309232 303853
rect 309296 303789 309312 303853
rect 309376 303789 309392 303853
rect 309456 303789 309462 303853
rect 309146 303773 309462 303789
rect 309146 303709 309152 303773
rect 309216 303709 309232 303773
rect 309296 303709 309312 303773
rect 309376 303709 309392 303773
rect 309456 303709 309462 303773
rect 527081 303786 527147 303789
rect 528553 303786 528619 303789
rect 527081 303784 528619 303786
rect 527081 303728 527086 303784
rect 527142 303728 528558 303784
rect 528614 303728 528619 303784
rect 527081 303726 528619 303728
rect 527081 303723 527147 303726
rect 528553 303723 528619 303726
rect 309146 303708 309462 303709
rect 524321 303650 524387 303653
rect 527265 303650 527331 303653
rect 524321 303648 527331 303650
rect 524321 303592 524326 303648
rect 524382 303592 527270 303648
rect 527326 303592 527331 303648
rect 524321 303590 527331 303592
rect 524321 303587 524387 303590
rect 527265 303587 527331 303590
rect 313365 303514 313431 303517
rect 317137 303514 317203 303517
rect 313365 303512 317203 303514
rect 313365 303456 313370 303512
rect 313426 303456 317142 303512
rect 317198 303456 317203 303512
rect 313365 303454 317203 303456
rect 313365 303451 313431 303454
rect 317137 303451 317203 303454
rect 515673 302834 515739 302837
rect 321510 302832 515739 302834
rect 321510 302776 515678 302832
rect 515734 302776 515739 302832
rect 321510 302774 515739 302776
rect 321510 302426 321570 302774
rect 515673 302771 515739 302774
rect 313230 302366 321570 302426
rect 306373 302154 306439 302157
rect 313230 302154 313290 302366
rect 522113 302290 522179 302293
rect 528645 302290 528711 302293
rect 580165 302290 580231 302293
rect 522113 302288 580231 302290
rect 522113 302232 522118 302288
rect 522174 302232 528650 302288
rect 528706 302232 580170 302288
rect 580226 302232 580231 302288
rect 522113 302230 580231 302232
rect 522113 302227 522179 302230
rect 528645 302227 528711 302230
rect 580165 302227 580231 302230
rect 306373 302152 313290 302154
rect 306373 302096 306378 302152
rect 306434 302096 313290 302152
rect 306373 302094 313290 302096
rect 306373 302091 306439 302094
rect 299197 302018 299263 302021
rect 317045 302018 317111 302021
rect 299197 302016 317111 302018
rect 299197 301960 299202 302016
rect 299258 301960 317050 302016
rect 317106 301960 317111 302016
rect 299197 301958 317111 301960
rect 299197 301955 299263 301958
rect 317045 301955 317111 301958
rect 302785 301882 302851 301885
rect 370497 301882 370563 301885
rect 302785 301880 370563 301882
rect 302785 301824 302790 301880
rect 302846 301824 370502 301880
rect 370558 301824 370563 301880
rect 302785 301822 370563 301824
rect 302785 301819 302851 301822
rect 370497 301819 370563 301822
rect 318241 301066 318307 301069
rect 318241 301064 518052 301066
rect 318241 301008 318246 301064
rect 318302 301008 518052 301064
rect 318241 301006 518052 301008
rect 318241 301003 318307 301006
rect 514753 299706 514819 299709
rect 514753 299704 518052 299706
rect 514753 299648 514758 299704
rect 514814 299648 518052 299704
rect 514753 299646 518052 299648
rect 514753 299643 514819 299646
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 464337 298346 464403 298349
rect 464337 298344 518052 298346
rect 464337 298288 464342 298344
rect 464398 298288 518052 298344
rect 464337 298286 518052 298288
rect 464337 298283 464403 298286
rect 377397 296986 377463 296989
rect 377397 296984 518052 296986
rect 377397 296928 377402 296984
rect 377458 296928 518052 296984
rect 377397 296926 518052 296928
rect 377397 296923 377463 296926
rect 515857 295626 515923 295629
rect 515857 295624 518052 295626
rect 515857 295568 515862 295624
rect 515918 295568 518052 295624
rect 515857 295566 518052 295568
rect 515857 295563 515923 295566
rect 295241 294538 295307 294541
rect 299473 294538 299539 294541
rect 295241 294536 299539 294538
rect 295241 294480 295246 294536
rect 295302 294480 299478 294536
rect 299534 294480 299539 294536
rect 295241 294478 299539 294480
rect 295241 294475 295307 294478
rect 299473 294475 299539 294478
rect 515581 294266 515647 294269
rect 515581 294264 518052 294266
rect 515581 294208 515586 294264
rect 515642 294208 518052 294264
rect 515581 294206 518052 294208
rect 515581 294203 515647 294206
rect -960 293028 480 293268
rect 515397 292906 515463 292909
rect 515397 292904 518052 292906
rect 515397 292848 515402 292904
rect 515458 292848 518052 292904
rect 515397 292846 518052 292848
rect 515397 292843 515463 292846
rect 515489 291546 515555 291549
rect 515489 291544 518052 291546
rect 515489 291488 515494 291544
rect 515550 291488 518052 291544
rect 515489 291486 518052 291488
rect 515489 291483 515555 291486
rect 529933 291002 529999 291005
rect 527804 291000 529999 291002
rect 527804 290944 529938 291000
rect 529994 290944 529999 291000
rect 527804 290942 529999 290944
rect 529933 290939 529999 290942
rect 384389 290186 384455 290189
rect 384389 290184 518052 290186
rect 384389 290128 384394 290184
rect 384450 290128 518052 290184
rect 384389 290126 518052 290128
rect 384389 290123 384455 290126
rect 309961 288826 310027 288829
rect 309961 288824 518052 288826
rect 309961 288768 309966 288824
rect 310022 288768 518052 288824
rect 309961 288766 518052 288768
rect 309961 288763 310027 288766
rect 311893 288418 311959 288421
rect 313733 288418 313799 288421
rect 311893 288416 313799 288418
rect 311893 288360 311898 288416
rect 311954 288360 313738 288416
rect 313794 288360 313799 288416
rect 311893 288358 313799 288360
rect 311893 288355 311959 288358
rect 313733 288355 313799 288358
rect 515673 287466 515739 287469
rect 515673 287464 518052 287466
rect 515673 287408 515678 287464
rect 515734 287408 518052 287464
rect 515673 287406 518052 287408
rect 515673 287403 515739 287406
rect 515581 286106 515647 286109
rect 515581 286104 518052 286106
rect 515581 286048 515586 286104
rect 515642 286048 518052 286104
rect 515581 286046 518052 286048
rect 515581 286043 515647 286046
rect 308121 285970 308187 285973
rect 312721 285970 312787 285973
rect 314469 285970 314535 285973
rect 308121 285968 314535 285970
rect 308121 285912 308126 285968
rect 308182 285912 312726 285968
rect 312782 285912 314474 285968
rect 314530 285912 314535 285968
rect 308121 285910 314535 285912
rect 308121 285907 308187 285910
rect 312721 285907 312787 285910
rect 314469 285907 314535 285910
rect 304809 285834 304875 285837
rect 312353 285834 312419 285837
rect 304809 285832 312419 285834
rect 304809 285776 304814 285832
rect 304870 285776 312358 285832
rect 312414 285776 312419 285832
rect 304809 285774 312419 285776
rect 304809 285771 304875 285774
rect 312353 285771 312419 285774
rect 312629 285698 312695 285701
rect 313825 285698 313891 285701
rect 312629 285696 313891 285698
rect 312629 285640 312634 285696
rect 312690 285640 313830 285696
rect 313886 285640 313891 285696
rect 312629 285638 313891 285640
rect 312629 285635 312695 285638
rect 313825 285635 313891 285638
rect 583520 285276 584960 285516
rect 514753 284746 514819 284749
rect 514753 284744 518052 284746
rect 514753 284688 514758 284744
rect 514814 284688 518052 284744
rect 514753 284686 518052 284688
rect 514753 284683 514819 284686
rect 295241 284474 295307 284477
rect 299473 284474 299539 284477
rect 295241 284472 299539 284474
rect 295241 284416 295246 284472
rect 295302 284416 299478 284472
rect 299534 284416 299539 284472
rect 295241 284414 299539 284416
rect 295241 284411 295307 284414
rect 299473 284411 299539 284414
rect 295241 284338 295307 284341
rect 298093 284338 298159 284341
rect 295241 284336 298202 284338
rect 295241 284280 295246 284336
rect 295302 284280 298098 284336
rect 298154 284280 298202 284336
rect 295241 284278 298202 284280
rect 295241 284275 295307 284278
rect 298093 284275 298202 284278
rect 298142 283389 298202 284275
rect 299473 283794 299539 283797
rect 304809 283794 304875 283797
rect 308121 283794 308187 283797
rect 299246 283792 299539 283794
rect 299246 283736 299478 283792
rect 299534 283736 299539 283792
rect 299246 283734 299539 283736
rect 298137 283384 298203 283389
rect 298137 283328 298142 283384
rect 298198 283328 298203 283384
rect 298137 283323 298203 283328
rect 299246 283386 299306 283734
rect 299473 283731 299539 283734
rect 304766 283792 304875 283794
rect 304766 283736 304814 283792
rect 304870 283736 304875 283792
rect 304766 283731 304875 283736
rect 308078 283792 308187 283794
rect 308078 283736 308126 283792
rect 308182 283736 308187 283792
rect 308078 283731 308187 283736
rect 304766 283389 304826 283731
rect 308078 283389 308138 283731
rect 299749 283386 299815 283389
rect 299246 283384 299815 283386
rect 299246 283328 299754 283384
rect 299810 283328 299815 283384
rect 299246 283326 299815 283328
rect 304766 283384 304837 283389
rect 304766 283328 304776 283384
rect 304832 283328 304837 283384
rect 304766 283326 304837 283328
rect 308078 283384 308154 283389
rect 308078 283328 308093 283384
rect 308149 283328 308154 283384
rect 308078 283326 308154 283328
rect 299749 283323 299815 283326
rect 304771 283323 304837 283326
rect 308088 283323 308154 283326
rect 317045 283386 317111 283389
rect 317045 283384 518052 283386
rect 317045 283328 317050 283384
rect 317106 283328 518052 283384
rect 317045 283326 518052 283328
rect 317045 283323 317111 283326
rect 309146 282999 309462 283000
rect 302146 282998 302462 282999
rect 302146 282934 302152 282998
rect 302216 282934 302232 282998
rect 302296 282934 302312 282998
rect 302376 282934 302392 282998
rect 302456 282934 302462 282998
rect 302146 282918 302462 282934
rect 302146 282854 302152 282918
rect 302216 282854 302232 282918
rect 302296 282854 302312 282918
rect 302376 282854 302392 282918
rect 302456 282854 302462 282918
rect 302146 282838 302462 282854
rect 302146 282774 302152 282838
rect 302216 282774 302232 282838
rect 302296 282774 302312 282838
rect 302376 282774 302392 282838
rect 302456 282774 302462 282838
rect 302146 282758 302462 282774
rect 302146 282694 302152 282758
rect 302216 282694 302232 282758
rect 302296 282694 302312 282758
rect 302376 282694 302392 282758
rect 302456 282694 302462 282758
rect 309146 282935 309152 282999
rect 309216 282935 309232 282999
rect 309296 282935 309312 282999
rect 309376 282935 309392 282999
rect 309456 282935 309462 282999
rect 309146 282919 309462 282935
rect 309146 282855 309152 282919
rect 309216 282855 309232 282919
rect 309296 282855 309312 282919
rect 309376 282855 309392 282919
rect 309456 282855 309462 282919
rect 309146 282839 309462 282855
rect 309146 282775 309152 282839
rect 309216 282775 309232 282839
rect 309296 282775 309312 282839
rect 309376 282775 309392 282839
rect 309456 282775 309462 282839
rect 309146 282759 309462 282775
rect 309146 282695 309152 282759
rect 309216 282695 309232 282759
rect 309296 282695 309312 282759
rect 309376 282695 309392 282759
rect 309456 282695 309462 282759
rect 309146 282694 309462 282695
rect 302146 282693 302462 282694
rect 303878 282237 304194 282238
rect 303878 282173 303884 282237
rect 303948 282173 303964 282237
rect 304028 282173 304044 282237
rect 304108 282173 304124 282237
rect 304188 282173 304194 282237
rect 303878 282157 304194 282173
rect 303878 282093 303884 282157
rect 303948 282093 303964 282157
rect 304028 282093 304044 282157
rect 304108 282093 304124 282157
rect 304188 282093 304194 282157
rect 303878 282077 304194 282093
rect 303878 282013 303884 282077
rect 303948 282013 303964 282077
rect 304028 282013 304044 282077
rect 304108 282013 304124 282077
rect 304188 282013 304194 282077
rect 303878 281997 304194 282013
rect 303878 281933 303884 281997
rect 303948 281933 303964 281997
rect 304028 281933 304044 281997
rect 304108 281933 304124 281997
rect 304188 281933 304194 281997
rect 303878 281917 304194 281933
rect 303878 281853 303884 281917
rect 303948 281853 303964 281917
rect 304028 281853 304044 281917
rect 304108 281853 304124 281917
rect 304188 281853 304194 281917
rect 303878 281837 304194 281853
rect 303878 281773 303884 281837
rect 303948 281773 303964 281837
rect 304028 281773 304044 281837
rect 304108 281773 304124 281837
rect 304188 281773 304194 281837
rect 303878 281757 304194 281773
rect 303878 281693 303884 281757
rect 303948 281693 303964 281757
rect 304028 281693 304044 281757
rect 304108 281693 304124 281757
rect 304188 281693 304194 281757
rect 303878 281677 304194 281693
rect 303878 281613 303884 281677
rect 303948 281613 303964 281677
rect 304028 281613 304044 281677
rect 304108 281613 304124 281677
rect 304188 281613 304194 281677
rect 310878 282182 311194 282183
rect 310878 282118 310884 282182
rect 310948 282118 310964 282182
rect 311028 282118 311044 282182
rect 311108 282118 311124 282182
rect 311188 282118 311194 282182
rect 382917 282162 382983 282165
rect 310878 282102 311194 282118
rect 310878 282038 310884 282102
rect 310948 282038 310964 282102
rect 311028 282038 311044 282102
rect 311108 282038 311124 282102
rect 311188 282038 311194 282102
rect 310878 282022 311194 282038
rect 315990 282160 382983 282162
rect 315990 282104 382922 282160
rect 382978 282104 382983 282160
rect 315990 282102 382983 282104
rect 310878 281958 310884 282022
rect 310948 281958 310964 282022
rect 311028 281958 311044 282022
rect 311108 281958 311124 282022
rect 311188 281958 311194 282022
rect 312537 282026 312603 282029
rect 315990 282026 316050 282102
rect 382917 282099 382983 282102
rect 312537 282024 316050 282026
rect 312537 281968 312542 282024
rect 312598 281968 316050 282024
rect 312537 281966 316050 281968
rect 515489 282026 515555 282029
rect 515489 282024 518052 282026
rect 515489 281968 515494 282024
rect 515550 281968 518052 282024
rect 515489 281966 518052 281968
rect 312537 281963 312603 281966
rect 515489 281963 515555 281966
rect 310878 281942 311194 281958
rect 310878 281878 310884 281942
rect 310948 281878 310964 281942
rect 311028 281878 311044 281942
rect 311108 281878 311124 281942
rect 311188 281878 311194 281942
rect 310878 281862 311194 281878
rect 310878 281798 310884 281862
rect 310948 281798 310964 281862
rect 311028 281798 311044 281862
rect 311108 281798 311124 281862
rect 311188 281798 311194 281862
rect 310878 281782 311194 281798
rect 310878 281718 310884 281782
rect 310948 281718 310964 281782
rect 311028 281718 311044 281782
rect 311108 281718 311124 281782
rect 311188 281718 311194 281782
rect 310878 281702 311194 281718
rect 310878 281638 310884 281702
rect 310948 281638 310964 281702
rect 311028 281638 311044 281702
rect 311108 281638 311124 281702
rect 311188 281638 311194 281702
rect 310878 281637 311194 281638
rect 303878 281612 304194 281613
rect 305729 281482 305795 281485
rect 373257 281482 373323 281485
rect 305729 281480 373323 281482
rect 305729 281424 305734 281480
rect 305790 281424 373262 281480
rect 373318 281424 373323 281480
rect 305729 281422 373323 281424
rect 305729 281419 305795 281422
rect 373257 281419 373323 281422
rect 299105 281346 299171 281349
rect 315757 281346 315823 281349
rect 299105 281344 315823 281346
rect 299105 281288 299110 281344
rect 299166 281288 315762 281344
rect 315818 281288 315823 281344
rect 299105 281286 315823 281288
rect 299105 281283 299171 281286
rect 315757 281283 315823 281286
rect 515397 280666 515463 280669
rect 515397 280664 518052 280666
rect 515397 280608 515402 280664
rect 515458 280608 518052 280664
rect 515397 280606 518052 280608
rect 515397 280603 515463 280606
rect -960 279972 480 280212
rect 308949 280122 309015 280125
rect 515673 280122 515739 280125
rect 308949 280120 515739 280122
rect 308949 280064 308954 280120
rect 309010 280064 515678 280120
rect 515734 280064 515739 280120
rect 308949 280062 515739 280064
rect 308949 280059 309015 280062
rect 515673 280059 515739 280062
rect 302417 279986 302483 279989
rect 326337 279986 326403 279989
rect 302417 279984 326403 279986
rect 302417 279928 302422 279984
rect 302478 279928 326342 279984
rect 326398 279928 326403 279984
rect 302417 279926 326403 279928
rect 302417 279923 302483 279926
rect 326337 279923 326403 279926
rect 518617 278898 518683 278901
rect 519537 278898 519603 278901
rect 518617 278896 519603 278898
rect 518617 278840 518622 278896
rect 518678 278840 519542 278896
rect 519598 278840 519603 278896
rect 518617 278838 519603 278840
rect 518617 278835 518683 278838
rect 519537 278835 519603 278838
rect 295241 277538 295307 277541
rect 298185 277538 298251 277541
rect 295241 277536 298251 277538
rect 295241 277480 295246 277536
rect 295302 277480 298190 277536
rect 298246 277480 298251 277536
rect 295241 277478 298251 277480
rect 295241 277475 295307 277478
rect 298185 277475 298251 277478
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 308765 265162 308831 265165
rect 308765 265160 312554 265162
rect 308765 265104 308770 265160
rect 308826 265104 312554 265160
rect 308765 265102 312554 265104
rect 308765 265099 308831 265102
rect 312494 265029 312554 265102
rect 295241 265026 295307 265029
rect 299473 265026 299539 265029
rect 295241 265024 299539 265026
rect 295241 264968 295246 265024
rect 295302 264968 299478 265024
rect 299534 264968 299539 265024
rect 295241 264966 299539 264968
rect 295241 264963 295307 264966
rect 299473 264963 299539 264966
rect 305085 265026 305151 265029
rect 312353 265026 312419 265029
rect 305085 265024 312419 265026
rect 305085 264968 305090 265024
rect 305146 264968 312358 265024
rect 312414 264968 312419 265024
rect 305085 264966 312419 264968
rect 312494 265026 312603 265029
rect 313273 265026 313339 265029
rect 312494 265024 313339 265026
rect 312494 264968 312542 265024
rect 312598 264968 313278 265024
rect 313334 264968 313339 265024
rect 312494 264966 313339 264968
rect 305085 264963 305151 264966
rect 312353 264963 312419 264966
rect 312537 264963 312603 264966
rect 313273 264963 313339 264966
rect 527081 264890 527147 264893
rect 528553 264890 528619 264893
rect 527081 264888 528619 264890
rect 527081 264832 527086 264888
rect 527142 264832 528558 264888
rect 528614 264832 528619 264888
rect 527081 264830 528619 264832
rect 527081 264827 527147 264830
rect 528553 264827 528619 264830
rect 524321 264618 524387 264621
rect 527265 264618 527331 264621
rect 524321 264616 527331 264618
rect 524321 264560 524326 264616
rect 524382 264560 527270 264616
rect 527326 264560 527331 264616
rect 524321 264558 527331 264560
rect 524321 264555 524387 264558
rect 527265 264555 527331 264558
rect 522113 264482 522179 264485
rect 528645 264482 528711 264485
rect 522113 264480 528711 264482
rect 522113 264424 522118 264480
rect 522174 264424 528650 264480
rect 528706 264424 528711 264480
rect 522113 264422 528711 264424
rect 522113 264419 522179 264422
rect 528645 264419 528711 264422
rect 519629 263666 519695 263669
rect 527817 263666 527883 263669
rect 519629 263664 527883 263666
rect 519629 263608 519634 263664
rect 519690 263608 527822 263664
rect 527878 263608 527883 263664
rect 519629 263606 527883 263608
rect 519629 263603 519695 263606
rect 527817 263603 527883 263606
rect 295149 262850 295215 262853
rect 298185 262850 298251 262853
rect 295149 262848 298251 262850
rect 295149 262792 295154 262848
rect 295210 262792 298190 262848
rect 298246 262792 298251 262848
rect 295149 262790 298251 262792
rect 295149 262787 295215 262790
rect 298185 262787 298251 262790
rect 302146 261998 302462 261999
rect 302146 261934 302152 261998
rect 302216 261934 302232 261998
rect 302296 261934 302312 261998
rect 302376 261934 302392 261998
rect 302456 261934 302462 261998
rect 302146 261918 302462 261934
rect 302146 261854 302152 261918
rect 302216 261854 302232 261918
rect 302296 261854 302312 261918
rect 302376 261854 302392 261918
rect 302456 261854 302462 261918
rect 302146 261838 302462 261854
rect 302146 261774 302152 261838
rect 302216 261774 302232 261838
rect 302296 261774 302312 261838
rect 302376 261774 302392 261838
rect 302456 261774 302462 261838
rect 302146 261758 302462 261774
rect 302146 261694 302152 261758
rect 302216 261694 302232 261758
rect 302296 261694 302312 261758
rect 302376 261694 302392 261758
rect 302456 261694 302462 261758
rect 302146 261693 302462 261694
rect 309146 261998 309462 261999
rect 309146 261934 309152 261998
rect 309216 261934 309232 261998
rect 309296 261934 309312 261998
rect 309376 261934 309392 261998
rect 309456 261934 309462 261998
rect 309146 261918 309462 261934
rect 309146 261854 309152 261918
rect 309216 261854 309232 261918
rect 309296 261854 309312 261918
rect 309376 261854 309392 261918
rect 309456 261854 309462 261918
rect 309146 261838 309462 261854
rect 309146 261774 309152 261838
rect 309216 261774 309232 261838
rect 309296 261774 309312 261838
rect 309376 261774 309392 261838
rect 309456 261774 309462 261838
rect 309146 261758 309462 261774
rect 309146 261694 309152 261758
rect 309216 261694 309232 261758
rect 309296 261694 309312 261758
rect 309376 261694 309392 261758
rect 309456 261694 309462 261758
rect 309146 261693 309462 261694
rect 312813 261626 312879 261629
rect 315757 261626 315823 261629
rect 312813 261624 315823 261626
rect 312813 261568 312818 261624
rect 312874 261568 315762 261624
rect 315818 261568 315823 261624
rect 312813 261566 315823 261568
rect 312813 261563 312879 261566
rect 315757 261563 315823 261566
rect 303878 261237 304194 261238
rect 303878 261173 303884 261237
rect 303948 261173 303964 261237
rect 304028 261173 304044 261237
rect 304108 261173 304124 261237
rect 304188 261173 304194 261237
rect 303878 261157 304194 261173
rect 303878 261093 303884 261157
rect 303948 261093 303964 261157
rect 304028 261093 304044 261157
rect 304108 261093 304124 261157
rect 304188 261093 304194 261157
rect 303878 261077 304194 261093
rect 303878 261013 303884 261077
rect 303948 261013 303964 261077
rect 304028 261013 304044 261077
rect 304108 261013 304124 261077
rect 304188 261013 304194 261077
rect 319437 261082 319503 261085
rect 319437 261080 518052 261082
rect 319437 261024 319442 261080
rect 319498 261024 518052 261080
rect 319437 261022 518052 261024
rect 319437 261019 319503 261022
rect 303878 260997 304194 261013
rect 303878 260933 303884 260997
rect 303948 260933 303964 260997
rect 304028 260933 304044 260997
rect 304108 260933 304124 260997
rect 304188 260933 304194 260997
rect 303878 260917 304194 260933
rect 303878 260853 303884 260917
rect 303948 260853 303964 260917
rect 304028 260853 304044 260917
rect 304108 260853 304124 260917
rect 304188 260853 304194 260917
rect 303878 260837 304194 260853
rect 303878 260773 303884 260837
rect 303948 260773 303964 260837
rect 304028 260773 304044 260837
rect 304108 260773 304124 260837
rect 304188 260773 304194 260837
rect 303878 260757 304194 260773
rect 303878 260693 303884 260757
rect 303948 260693 303964 260757
rect 304028 260693 304044 260757
rect 304108 260693 304124 260757
rect 304188 260693 304194 260757
rect 303878 260677 304194 260693
rect 303878 260613 303884 260677
rect 303948 260613 303964 260677
rect 304028 260613 304044 260677
rect 304108 260613 304124 260677
rect 304188 260613 304194 260677
rect 309501 260674 309567 260677
rect 309396 260672 309567 260674
rect 309396 260616 309506 260672
rect 309562 260616 309567 260672
rect 309396 260614 309567 260616
rect 303878 260612 304194 260613
rect 309501 260611 309567 260614
rect 305913 260538 305979 260541
rect 318425 260538 318491 260541
rect 305913 260536 318491 260538
rect 305913 260480 305918 260536
rect 305974 260480 318430 260536
rect 318486 260480 318491 260536
rect 305913 260478 318491 260480
rect 305913 260475 305979 260478
rect 318425 260475 318491 260478
rect 318057 259722 318123 259725
rect 318057 259720 518052 259722
rect 318057 259664 318062 259720
rect 318118 259664 518052 259720
rect 318057 259662 518052 259664
rect 318057 259659 318123 259662
rect 309501 259450 309567 259453
rect 515581 259450 515647 259453
rect 309501 259448 515647 259450
rect 309501 259392 309506 259448
rect 309562 259392 515586 259448
rect 515642 259392 515647 259448
rect 309501 259390 515647 259392
rect 309501 259387 309567 259390
rect 515581 259387 515647 259390
rect 299013 259314 299079 259317
rect 315665 259314 315731 259317
rect 299013 259312 315731 259314
rect 299013 259256 299018 259312
rect 299074 259256 315670 259312
rect 315726 259256 315731 259312
rect 299013 259254 315731 259256
rect 299013 259251 299079 259254
rect 315665 259251 315731 259254
rect 302601 259178 302667 259181
rect 314009 259178 314075 259181
rect 302601 259176 314075 259178
rect 302601 259120 302606 259176
rect 302662 259120 314014 259176
rect 314070 259120 314075 259176
rect 302601 259118 314075 259120
rect 302601 259115 302667 259118
rect 314009 259115 314075 259118
rect 583520 258756 584960 258996
rect 315297 258362 315363 258365
rect 315297 258360 518052 258362
rect 315297 258304 315302 258360
rect 315358 258304 518052 258360
rect 315297 258302 518052 258304
rect 315297 258299 315363 258302
rect 315481 257002 315547 257005
rect 315481 257000 518052 257002
rect 315481 256944 315486 257000
rect 315542 256944 518052 257000
rect 315481 256942 518052 256944
rect 315481 256939 315547 256942
rect 315573 255642 315639 255645
rect 315573 255640 518052 255642
rect 315573 255584 315578 255640
rect 315634 255584 518052 255640
rect 315573 255582 518052 255584
rect 315573 255579 315639 255582
rect 384297 254282 384363 254285
rect 384297 254280 518052 254282
rect -960 253996 480 254236
rect 384297 254224 384302 254280
rect 384358 254224 518052 254280
rect 384297 254222 518052 254224
rect 384297 254219 384363 254222
rect 381537 252922 381603 252925
rect 381537 252920 518052 252922
rect 381537 252864 381542 252920
rect 381598 252864 518052 252920
rect 381537 252862 518052 252864
rect 381537 252859 381603 252862
rect 314101 251562 314167 251565
rect 314101 251560 518052 251562
rect 314101 251504 314106 251560
rect 314162 251504 518052 251560
rect 314101 251502 518052 251504
rect 314101 251499 314167 251502
rect 529933 251018 529999 251021
rect 530577 251018 530643 251021
rect 527804 251016 530643 251018
rect 527804 250960 529938 251016
rect 529994 250960 530582 251016
rect 530638 250960 530643 251016
rect 527804 250958 530643 250960
rect 529933 250955 529999 250958
rect 530577 250955 530643 250958
rect 314193 250202 314259 250205
rect 314193 250200 518052 250202
rect 314193 250144 314198 250200
rect 314254 250144 518052 250200
rect 314193 250142 518052 250144
rect 314193 250139 314259 250142
rect 317137 248842 317203 248845
rect 317137 248840 518052 248842
rect 317137 248784 317142 248840
rect 317198 248784 518052 248840
rect 317137 248782 518052 248784
rect 317137 248779 317203 248782
rect 382917 247482 382983 247485
rect 382917 247480 518052 247482
rect 382917 247424 382922 247480
rect 382978 247424 518052 247480
rect 382917 247422 518052 247424
rect 382917 247419 382983 247422
rect 315757 246122 315823 246125
rect 315757 246120 518052 246122
rect 315757 246064 315762 246120
rect 315818 246064 518052 246120
rect 315757 246062 518052 246064
rect 315757 246059 315823 246062
rect 527817 245578 527883 245581
rect 583520 245578 584960 245668
rect 527817 245576 584960 245578
rect 527817 245520 527822 245576
rect 527878 245520 584960 245576
rect 527817 245518 584960 245520
rect 527817 245515 527883 245518
rect 583520 245428 584960 245518
rect 514753 244762 514819 244765
rect 514753 244760 518052 244762
rect 514753 244704 514758 244760
rect 514814 244704 518052 244760
rect 514753 244702 518052 244704
rect 514753 244699 514819 244702
rect 295241 243538 295307 243541
rect 300853 243538 300919 243541
rect 295241 243536 300919 243538
rect 295241 243480 295246 243536
rect 295302 243480 300858 243536
rect 300914 243480 300919 243536
rect 295241 243478 300919 243480
rect 295241 243475 295307 243478
rect 300853 243475 300919 243478
rect 304625 243402 304691 243405
rect 312077 243402 312143 243405
rect 312905 243402 312971 243405
rect 304625 243400 312971 243402
rect 304625 243344 304630 243400
rect 304686 243344 312082 243400
rect 312138 243344 312910 243400
rect 312966 243344 312971 243400
rect 304625 243342 312971 243344
rect 304625 243339 304691 243342
rect 312077 243339 312143 243342
rect 312905 243339 312971 243342
rect 515673 243402 515739 243405
rect 515673 243400 518052 243402
rect 515673 243344 515678 243400
rect 515734 243344 518052 243400
rect 515673 243342 518052 243344
rect 515673 243339 515739 243342
rect 296878 242084 297194 242085
rect 296878 242020 296884 242084
rect 296948 242020 296964 242084
rect 297028 242020 297044 242084
rect 297108 242020 297124 242084
rect 297188 242020 297194 242084
rect 296878 242004 297194 242020
rect 296878 241940 296884 242004
rect 296948 241940 296964 242004
rect 297028 241940 297044 242004
rect 297108 241940 297124 242004
rect 297188 241940 297194 242004
rect 296878 241924 297194 241940
rect 296878 241860 296884 241924
rect 296948 241860 296964 241924
rect 297028 241860 297044 241924
rect 297108 241860 297124 241924
rect 297188 241860 297194 241924
rect 303878 242084 304194 242085
rect 303878 242020 303884 242084
rect 303948 242020 303964 242084
rect 304028 242020 304044 242084
rect 304108 242020 304124 242084
rect 304188 242020 304194 242084
rect 303878 242004 304194 242020
rect 303878 241940 303884 242004
rect 303948 241940 303964 242004
rect 304028 241940 304044 242004
rect 304108 241940 304124 242004
rect 304188 241940 304194 242004
rect 303878 241924 304194 241940
rect 296878 241844 297194 241860
rect 296878 241780 296884 241844
rect 296948 241780 296964 241844
rect 297028 241780 297044 241844
rect 297108 241780 297124 241844
rect 297188 241780 297194 241844
rect 300853 241906 300919 241909
rect 300853 241904 300962 241906
rect 300853 241848 300858 241904
rect 300914 241848 300962 241904
rect 300853 241843 300962 241848
rect 296878 241779 297194 241780
rect 300902 241637 300962 241843
rect 303878 241860 303884 241924
rect 303948 241860 303964 241924
rect 304028 241860 304044 241924
rect 304108 241860 304124 241924
rect 304188 241860 304194 241924
rect 310878 242084 311194 242085
rect 310878 242020 310884 242084
rect 310948 242020 310964 242084
rect 311028 242020 311044 242084
rect 311108 242020 311124 242084
rect 311188 242020 311194 242084
rect 310878 242004 311194 242020
rect 310878 241940 310884 242004
rect 310948 241940 310964 242004
rect 311028 241940 311044 242004
rect 311108 241940 311124 242004
rect 311188 241940 311194 242004
rect 515581 242042 515647 242045
rect 515581 242040 518052 242042
rect 515581 241984 515586 242040
rect 515642 241984 518052 242040
rect 515581 241982 518052 241984
rect 515581 241979 515647 241982
rect 310878 241924 311194 241940
rect 304625 241906 304691 241909
rect 303878 241844 304194 241860
rect 303878 241780 303884 241844
rect 303948 241780 303964 241844
rect 304028 241780 304044 241844
rect 304108 241780 304124 241844
rect 304188 241780 304194 241844
rect 303878 241779 304194 241780
rect 304582 241904 304691 241906
rect 304582 241848 304630 241904
rect 304686 241848 304691 241904
rect 304582 241843 304691 241848
rect 310878 241860 310884 241924
rect 310948 241860 310964 241924
rect 311028 241860 311044 241924
rect 311108 241860 311124 241924
rect 311188 241860 311194 241924
rect 310878 241844 311194 241860
rect 300902 241632 301011 241637
rect 300902 241576 300950 241632
rect 301006 241576 301011 241632
rect 300902 241574 301011 241576
rect 300945 241571 301011 241574
rect 304582 241501 304642 241843
rect 310878 241780 310884 241844
rect 310948 241780 310964 241844
rect 311028 241780 311044 241844
rect 311108 241780 311124 241844
rect 311188 241780 311194 241844
rect 310878 241779 311194 241780
rect 304543 241496 304642 241501
rect 304543 241440 304548 241496
rect 304604 241440 304642 241496
rect 304543 241438 304642 241440
rect 304543 241435 304609 241438
rect -960 240940 480 241180
rect 295146 240999 295462 241000
rect 295146 240935 295152 240999
rect 295216 240935 295232 240999
rect 295296 240935 295312 240999
rect 295376 240935 295392 240999
rect 295456 240935 295462 240999
rect 295146 240919 295462 240935
rect 295146 240855 295152 240919
rect 295216 240855 295232 240919
rect 295296 240855 295312 240919
rect 295376 240855 295392 240919
rect 295456 240855 295462 240919
rect 295146 240839 295462 240855
rect 295146 240775 295152 240839
rect 295216 240775 295232 240839
rect 295296 240775 295312 240839
rect 295376 240775 295392 240839
rect 295456 240775 295462 240839
rect 295146 240759 295462 240775
rect 295146 240695 295152 240759
rect 295216 240695 295232 240759
rect 295296 240695 295312 240759
rect 295376 240695 295392 240759
rect 295456 240695 295462 240759
rect 295146 240694 295462 240695
rect 309146 240973 309462 240974
rect 309146 240909 309152 240973
rect 309216 240909 309232 240973
rect 309296 240909 309312 240973
rect 309376 240909 309392 240973
rect 309456 240909 309462 240973
rect 309146 240893 309462 240909
rect 309146 240829 309152 240893
rect 309216 240829 309232 240893
rect 309296 240829 309312 240893
rect 309376 240829 309392 240893
rect 309456 240829 309462 240893
rect 309146 240813 309462 240829
rect 309146 240749 309152 240813
rect 309216 240749 309232 240813
rect 309296 240749 309312 240813
rect 309376 240749 309392 240813
rect 309456 240749 309462 240813
rect 309146 240733 309462 240749
rect 309146 240669 309152 240733
rect 309216 240669 309232 240733
rect 309296 240669 309312 240733
rect 309376 240669 309392 240733
rect 309456 240669 309462 240733
rect 309146 240668 309462 240669
rect 402237 240682 402303 240685
rect 402237 240680 518052 240682
rect 402237 240624 402242 240680
rect 402298 240624 518052 240680
rect 402237 240622 518052 240624
rect 402237 240619 402303 240622
rect 310878 239912 311194 239913
rect 310878 239848 310884 239912
rect 310948 239848 310964 239912
rect 311028 239848 311044 239912
rect 311108 239848 311124 239912
rect 311188 239848 311194 239912
rect 310878 239832 311194 239848
rect 310878 239768 310884 239832
rect 310948 239768 310964 239832
rect 311028 239768 311044 239832
rect 311108 239768 311124 239832
rect 311188 239768 311194 239832
rect 310878 239752 311194 239768
rect 310878 239688 310884 239752
rect 310948 239688 310964 239752
rect 311028 239688 311044 239752
rect 311108 239688 311124 239752
rect 311188 239688 311194 239752
rect 310878 239672 311194 239688
rect 310878 239608 310884 239672
rect 310948 239608 310964 239672
rect 311028 239608 311044 239672
rect 311108 239608 311124 239672
rect 311188 239608 311194 239672
rect 310878 239607 311194 239608
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 309869 222730 309935 222733
rect 312537 222730 312603 222733
rect 309869 222728 312603 222730
rect 309869 222672 309874 222728
rect 309930 222672 312542 222728
rect 312598 222672 312603 222728
rect 309869 222670 312603 222672
rect 309869 222667 309935 222670
rect 312537 222667 312603 222670
rect 294873 222458 294939 222461
rect 305729 222458 305795 222461
rect 294873 222456 306390 222458
rect 294873 222400 294878 222456
rect 294934 222400 305734 222456
rect 305790 222400 306390 222456
rect 294873 222398 306390 222400
rect 294873 222395 294939 222398
rect 305729 222395 305795 222398
rect 306330 222322 306390 222398
rect 312077 222322 312143 222325
rect 306330 222320 312143 222322
rect 306330 222264 312082 222320
rect 312138 222264 312143 222320
rect 306330 222262 312143 222264
rect 312077 222259 312143 222262
rect 295057 221234 295123 221237
rect 295057 221232 300042 221234
rect 295057 221176 295062 221232
rect 295118 221176 300042 221232
rect 295057 221174 300042 221176
rect 295057 221171 295123 221174
rect 296878 221085 297194 221086
rect 296878 221021 296884 221085
rect 296948 221021 296964 221085
rect 297028 221021 297044 221085
rect 297108 221021 297124 221085
rect 297188 221021 297194 221085
rect 296878 221005 297194 221021
rect 296878 220941 296884 221005
rect 296948 220941 296964 221005
rect 297028 220941 297044 221005
rect 297108 220941 297124 221005
rect 297188 220941 297194 221005
rect 296878 220925 297194 220941
rect 296878 220861 296884 220925
rect 296948 220861 296964 220925
rect 297028 220861 297044 220925
rect 297108 220861 297124 220925
rect 297188 220861 297194 220925
rect 299982 220962 300042 221174
rect 303878 221085 304194 221086
rect 303878 221021 303884 221085
rect 303948 221021 303964 221085
rect 304028 221021 304044 221085
rect 304108 221021 304124 221085
rect 304188 221021 304194 221085
rect 303878 221005 304194 221021
rect 301313 220962 301379 220965
rect 299982 220960 301882 220962
rect 299982 220904 301318 220960
rect 301374 220904 301882 220960
rect 299982 220902 301882 220904
rect 301313 220899 301379 220902
rect 296878 220845 297194 220861
rect 296878 220781 296884 220845
rect 296948 220781 296964 220845
rect 297028 220781 297044 220845
rect 297108 220781 297124 220845
rect 297188 220781 297194 220845
rect 296878 220780 297194 220781
rect 301822 220693 301882 220902
rect 303878 220941 303884 221005
rect 303948 220941 303964 221005
rect 304028 220941 304044 221005
rect 304108 220941 304124 221005
rect 304188 220941 304194 221005
rect 310878 221085 311194 221086
rect 310878 221021 310884 221085
rect 310948 221021 310964 221085
rect 311028 221021 311044 221085
rect 311108 221021 311124 221085
rect 311188 221021 311194 221085
rect 310878 221005 311194 221021
rect 305729 220962 305795 220965
rect 309869 220962 309935 220965
rect 303878 220925 304194 220941
rect 303878 220861 303884 220925
rect 303948 220861 303964 220925
rect 304028 220861 304044 220925
rect 304108 220861 304124 220925
rect 304188 220861 304194 220925
rect 303878 220845 304194 220861
rect 303878 220781 303884 220845
rect 303948 220781 303964 220845
rect 304028 220781 304044 220845
rect 304108 220781 304124 220845
rect 304188 220781 304194 220845
rect 303878 220780 304194 220781
rect 305686 220960 305795 220962
rect 305686 220904 305734 220960
rect 305790 220904 305795 220960
rect 305686 220899 305795 220904
rect 309734 220960 309935 220962
rect 309734 220904 309874 220960
rect 309930 220904 309935 220960
rect 309734 220902 309935 220904
rect 305686 220693 305746 220899
rect 309734 220693 309794 220902
rect 309869 220899 309935 220902
rect 310878 220941 310884 221005
rect 310948 220941 310964 221005
rect 311028 220941 311044 221005
rect 311108 220941 311124 221005
rect 311188 220941 311194 221005
rect 310878 220925 311194 220941
rect 310878 220861 310884 220925
rect 310948 220861 310964 220925
rect 311028 220861 311044 220925
rect 311108 220861 311124 220925
rect 311188 220861 311194 220925
rect 310878 220845 311194 220861
rect 310878 220781 310884 220845
rect 310948 220781 310964 220845
rect 311028 220781 311044 220845
rect 311108 220781 311124 220845
rect 311188 220781 311194 220845
rect 310878 220780 311194 220781
rect 301822 220688 301931 220693
rect 301822 220632 301870 220688
rect 301926 220632 301931 220688
rect 301822 220630 301931 220632
rect 305686 220688 305795 220693
rect 305686 220632 305734 220688
rect 305790 220632 305795 220688
rect 305686 220630 305795 220632
rect 301865 220627 301931 220630
rect 305729 220627 305795 220630
rect 309685 220688 309794 220693
rect 309685 220632 309690 220688
rect 309746 220632 309794 220688
rect 309685 220630 309794 220632
rect 309685 220627 309751 220630
rect 295146 220000 295462 220001
rect 295146 219936 295152 220000
rect 295216 219936 295232 220000
rect 295296 219936 295312 220000
rect 295376 219936 295392 220000
rect 295456 219936 295462 220000
rect 295146 219920 295462 219936
rect 295146 219856 295152 219920
rect 295216 219856 295232 219920
rect 295296 219856 295312 219920
rect 295376 219856 295392 219920
rect 295456 219856 295462 219920
rect 295146 219840 295462 219856
rect 295146 219776 295152 219840
rect 295216 219776 295232 219840
rect 295296 219776 295312 219840
rect 295376 219776 295392 219840
rect 295456 219776 295462 219840
rect 295146 219760 295462 219776
rect 295146 219696 295152 219760
rect 295216 219696 295232 219760
rect 295296 219696 295312 219760
rect 295376 219696 295392 219760
rect 295456 219696 295462 219760
rect 295146 219695 295462 219696
rect 302146 219999 302462 220000
rect 302146 219935 302152 219999
rect 302216 219935 302232 219999
rect 302296 219935 302312 219999
rect 302376 219935 302392 219999
rect 302456 219935 302462 219999
rect 302146 219919 302462 219935
rect 302146 219855 302152 219919
rect 302216 219855 302232 219919
rect 302296 219855 302312 219919
rect 302376 219855 302392 219919
rect 302456 219855 302462 219919
rect 302146 219839 302462 219855
rect 302146 219775 302152 219839
rect 302216 219775 302232 219839
rect 302296 219775 302312 219839
rect 302376 219775 302392 219839
rect 302456 219775 302462 219839
rect 302146 219759 302462 219775
rect 302146 219695 302152 219759
rect 302216 219695 302232 219759
rect 302296 219695 302312 219759
rect 302376 219695 302392 219759
rect 302456 219695 302462 219759
rect 302146 219694 302462 219695
rect 309146 219999 309462 220000
rect 309146 219935 309152 219999
rect 309216 219935 309232 219999
rect 309296 219935 309312 219999
rect 309376 219935 309392 219999
rect 309456 219935 309462 219999
rect 309146 219919 309462 219935
rect 309146 219855 309152 219919
rect 309216 219855 309232 219919
rect 309296 219855 309312 219919
rect 309376 219855 309392 219919
rect 309456 219855 309462 219919
rect 309146 219839 309462 219855
rect 309146 219775 309152 219839
rect 309216 219775 309232 219839
rect 309296 219775 309312 219839
rect 309376 219775 309392 219839
rect 309456 219775 309462 219839
rect 309146 219759 309462 219775
rect 309146 219695 309152 219759
rect 309216 219695 309232 219759
rect 309296 219695 309312 219759
rect 309376 219695 309392 219759
rect 309456 219695 309462 219759
rect 309146 219694 309462 219695
rect 310998 219519 311144 219520
rect 310998 219455 311039 219519
rect 311103 219455 311144 219519
rect 310998 219454 311144 219455
rect 303918 219402 304064 219403
rect 303918 219338 303959 219402
rect 304023 219338 304064 219402
rect 303918 219337 304064 219338
rect 583520 218908 584960 219148
rect 314180 218726 321570 218786
rect 321510 218650 321570 218726
rect 515673 218650 515739 218653
rect 321510 218648 515739 218650
rect 321510 218592 515678 218648
rect 515734 218592 515739 218648
rect 321510 218590 515739 218592
rect 515673 218587 515739 218590
rect 307661 217970 307727 217973
rect 309593 217970 309659 217973
rect 315389 217970 315455 217973
rect 307661 217968 309659 217970
rect 307661 217912 307666 217968
rect 307722 217912 309598 217968
rect 309654 217912 309659 217968
rect 307661 217910 309659 217912
rect 307661 217907 307727 217910
rect 309593 217907 309659 217910
rect 310286 217968 315455 217970
rect 310286 217912 315394 217968
rect 315450 217912 315455 217968
rect 310286 217910 315455 217912
rect 299289 217834 299355 217837
rect 310286 217834 310346 217910
rect 315389 217907 315455 217910
rect 299289 217832 310346 217834
rect 299289 217776 299294 217832
rect 299350 217776 310346 217832
rect 299289 217774 310346 217776
rect 310421 217834 310487 217837
rect 317045 217834 317111 217837
rect 310421 217832 317111 217834
rect 310421 217776 310426 217832
rect 310482 217776 317050 217832
rect 317106 217776 317111 217832
rect 310421 217774 317111 217776
rect 299289 217771 299355 217774
rect 310421 217771 310487 217774
rect 317045 217771 317111 217774
rect 303153 217562 303219 217565
rect 347037 217562 347103 217565
rect 303153 217560 347103 217562
rect 303153 217504 303158 217560
rect 303214 217504 347042 217560
rect 347098 217504 347103 217560
rect 303153 217502 347103 217504
rect 303153 217499 303219 217502
rect 347037 217499 347103 217502
rect 306741 217426 306807 217429
rect 318333 217426 318399 217429
rect 306741 217424 318399 217426
rect 306741 217368 306746 217424
rect 306802 217368 318338 217424
rect 318394 217368 318399 217424
rect 306741 217366 318399 217368
rect 306741 217363 306807 217366
rect 318333 217363 318399 217366
rect 310421 216746 310487 216749
rect 313917 216746 313983 216749
rect 310421 216744 313983 216746
rect 310421 216688 310426 216744
rect 310482 216688 313922 216744
rect 313978 216688 313983 216744
rect 310421 216686 313983 216688
rect 310421 216683 310487 216686
rect 313917 216683 313983 216686
rect -960 214828 480 215068
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 294965 202874 295031 202877
rect 295241 202874 295307 202877
rect 294965 202872 295307 202874
rect 294965 202816 294970 202872
rect 295026 202816 295246 202872
rect 295302 202816 295307 202872
rect 294965 202814 295307 202816
rect 294965 202811 295031 202814
rect 295241 202811 295307 202814
rect 294873 202194 294939 202197
rect 303613 202194 303679 202197
rect 294873 202192 303679 202194
rect 294873 202136 294878 202192
rect 294934 202136 303618 202192
rect 303674 202136 303679 202192
rect 294873 202134 303679 202136
rect 294873 202131 294939 202134
rect 303613 202131 303679 202134
rect -960 201772 480 202012
rect 295057 201514 295123 201517
rect 300853 201514 300919 201517
rect 295057 201512 300919 201514
rect 295057 201456 295062 201512
rect 295118 201456 300858 201512
rect 300914 201456 300919 201512
rect 295057 201454 300919 201456
rect 295057 201451 295123 201454
rect 300853 201451 300919 201454
rect 303613 201514 303679 201517
rect 311157 201514 311223 201517
rect 303613 201512 311223 201514
rect 303613 201456 303618 201512
rect 303674 201456 311162 201512
rect 311218 201456 311223 201512
rect 303613 201454 311223 201456
rect 303613 201451 303679 201454
rect 311157 201451 311223 201454
rect 307661 200290 307727 200293
rect 307158 200288 307727 200290
rect 307158 200232 307666 200288
rect 307722 200232 307727 200288
rect 307158 200230 307727 200232
rect 300853 199882 300919 199885
rect 303613 199882 303679 199885
rect 300853 199880 300962 199882
rect 300853 199824 300858 199880
rect 300914 199824 300962 199880
rect 300853 199819 300962 199824
rect 303613 199880 303722 199882
rect 303613 199824 303618 199880
rect 303674 199824 303722 199880
rect 303613 199819 303722 199824
rect 300902 199613 300962 199819
rect 300853 199608 300962 199613
rect 300853 199552 300858 199608
rect 300914 199552 300962 199608
rect 300853 199550 300962 199552
rect 303662 199613 303722 199819
rect 303662 199608 303771 199613
rect 303662 199552 303710 199608
rect 303766 199552 303771 199608
rect 303662 199550 303771 199552
rect 307158 199610 307218 200230
rect 307661 200227 307727 200230
rect 307569 199610 307635 199613
rect 307158 199608 307635 199610
rect 307158 199552 307574 199608
rect 307630 199552 307635 199608
rect 307158 199550 307635 199552
rect 300853 199547 300919 199550
rect 303705 199547 303771 199550
rect 307569 199547 307635 199550
rect 515581 197706 515647 197709
rect 310868 197704 515647 197706
rect 310868 197648 515586 197704
rect 515642 197648 515647 197704
rect 310868 197646 515647 197648
rect 515581 197643 515647 197646
rect 304717 197298 304783 197301
rect 371877 197298 371943 197301
rect 304717 197296 371943 197298
rect 304717 197240 304722 197296
rect 304778 197240 371882 197296
rect 371938 197240 371943 197296
rect 304717 197238 371943 197240
rect 304717 197235 304783 197238
rect 371877 197235 371943 197238
rect 301681 197162 301747 197165
rect 316953 197162 317019 197165
rect 301681 197160 317019 197162
rect 301681 197104 301686 197160
rect 301742 197104 316958 197160
rect 317014 197104 317019 197160
rect 301681 197102 317019 197104
rect 301681 197099 301747 197102
rect 316953 197099 317019 197102
rect 307753 195938 307819 195941
rect 515489 195938 515555 195941
rect 307753 195936 515555 195938
rect 307753 195880 307758 195936
rect 307814 195880 515494 195936
rect 515550 195880 515555 195936
rect 307753 195878 515555 195880
rect 307753 195875 307819 195878
rect 515489 195875 515555 195878
rect 298645 195802 298711 195805
rect 316769 195802 316835 195805
rect 298645 195800 316835 195802
rect 298645 195744 298650 195800
rect 298706 195744 316774 195800
rect 316830 195744 316835 195800
rect 298645 195742 316835 195744
rect 298645 195739 298711 195742
rect 316769 195739 316835 195742
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 295057 181386 295123 181389
rect 304441 181386 304507 181389
rect 311157 181386 311223 181389
rect 371877 181386 371943 181389
rect 295057 181384 296730 181386
rect 295057 181328 295062 181384
rect 295118 181328 296730 181384
rect 295057 181326 296730 181328
rect 295057 181323 295123 181326
rect 296670 181114 296730 181326
rect 304441 181384 371943 181386
rect 304441 181328 304446 181384
rect 304502 181328 311162 181384
rect 311218 181328 371882 181384
rect 371938 181328 371943 181384
rect 304441 181326 371943 181328
rect 304441 181323 304507 181326
rect 311157 181323 311223 181326
rect 371877 181323 371943 181326
rect 300853 181114 300919 181117
rect 342897 181114 342963 181117
rect 296670 181112 342963 181114
rect 296670 181056 300858 181112
rect 300914 181056 342902 181112
rect 342958 181056 342963 181112
rect 296670 181054 342963 181056
rect 300853 181051 300919 181054
rect 342897 181051 342963 181054
rect 297265 180978 297331 180981
rect 311157 180978 311223 180981
rect 296670 180976 311223 180978
rect 296670 180920 297270 180976
rect 297326 180920 311162 180976
rect 311218 180920 311223 180976
rect 296670 180918 311223 180920
rect 295241 180842 295307 180845
rect 296670 180842 296730 180918
rect 297265 180915 297331 180918
rect 311157 180915 311223 180918
rect 295241 180840 296730 180842
rect 295241 180784 295246 180840
rect 295302 180784 296730 180840
rect 295241 180782 296730 180784
rect 295241 180779 295307 180782
rect 307661 179482 307727 179485
rect 580257 179482 580323 179485
rect 307158 179480 580323 179482
rect 307158 179424 307666 179480
rect 307722 179424 580262 179480
rect 580318 179424 580323 179480
rect 307158 179422 580323 179424
rect 296878 179285 297194 179286
rect 296878 179221 296884 179285
rect 296948 179221 296964 179285
rect 297028 179221 297044 179285
rect 297108 179221 297124 179285
rect 297188 179221 297194 179285
rect 296878 179205 297194 179221
rect 296878 179141 296884 179205
rect 296948 179141 296964 179205
rect 297028 179141 297044 179205
rect 297108 179141 297124 179205
rect 297188 179141 297194 179205
rect 296878 179125 297194 179141
rect 296878 179061 296884 179125
rect 296948 179061 296964 179125
rect 297028 179061 297044 179125
rect 297108 179061 297124 179125
rect 297188 179061 297194 179125
rect 303878 179285 304194 179286
rect 303878 179221 303884 179285
rect 303948 179221 303964 179285
rect 304028 179221 304044 179285
rect 304108 179221 304124 179285
rect 304188 179221 304194 179285
rect 303878 179205 304194 179221
rect 303878 179141 303884 179205
rect 303948 179141 303964 179205
rect 304028 179141 304044 179205
rect 304108 179141 304124 179205
rect 304188 179141 304194 179205
rect 303878 179125 304194 179141
rect 296878 179045 297194 179061
rect 296878 178981 296884 179045
rect 296948 178981 296964 179045
rect 297028 178981 297044 179045
rect 297108 178981 297124 179045
rect 297188 178981 297194 179045
rect 297265 179072 297331 179077
rect 297265 179016 297270 179072
rect 297326 179016 297331 179072
rect 297265 179011 297331 179016
rect 300853 179074 300919 179077
rect 300853 179072 300962 179074
rect 300853 179016 300858 179072
rect 300914 179016 300962 179072
rect 300853 179011 300962 179016
rect 296878 178980 297194 178981
rect 297268 178805 297328 179011
rect 300902 178805 300962 179011
rect 303878 179061 303884 179125
rect 303948 179061 303964 179125
rect 304028 179061 304044 179125
rect 304108 179061 304124 179125
rect 304188 179061 304194 179125
rect 304441 179074 304507 179077
rect 303878 179045 304194 179061
rect 303878 178981 303884 179045
rect 303948 178981 303964 179045
rect 304028 178981 304044 179045
rect 304108 178981 304124 179045
rect 304188 178981 304194 179045
rect 303878 178980 304194 178981
rect 304398 179072 304507 179074
rect 304398 179016 304446 179072
rect 304502 179016 304507 179072
rect 304398 179011 304507 179016
rect 297265 178800 297331 178805
rect 297265 178744 297270 178800
rect 297326 178744 297331 178800
rect 297265 178739 297331 178744
rect 300852 178800 300962 178805
rect 300852 178744 300857 178800
rect 300913 178744 300962 178800
rect 300852 178742 300962 178744
rect 303904 178802 303970 178805
rect 304398 178802 304458 179011
rect 307158 178805 307218 179422
rect 307661 179419 307727 179422
rect 580257 179419 580323 179422
rect 310882 179285 310958 179286
rect 310882 179221 310888 179285
rect 310952 179221 310958 179285
rect 310882 179205 310958 179221
rect 310882 179141 310888 179205
rect 310952 179141 310958 179205
rect 310882 179125 310958 179141
rect 310882 179061 310888 179125
rect 310952 179061 310958 179125
rect 310882 179045 310958 179061
rect 583520 179060 584960 179300
rect 310882 178981 310888 179045
rect 310952 178981 310958 179045
rect 310882 178980 310958 178981
rect 303904 178800 304458 178802
rect 303904 178744 303909 178800
rect 303965 178744 304458 178800
rect 303904 178742 304458 178744
rect 307109 178800 307218 178805
rect 307109 178744 307114 178800
rect 307170 178744 307218 178800
rect 307109 178742 307218 178744
rect 300852 178739 300918 178742
rect 303904 178739 303970 178742
rect 307109 178739 307175 178742
rect 295146 178199 295462 178200
rect 295146 178135 295152 178199
rect 295216 178135 295232 178199
rect 295296 178135 295312 178199
rect 295376 178135 295392 178199
rect 295456 178135 295462 178199
rect 295146 178119 295462 178135
rect 295146 178055 295152 178119
rect 295216 178055 295232 178119
rect 295296 178055 295312 178119
rect 295376 178055 295392 178119
rect 295456 178055 295462 178119
rect 295146 178039 295462 178055
rect 295146 177975 295152 178039
rect 295216 177975 295232 178039
rect 295296 177975 295312 178039
rect 295376 177975 295392 178039
rect 295456 177975 295462 178039
rect 295146 177959 295462 177975
rect 295146 177895 295152 177959
rect 295216 177895 295232 177959
rect 295296 177895 295312 177959
rect 295376 177895 295392 177959
rect 295456 177895 295462 177959
rect 295146 177894 295462 177895
rect 302146 178183 302462 178184
rect 302146 178119 302152 178183
rect 302216 178119 302232 178183
rect 302296 178119 302312 178183
rect 302376 178119 302392 178183
rect 302456 178119 302462 178183
rect 302146 178103 302462 178119
rect 302146 178039 302152 178103
rect 302216 178039 302232 178103
rect 302296 178039 302312 178103
rect 302376 178039 302392 178103
rect 302456 178039 302462 178103
rect 302146 178023 302462 178039
rect 302146 177959 302152 178023
rect 302216 177959 302232 178023
rect 302296 177959 302312 178023
rect 302376 177959 302392 178023
rect 302456 177959 302462 178023
rect 302146 177943 302462 177959
rect 302146 177879 302152 177943
rect 302216 177879 302232 177943
rect 302296 177879 302312 177943
rect 302376 177879 302392 177943
rect 302456 177879 302462 177943
rect 302146 177878 302462 177879
rect 309146 178183 309462 178184
rect 309146 178119 309152 178183
rect 309216 178119 309232 178183
rect 309296 178119 309312 178183
rect 309376 178119 309392 178183
rect 309456 178119 309462 178183
rect 309146 178103 309462 178119
rect 309146 178039 309152 178103
rect 309216 178039 309232 178103
rect 309296 178039 309312 178103
rect 309376 178039 309392 178103
rect 309456 178039 309462 178103
rect 309146 178023 309462 178039
rect 309146 177959 309152 178023
rect 309216 177959 309232 178023
rect 309296 177959 309312 178023
rect 309376 177959 309392 178023
rect 309456 177959 309462 178023
rect 309146 177943 309462 177959
rect 309146 177879 309152 177943
rect 309216 177879 309232 177943
rect 309296 177879 309312 177943
rect 309376 177879 309392 177943
rect 309456 177879 309462 177943
rect 309146 177878 309462 177879
rect 311525 177306 311591 177309
rect 580349 177306 580415 177309
rect 311525 177304 580415 177306
rect 311525 177248 311530 177304
rect 311586 177248 580354 177304
rect 580410 177248 580415 177304
rect 311525 177246 580415 177248
rect 311525 177243 311591 177246
rect 580349 177243 580415 177246
rect 402237 176898 402303 176901
rect 310868 176896 402303 176898
rect 310868 176840 402242 176896
rect 402298 176840 402303 176896
rect 310868 176838 402303 176840
rect 402237 176835 402303 176838
rect 307753 176626 307819 176629
rect 515397 176626 515463 176629
rect 307753 176624 515463 176626
rect 307753 176568 307758 176624
rect 307814 176568 515402 176624
rect 515458 176568 515463 176624
rect 307753 176566 515463 176568
rect 307753 176563 307819 176566
rect 515397 176563 515463 176566
rect 301681 176490 301747 176493
rect 318149 176490 318215 176493
rect 301681 176488 318215 176490
rect 301681 176432 301686 176488
rect 301742 176432 318154 176488
rect 318210 176432 318215 176488
rect 301681 176430 318215 176432
rect 301681 176427 301747 176430
rect 318149 176427 318215 176430
rect -960 175796 480 176036
rect 304717 175266 304783 175269
rect 329097 175266 329163 175269
rect 304717 175264 329163 175266
rect 304717 175208 304722 175264
rect 304778 175208 329102 175264
rect 329158 175208 329163 175264
rect 304717 175206 329163 175208
rect 304717 175203 304783 175206
rect 329097 175203 329163 175206
rect 298645 175130 298711 175133
rect 316677 175130 316743 175133
rect 298645 175128 316743 175130
rect 298645 175072 298650 175128
rect 298706 175072 316682 175128
rect 316738 175072 316743 175128
rect 298645 175070 316743 175072
rect 298645 175067 298711 175070
rect 316677 175067 316743 175070
rect 580349 165882 580415 165885
rect 583520 165882 584960 165972
rect 580349 165880 584960 165882
rect 580349 165824 580354 165880
rect 580410 165824 584960 165880
rect 580349 165822 584960 165824
rect 580349 165819 580415 165822
rect 583520 165732 584960 165822
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 580257 126034 580323 126037
rect 583520 126034 584960 126124
rect 580257 126032 584960 126034
rect 580257 125976 580262 126032
rect 580318 125976 584960 126032
rect 580257 125974 584960 125976
rect 580257 125971 580323 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 371877 86186 371943 86189
rect 583520 86186 584960 86276
rect 371877 86184 584960 86186
rect 371877 86128 371882 86184
rect 371938 86128 584960 86184
rect 371877 86126 584960 86128
rect 371877 86123 371943 86126
rect 583520 86036 584960 86126
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 342897 46338 342963 46341
rect 583520 46338 584960 46428
rect 342897 46336 584960 46338
rect 342897 46280 342902 46336
rect 342958 46280 584960 46336
rect 342897 46278 584960 46280
rect 342897 46275 342963 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 530577 19818 530643 19821
rect 583520 19818 584960 19908
rect 530577 19816 584960 19818
rect 530577 19760 530582 19816
rect 530638 19760 584960 19816
rect 530577 19758 584960 19760
rect 530577 19755 530643 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect 311157 6626 311223 6629
rect 583520 6626 584960 6716
rect 311157 6624 584960 6626
rect -960 6340 480 6580
rect 311157 6568 311162 6624
rect 311218 6568 584960 6624
rect 311157 6566 584960 6568
rect 311157 6563 311223 6566
rect 583520 6476 584960 6566
<< via3 >>
rect 296884 491650 296948 491654
rect 296884 491594 296888 491650
rect 296888 491594 296944 491650
rect 296944 491594 296948 491650
rect 296884 491590 296948 491594
rect 296964 491650 297028 491654
rect 296964 491594 296968 491650
rect 296968 491594 297024 491650
rect 297024 491594 297028 491650
rect 296964 491590 297028 491594
rect 297044 491650 297108 491654
rect 297044 491594 297048 491650
rect 297048 491594 297104 491650
rect 297104 491594 297108 491650
rect 297044 491590 297108 491594
rect 297124 491650 297188 491654
rect 297124 491594 297128 491650
rect 297128 491594 297184 491650
rect 297184 491594 297188 491650
rect 297124 491590 297188 491594
rect 296884 491570 296948 491574
rect 296884 491514 296888 491570
rect 296888 491514 296944 491570
rect 296944 491514 296948 491570
rect 296884 491510 296948 491514
rect 296964 491570 297028 491574
rect 296964 491514 296968 491570
rect 296968 491514 297024 491570
rect 297024 491514 297028 491570
rect 296964 491510 297028 491514
rect 297044 491570 297108 491574
rect 297044 491514 297048 491570
rect 297048 491514 297104 491570
rect 297104 491514 297108 491570
rect 297044 491510 297108 491514
rect 297124 491570 297188 491574
rect 297124 491514 297128 491570
rect 297128 491514 297184 491570
rect 297184 491514 297188 491570
rect 297124 491510 297188 491514
rect 296884 491490 296948 491494
rect 296884 491434 296888 491490
rect 296888 491434 296944 491490
rect 296944 491434 296948 491490
rect 296884 491430 296948 491434
rect 296964 491490 297028 491494
rect 296964 491434 296968 491490
rect 296968 491434 297024 491490
rect 297024 491434 297028 491490
rect 296964 491430 297028 491434
rect 297044 491490 297108 491494
rect 297044 491434 297048 491490
rect 297048 491434 297104 491490
rect 297104 491434 297108 491490
rect 297044 491430 297108 491434
rect 297124 491490 297188 491494
rect 297124 491434 297128 491490
rect 297128 491434 297184 491490
rect 297184 491434 297188 491490
rect 297124 491430 297188 491434
rect 296884 491410 296948 491414
rect 296884 491354 296888 491410
rect 296888 491354 296944 491410
rect 296944 491354 296948 491410
rect 296884 491350 296948 491354
rect 296964 491410 297028 491414
rect 296964 491354 296968 491410
rect 296968 491354 297024 491410
rect 297024 491354 297028 491410
rect 296964 491350 297028 491354
rect 297044 491410 297108 491414
rect 297044 491354 297048 491410
rect 297048 491354 297104 491410
rect 297104 491354 297108 491410
rect 297044 491350 297108 491354
rect 297124 491410 297188 491414
rect 297124 491354 297128 491410
rect 297128 491354 297184 491410
rect 297184 491354 297188 491410
rect 297124 491350 297188 491354
rect 303884 491650 303948 491654
rect 303884 491594 303888 491650
rect 303888 491594 303944 491650
rect 303944 491594 303948 491650
rect 303884 491590 303948 491594
rect 303964 491650 304028 491654
rect 303964 491594 303968 491650
rect 303968 491594 304024 491650
rect 304024 491594 304028 491650
rect 303964 491590 304028 491594
rect 304044 491650 304108 491654
rect 304044 491594 304048 491650
rect 304048 491594 304104 491650
rect 304104 491594 304108 491650
rect 304044 491590 304108 491594
rect 304124 491650 304188 491654
rect 304124 491594 304128 491650
rect 304128 491594 304184 491650
rect 304184 491594 304188 491650
rect 304124 491590 304188 491594
rect 303884 491570 303948 491574
rect 303884 491514 303888 491570
rect 303888 491514 303944 491570
rect 303944 491514 303948 491570
rect 303884 491510 303948 491514
rect 303964 491570 304028 491574
rect 303964 491514 303968 491570
rect 303968 491514 304024 491570
rect 304024 491514 304028 491570
rect 303964 491510 304028 491514
rect 304044 491570 304108 491574
rect 304044 491514 304048 491570
rect 304048 491514 304104 491570
rect 304104 491514 304108 491570
rect 304044 491510 304108 491514
rect 304124 491570 304188 491574
rect 304124 491514 304128 491570
rect 304128 491514 304184 491570
rect 304184 491514 304188 491570
rect 304124 491510 304188 491514
rect 303884 491490 303948 491494
rect 303884 491434 303888 491490
rect 303888 491434 303944 491490
rect 303944 491434 303948 491490
rect 303884 491430 303948 491434
rect 303964 491490 304028 491494
rect 303964 491434 303968 491490
rect 303968 491434 304024 491490
rect 304024 491434 304028 491490
rect 303964 491430 304028 491434
rect 304044 491490 304108 491494
rect 304044 491434 304048 491490
rect 304048 491434 304104 491490
rect 304104 491434 304108 491490
rect 304044 491430 304108 491434
rect 304124 491490 304188 491494
rect 304124 491434 304128 491490
rect 304128 491434 304184 491490
rect 304184 491434 304188 491490
rect 304124 491430 304188 491434
rect 310884 491650 310948 491654
rect 310884 491594 310888 491650
rect 310888 491594 310944 491650
rect 310944 491594 310948 491650
rect 310884 491590 310948 491594
rect 310964 491650 311028 491654
rect 310964 491594 310968 491650
rect 310968 491594 311024 491650
rect 311024 491594 311028 491650
rect 310964 491590 311028 491594
rect 311044 491650 311108 491654
rect 311044 491594 311048 491650
rect 311048 491594 311104 491650
rect 311104 491594 311108 491650
rect 311044 491590 311108 491594
rect 311124 491650 311188 491654
rect 311124 491594 311128 491650
rect 311128 491594 311184 491650
rect 311184 491594 311188 491650
rect 311124 491590 311188 491594
rect 310884 491570 310948 491574
rect 310884 491514 310888 491570
rect 310888 491514 310944 491570
rect 310944 491514 310948 491570
rect 310884 491510 310948 491514
rect 310964 491570 311028 491574
rect 310964 491514 310968 491570
rect 310968 491514 311024 491570
rect 311024 491514 311028 491570
rect 310964 491510 311028 491514
rect 311044 491570 311108 491574
rect 311044 491514 311048 491570
rect 311048 491514 311104 491570
rect 311104 491514 311108 491570
rect 311044 491510 311108 491514
rect 311124 491570 311188 491574
rect 311124 491514 311128 491570
rect 311128 491514 311184 491570
rect 311184 491514 311188 491570
rect 311124 491510 311188 491514
rect 303884 491410 303948 491414
rect 303884 491354 303888 491410
rect 303888 491354 303944 491410
rect 303944 491354 303948 491410
rect 303884 491350 303948 491354
rect 303964 491410 304028 491414
rect 303964 491354 303968 491410
rect 303968 491354 304024 491410
rect 304024 491354 304028 491410
rect 303964 491350 304028 491354
rect 304044 491410 304108 491414
rect 304044 491354 304048 491410
rect 304048 491354 304104 491410
rect 304104 491354 304108 491410
rect 304044 491350 304108 491354
rect 304124 491410 304188 491414
rect 304124 491354 304128 491410
rect 304128 491354 304184 491410
rect 304184 491354 304188 491410
rect 304124 491350 304188 491354
rect 310884 491490 310948 491494
rect 310884 491434 310888 491490
rect 310888 491434 310944 491490
rect 310944 491434 310948 491490
rect 310884 491430 310948 491434
rect 310964 491490 311028 491494
rect 310964 491434 310968 491490
rect 310968 491434 311024 491490
rect 311024 491434 311028 491490
rect 310964 491430 311028 491434
rect 311044 491490 311108 491494
rect 311044 491434 311048 491490
rect 311048 491434 311104 491490
rect 311104 491434 311108 491490
rect 311044 491430 311108 491434
rect 311124 491490 311188 491494
rect 311124 491434 311128 491490
rect 311128 491434 311184 491490
rect 311184 491434 311188 491490
rect 311124 491430 311188 491434
rect 310884 491410 310948 491414
rect 310884 491354 310888 491410
rect 310888 491354 310944 491410
rect 310944 491354 310948 491410
rect 310884 491350 310948 491354
rect 310964 491410 311028 491414
rect 310964 491354 310968 491410
rect 310968 491354 311024 491410
rect 311024 491354 311028 491410
rect 310964 491350 311028 491354
rect 311044 491410 311108 491414
rect 311044 491354 311048 491410
rect 311048 491354 311104 491410
rect 311104 491354 311108 491410
rect 311044 491350 311108 491354
rect 311124 491410 311188 491414
rect 311124 491354 311128 491410
rect 311128 491354 311184 491410
rect 311184 491354 311188 491410
rect 311124 491350 311188 491354
rect 295152 490534 295216 490538
rect 295152 490478 295156 490534
rect 295156 490478 295212 490534
rect 295212 490478 295216 490534
rect 295152 490474 295216 490478
rect 295232 490534 295296 490538
rect 295232 490478 295236 490534
rect 295236 490478 295292 490534
rect 295292 490478 295296 490534
rect 295232 490474 295296 490478
rect 295312 490534 295376 490538
rect 295312 490478 295316 490534
rect 295316 490478 295372 490534
rect 295372 490478 295376 490534
rect 295312 490474 295376 490478
rect 295392 490534 295456 490538
rect 295392 490478 295396 490534
rect 295396 490478 295452 490534
rect 295452 490478 295456 490534
rect 295392 490474 295456 490478
rect 295152 490454 295216 490458
rect 295152 490398 295156 490454
rect 295156 490398 295212 490454
rect 295212 490398 295216 490454
rect 295152 490394 295216 490398
rect 295232 490454 295296 490458
rect 295232 490398 295236 490454
rect 295236 490398 295292 490454
rect 295292 490398 295296 490454
rect 295232 490394 295296 490398
rect 295312 490454 295376 490458
rect 295312 490398 295316 490454
rect 295316 490398 295372 490454
rect 295372 490398 295376 490454
rect 295312 490394 295376 490398
rect 295392 490454 295456 490458
rect 295392 490398 295396 490454
rect 295396 490398 295452 490454
rect 295452 490398 295456 490454
rect 295392 490394 295456 490398
rect 295152 490374 295216 490378
rect 295152 490318 295156 490374
rect 295156 490318 295212 490374
rect 295212 490318 295216 490374
rect 295152 490314 295216 490318
rect 295232 490374 295296 490378
rect 295232 490318 295236 490374
rect 295236 490318 295292 490374
rect 295292 490318 295296 490374
rect 295232 490314 295296 490318
rect 295312 490374 295376 490378
rect 295312 490318 295316 490374
rect 295316 490318 295372 490374
rect 295372 490318 295376 490374
rect 295312 490314 295376 490318
rect 295392 490374 295456 490378
rect 295392 490318 295396 490374
rect 295396 490318 295452 490374
rect 295452 490318 295456 490374
rect 295392 490314 295456 490318
rect 303884 489478 303948 489482
rect 303884 489422 303888 489478
rect 303888 489422 303944 489478
rect 303944 489422 303948 489478
rect 303884 489418 303948 489422
rect 303964 489478 304028 489482
rect 303964 489422 303968 489478
rect 303968 489422 304024 489478
rect 304024 489422 304028 489478
rect 303964 489418 304028 489422
rect 304044 489478 304108 489482
rect 304044 489422 304048 489478
rect 304048 489422 304104 489478
rect 304104 489422 304108 489478
rect 304044 489418 304108 489422
rect 304124 489478 304188 489482
rect 304124 489422 304128 489478
rect 304128 489422 304184 489478
rect 304184 489422 304188 489478
rect 304124 489418 304188 489422
rect 303884 489398 303948 489402
rect 303884 489342 303888 489398
rect 303888 489342 303944 489398
rect 303944 489342 303948 489398
rect 303884 489338 303948 489342
rect 303964 489398 304028 489402
rect 303964 489342 303968 489398
rect 303968 489342 304024 489398
rect 304024 489342 304028 489398
rect 303964 489338 304028 489342
rect 304044 489398 304108 489402
rect 304044 489342 304048 489398
rect 304048 489342 304104 489398
rect 304104 489342 304108 489398
rect 304044 489338 304108 489342
rect 304124 489398 304188 489402
rect 304124 489342 304128 489398
rect 304128 489342 304184 489398
rect 304184 489342 304188 489398
rect 304124 489338 304188 489342
rect 303884 489318 303948 489322
rect 303884 489262 303888 489318
rect 303888 489262 303944 489318
rect 303944 489262 303948 489318
rect 303884 489258 303948 489262
rect 303964 489318 304028 489322
rect 303964 489262 303968 489318
rect 303968 489262 304024 489318
rect 304024 489262 304028 489318
rect 303964 489258 304028 489262
rect 304044 489318 304108 489322
rect 304044 489262 304048 489318
rect 304048 489262 304104 489318
rect 304104 489262 304108 489318
rect 304044 489258 304108 489262
rect 304124 489318 304188 489322
rect 304124 489262 304128 489318
rect 304128 489262 304184 489318
rect 304184 489262 304188 489318
rect 304124 489258 304188 489262
rect 303884 489238 303948 489242
rect 303884 489182 303888 489238
rect 303888 489182 303944 489238
rect 303944 489182 303948 489238
rect 303884 489178 303948 489182
rect 303964 489238 304028 489242
rect 303964 489182 303968 489238
rect 303968 489182 304024 489238
rect 304024 489182 304028 489238
rect 303964 489178 304028 489182
rect 304044 489238 304108 489242
rect 304044 489182 304048 489238
rect 304048 489182 304104 489238
rect 304104 489182 304108 489238
rect 304044 489178 304108 489182
rect 304124 489238 304188 489242
rect 304124 489182 304128 489238
rect 304128 489182 304184 489238
rect 304184 489182 304188 489238
rect 304124 489178 304188 489182
rect 310884 489478 310948 489482
rect 310884 489422 310888 489478
rect 310888 489422 310944 489478
rect 310944 489422 310948 489478
rect 310884 489418 310948 489422
rect 310964 489478 311028 489482
rect 310964 489422 310968 489478
rect 310968 489422 311024 489478
rect 311024 489422 311028 489478
rect 310964 489418 311028 489422
rect 311044 489478 311108 489482
rect 311044 489422 311048 489478
rect 311048 489422 311104 489478
rect 311104 489422 311108 489478
rect 311044 489418 311108 489422
rect 311124 489478 311188 489482
rect 311124 489422 311128 489478
rect 311128 489422 311184 489478
rect 311184 489422 311188 489478
rect 311124 489418 311188 489422
rect 310884 489398 310948 489402
rect 310884 489342 310888 489398
rect 310888 489342 310944 489398
rect 310944 489342 310948 489398
rect 310884 489338 310948 489342
rect 310964 489398 311028 489402
rect 310964 489342 310968 489398
rect 310968 489342 311024 489398
rect 311024 489342 311028 489398
rect 310964 489338 311028 489342
rect 311044 489398 311108 489402
rect 311044 489342 311048 489398
rect 311048 489342 311104 489398
rect 311104 489342 311108 489398
rect 311044 489338 311108 489342
rect 311124 489398 311188 489402
rect 311124 489342 311128 489398
rect 311128 489342 311184 489398
rect 311184 489342 311188 489398
rect 311124 489338 311188 489342
rect 310884 489318 310948 489322
rect 310884 489262 310888 489318
rect 310888 489262 310944 489318
rect 310944 489262 310948 489318
rect 310884 489258 310948 489262
rect 310964 489318 311028 489322
rect 310964 489262 310968 489318
rect 310968 489262 311024 489318
rect 311024 489262 311028 489318
rect 310964 489258 311028 489262
rect 311044 489318 311108 489322
rect 311044 489262 311048 489318
rect 311048 489262 311104 489318
rect 311104 489262 311108 489318
rect 311044 489258 311108 489262
rect 311124 489318 311188 489322
rect 311124 489262 311128 489318
rect 311128 489262 311184 489318
rect 311184 489262 311188 489318
rect 311124 489258 311188 489262
rect 310884 489238 310948 489242
rect 310884 489182 310888 489238
rect 310888 489182 310944 489238
rect 310944 489182 310948 489238
rect 310884 489178 310948 489182
rect 310964 489238 311028 489242
rect 310964 489182 310968 489238
rect 310968 489182 311024 489238
rect 311024 489182 311028 489238
rect 310964 489178 311028 489182
rect 311044 489238 311108 489242
rect 311044 489182 311048 489238
rect 311048 489182 311104 489238
rect 311104 489182 311108 489238
rect 311044 489178 311108 489182
rect 311124 489238 311188 489242
rect 311124 489182 311128 489238
rect 311128 489182 311184 489238
rect 311184 489182 311188 489238
rect 311124 489178 311188 489182
rect 296884 473110 296948 473114
rect 296884 473054 296888 473110
rect 296888 473054 296944 473110
rect 296944 473054 296948 473110
rect 296884 473050 296948 473054
rect 296964 473110 297028 473114
rect 296964 473054 296968 473110
rect 296968 473054 297024 473110
rect 297024 473054 297028 473110
rect 296964 473050 297028 473054
rect 297044 473110 297108 473114
rect 297044 473054 297048 473110
rect 297048 473054 297104 473110
rect 297104 473054 297108 473110
rect 297044 473050 297108 473054
rect 297124 473110 297188 473114
rect 297124 473054 297128 473110
rect 297128 473054 297184 473110
rect 297184 473054 297188 473110
rect 297124 473050 297188 473054
rect 296884 473030 296948 473034
rect 296884 472974 296888 473030
rect 296888 472974 296944 473030
rect 296944 472974 296948 473030
rect 296884 472970 296948 472974
rect 296964 473030 297028 473034
rect 296964 472974 296968 473030
rect 296968 472974 297024 473030
rect 297024 472974 297028 473030
rect 296964 472970 297028 472974
rect 297044 473030 297108 473034
rect 297044 472974 297048 473030
rect 297048 472974 297104 473030
rect 297104 472974 297108 473030
rect 297044 472970 297108 472974
rect 297124 473030 297188 473034
rect 297124 472974 297128 473030
rect 297128 472974 297184 473030
rect 297184 472974 297188 473030
rect 297124 472970 297188 472974
rect 303884 473110 303948 473114
rect 303884 473054 303888 473110
rect 303888 473054 303944 473110
rect 303944 473054 303948 473110
rect 303884 473050 303948 473054
rect 303964 473110 304028 473114
rect 303964 473054 303968 473110
rect 303968 473054 304024 473110
rect 304024 473054 304028 473110
rect 303964 473050 304028 473054
rect 304044 473110 304108 473114
rect 304044 473054 304048 473110
rect 304048 473054 304104 473110
rect 304104 473054 304108 473110
rect 304044 473050 304108 473054
rect 304124 473110 304188 473114
rect 304124 473054 304128 473110
rect 304128 473054 304184 473110
rect 304184 473054 304188 473110
rect 304124 473050 304188 473054
rect 296884 472950 296948 472954
rect 296884 472894 296888 472950
rect 296888 472894 296944 472950
rect 296944 472894 296948 472950
rect 296884 472890 296948 472894
rect 296964 472950 297028 472954
rect 296964 472894 296968 472950
rect 296968 472894 297024 472950
rect 297024 472894 297028 472950
rect 296964 472890 297028 472894
rect 297044 472950 297108 472954
rect 297044 472894 297048 472950
rect 297048 472894 297104 472950
rect 297104 472894 297108 472950
rect 297044 472890 297108 472894
rect 297124 472950 297188 472954
rect 297124 472894 297128 472950
rect 297128 472894 297184 472950
rect 297184 472894 297188 472950
rect 297124 472890 297188 472894
rect 303884 473030 303948 473034
rect 303884 472974 303888 473030
rect 303888 472974 303944 473030
rect 303944 472974 303948 473030
rect 303884 472970 303948 472974
rect 303964 473030 304028 473034
rect 303964 472974 303968 473030
rect 303968 472974 304024 473030
rect 304024 472974 304028 473030
rect 303964 472970 304028 472974
rect 304044 473030 304108 473034
rect 304044 472974 304048 473030
rect 304048 472974 304104 473030
rect 304104 472974 304108 473030
rect 304044 472970 304108 472974
rect 304124 473030 304188 473034
rect 304124 472974 304128 473030
rect 304128 472974 304184 473030
rect 304184 472974 304188 473030
rect 304124 472970 304188 472974
rect 296884 472870 296948 472874
rect 296884 472814 296888 472870
rect 296888 472814 296944 472870
rect 296944 472814 296948 472870
rect 296884 472810 296948 472814
rect 296964 472870 297028 472874
rect 296964 472814 296968 472870
rect 296968 472814 297024 472870
rect 297024 472814 297028 472870
rect 296964 472810 297028 472814
rect 297044 472870 297108 472874
rect 297044 472814 297048 472870
rect 297048 472814 297104 472870
rect 297104 472814 297108 472870
rect 297044 472810 297108 472814
rect 297124 472870 297188 472874
rect 297124 472814 297128 472870
rect 297128 472814 297184 472870
rect 297184 472814 297188 472870
rect 297124 472810 297188 472814
rect 303884 472950 303948 472954
rect 303884 472894 303888 472950
rect 303888 472894 303944 472950
rect 303944 472894 303948 472950
rect 303884 472890 303948 472894
rect 303964 472950 304028 472954
rect 303964 472894 303968 472950
rect 303968 472894 304024 472950
rect 304024 472894 304028 472950
rect 303964 472890 304028 472894
rect 304044 472950 304108 472954
rect 304044 472894 304048 472950
rect 304048 472894 304104 472950
rect 304104 472894 304108 472950
rect 304044 472890 304108 472894
rect 304124 472950 304188 472954
rect 304124 472894 304128 472950
rect 304128 472894 304184 472950
rect 304184 472894 304188 472950
rect 304124 472890 304188 472894
rect 303884 472870 303948 472874
rect 303884 472814 303888 472870
rect 303888 472814 303944 472870
rect 303944 472814 303948 472870
rect 303884 472810 303948 472814
rect 303964 472870 304028 472874
rect 303964 472814 303968 472870
rect 303968 472814 304024 472870
rect 304024 472814 304028 472870
rect 303964 472810 304028 472814
rect 304044 472870 304108 472874
rect 304044 472814 304048 472870
rect 304048 472814 304104 472870
rect 304104 472814 304108 472870
rect 304044 472810 304108 472814
rect 304124 472870 304188 472874
rect 304124 472814 304128 472870
rect 304128 472814 304184 472870
rect 304184 472814 304188 472870
rect 304124 472810 304188 472814
rect 310884 473110 310948 473114
rect 310884 473054 310888 473110
rect 310888 473054 310944 473110
rect 310944 473054 310948 473110
rect 310884 473050 310948 473054
rect 310964 473110 311028 473114
rect 310964 473054 310968 473110
rect 310968 473054 311024 473110
rect 311024 473054 311028 473110
rect 310964 473050 311028 473054
rect 311044 473110 311108 473114
rect 311044 473054 311048 473110
rect 311048 473054 311104 473110
rect 311104 473054 311108 473110
rect 311044 473050 311108 473054
rect 311124 473110 311188 473114
rect 311124 473054 311128 473110
rect 311128 473054 311184 473110
rect 311184 473054 311188 473110
rect 311124 473050 311188 473054
rect 310884 473030 310948 473034
rect 310884 472974 310888 473030
rect 310888 472974 310944 473030
rect 310944 472974 310948 473030
rect 310884 472970 310948 472974
rect 310964 473030 311028 473034
rect 310964 472974 310968 473030
rect 310968 472974 311024 473030
rect 311024 472974 311028 473030
rect 310964 472970 311028 472974
rect 311044 473030 311108 473034
rect 311044 472974 311048 473030
rect 311048 472974 311104 473030
rect 311104 472974 311108 473030
rect 311044 472970 311108 472974
rect 311124 473030 311188 473034
rect 311124 472974 311128 473030
rect 311128 472974 311184 473030
rect 311184 472974 311188 473030
rect 311124 472970 311188 472974
rect 310884 472950 310948 472954
rect 310884 472894 310888 472950
rect 310888 472894 310944 472950
rect 310944 472894 310948 472950
rect 310884 472890 310948 472894
rect 310964 472950 311028 472954
rect 310964 472894 310968 472950
rect 310968 472894 311024 472950
rect 311024 472894 311028 472950
rect 310964 472890 311028 472894
rect 311044 472950 311108 472954
rect 311044 472894 311048 472950
rect 311048 472894 311104 472950
rect 311104 472894 311108 472950
rect 311044 472890 311108 472894
rect 311124 472950 311188 472954
rect 311124 472894 311128 472950
rect 311128 472894 311184 472950
rect 311184 472894 311188 472950
rect 311124 472890 311188 472894
rect 310884 472870 310948 472874
rect 310884 472814 310888 472870
rect 310888 472814 310944 472870
rect 310944 472814 310948 472870
rect 310884 472810 310948 472814
rect 310964 472870 311028 472874
rect 310964 472814 310968 472870
rect 310968 472814 311024 472870
rect 311024 472814 311028 472870
rect 310964 472810 311028 472814
rect 311044 472870 311108 472874
rect 311044 472814 311048 472870
rect 311048 472814 311104 472870
rect 311104 472814 311108 472870
rect 311044 472810 311108 472814
rect 311124 472870 311188 472874
rect 311124 472814 311128 472870
rect 311128 472814 311184 472870
rect 311184 472814 311188 472870
rect 311124 472810 311188 472814
rect 302152 472009 302216 472013
rect 302152 471953 302156 472009
rect 302156 471953 302212 472009
rect 302212 471953 302216 472009
rect 302152 471949 302216 471953
rect 302232 472009 302296 472013
rect 302232 471953 302236 472009
rect 302236 471953 302292 472009
rect 302292 471953 302296 472009
rect 302232 471949 302296 471953
rect 302312 472009 302376 472013
rect 302312 471953 302316 472009
rect 302316 471953 302372 472009
rect 302372 471953 302376 472009
rect 302312 471949 302376 471953
rect 302392 472009 302456 472013
rect 302392 471953 302396 472009
rect 302396 471953 302452 472009
rect 302452 471953 302456 472009
rect 302392 471949 302456 471953
rect 302152 471929 302216 471933
rect 302152 471873 302156 471929
rect 302156 471873 302212 471929
rect 302212 471873 302216 471929
rect 302152 471869 302216 471873
rect 302232 471929 302296 471933
rect 302232 471873 302236 471929
rect 302236 471873 302292 471929
rect 302292 471873 302296 471929
rect 302232 471869 302296 471873
rect 302312 471929 302376 471933
rect 302312 471873 302316 471929
rect 302316 471873 302372 471929
rect 302372 471873 302376 471929
rect 302312 471869 302376 471873
rect 302392 471929 302456 471933
rect 302392 471873 302396 471929
rect 302396 471873 302452 471929
rect 302452 471873 302456 471929
rect 302392 471869 302456 471873
rect 302152 471849 302216 471853
rect 302152 471793 302156 471849
rect 302156 471793 302212 471849
rect 302212 471793 302216 471849
rect 302152 471789 302216 471793
rect 302232 471849 302296 471853
rect 302232 471793 302236 471849
rect 302236 471793 302292 471849
rect 302292 471793 302296 471849
rect 302232 471789 302296 471793
rect 302312 471849 302376 471853
rect 302312 471793 302316 471849
rect 302316 471793 302372 471849
rect 302372 471793 302376 471849
rect 302312 471789 302376 471793
rect 302392 471849 302456 471853
rect 302392 471793 302396 471849
rect 302396 471793 302452 471849
rect 302452 471793 302456 471849
rect 302392 471789 302456 471793
rect 302152 471769 302216 471773
rect 302152 471713 302156 471769
rect 302156 471713 302212 471769
rect 302212 471713 302216 471769
rect 302152 471709 302216 471713
rect 302232 471769 302296 471773
rect 302232 471713 302236 471769
rect 302236 471713 302292 471769
rect 302292 471713 302296 471769
rect 302232 471709 302296 471713
rect 302312 471769 302376 471773
rect 302312 471713 302316 471769
rect 302316 471713 302372 471769
rect 302372 471713 302376 471769
rect 302312 471709 302376 471713
rect 302392 471769 302456 471773
rect 302392 471713 302396 471769
rect 302396 471713 302452 471769
rect 302452 471713 302456 471769
rect 302392 471709 302456 471713
rect 309152 472009 309216 472013
rect 309152 471953 309156 472009
rect 309156 471953 309212 472009
rect 309212 471953 309216 472009
rect 309152 471949 309216 471953
rect 309232 472009 309296 472013
rect 309232 471953 309236 472009
rect 309236 471953 309292 472009
rect 309292 471953 309296 472009
rect 309232 471949 309296 471953
rect 309312 472009 309376 472013
rect 309312 471953 309316 472009
rect 309316 471953 309372 472009
rect 309372 471953 309376 472009
rect 309312 471949 309376 471953
rect 309392 472009 309456 472013
rect 309392 471953 309396 472009
rect 309396 471953 309452 472009
rect 309452 471953 309456 472009
rect 309392 471949 309456 471953
rect 309152 471929 309216 471933
rect 309152 471873 309156 471929
rect 309156 471873 309212 471929
rect 309212 471873 309216 471929
rect 309152 471869 309216 471873
rect 309232 471929 309296 471933
rect 309232 471873 309236 471929
rect 309236 471873 309292 471929
rect 309292 471873 309296 471929
rect 309232 471869 309296 471873
rect 309312 471929 309376 471933
rect 309312 471873 309316 471929
rect 309316 471873 309372 471929
rect 309372 471873 309376 471929
rect 309312 471869 309376 471873
rect 309392 471929 309456 471933
rect 309392 471873 309396 471929
rect 309396 471873 309452 471929
rect 309452 471873 309456 471929
rect 309392 471869 309456 471873
rect 309152 471849 309216 471853
rect 309152 471793 309156 471849
rect 309156 471793 309212 471849
rect 309212 471793 309216 471849
rect 309152 471789 309216 471793
rect 309232 471849 309296 471853
rect 309232 471793 309236 471849
rect 309236 471793 309292 471849
rect 309292 471793 309296 471849
rect 309232 471789 309296 471793
rect 309312 471849 309376 471853
rect 309312 471793 309316 471849
rect 309316 471793 309372 471849
rect 309372 471793 309376 471849
rect 309312 471789 309376 471793
rect 309392 471849 309456 471853
rect 309392 471793 309396 471849
rect 309396 471793 309452 471849
rect 309452 471793 309456 471849
rect 309392 471789 309456 471793
rect 309152 471769 309216 471773
rect 309152 471713 309156 471769
rect 309156 471713 309212 471769
rect 309212 471713 309216 471769
rect 309152 471709 309216 471713
rect 309232 471769 309296 471773
rect 309232 471713 309236 471769
rect 309236 471713 309292 471769
rect 309292 471713 309296 471769
rect 309232 471709 309296 471713
rect 309312 471769 309376 471773
rect 309312 471713 309316 471769
rect 309316 471713 309372 471769
rect 309372 471713 309376 471769
rect 309312 471709 309376 471713
rect 309392 471769 309456 471773
rect 309392 471713 309396 471769
rect 309396 471713 309452 471769
rect 309452 471713 309456 471769
rect 309392 471709 309456 471713
rect 296884 452054 296948 452058
rect 296884 451998 296888 452054
rect 296888 451998 296944 452054
rect 296944 451998 296948 452054
rect 296884 451994 296948 451998
rect 296964 452054 297028 452058
rect 296964 451998 296968 452054
rect 296968 451998 297024 452054
rect 297024 451998 297028 452054
rect 296964 451994 297028 451998
rect 297044 452054 297108 452058
rect 297044 451998 297048 452054
rect 297048 451998 297104 452054
rect 297104 451998 297108 452054
rect 297044 451994 297108 451998
rect 297124 452054 297188 452058
rect 297124 451998 297128 452054
rect 297128 451998 297184 452054
rect 297184 451998 297188 452054
rect 297124 451994 297188 451998
rect 296884 451974 296948 451978
rect 296884 451918 296888 451974
rect 296888 451918 296944 451974
rect 296944 451918 296948 451974
rect 296884 451914 296948 451918
rect 296964 451974 297028 451978
rect 296964 451918 296968 451974
rect 296968 451918 297024 451974
rect 297024 451918 297028 451974
rect 296964 451914 297028 451918
rect 297044 451974 297108 451978
rect 297044 451918 297048 451974
rect 297048 451918 297104 451974
rect 297104 451918 297108 451974
rect 297044 451914 297108 451918
rect 297124 451974 297188 451978
rect 297124 451918 297128 451974
rect 297128 451918 297184 451974
rect 297184 451918 297188 451974
rect 297124 451914 297188 451918
rect 296884 451894 296948 451898
rect 296884 451838 296888 451894
rect 296888 451838 296944 451894
rect 296944 451838 296948 451894
rect 296884 451834 296948 451838
rect 296964 451894 297028 451898
rect 296964 451838 296968 451894
rect 296968 451838 297024 451894
rect 297024 451838 297028 451894
rect 296964 451834 297028 451838
rect 297044 451894 297108 451898
rect 297044 451838 297048 451894
rect 297048 451838 297104 451894
rect 297104 451838 297108 451894
rect 297044 451834 297108 451838
rect 297124 451894 297188 451898
rect 297124 451838 297128 451894
rect 297128 451838 297184 451894
rect 297184 451838 297188 451894
rect 297124 451834 297188 451838
rect 296884 451814 296948 451818
rect 296884 451758 296888 451814
rect 296888 451758 296944 451814
rect 296944 451758 296948 451814
rect 296884 451754 296948 451758
rect 296964 451814 297028 451818
rect 296964 451758 296968 451814
rect 296968 451758 297024 451814
rect 297024 451758 297028 451814
rect 296964 451754 297028 451758
rect 297044 451814 297108 451818
rect 297044 451758 297048 451814
rect 297048 451758 297104 451814
rect 297104 451758 297108 451814
rect 297044 451754 297108 451758
rect 297124 451814 297188 451818
rect 297124 451758 297128 451814
rect 297128 451758 297184 451814
rect 297184 451758 297188 451814
rect 297124 451754 297188 451758
rect 296884 451734 296948 451738
rect 296884 451678 296888 451734
rect 296888 451678 296944 451734
rect 296944 451678 296948 451734
rect 296884 451674 296948 451678
rect 296964 451734 297028 451738
rect 296964 451678 296968 451734
rect 296968 451678 297024 451734
rect 297024 451678 297028 451734
rect 296964 451674 297028 451678
rect 297044 451734 297108 451738
rect 297044 451678 297048 451734
rect 297048 451678 297104 451734
rect 297104 451678 297108 451734
rect 297044 451674 297108 451678
rect 297124 451734 297188 451738
rect 297124 451678 297128 451734
rect 297128 451678 297184 451734
rect 297184 451678 297188 451734
rect 297124 451674 297188 451678
rect 296884 451654 296948 451658
rect 296884 451598 296888 451654
rect 296888 451598 296944 451654
rect 296944 451598 296948 451654
rect 296884 451594 296948 451598
rect 296964 451654 297028 451658
rect 296964 451598 296968 451654
rect 296968 451598 297024 451654
rect 297024 451598 297028 451654
rect 296964 451594 297028 451598
rect 297044 451654 297108 451658
rect 297044 451598 297048 451654
rect 297048 451598 297104 451654
rect 297104 451598 297108 451654
rect 297044 451594 297108 451598
rect 297124 451654 297188 451658
rect 297124 451598 297128 451654
rect 297128 451598 297184 451654
rect 297184 451598 297188 451654
rect 297124 451594 297188 451598
rect 296884 451574 296948 451578
rect 296884 451518 296888 451574
rect 296888 451518 296944 451574
rect 296944 451518 296948 451574
rect 296884 451514 296948 451518
rect 296964 451574 297028 451578
rect 296964 451518 296968 451574
rect 296968 451518 297024 451574
rect 297024 451518 297028 451574
rect 296964 451514 297028 451518
rect 297044 451574 297108 451578
rect 297044 451518 297048 451574
rect 297048 451518 297104 451574
rect 297104 451518 297108 451574
rect 297044 451514 297108 451518
rect 297124 451574 297188 451578
rect 297124 451518 297128 451574
rect 297128 451518 297184 451574
rect 297184 451518 297188 451574
rect 297124 451514 297188 451518
rect 296884 451494 296948 451498
rect 296884 451438 296888 451494
rect 296888 451438 296944 451494
rect 296944 451438 296948 451494
rect 296884 451434 296948 451438
rect 296964 451494 297028 451498
rect 296964 451438 296968 451494
rect 296968 451438 297024 451494
rect 297024 451438 297028 451494
rect 296964 451434 297028 451438
rect 297044 451494 297108 451498
rect 297044 451438 297048 451494
rect 297048 451438 297104 451494
rect 297104 451438 297108 451494
rect 297044 451434 297108 451438
rect 297124 451494 297188 451498
rect 297124 451438 297128 451494
rect 297128 451438 297184 451494
rect 297184 451438 297188 451494
rect 297124 451434 297188 451438
rect 296884 451414 296948 451418
rect 296884 451358 296888 451414
rect 296888 451358 296944 451414
rect 296944 451358 296948 451414
rect 296884 451354 296948 451358
rect 296964 451414 297028 451418
rect 296964 451358 296968 451414
rect 296968 451358 297024 451414
rect 297024 451358 297028 451414
rect 296964 451354 297028 451358
rect 297044 451414 297108 451418
rect 297044 451358 297048 451414
rect 297048 451358 297104 451414
rect 297104 451358 297108 451414
rect 297044 451354 297108 451358
rect 297124 451414 297188 451418
rect 297124 451358 297128 451414
rect 297128 451358 297184 451414
rect 297184 451358 297188 451414
rect 297124 451354 297188 451358
rect 296884 451334 296948 451338
rect 296884 451278 296888 451334
rect 296888 451278 296944 451334
rect 296944 451278 296948 451334
rect 296884 451274 296948 451278
rect 296964 451334 297028 451338
rect 296964 451278 296968 451334
rect 296968 451278 297024 451334
rect 297024 451278 297028 451334
rect 296964 451274 297028 451278
rect 297044 451334 297108 451338
rect 297044 451278 297048 451334
rect 297048 451278 297104 451334
rect 297104 451278 297108 451334
rect 297044 451274 297108 451278
rect 297124 451334 297188 451338
rect 297124 451278 297128 451334
rect 297128 451278 297184 451334
rect 297184 451278 297188 451334
rect 297124 451274 297188 451278
rect 303884 452054 303948 452058
rect 303884 451998 303888 452054
rect 303888 451998 303944 452054
rect 303944 451998 303948 452054
rect 303884 451994 303948 451998
rect 303964 452054 304028 452058
rect 303964 451998 303968 452054
rect 303968 451998 304024 452054
rect 304024 451998 304028 452054
rect 303964 451994 304028 451998
rect 304044 452054 304108 452058
rect 304044 451998 304048 452054
rect 304048 451998 304104 452054
rect 304104 451998 304108 452054
rect 304044 451994 304108 451998
rect 304124 452054 304188 452058
rect 304124 451998 304128 452054
rect 304128 451998 304184 452054
rect 304184 451998 304188 452054
rect 304124 451994 304188 451998
rect 303884 451974 303948 451978
rect 303884 451918 303888 451974
rect 303888 451918 303944 451974
rect 303944 451918 303948 451974
rect 303884 451914 303948 451918
rect 303964 451974 304028 451978
rect 303964 451918 303968 451974
rect 303968 451918 304024 451974
rect 304024 451918 304028 451974
rect 303964 451914 304028 451918
rect 304044 451974 304108 451978
rect 304044 451918 304048 451974
rect 304048 451918 304104 451974
rect 304104 451918 304108 451974
rect 304044 451914 304108 451918
rect 304124 451974 304188 451978
rect 304124 451918 304128 451974
rect 304128 451918 304184 451974
rect 304184 451918 304188 451974
rect 304124 451914 304188 451918
rect 303884 451894 303948 451898
rect 303884 451838 303888 451894
rect 303888 451838 303944 451894
rect 303944 451838 303948 451894
rect 303884 451834 303948 451838
rect 303964 451894 304028 451898
rect 303964 451838 303968 451894
rect 303968 451838 304024 451894
rect 304024 451838 304028 451894
rect 303964 451834 304028 451838
rect 304044 451894 304108 451898
rect 304044 451838 304048 451894
rect 304048 451838 304104 451894
rect 304104 451838 304108 451894
rect 304044 451834 304108 451838
rect 304124 451894 304188 451898
rect 304124 451838 304128 451894
rect 304128 451838 304184 451894
rect 304184 451838 304188 451894
rect 304124 451834 304188 451838
rect 303884 451814 303948 451818
rect 303884 451758 303888 451814
rect 303888 451758 303944 451814
rect 303944 451758 303948 451814
rect 303884 451754 303948 451758
rect 303964 451814 304028 451818
rect 303964 451758 303968 451814
rect 303968 451758 304024 451814
rect 304024 451758 304028 451814
rect 303964 451754 304028 451758
rect 304044 451814 304108 451818
rect 304044 451758 304048 451814
rect 304048 451758 304104 451814
rect 304104 451758 304108 451814
rect 304044 451754 304108 451758
rect 304124 451814 304188 451818
rect 304124 451758 304128 451814
rect 304128 451758 304184 451814
rect 304184 451758 304188 451814
rect 304124 451754 304188 451758
rect 310915 452054 310979 452058
rect 310915 451998 310919 452054
rect 310919 451998 310975 452054
rect 310975 451998 310979 452054
rect 310915 451994 310979 451998
rect 310995 452054 311059 452058
rect 310995 451998 310999 452054
rect 310999 451998 311055 452054
rect 311055 451998 311059 452054
rect 310995 451994 311059 451998
rect 310915 451974 310979 451978
rect 310915 451918 310919 451974
rect 310919 451918 310975 451974
rect 310975 451918 310979 451974
rect 310915 451914 310979 451918
rect 310995 451974 311059 451978
rect 310995 451918 310999 451974
rect 310999 451918 311055 451974
rect 311055 451918 311059 451974
rect 310995 451914 311059 451918
rect 310915 451894 310979 451898
rect 310915 451838 310919 451894
rect 310919 451838 310975 451894
rect 310975 451838 310979 451894
rect 310915 451834 310979 451838
rect 310995 451894 311059 451898
rect 310995 451838 310999 451894
rect 310999 451838 311055 451894
rect 311055 451838 311059 451894
rect 310995 451834 311059 451838
rect 303884 451734 303948 451738
rect 303884 451678 303888 451734
rect 303888 451678 303944 451734
rect 303944 451678 303948 451734
rect 303884 451674 303948 451678
rect 303964 451734 304028 451738
rect 303964 451678 303968 451734
rect 303968 451678 304024 451734
rect 304024 451678 304028 451734
rect 303964 451674 304028 451678
rect 304044 451734 304108 451738
rect 304044 451678 304048 451734
rect 304048 451678 304104 451734
rect 304104 451678 304108 451734
rect 304044 451674 304108 451678
rect 304124 451734 304188 451738
rect 304124 451678 304128 451734
rect 304128 451678 304184 451734
rect 304184 451678 304188 451734
rect 304124 451674 304188 451678
rect 310915 451814 310979 451818
rect 310915 451758 310919 451814
rect 310919 451758 310975 451814
rect 310975 451758 310979 451814
rect 310915 451754 310979 451758
rect 310995 451814 311059 451818
rect 310995 451758 310999 451814
rect 310999 451758 311055 451814
rect 311055 451758 311059 451814
rect 310995 451754 311059 451758
rect 303884 451654 303948 451658
rect 303884 451598 303888 451654
rect 303888 451598 303944 451654
rect 303944 451598 303948 451654
rect 303884 451594 303948 451598
rect 303964 451654 304028 451658
rect 303964 451598 303968 451654
rect 303968 451598 304024 451654
rect 304024 451598 304028 451654
rect 303964 451594 304028 451598
rect 304044 451654 304108 451658
rect 304044 451598 304048 451654
rect 304048 451598 304104 451654
rect 304104 451598 304108 451654
rect 304044 451594 304108 451598
rect 304124 451654 304188 451658
rect 304124 451598 304128 451654
rect 304128 451598 304184 451654
rect 304184 451598 304188 451654
rect 304124 451594 304188 451598
rect 303884 451574 303948 451578
rect 303884 451518 303888 451574
rect 303888 451518 303944 451574
rect 303944 451518 303948 451574
rect 303884 451514 303948 451518
rect 303964 451574 304028 451578
rect 303964 451518 303968 451574
rect 303968 451518 304024 451574
rect 304024 451518 304028 451574
rect 303964 451514 304028 451518
rect 304044 451574 304108 451578
rect 304044 451518 304048 451574
rect 304048 451518 304104 451574
rect 304104 451518 304108 451574
rect 304044 451514 304108 451518
rect 304124 451574 304188 451578
rect 304124 451518 304128 451574
rect 304128 451518 304184 451574
rect 304184 451518 304188 451574
rect 304124 451514 304188 451518
rect 303884 451494 303948 451498
rect 303884 451438 303888 451494
rect 303888 451438 303944 451494
rect 303944 451438 303948 451494
rect 303884 451434 303948 451438
rect 303964 451494 304028 451498
rect 303964 451438 303968 451494
rect 303968 451438 304024 451494
rect 304024 451438 304028 451494
rect 303964 451434 304028 451438
rect 304044 451494 304108 451498
rect 304044 451438 304048 451494
rect 304048 451438 304104 451494
rect 304104 451438 304108 451494
rect 304044 451434 304108 451438
rect 304124 451494 304188 451498
rect 304124 451438 304128 451494
rect 304128 451438 304184 451494
rect 304184 451438 304188 451494
rect 304124 451434 304188 451438
rect 310915 451734 310979 451738
rect 310915 451678 310919 451734
rect 310919 451678 310975 451734
rect 310975 451678 310979 451734
rect 310915 451674 310979 451678
rect 310995 451734 311059 451738
rect 310995 451678 310999 451734
rect 310999 451678 311055 451734
rect 311055 451678 311059 451734
rect 310995 451674 311059 451678
rect 310915 451654 310979 451658
rect 310915 451598 310919 451654
rect 310919 451598 310975 451654
rect 310975 451598 310979 451654
rect 310915 451594 310979 451598
rect 310995 451654 311059 451658
rect 310995 451598 310999 451654
rect 310999 451598 311055 451654
rect 311055 451598 311059 451654
rect 310995 451594 311059 451598
rect 310915 451574 310979 451578
rect 310915 451518 310919 451574
rect 310919 451518 310975 451574
rect 310975 451518 310979 451574
rect 310915 451514 310979 451518
rect 310995 451574 311059 451578
rect 310995 451518 310999 451574
rect 310999 451518 311055 451574
rect 311055 451518 311059 451574
rect 310995 451514 311059 451518
rect 310915 451494 310979 451498
rect 310915 451438 310919 451494
rect 310919 451438 310975 451494
rect 310975 451438 310979 451494
rect 310915 451434 310979 451438
rect 310995 451494 311059 451498
rect 310995 451438 310999 451494
rect 310999 451438 311055 451494
rect 311055 451438 311059 451494
rect 310995 451434 311059 451438
rect 303884 451414 303948 451418
rect 303884 451358 303888 451414
rect 303888 451358 303944 451414
rect 303944 451358 303948 451414
rect 303884 451354 303948 451358
rect 303964 451414 304028 451418
rect 303964 451358 303968 451414
rect 303968 451358 304024 451414
rect 304024 451358 304028 451414
rect 303964 451354 304028 451358
rect 304044 451414 304108 451418
rect 304044 451358 304048 451414
rect 304048 451358 304104 451414
rect 304104 451358 304108 451414
rect 304044 451354 304108 451358
rect 304124 451414 304188 451418
rect 304124 451358 304128 451414
rect 304128 451358 304184 451414
rect 304184 451358 304188 451414
rect 304124 451354 304188 451358
rect 303884 451334 303948 451338
rect 303884 451278 303888 451334
rect 303888 451278 303944 451334
rect 303944 451278 303948 451334
rect 303884 451274 303948 451278
rect 303964 451334 304028 451338
rect 303964 451278 303968 451334
rect 303968 451278 304024 451334
rect 304024 451278 304028 451334
rect 303964 451274 304028 451278
rect 304044 451334 304108 451338
rect 304044 451278 304048 451334
rect 304048 451278 304104 451334
rect 304104 451278 304108 451334
rect 304044 451274 304108 451278
rect 304124 451334 304188 451338
rect 304124 451278 304128 451334
rect 304128 451278 304184 451334
rect 304184 451278 304188 451334
rect 304124 451274 304188 451278
rect 310915 451414 310979 451418
rect 310915 451358 310919 451414
rect 310919 451358 310975 451414
rect 310975 451358 310979 451414
rect 310915 451354 310979 451358
rect 310995 451414 311059 451418
rect 310995 451358 310999 451414
rect 310999 451358 311055 451414
rect 311055 451358 311059 451414
rect 310995 451354 311059 451358
rect 310915 451334 310979 451338
rect 310915 451278 310919 451334
rect 310919 451278 310975 451334
rect 310975 451278 310979 451334
rect 310915 451274 310979 451278
rect 310995 451334 311059 451338
rect 310995 451278 310999 451334
rect 310999 451278 311055 451334
rect 311055 451278 311059 451334
rect 310995 451274 311059 451278
rect 310894 450177 310958 450181
rect 310894 450121 310898 450177
rect 310898 450121 310954 450177
rect 310954 450121 310958 450177
rect 310894 450117 310958 450121
rect 310974 450177 311038 450181
rect 310974 450121 310978 450177
rect 310978 450121 311034 450177
rect 311034 450121 311038 450177
rect 310974 450117 311038 450121
rect 311054 450177 311118 450181
rect 311054 450121 311058 450177
rect 311058 450121 311114 450177
rect 311114 450121 311118 450177
rect 311054 450117 311118 450121
rect 310894 450097 310958 450101
rect 310894 450041 310898 450097
rect 310898 450041 310954 450097
rect 310954 450041 310958 450097
rect 310894 450037 310958 450041
rect 310974 450097 311038 450101
rect 310974 450041 310978 450097
rect 310978 450041 311034 450097
rect 311034 450041 311038 450097
rect 310974 450037 311038 450041
rect 311054 450097 311118 450101
rect 311054 450041 311058 450097
rect 311058 450041 311114 450097
rect 311114 450041 311118 450097
rect 311054 450037 311118 450041
rect 310894 450017 310958 450021
rect 310894 449961 310898 450017
rect 310898 449961 310954 450017
rect 310954 449961 310958 450017
rect 310894 449957 310958 449961
rect 310974 450017 311038 450021
rect 310974 449961 310978 450017
rect 310978 449961 311034 450017
rect 311034 449961 311038 450017
rect 310974 449957 311038 449961
rect 311054 450017 311118 450021
rect 311054 449961 311058 450017
rect 311058 449961 311114 450017
rect 311114 449961 311118 450017
rect 311054 449957 311118 449961
rect 310894 449937 310958 449941
rect 310894 449881 310898 449937
rect 310898 449881 310954 449937
rect 310954 449881 310958 449937
rect 310894 449877 310958 449881
rect 310974 449937 311038 449941
rect 310974 449881 310978 449937
rect 310978 449881 311034 449937
rect 311034 449881 311038 449937
rect 310974 449877 311038 449881
rect 311054 449937 311118 449941
rect 311054 449881 311058 449937
rect 311058 449881 311114 449937
rect 311114 449881 311118 449937
rect 311054 449877 311118 449881
rect 310894 449857 310958 449861
rect 310894 449801 310898 449857
rect 310898 449801 310954 449857
rect 310954 449801 310958 449857
rect 310894 449797 310958 449801
rect 310974 449857 311038 449861
rect 310974 449801 310978 449857
rect 310978 449801 311034 449857
rect 311034 449801 311038 449857
rect 310974 449797 311038 449801
rect 311054 449857 311118 449861
rect 311054 449801 311058 449857
rect 311058 449801 311114 449857
rect 311114 449801 311118 449857
rect 311054 449797 311118 449801
rect 310894 449777 310958 449781
rect 310894 449721 310898 449777
rect 310898 449721 310954 449777
rect 310954 449721 310958 449777
rect 310894 449717 310958 449721
rect 310974 449777 311038 449781
rect 310974 449721 310978 449777
rect 310978 449721 311034 449777
rect 311034 449721 311038 449777
rect 310974 449717 311038 449721
rect 311054 449777 311118 449781
rect 311054 449721 311058 449777
rect 311058 449721 311114 449777
rect 311114 449721 311118 449777
rect 311054 449717 311118 449721
rect 310894 449697 310958 449701
rect 310894 449641 310898 449697
rect 310898 449641 310954 449697
rect 310954 449641 310958 449697
rect 310894 449637 310958 449641
rect 310974 449697 311038 449701
rect 310974 449641 310978 449697
rect 310978 449641 311034 449697
rect 311034 449641 311038 449697
rect 310974 449637 311038 449641
rect 311054 449697 311118 449701
rect 311054 449641 311058 449697
rect 311058 449641 311114 449697
rect 311114 449641 311118 449697
rect 311054 449637 311118 449641
rect 309187 429994 309251 429998
rect 309267 429994 309331 429998
rect 309347 429994 309411 429998
rect 309187 429938 309207 429994
rect 309207 429938 309231 429994
rect 309231 429938 309251 429994
rect 309267 429938 309287 429994
rect 309287 429938 309311 429994
rect 309311 429938 309331 429994
rect 309347 429938 309367 429994
rect 309367 429938 309391 429994
rect 309391 429938 309411 429994
rect 309187 429934 309251 429938
rect 309267 429934 309331 429938
rect 309347 429934 309411 429938
rect 309187 429914 309251 429918
rect 309267 429914 309331 429918
rect 309347 429914 309411 429918
rect 309187 429858 309207 429914
rect 309207 429858 309231 429914
rect 309231 429858 309251 429914
rect 309267 429858 309287 429914
rect 309287 429858 309311 429914
rect 309311 429858 309331 429914
rect 309347 429858 309367 429914
rect 309367 429858 309391 429914
rect 309391 429858 309411 429914
rect 309187 429854 309251 429858
rect 309267 429854 309331 429858
rect 309347 429854 309411 429858
rect 309187 429834 309251 429838
rect 309267 429834 309331 429838
rect 309347 429834 309411 429838
rect 309187 429778 309207 429834
rect 309207 429778 309231 429834
rect 309231 429778 309251 429834
rect 309267 429778 309287 429834
rect 309287 429778 309311 429834
rect 309311 429778 309331 429834
rect 309347 429778 309367 429834
rect 309367 429778 309391 429834
rect 309391 429778 309411 429834
rect 309187 429774 309251 429778
rect 309267 429774 309331 429778
rect 309347 429774 309411 429778
rect 309187 429754 309251 429758
rect 309267 429754 309331 429758
rect 309347 429754 309411 429758
rect 309187 429698 309207 429754
rect 309207 429698 309231 429754
rect 309231 429698 309251 429754
rect 309267 429698 309287 429754
rect 309287 429698 309311 429754
rect 309311 429698 309331 429754
rect 309347 429698 309367 429754
rect 309367 429698 309391 429754
rect 309391 429698 309411 429754
rect 309187 429694 309251 429698
rect 309267 429694 309331 429698
rect 309347 429694 309411 429698
rect 296884 410080 296948 410084
rect 296884 410024 296888 410080
rect 296888 410024 296944 410080
rect 296944 410024 296948 410080
rect 296884 410020 296948 410024
rect 296964 410080 297028 410084
rect 296964 410024 296968 410080
rect 296968 410024 297024 410080
rect 297024 410024 297028 410080
rect 296964 410020 297028 410024
rect 297044 410080 297108 410084
rect 297044 410024 297048 410080
rect 297048 410024 297104 410080
rect 297104 410024 297108 410080
rect 297044 410020 297108 410024
rect 297124 410080 297188 410084
rect 297124 410024 297128 410080
rect 297128 410024 297184 410080
rect 297184 410024 297188 410080
rect 297124 410020 297188 410024
rect 296884 410000 296948 410004
rect 296884 409944 296888 410000
rect 296888 409944 296944 410000
rect 296944 409944 296948 410000
rect 296884 409940 296948 409944
rect 296964 410000 297028 410004
rect 296964 409944 296968 410000
rect 296968 409944 297024 410000
rect 297024 409944 297028 410000
rect 296964 409940 297028 409944
rect 297044 410000 297108 410004
rect 297044 409944 297048 410000
rect 297048 409944 297104 410000
rect 297104 409944 297108 410000
rect 297044 409940 297108 409944
rect 297124 410000 297188 410004
rect 297124 409944 297128 410000
rect 297128 409944 297184 410000
rect 297184 409944 297188 410000
rect 297124 409940 297188 409944
rect 296884 409920 296948 409924
rect 296884 409864 296888 409920
rect 296888 409864 296944 409920
rect 296944 409864 296948 409920
rect 296884 409860 296948 409864
rect 296964 409920 297028 409924
rect 296964 409864 296968 409920
rect 296968 409864 297024 409920
rect 297024 409864 297028 409920
rect 296964 409860 297028 409864
rect 297044 409920 297108 409924
rect 297044 409864 297048 409920
rect 297048 409864 297104 409920
rect 297104 409864 297108 409920
rect 297044 409860 297108 409864
rect 297124 409920 297188 409924
rect 297124 409864 297128 409920
rect 297128 409864 297184 409920
rect 297184 409864 297188 409920
rect 297124 409860 297188 409864
rect 303884 410080 303948 410084
rect 303884 410024 303888 410080
rect 303888 410024 303944 410080
rect 303944 410024 303948 410080
rect 303884 410020 303948 410024
rect 303964 410080 304028 410084
rect 303964 410024 303968 410080
rect 303968 410024 304024 410080
rect 304024 410024 304028 410080
rect 303964 410020 304028 410024
rect 304044 410080 304108 410084
rect 304044 410024 304048 410080
rect 304048 410024 304104 410080
rect 304104 410024 304108 410080
rect 304044 410020 304108 410024
rect 304124 410080 304188 410084
rect 304124 410024 304128 410080
rect 304128 410024 304184 410080
rect 304184 410024 304188 410080
rect 304124 410020 304188 410024
rect 303884 410000 303948 410004
rect 303884 409944 303888 410000
rect 303888 409944 303944 410000
rect 303944 409944 303948 410000
rect 303884 409940 303948 409944
rect 303964 410000 304028 410004
rect 303964 409944 303968 410000
rect 303968 409944 304024 410000
rect 304024 409944 304028 410000
rect 303964 409940 304028 409944
rect 304044 410000 304108 410004
rect 304044 409944 304048 410000
rect 304048 409944 304104 410000
rect 304104 409944 304108 410000
rect 304044 409940 304108 409944
rect 304124 410000 304188 410004
rect 304124 409944 304128 410000
rect 304128 409944 304184 410000
rect 304184 409944 304188 410000
rect 304124 409940 304188 409944
rect 296884 409840 296948 409844
rect 296884 409784 296888 409840
rect 296888 409784 296944 409840
rect 296944 409784 296948 409840
rect 296884 409780 296948 409784
rect 296964 409840 297028 409844
rect 296964 409784 296968 409840
rect 296968 409784 297024 409840
rect 297024 409784 297028 409840
rect 296964 409780 297028 409784
rect 297044 409840 297108 409844
rect 297044 409784 297048 409840
rect 297048 409784 297104 409840
rect 297104 409784 297108 409840
rect 297044 409780 297108 409784
rect 297124 409840 297188 409844
rect 297124 409784 297128 409840
rect 297128 409784 297184 409840
rect 297184 409784 297188 409840
rect 297124 409780 297188 409784
rect 303884 409920 303948 409924
rect 303884 409864 303888 409920
rect 303888 409864 303944 409920
rect 303944 409864 303948 409920
rect 303884 409860 303948 409864
rect 303964 409920 304028 409924
rect 303964 409864 303968 409920
rect 303968 409864 304024 409920
rect 304024 409864 304028 409920
rect 303964 409860 304028 409864
rect 304044 409920 304108 409924
rect 304044 409864 304048 409920
rect 304048 409864 304104 409920
rect 304104 409864 304108 409920
rect 304044 409860 304108 409864
rect 304124 409920 304188 409924
rect 304124 409864 304128 409920
rect 304128 409864 304184 409920
rect 304184 409864 304188 409920
rect 304124 409860 304188 409864
rect 303884 409840 303948 409844
rect 303884 409784 303888 409840
rect 303888 409784 303944 409840
rect 303944 409784 303948 409840
rect 303884 409780 303948 409784
rect 303964 409840 304028 409844
rect 303964 409784 303968 409840
rect 303968 409784 304024 409840
rect 304024 409784 304028 409840
rect 303964 409780 304028 409784
rect 304044 409840 304108 409844
rect 304044 409784 304048 409840
rect 304048 409784 304104 409840
rect 304104 409784 304108 409840
rect 304044 409780 304108 409784
rect 304124 409840 304188 409844
rect 304124 409784 304128 409840
rect 304128 409784 304184 409840
rect 304184 409784 304188 409840
rect 304124 409780 304188 409784
rect 310884 410080 310948 410084
rect 310884 410024 310888 410080
rect 310888 410024 310944 410080
rect 310944 410024 310948 410080
rect 310884 410020 310948 410024
rect 310964 410080 311028 410084
rect 310964 410024 310968 410080
rect 310968 410024 311024 410080
rect 311024 410024 311028 410080
rect 310964 410020 311028 410024
rect 311044 410080 311108 410084
rect 311044 410024 311048 410080
rect 311048 410024 311104 410080
rect 311104 410024 311108 410080
rect 311044 410020 311108 410024
rect 311124 410080 311188 410084
rect 311124 410024 311128 410080
rect 311128 410024 311184 410080
rect 311184 410024 311188 410080
rect 311124 410020 311188 410024
rect 310884 410000 310948 410004
rect 310884 409944 310888 410000
rect 310888 409944 310944 410000
rect 310944 409944 310948 410000
rect 310884 409940 310948 409944
rect 310964 410000 311028 410004
rect 310964 409944 310968 410000
rect 310968 409944 311024 410000
rect 311024 409944 311028 410000
rect 310964 409940 311028 409944
rect 311044 410000 311108 410004
rect 311044 409944 311048 410000
rect 311048 409944 311104 410000
rect 311104 409944 311108 410000
rect 311044 409940 311108 409944
rect 311124 410000 311188 410004
rect 311124 409944 311128 410000
rect 311128 409944 311184 410000
rect 311184 409944 311188 410000
rect 311124 409940 311188 409944
rect 310884 409920 310948 409924
rect 310884 409864 310888 409920
rect 310888 409864 310944 409920
rect 310944 409864 310948 409920
rect 310884 409860 310948 409864
rect 310964 409920 311028 409924
rect 310964 409864 310968 409920
rect 310968 409864 311024 409920
rect 311024 409864 311028 409920
rect 310964 409860 311028 409864
rect 311044 409920 311108 409924
rect 311044 409864 311048 409920
rect 311048 409864 311104 409920
rect 311104 409864 311108 409920
rect 311044 409860 311108 409864
rect 311124 409920 311188 409924
rect 311124 409864 311128 409920
rect 311128 409864 311184 409920
rect 311184 409864 311188 409920
rect 311124 409860 311188 409864
rect 310884 409840 310948 409844
rect 310884 409784 310888 409840
rect 310888 409784 310944 409840
rect 310944 409784 310948 409840
rect 310884 409780 310948 409784
rect 310964 409840 311028 409844
rect 310964 409784 310968 409840
rect 310968 409784 311024 409840
rect 311024 409784 311028 409840
rect 310964 409780 311028 409784
rect 311044 409840 311108 409844
rect 311044 409784 311048 409840
rect 311048 409784 311104 409840
rect 311104 409784 311108 409840
rect 311044 409780 311108 409784
rect 311124 409840 311188 409844
rect 311124 409784 311128 409840
rect 311128 409784 311184 409840
rect 311184 409784 311188 409840
rect 311124 409780 311188 409784
rect 302152 408994 302216 408998
rect 302152 408938 302156 408994
rect 302156 408938 302212 408994
rect 302212 408938 302216 408994
rect 302152 408934 302216 408938
rect 302232 408994 302296 408998
rect 302232 408938 302236 408994
rect 302236 408938 302292 408994
rect 302292 408938 302296 408994
rect 302232 408934 302296 408938
rect 302312 408994 302376 408998
rect 302312 408938 302316 408994
rect 302316 408938 302372 408994
rect 302372 408938 302376 408994
rect 302312 408934 302376 408938
rect 302392 408994 302456 408998
rect 302392 408938 302396 408994
rect 302396 408938 302452 408994
rect 302452 408938 302456 408994
rect 302392 408934 302456 408938
rect 302152 408914 302216 408918
rect 302152 408858 302156 408914
rect 302156 408858 302212 408914
rect 302212 408858 302216 408914
rect 302152 408854 302216 408858
rect 302232 408914 302296 408918
rect 302232 408858 302236 408914
rect 302236 408858 302292 408914
rect 302292 408858 302296 408914
rect 302232 408854 302296 408858
rect 302312 408914 302376 408918
rect 302312 408858 302316 408914
rect 302316 408858 302372 408914
rect 302372 408858 302376 408914
rect 302312 408854 302376 408858
rect 302392 408914 302456 408918
rect 302392 408858 302396 408914
rect 302396 408858 302452 408914
rect 302452 408858 302456 408914
rect 302392 408854 302456 408858
rect 302152 408834 302216 408838
rect 302152 408778 302156 408834
rect 302156 408778 302212 408834
rect 302212 408778 302216 408834
rect 302152 408774 302216 408778
rect 302232 408834 302296 408838
rect 302232 408778 302236 408834
rect 302236 408778 302292 408834
rect 302292 408778 302296 408834
rect 302232 408774 302296 408778
rect 302312 408834 302376 408838
rect 302312 408778 302316 408834
rect 302316 408778 302372 408834
rect 302372 408778 302376 408834
rect 302312 408774 302376 408778
rect 302392 408834 302456 408838
rect 302392 408778 302396 408834
rect 302396 408778 302452 408834
rect 302452 408778 302456 408834
rect 302392 408774 302456 408778
rect 302152 408754 302216 408758
rect 302152 408698 302156 408754
rect 302156 408698 302212 408754
rect 302212 408698 302216 408754
rect 302152 408694 302216 408698
rect 302232 408754 302296 408758
rect 302232 408698 302236 408754
rect 302236 408698 302292 408754
rect 302292 408698 302296 408754
rect 302232 408694 302296 408698
rect 302312 408754 302376 408758
rect 302312 408698 302316 408754
rect 302316 408698 302372 408754
rect 302372 408698 302376 408754
rect 302312 408694 302376 408698
rect 302392 408754 302456 408758
rect 302392 408698 302396 408754
rect 302396 408698 302452 408754
rect 302452 408698 302456 408754
rect 302392 408694 302456 408698
rect 310884 407908 310948 407912
rect 310884 407852 310888 407908
rect 310888 407852 310944 407908
rect 310944 407852 310948 407908
rect 310884 407848 310948 407852
rect 310964 407908 311028 407912
rect 310964 407852 310968 407908
rect 310968 407852 311024 407908
rect 311024 407852 311028 407908
rect 310964 407848 311028 407852
rect 311044 407908 311108 407912
rect 311044 407852 311048 407908
rect 311048 407852 311104 407908
rect 311104 407852 311108 407908
rect 311044 407848 311108 407852
rect 311124 407908 311188 407912
rect 311124 407852 311128 407908
rect 311128 407852 311184 407908
rect 311184 407852 311188 407908
rect 311124 407848 311188 407852
rect 310884 407828 310948 407832
rect 310884 407772 310888 407828
rect 310888 407772 310944 407828
rect 310944 407772 310948 407828
rect 310884 407768 310948 407772
rect 310964 407828 311028 407832
rect 310964 407772 310968 407828
rect 310968 407772 311024 407828
rect 311024 407772 311028 407828
rect 310964 407768 311028 407772
rect 311044 407828 311108 407832
rect 311044 407772 311048 407828
rect 311048 407772 311104 407828
rect 311104 407772 311108 407828
rect 311044 407768 311108 407772
rect 311124 407828 311188 407832
rect 311124 407772 311128 407828
rect 311128 407772 311184 407828
rect 311184 407772 311188 407828
rect 311124 407768 311188 407772
rect 310884 407748 310948 407752
rect 310884 407692 310888 407748
rect 310888 407692 310944 407748
rect 310944 407692 310948 407748
rect 310884 407688 310948 407692
rect 310964 407748 311028 407752
rect 310964 407692 310968 407748
rect 310968 407692 311024 407748
rect 311024 407692 311028 407748
rect 310964 407688 311028 407692
rect 311044 407748 311108 407752
rect 311044 407692 311048 407748
rect 311048 407692 311104 407748
rect 311104 407692 311108 407748
rect 311044 407688 311108 407692
rect 311124 407748 311188 407752
rect 311124 407692 311128 407748
rect 311128 407692 311184 407748
rect 311184 407692 311188 407748
rect 311124 407688 311188 407692
rect 310884 407668 310948 407672
rect 310884 407612 310888 407668
rect 310888 407612 310944 407668
rect 310944 407612 310948 407668
rect 310884 407608 310948 407612
rect 310964 407668 311028 407672
rect 310964 407612 310968 407668
rect 310968 407612 311024 407668
rect 311024 407612 311028 407668
rect 310964 407608 311028 407612
rect 311044 407668 311108 407672
rect 311044 407612 311048 407668
rect 311048 407612 311104 407668
rect 311104 407612 311108 407668
rect 311044 407608 311108 407612
rect 311124 407668 311188 407672
rect 311124 407612 311128 407668
rect 311128 407612 311184 407668
rect 311184 407612 311188 407668
rect 311124 407608 311188 407612
rect 296884 389081 296948 389085
rect 296884 389025 296888 389081
rect 296888 389025 296944 389081
rect 296944 389025 296948 389081
rect 296884 389021 296948 389025
rect 296964 389081 297028 389085
rect 296964 389025 296968 389081
rect 296968 389025 297024 389081
rect 297024 389025 297028 389081
rect 296964 389021 297028 389025
rect 297044 389081 297108 389085
rect 297044 389025 297048 389081
rect 297048 389025 297104 389081
rect 297104 389025 297108 389081
rect 297044 389021 297108 389025
rect 297124 389081 297188 389085
rect 297124 389025 297128 389081
rect 297128 389025 297184 389081
rect 297184 389025 297188 389081
rect 297124 389021 297188 389025
rect 296884 389001 296948 389005
rect 296884 388945 296888 389001
rect 296888 388945 296944 389001
rect 296944 388945 296948 389001
rect 296884 388941 296948 388945
rect 296964 389001 297028 389005
rect 296964 388945 296968 389001
rect 296968 388945 297024 389001
rect 297024 388945 297028 389001
rect 296964 388941 297028 388945
rect 297044 389001 297108 389005
rect 297044 388945 297048 389001
rect 297048 388945 297104 389001
rect 297104 388945 297108 389001
rect 297044 388941 297108 388945
rect 297124 389001 297188 389005
rect 297124 388945 297128 389001
rect 297128 388945 297184 389001
rect 297184 388945 297188 389001
rect 297124 388941 297188 388945
rect 303884 389081 303948 389085
rect 303884 389025 303888 389081
rect 303888 389025 303944 389081
rect 303944 389025 303948 389081
rect 303884 389021 303948 389025
rect 303964 389081 304028 389085
rect 303964 389025 303968 389081
rect 303968 389025 304024 389081
rect 304024 389025 304028 389081
rect 303964 389021 304028 389025
rect 304044 389081 304108 389085
rect 304044 389025 304048 389081
rect 304048 389025 304104 389081
rect 304104 389025 304108 389081
rect 304044 389021 304108 389025
rect 304124 389081 304188 389085
rect 304124 389025 304128 389081
rect 304128 389025 304184 389081
rect 304184 389025 304188 389081
rect 304124 389021 304188 389025
rect 303884 389001 303948 389005
rect 303884 388945 303888 389001
rect 303888 388945 303944 389001
rect 303944 388945 303948 389001
rect 303884 388941 303948 388945
rect 303964 389001 304028 389005
rect 303964 388945 303968 389001
rect 303968 388945 304024 389001
rect 304024 388945 304028 389001
rect 303964 388941 304028 388945
rect 304044 389001 304108 389005
rect 304044 388945 304048 389001
rect 304048 388945 304104 389001
rect 304104 388945 304108 389001
rect 304044 388941 304108 388945
rect 304124 389001 304188 389005
rect 304124 388945 304128 389001
rect 304128 388945 304184 389001
rect 304184 388945 304188 389001
rect 304124 388941 304188 388945
rect 310884 389081 310948 389085
rect 310884 389025 310888 389081
rect 310888 389025 310944 389081
rect 310944 389025 310948 389081
rect 310884 389021 310948 389025
rect 310964 389081 311028 389085
rect 310964 389025 310968 389081
rect 310968 389025 311024 389081
rect 311024 389025 311028 389081
rect 310964 389021 311028 389025
rect 311044 389081 311108 389085
rect 311044 389025 311048 389081
rect 311048 389025 311104 389081
rect 311104 389025 311108 389081
rect 311044 389021 311108 389025
rect 311124 389081 311188 389085
rect 311124 389025 311128 389081
rect 311128 389025 311184 389081
rect 311184 389025 311188 389081
rect 311124 389021 311188 389025
rect 310884 389001 310948 389005
rect 310884 388945 310888 389001
rect 310888 388945 310944 389001
rect 310944 388945 310948 389001
rect 310884 388941 310948 388945
rect 310964 389001 311028 389005
rect 310964 388945 310968 389001
rect 310968 388945 311024 389001
rect 311024 388945 311028 389001
rect 310964 388941 311028 388945
rect 311044 389001 311108 389005
rect 311044 388945 311048 389001
rect 311048 388945 311104 389001
rect 311104 388945 311108 389001
rect 311044 388941 311108 388945
rect 311124 389001 311188 389005
rect 311124 388945 311128 389001
rect 311128 388945 311184 389001
rect 311184 388945 311188 389001
rect 311124 388941 311188 388945
rect 296884 388921 296948 388925
rect 296884 388865 296888 388921
rect 296888 388865 296944 388921
rect 296944 388865 296948 388921
rect 296884 388861 296948 388865
rect 296964 388921 297028 388925
rect 296964 388865 296968 388921
rect 296968 388865 297024 388921
rect 297024 388865 297028 388921
rect 296964 388861 297028 388865
rect 297044 388921 297108 388925
rect 297044 388865 297048 388921
rect 297048 388865 297104 388921
rect 297104 388865 297108 388921
rect 297044 388861 297108 388865
rect 297124 388921 297188 388925
rect 297124 388865 297128 388921
rect 297128 388865 297184 388921
rect 297184 388865 297188 388921
rect 297124 388861 297188 388865
rect 296884 388841 296948 388845
rect 296884 388785 296888 388841
rect 296888 388785 296944 388841
rect 296944 388785 296948 388841
rect 296884 388781 296948 388785
rect 296964 388841 297028 388845
rect 296964 388785 296968 388841
rect 296968 388785 297024 388841
rect 297024 388785 297028 388841
rect 296964 388781 297028 388785
rect 297044 388841 297108 388845
rect 297044 388785 297048 388841
rect 297048 388785 297104 388841
rect 297104 388785 297108 388841
rect 297044 388781 297108 388785
rect 297124 388841 297188 388845
rect 297124 388785 297128 388841
rect 297128 388785 297184 388841
rect 297184 388785 297188 388841
rect 297124 388781 297188 388785
rect 303884 388921 303948 388925
rect 303884 388865 303888 388921
rect 303888 388865 303944 388921
rect 303944 388865 303948 388921
rect 303884 388861 303948 388865
rect 303964 388921 304028 388925
rect 303964 388865 303968 388921
rect 303968 388865 304024 388921
rect 304024 388865 304028 388921
rect 303964 388861 304028 388865
rect 304044 388921 304108 388925
rect 304044 388865 304048 388921
rect 304048 388865 304104 388921
rect 304104 388865 304108 388921
rect 304044 388861 304108 388865
rect 304124 388921 304188 388925
rect 304124 388865 304128 388921
rect 304128 388865 304184 388921
rect 304184 388865 304188 388921
rect 304124 388861 304188 388865
rect 303884 388841 303948 388845
rect 303884 388785 303888 388841
rect 303888 388785 303944 388841
rect 303944 388785 303948 388841
rect 303884 388781 303948 388785
rect 303964 388841 304028 388845
rect 303964 388785 303968 388841
rect 303968 388785 304024 388841
rect 304024 388785 304028 388841
rect 303964 388781 304028 388785
rect 304044 388841 304108 388845
rect 304044 388785 304048 388841
rect 304048 388785 304104 388841
rect 304104 388785 304108 388841
rect 304044 388781 304108 388785
rect 304124 388841 304188 388845
rect 304124 388785 304128 388841
rect 304128 388785 304184 388841
rect 304184 388785 304188 388841
rect 304124 388781 304188 388785
rect 310884 388921 310948 388925
rect 310884 388865 310888 388921
rect 310888 388865 310944 388921
rect 310944 388865 310948 388921
rect 310884 388861 310948 388865
rect 310964 388921 311028 388925
rect 310964 388865 310968 388921
rect 310968 388865 311024 388921
rect 311024 388865 311028 388921
rect 310964 388861 311028 388865
rect 311044 388921 311108 388925
rect 311044 388865 311048 388921
rect 311048 388865 311104 388921
rect 311104 388865 311108 388921
rect 311044 388861 311108 388865
rect 311124 388921 311188 388925
rect 311124 388865 311128 388921
rect 311128 388865 311184 388921
rect 311184 388865 311188 388921
rect 311124 388861 311188 388865
rect 310884 388841 310948 388845
rect 310884 388785 310888 388841
rect 310888 388785 310944 388841
rect 310944 388785 310948 388841
rect 310884 388781 310948 388785
rect 310964 388841 311028 388845
rect 310964 388785 310968 388841
rect 310968 388785 311024 388841
rect 311024 388785 311028 388841
rect 310964 388781 311028 388785
rect 311044 388841 311108 388845
rect 311044 388785 311048 388841
rect 311048 388785 311104 388841
rect 311104 388785 311108 388841
rect 311044 388781 311108 388785
rect 311124 388841 311188 388845
rect 311124 388785 311128 388841
rect 311128 388785 311184 388841
rect 311184 388785 311188 388841
rect 311124 388781 311188 388785
rect 295152 387998 295216 388002
rect 295152 387942 295156 387998
rect 295156 387942 295212 387998
rect 295212 387942 295216 387998
rect 295152 387938 295216 387942
rect 295232 387998 295296 388002
rect 295232 387942 295236 387998
rect 295236 387942 295292 387998
rect 295292 387942 295296 387998
rect 295232 387938 295296 387942
rect 295312 387998 295376 388002
rect 295312 387942 295316 387998
rect 295316 387942 295372 387998
rect 295372 387942 295376 387998
rect 295312 387938 295376 387942
rect 295392 387998 295456 388002
rect 295392 387942 295396 387998
rect 295396 387942 295452 387998
rect 295452 387942 295456 387998
rect 295392 387938 295456 387942
rect 295152 387918 295216 387922
rect 295152 387862 295156 387918
rect 295156 387862 295212 387918
rect 295212 387862 295216 387918
rect 295152 387858 295216 387862
rect 295232 387918 295296 387922
rect 295232 387862 295236 387918
rect 295236 387862 295292 387918
rect 295292 387862 295296 387918
rect 295232 387858 295296 387862
rect 295312 387918 295376 387922
rect 295312 387862 295316 387918
rect 295316 387862 295372 387918
rect 295372 387862 295376 387918
rect 295312 387858 295376 387862
rect 295392 387918 295456 387922
rect 295392 387862 295396 387918
rect 295396 387862 295452 387918
rect 295452 387862 295456 387918
rect 295392 387858 295456 387862
rect 295152 387838 295216 387842
rect 295152 387782 295156 387838
rect 295156 387782 295212 387838
rect 295212 387782 295216 387838
rect 295152 387778 295216 387782
rect 295232 387838 295296 387842
rect 295232 387782 295236 387838
rect 295236 387782 295292 387838
rect 295292 387782 295296 387838
rect 295232 387778 295296 387782
rect 295312 387838 295376 387842
rect 295312 387782 295316 387838
rect 295316 387782 295372 387838
rect 295372 387782 295376 387838
rect 295312 387778 295376 387782
rect 295392 387838 295456 387842
rect 295392 387782 295396 387838
rect 295396 387782 295452 387838
rect 295452 387782 295456 387838
rect 295392 387778 295456 387782
rect 295152 387758 295216 387762
rect 295152 387702 295156 387758
rect 295156 387702 295212 387758
rect 295212 387702 295216 387758
rect 295152 387698 295216 387702
rect 295232 387758 295296 387762
rect 295232 387702 295236 387758
rect 295236 387702 295292 387758
rect 295292 387702 295296 387758
rect 295232 387698 295296 387702
rect 295312 387758 295376 387762
rect 295312 387702 295316 387758
rect 295316 387702 295372 387758
rect 295372 387702 295376 387758
rect 295312 387698 295376 387702
rect 295392 387758 295456 387762
rect 295392 387702 295396 387758
rect 295396 387702 295452 387758
rect 295452 387702 295456 387758
rect 295392 387698 295456 387702
rect 302152 387993 302216 387997
rect 302152 387937 302156 387993
rect 302156 387937 302212 387993
rect 302212 387937 302216 387993
rect 302152 387933 302216 387937
rect 302232 387993 302296 387997
rect 302232 387937 302236 387993
rect 302236 387937 302292 387993
rect 302292 387937 302296 387993
rect 302232 387933 302296 387937
rect 302312 387993 302376 387997
rect 302312 387937 302316 387993
rect 302316 387937 302372 387993
rect 302372 387937 302376 387993
rect 302312 387933 302376 387937
rect 302392 387993 302456 387997
rect 302392 387937 302396 387993
rect 302396 387937 302452 387993
rect 302452 387937 302456 387993
rect 302392 387933 302456 387937
rect 302152 387913 302216 387917
rect 302152 387857 302156 387913
rect 302156 387857 302212 387913
rect 302212 387857 302216 387913
rect 302152 387853 302216 387857
rect 302232 387913 302296 387917
rect 302232 387857 302236 387913
rect 302236 387857 302292 387913
rect 302292 387857 302296 387913
rect 302232 387853 302296 387857
rect 302312 387913 302376 387917
rect 302312 387857 302316 387913
rect 302316 387857 302372 387913
rect 302372 387857 302376 387913
rect 302312 387853 302376 387857
rect 302392 387913 302456 387917
rect 302392 387857 302396 387913
rect 302396 387857 302452 387913
rect 302452 387857 302456 387913
rect 302392 387853 302456 387857
rect 302152 387833 302216 387837
rect 302152 387777 302156 387833
rect 302156 387777 302212 387833
rect 302212 387777 302216 387833
rect 302152 387773 302216 387777
rect 302232 387833 302296 387837
rect 302232 387777 302236 387833
rect 302236 387777 302292 387833
rect 302292 387777 302296 387833
rect 302232 387773 302296 387777
rect 302312 387833 302376 387837
rect 302312 387777 302316 387833
rect 302316 387777 302372 387833
rect 302372 387777 302376 387833
rect 302312 387773 302376 387777
rect 302392 387833 302456 387837
rect 302392 387777 302396 387833
rect 302396 387777 302452 387833
rect 302452 387777 302456 387833
rect 302392 387773 302456 387777
rect 302152 387753 302216 387757
rect 302152 387697 302156 387753
rect 302156 387697 302212 387753
rect 302212 387697 302216 387753
rect 302152 387693 302216 387697
rect 302232 387753 302296 387757
rect 302232 387697 302236 387753
rect 302236 387697 302292 387753
rect 302292 387697 302296 387753
rect 302232 387693 302296 387697
rect 302312 387753 302376 387757
rect 302312 387697 302316 387753
rect 302316 387697 302372 387753
rect 302372 387697 302376 387753
rect 302312 387693 302376 387697
rect 302392 387753 302456 387757
rect 302392 387697 302396 387753
rect 302396 387697 302452 387753
rect 302452 387697 302456 387753
rect 302392 387693 302456 387697
rect 309152 387993 309216 387997
rect 309152 387937 309156 387993
rect 309156 387937 309212 387993
rect 309212 387937 309216 387993
rect 309152 387933 309216 387937
rect 309232 387993 309296 387997
rect 309232 387937 309236 387993
rect 309236 387937 309292 387993
rect 309292 387937 309296 387993
rect 309232 387933 309296 387937
rect 309312 387993 309376 387997
rect 309312 387937 309316 387993
rect 309316 387937 309372 387993
rect 309372 387937 309376 387993
rect 309312 387933 309376 387937
rect 309392 387993 309456 387997
rect 309392 387937 309396 387993
rect 309396 387937 309452 387993
rect 309452 387937 309456 387993
rect 309392 387933 309456 387937
rect 309152 387913 309216 387917
rect 309152 387857 309156 387913
rect 309156 387857 309212 387913
rect 309212 387857 309216 387913
rect 309152 387853 309216 387857
rect 309232 387913 309296 387917
rect 309232 387857 309236 387913
rect 309236 387857 309292 387913
rect 309292 387857 309296 387913
rect 309232 387853 309296 387857
rect 309312 387913 309376 387917
rect 309312 387857 309316 387913
rect 309316 387857 309372 387913
rect 309372 387857 309376 387913
rect 309312 387853 309376 387857
rect 309392 387913 309456 387917
rect 309392 387857 309396 387913
rect 309396 387857 309452 387913
rect 309452 387857 309456 387913
rect 309392 387853 309456 387857
rect 309152 387833 309216 387837
rect 309152 387777 309156 387833
rect 309156 387777 309212 387833
rect 309212 387777 309216 387833
rect 309152 387773 309216 387777
rect 309232 387833 309296 387837
rect 309232 387777 309236 387833
rect 309236 387777 309292 387833
rect 309292 387777 309296 387833
rect 309232 387773 309296 387777
rect 309312 387833 309376 387837
rect 309312 387777 309316 387833
rect 309316 387777 309372 387833
rect 309372 387777 309376 387833
rect 309312 387773 309376 387777
rect 309392 387833 309456 387837
rect 309392 387777 309396 387833
rect 309396 387777 309452 387833
rect 309452 387777 309456 387833
rect 309392 387773 309456 387777
rect 309152 387753 309216 387757
rect 309152 387697 309156 387753
rect 309156 387697 309212 387753
rect 309212 387697 309216 387753
rect 309152 387693 309216 387697
rect 309232 387753 309296 387757
rect 309232 387697 309236 387753
rect 309236 387697 309292 387753
rect 309292 387697 309296 387753
rect 309232 387693 309296 387697
rect 309312 387753 309376 387757
rect 309312 387697 309316 387753
rect 309316 387697 309372 387753
rect 309372 387697 309376 387753
rect 309312 387693 309376 387697
rect 309392 387753 309456 387757
rect 309392 387697 309396 387753
rect 309396 387697 309452 387753
rect 309452 387697 309456 387753
rect 309392 387693 309456 387697
rect 311040 387515 311104 387519
rect 311040 387459 311044 387515
rect 311044 387459 311100 387515
rect 311100 387459 311104 387515
rect 311040 387455 311104 387459
rect 303960 387398 304024 387402
rect 303960 387342 303964 387398
rect 303964 387342 304020 387398
rect 304020 387342 304024 387398
rect 303960 387338 304024 387342
rect 296884 347081 296948 347085
rect 296884 347025 296888 347081
rect 296888 347025 296944 347081
rect 296944 347025 296948 347081
rect 296884 347021 296948 347025
rect 296964 347081 297028 347085
rect 296964 347025 296968 347081
rect 296968 347025 297024 347081
rect 297024 347025 297028 347081
rect 296964 347021 297028 347025
rect 297044 347081 297108 347085
rect 297044 347025 297048 347081
rect 297048 347025 297104 347081
rect 297104 347025 297108 347081
rect 297044 347021 297108 347025
rect 297124 347081 297188 347085
rect 297124 347025 297128 347081
rect 297128 347025 297184 347081
rect 297184 347025 297188 347081
rect 297124 347021 297188 347025
rect 296884 347001 296948 347005
rect 296884 346945 296888 347001
rect 296888 346945 296944 347001
rect 296944 346945 296948 347001
rect 296884 346941 296948 346945
rect 296964 347001 297028 347005
rect 296964 346945 296968 347001
rect 296968 346945 297024 347001
rect 297024 346945 297028 347001
rect 296964 346941 297028 346945
rect 297044 347001 297108 347005
rect 297044 346945 297048 347001
rect 297048 346945 297104 347001
rect 297104 346945 297108 347001
rect 297044 346941 297108 346945
rect 297124 347001 297188 347005
rect 297124 346945 297128 347001
rect 297128 346945 297184 347001
rect 297184 346945 297188 347001
rect 297124 346941 297188 346945
rect 296884 346921 296948 346925
rect 296884 346865 296888 346921
rect 296888 346865 296944 346921
rect 296944 346865 296948 346921
rect 296884 346861 296948 346865
rect 296964 346921 297028 346925
rect 296964 346865 296968 346921
rect 296968 346865 297024 346921
rect 297024 346865 297028 346921
rect 296964 346861 297028 346865
rect 297044 346921 297108 346925
rect 297044 346865 297048 346921
rect 297048 346865 297104 346921
rect 297104 346865 297108 346921
rect 297044 346861 297108 346865
rect 297124 346921 297188 346925
rect 297124 346865 297128 346921
rect 297128 346865 297184 346921
rect 297184 346865 297188 346921
rect 297124 346861 297188 346865
rect 303884 347081 303948 347085
rect 303884 347025 303888 347081
rect 303888 347025 303944 347081
rect 303944 347025 303948 347081
rect 303884 347021 303948 347025
rect 303964 347081 304028 347085
rect 303964 347025 303968 347081
rect 303968 347025 304024 347081
rect 304024 347025 304028 347081
rect 303964 347021 304028 347025
rect 304044 347081 304108 347085
rect 304044 347025 304048 347081
rect 304048 347025 304104 347081
rect 304104 347025 304108 347081
rect 304044 347021 304108 347025
rect 304124 347081 304188 347085
rect 304124 347025 304128 347081
rect 304128 347025 304184 347081
rect 304184 347025 304188 347081
rect 304124 347021 304188 347025
rect 303884 347001 303948 347005
rect 303884 346945 303888 347001
rect 303888 346945 303944 347001
rect 303944 346945 303948 347001
rect 303884 346941 303948 346945
rect 303964 347001 304028 347005
rect 303964 346945 303968 347001
rect 303968 346945 304024 347001
rect 304024 346945 304028 347001
rect 303964 346941 304028 346945
rect 304044 347001 304108 347005
rect 304044 346945 304048 347001
rect 304048 346945 304104 347001
rect 304104 346945 304108 347001
rect 304044 346941 304108 346945
rect 304124 347001 304188 347005
rect 304124 346945 304128 347001
rect 304128 346945 304184 347001
rect 304184 346945 304188 347001
rect 304124 346941 304188 346945
rect 296884 346841 296948 346845
rect 296884 346785 296888 346841
rect 296888 346785 296944 346841
rect 296944 346785 296948 346841
rect 296884 346781 296948 346785
rect 296964 346841 297028 346845
rect 296964 346785 296968 346841
rect 296968 346785 297024 346841
rect 297024 346785 297028 346841
rect 296964 346781 297028 346785
rect 297044 346841 297108 346845
rect 297044 346785 297048 346841
rect 297048 346785 297104 346841
rect 297104 346785 297108 346841
rect 297044 346781 297108 346785
rect 297124 346841 297188 346845
rect 297124 346785 297128 346841
rect 297128 346785 297184 346841
rect 297184 346785 297188 346841
rect 297124 346781 297188 346785
rect 303884 346921 303948 346925
rect 303884 346865 303888 346921
rect 303888 346865 303944 346921
rect 303944 346865 303948 346921
rect 303884 346861 303948 346865
rect 303964 346921 304028 346925
rect 303964 346865 303968 346921
rect 303968 346865 304024 346921
rect 304024 346865 304028 346921
rect 303964 346861 304028 346865
rect 304044 346921 304108 346925
rect 304044 346865 304048 346921
rect 304048 346865 304104 346921
rect 304104 346865 304108 346921
rect 304044 346861 304108 346865
rect 304124 346921 304188 346925
rect 304124 346865 304128 346921
rect 304128 346865 304184 346921
rect 304184 346865 304188 346921
rect 304124 346861 304188 346865
rect 303884 346841 303948 346845
rect 303884 346785 303888 346841
rect 303888 346785 303944 346841
rect 303944 346785 303948 346841
rect 303884 346781 303948 346785
rect 303964 346841 304028 346845
rect 303964 346785 303968 346841
rect 303968 346785 304024 346841
rect 304024 346785 304028 346841
rect 303964 346781 304028 346785
rect 304044 346841 304108 346845
rect 304044 346785 304048 346841
rect 304048 346785 304104 346841
rect 304104 346785 304108 346841
rect 304044 346781 304108 346785
rect 304124 346841 304188 346845
rect 304124 346785 304128 346841
rect 304128 346785 304184 346841
rect 304184 346785 304188 346841
rect 304124 346781 304188 346785
rect 302152 345979 302216 345983
rect 302152 345923 302156 345979
rect 302156 345923 302212 345979
rect 302212 345923 302216 345979
rect 302152 345919 302216 345923
rect 302232 345979 302296 345983
rect 302232 345923 302236 345979
rect 302236 345923 302292 345979
rect 302292 345923 302296 345979
rect 302232 345919 302296 345923
rect 302312 345979 302376 345983
rect 302312 345923 302316 345979
rect 302316 345923 302372 345979
rect 302372 345923 302376 345979
rect 302312 345919 302376 345923
rect 302392 345979 302456 345983
rect 302392 345923 302396 345979
rect 302396 345923 302452 345979
rect 302452 345923 302456 345979
rect 302392 345919 302456 345923
rect 302152 345899 302216 345903
rect 302152 345843 302156 345899
rect 302156 345843 302212 345899
rect 302212 345843 302216 345899
rect 302152 345839 302216 345843
rect 302232 345899 302296 345903
rect 302232 345843 302236 345899
rect 302236 345843 302292 345899
rect 302292 345843 302296 345899
rect 302232 345839 302296 345843
rect 302312 345899 302376 345903
rect 302312 345843 302316 345899
rect 302316 345843 302372 345899
rect 302372 345843 302376 345899
rect 302312 345839 302376 345843
rect 302392 345899 302456 345903
rect 302392 345843 302396 345899
rect 302396 345843 302452 345899
rect 302452 345843 302456 345899
rect 302392 345839 302456 345843
rect 302152 345819 302216 345823
rect 302152 345763 302156 345819
rect 302156 345763 302212 345819
rect 302212 345763 302216 345819
rect 302152 345759 302216 345763
rect 302232 345819 302296 345823
rect 302232 345763 302236 345819
rect 302236 345763 302292 345819
rect 302292 345763 302296 345819
rect 302232 345759 302296 345763
rect 302312 345819 302376 345823
rect 302312 345763 302316 345819
rect 302316 345763 302372 345819
rect 302372 345763 302376 345819
rect 302312 345759 302376 345763
rect 302392 345819 302456 345823
rect 302392 345763 302396 345819
rect 302396 345763 302452 345819
rect 302452 345763 302456 345819
rect 302392 345759 302456 345763
rect 302152 345739 302216 345743
rect 302152 345683 302156 345739
rect 302156 345683 302212 345739
rect 302212 345683 302216 345739
rect 302152 345679 302216 345683
rect 302232 345739 302296 345743
rect 302232 345683 302236 345739
rect 302236 345683 302292 345739
rect 302292 345683 302296 345739
rect 302232 345679 302296 345683
rect 302312 345739 302376 345743
rect 302312 345683 302316 345739
rect 302316 345683 302372 345739
rect 302372 345683 302376 345739
rect 302312 345679 302376 345683
rect 302392 345739 302456 345743
rect 302392 345683 302396 345739
rect 302396 345683 302452 345739
rect 302452 345683 302456 345739
rect 302392 345679 302456 345683
rect 309152 345979 309216 345983
rect 309152 345923 309156 345979
rect 309156 345923 309212 345979
rect 309212 345923 309216 345979
rect 309152 345919 309216 345923
rect 309232 345979 309296 345983
rect 309232 345923 309236 345979
rect 309236 345923 309292 345979
rect 309292 345923 309296 345979
rect 309232 345919 309296 345923
rect 309312 345979 309376 345983
rect 309312 345923 309316 345979
rect 309316 345923 309372 345979
rect 309372 345923 309376 345979
rect 309312 345919 309376 345923
rect 309392 345979 309456 345983
rect 309392 345923 309396 345979
rect 309396 345923 309452 345979
rect 309452 345923 309456 345979
rect 309392 345919 309456 345923
rect 309152 345899 309216 345903
rect 309152 345843 309156 345899
rect 309156 345843 309212 345899
rect 309212 345843 309216 345899
rect 309152 345839 309216 345843
rect 309232 345899 309296 345903
rect 309232 345843 309236 345899
rect 309236 345843 309292 345899
rect 309292 345843 309296 345899
rect 309232 345839 309296 345843
rect 309312 345899 309376 345903
rect 309312 345843 309316 345899
rect 309316 345843 309372 345899
rect 309372 345843 309376 345899
rect 309312 345839 309376 345843
rect 309392 345899 309456 345903
rect 309392 345843 309396 345899
rect 309396 345843 309452 345899
rect 309452 345843 309456 345899
rect 309392 345839 309456 345843
rect 309152 345819 309216 345823
rect 309152 345763 309156 345819
rect 309156 345763 309212 345819
rect 309212 345763 309216 345819
rect 309152 345759 309216 345763
rect 309232 345819 309296 345823
rect 309232 345763 309236 345819
rect 309236 345763 309292 345819
rect 309292 345763 309296 345819
rect 309232 345759 309296 345763
rect 309312 345819 309376 345823
rect 309312 345763 309316 345819
rect 309316 345763 309372 345819
rect 309372 345763 309376 345819
rect 309312 345759 309376 345763
rect 309392 345819 309456 345823
rect 309392 345763 309396 345819
rect 309396 345763 309452 345819
rect 309452 345763 309456 345819
rect 309392 345759 309456 345763
rect 309152 345739 309216 345743
rect 309152 345683 309156 345739
rect 309156 345683 309212 345739
rect 309212 345683 309216 345739
rect 309152 345679 309216 345683
rect 309232 345739 309296 345743
rect 309232 345683 309236 345739
rect 309236 345683 309292 345739
rect 309292 345683 309296 345739
rect 309232 345679 309296 345683
rect 309312 345739 309376 345743
rect 309312 345683 309316 345739
rect 309316 345683 309372 345739
rect 309372 345683 309376 345739
rect 309312 345679 309376 345683
rect 309392 345739 309456 345743
rect 309392 345683 309396 345739
rect 309396 345683 309452 345739
rect 309452 345683 309456 345739
rect 309392 345679 309456 345683
rect 296884 326080 296948 326084
rect 296884 326024 296888 326080
rect 296888 326024 296944 326080
rect 296944 326024 296948 326080
rect 296884 326020 296948 326024
rect 296964 326080 297028 326084
rect 296964 326024 296968 326080
rect 296968 326024 297024 326080
rect 297024 326024 297028 326080
rect 296964 326020 297028 326024
rect 297044 326080 297108 326084
rect 297044 326024 297048 326080
rect 297048 326024 297104 326080
rect 297104 326024 297108 326080
rect 297044 326020 297108 326024
rect 297124 326080 297188 326084
rect 297124 326024 297128 326080
rect 297128 326024 297184 326080
rect 297184 326024 297188 326080
rect 297124 326020 297188 326024
rect 296884 326000 296948 326004
rect 296884 325944 296888 326000
rect 296888 325944 296944 326000
rect 296944 325944 296948 326000
rect 296884 325940 296948 325944
rect 296964 326000 297028 326004
rect 296964 325944 296968 326000
rect 296968 325944 297024 326000
rect 297024 325944 297028 326000
rect 296964 325940 297028 325944
rect 297044 326000 297108 326004
rect 297044 325944 297048 326000
rect 297048 325944 297104 326000
rect 297104 325944 297108 326000
rect 297044 325940 297108 325944
rect 297124 326000 297188 326004
rect 297124 325944 297128 326000
rect 297128 325944 297184 326000
rect 297184 325944 297188 326000
rect 297124 325940 297188 325944
rect 303884 326080 303948 326084
rect 303884 326024 303888 326080
rect 303888 326024 303944 326080
rect 303944 326024 303948 326080
rect 303884 326020 303948 326024
rect 303964 326080 304028 326084
rect 303964 326024 303968 326080
rect 303968 326024 304024 326080
rect 304024 326024 304028 326080
rect 303964 326020 304028 326024
rect 304044 326080 304108 326084
rect 304044 326024 304048 326080
rect 304048 326024 304104 326080
rect 304104 326024 304108 326080
rect 304044 326020 304108 326024
rect 304124 326080 304188 326084
rect 304124 326024 304128 326080
rect 304128 326024 304184 326080
rect 304184 326024 304188 326080
rect 304124 326020 304188 326024
rect 296884 325920 296948 325924
rect 296884 325864 296888 325920
rect 296888 325864 296944 325920
rect 296944 325864 296948 325920
rect 296884 325860 296948 325864
rect 296964 325920 297028 325924
rect 296964 325864 296968 325920
rect 296968 325864 297024 325920
rect 297024 325864 297028 325920
rect 296964 325860 297028 325864
rect 297044 325920 297108 325924
rect 297044 325864 297048 325920
rect 297048 325864 297104 325920
rect 297104 325864 297108 325920
rect 297044 325860 297108 325864
rect 297124 325920 297188 325924
rect 297124 325864 297128 325920
rect 297128 325864 297184 325920
rect 297184 325864 297188 325920
rect 297124 325860 297188 325864
rect 296884 325840 296948 325844
rect 296884 325784 296888 325840
rect 296888 325784 296944 325840
rect 296944 325784 296948 325840
rect 296884 325780 296948 325784
rect 296964 325840 297028 325844
rect 296964 325784 296968 325840
rect 296968 325784 297024 325840
rect 297024 325784 297028 325840
rect 296964 325780 297028 325784
rect 297044 325840 297108 325844
rect 297044 325784 297048 325840
rect 297048 325784 297104 325840
rect 297104 325784 297108 325840
rect 297044 325780 297108 325784
rect 297124 325840 297188 325844
rect 297124 325784 297128 325840
rect 297128 325784 297184 325840
rect 297184 325784 297188 325840
rect 297124 325780 297188 325784
rect 303884 326000 303948 326004
rect 303884 325944 303888 326000
rect 303888 325944 303944 326000
rect 303944 325944 303948 326000
rect 303884 325940 303948 325944
rect 303964 326000 304028 326004
rect 303964 325944 303968 326000
rect 303968 325944 304024 326000
rect 304024 325944 304028 326000
rect 303964 325940 304028 325944
rect 304044 326000 304108 326004
rect 304044 325944 304048 326000
rect 304048 325944 304104 326000
rect 304104 325944 304108 326000
rect 304044 325940 304108 325944
rect 304124 326000 304188 326004
rect 304124 325944 304128 326000
rect 304128 325944 304184 326000
rect 304184 325944 304188 326000
rect 304124 325940 304188 325944
rect 310884 326080 310948 326084
rect 310884 326024 310888 326080
rect 310888 326024 310944 326080
rect 310944 326024 310948 326080
rect 310884 326020 310948 326024
rect 310964 326080 311028 326084
rect 310964 326024 310968 326080
rect 310968 326024 311024 326080
rect 311024 326024 311028 326080
rect 310964 326020 311028 326024
rect 311044 326080 311108 326084
rect 311044 326024 311048 326080
rect 311048 326024 311104 326080
rect 311104 326024 311108 326080
rect 311044 326020 311108 326024
rect 311124 326080 311188 326084
rect 311124 326024 311128 326080
rect 311128 326024 311184 326080
rect 311184 326024 311188 326080
rect 311124 326020 311188 326024
rect 303884 325920 303948 325924
rect 303884 325864 303888 325920
rect 303888 325864 303944 325920
rect 303944 325864 303948 325920
rect 303884 325860 303948 325864
rect 303964 325920 304028 325924
rect 303964 325864 303968 325920
rect 303968 325864 304024 325920
rect 304024 325864 304028 325920
rect 303964 325860 304028 325864
rect 304044 325920 304108 325924
rect 304044 325864 304048 325920
rect 304048 325864 304104 325920
rect 304104 325864 304108 325920
rect 304044 325860 304108 325864
rect 304124 325920 304188 325924
rect 304124 325864 304128 325920
rect 304128 325864 304184 325920
rect 304184 325864 304188 325920
rect 304124 325860 304188 325864
rect 303884 325840 303948 325844
rect 303884 325784 303888 325840
rect 303888 325784 303944 325840
rect 303944 325784 303948 325840
rect 303884 325780 303948 325784
rect 303964 325840 304028 325844
rect 303964 325784 303968 325840
rect 303968 325784 304024 325840
rect 304024 325784 304028 325840
rect 303964 325780 304028 325784
rect 304044 325840 304108 325844
rect 304044 325784 304048 325840
rect 304048 325784 304104 325840
rect 304104 325784 304108 325840
rect 304044 325780 304108 325784
rect 304124 325840 304188 325844
rect 304124 325784 304128 325840
rect 304128 325784 304184 325840
rect 304184 325784 304188 325840
rect 304124 325780 304188 325784
rect 310884 326000 310948 326004
rect 310884 325944 310888 326000
rect 310888 325944 310944 326000
rect 310944 325944 310948 326000
rect 310884 325940 310948 325944
rect 310964 326000 311028 326004
rect 310964 325944 310968 326000
rect 310968 325944 311024 326000
rect 311024 325944 311028 326000
rect 310964 325940 311028 325944
rect 311044 326000 311108 326004
rect 311044 325944 311048 326000
rect 311048 325944 311104 326000
rect 311104 325944 311108 326000
rect 311044 325940 311108 325944
rect 311124 326000 311188 326004
rect 311124 325944 311128 326000
rect 311128 325944 311184 326000
rect 311184 325944 311188 326000
rect 311124 325940 311188 325944
rect 310884 325920 310948 325924
rect 310884 325864 310888 325920
rect 310888 325864 310944 325920
rect 310944 325864 310948 325920
rect 310884 325860 310948 325864
rect 310964 325920 311028 325924
rect 310964 325864 310968 325920
rect 310968 325864 311024 325920
rect 311024 325864 311028 325920
rect 310964 325860 311028 325864
rect 311044 325920 311108 325924
rect 311044 325864 311048 325920
rect 311048 325864 311104 325920
rect 311104 325864 311108 325920
rect 311044 325860 311108 325864
rect 311124 325920 311188 325924
rect 311124 325864 311128 325920
rect 311128 325864 311184 325920
rect 311184 325864 311188 325920
rect 311124 325860 311188 325864
rect 310884 325840 310948 325844
rect 310884 325784 310888 325840
rect 310888 325784 310944 325840
rect 310944 325784 310948 325840
rect 310884 325780 310948 325784
rect 310964 325840 311028 325844
rect 310964 325784 310968 325840
rect 310968 325784 311024 325840
rect 311024 325784 311028 325840
rect 310964 325780 311028 325784
rect 311044 325840 311108 325844
rect 311044 325784 311048 325840
rect 311048 325784 311104 325840
rect 311104 325784 311108 325840
rect 311044 325780 311108 325784
rect 311124 325840 311188 325844
rect 311124 325784 311128 325840
rect 311128 325784 311184 325840
rect 311184 325784 311188 325840
rect 311124 325780 311188 325784
rect 303884 323908 303948 323912
rect 303884 323852 303888 323908
rect 303888 323852 303944 323908
rect 303944 323852 303948 323908
rect 303884 323848 303948 323852
rect 303964 323908 304028 323912
rect 303964 323852 303968 323908
rect 303968 323852 304024 323908
rect 304024 323852 304028 323908
rect 303964 323848 304028 323852
rect 304044 323908 304108 323912
rect 304044 323852 304048 323908
rect 304048 323852 304104 323908
rect 304104 323852 304108 323908
rect 304044 323848 304108 323852
rect 304124 323908 304188 323912
rect 304124 323852 304128 323908
rect 304128 323852 304184 323908
rect 304184 323852 304188 323908
rect 304124 323848 304188 323852
rect 303884 323828 303948 323832
rect 303884 323772 303888 323828
rect 303888 323772 303944 323828
rect 303944 323772 303948 323828
rect 303884 323768 303948 323772
rect 303964 323828 304028 323832
rect 303964 323772 303968 323828
rect 303968 323772 304024 323828
rect 304024 323772 304028 323828
rect 303964 323768 304028 323772
rect 304044 323828 304108 323832
rect 304044 323772 304048 323828
rect 304048 323772 304104 323828
rect 304104 323772 304108 323828
rect 304044 323768 304108 323772
rect 304124 323828 304188 323832
rect 304124 323772 304128 323828
rect 304128 323772 304184 323828
rect 304184 323772 304188 323828
rect 304124 323768 304188 323772
rect 303884 323748 303948 323752
rect 303884 323692 303888 323748
rect 303888 323692 303944 323748
rect 303944 323692 303948 323748
rect 303884 323688 303948 323692
rect 303964 323748 304028 323752
rect 303964 323692 303968 323748
rect 303968 323692 304024 323748
rect 304024 323692 304028 323748
rect 303964 323688 304028 323692
rect 304044 323748 304108 323752
rect 304044 323692 304048 323748
rect 304048 323692 304104 323748
rect 304104 323692 304108 323748
rect 304044 323688 304108 323692
rect 304124 323748 304188 323752
rect 304124 323692 304128 323748
rect 304128 323692 304184 323748
rect 304184 323692 304188 323748
rect 304124 323688 304188 323692
rect 303884 323668 303948 323672
rect 303884 323612 303888 323668
rect 303888 323612 303944 323668
rect 303944 323612 303948 323668
rect 303884 323608 303948 323612
rect 303964 323668 304028 323672
rect 303964 323612 303968 323668
rect 303968 323612 304024 323668
rect 304024 323612 304028 323668
rect 303964 323608 304028 323612
rect 304044 323668 304108 323672
rect 304044 323612 304048 323668
rect 304048 323612 304104 323668
rect 304104 323612 304108 323668
rect 304044 323608 304108 323612
rect 304124 323668 304188 323672
rect 304124 323612 304128 323668
rect 304128 323612 304184 323668
rect 304184 323612 304188 323668
rect 304124 323608 304188 323612
rect 310884 323908 310948 323912
rect 310884 323852 310888 323908
rect 310888 323852 310944 323908
rect 310944 323852 310948 323908
rect 310884 323848 310948 323852
rect 310964 323908 311028 323912
rect 310964 323852 310968 323908
rect 310968 323852 311024 323908
rect 311024 323852 311028 323908
rect 310964 323848 311028 323852
rect 311044 323908 311108 323912
rect 311044 323852 311048 323908
rect 311048 323852 311104 323908
rect 311104 323852 311108 323908
rect 311044 323848 311108 323852
rect 311124 323908 311188 323912
rect 311124 323852 311128 323908
rect 311128 323852 311184 323908
rect 311184 323852 311188 323908
rect 311124 323848 311188 323852
rect 310884 323828 310948 323832
rect 310884 323772 310888 323828
rect 310888 323772 310944 323828
rect 310944 323772 310948 323828
rect 310884 323768 310948 323772
rect 310964 323828 311028 323832
rect 310964 323772 310968 323828
rect 310968 323772 311024 323828
rect 311024 323772 311028 323828
rect 310964 323768 311028 323772
rect 311044 323828 311108 323832
rect 311044 323772 311048 323828
rect 311048 323772 311104 323828
rect 311104 323772 311108 323828
rect 311044 323768 311108 323772
rect 311124 323828 311188 323832
rect 311124 323772 311128 323828
rect 311128 323772 311184 323828
rect 311184 323772 311188 323828
rect 311124 323768 311188 323772
rect 310884 323748 310948 323752
rect 310884 323692 310888 323748
rect 310888 323692 310944 323748
rect 310944 323692 310948 323748
rect 310884 323688 310948 323692
rect 310964 323748 311028 323752
rect 310964 323692 310968 323748
rect 310968 323692 311024 323748
rect 311024 323692 311028 323748
rect 310964 323688 311028 323692
rect 311044 323748 311108 323752
rect 311044 323692 311048 323748
rect 311048 323692 311104 323748
rect 311104 323692 311108 323748
rect 311044 323688 311108 323692
rect 311124 323748 311188 323752
rect 311124 323692 311128 323748
rect 311128 323692 311184 323748
rect 311184 323692 311188 323748
rect 311124 323688 311188 323692
rect 310884 323668 310948 323672
rect 310884 323612 310888 323668
rect 310888 323612 310944 323668
rect 310944 323612 310948 323668
rect 310884 323608 310948 323612
rect 310964 323668 311028 323672
rect 310964 323612 310968 323668
rect 310968 323612 311024 323668
rect 311024 323612 311028 323668
rect 310964 323608 311028 323612
rect 311044 323668 311108 323672
rect 311044 323612 311048 323668
rect 311048 323612 311104 323668
rect 311104 323612 311108 323668
rect 311044 323608 311108 323612
rect 311124 323668 311188 323672
rect 311124 323612 311128 323668
rect 311128 323612 311184 323668
rect 311184 323612 311188 323668
rect 311124 323608 311188 323612
rect 296884 305110 296948 305114
rect 296884 305054 296888 305110
rect 296888 305054 296944 305110
rect 296944 305054 296948 305110
rect 296884 305050 296948 305054
rect 296964 305110 297028 305114
rect 296964 305054 296968 305110
rect 296968 305054 297024 305110
rect 297024 305054 297028 305110
rect 296964 305050 297028 305054
rect 297044 305110 297108 305114
rect 297044 305054 297048 305110
rect 297048 305054 297104 305110
rect 297104 305054 297108 305110
rect 297044 305050 297108 305054
rect 297124 305110 297188 305114
rect 297124 305054 297128 305110
rect 297128 305054 297184 305110
rect 297184 305054 297188 305110
rect 297124 305050 297188 305054
rect 296884 305030 296948 305034
rect 296884 304974 296888 305030
rect 296888 304974 296944 305030
rect 296944 304974 296948 305030
rect 296884 304970 296948 304974
rect 296964 305030 297028 305034
rect 296964 304974 296968 305030
rect 296968 304974 297024 305030
rect 297024 304974 297028 305030
rect 296964 304970 297028 304974
rect 297044 305030 297108 305034
rect 297044 304974 297048 305030
rect 297048 304974 297104 305030
rect 297104 304974 297108 305030
rect 297044 304970 297108 304974
rect 297124 305030 297188 305034
rect 297124 304974 297128 305030
rect 297128 304974 297184 305030
rect 297184 304974 297188 305030
rect 297124 304970 297188 304974
rect 303884 305110 303948 305114
rect 303884 305054 303888 305110
rect 303888 305054 303944 305110
rect 303944 305054 303948 305110
rect 303884 305050 303948 305054
rect 303964 305110 304028 305114
rect 303964 305054 303968 305110
rect 303968 305054 304024 305110
rect 304024 305054 304028 305110
rect 303964 305050 304028 305054
rect 304044 305110 304108 305114
rect 304044 305054 304048 305110
rect 304048 305054 304104 305110
rect 304104 305054 304108 305110
rect 304044 305050 304108 305054
rect 304124 305110 304188 305114
rect 304124 305054 304128 305110
rect 304128 305054 304184 305110
rect 304184 305054 304188 305110
rect 304124 305050 304188 305054
rect 296884 304950 296948 304954
rect 296884 304894 296888 304950
rect 296888 304894 296944 304950
rect 296944 304894 296948 304950
rect 296884 304890 296948 304894
rect 296964 304950 297028 304954
rect 296964 304894 296968 304950
rect 296968 304894 297024 304950
rect 297024 304894 297028 304950
rect 296964 304890 297028 304894
rect 297044 304950 297108 304954
rect 297044 304894 297048 304950
rect 297048 304894 297104 304950
rect 297104 304894 297108 304950
rect 297044 304890 297108 304894
rect 297124 304950 297188 304954
rect 297124 304894 297128 304950
rect 297128 304894 297184 304950
rect 297184 304894 297188 304950
rect 297124 304890 297188 304894
rect 303884 305030 303948 305034
rect 303884 304974 303888 305030
rect 303888 304974 303944 305030
rect 303944 304974 303948 305030
rect 303884 304970 303948 304974
rect 303964 305030 304028 305034
rect 303964 304974 303968 305030
rect 303968 304974 304024 305030
rect 304024 304974 304028 305030
rect 303964 304970 304028 304974
rect 304044 305030 304108 305034
rect 304044 304974 304048 305030
rect 304048 304974 304104 305030
rect 304104 304974 304108 305030
rect 304044 304970 304108 304974
rect 304124 305030 304188 305034
rect 304124 304974 304128 305030
rect 304128 304974 304184 305030
rect 304184 304974 304188 305030
rect 304124 304970 304188 304974
rect 310884 305110 310948 305114
rect 310884 305054 310888 305110
rect 310888 305054 310944 305110
rect 310944 305054 310948 305110
rect 310884 305050 310948 305054
rect 310964 305110 311028 305114
rect 310964 305054 310968 305110
rect 310968 305054 311024 305110
rect 311024 305054 311028 305110
rect 310964 305050 311028 305054
rect 311044 305110 311108 305114
rect 311044 305054 311048 305110
rect 311048 305054 311104 305110
rect 311104 305054 311108 305110
rect 311044 305050 311108 305054
rect 311124 305110 311188 305114
rect 311124 305054 311128 305110
rect 311128 305054 311184 305110
rect 311184 305054 311188 305110
rect 311124 305050 311188 305054
rect 296884 304870 296948 304874
rect 296884 304814 296888 304870
rect 296888 304814 296944 304870
rect 296944 304814 296948 304870
rect 296884 304810 296948 304814
rect 296964 304870 297028 304874
rect 296964 304814 296968 304870
rect 296968 304814 297024 304870
rect 297024 304814 297028 304870
rect 296964 304810 297028 304814
rect 297044 304870 297108 304874
rect 297044 304814 297048 304870
rect 297048 304814 297104 304870
rect 297104 304814 297108 304870
rect 297044 304810 297108 304814
rect 297124 304870 297188 304874
rect 297124 304814 297128 304870
rect 297128 304814 297184 304870
rect 297184 304814 297188 304870
rect 297124 304810 297188 304814
rect 303884 304950 303948 304954
rect 303884 304894 303888 304950
rect 303888 304894 303944 304950
rect 303944 304894 303948 304950
rect 303884 304890 303948 304894
rect 303964 304950 304028 304954
rect 303964 304894 303968 304950
rect 303968 304894 304024 304950
rect 304024 304894 304028 304950
rect 303964 304890 304028 304894
rect 304044 304950 304108 304954
rect 304044 304894 304048 304950
rect 304048 304894 304104 304950
rect 304104 304894 304108 304950
rect 304044 304890 304108 304894
rect 304124 304950 304188 304954
rect 304124 304894 304128 304950
rect 304128 304894 304184 304950
rect 304184 304894 304188 304950
rect 304124 304890 304188 304894
rect 303884 304870 303948 304874
rect 303884 304814 303888 304870
rect 303888 304814 303944 304870
rect 303944 304814 303948 304870
rect 303884 304810 303948 304814
rect 303964 304870 304028 304874
rect 303964 304814 303968 304870
rect 303968 304814 304024 304870
rect 304024 304814 304028 304870
rect 303964 304810 304028 304814
rect 304044 304870 304108 304874
rect 304044 304814 304048 304870
rect 304048 304814 304104 304870
rect 304104 304814 304108 304870
rect 304044 304810 304108 304814
rect 304124 304870 304188 304874
rect 304124 304814 304128 304870
rect 304128 304814 304184 304870
rect 304184 304814 304188 304870
rect 304124 304810 304188 304814
rect 310884 305030 310948 305034
rect 310884 304974 310888 305030
rect 310888 304974 310944 305030
rect 310944 304974 310948 305030
rect 310884 304970 310948 304974
rect 310964 305030 311028 305034
rect 310964 304974 310968 305030
rect 310968 304974 311024 305030
rect 311024 304974 311028 305030
rect 310964 304970 311028 304974
rect 311044 305030 311108 305034
rect 311044 304974 311048 305030
rect 311048 304974 311104 305030
rect 311104 304974 311108 305030
rect 311044 304970 311108 304974
rect 311124 305030 311188 305034
rect 311124 304974 311128 305030
rect 311128 304974 311184 305030
rect 311184 304974 311188 305030
rect 311124 304970 311188 304974
rect 310884 304950 310948 304954
rect 310884 304894 310888 304950
rect 310888 304894 310944 304950
rect 310944 304894 310948 304950
rect 310884 304890 310948 304894
rect 310964 304950 311028 304954
rect 310964 304894 310968 304950
rect 310968 304894 311024 304950
rect 311024 304894 311028 304950
rect 310964 304890 311028 304894
rect 311044 304950 311108 304954
rect 311044 304894 311048 304950
rect 311048 304894 311104 304950
rect 311104 304894 311108 304950
rect 311044 304890 311108 304894
rect 311124 304950 311188 304954
rect 311124 304894 311128 304950
rect 311128 304894 311184 304950
rect 311184 304894 311188 304950
rect 311124 304890 311188 304894
rect 310884 304870 310948 304874
rect 310884 304814 310888 304870
rect 310888 304814 310944 304870
rect 310944 304814 310948 304870
rect 310884 304810 310948 304814
rect 310964 304870 311028 304874
rect 310964 304814 310968 304870
rect 310968 304814 311024 304870
rect 311024 304814 311028 304870
rect 310964 304810 311028 304814
rect 311044 304870 311108 304874
rect 311044 304814 311048 304870
rect 311048 304814 311104 304870
rect 311104 304814 311108 304870
rect 311044 304810 311108 304814
rect 311124 304870 311188 304874
rect 311124 304814 311128 304870
rect 311128 304814 311184 304870
rect 311184 304814 311188 304870
rect 311124 304810 311188 304814
rect 302152 304009 302216 304013
rect 302152 303953 302156 304009
rect 302156 303953 302212 304009
rect 302212 303953 302216 304009
rect 302152 303949 302216 303953
rect 302232 304009 302296 304013
rect 302232 303953 302236 304009
rect 302236 303953 302292 304009
rect 302292 303953 302296 304009
rect 302232 303949 302296 303953
rect 302312 304009 302376 304013
rect 302312 303953 302316 304009
rect 302316 303953 302372 304009
rect 302372 303953 302376 304009
rect 302312 303949 302376 303953
rect 302392 304009 302456 304013
rect 302392 303953 302396 304009
rect 302396 303953 302452 304009
rect 302452 303953 302456 304009
rect 302392 303949 302456 303953
rect 302152 303929 302216 303933
rect 302152 303873 302156 303929
rect 302156 303873 302212 303929
rect 302212 303873 302216 303929
rect 302152 303869 302216 303873
rect 302232 303929 302296 303933
rect 302232 303873 302236 303929
rect 302236 303873 302292 303929
rect 302292 303873 302296 303929
rect 302232 303869 302296 303873
rect 302312 303929 302376 303933
rect 302312 303873 302316 303929
rect 302316 303873 302372 303929
rect 302372 303873 302376 303929
rect 302312 303869 302376 303873
rect 302392 303929 302456 303933
rect 302392 303873 302396 303929
rect 302396 303873 302452 303929
rect 302452 303873 302456 303929
rect 302392 303869 302456 303873
rect 302152 303849 302216 303853
rect 302152 303793 302156 303849
rect 302156 303793 302212 303849
rect 302212 303793 302216 303849
rect 302152 303789 302216 303793
rect 302232 303849 302296 303853
rect 302232 303793 302236 303849
rect 302236 303793 302292 303849
rect 302292 303793 302296 303849
rect 302232 303789 302296 303793
rect 302312 303849 302376 303853
rect 302312 303793 302316 303849
rect 302316 303793 302372 303849
rect 302372 303793 302376 303849
rect 302312 303789 302376 303793
rect 302392 303849 302456 303853
rect 302392 303793 302396 303849
rect 302396 303793 302452 303849
rect 302452 303793 302456 303849
rect 302392 303789 302456 303793
rect 302152 303769 302216 303773
rect 302152 303713 302156 303769
rect 302156 303713 302212 303769
rect 302212 303713 302216 303769
rect 302152 303709 302216 303713
rect 302232 303769 302296 303773
rect 302232 303713 302236 303769
rect 302236 303713 302292 303769
rect 302292 303713 302296 303769
rect 302232 303709 302296 303713
rect 302312 303769 302376 303773
rect 302312 303713 302316 303769
rect 302316 303713 302372 303769
rect 302372 303713 302376 303769
rect 302312 303709 302376 303713
rect 302392 303769 302456 303773
rect 302392 303713 302396 303769
rect 302396 303713 302452 303769
rect 302452 303713 302456 303769
rect 302392 303709 302456 303713
rect 309152 304009 309216 304013
rect 309152 303953 309156 304009
rect 309156 303953 309212 304009
rect 309212 303953 309216 304009
rect 309152 303949 309216 303953
rect 309232 304009 309296 304013
rect 309232 303953 309236 304009
rect 309236 303953 309292 304009
rect 309292 303953 309296 304009
rect 309232 303949 309296 303953
rect 309312 304009 309376 304013
rect 309312 303953 309316 304009
rect 309316 303953 309372 304009
rect 309372 303953 309376 304009
rect 309312 303949 309376 303953
rect 309392 304009 309456 304013
rect 309392 303953 309396 304009
rect 309396 303953 309452 304009
rect 309452 303953 309456 304009
rect 309392 303949 309456 303953
rect 309152 303929 309216 303933
rect 309152 303873 309156 303929
rect 309156 303873 309212 303929
rect 309212 303873 309216 303929
rect 309152 303869 309216 303873
rect 309232 303929 309296 303933
rect 309232 303873 309236 303929
rect 309236 303873 309292 303929
rect 309292 303873 309296 303929
rect 309232 303869 309296 303873
rect 309312 303929 309376 303933
rect 309312 303873 309316 303929
rect 309316 303873 309372 303929
rect 309372 303873 309376 303929
rect 309312 303869 309376 303873
rect 309392 303929 309456 303933
rect 309392 303873 309396 303929
rect 309396 303873 309452 303929
rect 309452 303873 309456 303929
rect 309392 303869 309456 303873
rect 309152 303849 309216 303853
rect 309152 303793 309156 303849
rect 309156 303793 309212 303849
rect 309212 303793 309216 303849
rect 309152 303789 309216 303793
rect 309232 303849 309296 303853
rect 309232 303793 309236 303849
rect 309236 303793 309292 303849
rect 309292 303793 309296 303849
rect 309232 303789 309296 303793
rect 309312 303849 309376 303853
rect 309312 303793 309316 303849
rect 309316 303793 309372 303849
rect 309372 303793 309376 303849
rect 309312 303789 309376 303793
rect 309392 303849 309456 303853
rect 309392 303793 309396 303849
rect 309396 303793 309452 303849
rect 309452 303793 309456 303849
rect 309392 303789 309456 303793
rect 309152 303769 309216 303773
rect 309152 303713 309156 303769
rect 309156 303713 309212 303769
rect 309212 303713 309216 303769
rect 309152 303709 309216 303713
rect 309232 303769 309296 303773
rect 309232 303713 309236 303769
rect 309236 303713 309292 303769
rect 309292 303713 309296 303769
rect 309232 303709 309296 303713
rect 309312 303769 309376 303773
rect 309312 303713 309316 303769
rect 309316 303713 309372 303769
rect 309372 303713 309376 303769
rect 309312 303709 309376 303713
rect 309392 303769 309456 303773
rect 309392 303713 309396 303769
rect 309396 303713 309452 303769
rect 309452 303713 309456 303769
rect 309392 303709 309456 303713
rect 302152 282994 302216 282998
rect 302152 282938 302156 282994
rect 302156 282938 302212 282994
rect 302212 282938 302216 282994
rect 302152 282934 302216 282938
rect 302232 282994 302296 282998
rect 302232 282938 302236 282994
rect 302236 282938 302292 282994
rect 302292 282938 302296 282994
rect 302232 282934 302296 282938
rect 302312 282994 302376 282998
rect 302312 282938 302316 282994
rect 302316 282938 302372 282994
rect 302372 282938 302376 282994
rect 302312 282934 302376 282938
rect 302392 282994 302456 282998
rect 302392 282938 302396 282994
rect 302396 282938 302452 282994
rect 302452 282938 302456 282994
rect 302392 282934 302456 282938
rect 302152 282914 302216 282918
rect 302152 282858 302156 282914
rect 302156 282858 302212 282914
rect 302212 282858 302216 282914
rect 302152 282854 302216 282858
rect 302232 282914 302296 282918
rect 302232 282858 302236 282914
rect 302236 282858 302292 282914
rect 302292 282858 302296 282914
rect 302232 282854 302296 282858
rect 302312 282914 302376 282918
rect 302312 282858 302316 282914
rect 302316 282858 302372 282914
rect 302372 282858 302376 282914
rect 302312 282854 302376 282858
rect 302392 282914 302456 282918
rect 302392 282858 302396 282914
rect 302396 282858 302452 282914
rect 302452 282858 302456 282914
rect 302392 282854 302456 282858
rect 302152 282834 302216 282838
rect 302152 282778 302156 282834
rect 302156 282778 302212 282834
rect 302212 282778 302216 282834
rect 302152 282774 302216 282778
rect 302232 282834 302296 282838
rect 302232 282778 302236 282834
rect 302236 282778 302292 282834
rect 302292 282778 302296 282834
rect 302232 282774 302296 282778
rect 302312 282834 302376 282838
rect 302312 282778 302316 282834
rect 302316 282778 302372 282834
rect 302372 282778 302376 282834
rect 302312 282774 302376 282778
rect 302392 282834 302456 282838
rect 302392 282778 302396 282834
rect 302396 282778 302452 282834
rect 302452 282778 302456 282834
rect 302392 282774 302456 282778
rect 302152 282754 302216 282758
rect 302152 282698 302156 282754
rect 302156 282698 302212 282754
rect 302212 282698 302216 282754
rect 302152 282694 302216 282698
rect 302232 282754 302296 282758
rect 302232 282698 302236 282754
rect 302236 282698 302292 282754
rect 302292 282698 302296 282754
rect 302232 282694 302296 282698
rect 302312 282754 302376 282758
rect 302312 282698 302316 282754
rect 302316 282698 302372 282754
rect 302372 282698 302376 282754
rect 302312 282694 302376 282698
rect 302392 282754 302456 282758
rect 302392 282698 302396 282754
rect 302396 282698 302452 282754
rect 302452 282698 302456 282754
rect 302392 282694 302456 282698
rect 309152 282995 309216 282999
rect 309152 282939 309156 282995
rect 309156 282939 309212 282995
rect 309212 282939 309216 282995
rect 309152 282935 309216 282939
rect 309232 282995 309296 282999
rect 309232 282939 309236 282995
rect 309236 282939 309292 282995
rect 309292 282939 309296 282995
rect 309232 282935 309296 282939
rect 309312 282995 309376 282999
rect 309312 282939 309316 282995
rect 309316 282939 309372 282995
rect 309372 282939 309376 282995
rect 309312 282935 309376 282939
rect 309392 282995 309456 282999
rect 309392 282939 309396 282995
rect 309396 282939 309452 282995
rect 309452 282939 309456 282995
rect 309392 282935 309456 282939
rect 309152 282915 309216 282919
rect 309152 282859 309156 282915
rect 309156 282859 309212 282915
rect 309212 282859 309216 282915
rect 309152 282855 309216 282859
rect 309232 282915 309296 282919
rect 309232 282859 309236 282915
rect 309236 282859 309292 282915
rect 309292 282859 309296 282915
rect 309232 282855 309296 282859
rect 309312 282915 309376 282919
rect 309312 282859 309316 282915
rect 309316 282859 309372 282915
rect 309372 282859 309376 282915
rect 309312 282855 309376 282859
rect 309392 282915 309456 282919
rect 309392 282859 309396 282915
rect 309396 282859 309452 282915
rect 309452 282859 309456 282915
rect 309392 282855 309456 282859
rect 309152 282835 309216 282839
rect 309152 282779 309156 282835
rect 309156 282779 309212 282835
rect 309212 282779 309216 282835
rect 309152 282775 309216 282779
rect 309232 282835 309296 282839
rect 309232 282779 309236 282835
rect 309236 282779 309292 282835
rect 309292 282779 309296 282835
rect 309232 282775 309296 282779
rect 309312 282835 309376 282839
rect 309312 282779 309316 282835
rect 309316 282779 309372 282835
rect 309372 282779 309376 282835
rect 309312 282775 309376 282779
rect 309392 282835 309456 282839
rect 309392 282779 309396 282835
rect 309396 282779 309452 282835
rect 309452 282779 309456 282835
rect 309392 282775 309456 282779
rect 309152 282755 309216 282759
rect 309152 282699 309156 282755
rect 309156 282699 309212 282755
rect 309212 282699 309216 282755
rect 309152 282695 309216 282699
rect 309232 282755 309296 282759
rect 309232 282699 309236 282755
rect 309236 282699 309292 282755
rect 309292 282699 309296 282755
rect 309232 282695 309296 282699
rect 309312 282755 309376 282759
rect 309312 282699 309316 282755
rect 309316 282699 309372 282755
rect 309372 282699 309376 282755
rect 309312 282695 309376 282699
rect 309392 282755 309456 282759
rect 309392 282699 309396 282755
rect 309396 282699 309452 282755
rect 309452 282699 309456 282755
rect 309392 282695 309456 282699
rect 303884 282233 303948 282237
rect 303884 282177 303888 282233
rect 303888 282177 303944 282233
rect 303944 282177 303948 282233
rect 303884 282173 303948 282177
rect 303964 282233 304028 282237
rect 303964 282177 303968 282233
rect 303968 282177 304024 282233
rect 304024 282177 304028 282233
rect 303964 282173 304028 282177
rect 304044 282233 304108 282237
rect 304044 282177 304048 282233
rect 304048 282177 304104 282233
rect 304104 282177 304108 282233
rect 304044 282173 304108 282177
rect 304124 282233 304188 282237
rect 304124 282177 304128 282233
rect 304128 282177 304184 282233
rect 304184 282177 304188 282233
rect 304124 282173 304188 282177
rect 303884 282153 303948 282157
rect 303884 282097 303888 282153
rect 303888 282097 303944 282153
rect 303944 282097 303948 282153
rect 303884 282093 303948 282097
rect 303964 282153 304028 282157
rect 303964 282097 303968 282153
rect 303968 282097 304024 282153
rect 304024 282097 304028 282153
rect 303964 282093 304028 282097
rect 304044 282153 304108 282157
rect 304044 282097 304048 282153
rect 304048 282097 304104 282153
rect 304104 282097 304108 282153
rect 304044 282093 304108 282097
rect 304124 282153 304188 282157
rect 304124 282097 304128 282153
rect 304128 282097 304184 282153
rect 304184 282097 304188 282153
rect 304124 282093 304188 282097
rect 303884 282073 303948 282077
rect 303884 282017 303888 282073
rect 303888 282017 303944 282073
rect 303944 282017 303948 282073
rect 303884 282013 303948 282017
rect 303964 282073 304028 282077
rect 303964 282017 303968 282073
rect 303968 282017 304024 282073
rect 304024 282017 304028 282073
rect 303964 282013 304028 282017
rect 304044 282073 304108 282077
rect 304044 282017 304048 282073
rect 304048 282017 304104 282073
rect 304104 282017 304108 282073
rect 304044 282013 304108 282017
rect 304124 282073 304188 282077
rect 304124 282017 304128 282073
rect 304128 282017 304184 282073
rect 304184 282017 304188 282073
rect 304124 282013 304188 282017
rect 303884 281993 303948 281997
rect 303884 281937 303888 281993
rect 303888 281937 303944 281993
rect 303944 281937 303948 281993
rect 303884 281933 303948 281937
rect 303964 281993 304028 281997
rect 303964 281937 303968 281993
rect 303968 281937 304024 281993
rect 304024 281937 304028 281993
rect 303964 281933 304028 281937
rect 304044 281993 304108 281997
rect 304044 281937 304048 281993
rect 304048 281937 304104 281993
rect 304104 281937 304108 281993
rect 304044 281933 304108 281937
rect 304124 281993 304188 281997
rect 304124 281937 304128 281993
rect 304128 281937 304184 281993
rect 304184 281937 304188 281993
rect 304124 281933 304188 281937
rect 303884 281913 303948 281917
rect 303884 281857 303888 281913
rect 303888 281857 303944 281913
rect 303944 281857 303948 281913
rect 303884 281853 303948 281857
rect 303964 281913 304028 281917
rect 303964 281857 303968 281913
rect 303968 281857 304024 281913
rect 304024 281857 304028 281913
rect 303964 281853 304028 281857
rect 304044 281913 304108 281917
rect 304044 281857 304048 281913
rect 304048 281857 304104 281913
rect 304104 281857 304108 281913
rect 304044 281853 304108 281857
rect 304124 281913 304188 281917
rect 304124 281857 304128 281913
rect 304128 281857 304184 281913
rect 304184 281857 304188 281913
rect 304124 281853 304188 281857
rect 303884 281833 303948 281837
rect 303884 281777 303888 281833
rect 303888 281777 303944 281833
rect 303944 281777 303948 281833
rect 303884 281773 303948 281777
rect 303964 281833 304028 281837
rect 303964 281777 303968 281833
rect 303968 281777 304024 281833
rect 304024 281777 304028 281833
rect 303964 281773 304028 281777
rect 304044 281833 304108 281837
rect 304044 281777 304048 281833
rect 304048 281777 304104 281833
rect 304104 281777 304108 281833
rect 304044 281773 304108 281777
rect 304124 281833 304188 281837
rect 304124 281777 304128 281833
rect 304128 281777 304184 281833
rect 304184 281777 304188 281833
rect 304124 281773 304188 281777
rect 303884 281753 303948 281757
rect 303884 281697 303888 281753
rect 303888 281697 303944 281753
rect 303944 281697 303948 281753
rect 303884 281693 303948 281697
rect 303964 281753 304028 281757
rect 303964 281697 303968 281753
rect 303968 281697 304024 281753
rect 304024 281697 304028 281753
rect 303964 281693 304028 281697
rect 304044 281753 304108 281757
rect 304044 281697 304048 281753
rect 304048 281697 304104 281753
rect 304104 281697 304108 281753
rect 304044 281693 304108 281697
rect 304124 281753 304188 281757
rect 304124 281697 304128 281753
rect 304128 281697 304184 281753
rect 304184 281697 304188 281753
rect 304124 281693 304188 281697
rect 303884 281673 303948 281677
rect 303884 281617 303888 281673
rect 303888 281617 303944 281673
rect 303944 281617 303948 281673
rect 303884 281613 303948 281617
rect 303964 281673 304028 281677
rect 303964 281617 303968 281673
rect 303968 281617 304024 281673
rect 304024 281617 304028 281673
rect 303964 281613 304028 281617
rect 304044 281673 304108 281677
rect 304044 281617 304048 281673
rect 304048 281617 304104 281673
rect 304104 281617 304108 281673
rect 304044 281613 304108 281617
rect 304124 281673 304188 281677
rect 304124 281617 304128 281673
rect 304128 281617 304184 281673
rect 304184 281617 304188 281673
rect 304124 281613 304188 281617
rect 310884 282178 310948 282182
rect 310884 282122 310888 282178
rect 310888 282122 310944 282178
rect 310944 282122 310948 282178
rect 310884 282118 310948 282122
rect 310964 282178 311028 282182
rect 310964 282122 310968 282178
rect 310968 282122 311024 282178
rect 311024 282122 311028 282178
rect 310964 282118 311028 282122
rect 311044 282178 311108 282182
rect 311044 282122 311048 282178
rect 311048 282122 311104 282178
rect 311104 282122 311108 282178
rect 311044 282118 311108 282122
rect 311124 282178 311188 282182
rect 311124 282122 311128 282178
rect 311128 282122 311184 282178
rect 311184 282122 311188 282178
rect 311124 282118 311188 282122
rect 310884 282098 310948 282102
rect 310884 282042 310888 282098
rect 310888 282042 310944 282098
rect 310944 282042 310948 282098
rect 310884 282038 310948 282042
rect 310964 282098 311028 282102
rect 310964 282042 310968 282098
rect 310968 282042 311024 282098
rect 311024 282042 311028 282098
rect 310964 282038 311028 282042
rect 311044 282098 311108 282102
rect 311044 282042 311048 282098
rect 311048 282042 311104 282098
rect 311104 282042 311108 282098
rect 311044 282038 311108 282042
rect 311124 282098 311188 282102
rect 311124 282042 311128 282098
rect 311128 282042 311184 282098
rect 311184 282042 311188 282098
rect 311124 282038 311188 282042
rect 310884 282018 310948 282022
rect 310884 281962 310888 282018
rect 310888 281962 310944 282018
rect 310944 281962 310948 282018
rect 310884 281958 310948 281962
rect 310964 282018 311028 282022
rect 310964 281962 310968 282018
rect 310968 281962 311024 282018
rect 311024 281962 311028 282018
rect 310964 281958 311028 281962
rect 311044 282018 311108 282022
rect 311044 281962 311048 282018
rect 311048 281962 311104 282018
rect 311104 281962 311108 282018
rect 311044 281958 311108 281962
rect 311124 282018 311188 282022
rect 311124 281962 311128 282018
rect 311128 281962 311184 282018
rect 311184 281962 311188 282018
rect 311124 281958 311188 281962
rect 310884 281938 310948 281942
rect 310884 281882 310888 281938
rect 310888 281882 310944 281938
rect 310944 281882 310948 281938
rect 310884 281878 310948 281882
rect 310964 281938 311028 281942
rect 310964 281882 310968 281938
rect 310968 281882 311024 281938
rect 311024 281882 311028 281938
rect 310964 281878 311028 281882
rect 311044 281938 311108 281942
rect 311044 281882 311048 281938
rect 311048 281882 311104 281938
rect 311104 281882 311108 281938
rect 311044 281878 311108 281882
rect 311124 281938 311188 281942
rect 311124 281882 311128 281938
rect 311128 281882 311184 281938
rect 311184 281882 311188 281938
rect 311124 281878 311188 281882
rect 310884 281858 310948 281862
rect 310884 281802 310888 281858
rect 310888 281802 310944 281858
rect 310944 281802 310948 281858
rect 310884 281798 310948 281802
rect 310964 281858 311028 281862
rect 310964 281802 310968 281858
rect 310968 281802 311024 281858
rect 311024 281802 311028 281858
rect 310964 281798 311028 281802
rect 311044 281858 311108 281862
rect 311044 281802 311048 281858
rect 311048 281802 311104 281858
rect 311104 281802 311108 281858
rect 311044 281798 311108 281802
rect 311124 281858 311188 281862
rect 311124 281802 311128 281858
rect 311128 281802 311184 281858
rect 311184 281802 311188 281858
rect 311124 281798 311188 281802
rect 310884 281778 310948 281782
rect 310884 281722 310888 281778
rect 310888 281722 310944 281778
rect 310944 281722 310948 281778
rect 310884 281718 310948 281722
rect 310964 281778 311028 281782
rect 310964 281722 310968 281778
rect 310968 281722 311024 281778
rect 311024 281722 311028 281778
rect 310964 281718 311028 281722
rect 311044 281778 311108 281782
rect 311044 281722 311048 281778
rect 311048 281722 311104 281778
rect 311104 281722 311108 281778
rect 311044 281718 311108 281722
rect 311124 281778 311188 281782
rect 311124 281722 311128 281778
rect 311128 281722 311184 281778
rect 311184 281722 311188 281778
rect 311124 281718 311188 281722
rect 310884 281698 310948 281702
rect 310884 281642 310888 281698
rect 310888 281642 310944 281698
rect 310944 281642 310948 281698
rect 310884 281638 310948 281642
rect 310964 281698 311028 281702
rect 310964 281642 310968 281698
rect 310968 281642 311024 281698
rect 311024 281642 311028 281698
rect 310964 281638 311028 281642
rect 311044 281698 311108 281702
rect 311044 281642 311048 281698
rect 311048 281642 311104 281698
rect 311104 281642 311108 281698
rect 311044 281638 311108 281642
rect 311124 281698 311188 281702
rect 311124 281642 311128 281698
rect 311128 281642 311184 281698
rect 311184 281642 311188 281698
rect 311124 281638 311188 281642
rect 302152 261994 302216 261998
rect 302152 261938 302156 261994
rect 302156 261938 302212 261994
rect 302212 261938 302216 261994
rect 302152 261934 302216 261938
rect 302232 261994 302296 261998
rect 302232 261938 302236 261994
rect 302236 261938 302292 261994
rect 302292 261938 302296 261994
rect 302232 261934 302296 261938
rect 302312 261994 302376 261998
rect 302312 261938 302316 261994
rect 302316 261938 302372 261994
rect 302372 261938 302376 261994
rect 302312 261934 302376 261938
rect 302392 261994 302456 261998
rect 302392 261938 302396 261994
rect 302396 261938 302452 261994
rect 302452 261938 302456 261994
rect 302392 261934 302456 261938
rect 302152 261914 302216 261918
rect 302152 261858 302156 261914
rect 302156 261858 302212 261914
rect 302212 261858 302216 261914
rect 302152 261854 302216 261858
rect 302232 261914 302296 261918
rect 302232 261858 302236 261914
rect 302236 261858 302292 261914
rect 302292 261858 302296 261914
rect 302232 261854 302296 261858
rect 302312 261914 302376 261918
rect 302312 261858 302316 261914
rect 302316 261858 302372 261914
rect 302372 261858 302376 261914
rect 302312 261854 302376 261858
rect 302392 261914 302456 261918
rect 302392 261858 302396 261914
rect 302396 261858 302452 261914
rect 302452 261858 302456 261914
rect 302392 261854 302456 261858
rect 302152 261834 302216 261838
rect 302152 261778 302156 261834
rect 302156 261778 302212 261834
rect 302212 261778 302216 261834
rect 302152 261774 302216 261778
rect 302232 261834 302296 261838
rect 302232 261778 302236 261834
rect 302236 261778 302292 261834
rect 302292 261778 302296 261834
rect 302232 261774 302296 261778
rect 302312 261834 302376 261838
rect 302312 261778 302316 261834
rect 302316 261778 302372 261834
rect 302372 261778 302376 261834
rect 302312 261774 302376 261778
rect 302392 261834 302456 261838
rect 302392 261778 302396 261834
rect 302396 261778 302452 261834
rect 302452 261778 302456 261834
rect 302392 261774 302456 261778
rect 302152 261754 302216 261758
rect 302152 261698 302156 261754
rect 302156 261698 302212 261754
rect 302212 261698 302216 261754
rect 302152 261694 302216 261698
rect 302232 261754 302296 261758
rect 302232 261698 302236 261754
rect 302236 261698 302292 261754
rect 302292 261698 302296 261754
rect 302232 261694 302296 261698
rect 302312 261754 302376 261758
rect 302312 261698 302316 261754
rect 302316 261698 302372 261754
rect 302372 261698 302376 261754
rect 302312 261694 302376 261698
rect 302392 261754 302456 261758
rect 302392 261698 302396 261754
rect 302396 261698 302452 261754
rect 302452 261698 302456 261754
rect 302392 261694 302456 261698
rect 309152 261994 309216 261998
rect 309152 261938 309156 261994
rect 309156 261938 309212 261994
rect 309212 261938 309216 261994
rect 309152 261934 309216 261938
rect 309232 261994 309296 261998
rect 309232 261938 309236 261994
rect 309236 261938 309292 261994
rect 309292 261938 309296 261994
rect 309232 261934 309296 261938
rect 309312 261994 309376 261998
rect 309312 261938 309316 261994
rect 309316 261938 309372 261994
rect 309372 261938 309376 261994
rect 309312 261934 309376 261938
rect 309392 261994 309456 261998
rect 309392 261938 309396 261994
rect 309396 261938 309452 261994
rect 309452 261938 309456 261994
rect 309392 261934 309456 261938
rect 309152 261914 309216 261918
rect 309152 261858 309156 261914
rect 309156 261858 309212 261914
rect 309212 261858 309216 261914
rect 309152 261854 309216 261858
rect 309232 261914 309296 261918
rect 309232 261858 309236 261914
rect 309236 261858 309292 261914
rect 309292 261858 309296 261914
rect 309232 261854 309296 261858
rect 309312 261914 309376 261918
rect 309312 261858 309316 261914
rect 309316 261858 309372 261914
rect 309372 261858 309376 261914
rect 309312 261854 309376 261858
rect 309392 261914 309456 261918
rect 309392 261858 309396 261914
rect 309396 261858 309452 261914
rect 309452 261858 309456 261914
rect 309392 261854 309456 261858
rect 309152 261834 309216 261838
rect 309152 261778 309156 261834
rect 309156 261778 309212 261834
rect 309212 261778 309216 261834
rect 309152 261774 309216 261778
rect 309232 261834 309296 261838
rect 309232 261778 309236 261834
rect 309236 261778 309292 261834
rect 309292 261778 309296 261834
rect 309232 261774 309296 261778
rect 309312 261834 309376 261838
rect 309312 261778 309316 261834
rect 309316 261778 309372 261834
rect 309372 261778 309376 261834
rect 309312 261774 309376 261778
rect 309392 261834 309456 261838
rect 309392 261778 309396 261834
rect 309396 261778 309452 261834
rect 309452 261778 309456 261834
rect 309392 261774 309456 261778
rect 309152 261754 309216 261758
rect 309152 261698 309156 261754
rect 309156 261698 309212 261754
rect 309212 261698 309216 261754
rect 309152 261694 309216 261698
rect 309232 261754 309296 261758
rect 309232 261698 309236 261754
rect 309236 261698 309292 261754
rect 309292 261698 309296 261754
rect 309232 261694 309296 261698
rect 309312 261754 309376 261758
rect 309312 261698 309316 261754
rect 309316 261698 309372 261754
rect 309372 261698 309376 261754
rect 309312 261694 309376 261698
rect 309392 261754 309456 261758
rect 309392 261698 309396 261754
rect 309396 261698 309452 261754
rect 309452 261698 309456 261754
rect 309392 261694 309456 261698
rect 303884 261233 303948 261237
rect 303884 261177 303888 261233
rect 303888 261177 303944 261233
rect 303944 261177 303948 261233
rect 303884 261173 303948 261177
rect 303964 261233 304028 261237
rect 303964 261177 303968 261233
rect 303968 261177 304024 261233
rect 304024 261177 304028 261233
rect 303964 261173 304028 261177
rect 304044 261233 304108 261237
rect 304044 261177 304048 261233
rect 304048 261177 304104 261233
rect 304104 261177 304108 261233
rect 304044 261173 304108 261177
rect 304124 261233 304188 261237
rect 304124 261177 304128 261233
rect 304128 261177 304184 261233
rect 304184 261177 304188 261233
rect 304124 261173 304188 261177
rect 303884 261153 303948 261157
rect 303884 261097 303888 261153
rect 303888 261097 303944 261153
rect 303944 261097 303948 261153
rect 303884 261093 303948 261097
rect 303964 261153 304028 261157
rect 303964 261097 303968 261153
rect 303968 261097 304024 261153
rect 304024 261097 304028 261153
rect 303964 261093 304028 261097
rect 304044 261153 304108 261157
rect 304044 261097 304048 261153
rect 304048 261097 304104 261153
rect 304104 261097 304108 261153
rect 304044 261093 304108 261097
rect 304124 261153 304188 261157
rect 304124 261097 304128 261153
rect 304128 261097 304184 261153
rect 304184 261097 304188 261153
rect 304124 261093 304188 261097
rect 303884 261073 303948 261077
rect 303884 261017 303888 261073
rect 303888 261017 303944 261073
rect 303944 261017 303948 261073
rect 303884 261013 303948 261017
rect 303964 261073 304028 261077
rect 303964 261017 303968 261073
rect 303968 261017 304024 261073
rect 304024 261017 304028 261073
rect 303964 261013 304028 261017
rect 304044 261073 304108 261077
rect 304044 261017 304048 261073
rect 304048 261017 304104 261073
rect 304104 261017 304108 261073
rect 304044 261013 304108 261017
rect 304124 261073 304188 261077
rect 304124 261017 304128 261073
rect 304128 261017 304184 261073
rect 304184 261017 304188 261073
rect 304124 261013 304188 261017
rect 303884 260993 303948 260997
rect 303884 260937 303888 260993
rect 303888 260937 303944 260993
rect 303944 260937 303948 260993
rect 303884 260933 303948 260937
rect 303964 260993 304028 260997
rect 303964 260937 303968 260993
rect 303968 260937 304024 260993
rect 304024 260937 304028 260993
rect 303964 260933 304028 260937
rect 304044 260993 304108 260997
rect 304044 260937 304048 260993
rect 304048 260937 304104 260993
rect 304104 260937 304108 260993
rect 304044 260933 304108 260937
rect 304124 260993 304188 260997
rect 304124 260937 304128 260993
rect 304128 260937 304184 260993
rect 304184 260937 304188 260993
rect 304124 260933 304188 260937
rect 303884 260913 303948 260917
rect 303884 260857 303888 260913
rect 303888 260857 303944 260913
rect 303944 260857 303948 260913
rect 303884 260853 303948 260857
rect 303964 260913 304028 260917
rect 303964 260857 303968 260913
rect 303968 260857 304024 260913
rect 304024 260857 304028 260913
rect 303964 260853 304028 260857
rect 304044 260913 304108 260917
rect 304044 260857 304048 260913
rect 304048 260857 304104 260913
rect 304104 260857 304108 260913
rect 304044 260853 304108 260857
rect 304124 260913 304188 260917
rect 304124 260857 304128 260913
rect 304128 260857 304184 260913
rect 304184 260857 304188 260913
rect 304124 260853 304188 260857
rect 303884 260833 303948 260837
rect 303884 260777 303888 260833
rect 303888 260777 303944 260833
rect 303944 260777 303948 260833
rect 303884 260773 303948 260777
rect 303964 260833 304028 260837
rect 303964 260777 303968 260833
rect 303968 260777 304024 260833
rect 304024 260777 304028 260833
rect 303964 260773 304028 260777
rect 304044 260833 304108 260837
rect 304044 260777 304048 260833
rect 304048 260777 304104 260833
rect 304104 260777 304108 260833
rect 304044 260773 304108 260777
rect 304124 260833 304188 260837
rect 304124 260777 304128 260833
rect 304128 260777 304184 260833
rect 304184 260777 304188 260833
rect 304124 260773 304188 260777
rect 303884 260753 303948 260757
rect 303884 260697 303888 260753
rect 303888 260697 303944 260753
rect 303944 260697 303948 260753
rect 303884 260693 303948 260697
rect 303964 260753 304028 260757
rect 303964 260697 303968 260753
rect 303968 260697 304024 260753
rect 304024 260697 304028 260753
rect 303964 260693 304028 260697
rect 304044 260753 304108 260757
rect 304044 260697 304048 260753
rect 304048 260697 304104 260753
rect 304104 260697 304108 260753
rect 304044 260693 304108 260697
rect 304124 260753 304188 260757
rect 304124 260697 304128 260753
rect 304128 260697 304184 260753
rect 304184 260697 304188 260753
rect 304124 260693 304188 260697
rect 303884 260673 303948 260677
rect 303884 260617 303888 260673
rect 303888 260617 303944 260673
rect 303944 260617 303948 260673
rect 303884 260613 303948 260617
rect 303964 260673 304028 260677
rect 303964 260617 303968 260673
rect 303968 260617 304024 260673
rect 304024 260617 304028 260673
rect 303964 260613 304028 260617
rect 304044 260673 304108 260677
rect 304044 260617 304048 260673
rect 304048 260617 304104 260673
rect 304104 260617 304108 260673
rect 304044 260613 304108 260617
rect 304124 260673 304188 260677
rect 304124 260617 304128 260673
rect 304128 260617 304184 260673
rect 304184 260617 304188 260673
rect 304124 260613 304188 260617
rect 296884 242080 296948 242084
rect 296884 242024 296888 242080
rect 296888 242024 296944 242080
rect 296944 242024 296948 242080
rect 296884 242020 296948 242024
rect 296964 242080 297028 242084
rect 296964 242024 296968 242080
rect 296968 242024 297024 242080
rect 297024 242024 297028 242080
rect 296964 242020 297028 242024
rect 297044 242080 297108 242084
rect 297044 242024 297048 242080
rect 297048 242024 297104 242080
rect 297104 242024 297108 242080
rect 297044 242020 297108 242024
rect 297124 242080 297188 242084
rect 297124 242024 297128 242080
rect 297128 242024 297184 242080
rect 297184 242024 297188 242080
rect 297124 242020 297188 242024
rect 296884 242000 296948 242004
rect 296884 241944 296888 242000
rect 296888 241944 296944 242000
rect 296944 241944 296948 242000
rect 296884 241940 296948 241944
rect 296964 242000 297028 242004
rect 296964 241944 296968 242000
rect 296968 241944 297024 242000
rect 297024 241944 297028 242000
rect 296964 241940 297028 241944
rect 297044 242000 297108 242004
rect 297044 241944 297048 242000
rect 297048 241944 297104 242000
rect 297104 241944 297108 242000
rect 297044 241940 297108 241944
rect 297124 242000 297188 242004
rect 297124 241944 297128 242000
rect 297128 241944 297184 242000
rect 297184 241944 297188 242000
rect 297124 241940 297188 241944
rect 296884 241920 296948 241924
rect 296884 241864 296888 241920
rect 296888 241864 296944 241920
rect 296944 241864 296948 241920
rect 296884 241860 296948 241864
rect 296964 241920 297028 241924
rect 296964 241864 296968 241920
rect 296968 241864 297024 241920
rect 297024 241864 297028 241920
rect 296964 241860 297028 241864
rect 297044 241920 297108 241924
rect 297044 241864 297048 241920
rect 297048 241864 297104 241920
rect 297104 241864 297108 241920
rect 297044 241860 297108 241864
rect 297124 241920 297188 241924
rect 297124 241864 297128 241920
rect 297128 241864 297184 241920
rect 297184 241864 297188 241920
rect 297124 241860 297188 241864
rect 303884 242080 303948 242084
rect 303884 242024 303888 242080
rect 303888 242024 303944 242080
rect 303944 242024 303948 242080
rect 303884 242020 303948 242024
rect 303964 242080 304028 242084
rect 303964 242024 303968 242080
rect 303968 242024 304024 242080
rect 304024 242024 304028 242080
rect 303964 242020 304028 242024
rect 304044 242080 304108 242084
rect 304044 242024 304048 242080
rect 304048 242024 304104 242080
rect 304104 242024 304108 242080
rect 304044 242020 304108 242024
rect 304124 242080 304188 242084
rect 304124 242024 304128 242080
rect 304128 242024 304184 242080
rect 304184 242024 304188 242080
rect 304124 242020 304188 242024
rect 303884 242000 303948 242004
rect 303884 241944 303888 242000
rect 303888 241944 303944 242000
rect 303944 241944 303948 242000
rect 303884 241940 303948 241944
rect 303964 242000 304028 242004
rect 303964 241944 303968 242000
rect 303968 241944 304024 242000
rect 304024 241944 304028 242000
rect 303964 241940 304028 241944
rect 304044 242000 304108 242004
rect 304044 241944 304048 242000
rect 304048 241944 304104 242000
rect 304104 241944 304108 242000
rect 304044 241940 304108 241944
rect 304124 242000 304188 242004
rect 304124 241944 304128 242000
rect 304128 241944 304184 242000
rect 304184 241944 304188 242000
rect 304124 241940 304188 241944
rect 296884 241840 296948 241844
rect 296884 241784 296888 241840
rect 296888 241784 296944 241840
rect 296944 241784 296948 241840
rect 296884 241780 296948 241784
rect 296964 241840 297028 241844
rect 296964 241784 296968 241840
rect 296968 241784 297024 241840
rect 297024 241784 297028 241840
rect 296964 241780 297028 241784
rect 297044 241840 297108 241844
rect 297044 241784 297048 241840
rect 297048 241784 297104 241840
rect 297104 241784 297108 241840
rect 297044 241780 297108 241784
rect 297124 241840 297188 241844
rect 297124 241784 297128 241840
rect 297128 241784 297184 241840
rect 297184 241784 297188 241840
rect 297124 241780 297188 241784
rect 303884 241920 303948 241924
rect 303884 241864 303888 241920
rect 303888 241864 303944 241920
rect 303944 241864 303948 241920
rect 303884 241860 303948 241864
rect 303964 241920 304028 241924
rect 303964 241864 303968 241920
rect 303968 241864 304024 241920
rect 304024 241864 304028 241920
rect 303964 241860 304028 241864
rect 304044 241920 304108 241924
rect 304044 241864 304048 241920
rect 304048 241864 304104 241920
rect 304104 241864 304108 241920
rect 304044 241860 304108 241864
rect 304124 241920 304188 241924
rect 304124 241864 304128 241920
rect 304128 241864 304184 241920
rect 304184 241864 304188 241920
rect 304124 241860 304188 241864
rect 310884 242080 310948 242084
rect 310884 242024 310888 242080
rect 310888 242024 310944 242080
rect 310944 242024 310948 242080
rect 310884 242020 310948 242024
rect 310964 242080 311028 242084
rect 310964 242024 310968 242080
rect 310968 242024 311024 242080
rect 311024 242024 311028 242080
rect 310964 242020 311028 242024
rect 311044 242080 311108 242084
rect 311044 242024 311048 242080
rect 311048 242024 311104 242080
rect 311104 242024 311108 242080
rect 311044 242020 311108 242024
rect 311124 242080 311188 242084
rect 311124 242024 311128 242080
rect 311128 242024 311184 242080
rect 311184 242024 311188 242080
rect 311124 242020 311188 242024
rect 310884 242000 310948 242004
rect 310884 241944 310888 242000
rect 310888 241944 310944 242000
rect 310944 241944 310948 242000
rect 310884 241940 310948 241944
rect 310964 242000 311028 242004
rect 310964 241944 310968 242000
rect 310968 241944 311024 242000
rect 311024 241944 311028 242000
rect 310964 241940 311028 241944
rect 311044 242000 311108 242004
rect 311044 241944 311048 242000
rect 311048 241944 311104 242000
rect 311104 241944 311108 242000
rect 311044 241940 311108 241944
rect 311124 242000 311188 242004
rect 311124 241944 311128 242000
rect 311128 241944 311184 242000
rect 311184 241944 311188 242000
rect 311124 241940 311188 241944
rect 303884 241840 303948 241844
rect 303884 241784 303888 241840
rect 303888 241784 303944 241840
rect 303944 241784 303948 241840
rect 303884 241780 303948 241784
rect 303964 241840 304028 241844
rect 303964 241784 303968 241840
rect 303968 241784 304024 241840
rect 304024 241784 304028 241840
rect 303964 241780 304028 241784
rect 304044 241840 304108 241844
rect 304044 241784 304048 241840
rect 304048 241784 304104 241840
rect 304104 241784 304108 241840
rect 304044 241780 304108 241784
rect 304124 241840 304188 241844
rect 304124 241784 304128 241840
rect 304128 241784 304184 241840
rect 304184 241784 304188 241840
rect 304124 241780 304188 241784
rect 310884 241920 310948 241924
rect 310884 241864 310888 241920
rect 310888 241864 310944 241920
rect 310944 241864 310948 241920
rect 310884 241860 310948 241864
rect 310964 241920 311028 241924
rect 310964 241864 310968 241920
rect 310968 241864 311024 241920
rect 311024 241864 311028 241920
rect 310964 241860 311028 241864
rect 311044 241920 311108 241924
rect 311044 241864 311048 241920
rect 311048 241864 311104 241920
rect 311104 241864 311108 241920
rect 311044 241860 311108 241864
rect 311124 241920 311188 241924
rect 311124 241864 311128 241920
rect 311128 241864 311184 241920
rect 311184 241864 311188 241920
rect 311124 241860 311188 241864
rect 310884 241840 310948 241844
rect 310884 241784 310888 241840
rect 310888 241784 310944 241840
rect 310944 241784 310948 241840
rect 310884 241780 310948 241784
rect 310964 241840 311028 241844
rect 310964 241784 310968 241840
rect 310968 241784 311024 241840
rect 311024 241784 311028 241840
rect 310964 241780 311028 241784
rect 311044 241840 311108 241844
rect 311044 241784 311048 241840
rect 311048 241784 311104 241840
rect 311104 241784 311108 241840
rect 311044 241780 311108 241784
rect 311124 241840 311188 241844
rect 311124 241784 311128 241840
rect 311128 241784 311184 241840
rect 311184 241784 311188 241840
rect 311124 241780 311188 241784
rect 295152 240995 295216 240999
rect 295152 240939 295156 240995
rect 295156 240939 295212 240995
rect 295212 240939 295216 240995
rect 295152 240935 295216 240939
rect 295232 240995 295296 240999
rect 295232 240939 295236 240995
rect 295236 240939 295292 240995
rect 295292 240939 295296 240995
rect 295232 240935 295296 240939
rect 295312 240995 295376 240999
rect 295312 240939 295316 240995
rect 295316 240939 295372 240995
rect 295372 240939 295376 240995
rect 295312 240935 295376 240939
rect 295392 240995 295456 240999
rect 295392 240939 295396 240995
rect 295396 240939 295452 240995
rect 295452 240939 295456 240995
rect 295392 240935 295456 240939
rect 295152 240915 295216 240919
rect 295152 240859 295156 240915
rect 295156 240859 295212 240915
rect 295212 240859 295216 240915
rect 295152 240855 295216 240859
rect 295232 240915 295296 240919
rect 295232 240859 295236 240915
rect 295236 240859 295292 240915
rect 295292 240859 295296 240915
rect 295232 240855 295296 240859
rect 295312 240915 295376 240919
rect 295312 240859 295316 240915
rect 295316 240859 295372 240915
rect 295372 240859 295376 240915
rect 295312 240855 295376 240859
rect 295392 240915 295456 240919
rect 295392 240859 295396 240915
rect 295396 240859 295452 240915
rect 295452 240859 295456 240915
rect 295392 240855 295456 240859
rect 295152 240835 295216 240839
rect 295152 240779 295156 240835
rect 295156 240779 295212 240835
rect 295212 240779 295216 240835
rect 295152 240775 295216 240779
rect 295232 240835 295296 240839
rect 295232 240779 295236 240835
rect 295236 240779 295292 240835
rect 295292 240779 295296 240835
rect 295232 240775 295296 240779
rect 295312 240835 295376 240839
rect 295312 240779 295316 240835
rect 295316 240779 295372 240835
rect 295372 240779 295376 240835
rect 295312 240775 295376 240779
rect 295392 240835 295456 240839
rect 295392 240779 295396 240835
rect 295396 240779 295452 240835
rect 295452 240779 295456 240835
rect 295392 240775 295456 240779
rect 295152 240755 295216 240759
rect 295152 240699 295156 240755
rect 295156 240699 295212 240755
rect 295212 240699 295216 240755
rect 295152 240695 295216 240699
rect 295232 240755 295296 240759
rect 295232 240699 295236 240755
rect 295236 240699 295292 240755
rect 295292 240699 295296 240755
rect 295232 240695 295296 240699
rect 295312 240755 295376 240759
rect 295312 240699 295316 240755
rect 295316 240699 295372 240755
rect 295372 240699 295376 240755
rect 295312 240695 295376 240699
rect 295392 240755 295456 240759
rect 295392 240699 295396 240755
rect 295396 240699 295452 240755
rect 295452 240699 295456 240755
rect 295392 240695 295456 240699
rect 309152 240969 309216 240973
rect 309152 240913 309156 240969
rect 309156 240913 309212 240969
rect 309212 240913 309216 240969
rect 309152 240909 309216 240913
rect 309232 240969 309296 240973
rect 309232 240913 309236 240969
rect 309236 240913 309292 240969
rect 309292 240913 309296 240969
rect 309232 240909 309296 240913
rect 309312 240969 309376 240973
rect 309312 240913 309316 240969
rect 309316 240913 309372 240969
rect 309372 240913 309376 240969
rect 309312 240909 309376 240913
rect 309392 240969 309456 240973
rect 309392 240913 309396 240969
rect 309396 240913 309452 240969
rect 309452 240913 309456 240969
rect 309392 240909 309456 240913
rect 309152 240889 309216 240893
rect 309152 240833 309156 240889
rect 309156 240833 309212 240889
rect 309212 240833 309216 240889
rect 309152 240829 309216 240833
rect 309232 240889 309296 240893
rect 309232 240833 309236 240889
rect 309236 240833 309292 240889
rect 309292 240833 309296 240889
rect 309232 240829 309296 240833
rect 309312 240889 309376 240893
rect 309312 240833 309316 240889
rect 309316 240833 309372 240889
rect 309372 240833 309376 240889
rect 309312 240829 309376 240833
rect 309392 240889 309456 240893
rect 309392 240833 309396 240889
rect 309396 240833 309452 240889
rect 309452 240833 309456 240889
rect 309392 240829 309456 240833
rect 309152 240809 309216 240813
rect 309152 240753 309156 240809
rect 309156 240753 309212 240809
rect 309212 240753 309216 240809
rect 309152 240749 309216 240753
rect 309232 240809 309296 240813
rect 309232 240753 309236 240809
rect 309236 240753 309292 240809
rect 309292 240753 309296 240809
rect 309232 240749 309296 240753
rect 309312 240809 309376 240813
rect 309312 240753 309316 240809
rect 309316 240753 309372 240809
rect 309372 240753 309376 240809
rect 309312 240749 309376 240753
rect 309392 240809 309456 240813
rect 309392 240753 309396 240809
rect 309396 240753 309452 240809
rect 309452 240753 309456 240809
rect 309392 240749 309456 240753
rect 309152 240729 309216 240733
rect 309152 240673 309156 240729
rect 309156 240673 309212 240729
rect 309212 240673 309216 240729
rect 309152 240669 309216 240673
rect 309232 240729 309296 240733
rect 309232 240673 309236 240729
rect 309236 240673 309292 240729
rect 309292 240673 309296 240729
rect 309232 240669 309296 240673
rect 309312 240729 309376 240733
rect 309312 240673 309316 240729
rect 309316 240673 309372 240729
rect 309372 240673 309376 240729
rect 309312 240669 309376 240673
rect 309392 240729 309456 240733
rect 309392 240673 309396 240729
rect 309396 240673 309452 240729
rect 309452 240673 309456 240729
rect 309392 240669 309456 240673
rect 310884 239908 310948 239912
rect 310884 239852 310888 239908
rect 310888 239852 310944 239908
rect 310944 239852 310948 239908
rect 310884 239848 310948 239852
rect 310964 239908 311028 239912
rect 310964 239852 310968 239908
rect 310968 239852 311024 239908
rect 311024 239852 311028 239908
rect 310964 239848 311028 239852
rect 311044 239908 311108 239912
rect 311044 239852 311048 239908
rect 311048 239852 311104 239908
rect 311104 239852 311108 239908
rect 311044 239848 311108 239852
rect 311124 239908 311188 239912
rect 311124 239852 311128 239908
rect 311128 239852 311184 239908
rect 311184 239852 311188 239908
rect 311124 239848 311188 239852
rect 310884 239828 310948 239832
rect 310884 239772 310888 239828
rect 310888 239772 310944 239828
rect 310944 239772 310948 239828
rect 310884 239768 310948 239772
rect 310964 239828 311028 239832
rect 310964 239772 310968 239828
rect 310968 239772 311024 239828
rect 311024 239772 311028 239828
rect 310964 239768 311028 239772
rect 311044 239828 311108 239832
rect 311044 239772 311048 239828
rect 311048 239772 311104 239828
rect 311104 239772 311108 239828
rect 311044 239768 311108 239772
rect 311124 239828 311188 239832
rect 311124 239772 311128 239828
rect 311128 239772 311184 239828
rect 311184 239772 311188 239828
rect 311124 239768 311188 239772
rect 310884 239748 310948 239752
rect 310884 239692 310888 239748
rect 310888 239692 310944 239748
rect 310944 239692 310948 239748
rect 310884 239688 310948 239692
rect 310964 239748 311028 239752
rect 310964 239692 310968 239748
rect 310968 239692 311024 239748
rect 311024 239692 311028 239748
rect 310964 239688 311028 239692
rect 311044 239748 311108 239752
rect 311044 239692 311048 239748
rect 311048 239692 311104 239748
rect 311104 239692 311108 239748
rect 311044 239688 311108 239692
rect 311124 239748 311188 239752
rect 311124 239692 311128 239748
rect 311128 239692 311184 239748
rect 311184 239692 311188 239748
rect 311124 239688 311188 239692
rect 310884 239668 310948 239672
rect 310884 239612 310888 239668
rect 310888 239612 310944 239668
rect 310944 239612 310948 239668
rect 310884 239608 310948 239612
rect 310964 239668 311028 239672
rect 310964 239612 310968 239668
rect 310968 239612 311024 239668
rect 311024 239612 311028 239668
rect 310964 239608 311028 239612
rect 311044 239668 311108 239672
rect 311044 239612 311048 239668
rect 311048 239612 311104 239668
rect 311104 239612 311108 239668
rect 311044 239608 311108 239612
rect 311124 239668 311188 239672
rect 311124 239612 311128 239668
rect 311128 239612 311184 239668
rect 311184 239612 311188 239668
rect 311124 239608 311188 239612
rect 296884 221081 296948 221085
rect 296884 221025 296888 221081
rect 296888 221025 296944 221081
rect 296944 221025 296948 221081
rect 296884 221021 296948 221025
rect 296964 221081 297028 221085
rect 296964 221025 296968 221081
rect 296968 221025 297024 221081
rect 297024 221025 297028 221081
rect 296964 221021 297028 221025
rect 297044 221081 297108 221085
rect 297044 221025 297048 221081
rect 297048 221025 297104 221081
rect 297104 221025 297108 221081
rect 297044 221021 297108 221025
rect 297124 221081 297188 221085
rect 297124 221025 297128 221081
rect 297128 221025 297184 221081
rect 297184 221025 297188 221081
rect 297124 221021 297188 221025
rect 296884 221001 296948 221005
rect 296884 220945 296888 221001
rect 296888 220945 296944 221001
rect 296944 220945 296948 221001
rect 296884 220941 296948 220945
rect 296964 221001 297028 221005
rect 296964 220945 296968 221001
rect 296968 220945 297024 221001
rect 297024 220945 297028 221001
rect 296964 220941 297028 220945
rect 297044 221001 297108 221005
rect 297044 220945 297048 221001
rect 297048 220945 297104 221001
rect 297104 220945 297108 221001
rect 297044 220941 297108 220945
rect 297124 221001 297188 221005
rect 297124 220945 297128 221001
rect 297128 220945 297184 221001
rect 297184 220945 297188 221001
rect 297124 220941 297188 220945
rect 296884 220921 296948 220925
rect 296884 220865 296888 220921
rect 296888 220865 296944 220921
rect 296944 220865 296948 220921
rect 296884 220861 296948 220865
rect 296964 220921 297028 220925
rect 296964 220865 296968 220921
rect 296968 220865 297024 220921
rect 297024 220865 297028 220921
rect 296964 220861 297028 220865
rect 297044 220921 297108 220925
rect 297044 220865 297048 220921
rect 297048 220865 297104 220921
rect 297104 220865 297108 220921
rect 297044 220861 297108 220865
rect 297124 220921 297188 220925
rect 297124 220865 297128 220921
rect 297128 220865 297184 220921
rect 297184 220865 297188 220921
rect 297124 220861 297188 220865
rect 303884 221081 303948 221085
rect 303884 221025 303888 221081
rect 303888 221025 303944 221081
rect 303944 221025 303948 221081
rect 303884 221021 303948 221025
rect 303964 221081 304028 221085
rect 303964 221025 303968 221081
rect 303968 221025 304024 221081
rect 304024 221025 304028 221081
rect 303964 221021 304028 221025
rect 304044 221081 304108 221085
rect 304044 221025 304048 221081
rect 304048 221025 304104 221081
rect 304104 221025 304108 221081
rect 304044 221021 304108 221025
rect 304124 221081 304188 221085
rect 304124 221025 304128 221081
rect 304128 221025 304184 221081
rect 304184 221025 304188 221081
rect 304124 221021 304188 221025
rect 296884 220841 296948 220845
rect 296884 220785 296888 220841
rect 296888 220785 296944 220841
rect 296944 220785 296948 220841
rect 296884 220781 296948 220785
rect 296964 220841 297028 220845
rect 296964 220785 296968 220841
rect 296968 220785 297024 220841
rect 297024 220785 297028 220841
rect 296964 220781 297028 220785
rect 297044 220841 297108 220845
rect 297044 220785 297048 220841
rect 297048 220785 297104 220841
rect 297104 220785 297108 220841
rect 297044 220781 297108 220785
rect 297124 220841 297188 220845
rect 297124 220785 297128 220841
rect 297128 220785 297184 220841
rect 297184 220785 297188 220841
rect 297124 220781 297188 220785
rect 303884 221001 303948 221005
rect 303884 220945 303888 221001
rect 303888 220945 303944 221001
rect 303944 220945 303948 221001
rect 303884 220941 303948 220945
rect 303964 221001 304028 221005
rect 303964 220945 303968 221001
rect 303968 220945 304024 221001
rect 304024 220945 304028 221001
rect 303964 220941 304028 220945
rect 304044 221001 304108 221005
rect 304044 220945 304048 221001
rect 304048 220945 304104 221001
rect 304104 220945 304108 221001
rect 304044 220941 304108 220945
rect 304124 221001 304188 221005
rect 304124 220945 304128 221001
rect 304128 220945 304184 221001
rect 304184 220945 304188 221001
rect 304124 220941 304188 220945
rect 310884 221081 310948 221085
rect 310884 221025 310888 221081
rect 310888 221025 310944 221081
rect 310944 221025 310948 221081
rect 310884 221021 310948 221025
rect 310964 221081 311028 221085
rect 310964 221025 310968 221081
rect 310968 221025 311024 221081
rect 311024 221025 311028 221081
rect 310964 221021 311028 221025
rect 311044 221081 311108 221085
rect 311044 221025 311048 221081
rect 311048 221025 311104 221081
rect 311104 221025 311108 221081
rect 311044 221021 311108 221025
rect 311124 221081 311188 221085
rect 311124 221025 311128 221081
rect 311128 221025 311184 221081
rect 311184 221025 311188 221081
rect 311124 221021 311188 221025
rect 303884 220921 303948 220925
rect 303884 220865 303888 220921
rect 303888 220865 303944 220921
rect 303944 220865 303948 220921
rect 303884 220861 303948 220865
rect 303964 220921 304028 220925
rect 303964 220865 303968 220921
rect 303968 220865 304024 220921
rect 304024 220865 304028 220921
rect 303964 220861 304028 220865
rect 304044 220921 304108 220925
rect 304044 220865 304048 220921
rect 304048 220865 304104 220921
rect 304104 220865 304108 220921
rect 304044 220861 304108 220865
rect 304124 220921 304188 220925
rect 304124 220865 304128 220921
rect 304128 220865 304184 220921
rect 304184 220865 304188 220921
rect 304124 220861 304188 220865
rect 303884 220841 303948 220845
rect 303884 220785 303888 220841
rect 303888 220785 303944 220841
rect 303944 220785 303948 220841
rect 303884 220781 303948 220785
rect 303964 220841 304028 220845
rect 303964 220785 303968 220841
rect 303968 220785 304024 220841
rect 304024 220785 304028 220841
rect 303964 220781 304028 220785
rect 304044 220841 304108 220845
rect 304044 220785 304048 220841
rect 304048 220785 304104 220841
rect 304104 220785 304108 220841
rect 304044 220781 304108 220785
rect 304124 220841 304188 220845
rect 304124 220785 304128 220841
rect 304128 220785 304184 220841
rect 304184 220785 304188 220841
rect 304124 220781 304188 220785
rect 310884 221001 310948 221005
rect 310884 220945 310888 221001
rect 310888 220945 310944 221001
rect 310944 220945 310948 221001
rect 310884 220941 310948 220945
rect 310964 221001 311028 221005
rect 310964 220945 310968 221001
rect 310968 220945 311024 221001
rect 311024 220945 311028 221001
rect 310964 220941 311028 220945
rect 311044 221001 311108 221005
rect 311044 220945 311048 221001
rect 311048 220945 311104 221001
rect 311104 220945 311108 221001
rect 311044 220941 311108 220945
rect 311124 221001 311188 221005
rect 311124 220945 311128 221001
rect 311128 220945 311184 221001
rect 311184 220945 311188 221001
rect 311124 220941 311188 220945
rect 310884 220921 310948 220925
rect 310884 220865 310888 220921
rect 310888 220865 310944 220921
rect 310944 220865 310948 220921
rect 310884 220861 310948 220865
rect 310964 220921 311028 220925
rect 310964 220865 310968 220921
rect 310968 220865 311024 220921
rect 311024 220865 311028 220921
rect 310964 220861 311028 220865
rect 311044 220921 311108 220925
rect 311044 220865 311048 220921
rect 311048 220865 311104 220921
rect 311104 220865 311108 220921
rect 311044 220861 311108 220865
rect 311124 220921 311188 220925
rect 311124 220865 311128 220921
rect 311128 220865 311184 220921
rect 311184 220865 311188 220921
rect 311124 220861 311188 220865
rect 310884 220841 310948 220845
rect 310884 220785 310888 220841
rect 310888 220785 310944 220841
rect 310944 220785 310948 220841
rect 310884 220781 310948 220785
rect 310964 220841 311028 220845
rect 310964 220785 310968 220841
rect 310968 220785 311024 220841
rect 311024 220785 311028 220841
rect 310964 220781 311028 220785
rect 311044 220841 311108 220845
rect 311044 220785 311048 220841
rect 311048 220785 311104 220841
rect 311104 220785 311108 220841
rect 311044 220781 311108 220785
rect 311124 220841 311188 220845
rect 311124 220785 311128 220841
rect 311128 220785 311184 220841
rect 311184 220785 311188 220841
rect 311124 220781 311188 220785
rect 295152 219996 295216 220000
rect 295152 219940 295156 219996
rect 295156 219940 295212 219996
rect 295212 219940 295216 219996
rect 295152 219936 295216 219940
rect 295232 219996 295296 220000
rect 295232 219940 295236 219996
rect 295236 219940 295292 219996
rect 295292 219940 295296 219996
rect 295232 219936 295296 219940
rect 295312 219996 295376 220000
rect 295312 219940 295316 219996
rect 295316 219940 295372 219996
rect 295372 219940 295376 219996
rect 295312 219936 295376 219940
rect 295392 219996 295456 220000
rect 295392 219940 295396 219996
rect 295396 219940 295452 219996
rect 295452 219940 295456 219996
rect 295392 219936 295456 219940
rect 295152 219916 295216 219920
rect 295152 219860 295156 219916
rect 295156 219860 295212 219916
rect 295212 219860 295216 219916
rect 295152 219856 295216 219860
rect 295232 219916 295296 219920
rect 295232 219860 295236 219916
rect 295236 219860 295292 219916
rect 295292 219860 295296 219916
rect 295232 219856 295296 219860
rect 295312 219916 295376 219920
rect 295312 219860 295316 219916
rect 295316 219860 295372 219916
rect 295372 219860 295376 219916
rect 295312 219856 295376 219860
rect 295392 219916 295456 219920
rect 295392 219860 295396 219916
rect 295396 219860 295452 219916
rect 295452 219860 295456 219916
rect 295392 219856 295456 219860
rect 295152 219836 295216 219840
rect 295152 219780 295156 219836
rect 295156 219780 295212 219836
rect 295212 219780 295216 219836
rect 295152 219776 295216 219780
rect 295232 219836 295296 219840
rect 295232 219780 295236 219836
rect 295236 219780 295292 219836
rect 295292 219780 295296 219836
rect 295232 219776 295296 219780
rect 295312 219836 295376 219840
rect 295312 219780 295316 219836
rect 295316 219780 295372 219836
rect 295372 219780 295376 219836
rect 295312 219776 295376 219780
rect 295392 219836 295456 219840
rect 295392 219780 295396 219836
rect 295396 219780 295452 219836
rect 295452 219780 295456 219836
rect 295392 219776 295456 219780
rect 295152 219756 295216 219760
rect 295152 219700 295156 219756
rect 295156 219700 295212 219756
rect 295212 219700 295216 219756
rect 295152 219696 295216 219700
rect 295232 219756 295296 219760
rect 295232 219700 295236 219756
rect 295236 219700 295292 219756
rect 295292 219700 295296 219756
rect 295232 219696 295296 219700
rect 295312 219756 295376 219760
rect 295312 219700 295316 219756
rect 295316 219700 295372 219756
rect 295372 219700 295376 219756
rect 295312 219696 295376 219700
rect 295392 219756 295456 219760
rect 295392 219700 295396 219756
rect 295396 219700 295452 219756
rect 295452 219700 295456 219756
rect 295392 219696 295456 219700
rect 302152 219995 302216 219999
rect 302152 219939 302156 219995
rect 302156 219939 302212 219995
rect 302212 219939 302216 219995
rect 302152 219935 302216 219939
rect 302232 219995 302296 219999
rect 302232 219939 302236 219995
rect 302236 219939 302292 219995
rect 302292 219939 302296 219995
rect 302232 219935 302296 219939
rect 302312 219995 302376 219999
rect 302312 219939 302316 219995
rect 302316 219939 302372 219995
rect 302372 219939 302376 219995
rect 302312 219935 302376 219939
rect 302392 219995 302456 219999
rect 302392 219939 302396 219995
rect 302396 219939 302452 219995
rect 302452 219939 302456 219995
rect 302392 219935 302456 219939
rect 302152 219915 302216 219919
rect 302152 219859 302156 219915
rect 302156 219859 302212 219915
rect 302212 219859 302216 219915
rect 302152 219855 302216 219859
rect 302232 219915 302296 219919
rect 302232 219859 302236 219915
rect 302236 219859 302292 219915
rect 302292 219859 302296 219915
rect 302232 219855 302296 219859
rect 302312 219915 302376 219919
rect 302312 219859 302316 219915
rect 302316 219859 302372 219915
rect 302372 219859 302376 219915
rect 302312 219855 302376 219859
rect 302392 219915 302456 219919
rect 302392 219859 302396 219915
rect 302396 219859 302452 219915
rect 302452 219859 302456 219915
rect 302392 219855 302456 219859
rect 302152 219835 302216 219839
rect 302152 219779 302156 219835
rect 302156 219779 302212 219835
rect 302212 219779 302216 219835
rect 302152 219775 302216 219779
rect 302232 219835 302296 219839
rect 302232 219779 302236 219835
rect 302236 219779 302292 219835
rect 302292 219779 302296 219835
rect 302232 219775 302296 219779
rect 302312 219835 302376 219839
rect 302312 219779 302316 219835
rect 302316 219779 302372 219835
rect 302372 219779 302376 219835
rect 302312 219775 302376 219779
rect 302392 219835 302456 219839
rect 302392 219779 302396 219835
rect 302396 219779 302452 219835
rect 302452 219779 302456 219835
rect 302392 219775 302456 219779
rect 302152 219755 302216 219759
rect 302152 219699 302156 219755
rect 302156 219699 302212 219755
rect 302212 219699 302216 219755
rect 302152 219695 302216 219699
rect 302232 219755 302296 219759
rect 302232 219699 302236 219755
rect 302236 219699 302292 219755
rect 302292 219699 302296 219755
rect 302232 219695 302296 219699
rect 302312 219755 302376 219759
rect 302312 219699 302316 219755
rect 302316 219699 302372 219755
rect 302372 219699 302376 219755
rect 302312 219695 302376 219699
rect 302392 219755 302456 219759
rect 302392 219699 302396 219755
rect 302396 219699 302452 219755
rect 302452 219699 302456 219755
rect 302392 219695 302456 219699
rect 309152 219995 309216 219999
rect 309152 219939 309156 219995
rect 309156 219939 309212 219995
rect 309212 219939 309216 219995
rect 309152 219935 309216 219939
rect 309232 219995 309296 219999
rect 309232 219939 309236 219995
rect 309236 219939 309292 219995
rect 309292 219939 309296 219995
rect 309232 219935 309296 219939
rect 309312 219995 309376 219999
rect 309312 219939 309316 219995
rect 309316 219939 309372 219995
rect 309372 219939 309376 219995
rect 309312 219935 309376 219939
rect 309392 219995 309456 219999
rect 309392 219939 309396 219995
rect 309396 219939 309452 219995
rect 309452 219939 309456 219995
rect 309392 219935 309456 219939
rect 309152 219915 309216 219919
rect 309152 219859 309156 219915
rect 309156 219859 309212 219915
rect 309212 219859 309216 219915
rect 309152 219855 309216 219859
rect 309232 219915 309296 219919
rect 309232 219859 309236 219915
rect 309236 219859 309292 219915
rect 309292 219859 309296 219915
rect 309232 219855 309296 219859
rect 309312 219915 309376 219919
rect 309312 219859 309316 219915
rect 309316 219859 309372 219915
rect 309372 219859 309376 219915
rect 309312 219855 309376 219859
rect 309392 219915 309456 219919
rect 309392 219859 309396 219915
rect 309396 219859 309452 219915
rect 309452 219859 309456 219915
rect 309392 219855 309456 219859
rect 309152 219835 309216 219839
rect 309152 219779 309156 219835
rect 309156 219779 309212 219835
rect 309212 219779 309216 219835
rect 309152 219775 309216 219779
rect 309232 219835 309296 219839
rect 309232 219779 309236 219835
rect 309236 219779 309292 219835
rect 309292 219779 309296 219835
rect 309232 219775 309296 219779
rect 309312 219835 309376 219839
rect 309312 219779 309316 219835
rect 309316 219779 309372 219835
rect 309372 219779 309376 219835
rect 309312 219775 309376 219779
rect 309392 219835 309456 219839
rect 309392 219779 309396 219835
rect 309396 219779 309452 219835
rect 309452 219779 309456 219835
rect 309392 219775 309456 219779
rect 309152 219755 309216 219759
rect 309152 219699 309156 219755
rect 309156 219699 309212 219755
rect 309212 219699 309216 219755
rect 309152 219695 309216 219699
rect 309232 219755 309296 219759
rect 309232 219699 309236 219755
rect 309236 219699 309292 219755
rect 309292 219699 309296 219755
rect 309232 219695 309296 219699
rect 309312 219755 309376 219759
rect 309312 219699 309316 219755
rect 309316 219699 309372 219755
rect 309372 219699 309376 219755
rect 309312 219695 309376 219699
rect 309392 219755 309456 219759
rect 309392 219699 309396 219755
rect 309396 219699 309452 219755
rect 309452 219699 309456 219755
rect 309392 219695 309456 219699
rect 311039 219515 311103 219519
rect 311039 219459 311043 219515
rect 311043 219459 311099 219515
rect 311099 219459 311103 219515
rect 311039 219455 311103 219459
rect 303959 219398 304023 219402
rect 303959 219342 303963 219398
rect 303963 219342 304019 219398
rect 304019 219342 304023 219398
rect 303959 219338 304023 219342
rect 296884 179281 296948 179285
rect 296884 179225 296888 179281
rect 296888 179225 296944 179281
rect 296944 179225 296948 179281
rect 296884 179221 296948 179225
rect 296964 179281 297028 179285
rect 296964 179225 296968 179281
rect 296968 179225 297024 179281
rect 297024 179225 297028 179281
rect 296964 179221 297028 179225
rect 297044 179281 297108 179285
rect 297044 179225 297048 179281
rect 297048 179225 297104 179281
rect 297104 179225 297108 179281
rect 297044 179221 297108 179225
rect 297124 179281 297188 179285
rect 297124 179225 297128 179281
rect 297128 179225 297184 179281
rect 297184 179225 297188 179281
rect 297124 179221 297188 179225
rect 296884 179201 296948 179205
rect 296884 179145 296888 179201
rect 296888 179145 296944 179201
rect 296944 179145 296948 179201
rect 296884 179141 296948 179145
rect 296964 179201 297028 179205
rect 296964 179145 296968 179201
rect 296968 179145 297024 179201
rect 297024 179145 297028 179201
rect 296964 179141 297028 179145
rect 297044 179201 297108 179205
rect 297044 179145 297048 179201
rect 297048 179145 297104 179201
rect 297104 179145 297108 179201
rect 297044 179141 297108 179145
rect 297124 179201 297188 179205
rect 297124 179145 297128 179201
rect 297128 179145 297184 179201
rect 297184 179145 297188 179201
rect 297124 179141 297188 179145
rect 296884 179121 296948 179125
rect 296884 179065 296888 179121
rect 296888 179065 296944 179121
rect 296944 179065 296948 179121
rect 296884 179061 296948 179065
rect 296964 179121 297028 179125
rect 296964 179065 296968 179121
rect 296968 179065 297024 179121
rect 297024 179065 297028 179121
rect 296964 179061 297028 179065
rect 297044 179121 297108 179125
rect 297044 179065 297048 179121
rect 297048 179065 297104 179121
rect 297104 179065 297108 179121
rect 297044 179061 297108 179065
rect 297124 179121 297188 179125
rect 297124 179065 297128 179121
rect 297128 179065 297184 179121
rect 297184 179065 297188 179121
rect 297124 179061 297188 179065
rect 303884 179281 303948 179285
rect 303884 179225 303888 179281
rect 303888 179225 303944 179281
rect 303944 179225 303948 179281
rect 303884 179221 303948 179225
rect 303964 179281 304028 179285
rect 303964 179225 303968 179281
rect 303968 179225 304024 179281
rect 304024 179225 304028 179281
rect 303964 179221 304028 179225
rect 304044 179281 304108 179285
rect 304044 179225 304048 179281
rect 304048 179225 304104 179281
rect 304104 179225 304108 179281
rect 304044 179221 304108 179225
rect 304124 179281 304188 179285
rect 304124 179225 304128 179281
rect 304128 179225 304184 179281
rect 304184 179225 304188 179281
rect 304124 179221 304188 179225
rect 303884 179201 303948 179205
rect 303884 179145 303888 179201
rect 303888 179145 303944 179201
rect 303944 179145 303948 179201
rect 303884 179141 303948 179145
rect 303964 179201 304028 179205
rect 303964 179145 303968 179201
rect 303968 179145 304024 179201
rect 304024 179145 304028 179201
rect 303964 179141 304028 179145
rect 304044 179201 304108 179205
rect 304044 179145 304048 179201
rect 304048 179145 304104 179201
rect 304104 179145 304108 179201
rect 304044 179141 304108 179145
rect 304124 179201 304188 179205
rect 304124 179145 304128 179201
rect 304128 179145 304184 179201
rect 304184 179145 304188 179201
rect 304124 179141 304188 179145
rect 296884 179041 296948 179045
rect 296884 178985 296888 179041
rect 296888 178985 296944 179041
rect 296944 178985 296948 179041
rect 296884 178981 296948 178985
rect 296964 179041 297028 179045
rect 296964 178985 296968 179041
rect 296968 178985 297024 179041
rect 297024 178985 297028 179041
rect 296964 178981 297028 178985
rect 297044 179041 297108 179045
rect 297044 178985 297048 179041
rect 297048 178985 297104 179041
rect 297104 178985 297108 179041
rect 297044 178981 297108 178985
rect 297124 179041 297188 179045
rect 297124 178985 297128 179041
rect 297128 178985 297184 179041
rect 297184 178985 297188 179041
rect 297124 178981 297188 178985
rect 303884 179121 303948 179125
rect 303884 179065 303888 179121
rect 303888 179065 303944 179121
rect 303944 179065 303948 179121
rect 303884 179061 303948 179065
rect 303964 179121 304028 179125
rect 303964 179065 303968 179121
rect 303968 179065 304024 179121
rect 304024 179065 304028 179121
rect 303964 179061 304028 179065
rect 304044 179121 304108 179125
rect 304044 179065 304048 179121
rect 304048 179065 304104 179121
rect 304104 179065 304108 179121
rect 304044 179061 304108 179065
rect 304124 179121 304188 179125
rect 304124 179065 304128 179121
rect 304128 179065 304184 179121
rect 304184 179065 304188 179121
rect 304124 179061 304188 179065
rect 303884 179041 303948 179045
rect 303884 178985 303888 179041
rect 303888 178985 303944 179041
rect 303944 178985 303948 179041
rect 303884 178981 303948 178985
rect 303964 179041 304028 179045
rect 303964 178985 303968 179041
rect 303968 178985 304024 179041
rect 304024 178985 304028 179041
rect 303964 178981 304028 178985
rect 304044 179041 304108 179045
rect 304044 178985 304048 179041
rect 304048 178985 304104 179041
rect 304104 178985 304108 179041
rect 304044 178981 304108 178985
rect 304124 179041 304188 179045
rect 304124 178985 304128 179041
rect 304128 178985 304184 179041
rect 304184 178985 304188 179041
rect 304124 178981 304188 178985
rect 310888 179281 310952 179285
rect 310888 179225 310892 179281
rect 310892 179225 310948 179281
rect 310948 179225 310952 179281
rect 310888 179221 310952 179225
rect 310888 179201 310952 179205
rect 310888 179145 310892 179201
rect 310892 179145 310948 179201
rect 310948 179145 310952 179201
rect 310888 179141 310952 179145
rect 310888 179121 310952 179125
rect 310888 179065 310892 179121
rect 310892 179065 310948 179121
rect 310948 179065 310952 179121
rect 310888 179061 310952 179065
rect 310888 179041 310952 179045
rect 310888 178985 310892 179041
rect 310892 178985 310948 179041
rect 310948 178985 310952 179041
rect 310888 178981 310952 178985
rect 295152 178195 295216 178199
rect 295152 178139 295156 178195
rect 295156 178139 295212 178195
rect 295212 178139 295216 178195
rect 295152 178135 295216 178139
rect 295232 178195 295296 178199
rect 295232 178139 295236 178195
rect 295236 178139 295292 178195
rect 295292 178139 295296 178195
rect 295232 178135 295296 178139
rect 295312 178195 295376 178199
rect 295312 178139 295316 178195
rect 295316 178139 295372 178195
rect 295372 178139 295376 178195
rect 295312 178135 295376 178139
rect 295392 178195 295456 178199
rect 295392 178139 295396 178195
rect 295396 178139 295452 178195
rect 295452 178139 295456 178195
rect 295392 178135 295456 178139
rect 295152 178115 295216 178119
rect 295152 178059 295156 178115
rect 295156 178059 295212 178115
rect 295212 178059 295216 178115
rect 295152 178055 295216 178059
rect 295232 178115 295296 178119
rect 295232 178059 295236 178115
rect 295236 178059 295292 178115
rect 295292 178059 295296 178115
rect 295232 178055 295296 178059
rect 295312 178115 295376 178119
rect 295312 178059 295316 178115
rect 295316 178059 295372 178115
rect 295372 178059 295376 178115
rect 295312 178055 295376 178059
rect 295392 178115 295456 178119
rect 295392 178059 295396 178115
rect 295396 178059 295452 178115
rect 295452 178059 295456 178115
rect 295392 178055 295456 178059
rect 295152 178035 295216 178039
rect 295152 177979 295156 178035
rect 295156 177979 295212 178035
rect 295212 177979 295216 178035
rect 295152 177975 295216 177979
rect 295232 178035 295296 178039
rect 295232 177979 295236 178035
rect 295236 177979 295292 178035
rect 295292 177979 295296 178035
rect 295232 177975 295296 177979
rect 295312 178035 295376 178039
rect 295312 177979 295316 178035
rect 295316 177979 295372 178035
rect 295372 177979 295376 178035
rect 295312 177975 295376 177979
rect 295392 178035 295456 178039
rect 295392 177979 295396 178035
rect 295396 177979 295452 178035
rect 295452 177979 295456 178035
rect 295392 177975 295456 177979
rect 295152 177955 295216 177959
rect 295152 177899 295156 177955
rect 295156 177899 295212 177955
rect 295212 177899 295216 177955
rect 295152 177895 295216 177899
rect 295232 177955 295296 177959
rect 295232 177899 295236 177955
rect 295236 177899 295292 177955
rect 295292 177899 295296 177955
rect 295232 177895 295296 177899
rect 295312 177955 295376 177959
rect 295312 177899 295316 177955
rect 295316 177899 295372 177955
rect 295372 177899 295376 177955
rect 295312 177895 295376 177899
rect 295392 177955 295456 177959
rect 295392 177899 295396 177955
rect 295396 177899 295452 177955
rect 295452 177899 295456 177955
rect 295392 177895 295456 177899
rect 302152 178179 302216 178183
rect 302152 178123 302156 178179
rect 302156 178123 302212 178179
rect 302212 178123 302216 178179
rect 302152 178119 302216 178123
rect 302232 178179 302296 178183
rect 302232 178123 302236 178179
rect 302236 178123 302292 178179
rect 302292 178123 302296 178179
rect 302232 178119 302296 178123
rect 302312 178179 302376 178183
rect 302312 178123 302316 178179
rect 302316 178123 302372 178179
rect 302372 178123 302376 178179
rect 302312 178119 302376 178123
rect 302392 178179 302456 178183
rect 302392 178123 302396 178179
rect 302396 178123 302452 178179
rect 302452 178123 302456 178179
rect 302392 178119 302456 178123
rect 302152 178099 302216 178103
rect 302152 178043 302156 178099
rect 302156 178043 302212 178099
rect 302212 178043 302216 178099
rect 302152 178039 302216 178043
rect 302232 178099 302296 178103
rect 302232 178043 302236 178099
rect 302236 178043 302292 178099
rect 302292 178043 302296 178099
rect 302232 178039 302296 178043
rect 302312 178099 302376 178103
rect 302312 178043 302316 178099
rect 302316 178043 302372 178099
rect 302372 178043 302376 178099
rect 302312 178039 302376 178043
rect 302392 178099 302456 178103
rect 302392 178043 302396 178099
rect 302396 178043 302452 178099
rect 302452 178043 302456 178099
rect 302392 178039 302456 178043
rect 302152 178019 302216 178023
rect 302152 177963 302156 178019
rect 302156 177963 302212 178019
rect 302212 177963 302216 178019
rect 302152 177959 302216 177963
rect 302232 178019 302296 178023
rect 302232 177963 302236 178019
rect 302236 177963 302292 178019
rect 302292 177963 302296 178019
rect 302232 177959 302296 177963
rect 302312 178019 302376 178023
rect 302312 177963 302316 178019
rect 302316 177963 302372 178019
rect 302372 177963 302376 178019
rect 302312 177959 302376 177963
rect 302392 178019 302456 178023
rect 302392 177963 302396 178019
rect 302396 177963 302452 178019
rect 302452 177963 302456 178019
rect 302392 177959 302456 177963
rect 302152 177939 302216 177943
rect 302152 177883 302156 177939
rect 302156 177883 302212 177939
rect 302212 177883 302216 177939
rect 302152 177879 302216 177883
rect 302232 177939 302296 177943
rect 302232 177883 302236 177939
rect 302236 177883 302292 177939
rect 302292 177883 302296 177939
rect 302232 177879 302296 177883
rect 302312 177939 302376 177943
rect 302312 177883 302316 177939
rect 302316 177883 302372 177939
rect 302372 177883 302376 177939
rect 302312 177879 302376 177883
rect 302392 177939 302456 177943
rect 302392 177883 302396 177939
rect 302396 177883 302452 177939
rect 302452 177883 302456 177939
rect 302392 177879 302456 177883
rect 309152 178179 309216 178183
rect 309152 178123 309156 178179
rect 309156 178123 309212 178179
rect 309212 178123 309216 178179
rect 309152 178119 309216 178123
rect 309232 178179 309296 178183
rect 309232 178123 309236 178179
rect 309236 178123 309292 178179
rect 309292 178123 309296 178179
rect 309232 178119 309296 178123
rect 309312 178179 309376 178183
rect 309312 178123 309316 178179
rect 309316 178123 309372 178179
rect 309372 178123 309376 178179
rect 309312 178119 309376 178123
rect 309392 178179 309456 178183
rect 309392 178123 309396 178179
rect 309396 178123 309452 178179
rect 309452 178123 309456 178179
rect 309392 178119 309456 178123
rect 309152 178099 309216 178103
rect 309152 178043 309156 178099
rect 309156 178043 309212 178099
rect 309212 178043 309216 178099
rect 309152 178039 309216 178043
rect 309232 178099 309296 178103
rect 309232 178043 309236 178099
rect 309236 178043 309292 178099
rect 309292 178043 309296 178099
rect 309232 178039 309296 178043
rect 309312 178099 309376 178103
rect 309312 178043 309316 178099
rect 309316 178043 309372 178099
rect 309372 178043 309376 178099
rect 309312 178039 309376 178043
rect 309392 178099 309456 178103
rect 309392 178043 309396 178099
rect 309396 178043 309452 178099
rect 309452 178043 309456 178099
rect 309392 178039 309456 178043
rect 309152 178019 309216 178023
rect 309152 177963 309156 178019
rect 309156 177963 309212 178019
rect 309212 177963 309216 178019
rect 309152 177959 309216 177963
rect 309232 178019 309296 178023
rect 309232 177963 309236 178019
rect 309236 177963 309292 178019
rect 309292 177963 309296 178019
rect 309232 177959 309296 177963
rect 309312 178019 309376 178023
rect 309312 177963 309316 178019
rect 309316 177963 309372 178019
rect 309372 177963 309376 178019
rect 309312 177959 309376 177963
rect 309392 178019 309456 178023
rect 309392 177963 309396 178019
rect 309396 177963 309452 178019
rect 309452 177963 309456 178019
rect 309392 177959 309456 177963
rect 309152 177939 309216 177943
rect 309152 177883 309156 177939
rect 309156 177883 309212 177939
rect 309212 177883 309216 177939
rect 309152 177879 309216 177883
rect 309232 177939 309296 177943
rect 309232 177883 309236 177939
rect 309236 177883 309292 177939
rect 309292 177883 309296 177939
rect 309232 177879 309296 177883
rect 309312 177939 309376 177943
rect 309312 177883 309316 177939
rect 309316 177883 309372 177939
rect 309372 177883 309376 177939
rect 309312 177879 309376 177883
rect 309392 177939 309456 177943
rect 309392 177883 309396 177939
rect 309396 177883 309452 177939
rect 309452 177883 309456 177939
rect 309392 177879 309456 177883
<< metal4 >>
rect -4950 696561 -3538 707814
rect -4950 696325 -4842 696561
rect -4606 696325 -4522 696561
rect -4286 696325 -4202 696561
rect -3966 696325 -3882 696561
rect -3646 696325 -3538 696561
rect -4950 689561 -3538 696325
rect -4950 689325 -4842 689561
rect -4606 689325 -4522 689561
rect -4286 689325 -4202 689561
rect -3966 689325 -3882 689561
rect -3646 689325 -3538 689561
rect -4950 682561 -3538 689325
rect -4950 682325 -4842 682561
rect -4606 682325 -4522 682561
rect -4286 682325 -4202 682561
rect -3966 682325 -3882 682561
rect -3646 682325 -3538 682561
rect -4950 675561 -3538 682325
rect -4950 675325 -4842 675561
rect -4606 675325 -4522 675561
rect -4286 675325 -4202 675561
rect -3966 675325 -3882 675561
rect -3646 675325 -3538 675561
rect -4950 668561 -3538 675325
rect -4950 668325 -4842 668561
rect -4606 668325 -4522 668561
rect -4286 668325 -4202 668561
rect -3966 668325 -3882 668561
rect -3646 668325 -3538 668561
rect -4950 661561 -3538 668325
rect -4950 661325 -4842 661561
rect -4606 661325 -4522 661561
rect -4286 661325 -4202 661561
rect -3966 661325 -3882 661561
rect -3646 661325 -3538 661561
rect -4950 654561 -3538 661325
rect -4950 654325 -4842 654561
rect -4606 654325 -4522 654561
rect -4286 654325 -4202 654561
rect -3966 654325 -3882 654561
rect -3646 654325 -3538 654561
rect -4950 647561 -3538 654325
rect -4950 647325 -4842 647561
rect -4606 647325 -4522 647561
rect -4286 647325 -4202 647561
rect -3966 647325 -3882 647561
rect -3646 647325 -3538 647561
rect -4950 640561 -3538 647325
rect -4950 640325 -4842 640561
rect -4606 640325 -4522 640561
rect -4286 640325 -4202 640561
rect -3966 640325 -3882 640561
rect -3646 640325 -3538 640561
rect -4950 633561 -3538 640325
rect -4950 633325 -4842 633561
rect -4606 633325 -4522 633561
rect -4286 633325 -4202 633561
rect -3966 633325 -3882 633561
rect -3646 633325 -3538 633561
rect -4950 626561 -3538 633325
rect -4950 626325 -4842 626561
rect -4606 626325 -4522 626561
rect -4286 626325 -4202 626561
rect -3966 626325 -3882 626561
rect -3646 626325 -3538 626561
rect -4950 619561 -3538 626325
rect -4950 619325 -4842 619561
rect -4606 619325 -4522 619561
rect -4286 619325 -4202 619561
rect -3966 619325 -3882 619561
rect -3646 619325 -3538 619561
rect -4950 612561 -3538 619325
rect -4950 612325 -4842 612561
rect -4606 612325 -4522 612561
rect -4286 612325 -4202 612561
rect -3966 612325 -3882 612561
rect -3646 612325 -3538 612561
rect -4950 605561 -3538 612325
rect -4950 605325 -4842 605561
rect -4606 605325 -4522 605561
rect -4286 605325 -4202 605561
rect -3966 605325 -3882 605561
rect -3646 605325 -3538 605561
rect -4950 598561 -3538 605325
rect -4950 598325 -4842 598561
rect -4606 598325 -4522 598561
rect -4286 598325 -4202 598561
rect -3966 598325 -3882 598561
rect -3646 598325 -3538 598561
rect -4950 591561 -3538 598325
rect -4950 591325 -4842 591561
rect -4606 591325 -4522 591561
rect -4286 591325 -4202 591561
rect -3966 591325 -3882 591561
rect -3646 591325 -3538 591561
rect -4950 584561 -3538 591325
rect -4950 584325 -4842 584561
rect -4606 584325 -4522 584561
rect -4286 584325 -4202 584561
rect -3966 584325 -3882 584561
rect -3646 584325 -3538 584561
rect -4950 577561 -3538 584325
rect -4950 577325 -4842 577561
rect -4606 577325 -4522 577561
rect -4286 577325 -4202 577561
rect -3966 577325 -3882 577561
rect -3646 577325 -3538 577561
rect -4950 570561 -3538 577325
rect -4950 570325 -4842 570561
rect -4606 570325 -4522 570561
rect -4286 570325 -4202 570561
rect -3966 570325 -3882 570561
rect -3646 570325 -3538 570561
rect -4950 563561 -3538 570325
rect -4950 563325 -4842 563561
rect -4606 563325 -4522 563561
rect -4286 563325 -4202 563561
rect -3966 563325 -3882 563561
rect -3646 563325 -3538 563561
rect -4950 556561 -3538 563325
rect -4950 556325 -4842 556561
rect -4606 556325 -4522 556561
rect -4286 556325 -4202 556561
rect -3966 556325 -3882 556561
rect -3646 556325 -3538 556561
rect -4950 549561 -3538 556325
rect -4950 549325 -4842 549561
rect -4606 549325 -4522 549561
rect -4286 549325 -4202 549561
rect -3966 549325 -3882 549561
rect -3646 549325 -3538 549561
rect -4950 542561 -3538 549325
rect -4950 542325 -4842 542561
rect -4606 542325 -4522 542561
rect -4286 542325 -4202 542561
rect -3966 542325 -3882 542561
rect -3646 542325 -3538 542561
rect -4950 535561 -3538 542325
rect -4950 535325 -4842 535561
rect -4606 535325 -4522 535561
rect -4286 535325 -4202 535561
rect -3966 535325 -3882 535561
rect -3646 535325 -3538 535561
rect -4950 528561 -3538 535325
rect -4950 528325 -4842 528561
rect -4606 528325 -4522 528561
rect -4286 528325 -4202 528561
rect -3966 528325 -3882 528561
rect -3646 528325 -3538 528561
rect -4950 521561 -3538 528325
rect -4950 521325 -4842 521561
rect -4606 521325 -4522 521561
rect -4286 521325 -4202 521561
rect -3966 521325 -3882 521561
rect -3646 521325 -3538 521561
rect -4950 514561 -3538 521325
rect -4950 514325 -4842 514561
rect -4606 514325 -4522 514561
rect -4286 514325 -4202 514561
rect -3966 514325 -3882 514561
rect -3646 514325 -3538 514561
rect -4950 507561 -3538 514325
rect -4950 507325 -4842 507561
rect -4606 507325 -4522 507561
rect -4286 507325 -4202 507561
rect -3966 507325 -3882 507561
rect -3646 507325 -3538 507561
rect -4950 500561 -3538 507325
rect -4950 500325 -4842 500561
rect -4606 500325 -4522 500561
rect -4286 500325 -4202 500561
rect -3966 500325 -3882 500561
rect -3646 500325 -3538 500561
rect -4950 493561 -3538 500325
rect -4950 493325 -4842 493561
rect -4606 493325 -4522 493561
rect -4286 493325 -4202 493561
rect -3966 493325 -3882 493561
rect -3646 493325 -3538 493561
rect -4950 486561 -3538 493325
rect -4950 486325 -4842 486561
rect -4606 486325 -4522 486561
rect -4286 486325 -4202 486561
rect -3966 486325 -3882 486561
rect -3646 486325 -3538 486561
rect -4950 479561 -3538 486325
rect -4950 479325 -4842 479561
rect -4606 479325 -4522 479561
rect -4286 479325 -4202 479561
rect -3966 479325 -3882 479561
rect -3646 479325 -3538 479561
rect -4950 472561 -3538 479325
rect -4950 472325 -4842 472561
rect -4606 472325 -4522 472561
rect -4286 472325 -4202 472561
rect -3966 472325 -3882 472561
rect -3646 472325 -3538 472561
rect -4950 465561 -3538 472325
rect -4950 465325 -4842 465561
rect -4606 465325 -4522 465561
rect -4286 465325 -4202 465561
rect -3966 465325 -3882 465561
rect -3646 465325 -3538 465561
rect -4950 458561 -3538 465325
rect -4950 458325 -4842 458561
rect -4606 458325 -4522 458561
rect -4286 458325 -4202 458561
rect -3966 458325 -3882 458561
rect -3646 458325 -3538 458561
rect -4950 451561 -3538 458325
rect -4950 451325 -4842 451561
rect -4606 451325 -4522 451561
rect -4286 451325 -4202 451561
rect -3966 451325 -3882 451561
rect -3646 451325 -3538 451561
rect -4950 444561 -3538 451325
rect -4950 444325 -4842 444561
rect -4606 444325 -4522 444561
rect -4286 444325 -4202 444561
rect -3966 444325 -3882 444561
rect -3646 444325 -3538 444561
rect -4950 437561 -3538 444325
rect -4950 437325 -4842 437561
rect -4606 437325 -4522 437561
rect -4286 437325 -4202 437561
rect -3966 437325 -3882 437561
rect -3646 437325 -3538 437561
rect -4950 430561 -3538 437325
rect -4950 430325 -4842 430561
rect -4606 430325 -4522 430561
rect -4286 430325 -4202 430561
rect -3966 430325 -3882 430561
rect -3646 430325 -3538 430561
rect -4950 423561 -3538 430325
rect -4950 423325 -4842 423561
rect -4606 423325 -4522 423561
rect -4286 423325 -4202 423561
rect -3966 423325 -3882 423561
rect -3646 423325 -3538 423561
rect -4950 416561 -3538 423325
rect -4950 416325 -4842 416561
rect -4606 416325 -4522 416561
rect -4286 416325 -4202 416561
rect -3966 416325 -3882 416561
rect -3646 416325 -3538 416561
rect -4950 409561 -3538 416325
rect -4950 409325 -4842 409561
rect -4606 409325 -4522 409561
rect -4286 409325 -4202 409561
rect -3966 409325 -3882 409561
rect -3646 409325 -3538 409561
rect -4950 402561 -3538 409325
rect -4950 402325 -4842 402561
rect -4606 402325 -4522 402561
rect -4286 402325 -4202 402561
rect -3966 402325 -3882 402561
rect -3646 402325 -3538 402561
rect -4950 395561 -3538 402325
rect -4950 395325 -4842 395561
rect -4606 395325 -4522 395561
rect -4286 395325 -4202 395561
rect -3966 395325 -3882 395561
rect -3646 395325 -3538 395561
rect -4950 388561 -3538 395325
rect -4950 388325 -4842 388561
rect -4606 388325 -4522 388561
rect -4286 388325 -4202 388561
rect -3966 388325 -3882 388561
rect -3646 388325 -3538 388561
rect -4950 381561 -3538 388325
rect -4950 381325 -4842 381561
rect -4606 381325 -4522 381561
rect -4286 381325 -4202 381561
rect -3966 381325 -3882 381561
rect -3646 381325 -3538 381561
rect -4950 374561 -3538 381325
rect -4950 374325 -4842 374561
rect -4606 374325 -4522 374561
rect -4286 374325 -4202 374561
rect -3966 374325 -3882 374561
rect -3646 374325 -3538 374561
rect -4950 367561 -3538 374325
rect -4950 367325 -4842 367561
rect -4606 367325 -4522 367561
rect -4286 367325 -4202 367561
rect -3966 367325 -3882 367561
rect -3646 367325 -3538 367561
rect -4950 360561 -3538 367325
rect -4950 360325 -4842 360561
rect -4606 360325 -4522 360561
rect -4286 360325 -4202 360561
rect -3966 360325 -3882 360561
rect -3646 360325 -3538 360561
rect -4950 353561 -3538 360325
rect -4950 353325 -4842 353561
rect -4606 353325 -4522 353561
rect -4286 353325 -4202 353561
rect -3966 353325 -3882 353561
rect -3646 353325 -3538 353561
rect -4950 346561 -3538 353325
rect -4950 346325 -4842 346561
rect -4606 346325 -4522 346561
rect -4286 346325 -4202 346561
rect -3966 346325 -3882 346561
rect -3646 346325 -3538 346561
rect -4950 339561 -3538 346325
rect -4950 339325 -4842 339561
rect -4606 339325 -4522 339561
rect -4286 339325 -4202 339561
rect -3966 339325 -3882 339561
rect -3646 339325 -3538 339561
rect -4950 332561 -3538 339325
rect -4950 332325 -4842 332561
rect -4606 332325 -4522 332561
rect -4286 332325 -4202 332561
rect -3966 332325 -3882 332561
rect -3646 332325 -3538 332561
rect -4950 325561 -3538 332325
rect -4950 325325 -4842 325561
rect -4606 325325 -4522 325561
rect -4286 325325 -4202 325561
rect -3966 325325 -3882 325561
rect -3646 325325 -3538 325561
rect -4950 318561 -3538 325325
rect -4950 318325 -4842 318561
rect -4606 318325 -4522 318561
rect -4286 318325 -4202 318561
rect -3966 318325 -3882 318561
rect -3646 318325 -3538 318561
rect -4950 311561 -3538 318325
rect -4950 311325 -4842 311561
rect -4606 311325 -4522 311561
rect -4286 311325 -4202 311561
rect -3966 311325 -3882 311561
rect -3646 311325 -3538 311561
rect -4950 304561 -3538 311325
rect -4950 304325 -4842 304561
rect -4606 304325 -4522 304561
rect -4286 304325 -4202 304561
rect -3966 304325 -3882 304561
rect -3646 304325 -3538 304561
rect -4950 297561 -3538 304325
rect -4950 297325 -4842 297561
rect -4606 297325 -4522 297561
rect -4286 297325 -4202 297561
rect -3966 297325 -3882 297561
rect -3646 297325 -3538 297561
rect -4950 290561 -3538 297325
rect -4950 290325 -4842 290561
rect -4606 290325 -4522 290561
rect -4286 290325 -4202 290561
rect -3966 290325 -3882 290561
rect -3646 290325 -3538 290561
rect -4950 283561 -3538 290325
rect -4950 283325 -4842 283561
rect -4606 283325 -4522 283561
rect -4286 283325 -4202 283561
rect -3966 283325 -3882 283561
rect -3646 283325 -3538 283561
rect -4950 276561 -3538 283325
rect -4950 276325 -4842 276561
rect -4606 276325 -4522 276561
rect -4286 276325 -4202 276561
rect -3966 276325 -3882 276561
rect -3646 276325 -3538 276561
rect -4950 269561 -3538 276325
rect -4950 269325 -4842 269561
rect -4606 269325 -4522 269561
rect -4286 269325 -4202 269561
rect -3966 269325 -3882 269561
rect -3646 269325 -3538 269561
rect -4950 262561 -3538 269325
rect -4950 262325 -4842 262561
rect -4606 262325 -4522 262561
rect -4286 262325 -4202 262561
rect -3966 262325 -3882 262561
rect -3646 262325 -3538 262561
rect -4950 255561 -3538 262325
rect -4950 255325 -4842 255561
rect -4606 255325 -4522 255561
rect -4286 255325 -4202 255561
rect -3966 255325 -3882 255561
rect -3646 255325 -3538 255561
rect -4950 248561 -3538 255325
rect -4950 248325 -4842 248561
rect -4606 248325 -4522 248561
rect -4286 248325 -4202 248561
rect -3966 248325 -3882 248561
rect -3646 248325 -3538 248561
rect -4950 241561 -3538 248325
rect -4950 241325 -4842 241561
rect -4606 241325 -4522 241561
rect -4286 241325 -4202 241561
rect -3966 241325 -3882 241561
rect -3646 241325 -3538 241561
rect -4950 234561 -3538 241325
rect -4950 234325 -4842 234561
rect -4606 234325 -4522 234561
rect -4286 234325 -4202 234561
rect -3966 234325 -3882 234561
rect -3646 234325 -3538 234561
rect -4950 227561 -3538 234325
rect -4950 227325 -4842 227561
rect -4606 227325 -4522 227561
rect -4286 227325 -4202 227561
rect -3966 227325 -3882 227561
rect -3646 227325 -3538 227561
rect -4950 220561 -3538 227325
rect -4950 220325 -4842 220561
rect -4606 220325 -4522 220561
rect -4286 220325 -4202 220561
rect -3966 220325 -3882 220561
rect -3646 220325 -3538 220561
rect -4950 213561 -3538 220325
rect -4950 213325 -4842 213561
rect -4606 213325 -4522 213561
rect -4286 213325 -4202 213561
rect -3966 213325 -3882 213561
rect -3646 213325 -3538 213561
rect -4950 206561 -3538 213325
rect -4950 206325 -4842 206561
rect -4606 206325 -4522 206561
rect -4286 206325 -4202 206561
rect -3966 206325 -3882 206561
rect -3646 206325 -3538 206561
rect -4950 199561 -3538 206325
rect -4950 199325 -4842 199561
rect -4606 199325 -4522 199561
rect -4286 199325 -4202 199561
rect -3966 199325 -3882 199561
rect -3646 199325 -3538 199561
rect -4950 192561 -3538 199325
rect -4950 192325 -4842 192561
rect -4606 192325 -4522 192561
rect -4286 192325 -4202 192561
rect -3966 192325 -3882 192561
rect -3646 192325 -3538 192561
rect -4950 185561 -3538 192325
rect -4950 185325 -4842 185561
rect -4606 185325 -4522 185561
rect -4286 185325 -4202 185561
rect -3966 185325 -3882 185561
rect -3646 185325 -3538 185561
rect -4950 178561 -3538 185325
rect -4950 178325 -4842 178561
rect -4606 178325 -4522 178561
rect -4286 178325 -4202 178561
rect -3966 178325 -3882 178561
rect -3646 178325 -3538 178561
rect -4950 171561 -3538 178325
rect -4950 171325 -4842 171561
rect -4606 171325 -4522 171561
rect -4286 171325 -4202 171561
rect -3966 171325 -3882 171561
rect -3646 171325 -3538 171561
rect -4950 164561 -3538 171325
rect -4950 164325 -4842 164561
rect -4606 164325 -4522 164561
rect -4286 164325 -4202 164561
rect -3966 164325 -3882 164561
rect -3646 164325 -3538 164561
rect -4950 157561 -3538 164325
rect -4950 157325 -4842 157561
rect -4606 157325 -4522 157561
rect -4286 157325 -4202 157561
rect -3966 157325 -3882 157561
rect -3646 157325 -3538 157561
rect -4950 150561 -3538 157325
rect -4950 150325 -4842 150561
rect -4606 150325 -4522 150561
rect -4286 150325 -4202 150561
rect -3966 150325 -3882 150561
rect -3646 150325 -3538 150561
rect -4950 143561 -3538 150325
rect -4950 143325 -4842 143561
rect -4606 143325 -4522 143561
rect -4286 143325 -4202 143561
rect -3966 143325 -3882 143561
rect -3646 143325 -3538 143561
rect -4950 136561 -3538 143325
rect -4950 136325 -4842 136561
rect -4606 136325 -4522 136561
rect -4286 136325 -4202 136561
rect -3966 136325 -3882 136561
rect -3646 136325 -3538 136561
rect -4950 129561 -3538 136325
rect -4950 129325 -4842 129561
rect -4606 129325 -4522 129561
rect -4286 129325 -4202 129561
rect -3966 129325 -3882 129561
rect -3646 129325 -3538 129561
rect -4950 122561 -3538 129325
rect -4950 122325 -4842 122561
rect -4606 122325 -4522 122561
rect -4286 122325 -4202 122561
rect -3966 122325 -3882 122561
rect -3646 122325 -3538 122561
rect -4950 115561 -3538 122325
rect -4950 115325 -4842 115561
rect -4606 115325 -4522 115561
rect -4286 115325 -4202 115561
rect -3966 115325 -3882 115561
rect -3646 115325 -3538 115561
rect -4950 108561 -3538 115325
rect -4950 108325 -4842 108561
rect -4606 108325 -4522 108561
rect -4286 108325 -4202 108561
rect -3966 108325 -3882 108561
rect -3646 108325 -3538 108561
rect -4950 101561 -3538 108325
rect -4950 101325 -4842 101561
rect -4606 101325 -4522 101561
rect -4286 101325 -4202 101561
rect -3966 101325 -3882 101561
rect -3646 101325 -3538 101561
rect -4950 94561 -3538 101325
rect -4950 94325 -4842 94561
rect -4606 94325 -4522 94561
rect -4286 94325 -4202 94561
rect -3966 94325 -3882 94561
rect -3646 94325 -3538 94561
rect -4950 87561 -3538 94325
rect -4950 87325 -4842 87561
rect -4606 87325 -4522 87561
rect -4286 87325 -4202 87561
rect -3966 87325 -3882 87561
rect -3646 87325 -3538 87561
rect -4950 80561 -3538 87325
rect -4950 80325 -4842 80561
rect -4606 80325 -4522 80561
rect -4286 80325 -4202 80561
rect -3966 80325 -3882 80561
rect -3646 80325 -3538 80561
rect -4950 73561 -3538 80325
rect -4950 73325 -4842 73561
rect -4606 73325 -4522 73561
rect -4286 73325 -4202 73561
rect -3966 73325 -3882 73561
rect -3646 73325 -3538 73561
rect -4950 66561 -3538 73325
rect -4950 66325 -4842 66561
rect -4606 66325 -4522 66561
rect -4286 66325 -4202 66561
rect -3966 66325 -3882 66561
rect -3646 66325 -3538 66561
rect -4950 59561 -3538 66325
rect -4950 59325 -4842 59561
rect -4606 59325 -4522 59561
rect -4286 59325 -4202 59561
rect -3966 59325 -3882 59561
rect -3646 59325 -3538 59561
rect -4950 52561 -3538 59325
rect -4950 52325 -4842 52561
rect -4606 52325 -4522 52561
rect -4286 52325 -4202 52561
rect -3966 52325 -3882 52561
rect -3646 52325 -3538 52561
rect -4950 45561 -3538 52325
rect -4950 45325 -4842 45561
rect -4606 45325 -4522 45561
rect -4286 45325 -4202 45561
rect -3966 45325 -3882 45561
rect -3646 45325 -3538 45561
rect -4950 38561 -3538 45325
rect -4950 38325 -4842 38561
rect -4606 38325 -4522 38561
rect -4286 38325 -4202 38561
rect -3966 38325 -3882 38561
rect -3646 38325 -3538 38561
rect -4950 31561 -3538 38325
rect -4950 31325 -4842 31561
rect -4606 31325 -4522 31561
rect -4286 31325 -4202 31561
rect -3966 31325 -3882 31561
rect -3646 31325 -3538 31561
rect -4950 24561 -3538 31325
rect -4950 24325 -4842 24561
rect -4606 24325 -4522 24561
rect -4286 24325 -4202 24561
rect -3966 24325 -3882 24561
rect -3646 24325 -3538 24561
rect -4950 17561 -3538 24325
rect -4950 17325 -4842 17561
rect -4606 17325 -4522 17561
rect -4286 17325 -4202 17561
rect -3966 17325 -3882 17561
rect -3646 17325 -3538 17561
rect -4950 10561 -3538 17325
rect -4950 10325 -4842 10561
rect -4606 10325 -4522 10561
rect -4286 10325 -4202 10561
rect -3966 10325 -3882 10561
rect -3646 10325 -3538 10561
rect -4950 3561 -3538 10325
rect -4950 3325 -4842 3561
rect -4606 3325 -4522 3561
rect -4286 3325 -4202 3561
rect -3966 3325 -3882 3561
rect -3646 3325 -3538 3561
rect -4950 -3878 -3538 3325
rect -3198 705238 -1786 706062
rect -3198 705002 -2374 705238
rect -2138 705002 -2054 705238
rect -1818 705002 -1786 705238
rect -3198 704918 -1786 705002
rect -3198 704682 -2374 704918
rect -2138 704682 -2054 704918
rect -1818 704682 -1786 704918
rect -3198 695494 -1786 704682
rect -3198 695258 -3090 695494
rect -2854 695258 -2770 695494
rect -2534 695258 -2450 695494
rect -2214 695258 -2130 695494
rect -1894 695258 -1786 695494
rect -3198 688494 -1786 695258
rect -3198 688258 -3090 688494
rect -2854 688258 -2770 688494
rect -2534 688258 -2450 688494
rect -2214 688258 -2130 688494
rect -1894 688258 -1786 688494
rect -3198 681494 -1786 688258
rect -3198 681258 -3090 681494
rect -2854 681258 -2770 681494
rect -2534 681258 -2450 681494
rect -2214 681258 -2130 681494
rect -1894 681258 -1786 681494
rect -3198 674494 -1786 681258
rect -3198 674258 -3090 674494
rect -2854 674258 -2770 674494
rect -2534 674258 -2450 674494
rect -2214 674258 -2130 674494
rect -1894 674258 -1786 674494
rect -3198 667494 -1786 674258
rect -3198 667258 -3090 667494
rect -2854 667258 -2770 667494
rect -2534 667258 -2450 667494
rect -2214 667258 -2130 667494
rect -1894 667258 -1786 667494
rect -3198 660494 -1786 667258
rect -3198 660258 -3090 660494
rect -2854 660258 -2770 660494
rect -2534 660258 -2450 660494
rect -2214 660258 -2130 660494
rect -1894 660258 -1786 660494
rect -3198 653494 -1786 660258
rect -3198 653258 -3090 653494
rect -2854 653258 -2770 653494
rect -2534 653258 -2450 653494
rect -2214 653258 -2130 653494
rect -1894 653258 -1786 653494
rect -3198 646494 -1786 653258
rect -3198 646258 -3090 646494
rect -2854 646258 -2770 646494
rect -2534 646258 -2450 646494
rect -2214 646258 -2130 646494
rect -1894 646258 -1786 646494
rect -3198 639494 -1786 646258
rect -3198 639258 -3090 639494
rect -2854 639258 -2770 639494
rect -2534 639258 -2450 639494
rect -2214 639258 -2130 639494
rect -1894 639258 -1786 639494
rect -3198 632494 -1786 639258
rect -3198 632258 -3090 632494
rect -2854 632258 -2770 632494
rect -2534 632258 -2450 632494
rect -2214 632258 -2130 632494
rect -1894 632258 -1786 632494
rect -3198 625494 -1786 632258
rect -3198 625258 -3090 625494
rect -2854 625258 -2770 625494
rect -2534 625258 -2450 625494
rect -2214 625258 -2130 625494
rect -1894 625258 -1786 625494
rect -3198 618494 -1786 625258
rect -3198 618258 -3090 618494
rect -2854 618258 -2770 618494
rect -2534 618258 -2450 618494
rect -2214 618258 -2130 618494
rect -1894 618258 -1786 618494
rect -3198 611494 -1786 618258
rect -3198 611258 -3090 611494
rect -2854 611258 -2770 611494
rect -2534 611258 -2450 611494
rect -2214 611258 -2130 611494
rect -1894 611258 -1786 611494
rect -3198 604494 -1786 611258
rect -3198 604258 -3090 604494
rect -2854 604258 -2770 604494
rect -2534 604258 -2450 604494
rect -2214 604258 -2130 604494
rect -1894 604258 -1786 604494
rect -3198 597494 -1786 604258
rect -3198 597258 -3090 597494
rect -2854 597258 -2770 597494
rect -2534 597258 -2450 597494
rect -2214 597258 -2130 597494
rect -1894 597258 -1786 597494
rect -3198 590494 -1786 597258
rect -3198 590258 -3090 590494
rect -2854 590258 -2770 590494
rect -2534 590258 -2450 590494
rect -2214 590258 -2130 590494
rect -1894 590258 -1786 590494
rect -3198 583494 -1786 590258
rect -3198 583258 -3090 583494
rect -2854 583258 -2770 583494
rect -2534 583258 -2450 583494
rect -2214 583258 -2130 583494
rect -1894 583258 -1786 583494
rect -3198 576494 -1786 583258
rect -3198 576258 -3090 576494
rect -2854 576258 -2770 576494
rect -2534 576258 -2450 576494
rect -2214 576258 -2130 576494
rect -1894 576258 -1786 576494
rect -3198 569494 -1786 576258
rect -3198 569258 -3090 569494
rect -2854 569258 -2770 569494
rect -2534 569258 -2450 569494
rect -2214 569258 -2130 569494
rect -1894 569258 -1786 569494
rect -3198 562494 -1786 569258
rect -3198 562258 -3090 562494
rect -2854 562258 -2770 562494
rect -2534 562258 -2450 562494
rect -2214 562258 -2130 562494
rect -1894 562258 -1786 562494
rect -3198 555494 -1786 562258
rect -3198 555258 -3090 555494
rect -2854 555258 -2770 555494
rect -2534 555258 -2450 555494
rect -2214 555258 -2130 555494
rect -1894 555258 -1786 555494
rect -3198 548494 -1786 555258
rect -3198 548258 -3090 548494
rect -2854 548258 -2770 548494
rect -2534 548258 -2450 548494
rect -2214 548258 -2130 548494
rect -1894 548258 -1786 548494
rect -3198 541494 -1786 548258
rect -3198 541258 -3090 541494
rect -2854 541258 -2770 541494
rect -2534 541258 -2450 541494
rect -2214 541258 -2130 541494
rect -1894 541258 -1786 541494
rect -3198 534494 -1786 541258
rect -3198 534258 -3090 534494
rect -2854 534258 -2770 534494
rect -2534 534258 -2450 534494
rect -2214 534258 -2130 534494
rect -1894 534258 -1786 534494
rect -3198 527494 -1786 534258
rect -3198 527258 -3090 527494
rect -2854 527258 -2770 527494
rect -2534 527258 -2450 527494
rect -2214 527258 -2130 527494
rect -1894 527258 -1786 527494
rect -3198 520494 -1786 527258
rect -3198 520258 -3090 520494
rect -2854 520258 -2770 520494
rect -2534 520258 -2450 520494
rect -2214 520258 -2130 520494
rect -1894 520258 -1786 520494
rect -3198 513494 -1786 520258
rect -3198 513258 -3090 513494
rect -2854 513258 -2770 513494
rect -2534 513258 -2450 513494
rect -2214 513258 -2130 513494
rect -1894 513258 -1786 513494
rect -3198 506494 -1786 513258
rect -3198 506258 -3090 506494
rect -2854 506258 -2770 506494
rect -2534 506258 -2450 506494
rect -2214 506258 -2130 506494
rect -1894 506258 -1786 506494
rect -3198 499494 -1786 506258
rect -3198 499258 -3090 499494
rect -2854 499258 -2770 499494
rect -2534 499258 -2450 499494
rect -2214 499258 -2130 499494
rect -1894 499258 -1786 499494
rect -3198 492494 -1786 499258
rect -3198 492258 -3090 492494
rect -2854 492258 -2770 492494
rect -2534 492258 -2450 492494
rect -2214 492258 -2130 492494
rect -1894 492258 -1786 492494
rect -3198 485494 -1786 492258
rect -3198 485258 -3090 485494
rect -2854 485258 -2770 485494
rect -2534 485258 -2450 485494
rect -2214 485258 -2130 485494
rect -1894 485258 -1786 485494
rect -3198 478494 -1786 485258
rect -3198 478258 -3090 478494
rect -2854 478258 -2770 478494
rect -2534 478258 -2450 478494
rect -2214 478258 -2130 478494
rect -1894 478258 -1786 478494
rect -3198 471494 -1786 478258
rect -3198 471258 -3090 471494
rect -2854 471258 -2770 471494
rect -2534 471258 -2450 471494
rect -2214 471258 -2130 471494
rect -1894 471258 -1786 471494
rect -3198 464494 -1786 471258
rect -3198 464258 -3090 464494
rect -2854 464258 -2770 464494
rect -2534 464258 -2450 464494
rect -2214 464258 -2130 464494
rect -1894 464258 -1786 464494
rect -3198 457494 -1786 464258
rect -3198 457258 -3090 457494
rect -2854 457258 -2770 457494
rect -2534 457258 -2450 457494
rect -2214 457258 -2130 457494
rect -1894 457258 -1786 457494
rect -3198 450494 -1786 457258
rect -3198 450258 -3090 450494
rect -2854 450258 -2770 450494
rect -2534 450258 -2450 450494
rect -2214 450258 -2130 450494
rect -1894 450258 -1786 450494
rect -3198 443494 -1786 450258
rect -3198 443258 -3090 443494
rect -2854 443258 -2770 443494
rect -2534 443258 -2450 443494
rect -2214 443258 -2130 443494
rect -1894 443258 -1786 443494
rect -3198 436494 -1786 443258
rect -3198 436258 -3090 436494
rect -2854 436258 -2770 436494
rect -2534 436258 -2450 436494
rect -2214 436258 -2130 436494
rect -1894 436258 -1786 436494
rect -3198 429494 -1786 436258
rect -3198 429258 -3090 429494
rect -2854 429258 -2770 429494
rect -2534 429258 -2450 429494
rect -2214 429258 -2130 429494
rect -1894 429258 -1786 429494
rect -3198 422494 -1786 429258
rect -3198 422258 -3090 422494
rect -2854 422258 -2770 422494
rect -2534 422258 -2450 422494
rect -2214 422258 -2130 422494
rect -1894 422258 -1786 422494
rect -3198 415494 -1786 422258
rect -3198 415258 -3090 415494
rect -2854 415258 -2770 415494
rect -2534 415258 -2450 415494
rect -2214 415258 -2130 415494
rect -1894 415258 -1786 415494
rect -3198 408494 -1786 415258
rect -3198 408258 -3090 408494
rect -2854 408258 -2770 408494
rect -2534 408258 -2450 408494
rect -2214 408258 -2130 408494
rect -1894 408258 -1786 408494
rect -3198 401494 -1786 408258
rect -3198 401258 -3090 401494
rect -2854 401258 -2770 401494
rect -2534 401258 -2450 401494
rect -2214 401258 -2130 401494
rect -1894 401258 -1786 401494
rect -3198 394494 -1786 401258
rect -3198 394258 -3090 394494
rect -2854 394258 -2770 394494
rect -2534 394258 -2450 394494
rect -2214 394258 -2130 394494
rect -1894 394258 -1786 394494
rect -3198 387494 -1786 394258
rect -3198 387258 -3090 387494
rect -2854 387258 -2770 387494
rect -2534 387258 -2450 387494
rect -2214 387258 -2130 387494
rect -1894 387258 -1786 387494
rect -3198 380494 -1786 387258
rect -3198 380258 -3090 380494
rect -2854 380258 -2770 380494
rect -2534 380258 -2450 380494
rect -2214 380258 -2130 380494
rect -1894 380258 -1786 380494
rect -3198 373494 -1786 380258
rect -3198 373258 -3090 373494
rect -2854 373258 -2770 373494
rect -2534 373258 -2450 373494
rect -2214 373258 -2130 373494
rect -1894 373258 -1786 373494
rect -3198 366494 -1786 373258
rect -3198 366258 -3090 366494
rect -2854 366258 -2770 366494
rect -2534 366258 -2450 366494
rect -2214 366258 -2130 366494
rect -1894 366258 -1786 366494
rect -3198 359494 -1786 366258
rect -3198 359258 -3090 359494
rect -2854 359258 -2770 359494
rect -2534 359258 -2450 359494
rect -2214 359258 -2130 359494
rect -1894 359258 -1786 359494
rect -3198 352494 -1786 359258
rect -3198 352258 -3090 352494
rect -2854 352258 -2770 352494
rect -2534 352258 -2450 352494
rect -2214 352258 -2130 352494
rect -1894 352258 -1786 352494
rect -3198 345494 -1786 352258
rect -3198 345258 -3090 345494
rect -2854 345258 -2770 345494
rect -2534 345258 -2450 345494
rect -2214 345258 -2130 345494
rect -1894 345258 -1786 345494
rect -3198 338494 -1786 345258
rect -3198 338258 -3090 338494
rect -2854 338258 -2770 338494
rect -2534 338258 -2450 338494
rect -2214 338258 -2130 338494
rect -1894 338258 -1786 338494
rect -3198 331494 -1786 338258
rect -3198 331258 -3090 331494
rect -2854 331258 -2770 331494
rect -2534 331258 -2450 331494
rect -2214 331258 -2130 331494
rect -1894 331258 -1786 331494
rect -3198 324494 -1786 331258
rect -3198 324258 -3090 324494
rect -2854 324258 -2770 324494
rect -2534 324258 -2450 324494
rect -2214 324258 -2130 324494
rect -1894 324258 -1786 324494
rect -3198 317494 -1786 324258
rect -3198 317258 -3090 317494
rect -2854 317258 -2770 317494
rect -2534 317258 -2450 317494
rect -2214 317258 -2130 317494
rect -1894 317258 -1786 317494
rect -3198 310494 -1786 317258
rect -3198 310258 -3090 310494
rect -2854 310258 -2770 310494
rect -2534 310258 -2450 310494
rect -2214 310258 -2130 310494
rect -1894 310258 -1786 310494
rect -3198 303494 -1786 310258
rect -3198 303258 -3090 303494
rect -2854 303258 -2770 303494
rect -2534 303258 -2450 303494
rect -2214 303258 -2130 303494
rect -1894 303258 -1786 303494
rect -3198 296494 -1786 303258
rect -3198 296258 -3090 296494
rect -2854 296258 -2770 296494
rect -2534 296258 -2450 296494
rect -2214 296258 -2130 296494
rect -1894 296258 -1786 296494
rect -3198 289494 -1786 296258
rect -3198 289258 -3090 289494
rect -2854 289258 -2770 289494
rect -2534 289258 -2450 289494
rect -2214 289258 -2130 289494
rect -1894 289258 -1786 289494
rect -3198 282494 -1786 289258
rect -3198 282258 -3090 282494
rect -2854 282258 -2770 282494
rect -2534 282258 -2450 282494
rect -2214 282258 -2130 282494
rect -1894 282258 -1786 282494
rect -3198 275494 -1786 282258
rect -3198 275258 -3090 275494
rect -2854 275258 -2770 275494
rect -2534 275258 -2450 275494
rect -2214 275258 -2130 275494
rect -1894 275258 -1786 275494
rect -3198 268494 -1786 275258
rect -3198 268258 -3090 268494
rect -2854 268258 -2770 268494
rect -2534 268258 -2450 268494
rect -2214 268258 -2130 268494
rect -1894 268258 -1786 268494
rect -3198 261494 -1786 268258
rect -3198 261258 -3090 261494
rect -2854 261258 -2770 261494
rect -2534 261258 -2450 261494
rect -2214 261258 -2130 261494
rect -1894 261258 -1786 261494
rect -3198 254494 -1786 261258
rect -3198 254258 -3090 254494
rect -2854 254258 -2770 254494
rect -2534 254258 -2450 254494
rect -2214 254258 -2130 254494
rect -1894 254258 -1786 254494
rect -3198 247494 -1786 254258
rect -3198 247258 -3090 247494
rect -2854 247258 -2770 247494
rect -2534 247258 -2450 247494
rect -2214 247258 -2130 247494
rect -1894 247258 -1786 247494
rect -3198 240494 -1786 247258
rect -3198 240258 -3090 240494
rect -2854 240258 -2770 240494
rect -2534 240258 -2450 240494
rect -2214 240258 -2130 240494
rect -1894 240258 -1786 240494
rect -3198 233494 -1786 240258
rect -3198 233258 -3090 233494
rect -2854 233258 -2770 233494
rect -2534 233258 -2450 233494
rect -2214 233258 -2130 233494
rect -1894 233258 -1786 233494
rect -3198 226494 -1786 233258
rect -3198 226258 -3090 226494
rect -2854 226258 -2770 226494
rect -2534 226258 -2450 226494
rect -2214 226258 -2130 226494
rect -1894 226258 -1786 226494
rect -3198 219494 -1786 226258
rect -3198 219258 -3090 219494
rect -2854 219258 -2770 219494
rect -2534 219258 -2450 219494
rect -2214 219258 -2130 219494
rect -1894 219258 -1786 219494
rect -3198 212494 -1786 219258
rect -3198 212258 -3090 212494
rect -2854 212258 -2770 212494
rect -2534 212258 -2450 212494
rect -2214 212258 -2130 212494
rect -1894 212258 -1786 212494
rect -3198 205494 -1786 212258
rect -3198 205258 -3090 205494
rect -2854 205258 -2770 205494
rect -2534 205258 -2450 205494
rect -2214 205258 -2130 205494
rect -1894 205258 -1786 205494
rect -3198 198494 -1786 205258
rect -3198 198258 -3090 198494
rect -2854 198258 -2770 198494
rect -2534 198258 -2450 198494
rect -2214 198258 -2130 198494
rect -1894 198258 -1786 198494
rect -3198 191494 -1786 198258
rect -3198 191258 -3090 191494
rect -2854 191258 -2770 191494
rect -2534 191258 -2450 191494
rect -2214 191258 -2130 191494
rect -1894 191258 -1786 191494
rect -3198 184494 -1786 191258
rect -3198 184258 -3090 184494
rect -2854 184258 -2770 184494
rect -2534 184258 -2450 184494
rect -2214 184258 -2130 184494
rect -1894 184258 -1786 184494
rect -3198 177494 -1786 184258
rect -3198 177258 -3090 177494
rect -2854 177258 -2770 177494
rect -2534 177258 -2450 177494
rect -2214 177258 -2130 177494
rect -1894 177258 -1786 177494
rect -3198 170494 -1786 177258
rect -3198 170258 -3090 170494
rect -2854 170258 -2770 170494
rect -2534 170258 -2450 170494
rect -2214 170258 -2130 170494
rect -1894 170258 -1786 170494
rect -3198 163494 -1786 170258
rect -3198 163258 -3090 163494
rect -2854 163258 -2770 163494
rect -2534 163258 -2450 163494
rect -2214 163258 -2130 163494
rect -1894 163258 -1786 163494
rect -3198 156494 -1786 163258
rect -3198 156258 -3090 156494
rect -2854 156258 -2770 156494
rect -2534 156258 -2450 156494
rect -2214 156258 -2130 156494
rect -1894 156258 -1786 156494
rect -3198 149494 -1786 156258
rect -3198 149258 -3090 149494
rect -2854 149258 -2770 149494
rect -2534 149258 -2450 149494
rect -2214 149258 -2130 149494
rect -1894 149258 -1786 149494
rect -3198 142494 -1786 149258
rect -3198 142258 -3090 142494
rect -2854 142258 -2770 142494
rect -2534 142258 -2450 142494
rect -2214 142258 -2130 142494
rect -1894 142258 -1786 142494
rect -3198 135494 -1786 142258
rect -3198 135258 -3090 135494
rect -2854 135258 -2770 135494
rect -2534 135258 -2450 135494
rect -2214 135258 -2130 135494
rect -1894 135258 -1786 135494
rect -3198 128494 -1786 135258
rect -3198 128258 -3090 128494
rect -2854 128258 -2770 128494
rect -2534 128258 -2450 128494
rect -2214 128258 -2130 128494
rect -1894 128258 -1786 128494
rect -3198 121494 -1786 128258
rect -3198 121258 -3090 121494
rect -2854 121258 -2770 121494
rect -2534 121258 -2450 121494
rect -2214 121258 -2130 121494
rect -1894 121258 -1786 121494
rect -3198 114494 -1786 121258
rect -3198 114258 -3090 114494
rect -2854 114258 -2770 114494
rect -2534 114258 -2450 114494
rect -2214 114258 -2130 114494
rect -1894 114258 -1786 114494
rect -3198 107494 -1786 114258
rect -3198 107258 -3090 107494
rect -2854 107258 -2770 107494
rect -2534 107258 -2450 107494
rect -2214 107258 -2130 107494
rect -1894 107258 -1786 107494
rect -3198 100494 -1786 107258
rect -3198 100258 -3090 100494
rect -2854 100258 -2770 100494
rect -2534 100258 -2450 100494
rect -2214 100258 -2130 100494
rect -1894 100258 -1786 100494
rect -3198 93494 -1786 100258
rect -3198 93258 -3090 93494
rect -2854 93258 -2770 93494
rect -2534 93258 -2450 93494
rect -2214 93258 -2130 93494
rect -1894 93258 -1786 93494
rect -3198 86494 -1786 93258
rect -3198 86258 -3090 86494
rect -2854 86258 -2770 86494
rect -2534 86258 -2450 86494
rect -2214 86258 -2130 86494
rect -1894 86258 -1786 86494
rect -3198 79494 -1786 86258
rect -3198 79258 -3090 79494
rect -2854 79258 -2770 79494
rect -2534 79258 -2450 79494
rect -2214 79258 -2130 79494
rect -1894 79258 -1786 79494
rect -3198 72494 -1786 79258
rect -3198 72258 -3090 72494
rect -2854 72258 -2770 72494
rect -2534 72258 -2450 72494
rect -2214 72258 -2130 72494
rect -1894 72258 -1786 72494
rect -3198 65494 -1786 72258
rect -3198 65258 -3090 65494
rect -2854 65258 -2770 65494
rect -2534 65258 -2450 65494
rect -2214 65258 -2130 65494
rect -1894 65258 -1786 65494
rect -3198 58494 -1786 65258
rect -3198 58258 -3090 58494
rect -2854 58258 -2770 58494
rect -2534 58258 -2450 58494
rect -2214 58258 -2130 58494
rect -1894 58258 -1786 58494
rect -3198 51494 -1786 58258
rect -3198 51258 -3090 51494
rect -2854 51258 -2770 51494
rect -2534 51258 -2450 51494
rect -2214 51258 -2130 51494
rect -1894 51258 -1786 51494
rect -3198 44494 -1786 51258
rect -3198 44258 -3090 44494
rect -2854 44258 -2770 44494
rect -2534 44258 -2450 44494
rect -2214 44258 -2130 44494
rect -1894 44258 -1786 44494
rect -3198 37494 -1786 44258
rect -3198 37258 -3090 37494
rect -2854 37258 -2770 37494
rect -2534 37258 -2450 37494
rect -2214 37258 -2130 37494
rect -1894 37258 -1786 37494
rect -3198 30494 -1786 37258
rect -3198 30258 -3090 30494
rect -2854 30258 -2770 30494
rect -2534 30258 -2450 30494
rect -2214 30258 -2130 30494
rect -1894 30258 -1786 30494
rect -3198 23494 -1786 30258
rect -3198 23258 -3090 23494
rect -2854 23258 -2770 23494
rect -2534 23258 -2450 23494
rect -2214 23258 -2130 23494
rect -1894 23258 -1786 23494
rect -3198 16494 -1786 23258
rect -3198 16258 -3090 16494
rect -2854 16258 -2770 16494
rect -2534 16258 -2450 16494
rect -2214 16258 -2130 16494
rect -1894 16258 -1786 16494
rect -3198 9494 -1786 16258
rect -3198 9258 -3090 9494
rect -2854 9258 -2770 9494
rect -2534 9258 -2450 9494
rect -2214 9258 -2130 9494
rect -1894 9258 -1786 9494
rect -3198 2494 -1786 9258
rect -3198 2258 -3090 2494
rect -2854 2258 -2770 2494
rect -2534 2258 -2450 2494
rect -2214 2258 -2130 2494
rect -1894 2258 -1786 2494
rect -3198 -746 -1786 2258
rect -3198 -982 -2374 -746
rect -2138 -982 -2054 -746
rect -1818 -982 -1786 -746
rect -3198 -1066 -1786 -982
rect -3198 -1302 -2374 -1066
rect -2138 -1302 -2054 -1066
rect -1818 -1302 -1786 -1066
rect -3198 -2126 -1786 -1302
rect 1144 705238 1464 706230
rect 1144 705002 1186 705238
rect 1422 705002 1464 705238
rect 1144 704918 1464 705002
rect 1144 704682 1186 704918
rect 1422 704682 1464 704918
rect 1144 695494 1464 704682
rect 1144 695258 1186 695494
rect 1422 695258 1464 695494
rect 1144 688494 1464 695258
rect 1144 688258 1186 688494
rect 1422 688258 1464 688494
rect 1144 681494 1464 688258
rect 1144 681258 1186 681494
rect 1422 681258 1464 681494
rect 1144 674494 1464 681258
rect 1144 674258 1186 674494
rect 1422 674258 1464 674494
rect 1144 667494 1464 674258
rect 1144 667258 1186 667494
rect 1422 667258 1464 667494
rect 1144 660494 1464 667258
rect 1144 660258 1186 660494
rect 1422 660258 1464 660494
rect 1144 653494 1464 660258
rect 1144 653258 1186 653494
rect 1422 653258 1464 653494
rect 1144 646494 1464 653258
rect 1144 646258 1186 646494
rect 1422 646258 1464 646494
rect 1144 639494 1464 646258
rect 1144 639258 1186 639494
rect 1422 639258 1464 639494
rect 1144 632494 1464 639258
rect 1144 632258 1186 632494
rect 1422 632258 1464 632494
rect 1144 625494 1464 632258
rect 1144 625258 1186 625494
rect 1422 625258 1464 625494
rect 1144 618494 1464 625258
rect 1144 618258 1186 618494
rect 1422 618258 1464 618494
rect 1144 611494 1464 618258
rect 1144 611258 1186 611494
rect 1422 611258 1464 611494
rect 1144 604494 1464 611258
rect 1144 604258 1186 604494
rect 1422 604258 1464 604494
rect 1144 597494 1464 604258
rect 1144 597258 1186 597494
rect 1422 597258 1464 597494
rect 1144 590494 1464 597258
rect 1144 590258 1186 590494
rect 1422 590258 1464 590494
rect 1144 583494 1464 590258
rect 1144 583258 1186 583494
rect 1422 583258 1464 583494
rect 1144 576494 1464 583258
rect 1144 576258 1186 576494
rect 1422 576258 1464 576494
rect 1144 569494 1464 576258
rect 1144 569258 1186 569494
rect 1422 569258 1464 569494
rect 1144 562494 1464 569258
rect 1144 562258 1186 562494
rect 1422 562258 1464 562494
rect 1144 555494 1464 562258
rect 1144 555258 1186 555494
rect 1422 555258 1464 555494
rect 1144 548494 1464 555258
rect 1144 548258 1186 548494
rect 1422 548258 1464 548494
rect 1144 541494 1464 548258
rect 1144 541258 1186 541494
rect 1422 541258 1464 541494
rect 1144 534494 1464 541258
rect 1144 534258 1186 534494
rect 1422 534258 1464 534494
rect 1144 527494 1464 534258
rect 1144 527258 1186 527494
rect 1422 527258 1464 527494
rect 1144 520494 1464 527258
rect 1144 520258 1186 520494
rect 1422 520258 1464 520494
rect 1144 513494 1464 520258
rect 1144 513258 1186 513494
rect 1422 513258 1464 513494
rect 1144 506494 1464 513258
rect 1144 506258 1186 506494
rect 1422 506258 1464 506494
rect 1144 499494 1464 506258
rect 1144 499258 1186 499494
rect 1422 499258 1464 499494
rect 1144 492494 1464 499258
rect 1144 492258 1186 492494
rect 1422 492258 1464 492494
rect 1144 485494 1464 492258
rect 1144 485258 1186 485494
rect 1422 485258 1464 485494
rect 1144 478494 1464 485258
rect 1144 478258 1186 478494
rect 1422 478258 1464 478494
rect 1144 471494 1464 478258
rect 1144 471258 1186 471494
rect 1422 471258 1464 471494
rect 1144 464494 1464 471258
rect 1144 464258 1186 464494
rect 1422 464258 1464 464494
rect 1144 457494 1464 464258
rect 1144 457258 1186 457494
rect 1422 457258 1464 457494
rect 1144 450494 1464 457258
rect 1144 450258 1186 450494
rect 1422 450258 1464 450494
rect 1144 443494 1464 450258
rect 1144 443258 1186 443494
rect 1422 443258 1464 443494
rect 1144 436494 1464 443258
rect 1144 436258 1186 436494
rect 1422 436258 1464 436494
rect 1144 429494 1464 436258
rect 1144 429258 1186 429494
rect 1422 429258 1464 429494
rect 1144 422494 1464 429258
rect 1144 422258 1186 422494
rect 1422 422258 1464 422494
rect 1144 415494 1464 422258
rect 1144 415258 1186 415494
rect 1422 415258 1464 415494
rect 1144 408494 1464 415258
rect 1144 408258 1186 408494
rect 1422 408258 1464 408494
rect 1144 401494 1464 408258
rect 1144 401258 1186 401494
rect 1422 401258 1464 401494
rect 1144 394494 1464 401258
rect 1144 394258 1186 394494
rect 1422 394258 1464 394494
rect 1144 387494 1464 394258
rect 1144 387258 1186 387494
rect 1422 387258 1464 387494
rect 1144 380494 1464 387258
rect 1144 380258 1186 380494
rect 1422 380258 1464 380494
rect 1144 373494 1464 380258
rect 1144 373258 1186 373494
rect 1422 373258 1464 373494
rect 1144 366494 1464 373258
rect 1144 366258 1186 366494
rect 1422 366258 1464 366494
rect 1144 359494 1464 366258
rect 1144 359258 1186 359494
rect 1422 359258 1464 359494
rect 1144 352494 1464 359258
rect 1144 352258 1186 352494
rect 1422 352258 1464 352494
rect 1144 345494 1464 352258
rect 1144 345258 1186 345494
rect 1422 345258 1464 345494
rect 1144 338494 1464 345258
rect 1144 338258 1186 338494
rect 1422 338258 1464 338494
rect 1144 331494 1464 338258
rect 1144 331258 1186 331494
rect 1422 331258 1464 331494
rect 1144 324494 1464 331258
rect 1144 324258 1186 324494
rect 1422 324258 1464 324494
rect 1144 317494 1464 324258
rect 1144 317258 1186 317494
rect 1422 317258 1464 317494
rect 1144 310494 1464 317258
rect 1144 310258 1186 310494
rect 1422 310258 1464 310494
rect 1144 303494 1464 310258
rect 1144 303258 1186 303494
rect 1422 303258 1464 303494
rect 1144 296494 1464 303258
rect 1144 296258 1186 296494
rect 1422 296258 1464 296494
rect 1144 289494 1464 296258
rect 1144 289258 1186 289494
rect 1422 289258 1464 289494
rect 1144 282494 1464 289258
rect 1144 282258 1186 282494
rect 1422 282258 1464 282494
rect 1144 275494 1464 282258
rect 1144 275258 1186 275494
rect 1422 275258 1464 275494
rect 1144 268494 1464 275258
rect 1144 268258 1186 268494
rect 1422 268258 1464 268494
rect 1144 261494 1464 268258
rect 1144 261258 1186 261494
rect 1422 261258 1464 261494
rect 1144 254494 1464 261258
rect 1144 254258 1186 254494
rect 1422 254258 1464 254494
rect 1144 247494 1464 254258
rect 1144 247258 1186 247494
rect 1422 247258 1464 247494
rect 1144 240494 1464 247258
rect 1144 240258 1186 240494
rect 1422 240258 1464 240494
rect 1144 233494 1464 240258
rect 1144 233258 1186 233494
rect 1422 233258 1464 233494
rect 1144 226494 1464 233258
rect 1144 226258 1186 226494
rect 1422 226258 1464 226494
rect 1144 219494 1464 226258
rect 1144 219258 1186 219494
rect 1422 219258 1464 219494
rect 1144 212494 1464 219258
rect 1144 212258 1186 212494
rect 1422 212258 1464 212494
rect 1144 205494 1464 212258
rect 1144 205258 1186 205494
rect 1422 205258 1464 205494
rect 1144 198494 1464 205258
rect 1144 198258 1186 198494
rect 1422 198258 1464 198494
rect 1144 191494 1464 198258
rect 1144 191258 1186 191494
rect 1422 191258 1464 191494
rect 1144 184494 1464 191258
rect 1144 184258 1186 184494
rect 1422 184258 1464 184494
rect 1144 177494 1464 184258
rect 1144 177258 1186 177494
rect 1422 177258 1464 177494
rect 1144 170494 1464 177258
rect 1144 170258 1186 170494
rect 1422 170258 1464 170494
rect 1144 163494 1464 170258
rect 1144 163258 1186 163494
rect 1422 163258 1464 163494
rect 1144 156494 1464 163258
rect 1144 156258 1186 156494
rect 1422 156258 1464 156494
rect 1144 149494 1464 156258
rect 1144 149258 1186 149494
rect 1422 149258 1464 149494
rect 1144 142494 1464 149258
rect 1144 142258 1186 142494
rect 1422 142258 1464 142494
rect 1144 135494 1464 142258
rect 1144 135258 1186 135494
rect 1422 135258 1464 135494
rect 1144 128494 1464 135258
rect 1144 128258 1186 128494
rect 1422 128258 1464 128494
rect 1144 121494 1464 128258
rect 1144 121258 1186 121494
rect 1422 121258 1464 121494
rect 1144 114494 1464 121258
rect 1144 114258 1186 114494
rect 1422 114258 1464 114494
rect 1144 107494 1464 114258
rect 1144 107258 1186 107494
rect 1422 107258 1464 107494
rect 1144 100494 1464 107258
rect 1144 100258 1186 100494
rect 1422 100258 1464 100494
rect 1144 93494 1464 100258
rect 1144 93258 1186 93494
rect 1422 93258 1464 93494
rect 1144 86494 1464 93258
rect 1144 86258 1186 86494
rect 1422 86258 1464 86494
rect 1144 79494 1464 86258
rect 1144 79258 1186 79494
rect 1422 79258 1464 79494
rect 1144 72494 1464 79258
rect 1144 72258 1186 72494
rect 1422 72258 1464 72494
rect 1144 65494 1464 72258
rect 1144 65258 1186 65494
rect 1422 65258 1464 65494
rect 1144 58494 1464 65258
rect 1144 58258 1186 58494
rect 1422 58258 1464 58494
rect 1144 51494 1464 58258
rect 1144 51258 1186 51494
rect 1422 51258 1464 51494
rect 1144 44494 1464 51258
rect 1144 44258 1186 44494
rect 1422 44258 1464 44494
rect 1144 37494 1464 44258
rect 1144 37258 1186 37494
rect 1422 37258 1464 37494
rect 1144 30494 1464 37258
rect 1144 30258 1186 30494
rect 1422 30258 1464 30494
rect 1144 23494 1464 30258
rect 1144 23258 1186 23494
rect 1422 23258 1464 23494
rect 1144 16494 1464 23258
rect 1144 16258 1186 16494
rect 1422 16258 1464 16494
rect 1144 9494 1464 16258
rect 1144 9258 1186 9494
rect 1422 9258 1464 9494
rect 1144 2494 1464 9258
rect 1144 2258 1186 2494
rect 1422 2258 1464 2494
rect 1144 -746 1464 2258
rect 1144 -982 1186 -746
rect 1422 -982 1464 -746
rect 1144 -1066 1464 -982
rect 1144 -1302 1186 -1066
rect 1422 -1302 1464 -1066
rect 1144 -2294 1464 -1302
rect 2876 706198 3196 706230
rect 2876 705962 2918 706198
rect 3154 705962 3196 706198
rect 2876 705878 3196 705962
rect 2876 705642 2918 705878
rect 3154 705642 3196 705878
rect 2876 696561 3196 705642
rect 2876 696325 2918 696561
rect 3154 696325 3196 696561
rect 2876 689561 3196 696325
rect 2876 689325 2918 689561
rect 3154 689325 3196 689561
rect 2876 682561 3196 689325
rect 2876 682325 2918 682561
rect 3154 682325 3196 682561
rect 2876 675561 3196 682325
rect 2876 675325 2918 675561
rect 3154 675325 3196 675561
rect 2876 668561 3196 675325
rect 2876 668325 2918 668561
rect 3154 668325 3196 668561
rect 2876 661561 3196 668325
rect 2876 661325 2918 661561
rect 3154 661325 3196 661561
rect 2876 654561 3196 661325
rect 2876 654325 2918 654561
rect 3154 654325 3196 654561
rect 2876 647561 3196 654325
rect 2876 647325 2918 647561
rect 3154 647325 3196 647561
rect 2876 640561 3196 647325
rect 2876 640325 2918 640561
rect 3154 640325 3196 640561
rect 2876 633561 3196 640325
rect 2876 633325 2918 633561
rect 3154 633325 3196 633561
rect 2876 626561 3196 633325
rect 2876 626325 2918 626561
rect 3154 626325 3196 626561
rect 2876 619561 3196 626325
rect 2876 619325 2918 619561
rect 3154 619325 3196 619561
rect 2876 612561 3196 619325
rect 2876 612325 2918 612561
rect 3154 612325 3196 612561
rect 2876 605561 3196 612325
rect 2876 605325 2918 605561
rect 3154 605325 3196 605561
rect 2876 598561 3196 605325
rect 2876 598325 2918 598561
rect 3154 598325 3196 598561
rect 2876 591561 3196 598325
rect 2876 591325 2918 591561
rect 3154 591325 3196 591561
rect 2876 584561 3196 591325
rect 2876 584325 2918 584561
rect 3154 584325 3196 584561
rect 2876 577561 3196 584325
rect 2876 577325 2918 577561
rect 3154 577325 3196 577561
rect 2876 570561 3196 577325
rect 2876 570325 2918 570561
rect 3154 570325 3196 570561
rect 2876 563561 3196 570325
rect 2876 563325 2918 563561
rect 3154 563325 3196 563561
rect 2876 556561 3196 563325
rect 2876 556325 2918 556561
rect 3154 556325 3196 556561
rect 2876 549561 3196 556325
rect 2876 549325 2918 549561
rect 3154 549325 3196 549561
rect 2876 542561 3196 549325
rect 2876 542325 2918 542561
rect 3154 542325 3196 542561
rect 2876 535561 3196 542325
rect 2876 535325 2918 535561
rect 3154 535325 3196 535561
rect 2876 528561 3196 535325
rect 2876 528325 2918 528561
rect 3154 528325 3196 528561
rect 2876 521561 3196 528325
rect 2876 521325 2918 521561
rect 3154 521325 3196 521561
rect 2876 514561 3196 521325
rect 2876 514325 2918 514561
rect 3154 514325 3196 514561
rect 2876 507561 3196 514325
rect 2876 507325 2918 507561
rect 3154 507325 3196 507561
rect 2876 500561 3196 507325
rect 2876 500325 2918 500561
rect 3154 500325 3196 500561
rect 2876 493561 3196 500325
rect 2876 493325 2918 493561
rect 3154 493325 3196 493561
rect 2876 486561 3196 493325
rect 2876 486325 2918 486561
rect 3154 486325 3196 486561
rect 2876 479561 3196 486325
rect 2876 479325 2918 479561
rect 3154 479325 3196 479561
rect 2876 472561 3196 479325
rect 2876 472325 2918 472561
rect 3154 472325 3196 472561
rect 2876 465561 3196 472325
rect 2876 465325 2918 465561
rect 3154 465325 3196 465561
rect 2876 458561 3196 465325
rect 2876 458325 2918 458561
rect 3154 458325 3196 458561
rect 2876 451561 3196 458325
rect 2876 451325 2918 451561
rect 3154 451325 3196 451561
rect 2876 444561 3196 451325
rect 2876 444325 2918 444561
rect 3154 444325 3196 444561
rect 2876 437561 3196 444325
rect 2876 437325 2918 437561
rect 3154 437325 3196 437561
rect 2876 430561 3196 437325
rect 2876 430325 2918 430561
rect 3154 430325 3196 430561
rect 2876 423561 3196 430325
rect 2876 423325 2918 423561
rect 3154 423325 3196 423561
rect 2876 416561 3196 423325
rect 2876 416325 2918 416561
rect 3154 416325 3196 416561
rect 2876 409561 3196 416325
rect 2876 409325 2918 409561
rect 3154 409325 3196 409561
rect 2876 402561 3196 409325
rect 2876 402325 2918 402561
rect 3154 402325 3196 402561
rect 2876 395561 3196 402325
rect 2876 395325 2918 395561
rect 3154 395325 3196 395561
rect 2876 388561 3196 395325
rect 2876 388325 2918 388561
rect 3154 388325 3196 388561
rect 2876 381561 3196 388325
rect 2876 381325 2918 381561
rect 3154 381325 3196 381561
rect 2876 374561 3196 381325
rect 2876 374325 2918 374561
rect 3154 374325 3196 374561
rect 2876 367561 3196 374325
rect 2876 367325 2918 367561
rect 3154 367325 3196 367561
rect 2876 360561 3196 367325
rect 2876 360325 2918 360561
rect 3154 360325 3196 360561
rect 2876 353561 3196 360325
rect 2876 353325 2918 353561
rect 3154 353325 3196 353561
rect 2876 346561 3196 353325
rect 2876 346325 2918 346561
rect 3154 346325 3196 346561
rect 2876 339561 3196 346325
rect 2876 339325 2918 339561
rect 3154 339325 3196 339561
rect 2876 332561 3196 339325
rect 2876 332325 2918 332561
rect 3154 332325 3196 332561
rect 2876 325561 3196 332325
rect 2876 325325 2918 325561
rect 3154 325325 3196 325561
rect 2876 318561 3196 325325
rect 2876 318325 2918 318561
rect 3154 318325 3196 318561
rect 2876 311561 3196 318325
rect 2876 311325 2918 311561
rect 3154 311325 3196 311561
rect 2876 304561 3196 311325
rect 2876 304325 2918 304561
rect 3154 304325 3196 304561
rect 2876 297561 3196 304325
rect 2876 297325 2918 297561
rect 3154 297325 3196 297561
rect 2876 290561 3196 297325
rect 2876 290325 2918 290561
rect 3154 290325 3196 290561
rect 2876 283561 3196 290325
rect 2876 283325 2918 283561
rect 3154 283325 3196 283561
rect 2876 276561 3196 283325
rect 2876 276325 2918 276561
rect 3154 276325 3196 276561
rect 2876 269561 3196 276325
rect 2876 269325 2918 269561
rect 3154 269325 3196 269561
rect 2876 262561 3196 269325
rect 2876 262325 2918 262561
rect 3154 262325 3196 262561
rect 2876 255561 3196 262325
rect 2876 255325 2918 255561
rect 3154 255325 3196 255561
rect 2876 248561 3196 255325
rect 2876 248325 2918 248561
rect 3154 248325 3196 248561
rect 2876 241561 3196 248325
rect 2876 241325 2918 241561
rect 3154 241325 3196 241561
rect 2876 234561 3196 241325
rect 2876 234325 2918 234561
rect 3154 234325 3196 234561
rect 2876 227561 3196 234325
rect 2876 227325 2918 227561
rect 3154 227325 3196 227561
rect 2876 220561 3196 227325
rect 2876 220325 2918 220561
rect 3154 220325 3196 220561
rect 2876 213561 3196 220325
rect 2876 213325 2918 213561
rect 3154 213325 3196 213561
rect 2876 206561 3196 213325
rect 2876 206325 2918 206561
rect 3154 206325 3196 206561
rect 2876 199561 3196 206325
rect 2876 199325 2918 199561
rect 3154 199325 3196 199561
rect 2876 192561 3196 199325
rect 2876 192325 2918 192561
rect 3154 192325 3196 192561
rect 2876 185561 3196 192325
rect 2876 185325 2918 185561
rect 3154 185325 3196 185561
rect 2876 178561 3196 185325
rect 2876 178325 2918 178561
rect 3154 178325 3196 178561
rect 2876 171561 3196 178325
rect 2876 171325 2918 171561
rect 3154 171325 3196 171561
rect 2876 164561 3196 171325
rect 2876 164325 2918 164561
rect 3154 164325 3196 164561
rect 2876 157561 3196 164325
rect 2876 157325 2918 157561
rect 3154 157325 3196 157561
rect 2876 150561 3196 157325
rect 2876 150325 2918 150561
rect 3154 150325 3196 150561
rect 2876 143561 3196 150325
rect 2876 143325 2918 143561
rect 3154 143325 3196 143561
rect 2876 136561 3196 143325
rect 2876 136325 2918 136561
rect 3154 136325 3196 136561
rect 2876 129561 3196 136325
rect 2876 129325 2918 129561
rect 3154 129325 3196 129561
rect 2876 122561 3196 129325
rect 2876 122325 2918 122561
rect 3154 122325 3196 122561
rect 2876 115561 3196 122325
rect 2876 115325 2918 115561
rect 3154 115325 3196 115561
rect 2876 108561 3196 115325
rect 2876 108325 2918 108561
rect 3154 108325 3196 108561
rect 2876 101561 3196 108325
rect 2876 101325 2918 101561
rect 3154 101325 3196 101561
rect 2876 94561 3196 101325
rect 2876 94325 2918 94561
rect 3154 94325 3196 94561
rect 2876 87561 3196 94325
rect 2876 87325 2918 87561
rect 3154 87325 3196 87561
rect 2876 80561 3196 87325
rect 2876 80325 2918 80561
rect 3154 80325 3196 80561
rect 2876 73561 3196 80325
rect 2876 73325 2918 73561
rect 3154 73325 3196 73561
rect 2876 66561 3196 73325
rect 2876 66325 2918 66561
rect 3154 66325 3196 66561
rect 2876 59561 3196 66325
rect 2876 59325 2918 59561
rect 3154 59325 3196 59561
rect 2876 52561 3196 59325
rect 2876 52325 2918 52561
rect 3154 52325 3196 52561
rect 2876 45561 3196 52325
rect 2876 45325 2918 45561
rect 3154 45325 3196 45561
rect 2876 38561 3196 45325
rect 2876 38325 2918 38561
rect 3154 38325 3196 38561
rect 2876 31561 3196 38325
rect 2876 31325 2918 31561
rect 3154 31325 3196 31561
rect 2876 24561 3196 31325
rect 2876 24325 2918 24561
rect 3154 24325 3196 24561
rect 2876 17561 3196 24325
rect 2876 17325 2918 17561
rect 3154 17325 3196 17561
rect 2876 10561 3196 17325
rect 2876 10325 2918 10561
rect 3154 10325 3196 10561
rect 2876 3561 3196 10325
rect 2876 3325 2918 3561
rect 3154 3325 3196 3561
rect 2876 -1706 3196 3325
rect 2876 -1942 2918 -1706
rect 3154 -1942 3196 -1706
rect 2876 -2026 3196 -1942
rect 2876 -2262 2918 -2026
rect 3154 -2262 3196 -2026
rect 2876 -2294 3196 -2262
rect 8144 705238 8464 706230
rect 8144 705002 8186 705238
rect 8422 705002 8464 705238
rect 8144 704918 8464 705002
rect 8144 704682 8186 704918
rect 8422 704682 8464 704918
rect 8144 695494 8464 704682
rect 8144 695258 8186 695494
rect 8422 695258 8464 695494
rect 8144 688494 8464 695258
rect 8144 688258 8186 688494
rect 8422 688258 8464 688494
rect 8144 681494 8464 688258
rect 8144 681258 8186 681494
rect 8422 681258 8464 681494
rect 8144 674494 8464 681258
rect 8144 674258 8186 674494
rect 8422 674258 8464 674494
rect 8144 667494 8464 674258
rect 8144 667258 8186 667494
rect 8422 667258 8464 667494
rect 8144 660494 8464 667258
rect 8144 660258 8186 660494
rect 8422 660258 8464 660494
rect 8144 653494 8464 660258
rect 8144 653258 8186 653494
rect 8422 653258 8464 653494
rect 8144 646494 8464 653258
rect 8144 646258 8186 646494
rect 8422 646258 8464 646494
rect 8144 639494 8464 646258
rect 8144 639258 8186 639494
rect 8422 639258 8464 639494
rect 8144 632494 8464 639258
rect 8144 632258 8186 632494
rect 8422 632258 8464 632494
rect 8144 625494 8464 632258
rect 8144 625258 8186 625494
rect 8422 625258 8464 625494
rect 8144 618494 8464 625258
rect 8144 618258 8186 618494
rect 8422 618258 8464 618494
rect 8144 611494 8464 618258
rect 8144 611258 8186 611494
rect 8422 611258 8464 611494
rect 8144 604494 8464 611258
rect 8144 604258 8186 604494
rect 8422 604258 8464 604494
rect 8144 597494 8464 604258
rect 8144 597258 8186 597494
rect 8422 597258 8464 597494
rect 8144 590494 8464 597258
rect 8144 590258 8186 590494
rect 8422 590258 8464 590494
rect 8144 583494 8464 590258
rect 8144 583258 8186 583494
rect 8422 583258 8464 583494
rect 8144 576494 8464 583258
rect 8144 576258 8186 576494
rect 8422 576258 8464 576494
rect 8144 569494 8464 576258
rect 8144 569258 8186 569494
rect 8422 569258 8464 569494
rect 8144 562494 8464 569258
rect 8144 562258 8186 562494
rect 8422 562258 8464 562494
rect 8144 555494 8464 562258
rect 8144 555258 8186 555494
rect 8422 555258 8464 555494
rect 8144 548494 8464 555258
rect 8144 548258 8186 548494
rect 8422 548258 8464 548494
rect 8144 541494 8464 548258
rect 8144 541258 8186 541494
rect 8422 541258 8464 541494
rect 8144 534494 8464 541258
rect 8144 534258 8186 534494
rect 8422 534258 8464 534494
rect 8144 527494 8464 534258
rect 8144 527258 8186 527494
rect 8422 527258 8464 527494
rect 8144 520494 8464 527258
rect 8144 520258 8186 520494
rect 8422 520258 8464 520494
rect 8144 513494 8464 520258
rect 8144 513258 8186 513494
rect 8422 513258 8464 513494
rect 8144 506494 8464 513258
rect 8144 506258 8186 506494
rect 8422 506258 8464 506494
rect 8144 499494 8464 506258
rect 8144 499258 8186 499494
rect 8422 499258 8464 499494
rect 8144 492494 8464 499258
rect 8144 492258 8186 492494
rect 8422 492258 8464 492494
rect 8144 485494 8464 492258
rect 8144 485258 8186 485494
rect 8422 485258 8464 485494
rect 8144 478494 8464 485258
rect 8144 478258 8186 478494
rect 8422 478258 8464 478494
rect 8144 471494 8464 478258
rect 8144 471258 8186 471494
rect 8422 471258 8464 471494
rect 8144 464494 8464 471258
rect 8144 464258 8186 464494
rect 8422 464258 8464 464494
rect 8144 457494 8464 464258
rect 8144 457258 8186 457494
rect 8422 457258 8464 457494
rect 8144 450494 8464 457258
rect 8144 450258 8186 450494
rect 8422 450258 8464 450494
rect 8144 443494 8464 450258
rect 8144 443258 8186 443494
rect 8422 443258 8464 443494
rect 8144 436494 8464 443258
rect 8144 436258 8186 436494
rect 8422 436258 8464 436494
rect 8144 429494 8464 436258
rect 8144 429258 8186 429494
rect 8422 429258 8464 429494
rect 8144 422494 8464 429258
rect 8144 422258 8186 422494
rect 8422 422258 8464 422494
rect 8144 415494 8464 422258
rect 8144 415258 8186 415494
rect 8422 415258 8464 415494
rect 8144 408494 8464 415258
rect 8144 408258 8186 408494
rect 8422 408258 8464 408494
rect 8144 401494 8464 408258
rect 8144 401258 8186 401494
rect 8422 401258 8464 401494
rect 8144 394494 8464 401258
rect 8144 394258 8186 394494
rect 8422 394258 8464 394494
rect 8144 387494 8464 394258
rect 8144 387258 8186 387494
rect 8422 387258 8464 387494
rect 8144 380494 8464 387258
rect 8144 380258 8186 380494
rect 8422 380258 8464 380494
rect 8144 373494 8464 380258
rect 8144 373258 8186 373494
rect 8422 373258 8464 373494
rect 8144 366494 8464 373258
rect 8144 366258 8186 366494
rect 8422 366258 8464 366494
rect 8144 359494 8464 366258
rect 8144 359258 8186 359494
rect 8422 359258 8464 359494
rect 8144 352494 8464 359258
rect 8144 352258 8186 352494
rect 8422 352258 8464 352494
rect 8144 345494 8464 352258
rect 8144 345258 8186 345494
rect 8422 345258 8464 345494
rect 8144 338494 8464 345258
rect 8144 338258 8186 338494
rect 8422 338258 8464 338494
rect 8144 331494 8464 338258
rect 8144 331258 8186 331494
rect 8422 331258 8464 331494
rect 8144 324494 8464 331258
rect 8144 324258 8186 324494
rect 8422 324258 8464 324494
rect 8144 317494 8464 324258
rect 8144 317258 8186 317494
rect 8422 317258 8464 317494
rect 8144 310494 8464 317258
rect 8144 310258 8186 310494
rect 8422 310258 8464 310494
rect 8144 303494 8464 310258
rect 8144 303258 8186 303494
rect 8422 303258 8464 303494
rect 8144 296494 8464 303258
rect 8144 296258 8186 296494
rect 8422 296258 8464 296494
rect 8144 289494 8464 296258
rect 8144 289258 8186 289494
rect 8422 289258 8464 289494
rect 8144 282494 8464 289258
rect 8144 282258 8186 282494
rect 8422 282258 8464 282494
rect 8144 275494 8464 282258
rect 8144 275258 8186 275494
rect 8422 275258 8464 275494
rect 8144 268494 8464 275258
rect 8144 268258 8186 268494
rect 8422 268258 8464 268494
rect 8144 261494 8464 268258
rect 8144 261258 8186 261494
rect 8422 261258 8464 261494
rect 8144 254494 8464 261258
rect 8144 254258 8186 254494
rect 8422 254258 8464 254494
rect 8144 247494 8464 254258
rect 8144 247258 8186 247494
rect 8422 247258 8464 247494
rect 8144 240494 8464 247258
rect 8144 240258 8186 240494
rect 8422 240258 8464 240494
rect 8144 233494 8464 240258
rect 8144 233258 8186 233494
rect 8422 233258 8464 233494
rect 8144 226494 8464 233258
rect 8144 226258 8186 226494
rect 8422 226258 8464 226494
rect 8144 219494 8464 226258
rect 8144 219258 8186 219494
rect 8422 219258 8464 219494
rect 8144 212494 8464 219258
rect 8144 212258 8186 212494
rect 8422 212258 8464 212494
rect 8144 205494 8464 212258
rect 8144 205258 8186 205494
rect 8422 205258 8464 205494
rect 8144 198494 8464 205258
rect 8144 198258 8186 198494
rect 8422 198258 8464 198494
rect 8144 191494 8464 198258
rect 8144 191258 8186 191494
rect 8422 191258 8464 191494
rect 8144 184494 8464 191258
rect 8144 184258 8186 184494
rect 8422 184258 8464 184494
rect 8144 177494 8464 184258
rect 8144 177258 8186 177494
rect 8422 177258 8464 177494
rect 8144 170494 8464 177258
rect 8144 170258 8186 170494
rect 8422 170258 8464 170494
rect 8144 163494 8464 170258
rect 8144 163258 8186 163494
rect 8422 163258 8464 163494
rect 8144 156494 8464 163258
rect 8144 156258 8186 156494
rect 8422 156258 8464 156494
rect 8144 149494 8464 156258
rect 8144 149258 8186 149494
rect 8422 149258 8464 149494
rect 8144 142494 8464 149258
rect 8144 142258 8186 142494
rect 8422 142258 8464 142494
rect 8144 135494 8464 142258
rect 8144 135258 8186 135494
rect 8422 135258 8464 135494
rect 8144 128494 8464 135258
rect 8144 128258 8186 128494
rect 8422 128258 8464 128494
rect 8144 121494 8464 128258
rect 8144 121258 8186 121494
rect 8422 121258 8464 121494
rect 8144 114494 8464 121258
rect 8144 114258 8186 114494
rect 8422 114258 8464 114494
rect 8144 107494 8464 114258
rect 8144 107258 8186 107494
rect 8422 107258 8464 107494
rect 8144 100494 8464 107258
rect 8144 100258 8186 100494
rect 8422 100258 8464 100494
rect 8144 93494 8464 100258
rect 8144 93258 8186 93494
rect 8422 93258 8464 93494
rect 8144 86494 8464 93258
rect 8144 86258 8186 86494
rect 8422 86258 8464 86494
rect 8144 79494 8464 86258
rect 8144 79258 8186 79494
rect 8422 79258 8464 79494
rect 8144 72494 8464 79258
rect 8144 72258 8186 72494
rect 8422 72258 8464 72494
rect 8144 65494 8464 72258
rect 8144 65258 8186 65494
rect 8422 65258 8464 65494
rect 8144 58494 8464 65258
rect 8144 58258 8186 58494
rect 8422 58258 8464 58494
rect 8144 51494 8464 58258
rect 8144 51258 8186 51494
rect 8422 51258 8464 51494
rect 8144 44494 8464 51258
rect 8144 44258 8186 44494
rect 8422 44258 8464 44494
rect 8144 37494 8464 44258
rect 8144 37258 8186 37494
rect 8422 37258 8464 37494
rect 8144 30494 8464 37258
rect 8144 30258 8186 30494
rect 8422 30258 8464 30494
rect 8144 23494 8464 30258
rect 8144 23258 8186 23494
rect 8422 23258 8464 23494
rect 8144 16494 8464 23258
rect 8144 16258 8186 16494
rect 8422 16258 8464 16494
rect 8144 9494 8464 16258
rect 8144 9258 8186 9494
rect 8422 9258 8464 9494
rect 8144 2494 8464 9258
rect 8144 2258 8186 2494
rect 8422 2258 8464 2494
rect 8144 -746 8464 2258
rect 8144 -982 8186 -746
rect 8422 -982 8464 -746
rect 8144 -1066 8464 -982
rect 8144 -1302 8186 -1066
rect 8422 -1302 8464 -1066
rect 8144 -2294 8464 -1302
rect 9876 706198 10196 706230
rect 9876 705962 9918 706198
rect 10154 705962 10196 706198
rect 9876 705878 10196 705962
rect 9876 705642 9918 705878
rect 10154 705642 10196 705878
rect 9876 696561 10196 705642
rect 9876 696325 9918 696561
rect 10154 696325 10196 696561
rect 9876 689561 10196 696325
rect 9876 689325 9918 689561
rect 10154 689325 10196 689561
rect 9876 682561 10196 689325
rect 9876 682325 9918 682561
rect 10154 682325 10196 682561
rect 9876 675561 10196 682325
rect 9876 675325 9918 675561
rect 10154 675325 10196 675561
rect 9876 668561 10196 675325
rect 9876 668325 9918 668561
rect 10154 668325 10196 668561
rect 9876 661561 10196 668325
rect 9876 661325 9918 661561
rect 10154 661325 10196 661561
rect 9876 654561 10196 661325
rect 9876 654325 9918 654561
rect 10154 654325 10196 654561
rect 9876 647561 10196 654325
rect 9876 647325 9918 647561
rect 10154 647325 10196 647561
rect 9876 640561 10196 647325
rect 9876 640325 9918 640561
rect 10154 640325 10196 640561
rect 9876 633561 10196 640325
rect 9876 633325 9918 633561
rect 10154 633325 10196 633561
rect 9876 626561 10196 633325
rect 9876 626325 9918 626561
rect 10154 626325 10196 626561
rect 9876 619561 10196 626325
rect 9876 619325 9918 619561
rect 10154 619325 10196 619561
rect 9876 612561 10196 619325
rect 9876 612325 9918 612561
rect 10154 612325 10196 612561
rect 9876 605561 10196 612325
rect 9876 605325 9918 605561
rect 10154 605325 10196 605561
rect 9876 598561 10196 605325
rect 9876 598325 9918 598561
rect 10154 598325 10196 598561
rect 9876 591561 10196 598325
rect 9876 591325 9918 591561
rect 10154 591325 10196 591561
rect 9876 584561 10196 591325
rect 9876 584325 9918 584561
rect 10154 584325 10196 584561
rect 9876 577561 10196 584325
rect 9876 577325 9918 577561
rect 10154 577325 10196 577561
rect 9876 570561 10196 577325
rect 9876 570325 9918 570561
rect 10154 570325 10196 570561
rect 9876 563561 10196 570325
rect 9876 563325 9918 563561
rect 10154 563325 10196 563561
rect 9876 556561 10196 563325
rect 9876 556325 9918 556561
rect 10154 556325 10196 556561
rect 9876 549561 10196 556325
rect 9876 549325 9918 549561
rect 10154 549325 10196 549561
rect 9876 542561 10196 549325
rect 9876 542325 9918 542561
rect 10154 542325 10196 542561
rect 9876 535561 10196 542325
rect 9876 535325 9918 535561
rect 10154 535325 10196 535561
rect 9876 528561 10196 535325
rect 9876 528325 9918 528561
rect 10154 528325 10196 528561
rect 9876 521561 10196 528325
rect 9876 521325 9918 521561
rect 10154 521325 10196 521561
rect 9876 514561 10196 521325
rect 9876 514325 9918 514561
rect 10154 514325 10196 514561
rect 9876 507561 10196 514325
rect 9876 507325 9918 507561
rect 10154 507325 10196 507561
rect 9876 500561 10196 507325
rect 9876 500325 9918 500561
rect 10154 500325 10196 500561
rect 9876 493561 10196 500325
rect 9876 493325 9918 493561
rect 10154 493325 10196 493561
rect 9876 486561 10196 493325
rect 9876 486325 9918 486561
rect 10154 486325 10196 486561
rect 9876 479561 10196 486325
rect 9876 479325 9918 479561
rect 10154 479325 10196 479561
rect 9876 472561 10196 479325
rect 9876 472325 9918 472561
rect 10154 472325 10196 472561
rect 9876 465561 10196 472325
rect 9876 465325 9918 465561
rect 10154 465325 10196 465561
rect 9876 458561 10196 465325
rect 9876 458325 9918 458561
rect 10154 458325 10196 458561
rect 9876 451561 10196 458325
rect 9876 451325 9918 451561
rect 10154 451325 10196 451561
rect 9876 444561 10196 451325
rect 9876 444325 9918 444561
rect 10154 444325 10196 444561
rect 9876 437561 10196 444325
rect 9876 437325 9918 437561
rect 10154 437325 10196 437561
rect 9876 430561 10196 437325
rect 9876 430325 9918 430561
rect 10154 430325 10196 430561
rect 9876 423561 10196 430325
rect 9876 423325 9918 423561
rect 10154 423325 10196 423561
rect 9876 416561 10196 423325
rect 9876 416325 9918 416561
rect 10154 416325 10196 416561
rect 9876 409561 10196 416325
rect 9876 409325 9918 409561
rect 10154 409325 10196 409561
rect 9876 402561 10196 409325
rect 9876 402325 9918 402561
rect 10154 402325 10196 402561
rect 9876 395561 10196 402325
rect 9876 395325 9918 395561
rect 10154 395325 10196 395561
rect 9876 388561 10196 395325
rect 9876 388325 9918 388561
rect 10154 388325 10196 388561
rect 9876 381561 10196 388325
rect 9876 381325 9918 381561
rect 10154 381325 10196 381561
rect 9876 374561 10196 381325
rect 9876 374325 9918 374561
rect 10154 374325 10196 374561
rect 9876 367561 10196 374325
rect 9876 367325 9918 367561
rect 10154 367325 10196 367561
rect 9876 360561 10196 367325
rect 9876 360325 9918 360561
rect 10154 360325 10196 360561
rect 9876 353561 10196 360325
rect 9876 353325 9918 353561
rect 10154 353325 10196 353561
rect 9876 346561 10196 353325
rect 9876 346325 9918 346561
rect 10154 346325 10196 346561
rect 9876 339561 10196 346325
rect 9876 339325 9918 339561
rect 10154 339325 10196 339561
rect 9876 332561 10196 339325
rect 9876 332325 9918 332561
rect 10154 332325 10196 332561
rect 9876 325561 10196 332325
rect 9876 325325 9918 325561
rect 10154 325325 10196 325561
rect 9876 318561 10196 325325
rect 9876 318325 9918 318561
rect 10154 318325 10196 318561
rect 9876 311561 10196 318325
rect 9876 311325 9918 311561
rect 10154 311325 10196 311561
rect 9876 304561 10196 311325
rect 9876 304325 9918 304561
rect 10154 304325 10196 304561
rect 9876 297561 10196 304325
rect 9876 297325 9918 297561
rect 10154 297325 10196 297561
rect 9876 290561 10196 297325
rect 9876 290325 9918 290561
rect 10154 290325 10196 290561
rect 9876 283561 10196 290325
rect 9876 283325 9918 283561
rect 10154 283325 10196 283561
rect 9876 276561 10196 283325
rect 9876 276325 9918 276561
rect 10154 276325 10196 276561
rect 9876 269561 10196 276325
rect 9876 269325 9918 269561
rect 10154 269325 10196 269561
rect 9876 262561 10196 269325
rect 9876 262325 9918 262561
rect 10154 262325 10196 262561
rect 9876 255561 10196 262325
rect 9876 255325 9918 255561
rect 10154 255325 10196 255561
rect 9876 248561 10196 255325
rect 9876 248325 9918 248561
rect 10154 248325 10196 248561
rect 9876 241561 10196 248325
rect 9876 241325 9918 241561
rect 10154 241325 10196 241561
rect 9876 234561 10196 241325
rect 9876 234325 9918 234561
rect 10154 234325 10196 234561
rect 9876 227561 10196 234325
rect 9876 227325 9918 227561
rect 10154 227325 10196 227561
rect 9876 220561 10196 227325
rect 9876 220325 9918 220561
rect 10154 220325 10196 220561
rect 9876 213561 10196 220325
rect 9876 213325 9918 213561
rect 10154 213325 10196 213561
rect 9876 206561 10196 213325
rect 9876 206325 9918 206561
rect 10154 206325 10196 206561
rect 9876 199561 10196 206325
rect 9876 199325 9918 199561
rect 10154 199325 10196 199561
rect 9876 192561 10196 199325
rect 9876 192325 9918 192561
rect 10154 192325 10196 192561
rect 9876 185561 10196 192325
rect 9876 185325 9918 185561
rect 10154 185325 10196 185561
rect 9876 178561 10196 185325
rect 9876 178325 9918 178561
rect 10154 178325 10196 178561
rect 9876 171561 10196 178325
rect 9876 171325 9918 171561
rect 10154 171325 10196 171561
rect 9876 164561 10196 171325
rect 9876 164325 9918 164561
rect 10154 164325 10196 164561
rect 9876 157561 10196 164325
rect 9876 157325 9918 157561
rect 10154 157325 10196 157561
rect 9876 150561 10196 157325
rect 9876 150325 9918 150561
rect 10154 150325 10196 150561
rect 9876 143561 10196 150325
rect 9876 143325 9918 143561
rect 10154 143325 10196 143561
rect 9876 136561 10196 143325
rect 9876 136325 9918 136561
rect 10154 136325 10196 136561
rect 9876 129561 10196 136325
rect 9876 129325 9918 129561
rect 10154 129325 10196 129561
rect 9876 122561 10196 129325
rect 9876 122325 9918 122561
rect 10154 122325 10196 122561
rect 9876 115561 10196 122325
rect 9876 115325 9918 115561
rect 10154 115325 10196 115561
rect 9876 108561 10196 115325
rect 9876 108325 9918 108561
rect 10154 108325 10196 108561
rect 9876 101561 10196 108325
rect 9876 101325 9918 101561
rect 10154 101325 10196 101561
rect 9876 94561 10196 101325
rect 9876 94325 9918 94561
rect 10154 94325 10196 94561
rect 9876 87561 10196 94325
rect 9876 87325 9918 87561
rect 10154 87325 10196 87561
rect 9876 80561 10196 87325
rect 9876 80325 9918 80561
rect 10154 80325 10196 80561
rect 9876 73561 10196 80325
rect 9876 73325 9918 73561
rect 10154 73325 10196 73561
rect 9876 66561 10196 73325
rect 9876 66325 9918 66561
rect 10154 66325 10196 66561
rect 9876 59561 10196 66325
rect 9876 59325 9918 59561
rect 10154 59325 10196 59561
rect 9876 52561 10196 59325
rect 9876 52325 9918 52561
rect 10154 52325 10196 52561
rect 9876 45561 10196 52325
rect 9876 45325 9918 45561
rect 10154 45325 10196 45561
rect 9876 38561 10196 45325
rect 9876 38325 9918 38561
rect 10154 38325 10196 38561
rect 9876 31561 10196 38325
rect 9876 31325 9918 31561
rect 10154 31325 10196 31561
rect 9876 24561 10196 31325
rect 9876 24325 9918 24561
rect 10154 24325 10196 24561
rect 9876 17561 10196 24325
rect 9876 17325 9918 17561
rect 10154 17325 10196 17561
rect 9876 10561 10196 17325
rect 9876 10325 9918 10561
rect 10154 10325 10196 10561
rect 9876 3561 10196 10325
rect 9876 3325 9918 3561
rect 10154 3325 10196 3561
rect 9876 -1706 10196 3325
rect 9876 -1942 9918 -1706
rect 10154 -1942 10196 -1706
rect 9876 -2026 10196 -1942
rect 9876 -2262 9918 -2026
rect 10154 -2262 10196 -2026
rect 9876 -2294 10196 -2262
rect 15144 705238 15464 706230
rect 15144 705002 15186 705238
rect 15422 705002 15464 705238
rect 15144 704918 15464 705002
rect 15144 704682 15186 704918
rect 15422 704682 15464 704918
rect 15144 695494 15464 704682
rect 15144 695258 15186 695494
rect 15422 695258 15464 695494
rect 15144 688494 15464 695258
rect 15144 688258 15186 688494
rect 15422 688258 15464 688494
rect 15144 681494 15464 688258
rect 15144 681258 15186 681494
rect 15422 681258 15464 681494
rect 15144 674494 15464 681258
rect 15144 674258 15186 674494
rect 15422 674258 15464 674494
rect 15144 667494 15464 674258
rect 15144 667258 15186 667494
rect 15422 667258 15464 667494
rect 15144 660494 15464 667258
rect 15144 660258 15186 660494
rect 15422 660258 15464 660494
rect 15144 653494 15464 660258
rect 15144 653258 15186 653494
rect 15422 653258 15464 653494
rect 15144 646494 15464 653258
rect 15144 646258 15186 646494
rect 15422 646258 15464 646494
rect 15144 639494 15464 646258
rect 15144 639258 15186 639494
rect 15422 639258 15464 639494
rect 15144 632494 15464 639258
rect 15144 632258 15186 632494
rect 15422 632258 15464 632494
rect 15144 625494 15464 632258
rect 15144 625258 15186 625494
rect 15422 625258 15464 625494
rect 15144 618494 15464 625258
rect 15144 618258 15186 618494
rect 15422 618258 15464 618494
rect 15144 611494 15464 618258
rect 15144 611258 15186 611494
rect 15422 611258 15464 611494
rect 15144 604494 15464 611258
rect 15144 604258 15186 604494
rect 15422 604258 15464 604494
rect 15144 597494 15464 604258
rect 15144 597258 15186 597494
rect 15422 597258 15464 597494
rect 15144 590494 15464 597258
rect 15144 590258 15186 590494
rect 15422 590258 15464 590494
rect 15144 583494 15464 590258
rect 15144 583258 15186 583494
rect 15422 583258 15464 583494
rect 15144 576494 15464 583258
rect 15144 576258 15186 576494
rect 15422 576258 15464 576494
rect 15144 569494 15464 576258
rect 15144 569258 15186 569494
rect 15422 569258 15464 569494
rect 15144 562494 15464 569258
rect 15144 562258 15186 562494
rect 15422 562258 15464 562494
rect 15144 555494 15464 562258
rect 15144 555258 15186 555494
rect 15422 555258 15464 555494
rect 15144 548494 15464 555258
rect 15144 548258 15186 548494
rect 15422 548258 15464 548494
rect 15144 541494 15464 548258
rect 15144 541258 15186 541494
rect 15422 541258 15464 541494
rect 15144 534494 15464 541258
rect 15144 534258 15186 534494
rect 15422 534258 15464 534494
rect 15144 527494 15464 534258
rect 15144 527258 15186 527494
rect 15422 527258 15464 527494
rect 15144 520494 15464 527258
rect 15144 520258 15186 520494
rect 15422 520258 15464 520494
rect 15144 513494 15464 520258
rect 15144 513258 15186 513494
rect 15422 513258 15464 513494
rect 15144 506494 15464 513258
rect 15144 506258 15186 506494
rect 15422 506258 15464 506494
rect 15144 499494 15464 506258
rect 15144 499258 15186 499494
rect 15422 499258 15464 499494
rect 15144 492494 15464 499258
rect 15144 492258 15186 492494
rect 15422 492258 15464 492494
rect 15144 485494 15464 492258
rect 15144 485258 15186 485494
rect 15422 485258 15464 485494
rect 15144 478494 15464 485258
rect 15144 478258 15186 478494
rect 15422 478258 15464 478494
rect 15144 471494 15464 478258
rect 15144 471258 15186 471494
rect 15422 471258 15464 471494
rect 15144 464494 15464 471258
rect 15144 464258 15186 464494
rect 15422 464258 15464 464494
rect 15144 457494 15464 464258
rect 15144 457258 15186 457494
rect 15422 457258 15464 457494
rect 15144 450494 15464 457258
rect 15144 450258 15186 450494
rect 15422 450258 15464 450494
rect 15144 443494 15464 450258
rect 15144 443258 15186 443494
rect 15422 443258 15464 443494
rect 15144 436494 15464 443258
rect 15144 436258 15186 436494
rect 15422 436258 15464 436494
rect 15144 429494 15464 436258
rect 15144 429258 15186 429494
rect 15422 429258 15464 429494
rect 15144 422494 15464 429258
rect 15144 422258 15186 422494
rect 15422 422258 15464 422494
rect 15144 415494 15464 422258
rect 15144 415258 15186 415494
rect 15422 415258 15464 415494
rect 15144 408494 15464 415258
rect 15144 408258 15186 408494
rect 15422 408258 15464 408494
rect 15144 401494 15464 408258
rect 15144 401258 15186 401494
rect 15422 401258 15464 401494
rect 15144 394494 15464 401258
rect 15144 394258 15186 394494
rect 15422 394258 15464 394494
rect 15144 387494 15464 394258
rect 15144 387258 15186 387494
rect 15422 387258 15464 387494
rect 15144 380494 15464 387258
rect 15144 380258 15186 380494
rect 15422 380258 15464 380494
rect 15144 373494 15464 380258
rect 15144 373258 15186 373494
rect 15422 373258 15464 373494
rect 15144 366494 15464 373258
rect 15144 366258 15186 366494
rect 15422 366258 15464 366494
rect 15144 359494 15464 366258
rect 15144 359258 15186 359494
rect 15422 359258 15464 359494
rect 15144 352494 15464 359258
rect 15144 352258 15186 352494
rect 15422 352258 15464 352494
rect 15144 345494 15464 352258
rect 15144 345258 15186 345494
rect 15422 345258 15464 345494
rect 15144 338494 15464 345258
rect 15144 338258 15186 338494
rect 15422 338258 15464 338494
rect 15144 331494 15464 338258
rect 15144 331258 15186 331494
rect 15422 331258 15464 331494
rect 15144 324494 15464 331258
rect 15144 324258 15186 324494
rect 15422 324258 15464 324494
rect 15144 317494 15464 324258
rect 15144 317258 15186 317494
rect 15422 317258 15464 317494
rect 15144 310494 15464 317258
rect 15144 310258 15186 310494
rect 15422 310258 15464 310494
rect 15144 303494 15464 310258
rect 15144 303258 15186 303494
rect 15422 303258 15464 303494
rect 15144 296494 15464 303258
rect 15144 296258 15186 296494
rect 15422 296258 15464 296494
rect 15144 289494 15464 296258
rect 15144 289258 15186 289494
rect 15422 289258 15464 289494
rect 15144 282494 15464 289258
rect 15144 282258 15186 282494
rect 15422 282258 15464 282494
rect 15144 275494 15464 282258
rect 15144 275258 15186 275494
rect 15422 275258 15464 275494
rect 15144 268494 15464 275258
rect 15144 268258 15186 268494
rect 15422 268258 15464 268494
rect 15144 261494 15464 268258
rect 15144 261258 15186 261494
rect 15422 261258 15464 261494
rect 15144 254494 15464 261258
rect 15144 254258 15186 254494
rect 15422 254258 15464 254494
rect 15144 247494 15464 254258
rect 15144 247258 15186 247494
rect 15422 247258 15464 247494
rect 15144 240494 15464 247258
rect 15144 240258 15186 240494
rect 15422 240258 15464 240494
rect 15144 233494 15464 240258
rect 15144 233258 15186 233494
rect 15422 233258 15464 233494
rect 15144 226494 15464 233258
rect 15144 226258 15186 226494
rect 15422 226258 15464 226494
rect 15144 219494 15464 226258
rect 15144 219258 15186 219494
rect 15422 219258 15464 219494
rect 15144 212494 15464 219258
rect 15144 212258 15186 212494
rect 15422 212258 15464 212494
rect 15144 205494 15464 212258
rect 15144 205258 15186 205494
rect 15422 205258 15464 205494
rect 15144 198494 15464 205258
rect 15144 198258 15186 198494
rect 15422 198258 15464 198494
rect 15144 191494 15464 198258
rect 15144 191258 15186 191494
rect 15422 191258 15464 191494
rect 15144 184494 15464 191258
rect 15144 184258 15186 184494
rect 15422 184258 15464 184494
rect 15144 177494 15464 184258
rect 15144 177258 15186 177494
rect 15422 177258 15464 177494
rect 15144 170494 15464 177258
rect 15144 170258 15186 170494
rect 15422 170258 15464 170494
rect 15144 163494 15464 170258
rect 15144 163258 15186 163494
rect 15422 163258 15464 163494
rect 15144 156494 15464 163258
rect 15144 156258 15186 156494
rect 15422 156258 15464 156494
rect 15144 149494 15464 156258
rect 15144 149258 15186 149494
rect 15422 149258 15464 149494
rect 15144 142494 15464 149258
rect 15144 142258 15186 142494
rect 15422 142258 15464 142494
rect 15144 135494 15464 142258
rect 15144 135258 15186 135494
rect 15422 135258 15464 135494
rect 15144 128494 15464 135258
rect 15144 128258 15186 128494
rect 15422 128258 15464 128494
rect 15144 121494 15464 128258
rect 15144 121258 15186 121494
rect 15422 121258 15464 121494
rect 15144 114494 15464 121258
rect 15144 114258 15186 114494
rect 15422 114258 15464 114494
rect 15144 107494 15464 114258
rect 15144 107258 15186 107494
rect 15422 107258 15464 107494
rect 15144 100494 15464 107258
rect 15144 100258 15186 100494
rect 15422 100258 15464 100494
rect 15144 93494 15464 100258
rect 15144 93258 15186 93494
rect 15422 93258 15464 93494
rect 15144 86494 15464 93258
rect 15144 86258 15186 86494
rect 15422 86258 15464 86494
rect 15144 79494 15464 86258
rect 15144 79258 15186 79494
rect 15422 79258 15464 79494
rect 15144 72494 15464 79258
rect 15144 72258 15186 72494
rect 15422 72258 15464 72494
rect 15144 65494 15464 72258
rect 15144 65258 15186 65494
rect 15422 65258 15464 65494
rect 15144 58494 15464 65258
rect 15144 58258 15186 58494
rect 15422 58258 15464 58494
rect 15144 51494 15464 58258
rect 15144 51258 15186 51494
rect 15422 51258 15464 51494
rect 15144 44494 15464 51258
rect 15144 44258 15186 44494
rect 15422 44258 15464 44494
rect 15144 37494 15464 44258
rect 15144 37258 15186 37494
rect 15422 37258 15464 37494
rect 15144 30494 15464 37258
rect 15144 30258 15186 30494
rect 15422 30258 15464 30494
rect 15144 23494 15464 30258
rect 15144 23258 15186 23494
rect 15422 23258 15464 23494
rect 15144 16494 15464 23258
rect 15144 16258 15186 16494
rect 15422 16258 15464 16494
rect 15144 9494 15464 16258
rect 15144 9258 15186 9494
rect 15422 9258 15464 9494
rect 15144 2494 15464 9258
rect 15144 2258 15186 2494
rect 15422 2258 15464 2494
rect 15144 -746 15464 2258
rect 15144 -982 15186 -746
rect 15422 -982 15464 -746
rect 15144 -1066 15464 -982
rect 15144 -1302 15186 -1066
rect 15422 -1302 15464 -1066
rect 15144 -2294 15464 -1302
rect 16876 706198 17196 706230
rect 16876 705962 16918 706198
rect 17154 705962 17196 706198
rect 16876 705878 17196 705962
rect 16876 705642 16918 705878
rect 17154 705642 17196 705878
rect 16876 696561 17196 705642
rect 16876 696325 16918 696561
rect 17154 696325 17196 696561
rect 16876 689561 17196 696325
rect 16876 689325 16918 689561
rect 17154 689325 17196 689561
rect 16876 682561 17196 689325
rect 16876 682325 16918 682561
rect 17154 682325 17196 682561
rect 16876 675561 17196 682325
rect 16876 675325 16918 675561
rect 17154 675325 17196 675561
rect 16876 668561 17196 675325
rect 16876 668325 16918 668561
rect 17154 668325 17196 668561
rect 16876 661561 17196 668325
rect 16876 661325 16918 661561
rect 17154 661325 17196 661561
rect 16876 654561 17196 661325
rect 16876 654325 16918 654561
rect 17154 654325 17196 654561
rect 16876 647561 17196 654325
rect 16876 647325 16918 647561
rect 17154 647325 17196 647561
rect 16876 640561 17196 647325
rect 16876 640325 16918 640561
rect 17154 640325 17196 640561
rect 16876 633561 17196 640325
rect 16876 633325 16918 633561
rect 17154 633325 17196 633561
rect 16876 626561 17196 633325
rect 16876 626325 16918 626561
rect 17154 626325 17196 626561
rect 16876 619561 17196 626325
rect 16876 619325 16918 619561
rect 17154 619325 17196 619561
rect 16876 612561 17196 619325
rect 16876 612325 16918 612561
rect 17154 612325 17196 612561
rect 16876 605561 17196 612325
rect 16876 605325 16918 605561
rect 17154 605325 17196 605561
rect 16876 598561 17196 605325
rect 16876 598325 16918 598561
rect 17154 598325 17196 598561
rect 16876 591561 17196 598325
rect 16876 591325 16918 591561
rect 17154 591325 17196 591561
rect 16876 584561 17196 591325
rect 16876 584325 16918 584561
rect 17154 584325 17196 584561
rect 16876 577561 17196 584325
rect 16876 577325 16918 577561
rect 17154 577325 17196 577561
rect 16876 570561 17196 577325
rect 16876 570325 16918 570561
rect 17154 570325 17196 570561
rect 16876 563561 17196 570325
rect 16876 563325 16918 563561
rect 17154 563325 17196 563561
rect 16876 556561 17196 563325
rect 16876 556325 16918 556561
rect 17154 556325 17196 556561
rect 16876 549561 17196 556325
rect 16876 549325 16918 549561
rect 17154 549325 17196 549561
rect 16876 542561 17196 549325
rect 16876 542325 16918 542561
rect 17154 542325 17196 542561
rect 16876 535561 17196 542325
rect 16876 535325 16918 535561
rect 17154 535325 17196 535561
rect 16876 528561 17196 535325
rect 16876 528325 16918 528561
rect 17154 528325 17196 528561
rect 16876 521561 17196 528325
rect 16876 521325 16918 521561
rect 17154 521325 17196 521561
rect 16876 514561 17196 521325
rect 16876 514325 16918 514561
rect 17154 514325 17196 514561
rect 16876 507561 17196 514325
rect 16876 507325 16918 507561
rect 17154 507325 17196 507561
rect 16876 500561 17196 507325
rect 16876 500325 16918 500561
rect 17154 500325 17196 500561
rect 16876 493561 17196 500325
rect 16876 493325 16918 493561
rect 17154 493325 17196 493561
rect 16876 486561 17196 493325
rect 16876 486325 16918 486561
rect 17154 486325 17196 486561
rect 16876 479561 17196 486325
rect 16876 479325 16918 479561
rect 17154 479325 17196 479561
rect 16876 472561 17196 479325
rect 16876 472325 16918 472561
rect 17154 472325 17196 472561
rect 16876 465561 17196 472325
rect 16876 465325 16918 465561
rect 17154 465325 17196 465561
rect 16876 458561 17196 465325
rect 16876 458325 16918 458561
rect 17154 458325 17196 458561
rect 16876 451561 17196 458325
rect 16876 451325 16918 451561
rect 17154 451325 17196 451561
rect 16876 444561 17196 451325
rect 16876 444325 16918 444561
rect 17154 444325 17196 444561
rect 16876 437561 17196 444325
rect 16876 437325 16918 437561
rect 17154 437325 17196 437561
rect 16876 430561 17196 437325
rect 16876 430325 16918 430561
rect 17154 430325 17196 430561
rect 16876 423561 17196 430325
rect 16876 423325 16918 423561
rect 17154 423325 17196 423561
rect 16876 416561 17196 423325
rect 16876 416325 16918 416561
rect 17154 416325 17196 416561
rect 16876 409561 17196 416325
rect 16876 409325 16918 409561
rect 17154 409325 17196 409561
rect 16876 402561 17196 409325
rect 16876 402325 16918 402561
rect 17154 402325 17196 402561
rect 16876 395561 17196 402325
rect 16876 395325 16918 395561
rect 17154 395325 17196 395561
rect 16876 388561 17196 395325
rect 16876 388325 16918 388561
rect 17154 388325 17196 388561
rect 16876 381561 17196 388325
rect 16876 381325 16918 381561
rect 17154 381325 17196 381561
rect 16876 374561 17196 381325
rect 16876 374325 16918 374561
rect 17154 374325 17196 374561
rect 16876 367561 17196 374325
rect 16876 367325 16918 367561
rect 17154 367325 17196 367561
rect 16876 360561 17196 367325
rect 16876 360325 16918 360561
rect 17154 360325 17196 360561
rect 16876 353561 17196 360325
rect 16876 353325 16918 353561
rect 17154 353325 17196 353561
rect 16876 346561 17196 353325
rect 16876 346325 16918 346561
rect 17154 346325 17196 346561
rect 16876 339561 17196 346325
rect 16876 339325 16918 339561
rect 17154 339325 17196 339561
rect 16876 332561 17196 339325
rect 16876 332325 16918 332561
rect 17154 332325 17196 332561
rect 16876 325561 17196 332325
rect 16876 325325 16918 325561
rect 17154 325325 17196 325561
rect 16876 318561 17196 325325
rect 16876 318325 16918 318561
rect 17154 318325 17196 318561
rect 16876 311561 17196 318325
rect 16876 311325 16918 311561
rect 17154 311325 17196 311561
rect 16876 304561 17196 311325
rect 16876 304325 16918 304561
rect 17154 304325 17196 304561
rect 16876 297561 17196 304325
rect 16876 297325 16918 297561
rect 17154 297325 17196 297561
rect 16876 290561 17196 297325
rect 16876 290325 16918 290561
rect 17154 290325 17196 290561
rect 16876 283561 17196 290325
rect 16876 283325 16918 283561
rect 17154 283325 17196 283561
rect 16876 276561 17196 283325
rect 16876 276325 16918 276561
rect 17154 276325 17196 276561
rect 16876 269561 17196 276325
rect 16876 269325 16918 269561
rect 17154 269325 17196 269561
rect 16876 262561 17196 269325
rect 16876 262325 16918 262561
rect 17154 262325 17196 262561
rect 16876 255561 17196 262325
rect 16876 255325 16918 255561
rect 17154 255325 17196 255561
rect 16876 248561 17196 255325
rect 16876 248325 16918 248561
rect 17154 248325 17196 248561
rect 16876 241561 17196 248325
rect 16876 241325 16918 241561
rect 17154 241325 17196 241561
rect 16876 234561 17196 241325
rect 16876 234325 16918 234561
rect 17154 234325 17196 234561
rect 16876 227561 17196 234325
rect 16876 227325 16918 227561
rect 17154 227325 17196 227561
rect 16876 220561 17196 227325
rect 16876 220325 16918 220561
rect 17154 220325 17196 220561
rect 16876 213561 17196 220325
rect 16876 213325 16918 213561
rect 17154 213325 17196 213561
rect 16876 206561 17196 213325
rect 16876 206325 16918 206561
rect 17154 206325 17196 206561
rect 16876 199561 17196 206325
rect 16876 199325 16918 199561
rect 17154 199325 17196 199561
rect 16876 192561 17196 199325
rect 16876 192325 16918 192561
rect 17154 192325 17196 192561
rect 16876 185561 17196 192325
rect 16876 185325 16918 185561
rect 17154 185325 17196 185561
rect 16876 178561 17196 185325
rect 16876 178325 16918 178561
rect 17154 178325 17196 178561
rect 16876 171561 17196 178325
rect 16876 171325 16918 171561
rect 17154 171325 17196 171561
rect 16876 164561 17196 171325
rect 16876 164325 16918 164561
rect 17154 164325 17196 164561
rect 16876 157561 17196 164325
rect 16876 157325 16918 157561
rect 17154 157325 17196 157561
rect 16876 150561 17196 157325
rect 16876 150325 16918 150561
rect 17154 150325 17196 150561
rect 16876 143561 17196 150325
rect 16876 143325 16918 143561
rect 17154 143325 17196 143561
rect 16876 136561 17196 143325
rect 16876 136325 16918 136561
rect 17154 136325 17196 136561
rect 16876 129561 17196 136325
rect 16876 129325 16918 129561
rect 17154 129325 17196 129561
rect 16876 122561 17196 129325
rect 16876 122325 16918 122561
rect 17154 122325 17196 122561
rect 16876 115561 17196 122325
rect 16876 115325 16918 115561
rect 17154 115325 17196 115561
rect 16876 108561 17196 115325
rect 16876 108325 16918 108561
rect 17154 108325 17196 108561
rect 16876 101561 17196 108325
rect 16876 101325 16918 101561
rect 17154 101325 17196 101561
rect 16876 94561 17196 101325
rect 16876 94325 16918 94561
rect 17154 94325 17196 94561
rect 16876 87561 17196 94325
rect 16876 87325 16918 87561
rect 17154 87325 17196 87561
rect 16876 80561 17196 87325
rect 16876 80325 16918 80561
rect 17154 80325 17196 80561
rect 16876 73561 17196 80325
rect 16876 73325 16918 73561
rect 17154 73325 17196 73561
rect 16876 66561 17196 73325
rect 16876 66325 16918 66561
rect 17154 66325 17196 66561
rect 16876 59561 17196 66325
rect 16876 59325 16918 59561
rect 17154 59325 17196 59561
rect 16876 52561 17196 59325
rect 16876 52325 16918 52561
rect 17154 52325 17196 52561
rect 16876 45561 17196 52325
rect 16876 45325 16918 45561
rect 17154 45325 17196 45561
rect 16876 38561 17196 45325
rect 16876 38325 16918 38561
rect 17154 38325 17196 38561
rect 16876 31561 17196 38325
rect 16876 31325 16918 31561
rect 17154 31325 17196 31561
rect 16876 24561 17196 31325
rect 16876 24325 16918 24561
rect 17154 24325 17196 24561
rect 16876 17561 17196 24325
rect 16876 17325 16918 17561
rect 17154 17325 17196 17561
rect 16876 10561 17196 17325
rect 16876 10325 16918 10561
rect 17154 10325 17196 10561
rect 16876 3561 17196 10325
rect 16876 3325 16918 3561
rect 17154 3325 17196 3561
rect 16876 -1706 17196 3325
rect 16876 -1942 16918 -1706
rect 17154 -1942 17196 -1706
rect 16876 -2026 17196 -1942
rect 16876 -2262 16918 -2026
rect 17154 -2262 17196 -2026
rect 16876 -2294 17196 -2262
rect 22144 705238 22464 706230
rect 22144 705002 22186 705238
rect 22422 705002 22464 705238
rect 22144 704918 22464 705002
rect 22144 704682 22186 704918
rect 22422 704682 22464 704918
rect 22144 695494 22464 704682
rect 22144 695258 22186 695494
rect 22422 695258 22464 695494
rect 22144 688494 22464 695258
rect 22144 688258 22186 688494
rect 22422 688258 22464 688494
rect 22144 681494 22464 688258
rect 22144 681258 22186 681494
rect 22422 681258 22464 681494
rect 22144 674494 22464 681258
rect 22144 674258 22186 674494
rect 22422 674258 22464 674494
rect 22144 667494 22464 674258
rect 22144 667258 22186 667494
rect 22422 667258 22464 667494
rect 22144 660494 22464 667258
rect 22144 660258 22186 660494
rect 22422 660258 22464 660494
rect 22144 653494 22464 660258
rect 22144 653258 22186 653494
rect 22422 653258 22464 653494
rect 22144 646494 22464 653258
rect 22144 646258 22186 646494
rect 22422 646258 22464 646494
rect 22144 639494 22464 646258
rect 22144 639258 22186 639494
rect 22422 639258 22464 639494
rect 22144 632494 22464 639258
rect 22144 632258 22186 632494
rect 22422 632258 22464 632494
rect 22144 625494 22464 632258
rect 22144 625258 22186 625494
rect 22422 625258 22464 625494
rect 22144 618494 22464 625258
rect 22144 618258 22186 618494
rect 22422 618258 22464 618494
rect 22144 611494 22464 618258
rect 22144 611258 22186 611494
rect 22422 611258 22464 611494
rect 22144 604494 22464 611258
rect 22144 604258 22186 604494
rect 22422 604258 22464 604494
rect 22144 597494 22464 604258
rect 22144 597258 22186 597494
rect 22422 597258 22464 597494
rect 22144 590494 22464 597258
rect 22144 590258 22186 590494
rect 22422 590258 22464 590494
rect 22144 583494 22464 590258
rect 22144 583258 22186 583494
rect 22422 583258 22464 583494
rect 22144 576494 22464 583258
rect 22144 576258 22186 576494
rect 22422 576258 22464 576494
rect 22144 569494 22464 576258
rect 22144 569258 22186 569494
rect 22422 569258 22464 569494
rect 22144 562494 22464 569258
rect 22144 562258 22186 562494
rect 22422 562258 22464 562494
rect 22144 555494 22464 562258
rect 22144 555258 22186 555494
rect 22422 555258 22464 555494
rect 22144 548494 22464 555258
rect 22144 548258 22186 548494
rect 22422 548258 22464 548494
rect 22144 541494 22464 548258
rect 22144 541258 22186 541494
rect 22422 541258 22464 541494
rect 22144 534494 22464 541258
rect 22144 534258 22186 534494
rect 22422 534258 22464 534494
rect 22144 527494 22464 534258
rect 22144 527258 22186 527494
rect 22422 527258 22464 527494
rect 22144 520494 22464 527258
rect 22144 520258 22186 520494
rect 22422 520258 22464 520494
rect 22144 513494 22464 520258
rect 22144 513258 22186 513494
rect 22422 513258 22464 513494
rect 22144 506494 22464 513258
rect 22144 506258 22186 506494
rect 22422 506258 22464 506494
rect 22144 499494 22464 506258
rect 22144 499258 22186 499494
rect 22422 499258 22464 499494
rect 22144 492494 22464 499258
rect 22144 492258 22186 492494
rect 22422 492258 22464 492494
rect 22144 485494 22464 492258
rect 22144 485258 22186 485494
rect 22422 485258 22464 485494
rect 22144 478494 22464 485258
rect 22144 478258 22186 478494
rect 22422 478258 22464 478494
rect 22144 471494 22464 478258
rect 22144 471258 22186 471494
rect 22422 471258 22464 471494
rect 22144 464494 22464 471258
rect 22144 464258 22186 464494
rect 22422 464258 22464 464494
rect 22144 457494 22464 464258
rect 22144 457258 22186 457494
rect 22422 457258 22464 457494
rect 22144 450494 22464 457258
rect 22144 450258 22186 450494
rect 22422 450258 22464 450494
rect 22144 443494 22464 450258
rect 22144 443258 22186 443494
rect 22422 443258 22464 443494
rect 22144 436494 22464 443258
rect 22144 436258 22186 436494
rect 22422 436258 22464 436494
rect 22144 429494 22464 436258
rect 22144 429258 22186 429494
rect 22422 429258 22464 429494
rect 22144 422494 22464 429258
rect 22144 422258 22186 422494
rect 22422 422258 22464 422494
rect 22144 415494 22464 422258
rect 22144 415258 22186 415494
rect 22422 415258 22464 415494
rect 22144 408494 22464 415258
rect 22144 408258 22186 408494
rect 22422 408258 22464 408494
rect 22144 401494 22464 408258
rect 22144 401258 22186 401494
rect 22422 401258 22464 401494
rect 22144 394494 22464 401258
rect 22144 394258 22186 394494
rect 22422 394258 22464 394494
rect 22144 387494 22464 394258
rect 22144 387258 22186 387494
rect 22422 387258 22464 387494
rect 22144 380494 22464 387258
rect 22144 380258 22186 380494
rect 22422 380258 22464 380494
rect 22144 373494 22464 380258
rect 22144 373258 22186 373494
rect 22422 373258 22464 373494
rect 22144 366494 22464 373258
rect 22144 366258 22186 366494
rect 22422 366258 22464 366494
rect 22144 359494 22464 366258
rect 22144 359258 22186 359494
rect 22422 359258 22464 359494
rect 22144 352494 22464 359258
rect 22144 352258 22186 352494
rect 22422 352258 22464 352494
rect 22144 345494 22464 352258
rect 22144 345258 22186 345494
rect 22422 345258 22464 345494
rect 22144 338494 22464 345258
rect 22144 338258 22186 338494
rect 22422 338258 22464 338494
rect 22144 331494 22464 338258
rect 22144 331258 22186 331494
rect 22422 331258 22464 331494
rect 22144 324494 22464 331258
rect 22144 324258 22186 324494
rect 22422 324258 22464 324494
rect 22144 317494 22464 324258
rect 22144 317258 22186 317494
rect 22422 317258 22464 317494
rect 22144 310494 22464 317258
rect 22144 310258 22186 310494
rect 22422 310258 22464 310494
rect 22144 303494 22464 310258
rect 22144 303258 22186 303494
rect 22422 303258 22464 303494
rect 22144 296494 22464 303258
rect 22144 296258 22186 296494
rect 22422 296258 22464 296494
rect 22144 289494 22464 296258
rect 22144 289258 22186 289494
rect 22422 289258 22464 289494
rect 22144 282494 22464 289258
rect 22144 282258 22186 282494
rect 22422 282258 22464 282494
rect 22144 275494 22464 282258
rect 22144 275258 22186 275494
rect 22422 275258 22464 275494
rect 22144 268494 22464 275258
rect 22144 268258 22186 268494
rect 22422 268258 22464 268494
rect 22144 261494 22464 268258
rect 22144 261258 22186 261494
rect 22422 261258 22464 261494
rect 22144 254494 22464 261258
rect 22144 254258 22186 254494
rect 22422 254258 22464 254494
rect 22144 247494 22464 254258
rect 22144 247258 22186 247494
rect 22422 247258 22464 247494
rect 22144 240494 22464 247258
rect 22144 240258 22186 240494
rect 22422 240258 22464 240494
rect 22144 233494 22464 240258
rect 22144 233258 22186 233494
rect 22422 233258 22464 233494
rect 22144 226494 22464 233258
rect 22144 226258 22186 226494
rect 22422 226258 22464 226494
rect 22144 219494 22464 226258
rect 22144 219258 22186 219494
rect 22422 219258 22464 219494
rect 22144 212494 22464 219258
rect 22144 212258 22186 212494
rect 22422 212258 22464 212494
rect 22144 205494 22464 212258
rect 22144 205258 22186 205494
rect 22422 205258 22464 205494
rect 22144 198494 22464 205258
rect 22144 198258 22186 198494
rect 22422 198258 22464 198494
rect 22144 191494 22464 198258
rect 22144 191258 22186 191494
rect 22422 191258 22464 191494
rect 22144 184494 22464 191258
rect 22144 184258 22186 184494
rect 22422 184258 22464 184494
rect 22144 177494 22464 184258
rect 22144 177258 22186 177494
rect 22422 177258 22464 177494
rect 22144 170494 22464 177258
rect 22144 170258 22186 170494
rect 22422 170258 22464 170494
rect 22144 163494 22464 170258
rect 22144 163258 22186 163494
rect 22422 163258 22464 163494
rect 22144 156494 22464 163258
rect 22144 156258 22186 156494
rect 22422 156258 22464 156494
rect 22144 149494 22464 156258
rect 22144 149258 22186 149494
rect 22422 149258 22464 149494
rect 22144 142494 22464 149258
rect 22144 142258 22186 142494
rect 22422 142258 22464 142494
rect 22144 135494 22464 142258
rect 22144 135258 22186 135494
rect 22422 135258 22464 135494
rect 22144 128494 22464 135258
rect 22144 128258 22186 128494
rect 22422 128258 22464 128494
rect 22144 121494 22464 128258
rect 22144 121258 22186 121494
rect 22422 121258 22464 121494
rect 22144 114494 22464 121258
rect 22144 114258 22186 114494
rect 22422 114258 22464 114494
rect 22144 107494 22464 114258
rect 22144 107258 22186 107494
rect 22422 107258 22464 107494
rect 22144 100494 22464 107258
rect 22144 100258 22186 100494
rect 22422 100258 22464 100494
rect 22144 93494 22464 100258
rect 22144 93258 22186 93494
rect 22422 93258 22464 93494
rect 22144 86494 22464 93258
rect 22144 86258 22186 86494
rect 22422 86258 22464 86494
rect 22144 79494 22464 86258
rect 22144 79258 22186 79494
rect 22422 79258 22464 79494
rect 22144 72494 22464 79258
rect 22144 72258 22186 72494
rect 22422 72258 22464 72494
rect 22144 65494 22464 72258
rect 22144 65258 22186 65494
rect 22422 65258 22464 65494
rect 22144 58494 22464 65258
rect 22144 58258 22186 58494
rect 22422 58258 22464 58494
rect 22144 51494 22464 58258
rect 22144 51258 22186 51494
rect 22422 51258 22464 51494
rect 22144 44494 22464 51258
rect 22144 44258 22186 44494
rect 22422 44258 22464 44494
rect 22144 37494 22464 44258
rect 22144 37258 22186 37494
rect 22422 37258 22464 37494
rect 22144 30494 22464 37258
rect 22144 30258 22186 30494
rect 22422 30258 22464 30494
rect 22144 23494 22464 30258
rect 22144 23258 22186 23494
rect 22422 23258 22464 23494
rect 22144 16494 22464 23258
rect 22144 16258 22186 16494
rect 22422 16258 22464 16494
rect 22144 9494 22464 16258
rect 22144 9258 22186 9494
rect 22422 9258 22464 9494
rect 22144 2494 22464 9258
rect 22144 2258 22186 2494
rect 22422 2258 22464 2494
rect 22144 -746 22464 2258
rect 22144 -982 22186 -746
rect 22422 -982 22464 -746
rect 22144 -1066 22464 -982
rect 22144 -1302 22186 -1066
rect 22422 -1302 22464 -1066
rect 22144 -2294 22464 -1302
rect 23876 706198 24196 706230
rect 23876 705962 23918 706198
rect 24154 705962 24196 706198
rect 23876 705878 24196 705962
rect 23876 705642 23918 705878
rect 24154 705642 24196 705878
rect 23876 696561 24196 705642
rect 23876 696325 23918 696561
rect 24154 696325 24196 696561
rect 23876 689561 24196 696325
rect 23876 689325 23918 689561
rect 24154 689325 24196 689561
rect 23876 682561 24196 689325
rect 23876 682325 23918 682561
rect 24154 682325 24196 682561
rect 23876 675561 24196 682325
rect 23876 675325 23918 675561
rect 24154 675325 24196 675561
rect 23876 668561 24196 675325
rect 23876 668325 23918 668561
rect 24154 668325 24196 668561
rect 23876 661561 24196 668325
rect 23876 661325 23918 661561
rect 24154 661325 24196 661561
rect 23876 654561 24196 661325
rect 23876 654325 23918 654561
rect 24154 654325 24196 654561
rect 23876 647561 24196 654325
rect 23876 647325 23918 647561
rect 24154 647325 24196 647561
rect 23876 640561 24196 647325
rect 23876 640325 23918 640561
rect 24154 640325 24196 640561
rect 23876 633561 24196 640325
rect 23876 633325 23918 633561
rect 24154 633325 24196 633561
rect 23876 626561 24196 633325
rect 23876 626325 23918 626561
rect 24154 626325 24196 626561
rect 23876 619561 24196 626325
rect 23876 619325 23918 619561
rect 24154 619325 24196 619561
rect 23876 612561 24196 619325
rect 23876 612325 23918 612561
rect 24154 612325 24196 612561
rect 23876 605561 24196 612325
rect 23876 605325 23918 605561
rect 24154 605325 24196 605561
rect 23876 598561 24196 605325
rect 23876 598325 23918 598561
rect 24154 598325 24196 598561
rect 23876 591561 24196 598325
rect 23876 591325 23918 591561
rect 24154 591325 24196 591561
rect 23876 584561 24196 591325
rect 23876 584325 23918 584561
rect 24154 584325 24196 584561
rect 23876 577561 24196 584325
rect 23876 577325 23918 577561
rect 24154 577325 24196 577561
rect 23876 570561 24196 577325
rect 23876 570325 23918 570561
rect 24154 570325 24196 570561
rect 23876 563561 24196 570325
rect 23876 563325 23918 563561
rect 24154 563325 24196 563561
rect 23876 556561 24196 563325
rect 23876 556325 23918 556561
rect 24154 556325 24196 556561
rect 23876 549561 24196 556325
rect 23876 549325 23918 549561
rect 24154 549325 24196 549561
rect 23876 542561 24196 549325
rect 23876 542325 23918 542561
rect 24154 542325 24196 542561
rect 23876 535561 24196 542325
rect 23876 535325 23918 535561
rect 24154 535325 24196 535561
rect 23876 528561 24196 535325
rect 23876 528325 23918 528561
rect 24154 528325 24196 528561
rect 23876 521561 24196 528325
rect 23876 521325 23918 521561
rect 24154 521325 24196 521561
rect 23876 514561 24196 521325
rect 23876 514325 23918 514561
rect 24154 514325 24196 514561
rect 23876 507561 24196 514325
rect 23876 507325 23918 507561
rect 24154 507325 24196 507561
rect 23876 500561 24196 507325
rect 23876 500325 23918 500561
rect 24154 500325 24196 500561
rect 23876 493561 24196 500325
rect 23876 493325 23918 493561
rect 24154 493325 24196 493561
rect 23876 486561 24196 493325
rect 23876 486325 23918 486561
rect 24154 486325 24196 486561
rect 23876 479561 24196 486325
rect 23876 479325 23918 479561
rect 24154 479325 24196 479561
rect 23876 472561 24196 479325
rect 23876 472325 23918 472561
rect 24154 472325 24196 472561
rect 23876 465561 24196 472325
rect 23876 465325 23918 465561
rect 24154 465325 24196 465561
rect 23876 458561 24196 465325
rect 23876 458325 23918 458561
rect 24154 458325 24196 458561
rect 23876 451561 24196 458325
rect 23876 451325 23918 451561
rect 24154 451325 24196 451561
rect 23876 444561 24196 451325
rect 23876 444325 23918 444561
rect 24154 444325 24196 444561
rect 23876 437561 24196 444325
rect 23876 437325 23918 437561
rect 24154 437325 24196 437561
rect 23876 430561 24196 437325
rect 23876 430325 23918 430561
rect 24154 430325 24196 430561
rect 23876 423561 24196 430325
rect 23876 423325 23918 423561
rect 24154 423325 24196 423561
rect 23876 416561 24196 423325
rect 23876 416325 23918 416561
rect 24154 416325 24196 416561
rect 23876 409561 24196 416325
rect 23876 409325 23918 409561
rect 24154 409325 24196 409561
rect 23876 402561 24196 409325
rect 23876 402325 23918 402561
rect 24154 402325 24196 402561
rect 23876 395561 24196 402325
rect 23876 395325 23918 395561
rect 24154 395325 24196 395561
rect 23876 388561 24196 395325
rect 23876 388325 23918 388561
rect 24154 388325 24196 388561
rect 23876 381561 24196 388325
rect 23876 381325 23918 381561
rect 24154 381325 24196 381561
rect 23876 374561 24196 381325
rect 23876 374325 23918 374561
rect 24154 374325 24196 374561
rect 23876 367561 24196 374325
rect 23876 367325 23918 367561
rect 24154 367325 24196 367561
rect 23876 360561 24196 367325
rect 23876 360325 23918 360561
rect 24154 360325 24196 360561
rect 23876 353561 24196 360325
rect 23876 353325 23918 353561
rect 24154 353325 24196 353561
rect 23876 346561 24196 353325
rect 23876 346325 23918 346561
rect 24154 346325 24196 346561
rect 23876 339561 24196 346325
rect 23876 339325 23918 339561
rect 24154 339325 24196 339561
rect 23876 332561 24196 339325
rect 23876 332325 23918 332561
rect 24154 332325 24196 332561
rect 23876 325561 24196 332325
rect 23876 325325 23918 325561
rect 24154 325325 24196 325561
rect 23876 318561 24196 325325
rect 23876 318325 23918 318561
rect 24154 318325 24196 318561
rect 23876 311561 24196 318325
rect 23876 311325 23918 311561
rect 24154 311325 24196 311561
rect 23876 304561 24196 311325
rect 23876 304325 23918 304561
rect 24154 304325 24196 304561
rect 23876 297561 24196 304325
rect 23876 297325 23918 297561
rect 24154 297325 24196 297561
rect 23876 290561 24196 297325
rect 23876 290325 23918 290561
rect 24154 290325 24196 290561
rect 23876 283561 24196 290325
rect 23876 283325 23918 283561
rect 24154 283325 24196 283561
rect 23876 276561 24196 283325
rect 23876 276325 23918 276561
rect 24154 276325 24196 276561
rect 23876 269561 24196 276325
rect 23876 269325 23918 269561
rect 24154 269325 24196 269561
rect 23876 262561 24196 269325
rect 23876 262325 23918 262561
rect 24154 262325 24196 262561
rect 23876 255561 24196 262325
rect 23876 255325 23918 255561
rect 24154 255325 24196 255561
rect 23876 248561 24196 255325
rect 23876 248325 23918 248561
rect 24154 248325 24196 248561
rect 23876 241561 24196 248325
rect 23876 241325 23918 241561
rect 24154 241325 24196 241561
rect 23876 234561 24196 241325
rect 23876 234325 23918 234561
rect 24154 234325 24196 234561
rect 23876 227561 24196 234325
rect 23876 227325 23918 227561
rect 24154 227325 24196 227561
rect 23876 220561 24196 227325
rect 23876 220325 23918 220561
rect 24154 220325 24196 220561
rect 23876 213561 24196 220325
rect 23876 213325 23918 213561
rect 24154 213325 24196 213561
rect 23876 206561 24196 213325
rect 23876 206325 23918 206561
rect 24154 206325 24196 206561
rect 23876 199561 24196 206325
rect 23876 199325 23918 199561
rect 24154 199325 24196 199561
rect 23876 192561 24196 199325
rect 23876 192325 23918 192561
rect 24154 192325 24196 192561
rect 23876 185561 24196 192325
rect 23876 185325 23918 185561
rect 24154 185325 24196 185561
rect 23876 178561 24196 185325
rect 23876 178325 23918 178561
rect 24154 178325 24196 178561
rect 23876 171561 24196 178325
rect 23876 171325 23918 171561
rect 24154 171325 24196 171561
rect 23876 164561 24196 171325
rect 23876 164325 23918 164561
rect 24154 164325 24196 164561
rect 23876 157561 24196 164325
rect 23876 157325 23918 157561
rect 24154 157325 24196 157561
rect 23876 150561 24196 157325
rect 23876 150325 23918 150561
rect 24154 150325 24196 150561
rect 23876 143561 24196 150325
rect 23876 143325 23918 143561
rect 24154 143325 24196 143561
rect 23876 136561 24196 143325
rect 23876 136325 23918 136561
rect 24154 136325 24196 136561
rect 23876 129561 24196 136325
rect 23876 129325 23918 129561
rect 24154 129325 24196 129561
rect 23876 122561 24196 129325
rect 23876 122325 23918 122561
rect 24154 122325 24196 122561
rect 23876 115561 24196 122325
rect 23876 115325 23918 115561
rect 24154 115325 24196 115561
rect 23876 108561 24196 115325
rect 23876 108325 23918 108561
rect 24154 108325 24196 108561
rect 23876 101561 24196 108325
rect 23876 101325 23918 101561
rect 24154 101325 24196 101561
rect 23876 94561 24196 101325
rect 23876 94325 23918 94561
rect 24154 94325 24196 94561
rect 23876 87561 24196 94325
rect 23876 87325 23918 87561
rect 24154 87325 24196 87561
rect 23876 80561 24196 87325
rect 23876 80325 23918 80561
rect 24154 80325 24196 80561
rect 23876 73561 24196 80325
rect 23876 73325 23918 73561
rect 24154 73325 24196 73561
rect 23876 66561 24196 73325
rect 23876 66325 23918 66561
rect 24154 66325 24196 66561
rect 23876 59561 24196 66325
rect 23876 59325 23918 59561
rect 24154 59325 24196 59561
rect 23876 52561 24196 59325
rect 23876 52325 23918 52561
rect 24154 52325 24196 52561
rect 23876 45561 24196 52325
rect 23876 45325 23918 45561
rect 24154 45325 24196 45561
rect 23876 38561 24196 45325
rect 23876 38325 23918 38561
rect 24154 38325 24196 38561
rect 23876 31561 24196 38325
rect 23876 31325 23918 31561
rect 24154 31325 24196 31561
rect 23876 24561 24196 31325
rect 23876 24325 23918 24561
rect 24154 24325 24196 24561
rect 23876 17561 24196 24325
rect 23876 17325 23918 17561
rect 24154 17325 24196 17561
rect 23876 10561 24196 17325
rect 23876 10325 23918 10561
rect 24154 10325 24196 10561
rect 23876 3561 24196 10325
rect 23876 3325 23918 3561
rect 24154 3325 24196 3561
rect 23876 -1706 24196 3325
rect 23876 -1942 23918 -1706
rect 24154 -1942 24196 -1706
rect 23876 -2026 24196 -1942
rect 23876 -2262 23918 -2026
rect 24154 -2262 24196 -2026
rect 23876 -2294 24196 -2262
rect 29144 705238 29464 706230
rect 29144 705002 29186 705238
rect 29422 705002 29464 705238
rect 29144 704918 29464 705002
rect 29144 704682 29186 704918
rect 29422 704682 29464 704918
rect 29144 695494 29464 704682
rect 29144 695258 29186 695494
rect 29422 695258 29464 695494
rect 29144 688494 29464 695258
rect 29144 688258 29186 688494
rect 29422 688258 29464 688494
rect 29144 681494 29464 688258
rect 29144 681258 29186 681494
rect 29422 681258 29464 681494
rect 29144 674494 29464 681258
rect 29144 674258 29186 674494
rect 29422 674258 29464 674494
rect 29144 667494 29464 674258
rect 29144 667258 29186 667494
rect 29422 667258 29464 667494
rect 29144 660494 29464 667258
rect 29144 660258 29186 660494
rect 29422 660258 29464 660494
rect 29144 653494 29464 660258
rect 29144 653258 29186 653494
rect 29422 653258 29464 653494
rect 29144 646494 29464 653258
rect 29144 646258 29186 646494
rect 29422 646258 29464 646494
rect 29144 639494 29464 646258
rect 29144 639258 29186 639494
rect 29422 639258 29464 639494
rect 29144 632494 29464 639258
rect 29144 632258 29186 632494
rect 29422 632258 29464 632494
rect 29144 625494 29464 632258
rect 29144 625258 29186 625494
rect 29422 625258 29464 625494
rect 29144 618494 29464 625258
rect 29144 618258 29186 618494
rect 29422 618258 29464 618494
rect 29144 611494 29464 618258
rect 29144 611258 29186 611494
rect 29422 611258 29464 611494
rect 29144 604494 29464 611258
rect 29144 604258 29186 604494
rect 29422 604258 29464 604494
rect 29144 597494 29464 604258
rect 29144 597258 29186 597494
rect 29422 597258 29464 597494
rect 29144 590494 29464 597258
rect 29144 590258 29186 590494
rect 29422 590258 29464 590494
rect 29144 583494 29464 590258
rect 29144 583258 29186 583494
rect 29422 583258 29464 583494
rect 29144 576494 29464 583258
rect 29144 576258 29186 576494
rect 29422 576258 29464 576494
rect 29144 569494 29464 576258
rect 29144 569258 29186 569494
rect 29422 569258 29464 569494
rect 29144 562494 29464 569258
rect 29144 562258 29186 562494
rect 29422 562258 29464 562494
rect 29144 555494 29464 562258
rect 29144 555258 29186 555494
rect 29422 555258 29464 555494
rect 29144 548494 29464 555258
rect 29144 548258 29186 548494
rect 29422 548258 29464 548494
rect 29144 541494 29464 548258
rect 29144 541258 29186 541494
rect 29422 541258 29464 541494
rect 29144 534494 29464 541258
rect 29144 534258 29186 534494
rect 29422 534258 29464 534494
rect 29144 527494 29464 534258
rect 29144 527258 29186 527494
rect 29422 527258 29464 527494
rect 29144 520494 29464 527258
rect 29144 520258 29186 520494
rect 29422 520258 29464 520494
rect 29144 513494 29464 520258
rect 29144 513258 29186 513494
rect 29422 513258 29464 513494
rect 29144 506494 29464 513258
rect 29144 506258 29186 506494
rect 29422 506258 29464 506494
rect 29144 499494 29464 506258
rect 29144 499258 29186 499494
rect 29422 499258 29464 499494
rect 29144 492494 29464 499258
rect 29144 492258 29186 492494
rect 29422 492258 29464 492494
rect 29144 485494 29464 492258
rect 29144 485258 29186 485494
rect 29422 485258 29464 485494
rect 29144 478494 29464 485258
rect 29144 478258 29186 478494
rect 29422 478258 29464 478494
rect 29144 471494 29464 478258
rect 29144 471258 29186 471494
rect 29422 471258 29464 471494
rect 29144 464494 29464 471258
rect 29144 464258 29186 464494
rect 29422 464258 29464 464494
rect 29144 457494 29464 464258
rect 29144 457258 29186 457494
rect 29422 457258 29464 457494
rect 29144 450494 29464 457258
rect 29144 450258 29186 450494
rect 29422 450258 29464 450494
rect 29144 443494 29464 450258
rect 29144 443258 29186 443494
rect 29422 443258 29464 443494
rect 29144 436494 29464 443258
rect 29144 436258 29186 436494
rect 29422 436258 29464 436494
rect 29144 429494 29464 436258
rect 29144 429258 29186 429494
rect 29422 429258 29464 429494
rect 29144 422494 29464 429258
rect 29144 422258 29186 422494
rect 29422 422258 29464 422494
rect 29144 415494 29464 422258
rect 29144 415258 29186 415494
rect 29422 415258 29464 415494
rect 29144 408494 29464 415258
rect 29144 408258 29186 408494
rect 29422 408258 29464 408494
rect 29144 401494 29464 408258
rect 29144 401258 29186 401494
rect 29422 401258 29464 401494
rect 29144 394494 29464 401258
rect 29144 394258 29186 394494
rect 29422 394258 29464 394494
rect 29144 387494 29464 394258
rect 29144 387258 29186 387494
rect 29422 387258 29464 387494
rect 29144 380494 29464 387258
rect 29144 380258 29186 380494
rect 29422 380258 29464 380494
rect 29144 373494 29464 380258
rect 29144 373258 29186 373494
rect 29422 373258 29464 373494
rect 29144 366494 29464 373258
rect 29144 366258 29186 366494
rect 29422 366258 29464 366494
rect 29144 359494 29464 366258
rect 29144 359258 29186 359494
rect 29422 359258 29464 359494
rect 29144 352494 29464 359258
rect 29144 352258 29186 352494
rect 29422 352258 29464 352494
rect 29144 345494 29464 352258
rect 29144 345258 29186 345494
rect 29422 345258 29464 345494
rect 29144 338494 29464 345258
rect 29144 338258 29186 338494
rect 29422 338258 29464 338494
rect 29144 331494 29464 338258
rect 29144 331258 29186 331494
rect 29422 331258 29464 331494
rect 29144 324494 29464 331258
rect 29144 324258 29186 324494
rect 29422 324258 29464 324494
rect 29144 317494 29464 324258
rect 29144 317258 29186 317494
rect 29422 317258 29464 317494
rect 29144 310494 29464 317258
rect 29144 310258 29186 310494
rect 29422 310258 29464 310494
rect 29144 303494 29464 310258
rect 29144 303258 29186 303494
rect 29422 303258 29464 303494
rect 29144 296494 29464 303258
rect 29144 296258 29186 296494
rect 29422 296258 29464 296494
rect 29144 289494 29464 296258
rect 29144 289258 29186 289494
rect 29422 289258 29464 289494
rect 29144 282494 29464 289258
rect 29144 282258 29186 282494
rect 29422 282258 29464 282494
rect 29144 275494 29464 282258
rect 29144 275258 29186 275494
rect 29422 275258 29464 275494
rect 29144 268494 29464 275258
rect 29144 268258 29186 268494
rect 29422 268258 29464 268494
rect 29144 261494 29464 268258
rect 29144 261258 29186 261494
rect 29422 261258 29464 261494
rect 29144 254494 29464 261258
rect 29144 254258 29186 254494
rect 29422 254258 29464 254494
rect 29144 247494 29464 254258
rect 29144 247258 29186 247494
rect 29422 247258 29464 247494
rect 29144 240494 29464 247258
rect 29144 240258 29186 240494
rect 29422 240258 29464 240494
rect 29144 233494 29464 240258
rect 29144 233258 29186 233494
rect 29422 233258 29464 233494
rect 29144 226494 29464 233258
rect 29144 226258 29186 226494
rect 29422 226258 29464 226494
rect 29144 219494 29464 226258
rect 29144 219258 29186 219494
rect 29422 219258 29464 219494
rect 29144 212494 29464 219258
rect 29144 212258 29186 212494
rect 29422 212258 29464 212494
rect 29144 205494 29464 212258
rect 29144 205258 29186 205494
rect 29422 205258 29464 205494
rect 29144 198494 29464 205258
rect 29144 198258 29186 198494
rect 29422 198258 29464 198494
rect 29144 191494 29464 198258
rect 29144 191258 29186 191494
rect 29422 191258 29464 191494
rect 29144 184494 29464 191258
rect 29144 184258 29186 184494
rect 29422 184258 29464 184494
rect 29144 177494 29464 184258
rect 29144 177258 29186 177494
rect 29422 177258 29464 177494
rect 29144 170494 29464 177258
rect 29144 170258 29186 170494
rect 29422 170258 29464 170494
rect 29144 163494 29464 170258
rect 29144 163258 29186 163494
rect 29422 163258 29464 163494
rect 29144 156494 29464 163258
rect 29144 156258 29186 156494
rect 29422 156258 29464 156494
rect 29144 149494 29464 156258
rect 29144 149258 29186 149494
rect 29422 149258 29464 149494
rect 29144 142494 29464 149258
rect 29144 142258 29186 142494
rect 29422 142258 29464 142494
rect 29144 135494 29464 142258
rect 29144 135258 29186 135494
rect 29422 135258 29464 135494
rect 29144 128494 29464 135258
rect 29144 128258 29186 128494
rect 29422 128258 29464 128494
rect 29144 121494 29464 128258
rect 29144 121258 29186 121494
rect 29422 121258 29464 121494
rect 29144 114494 29464 121258
rect 29144 114258 29186 114494
rect 29422 114258 29464 114494
rect 29144 107494 29464 114258
rect 29144 107258 29186 107494
rect 29422 107258 29464 107494
rect 29144 100494 29464 107258
rect 29144 100258 29186 100494
rect 29422 100258 29464 100494
rect 29144 93494 29464 100258
rect 29144 93258 29186 93494
rect 29422 93258 29464 93494
rect 29144 86494 29464 93258
rect 29144 86258 29186 86494
rect 29422 86258 29464 86494
rect 29144 79494 29464 86258
rect 29144 79258 29186 79494
rect 29422 79258 29464 79494
rect 29144 72494 29464 79258
rect 29144 72258 29186 72494
rect 29422 72258 29464 72494
rect 29144 65494 29464 72258
rect 29144 65258 29186 65494
rect 29422 65258 29464 65494
rect 29144 58494 29464 65258
rect 29144 58258 29186 58494
rect 29422 58258 29464 58494
rect 29144 51494 29464 58258
rect 29144 51258 29186 51494
rect 29422 51258 29464 51494
rect 29144 44494 29464 51258
rect 29144 44258 29186 44494
rect 29422 44258 29464 44494
rect 29144 37494 29464 44258
rect 29144 37258 29186 37494
rect 29422 37258 29464 37494
rect 29144 30494 29464 37258
rect 29144 30258 29186 30494
rect 29422 30258 29464 30494
rect 29144 23494 29464 30258
rect 29144 23258 29186 23494
rect 29422 23258 29464 23494
rect 29144 16494 29464 23258
rect 29144 16258 29186 16494
rect 29422 16258 29464 16494
rect 29144 9494 29464 16258
rect 29144 9258 29186 9494
rect 29422 9258 29464 9494
rect 29144 2494 29464 9258
rect 29144 2258 29186 2494
rect 29422 2258 29464 2494
rect 29144 -746 29464 2258
rect 29144 -982 29186 -746
rect 29422 -982 29464 -746
rect 29144 -1066 29464 -982
rect 29144 -1302 29186 -1066
rect 29422 -1302 29464 -1066
rect 29144 -2294 29464 -1302
rect 30876 706198 31196 706230
rect 30876 705962 30918 706198
rect 31154 705962 31196 706198
rect 30876 705878 31196 705962
rect 30876 705642 30918 705878
rect 31154 705642 31196 705878
rect 30876 696561 31196 705642
rect 30876 696325 30918 696561
rect 31154 696325 31196 696561
rect 30876 689561 31196 696325
rect 30876 689325 30918 689561
rect 31154 689325 31196 689561
rect 30876 682561 31196 689325
rect 30876 682325 30918 682561
rect 31154 682325 31196 682561
rect 30876 675561 31196 682325
rect 30876 675325 30918 675561
rect 31154 675325 31196 675561
rect 30876 668561 31196 675325
rect 30876 668325 30918 668561
rect 31154 668325 31196 668561
rect 30876 661561 31196 668325
rect 30876 661325 30918 661561
rect 31154 661325 31196 661561
rect 30876 654561 31196 661325
rect 30876 654325 30918 654561
rect 31154 654325 31196 654561
rect 30876 647561 31196 654325
rect 30876 647325 30918 647561
rect 31154 647325 31196 647561
rect 30876 640561 31196 647325
rect 30876 640325 30918 640561
rect 31154 640325 31196 640561
rect 30876 633561 31196 640325
rect 30876 633325 30918 633561
rect 31154 633325 31196 633561
rect 30876 626561 31196 633325
rect 30876 626325 30918 626561
rect 31154 626325 31196 626561
rect 30876 619561 31196 626325
rect 30876 619325 30918 619561
rect 31154 619325 31196 619561
rect 30876 612561 31196 619325
rect 30876 612325 30918 612561
rect 31154 612325 31196 612561
rect 30876 605561 31196 612325
rect 30876 605325 30918 605561
rect 31154 605325 31196 605561
rect 30876 598561 31196 605325
rect 30876 598325 30918 598561
rect 31154 598325 31196 598561
rect 30876 591561 31196 598325
rect 30876 591325 30918 591561
rect 31154 591325 31196 591561
rect 30876 584561 31196 591325
rect 30876 584325 30918 584561
rect 31154 584325 31196 584561
rect 30876 577561 31196 584325
rect 30876 577325 30918 577561
rect 31154 577325 31196 577561
rect 30876 570561 31196 577325
rect 30876 570325 30918 570561
rect 31154 570325 31196 570561
rect 30876 563561 31196 570325
rect 30876 563325 30918 563561
rect 31154 563325 31196 563561
rect 30876 556561 31196 563325
rect 30876 556325 30918 556561
rect 31154 556325 31196 556561
rect 30876 549561 31196 556325
rect 30876 549325 30918 549561
rect 31154 549325 31196 549561
rect 30876 542561 31196 549325
rect 30876 542325 30918 542561
rect 31154 542325 31196 542561
rect 30876 535561 31196 542325
rect 30876 535325 30918 535561
rect 31154 535325 31196 535561
rect 30876 528561 31196 535325
rect 30876 528325 30918 528561
rect 31154 528325 31196 528561
rect 30876 521561 31196 528325
rect 30876 521325 30918 521561
rect 31154 521325 31196 521561
rect 30876 514561 31196 521325
rect 30876 514325 30918 514561
rect 31154 514325 31196 514561
rect 30876 507561 31196 514325
rect 30876 507325 30918 507561
rect 31154 507325 31196 507561
rect 30876 500561 31196 507325
rect 30876 500325 30918 500561
rect 31154 500325 31196 500561
rect 30876 493561 31196 500325
rect 30876 493325 30918 493561
rect 31154 493325 31196 493561
rect 30876 486561 31196 493325
rect 30876 486325 30918 486561
rect 31154 486325 31196 486561
rect 30876 479561 31196 486325
rect 30876 479325 30918 479561
rect 31154 479325 31196 479561
rect 30876 472561 31196 479325
rect 30876 472325 30918 472561
rect 31154 472325 31196 472561
rect 30876 465561 31196 472325
rect 30876 465325 30918 465561
rect 31154 465325 31196 465561
rect 30876 458561 31196 465325
rect 30876 458325 30918 458561
rect 31154 458325 31196 458561
rect 30876 451561 31196 458325
rect 30876 451325 30918 451561
rect 31154 451325 31196 451561
rect 30876 444561 31196 451325
rect 30876 444325 30918 444561
rect 31154 444325 31196 444561
rect 30876 437561 31196 444325
rect 30876 437325 30918 437561
rect 31154 437325 31196 437561
rect 30876 430561 31196 437325
rect 30876 430325 30918 430561
rect 31154 430325 31196 430561
rect 30876 423561 31196 430325
rect 30876 423325 30918 423561
rect 31154 423325 31196 423561
rect 30876 416561 31196 423325
rect 30876 416325 30918 416561
rect 31154 416325 31196 416561
rect 30876 409561 31196 416325
rect 30876 409325 30918 409561
rect 31154 409325 31196 409561
rect 30876 402561 31196 409325
rect 30876 402325 30918 402561
rect 31154 402325 31196 402561
rect 30876 395561 31196 402325
rect 30876 395325 30918 395561
rect 31154 395325 31196 395561
rect 30876 388561 31196 395325
rect 30876 388325 30918 388561
rect 31154 388325 31196 388561
rect 30876 381561 31196 388325
rect 30876 381325 30918 381561
rect 31154 381325 31196 381561
rect 30876 374561 31196 381325
rect 30876 374325 30918 374561
rect 31154 374325 31196 374561
rect 30876 367561 31196 374325
rect 30876 367325 30918 367561
rect 31154 367325 31196 367561
rect 30876 360561 31196 367325
rect 30876 360325 30918 360561
rect 31154 360325 31196 360561
rect 30876 353561 31196 360325
rect 30876 353325 30918 353561
rect 31154 353325 31196 353561
rect 30876 346561 31196 353325
rect 30876 346325 30918 346561
rect 31154 346325 31196 346561
rect 30876 339561 31196 346325
rect 30876 339325 30918 339561
rect 31154 339325 31196 339561
rect 30876 332561 31196 339325
rect 30876 332325 30918 332561
rect 31154 332325 31196 332561
rect 30876 325561 31196 332325
rect 30876 325325 30918 325561
rect 31154 325325 31196 325561
rect 30876 318561 31196 325325
rect 30876 318325 30918 318561
rect 31154 318325 31196 318561
rect 30876 311561 31196 318325
rect 30876 311325 30918 311561
rect 31154 311325 31196 311561
rect 30876 304561 31196 311325
rect 30876 304325 30918 304561
rect 31154 304325 31196 304561
rect 30876 297561 31196 304325
rect 30876 297325 30918 297561
rect 31154 297325 31196 297561
rect 30876 290561 31196 297325
rect 30876 290325 30918 290561
rect 31154 290325 31196 290561
rect 30876 283561 31196 290325
rect 30876 283325 30918 283561
rect 31154 283325 31196 283561
rect 30876 276561 31196 283325
rect 30876 276325 30918 276561
rect 31154 276325 31196 276561
rect 30876 269561 31196 276325
rect 30876 269325 30918 269561
rect 31154 269325 31196 269561
rect 30876 262561 31196 269325
rect 30876 262325 30918 262561
rect 31154 262325 31196 262561
rect 30876 255561 31196 262325
rect 30876 255325 30918 255561
rect 31154 255325 31196 255561
rect 30876 248561 31196 255325
rect 30876 248325 30918 248561
rect 31154 248325 31196 248561
rect 30876 241561 31196 248325
rect 30876 241325 30918 241561
rect 31154 241325 31196 241561
rect 30876 234561 31196 241325
rect 30876 234325 30918 234561
rect 31154 234325 31196 234561
rect 30876 227561 31196 234325
rect 30876 227325 30918 227561
rect 31154 227325 31196 227561
rect 30876 220561 31196 227325
rect 30876 220325 30918 220561
rect 31154 220325 31196 220561
rect 30876 213561 31196 220325
rect 30876 213325 30918 213561
rect 31154 213325 31196 213561
rect 30876 206561 31196 213325
rect 30876 206325 30918 206561
rect 31154 206325 31196 206561
rect 30876 199561 31196 206325
rect 30876 199325 30918 199561
rect 31154 199325 31196 199561
rect 30876 192561 31196 199325
rect 30876 192325 30918 192561
rect 31154 192325 31196 192561
rect 30876 185561 31196 192325
rect 30876 185325 30918 185561
rect 31154 185325 31196 185561
rect 30876 178561 31196 185325
rect 30876 178325 30918 178561
rect 31154 178325 31196 178561
rect 30876 171561 31196 178325
rect 30876 171325 30918 171561
rect 31154 171325 31196 171561
rect 30876 164561 31196 171325
rect 30876 164325 30918 164561
rect 31154 164325 31196 164561
rect 30876 157561 31196 164325
rect 30876 157325 30918 157561
rect 31154 157325 31196 157561
rect 30876 150561 31196 157325
rect 30876 150325 30918 150561
rect 31154 150325 31196 150561
rect 30876 143561 31196 150325
rect 30876 143325 30918 143561
rect 31154 143325 31196 143561
rect 30876 136561 31196 143325
rect 30876 136325 30918 136561
rect 31154 136325 31196 136561
rect 30876 129561 31196 136325
rect 30876 129325 30918 129561
rect 31154 129325 31196 129561
rect 30876 122561 31196 129325
rect 30876 122325 30918 122561
rect 31154 122325 31196 122561
rect 30876 115561 31196 122325
rect 30876 115325 30918 115561
rect 31154 115325 31196 115561
rect 30876 108561 31196 115325
rect 30876 108325 30918 108561
rect 31154 108325 31196 108561
rect 30876 101561 31196 108325
rect 30876 101325 30918 101561
rect 31154 101325 31196 101561
rect 30876 94561 31196 101325
rect 30876 94325 30918 94561
rect 31154 94325 31196 94561
rect 30876 87561 31196 94325
rect 30876 87325 30918 87561
rect 31154 87325 31196 87561
rect 30876 80561 31196 87325
rect 30876 80325 30918 80561
rect 31154 80325 31196 80561
rect 30876 73561 31196 80325
rect 30876 73325 30918 73561
rect 31154 73325 31196 73561
rect 30876 66561 31196 73325
rect 30876 66325 30918 66561
rect 31154 66325 31196 66561
rect 30876 59561 31196 66325
rect 30876 59325 30918 59561
rect 31154 59325 31196 59561
rect 30876 52561 31196 59325
rect 30876 52325 30918 52561
rect 31154 52325 31196 52561
rect 30876 45561 31196 52325
rect 30876 45325 30918 45561
rect 31154 45325 31196 45561
rect 30876 38561 31196 45325
rect 30876 38325 30918 38561
rect 31154 38325 31196 38561
rect 30876 31561 31196 38325
rect 30876 31325 30918 31561
rect 31154 31325 31196 31561
rect 30876 24561 31196 31325
rect 30876 24325 30918 24561
rect 31154 24325 31196 24561
rect 30876 17561 31196 24325
rect 30876 17325 30918 17561
rect 31154 17325 31196 17561
rect 30876 10561 31196 17325
rect 30876 10325 30918 10561
rect 31154 10325 31196 10561
rect 30876 3561 31196 10325
rect 30876 3325 30918 3561
rect 31154 3325 31196 3561
rect 30876 -1706 31196 3325
rect 30876 -1942 30918 -1706
rect 31154 -1942 31196 -1706
rect 30876 -2026 31196 -1942
rect 30876 -2262 30918 -2026
rect 31154 -2262 31196 -2026
rect 30876 -2294 31196 -2262
rect 36144 705238 36464 706230
rect 36144 705002 36186 705238
rect 36422 705002 36464 705238
rect 36144 704918 36464 705002
rect 36144 704682 36186 704918
rect 36422 704682 36464 704918
rect 36144 695494 36464 704682
rect 36144 695258 36186 695494
rect 36422 695258 36464 695494
rect 36144 688494 36464 695258
rect 36144 688258 36186 688494
rect 36422 688258 36464 688494
rect 36144 681494 36464 688258
rect 36144 681258 36186 681494
rect 36422 681258 36464 681494
rect 36144 674494 36464 681258
rect 36144 674258 36186 674494
rect 36422 674258 36464 674494
rect 36144 667494 36464 674258
rect 36144 667258 36186 667494
rect 36422 667258 36464 667494
rect 36144 660494 36464 667258
rect 36144 660258 36186 660494
rect 36422 660258 36464 660494
rect 36144 653494 36464 660258
rect 36144 653258 36186 653494
rect 36422 653258 36464 653494
rect 36144 646494 36464 653258
rect 36144 646258 36186 646494
rect 36422 646258 36464 646494
rect 36144 639494 36464 646258
rect 36144 639258 36186 639494
rect 36422 639258 36464 639494
rect 36144 632494 36464 639258
rect 36144 632258 36186 632494
rect 36422 632258 36464 632494
rect 36144 625494 36464 632258
rect 36144 625258 36186 625494
rect 36422 625258 36464 625494
rect 36144 618494 36464 625258
rect 36144 618258 36186 618494
rect 36422 618258 36464 618494
rect 36144 611494 36464 618258
rect 36144 611258 36186 611494
rect 36422 611258 36464 611494
rect 36144 604494 36464 611258
rect 36144 604258 36186 604494
rect 36422 604258 36464 604494
rect 36144 597494 36464 604258
rect 36144 597258 36186 597494
rect 36422 597258 36464 597494
rect 36144 590494 36464 597258
rect 36144 590258 36186 590494
rect 36422 590258 36464 590494
rect 36144 583494 36464 590258
rect 36144 583258 36186 583494
rect 36422 583258 36464 583494
rect 36144 576494 36464 583258
rect 36144 576258 36186 576494
rect 36422 576258 36464 576494
rect 36144 569494 36464 576258
rect 36144 569258 36186 569494
rect 36422 569258 36464 569494
rect 36144 562494 36464 569258
rect 36144 562258 36186 562494
rect 36422 562258 36464 562494
rect 36144 555494 36464 562258
rect 36144 555258 36186 555494
rect 36422 555258 36464 555494
rect 36144 548494 36464 555258
rect 36144 548258 36186 548494
rect 36422 548258 36464 548494
rect 36144 541494 36464 548258
rect 36144 541258 36186 541494
rect 36422 541258 36464 541494
rect 36144 534494 36464 541258
rect 36144 534258 36186 534494
rect 36422 534258 36464 534494
rect 36144 527494 36464 534258
rect 36144 527258 36186 527494
rect 36422 527258 36464 527494
rect 36144 520494 36464 527258
rect 36144 520258 36186 520494
rect 36422 520258 36464 520494
rect 36144 513494 36464 520258
rect 36144 513258 36186 513494
rect 36422 513258 36464 513494
rect 36144 506494 36464 513258
rect 36144 506258 36186 506494
rect 36422 506258 36464 506494
rect 36144 499494 36464 506258
rect 36144 499258 36186 499494
rect 36422 499258 36464 499494
rect 36144 492494 36464 499258
rect 36144 492258 36186 492494
rect 36422 492258 36464 492494
rect 36144 485494 36464 492258
rect 36144 485258 36186 485494
rect 36422 485258 36464 485494
rect 36144 478494 36464 485258
rect 36144 478258 36186 478494
rect 36422 478258 36464 478494
rect 36144 471494 36464 478258
rect 36144 471258 36186 471494
rect 36422 471258 36464 471494
rect 36144 464494 36464 471258
rect 36144 464258 36186 464494
rect 36422 464258 36464 464494
rect 36144 457494 36464 464258
rect 36144 457258 36186 457494
rect 36422 457258 36464 457494
rect 36144 450494 36464 457258
rect 36144 450258 36186 450494
rect 36422 450258 36464 450494
rect 36144 443494 36464 450258
rect 36144 443258 36186 443494
rect 36422 443258 36464 443494
rect 36144 436494 36464 443258
rect 36144 436258 36186 436494
rect 36422 436258 36464 436494
rect 36144 429494 36464 436258
rect 36144 429258 36186 429494
rect 36422 429258 36464 429494
rect 36144 422494 36464 429258
rect 36144 422258 36186 422494
rect 36422 422258 36464 422494
rect 36144 415494 36464 422258
rect 36144 415258 36186 415494
rect 36422 415258 36464 415494
rect 36144 408494 36464 415258
rect 36144 408258 36186 408494
rect 36422 408258 36464 408494
rect 36144 401494 36464 408258
rect 36144 401258 36186 401494
rect 36422 401258 36464 401494
rect 36144 394494 36464 401258
rect 36144 394258 36186 394494
rect 36422 394258 36464 394494
rect 36144 387494 36464 394258
rect 36144 387258 36186 387494
rect 36422 387258 36464 387494
rect 36144 380494 36464 387258
rect 36144 380258 36186 380494
rect 36422 380258 36464 380494
rect 36144 373494 36464 380258
rect 36144 373258 36186 373494
rect 36422 373258 36464 373494
rect 36144 366494 36464 373258
rect 36144 366258 36186 366494
rect 36422 366258 36464 366494
rect 36144 359494 36464 366258
rect 36144 359258 36186 359494
rect 36422 359258 36464 359494
rect 36144 352494 36464 359258
rect 36144 352258 36186 352494
rect 36422 352258 36464 352494
rect 36144 345494 36464 352258
rect 36144 345258 36186 345494
rect 36422 345258 36464 345494
rect 36144 338494 36464 345258
rect 36144 338258 36186 338494
rect 36422 338258 36464 338494
rect 36144 331494 36464 338258
rect 36144 331258 36186 331494
rect 36422 331258 36464 331494
rect 36144 324494 36464 331258
rect 36144 324258 36186 324494
rect 36422 324258 36464 324494
rect 36144 317494 36464 324258
rect 36144 317258 36186 317494
rect 36422 317258 36464 317494
rect 36144 310494 36464 317258
rect 36144 310258 36186 310494
rect 36422 310258 36464 310494
rect 36144 303494 36464 310258
rect 36144 303258 36186 303494
rect 36422 303258 36464 303494
rect 36144 296494 36464 303258
rect 36144 296258 36186 296494
rect 36422 296258 36464 296494
rect 36144 289494 36464 296258
rect 36144 289258 36186 289494
rect 36422 289258 36464 289494
rect 36144 282494 36464 289258
rect 36144 282258 36186 282494
rect 36422 282258 36464 282494
rect 36144 275494 36464 282258
rect 36144 275258 36186 275494
rect 36422 275258 36464 275494
rect 36144 268494 36464 275258
rect 36144 268258 36186 268494
rect 36422 268258 36464 268494
rect 36144 261494 36464 268258
rect 36144 261258 36186 261494
rect 36422 261258 36464 261494
rect 36144 254494 36464 261258
rect 36144 254258 36186 254494
rect 36422 254258 36464 254494
rect 36144 247494 36464 254258
rect 36144 247258 36186 247494
rect 36422 247258 36464 247494
rect 36144 240494 36464 247258
rect 36144 240258 36186 240494
rect 36422 240258 36464 240494
rect 36144 233494 36464 240258
rect 36144 233258 36186 233494
rect 36422 233258 36464 233494
rect 36144 226494 36464 233258
rect 36144 226258 36186 226494
rect 36422 226258 36464 226494
rect 36144 219494 36464 226258
rect 36144 219258 36186 219494
rect 36422 219258 36464 219494
rect 36144 212494 36464 219258
rect 36144 212258 36186 212494
rect 36422 212258 36464 212494
rect 36144 205494 36464 212258
rect 36144 205258 36186 205494
rect 36422 205258 36464 205494
rect 36144 198494 36464 205258
rect 36144 198258 36186 198494
rect 36422 198258 36464 198494
rect 36144 191494 36464 198258
rect 36144 191258 36186 191494
rect 36422 191258 36464 191494
rect 36144 184494 36464 191258
rect 36144 184258 36186 184494
rect 36422 184258 36464 184494
rect 36144 177494 36464 184258
rect 36144 177258 36186 177494
rect 36422 177258 36464 177494
rect 36144 170494 36464 177258
rect 36144 170258 36186 170494
rect 36422 170258 36464 170494
rect 36144 163494 36464 170258
rect 36144 163258 36186 163494
rect 36422 163258 36464 163494
rect 36144 156494 36464 163258
rect 36144 156258 36186 156494
rect 36422 156258 36464 156494
rect 36144 149494 36464 156258
rect 36144 149258 36186 149494
rect 36422 149258 36464 149494
rect 36144 142494 36464 149258
rect 36144 142258 36186 142494
rect 36422 142258 36464 142494
rect 36144 135494 36464 142258
rect 36144 135258 36186 135494
rect 36422 135258 36464 135494
rect 36144 128494 36464 135258
rect 36144 128258 36186 128494
rect 36422 128258 36464 128494
rect 36144 121494 36464 128258
rect 36144 121258 36186 121494
rect 36422 121258 36464 121494
rect 36144 114494 36464 121258
rect 36144 114258 36186 114494
rect 36422 114258 36464 114494
rect 36144 107494 36464 114258
rect 36144 107258 36186 107494
rect 36422 107258 36464 107494
rect 36144 100494 36464 107258
rect 36144 100258 36186 100494
rect 36422 100258 36464 100494
rect 36144 93494 36464 100258
rect 36144 93258 36186 93494
rect 36422 93258 36464 93494
rect 36144 86494 36464 93258
rect 36144 86258 36186 86494
rect 36422 86258 36464 86494
rect 36144 79494 36464 86258
rect 36144 79258 36186 79494
rect 36422 79258 36464 79494
rect 36144 72494 36464 79258
rect 36144 72258 36186 72494
rect 36422 72258 36464 72494
rect 36144 65494 36464 72258
rect 36144 65258 36186 65494
rect 36422 65258 36464 65494
rect 36144 58494 36464 65258
rect 36144 58258 36186 58494
rect 36422 58258 36464 58494
rect 36144 51494 36464 58258
rect 36144 51258 36186 51494
rect 36422 51258 36464 51494
rect 36144 44494 36464 51258
rect 36144 44258 36186 44494
rect 36422 44258 36464 44494
rect 36144 37494 36464 44258
rect 36144 37258 36186 37494
rect 36422 37258 36464 37494
rect 36144 30494 36464 37258
rect 36144 30258 36186 30494
rect 36422 30258 36464 30494
rect 36144 23494 36464 30258
rect 36144 23258 36186 23494
rect 36422 23258 36464 23494
rect 36144 16494 36464 23258
rect 36144 16258 36186 16494
rect 36422 16258 36464 16494
rect 36144 9494 36464 16258
rect 36144 9258 36186 9494
rect 36422 9258 36464 9494
rect 36144 2494 36464 9258
rect 36144 2258 36186 2494
rect 36422 2258 36464 2494
rect 36144 -746 36464 2258
rect 36144 -982 36186 -746
rect 36422 -982 36464 -746
rect 36144 -1066 36464 -982
rect 36144 -1302 36186 -1066
rect 36422 -1302 36464 -1066
rect 36144 -2294 36464 -1302
rect 37876 706198 38196 706230
rect 37876 705962 37918 706198
rect 38154 705962 38196 706198
rect 37876 705878 38196 705962
rect 37876 705642 37918 705878
rect 38154 705642 38196 705878
rect 37876 696561 38196 705642
rect 37876 696325 37918 696561
rect 38154 696325 38196 696561
rect 37876 689561 38196 696325
rect 37876 689325 37918 689561
rect 38154 689325 38196 689561
rect 37876 682561 38196 689325
rect 37876 682325 37918 682561
rect 38154 682325 38196 682561
rect 37876 675561 38196 682325
rect 37876 675325 37918 675561
rect 38154 675325 38196 675561
rect 37876 668561 38196 675325
rect 37876 668325 37918 668561
rect 38154 668325 38196 668561
rect 37876 661561 38196 668325
rect 37876 661325 37918 661561
rect 38154 661325 38196 661561
rect 37876 654561 38196 661325
rect 37876 654325 37918 654561
rect 38154 654325 38196 654561
rect 37876 647561 38196 654325
rect 37876 647325 37918 647561
rect 38154 647325 38196 647561
rect 37876 640561 38196 647325
rect 37876 640325 37918 640561
rect 38154 640325 38196 640561
rect 37876 633561 38196 640325
rect 37876 633325 37918 633561
rect 38154 633325 38196 633561
rect 37876 626561 38196 633325
rect 37876 626325 37918 626561
rect 38154 626325 38196 626561
rect 37876 619561 38196 626325
rect 37876 619325 37918 619561
rect 38154 619325 38196 619561
rect 37876 612561 38196 619325
rect 37876 612325 37918 612561
rect 38154 612325 38196 612561
rect 37876 605561 38196 612325
rect 37876 605325 37918 605561
rect 38154 605325 38196 605561
rect 37876 598561 38196 605325
rect 37876 598325 37918 598561
rect 38154 598325 38196 598561
rect 37876 591561 38196 598325
rect 37876 591325 37918 591561
rect 38154 591325 38196 591561
rect 37876 584561 38196 591325
rect 37876 584325 37918 584561
rect 38154 584325 38196 584561
rect 37876 577561 38196 584325
rect 37876 577325 37918 577561
rect 38154 577325 38196 577561
rect 37876 570561 38196 577325
rect 37876 570325 37918 570561
rect 38154 570325 38196 570561
rect 37876 563561 38196 570325
rect 37876 563325 37918 563561
rect 38154 563325 38196 563561
rect 37876 556561 38196 563325
rect 37876 556325 37918 556561
rect 38154 556325 38196 556561
rect 37876 549561 38196 556325
rect 37876 549325 37918 549561
rect 38154 549325 38196 549561
rect 37876 542561 38196 549325
rect 37876 542325 37918 542561
rect 38154 542325 38196 542561
rect 37876 535561 38196 542325
rect 37876 535325 37918 535561
rect 38154 535325 38196 535561
rect 37876 528561 38196 535325
rect 37876 528325 37918 528561
rect 38154 528325 38196 528561
rect 37876 521561 38196 528325
rect 37876 521325 37918 521561
rect 38154 521325 38196 521561
rect 37876 514561 38196 521325
rect 37876 514325 37918 514561
rect 38154 514325 38196 514561
rect 37876 507561 38196 514325
rect 37876 507325 37918 507561
rect 38154 507325 38196 507561
rect 37876 500561 38196 507325
rect 37876 500325 37918 500561
rect 38154 500325 38196 500561
rect 37876 493561 38196 500325
rect 37876 493325 37918 493561
rect 38154 493325 38196 493561
rect 37876 486561 38196 493325
rect 37876 486325 37918 486561
rect 38154 486325 38196 486561
rect 37876 479561 38196 486325
rect 37876 479325 37918 479561
rect 38154 479325 38196 479561
rect 37876 472561 38196 479325
rect 37876 472325 37918 472561
rect 38154 472325 38196 472561
rect 37876 465561 38196 472325
rect 37876 465325 37918 465561
rect 38154 465325 38196 465561
rect 37876 458561 38196 465325
rect 37876 458325 37918 458561
rect 38154 458325 38196 458561
rect 37876 451561 38196 458325
rect 37876 451325 37918 451561
rect 38154 451325 38196 451561
rect 37876 444561 38196 451325
rect 37876 444325 37918 444561
rect 38154 444325 38196 444561
rect 37876 437561 38196 444325
rect 37876 437325 37918 437561
rect 38154 437325 38196 437561
rect 37876 430561 38196 437325
rect 37876 430325 37918 430561
rect 38154 430325 38196 430561
rect 37876 423561 38196 430325
rect 37876 423325 37918 423561
rect 38154 423325 38196 423561
rect 37876 416561 38196 423325
rect 37876 416325 37918 416561
rect 38154 416325 38196 416561
rect 37876 409561 38196 416325
rect 37876 409325 37918 409561
rect 38154 409325 38196 409561
rect 37876 402561 38196 409325
rect 37876 402325 37918 402561
rect 38154 402325 38196 402561
rect 37876 395561 38196 402325
rect 37876 395325 37918 395561
rect 38154 395325 38196 395561
rect 37876 388561 38196 395325
rect 37876 388325 37918 388561
rect 38154 388325 38196 388561
rect 37876 381561 38196 388325
rect 37876 381325 37918 381561
rect 38154 381325 38196 381561
rect 37876 374561 38196 381325
rect 37876 374325 37918 374561
rect 38154 374325 38196 374561
rect 37876 367561 38196 374325
rect 37876 367325 37918 367561
rect 38154 367325 38196 367561
rect 37876 360561 38196 367325
rect 37876 360325 37918 360561
rect 38154 360325 38196 360561
rect 37876 353561 38196 360325
rect 37876 353325 37918 353561
rect 38154 353325 38196 353561
rect 37876 346561 38196 353325
rect 37876 346325 37918 346561
rect 38154 346325 38196 346561
rect 37876 339561 38196 346325
rect 37876 339325 37918 339561
rect 38154 339325 38196 339561
rect 37876 332561 38196 339325
rect 37876 332325 37918 332561
rect 38154 332325 38196 332561
rect 37876 325561 38196 332325
rect 37876 325325 37918 325561
rect 38154 325325 38196 325561
rect 37876 318561 38196 325325
rect 37876 318325 37918 318561
rect 38154 318325 38196 318561
rect 37876 311561 38196 318325
rect 37876 311325 37918 311561
rect 38154 311325 38196 311561
rect 37876 304561 38196 311325
rect 37876 304325 37918 304561
rect 38154 304325 38196 304561
rect 37876 297561 38196 304325
rect 37876 297325 37918 297561
rect 38154 297325 38196 297561
rect 37876 290561 38196 297325
rect 37876 290325 37918 290561
rect 38154 290325 38196 290561
rect 37876 283561 38196 290325
rect 37876 283325 37918 283561
rect 38154 283325 38196 283561
rect 37876 276561 38196 283325
rect 37876 276325 37918 276561
rect 38154 276325 38196 276561
rect 37876 269561 38196 276325
rect 37876 269325 37918 269561
rect 38154 269325 38196 269561
rect 37876 262561 38196 269325
rect 37876 262325 37918 262561
rect 38154 262325 38196 262561
rect 37876 255561 38196 262325
rect 37876 255325 37918 255561
rect 38154 255325 38196 255561
rect 37876 248561 38196 255325
rect 37876 248325 37918 248561
rect 38154 248325 38196 248561
rect 37876 241561 38196 248325
rect 37876 241325 37918 241561
rect 38154 241325 38196 241561
rect 37876 234561 38196 241325
rect 37876 234325 37918 234561
rect 38154 234325 38196 234561
rect 37876 227561 38196 234325
rect 37876 227325 37918 227561
rect 38154 227325 38196 227561
rect 37876 220561 38196 227325
rect 37876 220325 37918 220561
rect 38154 220325 38196 220561
rect 37876 213561 38196 220325
rect 37876 213325 37918 213561
rect 38154 213325 38196 213561
rect 37876 206561 38196 213325
rect 37876 206325 37918 206561
rect 38154 206325 38196 206561
rect 37876 199561 38196 206325
rect 37876 199325 37918 199561
rect 38154 199325 38196 199561
rect 37876 192561 38196 199325
rect 37876 192325 37918 192561
rect 38154 192325 38196 192561
rect 37876 185561 38196 192325
rect 37876 185325 37918 185561
rect 38154 185325 38196 185561
rect 37876 178561 38196 185325
rect 37876 178325 37918 178561
rect 38154 178325 38196 178561
rect 37876 171561 38196 178325
rect 37876 171325 37918 171561
rect 38154 171325 38196 171561
rect 37876 164561 38196 171325
rect 37876 164325 37918 164561
rect 38154 164325 38196 164561
rect 37876 157561 38196 164325
rect 37876 157325 37918 157561
rect 38154 157325 38196 157561
rect 37876 150561 38196 157325
rect 37876 150325 37918 150561
rect 38154 150325 38196 150561
rect 37876 143561 38196 150325
rect 37876 143325 37918 143561
rect 38154 143325 38196 143561
rect 37876 136561 38196 143325
rect 37876 136325 37918 136561
rect 38154 136325 38196 136561
rect 37876 129561 38196 136325
rect 37876 129325 37918 129561
rect 38154 129325 38196 129561
rect 37876 122561 38196 129325
rect 37876 122325 37918 122561
rect 38154 122325 38196 122561
rect 37876 115561 38196 122325
rect 37876 115325 37918 115561
rect 38154 115325 38196 115561
rect 37876 108561 38196 115325
rect 37876 108325 37918 108561
rect 38154 108325 38196 108561
rect 37876 101561 38196 108325
rect 37876 101325 37918 101561
rect 38154 101325 38196 101561
rect 37876 94561 38196 101325
rect 37876 94325 37918 94561
rect 38154 94325 38196 94561
rect 37876 87561 38196 94325
rect 37876 87325 37918 87561
rect 38154 87325 38196 87561
rect 37876 80561 38196 87325
rect 37876 80325 37918 80561
rect 38154 80325 38196 80561
rect 37876 73561 38196 80325
rect 37876 73325 37918 73561
rect 38154 73325 38196 73561
rect 37876 66561 38196 73325
rect 37876 66325 37918 66561
rect 38154 66325 38196 66561
rect 37876 59561 38196 66325
rect 37876 59325 37918 59561
rect 38154 59325 38196 59561
rect 37876 52561 38196 59325
rect 37876 52325 37918 52561
rect 38154 52325 38196 52561
rect 37876 45561 38196 52325
rect 37876 45325 37918 45561
rect 38154 45325 38196 45561
rect 37876 38561 38196 45325
rect 37876 38325 37918 38561
rect 38154 38325 38196 38561
rect 37876 31561 38196 38325
rect 37876 31325 37918 31561
rect 38154 31325 38196 31561
rect 37876 24561 38196 31325
rect 37876 24325 37918 24561
rect 38154 24325 38196 24561
rect 37876 17561 38196 24325
rect 37876 17325 37918 17561
rect 38154 17325 38196 17561
rect 37876 10561 38196 17325
rect 37876 10325 37918 10561
rect 38154 10325 38196 10561
rect 37876 3561 38196 10325
rect 37876 3325 37918 3561
rect 38154 3325 38196 3561
rect 37876 -1706 38196 3325
rect 37876 -1942 37918 -1706
rect 38154 -1942 38196 -1706
rect 37876 -2026 38196 -1942
rect 37876 -2262 37918 -2026
rect 38154 -2262 38196 -2026
rect 37876 -2294 38196 -2262
rect 43144 705238 43464 706230
rect 43144 705002 43186 705238
rect 43422 705002 43464 705238
rect 43144 704918 43464 705002
rect 43144 704682 43186 704918
rect 43422 704682 43464 704918
rect 43144 695494 43464 704682
rect 43144 695258 43186 695494
rect 43422 695258 43464 695494
rect 43144 688494 43464 695258
rect 43144 688258 43186 688494
rect 43422 688258 43464 688494
rect 43144 681494 43464 688258
rect 43144 681258 43186 681494
rect 43422 681258 43464 681494
rect 43144 674494 43464 681258
rect 43144 674258 43186 674494
rect 43422 674258 43464 674494
rect 43144 667494 43464 674258
rect 43144 667258 43186 667494
rect 43422 667258 43464 667494
rect 43144 660494 43464 667258
rect 43144 660258 43186 660494
rect 43422 660258 43464 660494
rect 43144 653494 43464 660258
rect 43144 653258 43186 653494
rect 43422 653258 43464 653494
rect 43144 646494 43464 653258
rect 43144 646258 43186 646494
rect 43422 646258 43464 646494
rect 43144 639494 43464 646258
rect 43144 639258 43186 639494
rect 43422 639258 43464 639494
rect 43144 632494 43464 639258
rect 43144 632258 43186 632494
rect 43422 632258 43464 632494
rect 43144 625494 43464 632258
rect 43144 625258 43186 625494
rect 43422 625258 43464 625494
rect 43144 618494 43464 625258
rect 43144 618258 43186 618494
rect 43422 618258 43464 618494
rect 43144 611494 43464 618258
rect 43144 611258 43186 611494
rect 43422 611258 43464 611494
rect 43144 604494 43464 611258
rect 43144 604258 43186 604494
rect 43422 604258 43464 604494
rect 43144 597494 43464 604258
rect 43144 597258 43186 597494
rect 43422 597258 43464 597494
rect 43144 590494 43464 597258
rect 43144 590258 43186 590494
rect 43422 590258 43464 590494
rect 43144 583494 43464 590258
rect 43144 583258 43186 583494
rect 43422 583258 43464 583494
rect 43144 576494 43464 583258
rect 43144 576258 43186 576494
rect 43422 576258 43464 576494
rect 43144 569494 43464 576258
rect 43144 569258 43186 569494
rect 43422 569258 43464 569494
rect 43144 562494 43464 569258
rect 43144 562258 43186 562494
rect 43422 562258 43464 562494
rect 43144 555494 43464 562258
rect 43144 555258 43186 555494
rect 43422 555258 43464 555494
rect 43144 548494 43464 555258
rect 43144 548258 43186 548494
rect 43422 548258 43464 548494
rect 43144 541494 43464 548258
rect 43144 541258 43186 541494
rect 43422 541258 43464 541494
rect 43144 534494 43464 541258
rect 43144 534258 43186 534494
rect 43422 534258 43464 534494
rect 43144 527494 43464 534258
rect 43144 527258 43186 527494
rect 43422 527258 43464 527494
rect 43144 520494 43464 527258
rect 43144 520258 43186 520494
rect 43422 520258 43464 520494
rect 43144 513494 43464 520258
rect 43144 513258 43186 513494
rect 43422 513258 43464 513494
rect 43144 506494 43464 513258
rect 43144 506258 43186 506494
rect 43422 506258 43464 506494
rect 43144 499494 43464 506258
rect 43144 499258 43186 499494
rect 43422 499258 43464 499494
rect 43144 492494 43464 499258
rect 43144 492258 43186 492494
rect 43422 492258 43464 492494
rect 43144 485494 43464 492258
rect 43144 485258 43186 485494
rect 43422 485258 43464 485494
rect 43144 478494 43464 485258
rect 43144 478258 43186 478494
rect 43422 478258 43464 478494
rect 43144 471494 43464 478258
rect 43144 471258 43186 471494
rect 43422 471258 43464 471494
rect 43144 464494 43464 471258
rect 43144 464258 43186 464494
rect 43422 464258 43464 464494
rect 43144 457494 43464 464258
rect 43144 457258 43186 457494
rect 43422 457258 43464 457494
rect 43144 450494 43464 457258
rect 43144 450258 43186 450494
rect 43422 450258 43464 450494
rect 43144 443494 43464 450258
rect 43144 443258 43186 443494
rect 43422 443258 43464 443494
rect 43144 436494 43464 443258
rect 43144 436258 43186 436494
rect 43422 436258 43464 436494
rect 43144 429494 43464 436258
rect 43144 429258 43186 429494
rect 43422 429258 43464 429494
rect 43144 422494 43464 429258
rect 43144 422258 43186 422494
rect 43422 422258 43464 422494
rect 43144 415494 43464 422258
rect 43144 415258 43186 415494
rect 43422 415258 43464 415494
rect 43144 408494 43464 415258
rect 43144 408258 43186 408494
rect 43422 408258 43464 408494
rect 43144 401494 43464 408258
rect 43144 401258 43186 401494
rect 43422 401258 43464 401494
rect 43144 394494 43464 401258
rect 43144 394258 43186 394494
rect 43422 394258 43464 394494
rect 43144 387494 43464 394258
rect 43144 387258 43186 387494
rect 43422 387258 43464 387494
rect 43144 380494 43464 387258
rect 43144 380258 43186 380494
rect 43422 380258 43464 380494
rect 43144 373494 43464 380258
rect 43144 373258 43186 373494
rect 43422 373258 43464 373494
rect 43144 366494 43464 373258
rect 43144 366258 43186 366494
rect 43422 366258 43464 366494
rect 43144 359494 43464 366258
rect 43144 359258 43186 359494
rect 43422 359258 43464 359494
rect 43144 352494 43464 359258
rect 43144 352258 43186 352494
rect 43422 352258 43464 352494
rect 43144 345494 43464 352258
rect 43144 345258 43186 345494
rect 43422 345258 43464 345494
rect 43144 338494 43464 345258
rect 43144 338258 43186 338494
rect 43422 338258 43464 338494
rect 43144 331494 43464 338258
rect 43144 331258 43186 331494
rect 43422 331258 43464 331494
rect 43144 324494 43464 331258
rect 43144 324258 43186 324494
rect 43422 324258 43464 324494
rect 43144 317494 43464 324258
rect 43144 317258 43186 317494
rect 43422 317258 43464 317494
rect 43144 310494 43464 317258
rect 43144 310258 43186 310494
rect 43422 310258 43464 310494
rect 43144 303494 43464 310258
rect 43144 303258 43186 303494
rect 43422 303258 43464 303494
rect 43144 296494 43464 303258
rect 43144 296258 43186 296494
rect 43422 296258 43464 296494
rect 43144 289494 43464 296258
rect 43144 289258 43186 289494
rect 43422 289258 43464 289494
rect 43144 282494 43464 289258
rect 43144 282258 43186 282494
rect 43422 282258 43464 282494
rect 43144 275494 43464 282258
rect 43144 275258 43186 275494
rect 43422 275258 43464 275494
rect 43144 268494 43464 275258
rect 43144 268258 43186 268494
rect 43422 268258 43464 268494
rect 43144 261494 43464 268258
rect 43144 261258 43186 261494
rect 43422 261258 43464 261494
rect 43144 254494 43464 261258
rect 43144 254258 43186 254494
rect 43422 254258 43464 254494
rect 43144 247494 43464 254258
rect 43144 247258 43186 247494
rect 43422 247258 43464 247494
rect 43144 240494 43464 247258
rect 43144 240258 43186 240494
rect 43422 240258 43464 240494
rect 43144 233494 43464 240258
rect 43144 233258 43186 233494
rect 43422 233258 43464 233494
rect 43144 226494 43464 233258
rect 43144 226258 43186 226494
rect 43422 226258 43464 226494
rect 43144 219494 43464 226258
rect 43144 219258 43186 219494
rect 43422 219258 43464 219494
rect 43144 212494 43464 219258
rect 43144 212258 43186 212494
rect 43422 212258 43464 212494
rect 43144 205494 43464 212258
rect 43144 205258 43186 205494
rect 43422 205258 43464 205494
rect 43144 198494 43464 205258
rect 43144 198258 43186 198494
rect 43422 198258 43464 198494
rect 43144 191494 43464 198258
rect 43144 191258 43186 191494
rect 43422 191258 43464 191494
rect 43144 184494 43464 191258
rect 43144 184258 43186 184494
rect 43422 184258 43464 184494
rect 43144 177494 43464 184258
rect 43144 177258 43186 177494
rect 43422 177258 43464 177494
rect 43144 170494 43464 177258
rect 43144 170258 43186 170494
rect 43422 170258 43464 170494
rect 43144 163494 43464 170258
rect 43144 163258 43186 163494
rect 43422 163258 43464 163494
rect 43144 156494 43464 163258
rect 43144 156258 43186 156494
rect 43422 156258 43464 156494
rect 43144 149494 43464 156258
rect 43144 149258 43186 149494
rect 43422 149258 43464 149494
rect 43144 142494 43464 149258
rect 43144 142258 43186 142494
rect 43422 142258 43464 142494
rect 43144 135494 43464 142258
rect 43144 135258 43186 135494
rect 43422 135258 43464 135494
rect 43144 128494 43464 135258
rect 43144 128258 43186 128494
rect 43422 128258 43464 128494
rect 43144 121494 43464 128258
rect 43144 121258 43186 121494
rect 43422 121258 43464 121494
rect 43144 114494 43464 121258
rect 43144 114258 43186 114494
rect 43422 114258 43464 114494
rect 43144 107494 43464 114258
rect 43144 107258 43186 107494
rect 43422 107258 43464 107494
rect 43144 100494 43464 107258
rect 43144 100258 43186 100494
rect 43422 100258 43464 100494
rect 43144 93494 43464 100258
rect 43144 93258 43186 93494
rect 43422 93258 43464 93494
rect 43144 86494 43464 93258
rect 43144 86258 43186 86494
rect 43422 86258 43464 86494
rect 43144 79494 43464 86258
rect 43144 79258 43186 79494
rect 43422 79258 43464 79494
rect 43144 72494 43464 79258
rect 43144 72258 43186 72494
rect 43422 72258 43464 72494
rect 43144 65494 43464 72258
rect 43144 65258 43186 65494
rect 43422 65258 43464 65494
rect 43144 58494 43464 65258
rect 43144 58258 43186 58494
rect 43422 58258 43464 58494
rect 43144 51494 43464 58258
rect 43144 51258 43186 51494
rect 43422 51258 43464 51494
rect 43144 44494 43464 51258
rect 43144 44258 43186 44494
rect 43422 44258 43464 44494
rect 43144 37494 43464 44258
rect 43144 37258 43186 37494
rect 43422 37258 43464 37494
rect 43144 30494 43464 37258
rect 43144 30258 43186 30494
rect 43422 30258 43464 30494
rect 43144 23494 43464 30258
rect 43144 23258 43186 23494
rect 43422 23258 43464 23494
rect 43144 16494 43464 23258
rect 43144 16258 43186 16494
rect 43422 16258 43464 16494
rect 43144 9494 43464 16258
rect 43144 9258 43186 9494
rect 43422 9258 43464 9494
rect 43144 2494 43464 9258
rect 43144 2258 43186 2494
rect 43422 2258 43464 2494
rect 43144 -746 43464 2258
rect 43144 -982 43186 -746
rect 43422 -982 43464 -746
rect 43144 -1066 43464 -982
rect 43144 -1302 43186 -1066
rect 43422 -1302 43464 -1066
rect 43144 -2294 43464 -1302
rect 44876 706198 45196 706230
rect 44876 705962 44918 706198
rect 45154 705962 45196 706198
rect 44876 705878 45196 705962
rect 44876 705642 44918 705878
rect 45154 705642 45196 705878
rect 44876 696561 45196 705642
rect 44876 696325 44918 696561
rect 45154 696325 45196 696561
rect 44876 689561 45196 696325
rect 44876 689325 44918 689561
rect 45154 689325 45196 689561
rect 44876 682561 45196 689325
rect 44876 682325 44918 682561
rect 45154 682325 45196 682561
rect 44876 675561 45196 682325
rect 44876 675325 44918 675561
rect 45154 675325 45196 675561
rect 44876 668561 45196 675325
rect 44876 668325 44918 668561
rect 45154 668325 45196 668561
rect 44876 661561 45196 668325
rect 44876 661325 44918 661561
rect 45154 661325 45196 661561
rect 44876 654561 45196 661325
rect 44876 654325 44918 654561
rect 45154 654325 45196 654561
rect 44876 647561 45196 654325
rect 44876 647325 44918 647561
rect 45154 647325 45196 647561
rect 44876 640561 45196 647325
rect 44876 640325 44918 640561
rect 45154 640325 45196 640561
rect 44876 633561 45196 640325
rect 44876 633325 44918 633561
rect 45154 633325 45196 633561
rect 44876 626561 45196 633325
rect 44876 626325 44918 626561
rect 45154 626325 45196 626561
rect 44876 619561 45196 626325
rect 44876 619325 44918 619561
rect 45154 619325 45196 619561
rect 44876 612561 45196 619325
rect 44876 612325 44918 612561
rect 45154 612325 45196 612561
rect 44876 605561 45196 612325
rect 44876 605325 44918 605561
rect 45154 605325 45196 605561
rect 44876 598561 45196 605325
rect 44876 598325 44918 598561
rect 45154 598325 45196 598561
rect 44876 591561 45196 598325
rect 44876 591325 44918 591561
rect 45154 591325 45196 591561
rect 44876 584561 45196 591325
rect 44876 584325 44918 584561
rect 45154 584325 45196 584561
rect 44876 577561 45196 584325
rect 44876 577325 44918 577561
rect 45154 577325 45196 577561
rect 44876 570561 45196 577325
rect 44876 570325 44918 570561
rect 45154 570325 45196 570561
rect 44876 563561 45196 570325
rect 44876 563325 44918 563561
rect 45154 563325 45196 563561
rect 44876 556561 45196 563325
rect 44876 556325 44918 556561
rect 45154 556325 45196 556561
rect 44876 549561 45196 556325
rect 44876 549325 44918 549561
rect 45154 549325 45196 549561
rect 44876 542561 45196 549325
rect 44876 542325 44918 542561
rect 45154 542325 45196 542561
rect 44876 535561 45196 542325
rect 44876 535325 44918 535561
rect 45154 535325 45196 535561
rect 44876 528561 45196 535325
rect 44876 528325 44918 528561
rect 45154 528325 45196 528561
rect 44876 521561 45196 528325
rect 44876 521325 44918 521561
rect 45154 521325 45196 521561
rect 44876 514561 45196 521325
rect 44876 514325 44918 514561
rect 45154 514325 45196 514561
rect 44876 507561 45196 514325
rect 44876 507325 44918 507561
rect 45154 507325 45196 507561
rect 44876 500561 45196 507325
rect 44876 500325 44918 500561
rect 45154 500325 45196 500561
rect 44876 493561 45196 500325
rect 44876 493325 44918 493561
rect 45154 493325 45196 493561
rect 44876 486561 45196 493325
rect 44876 486325 44918 486561
rect 45154 486325 45196 486561
rect 44876 479561 45196 486325
rect 44876 479325 44918 479561
rect 45154 479325 45196 479561
rect 44876 472561 45196 479325
rect 44876 472325 44918 472561
rect 45154 472325 45196 472561
rect 44876 465561 45196 472325
rect 44876 465325 44918 465561
rect 45154 465325 45196 465561
rect 44876 458561 45196 465325
rect 44876 458325 44918 458561
rect 45154 458325 45196 458561
rect 44876 451561 45196 458325
rect 44876 451325 44918 451561
rect 45154 451325 45196 451561
rect 44876 444561 45196 451325
rect 44876 444325 44918 444561
rect 45154 444325 45196 444561
rect 44876 437561 45196 444325
rect 44876 437325 44918 437561
rect 45154 437325 45196 437561
rect 44876 430561 45196 437325
rect 44876 430325 44918 430561
rect 45154 430325 45196 430561
rect 44876 423561 45196 430325
rect 44876 423325 44918 423561
rect 45154 423325 45196 423561
rect 44876 416561 45196 423325
rect 44876 416325 44918 416561
rect 45154 416325 45196 416561
rect 44876 409561 45196 416325
rect 44876 409325 44918 409561
rect 45154 409325 45196 409561
rect 44876 402561 45196 409325
rect 44876 402325 44918 402561
rect 45154 402325 45196 402561
rect 44876 395561 45196 402325
rect 44876 395325 44918 395561
rect 45154 395325 45196 395561
rect 44876 388561 45196 395325
rect 44876 388325 44918 388561
rect 45154 388325 45196 388561
rect 44876 381561 45196 388325
rect 44876 381325 44918 381561
rect 45154 381325 45196 381561
rect 44876 374561 45196 381325
rect 44876 374325 44918 374561
rect 45154 374325 45196 374561
rect 44876 367561 45196 374325
rect 44876 367325 44918 367561
rect 45154 367325 45196 367561
rect 44876 360561 45196 367325
rect 44876 360325 44918 360561
rect 45154 360325 45196 360561
rect 44876 353561 45196 360325
rect 44876 353325 44918 353561
rect 45154 353325 45196 353561
rect 44876 346561 45196 353325
rect 44876 346325 44918 346561
rect 45154 346325 45196 346561
rect 44876 339561 45196 346325
rect 44876 339325 44918 339561
rect 45154 339325 45196 339561
rect 44876 332561 45196 339325
rect 44876 332325 44918 332561
rect 45154 332325 45196 332561
rect 44876 325561 45196 332325
rect 44876 325325 44918 325561
rect 45154 325325 45196 325561
rect 44876 318561 45196 325325
rect 44876 318325 44918 318561
rect 45154 318325 45196 318561
rect 44876 311561 45196 318325
rect 44876 311325 44918 311561
rect 45154 311325 45196 311561
rect 44876 304561 45196 311325
rect 44876 304325 44918 304561
rect 45154 304325 45196 304561
rect 44876 297561 45196 304325
rect 44876 297325 44918 297561
rect 45154 297325 45196 297561
rect 44876 290561 45196 297325
rect 44876 290325 44918 290561
rect 45154 290325 45196 290561
rect 44876 283561 45196 290325
rect 44876 283325 44918 283561
rect 45154 283325 45196 283561
rect 44876 276561 45196 283325
rect 44876 276325 44918 276561
rect 45154 276325 45196 276561
rect 44876 269561 45196 276325
rect 44876 269325 44918 269561
rect 45154 269325 45196 269561
rect 44876 262561 45196 269325
rect 44876 262325 44918 262561
rect 45154 262325 45196 262561
rect 44876 255561 45196 262325
rect 44876 255325 44918 255561
rect 45154 255325 45196 255561
rect 44876 248561 45196 255325
rect 44876 248325 44918 248561
rect 45154 248325 45196 248561
rect 44876 241561 45196 248325
rect 44876 241325 44918 241561
rect 45154 241325 45196 241561
rect 44876 234561 45196 241325
rect 44876 234325 44918 234561
rect 45154 234325 45196 234561
rect 44876 227561 45196 234325
rect 44876 227325 44918 227561
rect 45154 227325 45196 227561
rect 44876 220561 45196 227325
rect 44876 220325 44918 220561
rect 45154 220325 45196 220561
rect 44876 213561 45196 220325
rect 44876 213325 44918 213561
rect 45154 213325 45196 213561
rect 44876 206561 45196 213325
rect 44876 206325 44918 206561
rect 45154 206325 45196 206561
rect 44876 199561 45196 206325
rect 44876 199325 44918 199561
rect 45154 199325 45196 199561
rect 44876 192561 45196 199325
rect 44876 192325 44918 192561
rect 45154 192325 45196 192561
rect 44876 185561 45196 192325
rect 44876 185325 44918 185561
rect 45154 185325 45196 185561
rect 44876 178561 45196 185325
rect 44876 178325 44918 178561
rect 45154 178325 45196 178561
rect 44876 171561 45196 178325
rect 44876 171325 44918 171561
rect 45154 171325 45196 171561
rect 44876 164561 45196 171325
rect 44876 164325 44918 164561
rect 45154 164325 45196 164561
rect 44876 157561 45196 164325
rect 44876 157325 44918 157561
rect 45154 157325 45196 157561
rect 44876 150561 45196 157325
rect 44876 150325 44918 150561
rect 45154 150325 45196 150561
rect 44876 143561 45196 150325
rect 44876 143325 44918 143561
rect 45154 143325 45196 143561
rect 44876 136561 45196 143325
rect 44876 136325 44918 136561
rect 45154 136325 45196 136561
rect 44876 129561 45196 136325
rect 44876 129325 44918 129561
rect 45154 129325 45196 129561
rect 44876 122561 45196 129325
rect 44876 122325 44918 122561
rect 45154 122325 45196 122561
rect 44876 115561 45196 122325
rect 44876 115325 44918 115561
rect 45154 115325 45196 115561
rect 44876 108561 45196 115325
rect 44876 108325 44918 108561
rect 45154 108325 45196 108561
rect 44876 101561 45196 108325
rect 44876 101325 44918 101561
rect 45154 101325 45196 101561
rect 44876 94561 45196 101325
rect 44876 94325 44918 94561
rect 45154 94325 45196 94561
rect 44876 87561 45196 94325
rect 44876 87325 44918 87561
rect 45154 87325 45196 87561
rect 44876 80561 45196 87325
rect 44876 80325 44918 80561
rect 45154 80325 45196 80561
rect 44876 73561 45196 80325
rect 44876 73325 44918 73561
rect 45154 73325 45196 73561
rect 44876 66561 45196 73325
rect 44876 66325 44918 66561
rect 45154 66325 45196 66561
rect 44876 59561 45196 66325
rect 44876 59325 44918 59561
rect 45154 59325 45196 59561
rect 44876 52561 45196 59325
rect 44876 52325 44918 52561
rect 45154 52325 45196 52561
rect 44876 45561 45196 52325
rect 44876 45325 44918 45561
rect 45154 45325 45196 45561
rect 44876 38561 45196 45325
rect 44876 38325 44918 38561
rect 45154 38325 45196 38561
rect 44876 31561 45196 38325
rect 44876 31325 44918 31561
rect 45154 31325 45196 31561
rect 44876 24561 45196 31325
rect 44876 24325 44918 24561
rect 45154 24325 45196 24561
rect 44876 17561 45196 24325
rect 44876 17325 44918 17561
rect 45154 17325 45196 17561
rect 44876 10561 45196 17325
rect 44876 10325 44918 10561
rect 45154 10325 45196 10561
rect 44876 3561 45196 10325
rect 44876 3325 44918 3561
rect 45154 3325 45196 3561
rect 44876 -1706 45196 3325
rect 44876 -1942 44918 -1706
rect 45154 -1942 45196 -1706
rect 44876 -2026 45196 -1942
rect 44876 -2262 44918 -2026
rect 45154 -2262 45196 -2026
rect 44876 -2294 45196 -2262
rect 50144 705238 50464 706230
rect 50144 705002 50186 705238
rect 50422 705002 50464 705238
rect 50144 704918 50464 705002
rect 50144 704682 50186 704918
rect 50422 704682 50464 704918
rect 50144 695494 50464 704682
rect 50144 695258 50186 695494
rect 50422 695258 50464 695494
rect 50144 688494 50464 695258
rect 50144 688258 50186 688494
rect 50422 688258 50464 688494
rect 50144 681494 50464 688258
rect 50144 681258 50186 681494
rect 50422 681258 50464 681494
rect 50144 674494 50464 681258
rect 50144 674258 50186 674494
rect 50422 674258 50464 674494
rect 50144 667494 50464 674258
rect 50144 667258 50186 667494
rect 50422 667258 50464 667494
rect 50144 660494 50464 667258
rect 50144 660258 50186 660494
rect 50422 660258 50464 660494
rect 50144 653494 50464 660258
rect 50144 653258 50186 653494
rect 50422 653258 50464 653494
rect 50144 646494 50464 653258
rect 50144 646258 50186 646494
rect 50422 646258 50464 646494
rect 50144 639494 50464 646258
rect 50144 639258 50186 639494
rect 50422 639258 50464 639494
rect 50144 632494 50464 639258
rect 50144 632258 50186 632494
rect 50422 632258 50464 632494
rect 50144 625494 50464 632258
rect 50144 625258 50186 625494
rect 50422 625258 50464 625494
rect 50144 618494 50464 625258
rect 50144 618258 50186 618494
rect 50422 618258 50464 618494
rect 50144 611494 50464 618258
rect 50144 611258 50186 611494
rect 50422 611258 50464 611494
rect 50144 604494 50464 611258
rect 50144 604258 50186 604494
rect 50422 604258 50464 604494
rect 50144 597494 50464 604258
rect 50144 597258 50186 597494
rect 50422 597258 50464 597494
rect 50144 590494 50464 597258
rect 50144 590258 50186 590494
rect 50422 590258 50464 590494
rect 50144 583494 50464 590258
rect 50144 583258 50186 583494
rect 50422 583258 50464 583494
rect 50144 576494 50464 583258
rect 50144 576258 50186 576494
rect 50422 576258 50464 576494
rect 50144 569494 50464 576258
rect 50144 569258 50186 569494
rect 50422 569258 50464 569494
rect 50144 562494 50464 569258
rect 50144 562258 50186 562494
rect 50422 562258 50464 562494
rect 50144 555494 50464 562258
rect 50144 555258 50186 555494
rect 50422 555258 50464 555494
rect 50144 548494 50464 555258
rect 50144 548258 50186 548494
rect 50422 548258 50464 548494
rect 50144 541494 50464 548258
rect 50144 541258 50186 541494
rect 50422 541258 50464 541494
rect 50144 534494 50464 541258
rect 50144 534258 50186 534494
rect 50422 534258 50464 534494
rect 50144 527494 50464 534258
rect 50144 527258 50186 527494
rect 50422 527258 50464 527494
rect 50144 520494 50464 527258
rect 50144 520258 50186 520494
rect 50422 520258 50464 520494
rect 50144 513494 50464 520258
rect 50144 513258 50186 513494
rect 50422 513258 50464 513494
rect 50144 506494 50464 513258
rect 50144 506258 50186 506494
rect 50422 506258 50464 506494
rect 50144 499494 50464 506258
rect 50144 499258 50186 499494
rect 50422 499258 50464 499494
rect 50144 492494 50464 499258
rect 50144 492258 50186 492494
rect 50422 492258 50464 492494
rect 50144 485494 50464 492258
rect 50144 485258 50186 485494
rect 50422 485258 50464 485494
rect 50144 478494 50464 485258
rect 50144 478258 50186 478494
rect 50422 478258 50464 478494
rect 50144 471494 50464 478258
rect 50144 471258 50186 471494
rect 50422 471258 50464 471494
rect 50144 464494 50464 471258
rect 50144 464258 50186 464494
rect 50422 464258 50464 464494
rect 50144 457494 50464 464258
rect 50144 457258 50186 457494
rect 50422 457258 50464 457494
rect 50144 450494 50464 457258
rect 50144 450258 50186 450494
rect 50422 450258 50464 450494
rect 50144 443494 50464 450258
rect 50144 443258 50186 443494
rect 50422 443258 50464 443494
rect 50144 436494 50464 443258
rect 50144 436258 50186 436494
rect 50422 436258 50464 436494
rect 50144 429494 50464 436258
rect 50144 429258 50186 429494
rect 50422 429258 50464 429494
rect 50144 422494 50464 429258
rect 50144 422258 50186 422494
rect 50422 422258 50464 422494
rect 50144 415494 50464 422258
rect 50144 415258 50186 415494
rect 50422 415258 50464 415494
rect 50144 408494 50464 415258
rect 50144 408258 50186 408494
rect 50422 408258 50464 408494
rect 50144 401494 50464 408258
rect 50144 401258 50186 401494
rect 50422 401258 50464 401494
rect 50144 394494 50464 401258
rect 50144 394258 50186 394494
rect 50422 394258 50464 394494
rect 50144 387494 50464 394258
rect 50144 387258 50186 387494
rect 50422 387258 50464 387494
rect 50144 380494 50464 387258
rect 50144 380258 50186 380494
rect 50422 380258 50464 380494
rect 50144 373494 50464 380258
rect 50144 373258 50186 373494
rect 50422 373258 50464 373494
rect 50144 366494 50464 373258
rect 50144 366258 50186 366494
rect 50422 366258 50464 366494
rect 50144 359494 50464 366258
rect 50144 359258 50186 359494
rect 50422 359258 50464 359494
rect 50144 352494 50464 359258
rect 50144 352258 50186 352494
rect 50422 352258 50464 352494
rect 50144 345494 50464 352258
rect 50144 345258 50186 345494
rect 50422 345258 50464 345494
rect 50144 338494 50464 345258
rect 50144 338258 50186 338494
rect 50422 338258 50464 338494
rect 50144 331494 50464 338258
rect 50144 331258 50186 331494
rect 50422 331258 50464 331494
rect 50144 324494 50464 331258
rect 50144 324258 50186 324494
rect 50422 324258 50464 324494
rect 50144 317494 50464 324258
rect 50144 317258 50186 317494
rect 50422 317258 50464 317494
rect 50144 310494 50464 317258
rect 50144 310258 50186 310494
rect 50422 310258 50464 310494
rect 50144 303494 50464 310258
rect 50144 303258 50186 303494
rect 50422 303258 50464 303494
rect 50144 296494 50464 303258
rect 50144 296258 50186 296494
rect 50422 296258 50464 296494
rect 50144 289494 50464 296258
rect 50144 289258 50186 289494
rect 50422 289258 50464 289494
rect 50144 282494 50464 289258
rect 50144 282258 50186 282494
rect 50422 282258 50464 282494
rect 50144 275494 50464 282258
rect 50144 275258 50186 275494
rect 50422 275258 50464 275494
rect 50144 268494 50464 275258
rect 50144 268258 50186 268494
rect 50422 268258 50464 268494
rect 50144 261494 50464 268258
rect 50144 261258 50186 261494
rect 50422 261258 50464 261494
rect 50144 254494 50464 261258
rect 50144 254258 50186 254494
rect 50422 254258 50464 254494
rect 50144 247494 50464 254258
rect 50144 247258 50186 247494
rect 50422 247258 50464 247494
rect 50144 240494 50464 247258
rect 50144 240258 50186 240494
rect 50422 240258 50464 240494
rect 50144 233494 50464 240258
rect 50144 233258 50186 233494
rect 50422 233258 50464 233494
rect 50144 226494 50464 233258
rect 50144 226258 50186 226494
rect 50422 226258 50464 226494
rect 50144 219494 50464 226258
rect 50144 219258 50186 219494
rect 50422 219258 50464 219494
rect 50144 212494 50464 219258
rect 50144 212258 50186 212494
rect 50422 212258 50464 212494
rect 50144 205494 50464 212258
rect 50144 205258 50186 205494
rect 50422 205258 50464 205494
rect 50144 198494 50464 205258
rect 50144 198258 50186 198494
rect 50422 198258 50464 198494
rect 50144 191494 50464 198258
rect 50144 191258 50186 191494
rect 50422 191258 50464 191494
rect 50144 184494 50464 191258
rect 50144 184258 50186 184494
rect 50422 184258 50464 184494
rect 50144 177494 50464 184258
rect 50144 177258 50186 177494
rect 50422 177258 50464 177494
rect 50144 170494 50464 177258
rect 50144 170258 50186 170494
rect 50422 170258 50464 170494
rect 50144 163494 50464 170258
rect 50144 163258 50186 163494
rect 50422 163258 50464 163494
rect 50144 156494 50464 163258
rect 50144 156258 50186 156494
rect 50422 156258 50464 156494
rect 50144 149494 50464 156258
rect 50144 149258 50186 149494
rect 50422 149258 50464 149494
rect 50144 142494 50464 149258
rect 50144 142258 50186 142494
rect 50422 142258 50464 142494
rect 50144 135494 50464 142258
rect 50144 135258 50186 135494
rect 50422 135258 50464 135494
rect 50144 128494 50464 135258
rect 50144 128258 50186 128494
rect 50422 128258 50464 128494
rect 50144 121494 50464 128258
rect 50144 121258 50186 121494
rect 50422 121258 50464 121494
rect 50144 114494 50464 121258
rect 50144 114258 50186 114494
rect 50422 114258 50464 114494
rect 50144 107494 50464 114258
rect 50144 107258 50186 107494
rect 50422 107258 50464 107494
rect 50144 100494 50464 107258
rect 50144 100258 50186 100494
rect 50422 100258 50464 100494
rect 50144 93494 50464 100258
rect 50144 93258 50186 93494
rect 50422 93258 50464 93494
rect 50144 86494 50464 93258
rect 50144 86258 50186 86494
rect 50422 86258 50464 86494
rect 50144 79494 50464 86258
rect 50144 79258 50186 79494
rect 50422 79258 50464 79494
rect 50144 72494 50464 79258
rect 50144 72258 50186 72494
rect 50422 72258 50464 72494
rect 50144 65494 50464 72258
rect 50144 65258 50186 65494
rect 50422 65258 50464 65494
rect 50144 58494 50464 65258
rect 50144 58258 50186 58494
rect 50422 58258 50464 58494
rect 50144 51494 50464 58258
rect 50144 51258 50186 51494
rect 50422 51258 50464 51494
rect 50144 44494 50464 51258
rect 50144 44258 50186 44494
rect 50422 44258 50464 44494
rect 50144 37494 50464 44258
rect 50144 37258 50186 37494
rect 50422 37258 50464 37494
rect 50144 30494 50464 37258
rect 50144 30258 50186 30494
rect 50422 30258 50464 30494
rect 50144 23494 50464 30258
rect 50144 23258 50186 23494
rect 50422 23258 50464 23494
rect 50144 16494 50464 23258
rect 50144 16258 50186 16494
rect 50422 16258 50464 16494
rect 50144 9494 50464 16258
rect 50144 9258 50186 9494
rect 50422 9258 50464 9494
rect 50144 2494 50464 9258
rect 50144 2258 50186 2494
rect 50422 2258 50464 2494
rect 50144 -746 50464 2258
rect 50144 -982 50186 -746
rect 50422 -982 50464 -746
rect 50144 -1066 50464 -982
rect 50144 -1302 50186 -1066
rect 50422 -1302 50464 -1066
rect 50144 -2294 50464 -1302
rect 51876 706198 52196 706230
rect 51876 705962 51918 706198
rect 52154 705962 52196 706198
rect 51876 705878 52196 705962
rect 51876 705642 51918 705878
rect 52154 705642 52196 705878
rect 51876 696561 52196 705642
rect 51876 696325 51918 696561
rect 52154 696325 52196 696561
rect 51876 689561 52196 696325
rect 51876 689325 51918 689561
rect 52154 689325 52196 689561
rect 51876 682561 52196 689325
rect 51876 682325 51918 682561
rect 52154 682325 52196 682561
rect 51876 675561 52196 682325
rect 51876 675325 51918 675561
rect 52154 675325 52196 675561
rect 51876 668561 52196 675325
rect 51876 668325 51918 668561
rect 52154 668325 52196 668561
rect 51876 661561 52196 668325
rect 51876 661325 51918 661561
rect 52154 661325 52196 661561
rect 51876 654561 52196 661325
rect 51876 654325 51918 654561
rect 52154 654325 52196 654561
rect 51876 647561 52196 654325
rect 51876 647325 51918 647561
rect 52154 647325 52196 647561
rect 51876 640561 52196 647325
rect 51876 640325 51918 640561
rect 52154 640325 52196 640561
rect 51876 633561 52196 640325
rect 51876 633325 51918 633561
rect 52154 633325 52196 633561
rect 51876 626561 52196 633325
rect 51876 626325 51918 626561
rect 52154 626325 52196 626561
rect 51876 619561 52196 626325
rect 51876 619325 51918 619561
rect 52154 619325 52196 619561
rect 51876 612561 52196 619325
rect 51876 612325 51918 612561
rect 52154 612325 52196 612561
rect 51876 605561 52196 612325
rect 51876 605325 51918 605561
rect 52154 605325 52196 605561
rect 51876 598561 52196 605325
rect 51876 598325 51918 598561
rect 52154 598325 52196 598561
rect 51876 591561 52196 598325
rect 51876 591325 51918 591561
rect 52154 591325 52196 591561
rect 51876 584561 52196 591325
rect 51876 584325 51918 584561
rect 52154 584325 52196 584561
rect 51876 577561 52196 584325
rect 51876 577325 51918 577561
rect 52154 577325 52196 577561
rect 51876 570561 52196 577325
rect 51876 570325 51918 570561
rect 52154 570325 52196 570561
rect 51876 563561 52196 570325
rect 51876 563325 51918 563561
rect 52154 563325 52196 563561
rect 51876 556561 52196 563325
rect 51876 556325 51918 556561
rect 52154 556325 52196 556561
rect 51876 549561 52196 556325
rect 51876 549325 51918 549561
rect 52154 549325 52196 549561
rect 51876 542561 52196 549325
rect 51876 542325 51918 542561
rect 52154 542325 52196 542561
rect 51876 535561 52196 542325
rect 51876 535325 51918 535561
rect 52154 535325 52196 535561
rect 51876 528561 52196 535325
rect 51876 528325 51918 528561
rect 52154 528325 52196 528561
rect 51876 521561 52196 528325
rect 51876 521325 51918 521561
rect 52154 521325 52196 521561
rect 51876 514561 52196 521325
rect 51876 514325 51918 514561
rect 52154 514325 52196 514561
rect 51876 507561 52196 514325
rect 51876 507325 51918 507561
rect 52154 507325 52196 507561
rect 51876 500561 52196 507325
rect 51876 500325 51918 500561
rect 52154 500325 52196 500561
rect 51876 493561 52196 500325
rect 51876 493325 51918 493561
rect 52154 493325 52196 493561
rect 51876 486561 52196 493325
rect 51876 486325 51918 486561
rect 52154 486325 52196 486561
rect 51876 479561 52196 486325
rect 51876 479325 51918 479561
rect 52154 479325 52196 479561
rect 51876 472561 52196 479325
rect 51876 472325 51918 472561
rect 52154 472325 52196 472561
rect 51876 465561 52196 472325
rect 51876 465325 51918 465561
rect 52154 465325 52196 465561
rect 51876 458561 52196 465325
rect 51876 458325 51918 458561
rect 52154 458325 52196 458561
rect 51876 451561 52196 458325
rect 51876 451325 51918 451561
rect 52154 451325 52196 451561
rect 51876 444561 52196 451325
rect 51876 444325 51918 444561
rect 52154 444325 52196 444561
rect 51876 437561 52196 444325
rect 51876 437325 51918 437561
rect 52154 437325 52196 437561
rect 51876 430561 52196 437325
rect 51876 430325 51918 430561
rect 52154 430325 52196 430561
rect 51876 423561 52196 430325
rect 51876 423325 51918 423561
rect 52154 423325 52196 423561
rect 51876 416561 52196 423325
rect 51876 416325 51918 416561
rect 52154 416325 52196 416561
rect 51876 409561 52196 416325
rect 51876 409325 51918 409561
rect 52154 409325 52196 409561
rect 51876 402561 52196 409325
rect 51876 402325 51918 402561
rect 52154 402325 52196 402561
rect 51876 395561 52196 402325
rect 51876 395325 51918 395561
rect 52154 395325 52196 395561
rect 51876 388561 52196 395325
rect 51876 388325 51918 388561
rect 52154 388325 52196 388561
rect 51876 381561 52196 388325
rect 51876 381325 51918 381561
rect 52154 381325 52196 381561
rect 51876 374561 52196 381325
rect 51876 374325 51918 374561
rect 52154 374325 52196 374561
rect 51876 367561 52196 374325
rect 51876 367325 51918 367561
rect 52154 367325 52196 367561
rect 51876 360561 52196 367325
rect 51876 360325 51918 360561
rect 52154 360325 52196 360561
rect 51876 353561 52196 360325
rect 51876 353325 51918 353561
rect 52154 353325 52196 353561
rect 51876 346561 52196 353325
rect 51876 346325 51918 346561
rect 52154 346325 52196 346561
rect 51876 339561 52196 346325
rect 51876 339325 51918 339561
rect 52154 339325 52196 339561
rect 51876 332561 52196 339325
rect 51876 332325 51918 332561
rect 52154 332325 52196 332561
rect 51876 325561 52196 332325
rect 51876 325325 51918 325561
rect 52154 325325 52196 325561
rect 51876 318561 52196 325325
rect 51876 318325 51918 318561
rect 52154 318325 52196 318561
rect 51876 311561 52196 318325
rect 51876 311325 51918 311561
rect 52154 311325 52196 311561
rect 51876 304561 52196 311325
rect 51876 304325 51918 304561
rect 52154 304325 52196 304561
rect 51876 297561 52196 304325
rect 51876 297325 51918 297561
rect 52154 297325 52196 297561
rect 51876 290561 52196 297325
rect 51876 290325 51918 290561
rect 52154 290325 52196 290561
rect 51876 283561 52196 290325
rect 51876 283325 51918 283561
rect 52154 283325 52196 283561
rect 51876 276561 52196 283325
rect 51876 276325 51918 276561
rect 52154 276325 52196 276561
rect 51876 269561 52196 276325
rect 51876 269325 51918 269561
rect 52154 269325 52196 269561
rect 51876 262561 52196 269325
rect 51876 262325 51918 262561
rect 52154 262325 52196 262561
rect 51876 255561 52196 262325
rect 51876 255325 51918 255561
rect 52154 255325 52196 255561
rect 51876 248561 52196 255325
rect 51876 248325 51918 248561
rect 52154 248325 52196 248561
rect 51876 241561 52196 248325
rect 51876 241325 51918 241561
rect 52154 241325 52196 241561
rect 51876 234561 52196 241325
rect 51876 234325 51918 234561
rect 52154 234325 52196 234561
rect 51876 227561 52196 234325
rect 51876 227325 51918 227561
rect 52154 227325 52196 227561
rect 51876 220561 52196 227325
rect 51876 220325 51918 220561
rect 52154 220325 52196 220561
rect 51876 213561 52196 220325
rect 51876 213325 51918 213561
rect 52154 213325 52196 213561
rect 51876 206561 52196 213325
rect 51876 206325 51918 206561
rect 52154 206325 52196 206561
rect 51876 199561 52196 206325
rect 51876 199325 51918 199561
rect 52154 199325 52196 199561
rect 51876 192561 52196 199325
rect 51876 192325 51918 192561
rect 52154 192325 52196 192561
rect 51876 185561 52196 192325
rect 51876 185325 51918 185561
rect 52154 185325 52196 185561
rect 51876 178561 52196 185325
rect 51876 178325 51918 178561
rect 52154 178325 52196 178561
rect 51876 171561 52196 178325
rect 51876 171325 51918 171561
rect 52154 171325 52196 171561
rect 51876 164561 52196 171325
rect 51876 164325 51918 164561
rect 52154 164325 52196 164561
rect 51876 157561 52196 164325
rect 51876 157325 51918 157561
rect 52154 157325 52196 157561
rect 51876 150561 52196 157325
rect 51876 150325 51918 150561
rect 52154 150325 52196 150561
rect 51876 143561 52196 150325
rect 51876 143325 51918 143561
rect 52154 143325 52196 143561
rect 51876 136561 52196 143325
rect 51876 136325 51918 136561
rect 52154 136325 52196 136561
rect 51876 129561 52196 136325
rect 51876 129325 51918 129561
rect 52154 129325 52196 129561
rect 51876 122561 52196 129325
rect 51876 122325 51918 122561
rect 52154 122325 52196 122561
rect 51876 115561 52196 122325
rect 51876 115325 51918 115561
rect 52154 115325 52196 115561
rect 51876 108561 52196 115325
rect 51876 108325 51918 108561
rect 52154 108325 52196 108561
rect 51876 101561 52196 108325
rect 51876 101325 51918 101561
rect 52154 101325 52196 101561
rect 51876 94561 52196 101325
rect 51876 94325 51918 94561
rect 52154 94325 52196 94561
rect 51876 87561 52196 94325
rect 51876 87325 51918 87561
rect 52154 87325 52196 87561
rect 51876 80561 52196 87325
rect 51876 80325 51918 80561
rect 52154 80325 52196 80561
rect 51876 73561 52196 80325
rect 51876 73325 51918 73561
rect 52154 73325 52196 73561
rect 51876 66561 52196 73325
rect 51876 66325 51918 66561
rect 52154 66325 52196 66561
rect 51876 59561 52196 66325
rect 51876 59325 51918 59561
rect 52154 59325 52196 59561
rect 51876 52561 52196 59325
rect 51876 52325 51918 52561
rect 52154 52325 52196 52561
rect 51876 45561 52196 52325
rect 51876 45325 51918 45561
rect 52154 45325 52196 45561
rect 51876 38561 52196 45325
rect 51876 38325 51918 38561
rect 52154 38325 52196 38561
rect 51876 31561 52196 38325
rect 51876 31325 51918 31561
rect 52154 31325 52196 31561
rect 51876 24561 52196 31325
rect 51876 24325 51918 24561
rect 52154 24325 52196 24561
rect 51876 17561 52196 24325
rect 51876 17325 51918 17561
rect 52154 17325 52196 17561
rect 51876 10561 52196 17325
rect 51876 10325 51918 10561
rect 52154 10325 52196 10561
rect 51876 3561 52196 10325
rect 51876 3325 51918 3561
rect 52154 3325 52196 3561
rect 51876 -1706 52196 3325
rect 51876 -1942 51918 -1706
rect 52154 -1942 52196 -1706
rect 51876 -2026 52196 -1942
rect 51876 -2262 51918 -2026
rect 52154 -2262 52196 -2026
rect 51876 -2294 52196 -2262
rect 57144 705238 57464 706230
rect 57144 705002 57186 705238
rect 57422 705002 57464 705238
rect 57144 704918 57464 705002
rect 57144 704682 57186 704918
rect 57422 704682 57464 704918
rect 57144 695494 57464 704682
rect 57144 695258 57186 695494
rect 57422 695258 57464 695494
rect 57144 688494 57464 695258
rect 57144 688258 57186 688494
rect 57422 688258 57464 688494
rect 57144 681494 57464 688258
rect 57144 681258 57186 681494
rect 57422 681258 57464 681494
rect 57144 674494 57464 681258
rect 57144 674258 57186 674494
rect 57422 674258 57464 674494
rect 57144 667494 57464 674258
rect 57144 667258 57186 667494
rect 57422 667258 57464 667494
rect 57144 660494 57464 667258
rect 57144 660258 57186 660494
rect 57422 660258 57464 660494
rect 57144 653494 57464 660258
rect 57144 653258 57186 653494
rect 57422 653258 57464 653494
rect 57144 646494 57464 653258
rect 57144 646258 57186 646494
rect 57422 646258 57464 646494
rect 57144 639494 57464 646258
rect 57144 639258 57186 639494
rect 57422 639258 57464 639494
rect 57144 632494 57464 639258
rect 57144 632258 57186 632494
rect 57422 632258 57464 632494
rect 57144 625494 57464 632258
rect 57144 625258 57186 625494
rect 57422 625258 57464 625494
rect 57144 618494 57464 625258
rect 57144 618258 57186 618494
rect 57422 618258 57464 618494
rect 57144 611494 57464 618258
rect 57144 611258 57186 611494
rect 57422 611258 57464 611494
rect 57144 604494 57464 611258
rect 57144 604258 57186 604494
rect 57422 604258 57464 604494
rect 57144 597494 57464 604258
rect 57144 597258 57186 597494
rect 57422 597258 57464 597494
rect 57144 590494 57464 597258
rect 57144 590258 57186 590494
rect 57422 590258 57464 590494
rect 57144 583494 57464 590258
rect 57144 583258 57186 583494
rect 57422 583258 57464 583494
rect 57144 576494 57464 583258
rect 57144 576258 57186 576494
rect 57422 576258 57464 576494
rect 57144 569494 57464 576258
rect 57144 569258 57186 569494
rect 57422 569258 57464 569494
rect 57144 562494 57464 569258
rect 57144 562258 57186 562494
rect 57422 562258 57464 562494
rect 57144 555494 57464 562258
rect 57144 555258 57186 555494
rect 57422 555258 57464 555494
rect 57144 548494 57464 555258
rect 57144 548258 57186 548494
rect 57422 548258 57464 548494
rect 57144 541494 57464 548258
rect 57144 541258 57186 541494
rect 57422 541258 57464 541494
rect 57144 534494 57464 541258
rect 57144 534258 57186 534494
rect 57422 534258 57464 534494
rect 57144 527494 57464 534258
rect 57144 527258 57186 527494
rect 57422 527258 57464 527494
rect 57144 520494 57464 527258
rect 57144 520258 57186 520494
rect 57422 520258 57464 520494
rect 57144 513494 57464 520258
rect 57144 513258 57186 513494
rect 57422 513258 57464 513494
rect 57144 506494 57464 513258
rect 57144 506258 57186 506494
rect 57422 506258 57464 506494
rect 57144 499494 57464 506258
rect 57144 499258 57186 499494
rect 57422 499258 57464 499494
rect 57144 492494 57464 499258
rect 57144 492258 57186 492494
rect 57422 492258 57464 492494
rect 57144 485494 57464 492258
rect 57144 485258 57186 485494
rect 57422 485258 57464 485494
rect 57144 478494 57464 485258
rect 57144 478258 57186 478494
rect 57422 478258 57464 478494
rect 57144 471494 57464 478258
rect 57144 471258 57186 471494
rect 57422 471258 57464 471494
rect 57144 464494 57464 471258
rect 57144 464258 57186 464494
rect 57422 464258 57464 464494
rect 57144 457494 57464 464258
rect 57144 457258 57186 457494
rect 57422 457258 57464 457494
rect 57144 450494 57464 457258
rect 57144 450258 57186 450494
rect 57422 450258 57464 450494
rect 57144 443494 57464 450258
rect 57144 443258 57186 443494
rect 57422 443258 57464 443494
rect 57144 436494 57464 443258
rect 57144 436258 57186 436494
rect 57422 436258 57464 436494
rect 57144 429494 57464 436258
rect 57144 429258 57186 429494
rect 57422 429258 57464 429494
rect 57144 422494 57464 429258
rect 57144 422258 57186 422494
rect 57422 422258 57464 422494
rect 57144 415494 57464 422258
rect 57144 415258 57186 415494
rect 57422 415258 57464 415494
rect 57144 408494 57464 415258
rect 57144 408258 57186 408494
rect 57422 408258 57464 408494
rect 57144 401494 57464 408258
rect 57144 401258 57186 401494
rect 57422 401258 57464 401494
rect 57144 394494 57464 401258
rect 57144 394258 57186 394494
rect 57422 394258 57464 394494
rect 57144 387494 57464 394258
rect 57144 387258 57186 387494
rect 57422 387258 57464 387494
rect 57144 380494 57464 387258
rect 57144 380258 57186 380494
rect 57422 380258 57464 380494
rect 57144 373494 57464 380258
rect 57144 373258 57186 373494
rect 57422 373258 57464 373494
rect 57144 366494 57464 373258
rect 57144 366258 57186 366494
rect 57422 366258 57464 366494
rect 57144 359494 57464 366258
rect 57144 359258 57186 359494
rect 57422 359258 57464 359494
rect 57144 352494 57464 359258
rect 57144 352258 57186 352494
rect 57422 352258 57464 352494
rect 57144 345494 57464 352258
rect 57144 345258 57186 345494
rect 57422 345258 57464 345494
rect 57144 338494 57464 345258
rect 57144 338258 57186 338494
rect 57422 338258 57464 338494
rect 57144 331494 57464 338258
rect 57144 331258 57186 331494
rect 57422 331258 57464 331494
rect 57144 324494 57464 331258
rect 57144 324258 57186 324494
rect 57422 324258 57464 324494
rect 57144 317494 57464 324258
rect 57144 317258 57186 317494
rect 57422 317258 57464 317494
rect 57144 310494 57464 317258
rect 57144 310258 57186 310494
rect 57422 310258 57464 310494
rect 57144 303494 57464 310258
rect 57144 303258 57186 303494
rect 57422 303258 57464 303494
rect 57144 296494 57464 303258
rect 57144 296258 57186 296494
rect 57422 296258 57464 296494
rect 57144 289494 57464 296258
rect 57144 289258 57186 289494
rect 57422 289258 57464 289494
rect 57144 282494 57464 289258
rect 57144 282258 57186 282494
rect 57422 282258 57464 282494
rect 57144 275494 57464 282258
rect 57144 275258 57186 275494
rect 57422 275258 57464 275494
rect 57144 268494 57464 275258
rect 57144 268258 57186 268494
rect 57422 268258 57464 268494
rect 57144 261494 57464 268258
rect 57144 261258 57186 261494
rect 57422 261258 57464 261494
rect 57144 254494 57464 261258
rect 57144 254258 57186 254494
rect 57422 254258 57464 254494
rect 57144 247494 57464 254258
rect 57144 247258 57186 247494
rect 57422 247258 57464 247494
rect 57144 240494 57464 247258
rect 57144 240258 57186 240494
rect 57422 240258 57464 240494
rect 57144 233494 57464 240258
rect 57144 233258 57186 233494
rect 57422 233258 57464 233494
rect 57144 226494 57464 233258
rect 57144 226258 57186 226494
rect 57422 226258 57464 226494
rect 57144 219494 57464 226258
rect 57144 219258 57186 219494
rect 57422 219258 57464 219494
rect 57144 212494 57464 219258
rect 57144 212258 57186 212494
rect 57422 212258 57464 212494
rect 57144 205494 57464 212258
rect 57144 205258 57186 205494
rect 57422 205258 57464 205494
rect 57144 198494 57464 205258
rect 57144 198258 57186 198494
rect 57422 198258 57464 198494
rect 57144 191494 57464 198258
rect 57144 191258 57186 191494
rect 57422 191258 57464 191494
rect 57144 184494 57464 191258
rect 57144 184258 57186 184494
rect 57422 184258 57464 184494
rect 57144 177494 57464 184258
rect 57144 177258 57186 177494
rect 57422 177258 57464 177494
rect 57144 170494 57464 177258
rect 57144 170258 57186 170494
rect 57422 170258 57464 170494
rect 57144 163494 57464 170258
rect 57144 163258 57186 163494
rect 57422 163258 57464 163494
rect 57144 156494 57464 163258
rect 57144 156258 57186 156494
rect 57422 156258 57464 156494
rect 57144 149494 57464 156258
rect 57144 149258 57186 149494
rect 57422 149258 57464 149494
rect 57144 142494 57464 149258
rect 57144 142258 57186 142494
rect 57422 142258 57464 142494
rect 57144 135494 57464 142258
rect 57144 135258 57186 135494
rect 57422 135258 57464 135494
rect 57144 128494 57464 135258
rect 57144 128258 57186 128494
rect 57422 128258 57464 128494
rect 57144 121494 57464 128258
rect 57144 121258 57186 121494
rect 57422 121258 57464 121494
rect 57144 114494 57464 121258
rect 57144 114258 57186 114494
rect 57422 114258 57464 114494
rect 57144 107494 57464 114258
rect 57144 107258 57186 107494
rect 57422 107258 57464 107494
rect 57144 100494 57464 107258
rect 57144 100258 57186 100494
rect 57422 100258 57464 100494
rect 57144 93494 57464 100258
rect 57144 93258 57186 93494
rect 57422 93258 57464 93494
rect 57144 86494 57464 93258
rect 57144 86258 57186 86494
rect 57422 86258 57464 86494
rect 57144 79494 57464 86258
rect 57144 79258 57186 79494
rect 57422 79258 57464 79494
rect 57144 72494 57464 79258
rect 57144 72258 57186 72494
rect 57422 72258 57464 72494
rect 57144 65494 57464 72258
rect 57144 65258 57186 65494
rect 57422 65258 57464 65494
rect 57144 58494 57464 65258
rect 57144 58258 57186 58494
rect 57422 58258 57464 58494
rect 57144 51494 57464 58258
rect 57144 51258 57186 51494
rect 57422 51258 57464 51494
rect 57144 44494 57464 51258
rect 57144 44258 57186 44494
rect 57422 44258 57464 44494
rect 57144 37494 57464 44258
rect 57144 37258 57186 37494
rect 57422 37258 57464 37494
rect 57144 30494 57464 37258
rect 57144 30258 57186 30494
rect 57422 30258 57464 30494
rect 57144 23494 57464 30258
rect 57144 23258 57186 23494
rect 57422 23258 57464 23494
rect 57144 16494 57464 23258
rect 57144 16258 57186 16494
rect 57422 16258 57464 16494
rect 57144 9494 57464 16258
rect 57144 9258 57186 9494
rect 57422 9258 57464 9494
rect 57144 2494 57464 9258
rect 57144 2258 57186 2494
rect 57422 2258 57464 2494
rect 57144 -746 57464 2258
rect 57144 -982 57186 -746
rect 57422 -982 57464 -746
rect 57144 -1066 57464 -982
rect 57144 -1302 57186 -1066
rect 57422 -1302 57464 -1066
rect 57144 -2294 57464 -1302
rect 58876 706198 59196 706230
rect 58876 705962 58918 706198
rect 59154 705962 59196 706198
rect 58876 705878 59196 705962
rect 58876 705642 58918 705878
rect 59154 705642 59196 705878
rect 58876 696561 59196 705642
rect 58876 696325 58918 696561
rect 59154 696325 59196 696561
rect 58876 689561 59196 696325
rect 58876 689325 58918 689561
rect 59154 689325 59196 689561
rect 58876 682561 59196 689325
rect 58876 682325 58918 682561
rect 59154 682325 59196 682561
rect 58876 675561 59196 682325
rect 58876 675325 58918 675561
rect 59154 675325 59196 675561
rect 58876 668561 59196 675325
rect 58876 668325 58918 668561
rect 59154 668325 59196 668561
rect 58876 661561 59196 668325
rect 58876 661325 58918 661561
rect 59154 661325 59196 661561
rect 58876 654561 59196 661325
rect 58876 654325 58918 654561
rect 59154 654325 59196 654561
rect 58876 647561 59196 654325
rect 58876 647325 58918 647561
rect 59154 647325 59196 647561
rect 58876 640561 59196 647325
rect 58876 640325 58918 640561
rect 59154 640325 59196 640561
rect 58876 633561 59196 640325
rect 58876 633325 58918 633561
rect 59154 633325 59196 633561
rect 58876 626561 59196 633325
rect 58876 626325 58918 626561
rect 59154 626325 59196 626561
rect 58876 619561 59196 626325
rect 58876 619325 58918 619561
rect 59154 619325 59196 619561
rect 58876 612561 59196 619325
rect 58876 612325 58918 612561
rect 59154 612325 59196 612561
rect 58876 605561 59196 612325
rect 58876 605325 58918 605561
rect 59154 605325 59196 605561
rect 58876 598561 59196 605325
rect 58876 598325 58918 598561
rect 59154 598325 59196 598561
rect 58876 591561 59196 598325
rect 58876 591325 58918 591561
rect 59154 591325 59196 591561
rect 58876 584561 59196 591325
rect 58876 584325 58918 584561
rect 59154 584325 59196 584561
rect 58876 577561 59196 584325
rect 58876 577325 58918 577561
rect 59154 577325 59196 577561
rect 58876 570561 59196 577325
rect 58876 570325 58918 570561
rect 59154 570325 59196 570561
rect 58876 563561 59196 570325
rect 58876 563325 58918 563561
rect 59154 563325 59196 563561
rect 58876 556561 59196 563325
rect 58876 556325 58918 556561
rect 59154 556325 59196 556561
rect 58876 549561 59196 556325
rect 58876 549325 58918 549561
rect 59154 549325 59196 549561
rect 58876 542561 59196 549325
rect 58876 542325 58918 542561
rect 59154 542325 59196 542561
rect 58876 535561 59196 542325
rect 58876 535325 58918 535561
rect 59154 535325 59196 535561
rect 58876 528561 59196 535325
rect 58876 528325 58918 528561
rect 59154 528325 59196 528561
rect 58876 521561 59196 528325
rect 58876 521325 58918 521561
rect 59154 521325 59196 521561
rect 58876 514561 59196 521325
rect 58876 514325 58918 514561
rect 59154 514325 59196 514561
rect 58876 507561 59196 514325
rect 58876 507325 58918 507561
rect 59154 507325 59196 507561
rect 58876 500561 59196 507325
rect 58876 500325 58918 500561
rect 59154 500325 59196 500561
rect 58876 493561 59196 500325
rect 58876 493325 58918 493561
rect 59154 493325 59196 493561
rect 58876 486561 59196 493325
rect 58876 486325 58918 486561
rect 59154 486325 59196 486561
rect 58876 479561 59196 486325
rect 58876 479325 58918 479561
rect 59154 479325 59196 479561
rect 58876 472561 59196 479325
rect 58876 472325 58918 472561
rect 59154 472325 59196 472561
rect 58876 465561 59196 472325
rect 58876 465325 58918 465561
rect 59154 465325 59196 465561
rect 58876 458561 59196 465325
rect 58876 458325 58918 458561
rect 59154 458325 59196 458561
rect 58876 451561 59196 458325
rect 58876 451325 58918 451561
rect 59154 451325 59196 451561
rect 58876 444561 59196 451325
rect 58876 444325 58918 444561
rect 59154 444325 59196 444561
rect 58876 437561 59196 444325
rect 58876 437325 58918 437561
rect 59154 437325 59196 437561
rect 58876 430561 59196 437325
rect 58876 430325 58918 430561
rect 59154 430325 59196 430561
rect 58876 423561 59196 430325
rect 58876 423325 58918 423561
rect 59154 423325 59196 423561
rect 58876 416561 59196 423325
rect 58876 416325 58918 416561
rect 59154 416325 59196 416561
rect 58876 409561 59196 416325
rect 58876 409325 58918 409561
rect 59154 409325 59196 409561
rect 58876 402561 59196 409325
rect 58876 402325 58918 402561
rect 59154 402325 59196 402561
rect 58876 395561 59196 402325
rect 58876 395325 58918 395561
rect 59154 395325 59196 395561
rect 58876 388561 59196 395325
rect 58876 388325 58918 388561
rect 59154 388325 59196 388561
rect 58876 381561 59196 388325
rect 58876 381325 58918 381561
rect 59154 381325 59196 381561
rect 58876 374561 59196 381325
rect 58876 374325 58918 374561
rect 59154 374325 59196 374561
rect 58876 367561 59196 374325
rect 58876 367325 58918 367561
rect 59154 367325 59196 367561
rect 58876 360561 59196 367325
rect 58876 360325 58918 360561
rect 59154 360325 59196 360561
rect 58876 353561 59196 360325
rect 58876 353325 58918 353561
rect 59154 353325 59196 353561
rect 58876 346561 59196 353325
rect 58876 346325 58918 346561
rect 59154 346325 59196 346561
rect 58876 339561 59196 346325
rect 58876 339325 58918 339561
rect 59154 339325 59196 339561
rect 58876 332561 59196 339325
rect 58876 332325 58918 332561
rect 59154 332325 59196 332561
rect 58876 325561 59196 332325
rect 58876 325325 58918 325561
rect 59154 325325 59196 325561
rect 58876 318561 59196 325325
rect 58876 318325 58918 318561
rect 59154 318325 59196 318561
rect 58876 311561 59196 318325
rect 58876 311325 58918 311561
rect 59154 311325 59196 311561
rect 58876 304561 59196 311325
rect 58876 304325 58918 304561
rect 59154 304325 59196 304561
rect 58876 297561 59196 304325
rect 58876 297325 58918 297561
rect 59154 297325 59196 297561
rect 58876 290561 59196 297325
rect 58876 290325 58918 290561
rect 59154 290325 59196 290561
rect 58876 283561 59196 290325
rect 58876 283325 58918 283561
rect 59154 283325 59196 283561
rect 58876 276561 59196 283325
rect 58876 276325 58918 276561
rect 59154 276325 59196 276561
rect 58876 269561 59196 276325
rect 58876 269325 58918 269561
rect 59154 269325 59196 269561
rect 58876 262561 59196 269325
rect 58876 262325 58918 262561
rect 59154 262325 59196 262561
rect 58876 255561 59196 262325
rect 58876 255325 58918 255561
rect 59154 255325 59196 255561
rect 58876 248561 59196 255325
rect 58876 248325 58918 248561
rect 59154 248325 59196 248561
rect 58876 241561 59196 248325
rect 58876 241325 58918 241561
rect 59154 241325 59196 241561
rect 58876 234561 59196 241325
rect 58876 234325 58918 234561
rect 59154 234325 59196 234561
rect 58876 227561 59196 234325
rect 58876 227325 58918 227561
rect 59154 227325 59196 227561
rect 58876 220561 59196 227325
rect 58876 220325 58918 220561
rect 59154 220325 59196 220561
rect 58876 213561 59196 220325
rect 58876 213325 58918 213561
rect 59154 213325 59196 213561
rect 58876 206561 59196 213325
rect 58876 206325 58918 206561
rect 59154 206325 59196 206561
rect 58876 199561 59196 206325
rect 58876 199325 58918 199561
rect 59154 199325 59196 199561
rect 58876 192561 59196 199325
rect 58876 192325 58918 192561
rect 59154 192325 59196 192561
rect 58876 185561 59196 192325
rect 58876 185325 58918 185561
rect 59154 185325 59196 185561
rect 58876 178561 59196 185325
rect 58876 178325 58918 178561
rect 59154 178325 59196 178561
rect 58876 171561 59196 178325
rect 58876 171325 58918 171561
rect 59154 171325 59196 171561
rect 58876 164561 59196 171325
rect 58876 164325 58918 164561
rect 59154 164325 59196 164561
rect 58876 157561 59196 164325
rect 58876 157325 58918 157561
rect 59154 157325 59196 157561
rect 58876 150561 59196 157325
rect 58876 150325 58918 150561
rect 59154 150325 59196 150561
rect 58876 143561 59196 150325
rect 58876 143325 58918 143561
rect 59154 143325 59196 143561
rect 58876 136561 59196 143325
rect 58876 136325 58918 136561
rect 59154 136325 59196 136561
rect 58876 129561 59196 136325
rect 58876 129325 58918 129561
rect 59154 129325 59196 129561
rect 58876 122561 59196 129325
rect 58876 122325 58918 122561
rect 59154 122325 59196 122561
rect 58876 115561 59196 122325
rect 58876 115325 58918 115561
rect 59154 115325 59196 115561
rect 58876 108561 59196 115325
rect 58876 108325 58918 108561
rect 59154 108325 59196 108561
rect 58876 101561 59196 108325
rect 58876 101325 58918 101561
rect 59154 101325 59196 101561
rect 58876 94561 59196 101325
rect 58876 94325 58918 94561
rect 59154 94325 59196 94561
rect 58876 87561 59196 94325
rect 58876 87325 58918 87561
rect 59154 87325 59196 87561
rect 58876 80561 59196 87325
rect 58876 80325 58918 80561
rect 59154 80325 59196 80561
rect 58876 73561 59196 80325
rect 58876 73325 58918 73561
rect 59154 73325 59196 73561
rect 58876 66561 59196 73325
rect 58876 66325 58918 66561
rect 59154 66325 59196 66561
rect 58876 59561 59196 66325
rect 58876 59325 58918 59561
rect 59154 59325 59196 59561
rect 58876 52561 59196 59325
rect 58876 52325 58918 52561
rect 59154 52325 59196 52561
rect 58876 45561 59196 52325
rect 58876 45325 58918 45561
rect 59154 45325 59196 45561
rect 58876 38561 59196 45325
rect 58876 38325 58918 38561
rect 59154 38325 59196 38561
rect 58876 31561 59196 38325
rect 58876 31325 58918 31561
rect 59154 31325 59196 31561
rect 58876 24561 59196 31325
rect 58876 24325 58918 24561
rect 59154 24325 59196 24561
rect 58876 17561 59196 24325
rect 58876 17325 58918 17561
rect 59154 17325 59196 17561
rect 58876 10561 59196 17325
rect 58876 10325 58918 10561
rect 59154 10325 59196 10561
rect 58876 3561 59196 10325
rect 58876 3325 58918 3561
rect 59154 3325 59196 3561
rect 58876 -1706 59196 3325
rect 58876 -1942 58918 -1706
rect 59154 -1942 59196 -1706
rect 58876 -2026 59196 -1942
rect 58876 -2262 58918 -2026
rect 59154 -2262 59196 -2026
rect 58876 -2294 59196 -2262
rect 64144 705238 64464 706230
rect 64144 705002 64186 705238
rect 64422 705002 64464 705238
rect 64144 704918 64464 705002
rect 64144 704682 64186 704918
rect 64422 704682 64464 704918
rect 64144 695494 64464 704682
rect 64144 695258 64186 695494
rect 64422 695258 64464 695494
rect 64144 688494 64464 695258
rect 64144 688258 64186 688494
rect 64422 688258 64464 688494
rect 64144 681494 64464 688258
rect 64144 681258 64186 681494
rect 64422 681258 64464 681494
rect 64144 674494 64464 681258
rect 64144 674258 64186 674494
rect 64422 674258 64464 674494
rect 64144 667494 64464 674258
rect 64144 667258 64186 667494
rect 64422 667258 64464 667494
rect 64144 660494 64464 667258
rect 64144 660258 64186 660494
rect 64422 660258 64464 660494
rect 64144 653494 64464 660258
rect 64144 653258 64186 653494
rect 64422 653258 64464 653494
rect 64144 646494 64464 653258
rect 64144 646258 64186 646494
rect 64422 646258 64464 646494
rect 64144 639494 64464 646258
rect 64144 639258 64186 639494
rect 64422 639258 64464 639494
rect 64144 632494 64464 639258
rect 64144 632258 64186 632494
rect 64422 632258 64464 632494
rect 64144 625494 64464 632258
rect 64144 625258 64186 625494
rect 64422 625258 64464 625494
rect 64144 618494 64464 625258
rect 64144 618258 64186 618494
rect 64422 618258 64464 618494
rect 64144 611494 64464 618258
rect 64144 611258 64186 611494
rect 64422 611258 64464 611494
rect 64144 604494 64464 611258
rect 64144 604258 64186 604494
rect 64422 604258 64464 604494
rect 64144 597494 64464 604258
rect 64144 597258 64186 597494
rect 64422 597258 64464 597494
rect 64144 590494 64464 597258
rect 64144 590258 64186 590494
rect 64422 590258 64464 590494
rect 64144 583494 64464 590258
rect 64144 583258 64186 583494
rect 64422 583258 64464 583494
rect 64144 576494 64464 583258
rect 64144 576258 64186 576494
rect 64422 576258 64464 576494
rect 64144 569494 64464 576258
rect 64144 569258 64186 569494
rect 64422 569258 64464 569494
rect 64144 562494 64464 569258
rect 64144 562258 64186 562494
rect 64422 562258 64464 562494
rect 64144 555494 64464 562258
rect 64144 555258 64186 555494
rect 64422 555258 64464 555494
rect 64144 548494 64464 555258
rect 64144 548258 64186 548494
rect 64422 548258 64464 548494
rect 64144 541494 64464 548258
rect 64144 541258 64186 541494
rect 64422 541258 64464 541494
rect 64144 534494 64464 541258
rect 64144 534258 64186 534494
rect 64422 534258 64464 534494
rect 64144 527494 64464 534258
rect 64144 527258 64186 527494
rect 64422 527258 64464 527494
rect 64144 520494 64464 527258
rect 64144 520258 64186 520494
rect 64422 520258 64464 520494
rect 64144 513494 64464 520258
rect 64144 513258 64186 513494
rect 64422 513258 64464 513494
rect 64144 506494 64464 513258
rect 64144 506258 64186 506494
rect 64422 506258 64464 506494
rect 64144 499494 64464 506258
rect 64144 499258 64186 499494
rect 64422 499258 64464 499494
rect 64144 492494 64464 499258
rect 64144 492258 64186 492494
rect 64422 492258 64464 492494
rect 64144 485494 64464 492258
rect 64144 485258 64186 485494
rect 64422 485258 64464 485494
rect 64144 478494 64464 485258
rect 64144 478258 64186 478494
rect 64422 478258 64464 478494
rect 64144 471494 64464 478258
rect 64144 471258 64186 471494
rect 64422 471258 64464 471494
rect 64144 464494 64464 471258
rect 64144 464258 64186 464494
rect 64422 464258 64464 464494
rect 64144 457494 64464 464258
rect 64144 457258 64186 457494
rect 64422 457258 64464 457494
rect 64144 450494 64464 457258
rect 64144 450258 64186 450494
rect 64422 450258 64464 450494
rect 64144 443494 64464 450258
rect 64144 443258 64186 443494
rect 64422 443258 64464 443494
rect 64144 436494 64464 443258
rect 64144 436258 64186 436494
rect 64422 436258 64464 436494
rect 64144 429494 64464 436258
rect 64144 429258 64186 429494
rect 64422 429258 64464 429494
rect 64144 422494 64464 429258
rect 64144 422258 64186 422494
rect 64422 422258 64464 422494
rect 64144 415494 64464 422258
rect 64144 415258 64186 415494
rect 64422 415258 64464 415494
rect 64144 408494 64464 415258
rect 64144 408258 64186 408494
rect 64422 408258 64464 408494
rect 64144 401494 64464 408258
rect 64144 401258 64186 401494
rect 64422 401258 64464 401494
rect 64144 394494 64464 401258
rect 64144 394258 64186 394494
rect 64422 394258 64464 394494
rect 64144 387494 64464 394258
rect 64144 387258 64186 387494
rect 64422 387258 64464 387494
rect 64144 380494 64464 387258
rect 64144 380258 64186 380494
rect 64422 380258 64464 380494
rect 64144 373494 64464 380258
rect 64144 373258 64186 373494
rect 64422 373258 64464 373494
rect 64144 366494 64464 373258
rect 64144 366258 64186 366494
rect 64422 366258 64464 366494
rect 64144 359494 64464 366258
rect 64144 359258 64186 359494
rect 64422 359258 64464 359494
rect 64144 352494 64464 359258
rect 64144 352258 64186 352494
rect 64422 352258 64464 352494
rect 64144 345494 64464 352258
rect 64144 345258 64186 345494
rect 64422 345258 64464 345494
rect 64144 338494 64464 345258
rect 64144 338258 64186 338494
rect 64422 338258 64464 338494
rect 64144 331494 64464 338258
rect 64144 331258 64186 331494
rect 64422 331258 64464 331494
rect 64144 324494 64464 331258
rect 64144 324258 64186 324494
rect 64422 324258 64464 324494
rect 64144 317494 64464 324258
rect 64144 317258 64186 317494
rect 64422 317258 64464 317494
rect 64144 310494 64464 317258
rect 64144 310258 64186 310494
rect 64422 310258 64464 310494
rect 64144 303494 64464 310258
rect 64144 303258 64186 303494
rect 64422 303258 64464 303494
rect 64144 296494 64464 303258
rect 64144 296258 64186 296494
rect 64422 296258 64464 296494
rect 64144 289494 64464 296258
rect 64144 289258 64186 289494
rect 64422 289258 64464 289494
rect 64144 282494 64464 289258
rect 64144 282258 64186 282494
rect 64422 282258 64464 282494
rect 64144 275494 64464 282258
rect 64144 275258 64186 275494
rect 64422 275258 64464 275494
rect 64144 268494 64464 275258
rect 64144 268258 64186 268494
rect 64422 268258 64464 268494
rect 64144 261494 64464 268258
rect 64144 261258 64186 261494
rect 64422 261258 64464 261494
rect 64144 254494 64464 261258
rect 64144 254258 64186 254494
rect 64422 254258 64464 254494
rect 64144 247494 64464 254258
rect 64144 247258 64186 247494
rect 64422 247258 64464 247494
rect 64144 240494 64464 247258
rect 64144 240258 64186 240494
rect 64422 240258 64464 240494
rect 64144 233494 64464 240258
rect 64144 233258 64186 233494
rect 64422 233258 64464 233494
rect 64144 226494 64464 233258
rect 64144 226258 64186 226494
rect 64422 226258 64464 226494
rect 64144 219494 64464 226258
rect 64144 219258 64186 219494
rect 64422 219258 64464 219494
rect 64144 212494 64464 219258
rect 64144 212258 64186 212494
rect 64422 212258 64464 212494
rect 64144 205494 64464 212258
rect 64144 205258 64186 205494
rect 64422 205258 64464 205494
rect 64144 198494 64464 205258
rect 64144 198258 64186 198494
rect 64422 198258 64464 198494
rect 64144 191494 64464 198258
rect 64144 191258 64186 191494
rect 64422 191258 64464 191494
rect 64144 184494 64464 191258
rect 64144 184258 64186 184494
rect 64422 184258 64464 184494
rect 64144 177494 64464 184258
rect 64144 177258 64186 177494
rect 64422 177258 64464 177494
rect 64144 170494 64464 177258
rect 64144 170258 64186 170494
rect 64422 170258 64464 170494
rect 64144 163494 64464 170258
rect 64144 163258 64186 163494
rect 64422 163258 64464 163494
rect 64144 156494 64464 163258
rect 64144 156258 64186 156494
rect 64422 156258 64464 156494
rect 64144 149494 64464 156258
rect 64144 149258 64186 149494
rect 64422 149258 64464 149494
rect 64144 142494 64464 149258
rect 64144 142258 64186 142494
rect 64422 142258 64464 142494
rect 64144 135494 64464 142258
rect 64144 135258 64186 135494
rect 64422 135258 64464 135494
rect 64144 128494 64464 135258
rect 64144 128258 64186 128494
rect 64422 128258 64464 128494
rect 64144 121494 64464 128258
rect 64144 121258 64186 121494
rect 64422 121258 64464 121494
rect 64144 114494 64464 121258
rect 64144 114258 64186 114494
rect 64422 114258 64464 114494
rect 64144 107494 64464 114258
rect 64144 107258 64186 107494
rect 64422 107258 64464 107494
rect 64144 100494 64464 107258
rect 64144 100258 64186 100494
rect 64422 100258 64464 100494
rect 64144 93494 64464 100258
rect 64144 93258 64186 93494
rect 64422 93258 64464 93494
rect 64144 86494 64464 93258
rect 64144 86258 64186 86494
rect 64422 86258 64464 86494
rect 64144 79494 64464 86258
rect 64144 79258 64186 79494
rect 64422 79258 64464 79494
rect 64144 72494 64464 79258
rect 64144 72258 64186 72494
rect 64422 72258 64464 72494
rect 64144 65494 64464 72258
rect 64144 65258 64186 65494
rect 64422 65258 64464 65494
rect 64144 58494 64464 65258
rect 64144 58258 64186 58494
rect 64422 58258 64464 58494
rect 64144 51494 64464 58258
rect 64144 51258 64186 51494
rect 64422 51258 64464 51494
rect 64144 44494 64464 51258
rect 64144 44258 64186 44494
rect 64422 44258 64464 44494
rect 64144 37494 64464 44258
rect 64144 37258 64186 37494
rect 64422 37258 64464 37494
rect 64144 30494 64464 37258
rect 64144 30258 64186 30494
rect 64422 30258 64464 30494
rect 64144 23494 64464 30258
rect 64144 23258 64186 23494
rect 64422 23258 64464 23494
rect 64144 16494 64464 23258
rect 64144 16258 64186 16494
rect 64422 16258 64464 16494
rect 64144 9494 64464 16258
rect 64144 9258 64186 9494
rect 64422 9258 64464 9494
rect 64144 2494 64464 9258
rect 64144 2258 64186 2494
rect 64422 2258 64464 2494
rect 64144 -746 64464 2258
rect 64144 -982 64186 -746
rect 64422 -982 64464 -746
rect 64144 -1066 64464 -982
rect 64144 -1302 64186 -1066
rect 64422 -1302 64464 -1066
rect 64144 -2294 64464 -1302
rect 65876 706198 66196 706230
rect 65876 705962 65918 706198
rect 66154 705962 66196 706198
rect 65876 705878 66196 705962
rect 65876 705642 65918 705878
rect 66154 705642 66196 705878
rect 65876 696561 66196 705642
rect 65876 696325 65918 696561
rect 66154 696325 66196 696561
rect 65876 689561 66196 696325
rect 65876 689325 65918 689561
rect 66154 689325 66196 689561
rect 65876 682561 66196 689325
rect 65876 682325 65918 682561
rect 66154 682325 66196 682561
rect 65876 675561 66196 682325
rect 65876 675325 65918 675561
rect 66154 675325 66196 675561
rect 65876 668561 66196 675325
rect 65876 668325 65918 668561
rect 66154 668325 66196 668561
rect 65876 661561 66196 668325
rect 65876 661325 65918 661561
rect 66154 661325 66196 661561
rect 65876 654561 66196 661325
rect 65876 654325 65918 654561
rect 66154 654325 66196 654561
rect 65876 647561 66196 654325
rect 65876 647325 65918 647561
rect 66154 647325 66196 647561
rect 65876 640561 66196 647325
rect 65876 640325 65918 640561
rect 66154 640325 66196 640561
rect 65876 633561 66196 640325
rect 65876 633325 65918 633561
rect 66154 633325 66196 633561
rect 65876 626561 66196 633325
rect 65876 626325 65918 626561
rect 66154 626325 66196 626561
rect 65876 619561 66196 626325
rect 65876 619325 65918 619561
rect 66154 619325 66196 619561
rect 65876 612561 66196 619325
rect 65876 612325 65918 612561
rect 66154 612325 66196 612561
rect 65876 605561 66196 612325
rect 65876 605325 65918 605561
rect 66154 605325 66196 605561
rect 65876 598561 66196 605325
rect 65876 598325 65918 598561
rect 66154 598325 66196 598561
rect 65876 591561 66196 598325
rect 65876 591325 65918 591561
rect 66154 591325 66196 591561
rect 65876 584561 66196 591325
rect 65876 584325 65918 584561
rect 66154 584325 66196 584561
rect 65876 577561 66196 584325
rect 65876 577325 65918 577561
rect 66154 577325 66196 577561
rect 65876 570561 66196 577325
rect 65876 570325 65918 570561
rect 66154 570325 66196 570561
rect 65876 563561 66196 570325
rect 65876 563325 65918 563561
rect 66154 563325 66196 563561
rect 65876 556561 66196 563325
rect 65876 556325 65918 556561
rect 66154 556325 66196 556561
rect 65876 549561 66196 556325
rect 65876 549325 65918 549561
rect 66154 549325 66196 549561
rect 65876 542561 66196 549325
rect 65876 542325 65918 542561
rect 66154 542325 66196 542561
rect 65876 535561 66196 542325
rect 65876 535325 65918 535561
rect 66154 535325 66196 535561
rect 65876 528561 66196 535325
rect 65876 528325 65918 528561
rect 66154 528325 66196 528561
rect 65876 521561 66196 528325
rect 65876 521325 65918 521561
rect 66154 521325 66196 521561
rect 65876 514561 66196 521325
rect 65876 514325 65918 514561
rect 66154 514325 66196 514561
rect 65876 507561 66196 514325
rect 65876 507325 65918 507561
rect 66154 507325 66196 507561
rect 65876 500561 66196 507325
rect 65876 500325 65918 500561
rect 66154 500325 66196 500561
rect 65876 493561 66196 500325
rect 65876 493325 65918 493561
rect 66154 493325 66196 493561
rect 65876 486561 66196 493325
rect 65876 486325 65918 486561
rect 66154 486325 66196 486561
rect 65876 479561 66196 486325
rect 65876 479325 65918 479561
rect 66154 479325 66196 479561
rect 65876 472561 66196 479325
rect 65876 472325 65918 472561
rect 66154 472325 66196 472561
rect 65876 465561 66196 472325
rect 65876 465325 65918 465561
rect 66154 465325 66196 465561
rect 65876 458561 66196 465325
rect 65876 458325 65918 458561
rect 66154 458325 66196 458561
rect 65876 451561 66196 458325
rect 65876 451325 65918 451561
rect 66154 451325 66196 451561
rect 65876 444561 66196 451325
rect 65876 444325 65918 444561
rect 66154 444325 66196 444561
rect 65876 437561 66196 444325
rect 65876 437325 65918 437561
rect 66154 437325 66196 437561
rect 65876 430561 66196 437325
rect 65876 430325 65918 430561
rect 66154 430325 66196 430561
rect 65876 423561 66196 430325
rect 65876 423325 65918 423561
rect 66154 423325 66196 423561
rect 65876 416561 66196 423325
rect 65876 416325 65918 416561
rect 66154 416325 66196 416561
rect 65876 409561 66196 416325
rect 65876 409325 65918 409561
rect 66154 409325 66196 409561
rect 65876 402561 66196 409325
rect 65876 402325 65918 402561
rect 66154 402325 66196 402561
rect 65876 395561 66196 402325
rect 65876 395325 65918 395561
rect 66154 395325 66196 395561
rect 65876 388561 66196 395325
rect 65876 388325 65918 388561
rect 66154 388325 66196 388561
rect 65876 381561 66196 388325
rect 65876 381325 65918 381561
rect 66154 381325 66196 381561
rect 65876 374561 66196 381325
rect 65876 374325 65918 374561
rect 66154 374325 66196 374561
rect 65876 367561 66196 374325
rect 65876 367325 65918 367561
rect 66154 367325 66196 367561
rect 65876 360561 66196 367325
rect 65876 360325 65918 360561
rect 66154 360325 66196 360561
rect 65876 353561 66196 360325
rect 65876 353325 65918 353561
rect 66154 353325 66196 353561
rect 65876 346561 66196 353325
rect 65876 346325 65918 346561
rect 66154 346325 66196 346561
rect 65876 339561 66196 346325
rect 65876 339325 65918 339561
rect 66154 339325 66196 339561
rect 65876 332561 66196 339325
rect 65876 332325 65918 332561
rect 66154 332325 66196 332561
rect 65876 325561 66196 332325
rect 65876 325325 65918 325561
rect 66154 325325 66196 325561
rect 65876 318561 66196 325325
rect 65876 318325 65918 318561
rect 66154 318325 66196 318561
rect 65876 311561 66196 318325
rect 65876 311325 65918 311561
rect 66154 311325 66196 311561
rect 65876 304561 66196 311325
rect 65876 304325 65918 304561
rect 66154 304325 66196 304561
rect 65876 297561 66196 304325
rect 65876 297325 65918 297561
rect 66154 297325 66196 297561
rect 65876 290561 66196 297325
rect 65876 290325 65918 290561
rect 66154 290325 66196 290561
rect 65876 283561 66196 290325
rect 65876 283325 65918 283561
rect 66154 283325 66196 283561
rect 65876 276561 66196 283325
rect 65876 276325 65918 276561
rect 66154 276325 66196 276561
rect 65876 269561 66196 276325
rect 65876 269325 65918 269561
rect 66154 269325 66196 269561
rect 65876 262561 66196 269325
rect 65876 262325 65918 262561
rect 66154 262325 66196 262561
rect 65876 255561 66196 262325
rect 65876 255325 65918 255561
rect 66154 255325 66196 255561
rect 65876 248561 66196 255325
rect 65876 248325 65918 248561
rect 66154 248325 66196 248561
rect 65876 241561 66196 248325
rect 65876 241325 65918 241561
rect 66154 241325 66196 241561
rect 65876 234561 66196 241325
rect 65876 234325 65918 234561
rect 66154 234325 66196 234561
rect 65876 227561 66196 234325
rect 65876 227325 65918 227561
rect 66154 227325 66196 227561
rect 65876 220561 66196 227325
rect 65876 220325 65918 220561
rect 66154 220325 66196 220561
rect 65876 213561 66196 220325
rect 65876 213325 65918 213561
rect 66154 213325 66196 213561
rect 65876 206561 66196 213325
rect 65876 206325 65918 206561
rect 66154 206325 66196 206561
rect 65876 199561 66196 206325
rect 65876 199325 65918 199561
rect 66154 199325 66196 199561
rect 65876 192561 66196 199325
rect 65876 192325 65918 192561
rect 66154 192325 66196 192561
rect 65876 185561 66196 192325
rect 65876 185325 65918 185561
rect 66154 185325 66196 185561
rect 65876 178561 66196 185325
rect 65876 178325 65918 178561
rect 66154 178325 66196 178561
rect 65876 171561 66196 178325
rect 65876 171325 65918 171561
rect 66154 171325 66196 171561
rect 65876 164561 66196 171325
rect 65876 164325 65918 164561
rect 66154 164325 66196 164561
rect 65876 157561 66196 164325
rect 65876 157325 65918 157561
rect 66154 157325 66196 157561
rect 65876 150561 66196 157325
rect 65876 150325 65918 150561
rect 66154 150325 66196 150561
rect 65876 143561 66196 150325
rect 65876 143325 65918 143561
rect 66154 143325 66196 143561
rect 65876 136561 66196 143325
rect 65876 136325 65918 136561
rect 66154 136325 66196 136561
rect 65876 129561 66196 136325
rect 65876 129325 65918 129561
rect 66154 129325 66196 129561
rect 65876 122561 66196 129325
rect 65876 122325 65918 122561
rect 66154 122325 66196 122561
rect 65876 115561 66196 122325
rect 65876 115325 65918 115561
rect 66154 115325 66196 115561
rect 65876 108561 66196 115325
rect 65876 108325 65918 108561
rect 66154 108325 66196 108561
rect 65876 101561 66196 108325
rect 65876 101325 65918 101561
rect 66154 101325 66196 101561
rect 65876 94561 66196 101325
rect 65876 94325 65918 94561
rect 66154 94325 66196 94561
rect 65876 87561 66196 94325
rect 65876 87325 65918 87561
rect 66154 87325 66196 87561
rect 65876 80561 66196 87325
rect 65876 80325 65918 80561
rect 66154 80325 66196 80561
rect 65876 73561 66196 80325
rect 65876 73325 65918 73561
rect 66154 73325 66196 73561
rect 65876 66561 66196 73325
rect 65876 66325 65918 66561
rect 66154 66325 66196 66561
rect 65876 59561 66196 66325
rect 65876 59325 65918 59561
rect 66154 59325 66196 59561
rect 65876 52561 66196 59325
rect 65876 52325 65918 52561
rect 66154 52325 66196 52561
rect 65876 45561 66196 52325
rect 65876 45325 65918 45561
rect 66154 45325 66196 45561
rect 65876 38561 66196 45325
rect 65876 38325 65918 38561
rect 66154 38325 66196 38561
rect 65876 31561 66196 38325
rect 65876 31325 65918 31561
rect 66154 31325 66196 31561
rect 65876 24561 66196 31325
rect 65876 24325 65918 24561
rect 66154 24325 66196 24561
rect 65876 17561 66196 24325
rect 65876 17325 65918 17561
rect 66154 17325 66196 17561
rect 65876 10561 66196 17325
rect 65876 10325 65918 10561
rect 66154 10325 66196 10561
rect 65876 3561 66196 10325
rect 65876 3325 65918 3561
rect 66154 3325 66196 3561
rect 65876 -1706 66196 3325
rect 65876 -1942 65918 -1706
rect 66154 -1942 66196 -1706
rect 65876 -2026 66196 -1942
rect 65876 -2262 65918 -2026
rect 66154 -2262 66196 -2026
rect 65876 -2294 66196 -2262
rect 71144 705238 71464 706230
rect 71144 705002 71186 705238
rect 71422 705002 71464 705238
rect 71144 704918 71464 705002
rect 71144 704682 71186 704918
rect 71422 704682 71464 704918
rect 71144 695494 71464 704682
rect 71144 695258 71186 695494
rect 71422 695258 71464 695494
rect 71144 688494 71464 695258
rect 71144 688258 71186 688494
rect 71422 688258 71464 688494
rect 71144 681494 71464 688258
rect 71144 681258 71186 681494
rect 71422 681258 71464 681494
rect 71144 674494 71464 681258
rect 71144 674258 71186 674494
rect 71422 674258 71464 674494
rect 71144 667494 71464 674258
rect 71144 667258 71186 667494
rect 71422 667258 71464 667494
rect 71144 660494 71464 667258
rect 71144 660258 71186 660494
rect 71422 660258 71464 660494
rect 71144 653494 71464 660258
rect 71144 653258 71186 653494
rect 71422 653258 71464 653494
rect 71144 646494 71464 653258
rect 71144 646258 71186 646494
rect 71422 646258 71464 646494
rect 71144 639494 71464 646258
rect 71144 639258 71186 639494
rect 71422 639258 71464 639494
rect 71144 632494 71464 639258
rect 71144 632258 71186 632494
rect 71422 632258 71464 632494
rect 71144 625494 71464 632258
rect 71144 625258 71186 625494
rect 71422 625258 71464 625494
rect 71144 618494 71464 625258
rect 71144 618258 71186 618494
rect 71422 618258 71464 618494
rect 71144 611494 71464 618258
rect 71144 611258 71186 611494
rect 71422 611258 71464 611494
rect 71144 604494 71464 611258
rect 71144 604258 71186 604494
rect 71422 604258 71464 604494
rect 71144 597494 71464 604258
rect 71144 597258 71186 597494
rect 71422 597258 71464 597494
rect 71144 590494 71464 597258
rect 71144 590258 71186 590494
rect 71422 590258 71464 590494
rect 71144 583494 71464 590258
rect 71144 583258 71186 583494
rect 71422 583258 71464 583494
rect 71144 576494 71464 583258
rect 71144 576258 71186 576494
rect 71422 576258 71464 576494
rect 71144 569494 71464 576258
rect 71144 569258 71186 569494
rect 71422 569258 71464 569494
rect 71144 562494 71464 569258
rect 71144 562258 71186 562494
rect 71422 562258 71464 562494
rect 71144 555494 71464 562258
rect 71144 555258 71186 555494
rect 71422 555258 71464 555494
rect 71144 548494 71464 555258
rect 71144 548258 71186 548494
rect 71422 548258 71464 548494
rect 71144 541494 71464 548258
rect 71144 541258 71186 541494
rect 71422 541258 71464 541494
rect 71144 534494 71464 541258
rect 71144 534258 71186 534494
rect 71422 534258 71464 534494
rect 71144 527494 71464 534258
rect 71144 527258 71186 527494
rect 71422 527258 71464 527494
rect 71144 520494 71464 527258
rect 71144 520258 71186 520494
rect 71422 520258 71464 520494
rect 71144 513494 71464 520258
rect 71144 513258 71186 513494
rect 71422 513258 71464 513494
rect 71144 506494 71464 513258
rect 71144 506258 71186 506494
rect 71422 506258 71464 506494
rect 71144 499494 71464 506258
rect 71144 499258 71186 499494
rect 71422 499258 71464 499494
rect 71144 492494 71464 499258
rect 71144 492258 71186 492494
rect 71422 492258 71464 492494
rect 71144 485494 71464 492258
rect 71144 485258 71186 485494
rect 71422 485258 71464 485494
rect 71144 478494 71464 485258
rect 71144 478258 71186 478494
rect 71422 478258 71464 478494
rect 71144 471494 71464 478258
rect 71144 471258 71186 471494
rect 71422 471258 71464 471494
rect 71144 464494 71464 471258
rect 71144 464258 71186 464494
rect 71422 464258 71464 464494
rect 71144 457494 71464 464258
rect 71144 457258 71186 457494
rect 71422 457258 71464 457494
rect 71144 450494 71464 457258
rect 71144 450258 71186 450494
rect 71422 450258 71464 450494
rect 71144 443494 71464 450258
rect 71144 443258 71186 443494
rect 71422 443258 71464 443494
rect 71144 436494 71464 443258
rect 71144 436258 71186 436494
rect 71422 436258 71464 436494
rect 71144 429494 71464 436258
rect 71144 429258 71186 429494
rect 71422 429258 71464 429494
rect 71144 422494 71464 429258
rect 71144 422258 71186 422494
rect 71422 422258 71464 422494
rect 71144 415494 71464 422258
rect 71144 415258 71186 415494
rect 71422 415258 71464 415494
rect 71144 408494 71464 415258
rect 71144 408258 71186 408494
rect 71422 408258 71464 408494
rect 71144 401494 71464 408258
rect 71144 401258 71186 401494
rect 71422 401258 71464 401494
rect 71144 394494 71464 401258
rect 71144 394258 71186 394494
rect 71422 394258 71464 394494
rect 71144 387494 71464 394258
rect 71144 387258 71186 387494
rect 71422 387258 71464 387494
rect 71144 380494 71464 387258
rect 71144 380258 71186 380494
rect 71422 380258 71464 380494
rect 71144 373494 71464 380258
rect 71144 373258 71186 373494
rect 71422 373258 71464 373494
rect 71144 366494 71464 373258
rect 71144 366258 71186 366494
rect 71422 366258 71464 366494
rect 71144 359494 71464 366258
rect 71144 359258 71186 359494
rect 71422 359258 71464 359494
rect 71144 352494 71464 359258
rect 71144 352258 71186 352494
rect 71422 352258 71464 352494
rect 71144 345494 71464 352258
rect 71144 345258 71186 345494
rect 71422 345258 71464 345494
rect 71144 338494 71464 345258
rect 71144 338258 71186 338494
rect 71422 338258 71464 338494
rect 71144 331494 71464 338258
rect 71144 331258 71186 331494
rect 71422 331258 71464 331494
rect 71144 324494 71464 331258
rect 71144 324258 71186 324494
rect 71422 324258 71464 324494
rect 71144 317494 71464 324258
rect 71144 317258 71186 317494
rect 71422 317258 71464 317494
rect 71144 310494 71464 317258
rect 71144 310258 71186 310494
rect 71422 310258 71464 310494
rect 71144 303494 71464 310258
rect 71144 303258 71186 303494
rect 71422 303258 71464 303494
rect 71144 296494 71464 303258
rect 71144 296258 71186 296494
rect 71422 296258 71464 296494
rect 71144 289494 71464 296258
rect 71144 289258 71186 289494
rect 71422 289258 71464 289494
rect 71144 282494 71464 289258
rect 71144 282258 71186 282494
rect 71422 282258 71464 282494
rect 71144 275494 71464 282258
rect 71144 275258 71186 275494
rect 71422 275258 71464 275494
rect 71144 268494 71464 275258
rect 71144 268258 71186 268494
rect 71422 268258 71464 268494
rect 71144 261494 71464 268258
rect 71144 261258 71186 261494
rect 71422 261258 71464 261494
rect 71144 254494 71464 261258
rect 71144 254258 71186 254494
rect 71422 254258 71464 254494
rect 71144 247494 71464 254258
rect 71144 247258 71186 247494
rect 71422 247258 71464 247494
rect 71144 240494 71464 247258
rect 71144 240258 71186 240494
rect 71422 240258 71464 240494
rect 71144 233494 71464 240258
rect 71144 233258 71186 233494
rect 71422 233258 71464 233494
rect 71144 226494 71464 233258
rect 71144 226258 71186 226494
rect 71422 226258 71464 226494
rect 71144 219494 71464 226258
rect 71144 219258 71186 219494
rect 71422 219258 71464 219494
rect 71144 212494 71464 219258
rect 71144 212258 71186 212494
rect 71422 212258 71464 212494
rect 71144 205494 71464 212258
rect 71144 205258 71186 205494
rect 71422 205258 71464 205494
rect 71144 198494 71464 205258
rect 71144 198258 71186 198494
rect 71422 198258 71464 198494
rect 71144 191494 71464 198258
rect 71144 191258 71186 191494
rect 71422 191258 71464 191494
rect 71144 184494 71464 191258
rect 71144 184258 71186 184494
rect 71422 184258 71464 184494
rect 71144 177494 71464 184258
rect 71144 177258 71186 177494
rect 71422 177258 71464 177494
rect 71144 170494 71464 177258
rect 71144 170258 71186 170494
rect 71422 170258 71464 170494
rect 71144 163494 71464 170258
rect 71144 163258 71186 163494
rect 71422 163258 71464 163494
rect 71144 156494 71464 163258
rect 71144 156258 71186 156494
rect 71422 156258 71464 156494
rect 71144 149494 71464 156258
rect 71144 149258 71186 149494
rect 71422 149258 71464 149494
rect 71144 142494 71464 149258
rect 71144 142258 71186 142494
rect 71422 142258 71464 142494
rect 71144 135494 71464 142258
rect 71144 135258 71186 135494
rect 71422 135258 71464 135494
rect 71144 128494 71464 135258
rect 71144 128258 71186 128494
rect 71422 128258 71464 128494
rect 71144 121494 71464 128258
rect 71144 121258 71186 121494
rect 71422 121258 71464 121494
rect 71144 114494 71464 121258
rect 71144 114258 71186 114494
rect 71422 114258 71464 114494
rect 71144 107494 71464 114258
rect 71144 107258 71186 107494
rect 71422 107258 71464 107494
rect 71144 100494 71464 107258
rect 71144 100258 71186 100494
rect 71422 100258 71464 100494
rect 71144 93494 71464 100258
rect 71144 93258 71186 93494
rect 71422 93258 71464 93494
rect 71144 86494 71464 93258
rect 71144 86258 71186 86494
rect 71422 86258 71464 86494
rect 71144 79494 71464 86258
rect 71144 79258 71186 79494
rect 71422 79258 71464 79494
rect 71144 72494 71464 79258
rect 71144 72258 71186 72494
rect 71422 72258 71464 72494
rect 71144 65494 71464 72258
rect 71144 65258 71186 65494
rect 71422 65258 71464 65494
rect 71144 58494 71464 65258
rect 71144 58258 71186 58494
rect 71422 58258 71464 58494
rect 71144 51494 71464 58258
rect 71144 51258 71186 51494
rect 71422 51258 71464 51494
rect 71144 44494 71464 51258
rect 71144 44258 71186 44494
rect 71422 44258 71464 44494
rect 71144 37494 71464 44258
rect 71144 37258 71186 37494
rect 71422 37258 71464 37494
rect 71144 30494 71464 37258
rect 71144 30258 71186 30494
rect 71422 30258 71464 30494
rect 71144 23494 71464 30258
rect 71144 23258 71186 23494
rect 71422 23258 71464 23494
rect 71144 16494 71464 23258
rect 71144 16258 71186 16494
rect 71422 16258 71464 16494
rect 71144 9494 71464 16258
rect 71144 9258 71186 9494
rect 71422 9258 71464 9494
rect 71144 2494 71464 9258
rect 71144 2258 71186 2494
rect 71422 2258 71464 2494
rect 71144 -746 71464 2258
rect 71144 -982 71186 -746
rect 71422 -982 71464 -746
rect 71144 -1066 71464 -982
rect 71144 -1302 71186 -1066
rect 71422 -1302 71464 -1066
rect 71144 -2294 71464 -1302
rect 72876 706198 73196 706230
rect 72876 705962 72918 706198
rect 73154 705962 73196 706198
rect 72876 705878 73196 705962
rect 72876 705642 72918 705878
rect 73154 705642 73196 705878
rect 72876 696561 73196 705642
rect 72876 696325 72918 696561
rect 73154 696325 73196 696561
rect 72876 689561 73196 696325
rect 72876 689325 72918 689561
rect 73154 689325 73196 689561
rect 72876 682561 73196 689325
rect 72876 682325 72918 682561
rect 73154 682325 73196 682561
rect 72876 675561 73196 682325
rect 72876 675325 72918 675561
rect 73154 675325 73196 675561
rect 72876 668561 73196 675325
rect 72876 668325 72918 668561
rect 73154 668325 73196 668561
rect 72876 661561 73196 668325
rect 72876 661325 72918 661561
rect 73154 661325 73196 661561
rect 72876 654561 73196 661325
rect 72876 654325 72918 654561
rect 73154 654325 73196 654561
rect 72876 647561 73196 654325
rect 72876 647325 72918 647561
rect 73154 647325 73196 647561
rect 72876 640561 73196 647325
rect 72876 640325 72918 640561
rect 73154 640325 73196 640561
rect 72876 633561 73196 640325
rect 72876 633325 72918 633561
rect 73154 633325 73196 633561
rect 72876 626561 73196 633325
rect 72876 626325 72918 626561
rect 73154 626325 73196 626561
rect 72876 619561 73196 626325
rect 72876 619325 72918 619561
rect 73154 619325 73196 619561
rect 72876 612561 73196 619325
rect 72876 612325 72918 612561
rect 73154 612325 73196 612561
rect 72876 605561 73196 612325
rect 72876 605325 72918 605561
rect 73154 605325 73196 605561
rect 72876 598561 73196 605325
rect 72876 598325 72918 598561
rect 73154 598325 73196 598561
rect 72876 591561 73196 598325
rect 72876 591325 72918 591561
rect 73154 591325 73196 591561
rect 72876 584561 73196 591325
rect 72876 584325 72918 584561
rect 73154 584325 73196 584561
rect 72876 577561 73196 584325
rect 72876 577325 72918 577561
rect 73154 577325 73196 577561
rect 72876 570561 73196 577325
rect 72876 570325 72918 570561
rect 73154 570325 73196 570561
rect 72876 563561 73196 570325
rect 72876 563325 72918 563561
rect 73154 563325 73196 563561
rect 72876 556561 73196 563325
rect 72876 556325 72918 556561
rect 73154 556325 73196 556561
rect 72876 549561 73196 556325
rect 72876 549325 72918 549561
rect 73154 549325 73196 549561
rect 72876 542561 73196 549325
rect 72876 542325 72918 542561
rect 73154 542325 73196 542561
rect 72876 535561 73196 542325
rect 72876 535325 72918 535561
rect 73154 535325 73196 535561
rect 72876 528561 73196 535325
rect 72876 528325 72918 528561
rect 73154 528325 73196 528561
rect 72876 521561 73196 528325
rect 72876 521325 72918 521561
rect 73154 521325 73196 521561
rect 72876 514561 73196 521325
rect 72876 514325 72918 514561
rect 73154 514325 73196 514561
rect 72876 507561 73196 514325
rect 72876 507325 72918 507561
rect 73154 507325 73196 507561
rect 72876 500561 73196 507325
rect 72876 500325 72918 500561
rect 73154 500325 73196 500561
rect 72876 493561 73196 500325
rect 72876 493325 72918 493561
rect 73154 493325 73196 493561
rect 72876 486561 73196 493325
rect 72876 486325 72918 486561
rect 73154 486325 73196 486561
rect 72876 479561 73196 486325
rect 72876 479325 72918 479561
rect 73154 479325 73196 479561
rect 72876 472561 73196 479325
rect 72876 472325 72918 472561
rect 73154 472325 73196 472561
rect 72876 465561 73196 472325
rect 72876 465325 72918 465561
rect 73154 465325 73196 465561
rect 72876 458561 73196 465325
rect 72876 458325 72918 458561
rect 73154 458325 73196 458561
rect 72876 451561 73196 458325
rect 72876 451325 72918 451561
rect 73154 451325 73196 451561
rect 72876 444561 73196 451325
rect 72876 444325 72918 444561
rect 73154 444325 73196 444561
rect 72876 437561 73196 444325
rect 72876 437325 72918 437561
rect 73154 437325 73196 437561
rect 72876 430561 73196 437325
rect 72876 430325 72918 430561
rect 73154 430325 73196 430561
rect 72876 423561 73196 430325
rect 72876 423325 72918 423561
rect 73154 423325 73196 423561
rect 72876 416561 73196 423325
rect 72876 416325 72918 416561
rect 73154 416325 73196 416561
rect 72876 409561 73196 416325
rect 72876 409325 72918 409561
rect 73154 409325 73196 409561
rect 72876 402561 73196 409325
rect 72876 402325 72918 402561
rect 73154 402325 73196 402561
rect 72876 395561 73196 402325
rect 72876 395325 72918 395561
rect 73154 395325 73196 395561
rect 72876 388561 73196 395325
rect 72876 388325 72918 388561
rect 73154 388325 73196 388561
rect 72876 381561 73196 388325
rect 72876 381325 72918 381561
rect 73154 381325 73196 381561
rect 72876 374561 73196 381325
rect 72876 374325 72918 374561
rect 73154 374325 73196 374561
rect 72876 367561 73196 374325
rect 72876 367325 72918 367561
rect 73154 367325 73196 367561
rect 72876 360561 73196 367325
rect 72876 360325 72918 360561
rect 73154 360325 73196 360561
rect 72876 353561 73196 360325
rect 72876 353325 72918 353561
rect 73154 353325 73196 353561
rect 72876 346561 73196 353325
rect 72876 346325 72918 346561
rect 73154 346325 73196 346561
rect 72876 339561 73196 346325
rect 72876 339325 72918 339561
rect 73154 339325 73196 339561
rect 72876 332561 73196 339325
rect 72876 332325 72918 332561
rect 73154 332325 73196 332561
rect 72876 325561 73196 332325
rect 72876 325325 72918 325561
rect 73154 325325 73196 325561
rect 72876 318561 73196 325325
rect 72876 318325 72918 318561
rect 73154 318325 73196 318561
rect 72876 311561 73196 318325
rect 72876 311325 72918 311561
rect 73154 311325 73196 311561
rect 72876 304561 73196 311325
rect 72876 304325 72918 304561
rect 73154 304325 73196 304561
rect 72876 297561 73196 304325
rect 72876 297325 72918 297561
rect 73154 297325 73196 297561
rect 72876 290561 73196 297325
rect 72876 290325 72918 290561
rect 73154 290325 73196 290561
rect 72876 283561 73196 290325
rect 72876 283325 72918 283561
rect 73154 283325 73196 283561
rect 72876 276561 73196 283325
rect 72876 276325 72918 276561
rect 73154 276325 73196 276561
rect 72876 269561 73196 276325
rect 72876 269325 72918 269561
rect 73154 269325 73196 269561
rect 72876 262561 73196 269325
rect 72876 262325 72918 262561
rect 73154 262325 73196 262561
rect 72876 255561 73196 262325
rect 72876 255325 72918 255561
rect 73154 255325 73196 255561
rect 72876 248561 73196 255325
rect 72876 248325 72918 248561
rect 73154 248325 73196 248561
rect 72876 241561 73196 248325
rect 72876 241325 72918 241561
rect 73154 241325 73196 241561
rect 72876 234561 73196 241325
rect 72876 234325 72918 234561
rect 73154 234325 73196 234561
rect 72876 227561 73196 234325
rect 72876 227325 72918 227561
rect 73154 227325 73196 227561
rect 72876 220561 73196 227325
rect 72876 220325 72918 220561
rect 73154 220325 73196 220561
rect 72876 213561 73196 220325
rect 72876 213325 72918 213561
rect 73154 213325 73196 213561
rect 72876 206561 73196 213325
rect 72876 206325 72918 206561
rect 73154 206325 73196 206561
rect 72876 199561 73196 206325
rect 72876 199325 72918 199561
rect 73154 199325 73196 199561
rect 72876 192561 73196 199325
rect 72876 192325 72918 192561
rect 73154 192325 73196 192561
rect 72876 185561 73196 192325
rect 72876 185325 72918 185561
rect 73154 185325 73196 185561
rect 72876 178561 73196 185325
rect 72876 178325 72918 178561
rect 73154 178325 73196 178561
rect 72876 171561 73196 178325
rect 72876 171325 72918 171561
rect 73154 171325 73196 171561
rect 72876 164561 73196 171325
rect 72876 164325 72918 164561
rect 73154 164325 73196 164561
rect 72876 157561 73196 164325
rect 72876 157325 72918 157561
rect 73154 157325 73196 157561
rect 72876 150561 73196 157325
rect 72876 150325 72918 150561
rect 73154 150325 73196 150561
rect 72876 143561 73196 150325
rect 72876 143325 72918 143561
rect 73154 143325 73196 143561
rect 72876 136561 73196 143325
rect 72876 136325 72918 136561
rect 73154 136325 73196 136561
rect 72876 129561 73196 136325
rect 72876 129325 72918 129561
rect 73154 129325 73196 129561
rect 72876 122561 73196 129325
rect 72876 122325 72918 122561
rect 73154 122325 73196 122561
rect 72876 115561 73196 122325
rect 72876 115325 72918 115561
rect 73154 115325 73196 115561
rect 72876 108561 73196 115325
rect 72876 108325 72918 108561
rect 73154 108325 73196 108561
rect 72876 101561 73196 108325
rect 72876 101325 72918 101561
rect 73154 101325 73196 101561
rect 72876 94561 73196 101325
rect 72876 94325 72918 94561
rect 73154 94325 73196 94561
rect 72876 87561 73196 94325
rect 72876 87325 72918 87561
rect 73154 87325 73196 87561
rect 72876 80561 73196 87325
rect 72876 80325 72918 80561
rect 73154 80325 73196 80561
rect 72876 73561 73196 80325
rect 72876 73325 72918 73561
rect 73154 73325 73196 73561
rect 72876 66561 73196 73325
rect 72876 66325 72918 66561
rect 73154 66325 73196 66561
rect 72876 59561 73196 66325
rect 72876 59325 72918 59561
rect 73154 59325 73196 59561
rect 72876 52561 73196 59325
rect 72876 52325 72918 52561
rect 73154 52325 73196 52561
rect 72876 45561 73196 52325
rect 72876 45325 72918 45561
rect 73154 45325 73196 45561
rect 72876 38561 73196 45325
rect 72876 38325 72918 38561
rect 73154 38325 73196 38561
rect 72876 31561 73196 38325
rect 72876 31325 72918 31561
rect 73154 31325 73196 31561
rect 72876 24561 73196 31325
rect 72876 24325 72918 24561
rect 73154 24325 73196 24561
rect 72876 17561 73196 24325
rect 72876 17325 72918 17561
rect 73154 17325 73196 17561
rect 72876 10561 73196 17325
rect 72876 10325 72918 10561
rect 73154 10325 73196 10561
rect 72876 3561 73196 10325
rect 72876 3325 72918 3561
rect 73154 3325 73196 3561
rect 72876 -1706 73196 3325
rect 72876 -1942 72918 -1706
rect 73154 -1942 73196 -1706
rect 72876 -2026 73196 -1942
rect 72876 -2262 72918 -2026
rect 73154 -2262 73196 -2026
rect 72876 -2294 73196 -2262
rect 78144 705238 78464 706230
rect 78144 705002 78186 705238
rect 78422 705002 78464 705238
rect 78144 704918 78464 705002
rect 78144 704682 78186 704918
rect 78422 704682 78464 704918
rect 78144 695494 78464 704682
rect 78144 695258 78186 695494
rect 78422 695258 78464 695494
rect 78144 688494 78464 695258
rect 78144 688258 78186 688494
rect 78422 688258 78464 688494
rect 78144 681494 78464 688258
rect 78144 681258 78186 681494
rect 78422 681258 78464 681494
rect 78144 674494 78464 681258
rect 78144 674258 78186 674494
rect 78422 674258 78464 674494
rect 78144 667494 78464 674258
rect 78144 667258 78186 667494
rect 78422 667258 78464 667494
rect 78144 660494 78464 667258
rect 78144 660258 78186 660494
rect 78422 660258 78464 660494
rect 78144 653494 78464 660258
rect 78144 653258 78186 653494
rect 78422 653258 78464 653494
rect 78144 646494 78464 653258
rect 78144 646258 78186 646494
rect 78422 646258 78464 646494
rect 78144 639494 78464 646258
rect 78144 639258 78186 639494
rect 78422 639258 78464 639494
rect 78144 632494 78464 639258
rect 78144 632258 78186 632494
rect 78422 632258 78464 632494
rect 78144 625494 78464 632258
rect 78144 625258 78186 625494
rect 78422 625258 78464 625494
rect 78144 618494 78464 625258
rect 78144 618258 78186 618494
rect 78422 618258 78464 618494
rect 78144 611494 78464 618258
rect 78144 611258 78186 611494
rect 78422 611258 78464 611494
rect 78144 604494 78464 611258
rect 78144 604258 78186 604494
rect 78422 604258 78464 604494
rect 78144 597494 78464 604258
rect 78144 597258 78186 597494
rect 78422 597258 78464 597494
rect 78144 590494 78464 597258
rect 78144 590258 78186 590494
rect 78422 590258 78464 590494
rect 78144 583494 78464 590258
rect 78144 583258 78186 583494
rect 78422 583258 78464 583494
rect 78144 576494 78464 583258
rect 78144 576258 78186 576494
rect 78422 576258 78464 576494
rect 78144 569494 78464 576258
rect 78144 569258 78186 569494
rect 78422 569258 78464 569494
rect 78144 562494 78464 569258
rect 78144 562258 78186 562494
rect 78422 562258 78464 562494
rect 78144 555494 78464 562258
rect 78144 555258 78186 555494
rect 78422 555258 78464 555494
rect 78144 548494 78464 555258
rect 78144 548258 78186 548494
rect 78422 548258 78464 548494
rect 78144 541494 78464 548258
rect 78144 541258 78186 541494
rect 78422 541258 78464 541494
rect 78144 534494 78464 541258
rect 78144 534258 78186 534494
rect 78422 534258 78464 534494
rect 78144 527494 78464 534258
rect 78144 527258 78186 527494
rect 78422 527258 78464 527494
rect 78144 520494 78464 527258
rect 78144 520258 78186 520494
rect 78422 520258 78464 520494
rect 78144 513494 78464 520258
rect 78144 513258 78186 513494
rect 78422 513258 78464 513494
rect 78144 506494 78464 513258
rect 78144 506258 78186 506494
rect 78422 506258 78464 506494
rect 78144 499494 78464 506258
rect 78144 499258 78186 499494
rect 78422 499258 78464 499494
rect 78144 492494 78464 499258
rect 78144 492258 78186 492494
rect 78422 492258 78464 492494
rect 78144 485494 78464 492258
rect 78144 485258 78186 485494
rect 78422 485258 78464 485494
rect 78144 478494 78464 485258
rect 78144 478258 78186 478494
rect 78422 478258 78464 478494
rect 78144 471494 78464 478258
rect 78144 471258 78186 471494
rect 78422 471258 78464 471494
rect 78144 464494 78464 471258
rect 78144 464258 78186 464494
rect 78422 464258 78464 464494
rect 78144 457494 78464 464258
rect 78144 457258 78186 457494
rect 78422 457258 78464 457494
rect 78144 450494 78464 457258
rect 78144 450258 78186 450494
rect 78422 450258 78464 450494
rect 78144 443494 78464 450258
rect 78144 443258 78186 443494
rect 78422 443258 78464 443494
rect 78144 436494 78464 443258
rect 78144 436258 78186 436494
rect 78422 436258 78464 436494
rect 78144 429494 78464 436258
rect 78144 429258 78186 429494
rect 78422 429258 78464 429494
rect 78144 422494 78464 429258
rect 78144 422258 78186 422494
rect 78422 422258 78464 422494
rect 78144 415494 78464 422258
rect 78144 415258 78186 415494
rect 78422 415258 78464 415494
rect 78144 408494 78464 415258
rect 78144 408258 78186 408494
rect 78422 408258 78464 408494
rect 78144 401494 78464 408258
rect 78144 401258 78186 401494
rect 78422 401258 78464 401494
rect 78144 394494 78464 401258
rect 78144 394258 78186 394494
rect 78422 394258 78464 394494
rect 78144 387494 78464 394258
rect 78144 387258 78186 387494
rect 78422 387258 78464 387494
rect 78144 380494 78464 387258
rect 78144 380258 78186 380494
rect 78422 380258 78464 380494
rect 78144 373494 78464 380258
rect 78144 373258 78186 373494
rect 78422 373258 78464 373494
rect 78144 366494 78464 373258
rect 78144 366258 78186 366494
rect 78422 366258 78464 366494
rect 78144 359494 78464 366258
rect 78144 359258 78186 359494
rect 78422 359258 78464 359494
rect 78144 352494 78464 359258
rect 78144 352258 78186 352494
rect 78422 352258 78464 352494
rect 78144 345494 78464 352258
rect 78144 345258 78186 345494
rect 78422 345258 78464 345494
rect 78144 338494 78464 345258
rect 78144 338258 78186 338494
rect 78422 338258 78464 338494
rect 78144 331494 78464 338258
rect 78144 331258 78186 331494
rect 78422 331258 78464 331494
rect 78144 324494 78464 331258
rect 78144 324258 78186 324494
rect 78422 324258 78464 324494
rect 78144 317494 78464 324258
rect 78144 317258 78186 317494
rect 78422 317258 78464 317494
rect 78144 310494 78464 317258
rect 78144 310258 78186 310494
rect 78422 310258 78464 310494
rect 78144 303494 78464 310258
rect 78144 303258 78186 303494
rect 78422 303258 78464 303494
rect 78144 296494 78464 303258
rect 78144 296258 78186 296494
rect 78422 296258 78464 296494
rect 78144 289494 78464 296258
rect 78144 289258 78186 289494
rect 78422 289258 78464 289494
rect 78144 282494 78464 289258
rect 78144 282258 78186 282494
rect 78422 282258 78464 282494
rect 78144 275494 78464 282258
rect 78144 275258 78186 275494
rect 78422 275258 78464 275494
rect 78144 268494 78464 275258
rect 78144 268258 78186 268494
rect 78422 268258 78464 268494
rect 78144 261494 78464 268258
rect 78144 261258 78186 261494
rect 78422 261258 78464 261494
rect 78144 254494 78464 261258
rect 78144 254258 78186 254494
rect 78422 254258 78464 254494
rect 78144 247494 78464 254258
rect 78144 247258 78186 247494
rect 78422 247258 78464 247494
rect 78144 240494 78464 247258
rect 78144 240258 78186 240494
rect 78422 240258 78464 240494
rect 78144 233494 78464 240258
rect 78144 233258 78186 233494
rect 78422 233258 78464 233494
rect 78144 226494 78464 233258
rect 78144 226258 78186 226494
rect 78422 226258 78464 226494
rect 78144 219494 78464 226258
rect 78144 219258 78186 219494
rect 78422 219258 78464 219494
rect 78144 212494 78464 219258
rect 78144 212258 78186 212494
rect 78422 212258 78464 212494
rect 78144 205494 78464 212258
rect 78144 205258 78186 205494
rect 78422 205258 78464 205494
rect 78144 198494 78464 205258
rect 78144 198258 78186 198494
rect 78422 198258 78464 198494
rect 78144 191494 78464 198258
rect 78144 191258 78186 191494
rect 78422 191258 78464 191494
rect 78144 184494 78464 191258
rect 78144 184258 78186 184494
rect 78422 184258 78464 184494
rect 78144 177494 78464 184258
rect 78144 177258 78186 177494
rect 78422 177258 78464 177494
rect 78144 170494 78464 177258
rect 78144 170258 78186 170494
rect 78422 170258 78464 170494
rect 78144 163494 78464 170258
rect 78144 163258 78186 163494
rect 78422 163258 78464 163494
rect 78144 156494 78464 163258
rect 78144 156258 78186 156494
rect 78422 156258 78464 156494
rect 78144 149494 78464 156258
rect 78144 149258 78186 149494
rect 78422 149258 78464 149494
rect 78144 142494 78464 149258
rect 78144 142258 78186 142494
rect 78422 142258 78464 142494
rect 78144 135494 78464 142258
rect 78144 135258 78186 135494
rect 78422 135258 78464 135494
rect 78144 128494 78464 135258
rect 78144 128258 78186 128494
rect 78422 128258 78464 128494
rect 78144 121494 78464 128258
rect 78144 121258 78186 121494
rect 78422 121258 78464 121494
rect 78144 114494 78464 121258
rect 78144 114258 78186 114494
rect 78422 114258 78464 114494
rect 78144 107494 78464 114258
rect 78144 107258 78186 107494
rect 78422 107258 78464 107494
rect 78144 100494 78464 107258
rect 78144 100258 78186 100494
rect 78422 100258 78464 100494
rect 78144 93494 78464 100258
rect 78144 93258 78186 93494
rect 78422 93258 78464 93494
rect 78144 86494 78464 93258
rect 78144 86258 78186 86494
rect 78422 86258 78464 86494
rect 78144 79494 78464 86258
rect 78144 79258 78186 79494
rect 78422 79258 78464 79494
rect 78144 72494 78464 79258
rect 78144 72258 78186 72494
rect 78422 72258 78464 72494
rect 78144 65494 78464 72258
rect 78144 65258 78186 65494
rect 78422 65258 78464 65494
rect 78144 58494 78464 65258
rect 78144 58258 78186 58494
rect 78422 58258 78464 58494
rect 78144 51494 78464 58258
rect 78144 51258 78186 51494
rect 78422 51258 78464 51494
rect 78144 44494 78464 51258
rect 78144 44258 78186 44494
rect 78422 44258 78464 44494
rect 78144 37494 78464 44258
rect 78144 37258 78186 37494
rect 78422 37258 78464 37494
rect 78144 30494 78464 37258
rect 78144 30258 78186 30494
rect 78422 30258 78464 30494
rect 78144 23494 78464 30258
rect 78144 23258 78186 23494
rect 78422 23258 78464 23494
rect 78144 16494 78464 23258
rect 78144 16258 78186 16494
rect 78422 16258 78464 16494
rect 78144 9494 78464 16258
rect 78144 9258 78186 9494
rect 78422 9258 78464 9494
rect 78144 2494 78464 9258
rect 78144 2258 78186 2494
rect 78422 2258 78464 2494
rect 78144 -746 78464 2258
rect 78144 -982 78186 -746
rect 78422 -982 78464 -746
rect 78144 -1066 78464 -982
rect 78144 -1302 78186 -1066
rect 78422 -1302 78464 -1066
rect 78144 -2294 78464 -1302
rect 79876 706198 80196 706230
rect 79876 705962 79918 706198
rect 80154 705962 80196 706198
rect 79876 705878 80196 705962
rect 79876 705642 79918 705878
rect 80154 705642 80196 705878
rect 79876 696561 80196 705642
rect 79876 696325 79918 696561
rect 80154 696325 80196 696561
rect 79876 689561 80196 696325
rect 79876 689325 79918 689561
rect 80154 689325 80196 689561
rect 79876 682561 80196 689325
rect 79876 682325 79918 682561
rect 80154 682325 80196 682561
rect 79876 675561 80196 682325
rect 79876 675325 79918 675561
rect 80154 675325 80196 675561
rect 79876 668561 80196 675325
rect 79876 668325 79918 668561
rect 80154 668325 80196 668561
rect 79876 661561 80196 668325
rect 79876 661325 79918 661561
rect 80154 661325 80196 661561
rect 79876 654561 80196 661325
rect 79876 654325 79918 654561
rect 80154 654325 80196 654561
rect 79876 647561 80196 654325
rect 79876 647325 79918 647561
rect 80154 647325 80196 647561
rect 79876 640561 80196 647325
rect 79876 640325 79918 640561
rect 80154 640325 80196 640561
rect 79876 633561 80196 640325
rect 79876 633325 79918 633561
rect 80154 633325 80196 633561
rect 79876 626561 80196 633325
rect 79876 626325 79918 626561
rect 80154 626325 80196 626561
rect 79876 619561 80196 626325
rect 79876 619325 79918 619561
rect 80154 619325 80196 619561
rect 79876 612561 80196 619325
rect 79876 612325 79918 612561
rect 80154 612325 80196 612561
rect 79876 605561 80196 612325
rect 79876 605325 79918 605561
rect 80154 605325 80196 605561
rect 79876 598561 80196 605325
rect 79876 598325 79918 598561
rect 80154 598325 80196 598561
rect 79876 591561 80196 598325
rect 79876 591325 79918 591561
rect 80154 591325 80196 591561
rect 79876 584561 80196 591325
rect 79876 584325 79918 584561
rect 80154 584325 80196 584561
rect 79876 577561 80196 584325
rect 79876 577325 79918 577561
rect 80154 577325 80196 577561
rect 79876 570561 80196 577325
rect 79876 570325 79918 570561
rect 80154 570325 80196 570561
rect 79876 563561 80196 570325
rect 79876 563325 79918 563561
rect 80154 563325 80196 563561
rect 79876 556561 80196 563325
rect 79876 556325 79918 556561
rect 80154 556325 80196 556561
rect 79876 549561 80196 556325
rect 79876 549325 79918 549561
rect 80154 549325 80196 549561
rect 79876 542561 80196 549325
rect 79876 542325 79918 542561
rect 80154 542325 80196 542561
rect 79876 535561 80196 542325
rect 79876 535325 79918 535561
rect 80154 535325 80196 535561
rect 79876 528561 80196 535325
rect 79876 528325 79918 528561
rect 80154 528325 80196 528561
rect 79876 521561 80196 528325
rect 79876 521325 79918 521561
rect 80154 521325 80196 521561
rect 79876 514561 80196 521325
rect 79876 514325 79918 514561
rect 80154 514325 80196 514561
rect 79876 507561 80196 514325
rect 79876 507325 79918 507561
rect 80154 507325 80196 507561
rect 79876 500561 80196 507325
rect 79876 500325 79918 500561
rect 80154 500325 80196 500561
rect 79876 493561 80196 500325
rect 79876 493325 79918 493561
rect 80154 493325 80196 493561
rect 79876 486561 80196 493325
rect 79876 486325 79918 486561
rect 80154 486325 80196 486561
rect 79876 479561 80196 486325
rect 79876 479325 79918 479561
rect 80154 479325 80196 479561
rect 79876 472561 80196 479325
rect 79876 472325 79918 472561
rect 80154 472325 80196 472561
rect 79876 465561 80196 472325
rect 79876 465325 79918 465561
rect 80154 465325 80196 465561
rect 79876 458561 80196 465325
rect 79876 458325 79918 458561
rect 80154 458325 80196 458561
rect 79876 451561 80196 458325
rect 79876 451325 79918 451561
rect 80154 451325 80196 451561
rect 79876 444561 80196 451325
rect 79876 444325 79918 444561
rect 80154 444325 80196 444561
rect 79876 437561 80196 444325
rect 79876 437325 79918 437561
rect 80154 437325 80196 437561
rect 79876 430561 80196 437325
rect 79876 430325 79918 430561
rect 80154 430325 80196 430561
rect 79876 423561 80196 430325
rect 79876 423325 79918 423561
rect 80154 423325 80196 423561
rect 79876 416561 80196 423325
rect 79876 416325 79918 416561
rect 80154 416325 80196 416561
rect 79876 409561 80196 416325
rect 79876 409325 79918 409561
rect 80154 409325 80196 409561
rect 79876 402561 80196 409325
rect 79876 402325 79918 402561
rect 80154 402325 80196 402561
rect 79876 395561 80196 402325
rect 79876 395325 79918 395561
rect 80154 395325 80196 395561
rect 79876 388561 80196 395325
rect 79876 388325 79918 388561
rect 80154 388325 80196 388561
rect 79876 381561 80196 388325
rect 79876 381325 79918 381561
rect 80154 381325 80196 381561
rect 79876 374561 80196 381325
rect 79876 374325 79918 374561
rect 80154 374325 80196 374561
rect 79876 367561 80196 374325
rect 79876 367325 79918 367561
rect 80154 367325 80196 367561
rect 79876 360561 80196 367325
rect 79876 360325 79918 360561
rect 80154 360325 80196 360561
rect 79876 353561 80196 360325
rect 79876 353325 79918 353561
rect 80154 353325 80196 353561
rect 79876 346561 80196 353325
rect 79876 346325 79918 346561
rect 80154 346325 80196 346561
rect 79876 339561 80196 346325
rect 79876 339325 79918 339561
rect 80154 339325 80196 339561
rect 79876 332561 80196 339325
rect 79876 332325 79918 332561
rect 80154 332325 80196 332561
rect 79876 325561 80196 332325
rect 79876 325325 79918 325561
rect 80154 325325 80196 325561
rect 79876 318561 80196 325325
rect 79876 318325 79918 318561
rect 80154 318325 80196 318561
rect 79876 311561 80196 318325
rect 79876 311325 79918 311561
rect 80154 311325 80196 311561
rect 79876 304561 80196 311325
rect 79876 304325 79918 304561
rect 80154 304325 80196 304561
rect 79876 297561 80196 304325
rect 79876 297325 79918 297561
rect 80154 297325 80196 297561
rect 79876 290561 80196 297325
rect 79876 290325 79918 290561
rect 80154 290325 80196 290561
rect 79876 283561 80196 290325
rect 79876 283325 79918 283561
rect 80154 283325 80196 283561
rect 79876 276561 80196 283325
rect 79876 276325 79918 276561
rect 80154 276325 80196 276561
rect 79876 269561 80196 276325
rect 79876 269325 79918 269561
rect 80154 269325 80196 269561
rect 79876 262561 80196 269325
rect 79876 262325 79918 262561
rect 80154 262325 80196 262561
rect 79876 255561 80196 262325
rect 79876 255325 79918 255561
rect 80154 255325 80196 255561
rect 79876 248561 80196 255325
rect 79876 248325 79918 248561
rect 80154 248325 80196 248561
rect 79876 241561 80196 248325
rect 79876 241325 79918 241561
rect 80154 241325 80196 241561
rect 79876 234561 80196 241325
rect 79876 234325 79918 234561
rect 80154 234325 80196 234561
rect 79876 227561 80196 234325
rect 79876 227325 79918 227561
rect 80154 227325 80196 227561
rect 79876 220561 80196 227325
rect 79876 220325 79918 220561
rect 80154 220325 80196 220561
rect 79876 213561 80196 220325
rect 79876 213325 79918 213561
rect 80154 213325 80196 213561
rect 79876 206561 80196 213325
rect 79876 206325 79918 206561
rect 80154 206325 80196 206561
rect 79876 199561 80196 206325
rect 79876 199325 79918 199561
rect 80154 199325 80196 199561
rect 79876 192561 80196 199325
rect 79876 192325 79918 192561
rect 80154 192325 80196 192561
rect 79876 185561 80196 192325
rect 79876 185325 79918 185561
rect 80154 185325 80196 185561
rect 79876 178561 80196 185325
rect 79876 178325 79918 178561
rect 80154 178325 80196 178561
rect 79876 171561 80196 178325
rect 79876 171325 79918 171561
rect 80154 171325 80196 171561
rect 79876 164561 80196 171325
rect 79876 164325 79918 164561
rect 80154 164325 80196 164561
rect 79876 157561 80196 164325
rect 79876 157325 79918 157561
rect 80154 157325 80196 157561
rect 79876 150561 80196 157325
rect 79876 150325 79918 150561
rect 80154 150325 80196 150561
rect 79876 143561 80196 150325
rect 79876 143325 79918 143561
rect 80154 143325 80196 143561
rect 79876 136561 80196 143325
rect 79876 136325 79918 136561
rect 80154 136325 80196 136561
rect 79876 129561 80196 136325
rect 79876 129325 79918 129561
rect 80154 129325 80196 129561
rect 79876 122561 80196 129325
rect 79876 122325 79918 122561
rect 80154 122325 80196 122561
rect 79876 115561 80196 122325
rect 79876 115325 79918 115561
rect 80154 115325 80196 115561
rect 79876 108561 80196 115325
rect 79876 108325 79918 108561
rect 80154 108325 80196 108561
rect 79876 101561 80196 108325
rect 79876 101325 79918 101561
rect 80154 101325 80196 101561
rect 79876 94561 80196 101325
rect 79876 94325 79918 94561
rect 80154 94325 80196 94561
rect 79876 87561 80196 94325
rect 79876 87325 79918 87561
rect 80154 87325 80196 87561
rect 79876 80561 80196 87325
rect 79876 80325 79918 80561
rect 80154 80325 80196 80561
rect 79876 73561 80196 80325
rect 79876 73325 79918 73561
rect 80154 73325 80196 73561
rect 79876 66561 80196 73325
rect 79876 66325 79918 66561
rect 80154 66325 80196 66561
rect 79876 59561 80196 66325
rect 79876 59325 79918 59561
rect 80154 59325 80196 59561
rect 79876 52561 80196 59325
rect 79876 52325 79918 52561
rect 80154 52325 80196 52561
rect 79876 45561 80196 52325
rect 79876 45325 79918 45561
rect 80154 45325 80196 45561
rect 79876 38561 80196 45325
rect 79876 38325 79918 38561
rect 80154 38325 80196 38561
rect 79876 31561 80196 38325
rect 79876 31325 79918 31561
rect 80154 31325 80196 31561
rect 79876 24561 80196 31325
rect 79876 24325 79918 24561
rect 80154 24325 80196 24561
rect 79876 17561 80196 24325
rect 79876 17325 79918 17561
rect 80154 17325 80196 17561
rect 79876 10561 80196 17325
rect 79876 10325 79918 10561
rect 80154 10325 80196 10561
rect 79876 3561 80196 10325
rect 79876 3325 79918 3561
rect 80154 3325 80196 3561
rect 79876 -1706 80196 3325
rect 79876 -1942 79918 -1706
rect 80154 -1942 80196 -1706
rect 79876 -2026 80196 -1942
rect 79876 -2262 79918 -2026
rect 80154 -2262 80196 -2026
rect 79876 -2294 80196 -2262
rect 85144 705238 85464 706230
rect 85144 705002 85186 705238
rect 85422 705002 85464 705238
rect 85144 704918 85464 705002
rect 85144 704682 85186 704918
rect 85422 704682 85464 704918
rect 85144 695494 85464 704682
rect 85144 695258 85186 695494
rect 85422 695258 85464 695494
rect 85144 688494 85464 695258
rect 85144 688258 85186 688494
rect 85422 688258 85464 688494
rect 85144 681494 85464 688258
rect 85144 681258 85186 681494
rect 85422 681258 85464 681494
rect 85144 674494 85464 681258
rect 85144 674258 85186 674494
rect 85422 674258 85464 674494
rect 85144 667494 85464 674258
rect 85144 667258 85186 667494
rect 85422 667258 85464 667494
rect 85144 660494 85464 667258
rect 85144 660258 85186 660494
rect 85422 660258 85464 660494
rect 85144 653494 85464 660258
rect 85144 653258 85186 653494
rect 85422 653258 85464 653494
rect 85144 646494 85464 653258
rect 85144 646258 85186 646494
rect 85422 646258 85464 646494
rect 85144 639494 85464 646258
rect 85144 639258 85186 639494
rect 85422 639258 85464 639494
rect 85144 632494 85464 639258
rect 85144 632258 85186 632494
rect 85422 632258 85464 632494
rect 85144 625494 85464 632258
rect 85144 625258 85186 625494
rect 85422 625258 85464 625494
rect 85144 618494 85464 625258
rect 85144 618258 85186 618494
rect 85422 618258 85464 618494
rect 85144 611494 85464 618258
rect 85144 611258 85186 611494
rect 85422 611258 85464 611494
rect 85144 604494 85464 611258
rect 85144 604258 85186 604494
rect 85422 604258 85464 604494
rect 85144 597494 85464 604258
rect 85144 597258 85186 597494
rect 85422 597258 85464 597494
rect 85144 590494 85464 597258
rect 85144 590258 85186 590494
rect 85422 590258 85464 590494
rect 85144 583494 85464 590258
rect 85144 583258 85186 583494
rect 85422 583258 85464 583494
rect 85144 576494 85464 583258
rect 85144 576258 85186 576494
rect 85422 576258 85464 576494
rect 85144 569494 85464 576258
rect 85144 569258 85186 569494
rect 85422 569258 85464 569494
rect 85144 562494 85464 569258
rect 85144 562258 85186 562494
rect 85422 562258 85464 562494
rect 85144 555494 85464 562258
rect 85144 555258 85186 555494
rect 85422 555258 85464 555494
rect 85144 548494 85464 555258
rect 85144 548258 85186 548494
rect 85422 548258 85464 548494
rect 85144 541494 85464 548258
rect 85144 541258 85186 541494
rect 85422 541258 85464 541494
rect 85144 534494 85464 541258
rect 85144 534258 85186 534494
rect 85422 534258 85464 534494
rect 85144 527494 85464 534258
rect 85144 527258 85186 527494
rect 85422 527258 85464 527494
rect 85144 520494 85464 527258
rect 85144 520258 85186 520494
rect 85422 520258 85464 520494
rect 85144 513494 85464 520258
rect 85144 513258 85186 513494
rect 85422 513258 85464 513494
rect 85144 506494 85464 513258
rect 85144 506258 85186 506494
rect 85422 506258 85464 506494
rect 85144 499494 85464 506258
rect 85144 499258 85186 499494
rect 85422 499258 85464 499494
rect 85144 492494 85464 499258
rect 85144 492258 85186 492494
rect 85422 492258 85464 492494
rect 85144 485494 85464 492258
rect 85144 485258 85186 485494
rect 85422 485258 85464 485494
rect 85144 478494 85464 485258
rect 85144 478258 85186 478494
rect 85422 478258 85464 478494
rect 85144 471494 85464 478258
rect 85144 471258 85186 471494
rect 85422 471258 85464 471494
rect 85144 464494 85464 471258
rect 85144 464258 85186 464494
rect 85422 464258 85464 464494
rect 85144 457494 85464 464258
rect 85144 457258 85186 457494
rect 85422 457258 85464 457494
rect 85144 450494 85464 457258
rect 85144 450258 85186 450494
rect 85422 450258 85464 450494
rect 85144 443494 85464 450258
rect 85144 443258 85186 443494
rect 85422 443258 85464 443494
rect 85144 436494 85464 443258
rect 85144 436258 85186 436494
rect 85422 436258 85464 436494
rect 85144 429494 85464 436258
rect 85144 429258 85186 429494
rect 85422 429258 85464 429494
rect 85144 422494 85464 429258
rect 85144 422258 85186 422494
rect 85422 422258 85464 422494
rect 85144 415494 85464 422258
rect 85144 415258 85186 415494
rect 85422 415258 85464 415494
rect 85144 408494 85464 415258
rect 85144 408258 85186 408494
rect 85422 408258 85464 408494
rect 85144 401494 85464 408258
rect 85144 401258 85186 401494
rect 85422 401258 85464 401494
rect 85144 394494 85464 401258
rect 85144 394258 85186 394494
rect 85422 394258 85464 394494
rect 85144 387494 85464 394258
rect 85144 387258 85186 387494
rect 85422 387258 85464 387494
rect 85144 380494 85464 387258
rect 85144 380258 85186 380494
rect 85422 380258 85464 380494
rect 85144 373494 85464 380258
rect 85144 373258 85186 373494
rect 85422 373258 85464 373494
rect 85144 366494 85464 373258
rect 85144 366258 85186 366494
rect 85422 366258 85464 366494
rect 85144 359494 85464 366258
rect 85144 359258 85186 359494
rect 85422 359258 85464 359494
rect 85144 352494 85464 359258
rect 85144 352258 85186 352494
rect 85422 352258 85464 352494
rect 85144 345494 85464 352258
rect 85144 345258 85186 345494
rect 85422 345258 85464 345494
rect 85144 338494 85464 345258
rect 85144 338258 85186 338494
rect 85422 338258 85464 338494
rect 85144 331494 85464 338258
rect 85144 331258 85186 331494
rect 85422 331258 85464 331494
rect 85144 324494 85464 331258
rect 85144 324258 85186 324494
rect 85422 324258 85464 324494
rect 85144 317494 85464 324258
rect 85144 317258 85186 317494
rect 85422 317258 85464 317494
rect 85144 310494 85464 317258
rect 85144 310258 85186 310494
rect 85422 310258 85464 310494
rect 85144 303494 85464 310258
rect 85144 303258 85186 303494
rect 85422 303258 85464 303494
rect 85144 296494 85464 303258
rect 85144 296258 85186 296494
rect 85422 296258 85464 296494
rect 85144 289494 85464 296258
rect 85144 289258 85186 289494
rect 85422 289258 85464 289494
rect 85144 282494 85464 289258
rect 85144 282258 85186 282494
rect 85422 282258 85464 282494
rect 85144 275494 85464 282258
rect 85144 275258 85186 275494
rect 85422 275258 85464 275494
rect 85144 268494 85464 275258
rect 85144 268258 85186 268494
rect 85422 268258 85464 268494
rect 85144 261494 85464 268258
rect 85144 261258 85186 261494
rect 85422 261258 85464 261494
rect 85144 254494 85464 261258
rect 85144 254258 85186 254494
rect 85422 254258 85464 254494
rect 85144 247494 85464 254258
rect 85144 247258 85186 247494
rect 85422 247258 85464 247494
rect 85144 240494 85464 247258
rect 85144 240258 85186 240494
rect 85422 240258 85464 240494
rect 85144 233494 85464 240258
rect 85144 233258 85186 233494
rect 85422 233258 85464 233494
rect 85144 226494 85464 233258
rect 85144 226258 85186 226494
rect 85422 226258 85464 226494
rect 85144 219494 85464 226258
rect 85144 219258 85186 219494
rect 85422 219258 85464 219494
rect 85144 212494 85464 219258
rect 85144 212258 85186 212494
rect 85422 212258 85464 212494
rect 85144 205494 85464 212258
rect 85144 205258 85186 205494
rect 85422 205258 85464 205494
rect 85144 198494 85464 205258
rect 85144 198258 85186 198494
rect 85422 198258 85464 198494
rect 85144 191494 85464 198258
rect 85144 191258 85186 191494
rect 85422 191258 85464 191494
rect 85144 184494 85464 191258
rect 85144 184258 85186 184494
rect 85422 184258 85464 184494
rect 85144 177494 85464 184258
rect 85144 177258 85186 177494
rect 85422 177258 85464 177494
rect 85144 170494 85464 177258
rect 85144 170258 85186 170494
rect 85422 170258 85464 170494
rect 85144 163494 85464 170258
rect 85144 163258 85186 163494
rect 85422 163258 85464 163494
rect 85144 156494 85464 163258
rect 85144 156258 85186 156494
rect 85422 156258 85464 156494
rect 85144 149494 85464 156258
rect 85144 149258 85186 149494
rect 85422 149258 85464 149494
rect 85144 142494 85464 149258
rect 85144 142258 85186 142494
rect 85422 142258 85464 142494
rect 85144 135494 85464 142258
rect 85144 135258 85186 135494
rect 85422 135258 85464 135494
rect 85144 128494 85464 135258
rect 85144 128258 85186 128494
rect 85422 128258 85464 128494
rect 85144 121494 85464 128258
rect 85144 121258 85186 121494
rect 85422 121258 85464 121494
rect 85144 114494 85464 121258
rect 85144 114258 85186 114494
rect 85422 114258 85464 114494
rect 85144 107494 85464 114258
rect 85144 107258 85186 107494
rect 85422 107258 85464 107494
rect 85144 100494 85464 107258
rect 85144 100258 85186 100494
rect 85422 100258 85464 100494
rect 85144 93494 85464 100258
rect 85144 93258 85186 93494
rect 85422 93258 85464 93494
rect 85144 86494 85464 93258
rect 85144 86258 85186 86494
rect 85422 86258 85464 86494
rect 85144 79494 85464 86258
rect 85144 79258 85186 79494
rect 85422 79258 85464 79494
rect 85144 72494 85464 79258
rect 85144 72258 85186 72494
rect 85422 72258 85464 72494
rect 85144 65494 85464 72258
rect 85144 65258 85186 65494
rect 85422 65258 85464 65494
rect 85144 58494 85464 65258
rect 85144 58258 85186 58494
rect 85422 58258 85464 58494
rect 85144 51494 85464 58258
rect 85144 51258 85186 51494
rect 85422 51258 85464 51494
rect 85144 44494 85464 51258
rect 85144 44258 85186 44494
rect 85422 44258 85464 44494
rect 85144 37494 85464 44258
rect 85144 37258 85186 37494
rect 85422 37258 85464 37494
rect 85144 30494 85464 37258
rect 85144 30258 85186 30494
rect 85422 30258 85464 30494
rect 85144 23494 85464 30258
rect 85144 23258 85186 23494
rect 85422 23258 85464 23494
rect 85144 16494 85464 23258
rect 85144 16258 85186 16494
rect 85422 16258 85464 16494
rect 85144 9494 85464 16258
rect 85144 9258 85186 9494
rect 85422 9258 85464 9494
rect 85144 2494 85464 9258
rect 85144 2258 85186 2494
rect 85422 2258 85464 2494
rect 85144 -746 85464 2258
rect 85144 -982 85186 -746
rect 85422 -982 85464 -746
rect 85144 -1066 85464 -982
rect 85144 -1302 85186 -1066
rect 85422 -1302 85464 -1066
rect 85144 -2294 85464 -1302
rect 86876 706198 87196 706230
rect 86876 705962 86918 706198
rect 87154 705962 87196 706198
rect 86876 705878 87196 705962
rect 86876 705642 86918 705878
rect 87154 705642 87196 705878
rect 86876 696561 87196 705642
rect 86876 696325 86918 696561
rect 87154 696325 87196 696561
rect 86876 689561 87196 696325
rect 86876 689325 86918 689561
rect 87154 689325 87196 689561
rect 86876 682561 87196 689325
rect 86876 682325 86918 682561
rect 87154 682325 87196 682561
rect 86876 675561 87196 682325
rect 86876 675325 86918 675561
rect 87154 675325 87196 675561
rect 86876 668561 87196 675325
rect 86876 668325 86918 668561
rect 87154 668325 87196 668561
rect 86876 661561 87196 668325
rect 86876 661325 86918 661561
rect 87154 661325 87196 661561
rect 86876 654561 87196 661325
rect 86876 654325 86918 654561
rect 87154 654325 87196 654561
rect 86876 647561 87196 654325
rect 86876 647325 86918 647561
rect 87154 647325 87196 647561
rect 86876 640561 87196 647325
rect 86876 640325 86918 640561
rect 87154 640325 87196 640561
rect 86876 633561 87196 640325
rect 86876 633325 86918 633561
rect 87154 633325 87196 633561
rect 86876 626561 87196 633325
rect 86876 626325 86918 626561
rect 87154 626325 87196 626561
rect 86876 619561 87196 626325
rect 86876 619325 86918 619561
rect 87154 619325 87196 619561
rect 86876 612561 87196 619325
rect 86876 612325 86918 612561
rect 87154 612325 87196 612561
rect 86876 605561 87196 612325
rect 86876 605325 86918 605561
rect 87154 605325 87196 605561
rect 86876 598561 87196 605325
rect 86876 598325 86918 598561
rect 87154 598325 87196 598561
rect 86876 591561 87196 598325
rect 86876 591325 86918 591561
rect 87154 591325 87196 591561
rect 86876 584561 87196 591325
rect 86876 584325 86918 584561
rect 87154 584325 87196 584561
rect 86876 577561 87196 584325
rect 86876 577325 86918 577561
rect 87154 577325 87196 577561
rect 86876 570561 87196 577325
rect 86876 570325 86918 570561
rect 87154 570325 87196 570561
rect 86876 563561 87196 570325
rect 86876 563325 86918 563561
rect 87154 563325 87196 563561
rect 86876 556561 87196 563325
rect 86876 556325 86918 556561
rect 87154 556325 87196 556561
rect 86876 549561 87196 556325
rect 86876 549325 86918 549561
rect 87154 549325 87196 549561
rect 86876 542561 87196 549325
rect 86876 542325 86918 542561
rect 87154 542325 87196 542561
rect 86876 535561 87196 542325
rect 86876 535325 86918 535561
rect 87154 535325 87196 535561
rect 86876 528561 87196 535325
rect 86876 528325 86918 528561
rect 87154 528325 87196 528561
rect 86876 521561 87196 528325
rect 86876 521325 86918 521561
rect 87154 521325 87196 521561
rect 86876 514561 87196 521325
rect 86876 514325 86918 514561
rect 87154 514325 87196 514561
rect 86876 507561 87196 514325
rect 86876 507325 86918 507561
rect 87154 507325 87196 507561
rect 86876 500561 87196 507325
rect 86876 500325 86918 500561
rect 87154 500325 87196 500561
rect 86876 493561 87196 500325
rect 86876 493325 86918 493561
rect 87154 493325 87196 493561
rect 86876 486561 87196 493325
rect 86876 486325 86918 486561
rect 87154 486325 87196 486561
rect 86876 479561 87196 486325
rect 86876 479325 86918 479561
rect 87154 479325 87196 479561
rect 86876 472561 87196 479325
rect 86876 472325 86918 472561
rect 87154 472325 87196 472561
rect 86876 465561 87196 472325
rect 86876 465325 86918 465561
rect 87154 465325 87196 465561
rect 86876 458561 87196 465325
rect 86876 458325 86918 458561
rect 87154 458325 87196 458561
rect 86876 451561 87196 458325
rect 86876 451325 86918 451561
rect 87154 451325 87196 451561
rect 86876 444561 87196 451325
rect 86876 444325 86918 444561
rect 87154 444325 87196 444561
rect 86876 437561 87196 444325
rect 86876 437325 86918 437561
rect 87154 437325 87196 437561
rect 86876 430561 87196 437325
rect 86876 430325 86918 430561
rect 87154 430325 87196 430561
rect 86876 423561 87196 430325
rect 86876 423325 86918 423561
rect 87154 423325 87196 423561
rect 86876 416561 87196 423325
rect 86876 416325 86918 416561
rect 87154 416325 87196 416561
rect 86876 409561 87196 416325
rect 86876 409325 86918 409561
rect 87154 409325 87196 409561
rect 86876 402561 87196 409325
rect 86876 402325 86918 402561
rect 87154 402325 87196 402561
rect 86876 395561 87196 402325
rect 86876 395325 86918 395561
rect 87154 395325 87196 395561
rect 86876 388561 87196 395325
rect 86876 388325 86918 388561
rect 87154 388325 87196 388561
rect 86876 381561 87196 388325
rect 86876 381325 86918 381561
rect 87154 381325 87196 381561
rect 86876 374561 87196 381325
rect 86876 374325 86918 374561
rect 87154 374325 87196 374561
rect 86876 367561 87196 374325
rect 86876 367325 86918 367561
rect 87154 367325 87196 367561
rect 86876 360561 87196 367325
rect 86876 360325 86918 360561
rect 87154 360325 87196 360561
rect 86876 353561 87196 360325
rect 86876 353325 86918 353561
rect 87154 353325 87196 353561
rect 86876 346561 87196 353325
rect 86876 346325 86918 346561
rect 87154 346325 87196 346561
rect 86876 339561 87196 346325
rect 86876 339325 86918 339561
rect 87154 339325 87196 339561
rect 86876 332561 87196 339325
rect 86876 332325 86918 332561
rect 87154 332325 87196 332561
rect 86876 325561 87196 332325
rect 86876 325325 86918 325561
rect 87154 325325 87196 325561
rect 86876 318561 87196 325325
rect 86876 318325 86918 318561
rect 87154 318325 87196 318561
rect 86876 311561 87196 318325
rect 86876 311325 86918 311561
rect 87154 311325 87196 311561
rect 86876 304561 87196 311325
rect 86876 304325 86918 304561
rect 87154 304325 87196 304561
rect 86876 297561 87196 304325
rect 86876 297325 86918 297561
rect 87154 297325 87196 297561
rect 86876 290561 87196 297325
rect 86876 290325 86918 290561
rect 87154 290325 87196 290561
rect 86876 283561 87196 290325
rect 86876 283325 86918 283561
rect 87154 283325 87196 283561
rect 86876 276561 87196 283325
rect 86876 276325 86918 276561
rect 87154 276325 87196 276561
rect 86876 269561 87196 276325
rect 86876 269325 86918 269561
rect 87154 269325 87196 269561
rect 86876 262561 87196 269325
rect 86876 262325 86918 262561
rect 87154 262325 87196 262561
rect 86876 255561 87196 262325
rect 86876 255325 86918 255561
rect 87154 255325 87196 255561
rect 86876 248561 87196 255325
rect 86876 248325 86918 248561
rect 87154 248325 87196 248561
rect 86876 241561 87196 248325
rect 86876 241325 86918 241561
rect 87154 241325 87196 241561
rect 86876 234561 87196 241325
rect 86876 234325 86918 234561
rect 87154 234325 87196 234561
rect 86876 227561 87196 234325
rect 86876 227325 86918 227561
rect 87154 227325 87196 227561
rect 86876 220561 87196 227325
rect 86876 220325 86918 220561
rect 87154 220325 87196 220561
rect 86876 213561 87196 220325
rect 86876 213325 86918 213561
rect 87154 213325 87196 213561
rect 86876 206561 87196 213325
rect 86876 206325 86918 206561
rect 87154 206325 87196 206561
rect 86876 199561 87196 206325
rect 86876 199325 86918 199561
rect 87154 199325 87196 199561
rect 86876 192561 87196 199325
rect 86876 192325 86918 192561
rect 87154 192325 87196 192561
rect 86876 185561 87196 192325
rect 86876 185325 86918 185561
rect 87154 185325 87196 185561
rect 86876 178561 87196 185325
rect 86876 178325 86918 178561
rect 87154 178325 87196 178561
rect 86876 171561 87196 178325
rect 86876 171325 86918 171561
rect 87154 171325 87196 171561
rect 86876 164561 87196 171325
rect 86876 164325 86918 164561
rect 87154 164325 87196 164561
rect 86876 157561 87196 164325
rect 86876 157325 86918 157561
rect 87154 157325 87196 157561
rect 86876 150561 87196 157325
rect 86876 150325 86918 150561
rect 87154 150325 87196 150561
rect 86876 143561 87196 150325
rect 86876 143325 86918 143561
rect 87154 143325 87196 143561
rect 86876 136561 87196 143325
rect 86876 136325 86918 136561
rect 87154 136325 87196 136561
rect 86876 129561 87196 136325
rect 86876 129325 86918 129561
rect 87154 129325 87196 129561
rect 86876 122561 87196 129325
rect 86876 122325 86918 122561
rect 87154 122325 87196 122561
rect 86876 115561 87196 122325
rect 86876 115325 86918 115561
rect 87154 115325 87196 115561
rect 86876 108561 87196 115325
rect 86876 108325 86918 108561
rect 87154 108325 87196 108561
rect 86876 101561 87196 108325
rect 86876 101325 86918 101561
rect 87154 101325 87196 101561
rect 86876 94561 87196 101325
rect 86876 94325 86918 94561
rect 87154 94325 87196 94561
rect 86876 87561 87196 94325
rect 86876 87325 86918 87561
rect 87154 87325 87196 87561
rect 86876 80561 87196 87325
rect 86876 80325 86918 80561
rect 87154 80325 87196 80561
rect 86876 73561 87196 80325
rect 86876 73325 86918 73561
rect 87154 73325 87196 73561
rect 86876 66561 87196 73325
rect 86876 66325 86918 66561
rect 87154 66325 87196 66561
rect 86876 59561 87196 66325
rect 86876 59325 86918 59561
rect 87154 59325 87196 59561
rect 86876 52561 87196 59325
rect 86876 52325 86918 52561
rect 87154 52325 87196 52561
rect 86876 45561 87196 52325
rect 86876 45325 86918 45561
rect 87154 45325 87196 45561
rect 86876 38561 87196 45325
rect 86876 38325 86918 38561
rect 87154 38325 87196 38561
rect 86876 31561 87196 38325
rect 86876 31325 86918 31561
rect 87154 31325 87196 31561
rect 86876 24561 87196 31325
rect 86876 24325 86918 24561
rect 87154 24325 87196 24561
rect 86876 17561 87196 24325
rect 86876 17325 86918 17561
rect 87154 17325 87196 17561
rect 86876 10561 87196 17325
rect 86876 10325 86918 10561
rect 87154 10325 87196 10561
rect 86876 3561 87196 10325
rect 86876 3325 86918 3561
rect 87154 3325 87196 3561
rect 86876 -1706 87196 3325
rect 86876 -1942 86918 -1706
rect 87154 -1942 87196 -1706
rect 86876 -2026 87196 -1942
rect 86876 -2262 86918 -2026
rect 87154 -2262 87196 -2026
rect 86876 -2294 87196 -2262
rect 92144 705238 92464 706230
rect 92144 705002 92186 705238
rect 92422 705002 92464 705238
rect 92144 704918 92464 705002
rect 92144 704682 92186 704918
rect 92422 704682 92464 704918
rect 92144 695494 92464 704682
rect 92144 695258 92186 695494
rect 92422 695258 92464 695494
rect 92144 688494 92464 695258
rect 92144 688258 92186 688494
rect 92422 688258 92464 688494
rect 92144 681494 92464 688258
rect 92144 681258 92186 681494
rect 92422 681258 92464 681494
rect 92144 674494 92464 681258
rect 92144 674258 92186 674494
rect 92422 674258 92464 674494
rect 92144 667494 92464 674258
rect 92144 667258 92186 667494
rect 92422 667258 92464 667494
rect 92144 660494 92464 667258
rect 92144 660258 92186 660494
rect 92422 660258 92464 660494
rect 92144 653494 92464 660258
rect 92144 653258 92186 653494
rect 92422 653258 92464 653494
rect 92144 646494 92464 653258
rect 92144 646258 92186 646494
rect 92422 646258 92464 646494
rect 92144 639494 92464 646258
rect 92144 639258 92186 639494
rect 92422 639258 92464 639494
rect 92144 632494 92464 639258
rect 92144 632258 92186 632494
rect 92422 632258 92464 632494
rect 92144 625494 92464 632258
rect 92144 625258 92186 625494
rect 92422 625258 92464 625494
rect 92144 618494 92464 625258
rect 92144 618258 92186 618494
rect 92422 618258 92464 618494
rect 92144 611494 92464 618258
rect 92144 611258 92186 611494
rect 92422 611258 92464 611494
rect 92144 604494 92464 611258
rect 92144 604258 92186 604494
rect 92422 604258 92464 604494
rect 92144 597494 92464 604258
rect 92144 597258 92186 597494
rect 92422 597258 92464 597494
rect 92144 590494 92464 597258
rect 92144 590258 92186 590494
rect 92422 590258 92464 590494
rect 92144 583494 92464 590258
rect 92144 583258 92186 583494
rect 92422 583258 92464 583494
rect 92144 576494 92464 583258
rect 92144 576258 92186 576494
rect 92422 576258 92464 576494
rect 92144 569494 92464 576258
rect 92144 569258 92186 569494
rect 92422 569258 92464 569494
rect 92144 562494 92464 569258
rect 92144 562258 92186 562494
rect 92422 562258 92464 562494
rect 92144 555494 92464 562258
rect 92144 555258 92186 555494
rect 92422 555258 92464 555494
rect 92144 548494 92464 555258
rect 92144 548258 92186 548494
rect 92422 548258 92464 548494
rect 92144 541494 92464 548258
rect 92144 541258 92186 541494
rect 92422 541258 92464 541494
rect 92144 534494 92464 541258
rect 92144 534258 92186 534494
rect 92422 534258 92464 534494
rect 92144 527494 92464 534258
rect 92144 527258 92186 527494
rect 92422 527258 92464 527494
rect 92144 520494 92464 527258
rect 92144 520258 92186 520494
rect 92422 520258 92464 520494
rect 92144 513494 92464 520258
rect 92144 513258 92186 513494
rect 92422 513258 92464 513494
rect 92144 506494 92464 513258
rect 92144 506258 92186 506494
rect 92422 506258 92464 506494
rect 92144 499494 92464 506258
rect 92144 499258 92186 499494
rect 92422 499258 92464 499494
rect 92144 492494 92464 499258
rect 92144 492258 92186 492494
rect 92422 492258 92464 492494
rect 92144 485494 92464 492258
rect 92144 485258 92186 485494
rect 92422 485258 92464 485494
rect 92144 478494 92464 485258
rect 92144 478258 92186 478494
rect 92422 478258 92464 478494
rect 92144 471494 92464 478258
rect 92144 471258 92186 471494
rect 92422 471258 92464 471494
rect 92144 464494 92464 471258
rect 92144 464258 92186 464494
rect 92422 464258 92464 464494
rect 92144 457494 92464 464258
rect 92144 457258 92186 457494
rect 92422 457258 92464 457494
rect 92144 450494 92464 457258
rect 92144 450258 92186 450494
rect 92422 450258 92464 450494
rect 92144 443494 92464 450258
rect 92144 443258 92186 443494
rect 92422 443258 92464 443494
rect 92144 436494 92464 443258
rect 92144 436258 92186 436494
rect 92422 436258 92464 436494
rect 92144 429494 92464 436258
rect 92144 429258 92186 429494
rect 92422 429258 92464 429494
rect 92144 422494 92464 429258
rect 92144 422258 92186 422494
rect 92422 422258 92464 422494
rect 92144 415494 92464 422258
rect 92144 415258 92186 415494
rect 92422 415258 92464 415494
rect 92144 408494 92464 415258
rect 92144 408258 92186 408494
rect 92422 408258 92464 408494
rect 92144 401494 92464 408258
rect 92144 401258 92186 401494
rect 92422 401258 92464 401494
rect 92144 394494 92464 401258
rect 92144 394258 92186 394494
rect 92422 394258 92464 394494
rect 92144 387494 92464 394258
rect 92144 387258 92186 387494
rect 92422 387258 92464 387494
rect 92144 380494 92464 387258
rect 92144 380258 92186 380494
rect 92422 380258 92464 380494
rect 92144 373494 92464 380258
rect 92144 373258 92186 373494
rect 92422 373258 92464 373494
rect 92144 366494 92464 373258
rect 92144 366258 92186 366494
rect 92422 366258 92464 366494
rect 92144 359494 92464 366258
rect 92144 359258 92186 359494
rect 92422 359258 92464 359494
rect 92144 352494 92464 359258
rect 92144 352258 92186 352494
rect 92422 352258 92464 352494
rect 92144 345494 92464 352258
rect 92144 345258 92186 345494
rect 92422 345258 92464 345494
rect 92144 338494 92464 345258
rect 92144 338258 92186 338494
rect 92422 338258 92464 338494
rect 92144 331494 92464 338258
rect 92144 331258 92186 331494
rect 92422 331258 92464 331494
rect 92144 324494 92464 331258
rect 92144 324258 92186 324494
rect 92422 324258 92464 324494
rect 92144 317494 92464 324258
rect 92144 317258 92186 317494
rect 92422 317258 92464 317494
rect 92144 310494 92464 317258
rect 92144 310258 92186 310494
rect 92422 310258 92464 310494
rect 92144 303494 92464 310258
rect 92144 303258 92186 303494
rect 92422 303258 92464 303494
rect 92144 296494 92464 303258
rect 92144 296258 92186 296494
rect 92422 296258 92464 296494
rect 92144 289494 92464 296258
rect 92144 289258 92186 289494
rect 92422 289258 92464 289494
rect 92144 282494 92464 289258
rect 92144 282258 92186 282494
rect 92422 282258 92464 282494
rect 92144 275494 92464 282258
rect 92144 275258 92186 275494
rect 92422 275258 92464 275494
rect 92144 268494 92464 275258
rect 92144 268258 92186 268494
rect 92422 268258 92464 268494
rect 92144 261494 92464 268258
rect 92144 261258 92186 261494
rect 92422 261258 92464 261494
rect 92144 254494 92464 261258
rect 92144 254258 92186 254494
rect 92422 254258 92464 254494
rect 92144 247494 92464 254258
rect 92144 247258 92186 247494
rect 92422 247258 92464 247494
rect 92144 240494 92464 247258
rect 92144 240258 92186 240494
rect 92422 240258 92464 240494
rect 92144 233494 92464 240258
rect 92144 233258 92186 233494
rect 92422 233258 92464 233494
rect 92144 226494 92464 233258
rect 92144 226258 92186 226494
rect 92422 226258 92464 226494
rect 92144 219494 92464 226258
rect 92144 219258 92186 219494
rect 92422 219258 92464 219494
rect 92144 212494 92464 219258
rect 92144 212258 92186 212494
rect 92422 212258 92464 212494
rect 92144 205494 92464 212258
rect 92144 205258 92186 205494
rect 92422 205258 92464 205494
rect 92144 198494 92464 205258
rect 92144 198258 92186 198494
rect 92422 198258 92464 198494
rect 92144 191494 92464 198258
rect 92144 191258 92186 191494
rect 92422 191258 92464 191494
rect 92144 184494 92464 191258
rect 92144 184258 92186 184494
rect 92422 184258 92464 184494
rect 92144 177494 92464 184258
rect 92144 177258 92186 177494
rect 92422 177258 92464 177494
rect 92144 170494 92464 177258
rect 92144 170258 92186 170494
rect 92422 170258 92464 170494
rect 92144 163494 92464 170258
rect 92144 163258 92186 163494
rect 92422 163258 92464 163494
rect 92144 156494 92464 163258
rect 92144 156258 92186 156494
rect 92422 156258 92464 156494
rect 92144 149494 92464 156258
rect 92144 149258 92186 149494
rect 92422 149258 92464 149494
rect 92144 142494 92464 149258
rect 92144 142258 92186 142494
rect 92422 142258 92464 142494
rect 92144 135494 92464 142258
rect 92144 135258 92186 135494
rect 92422 135258 92464 135494
rect 92144 128494 92464 135258
rect 92144 128258 92186 128494
rect 92422 128258 92464 128494
rect 92144 121494 92464 128258
rect 92144 121258 92186 121494
rect 92422 121258 92464 121494
rect 92144 114494 92464 121258
rect 92144 114258 92186 114494
rect 92422 114258 92464 114494
rect 92144 107494 92464 114258
rect 92144 107258 92186 107494
rect 92422 107258 92464 107494
rect 92144 100494 92464 107258
rect 92144 100258 92186 100494
rect 92422 100258 92464 100494
rect 92144 93494 92464 100258
rect 92144 93258 92186 93494
rect 92422 93258 92464 93494
rect 92144 86494 92464 93258
rect 92144 86258 92186 86494
rect 92422 86258 92464 86494
rect 92144 79494 92464 86258
rect 92144 79258 92186 79494
rect 92422 79258 92464 79494
rect 92144 72494 92464 79258
rect 92144 72258 92186 72494
rect 92422 72258 92464 72494
rect 92144 65494 92464 72258
rect 92144 65258 92186 65494
rect 92422 65258 92464 65494
rect 92144 58494 92464 65258
rect 92144 58258 92186 58494
rect 92422 58258 92464 58494
rect 92144 51494 92464 58258
rect 92144 51258 92186 51494
rect 92422 51258 92464 51494
rect 92144 44494 92464 51258
rect 92144 44258 92186 44494
rect 92422 44258 92464 44494
rect 92144 37494 92464 44258
rect 92144 37258 92186 37494
rect 92422 37258 92464 37494
rect 92144 30494 92464 37258
rect 92144 30258 92186 30494
rect 92422 30258 92464 30494
rect 92144 23494 92464 30258
rect 92144 23258 92186 23494
rect 92422 23258 92464 23494
rect 92144 16494 92464 23258
rect 92144 16258 92186 16494
rect 92422 16258 92464 16494
rect 92144 9494 92464 16258
rect 92144 9258 92186 9494
rect 92422 9258 92464 9494
rect 92144 2494 92464 9258
rect 92144 2258 92186 2494
rect 92422 2258 92464 2494
rect 92144 -746 92464 2258
rect 92144 -982 92186 -746
rect 92422 -982 92464 -746
rect 92144 -1066 92464 -982
rect 92144 -1302 92186 -1066
rect 92422 -1302 92464 -1066
rect 92144 -2294 92464 -1302
rect 93876 706198 94196 706230
rect 93876 705962 93918 706198
rect 94154 705962 94196 706198
rect 93876 705878 94196 705962
rect 93876 705642 93918 705878
rect 94154 705642 94196 705878
rect 93876 696561 94196 705642
rect 93876 696325 93918 696561
rect 94154 696325 94196 696561
rect 93876 689561 94196 696325
rect 93876 689325 93918 689561
rect 94154 689325 94196 689561
rect 93876 682561 94196 689325
rect 93876 682325 93918 682561
rect 94154 682325 94196 682561
rect 93876 675561 94196 682325
rect 93876 675325 93918 675561
rect 94154 675325 94196 675561
rect 93876 668561 94196 675325
rect 93876 668325 93918 668561
rect 94154 668325 94196 668561
rect 93876 661561 94196 668325
rect 93876 661325 93918 661561
rect 94154 661325 94196 661561
rect 93876 654561 94196 661325
rect 93876 654325 93918 654561
rect 94154 654325 94196 654561
rect 93876 647561 94196 654325
rect 93876 647325 93918 647561
rect 94154 647325 94196 647561
rect 93876 640561 94196 647325
rect 93876 640325 93918 640561
rect 94154 640325 94196 640561
rect 93876 633561 94196 640325
rect 93876 633325 93918 633561
rect 94154 633325 94196 633561
rect 93876 626561 94196 633325
rect 93876 626325 93918 626561
rect 94154 626325 94196 626561
rect 93876 619561 94196 626325
rect 93876 619325 93918 619561
rect 94154 619325 94196 619561
rect 93876 612561 94196 619325
rect 93876 612325 93918 612561
rect 94154 612325 94196 612561
rect 93876 605561 94196 612325
rect 93876 605325 93918 605561
rect 94154 605325 94196 605561
rect 93876 598561 94196 605325
rect 93876 598325 93918 598561
rect 94154 598325 94196 598561
rect 93876 591561 94196 598325
rect 93876 591325 93918 591561
rect 94154 591325 94196 591561
rect 93876 584561 94196 591325
rect 93876 584325 93918 584561
rect 94154 584325 94196 584561
rect 93876 577561 94196 584325
rect 93876 577325 93918 577561
rect 94154 577325 94196 577561
rect 93876 570561 94196 577325
rect 93876 570325 93918 570561
rect 94154 570325 94196 570561
rect 93876 563561 94196 570325
rect 93876 563325 93918 563561
rect 94154 563325 94196 563561
rect 93876 556561 94196 563325
rect 93876 556325 93918 556561
rect 94154 556325 94196 556561
rect 93876 549561 94196 556325
rect 93876 549325 93918 549561
rect 94154 549325 94196 549561
rect 93876 542561 94196 549325
rect 93876 542325 93918 542561
rect 94154 542325 94196 542561
rect 93876 535561 94196 542325
rect 93876 535325 93918 535561
rect 94154 535325 94196 535561
rect 93876 528561 94196 535325
rect 93876 528325 93918 528561
rect 94154 528325 94196 528561
rect 93876 521561 94196 528325
rect 93876 521325 93918 521561
rect 94154 521325 94196 521561
rect 93876 514561 94196 521325
rect 93876 514325 93918 514561
rect 94154 514325 94196 514561
rect 93876 507561 94196 514325
rect 93876 507325 93918 507561
rect 94154 507325 94196 507561
rect 93876 500561 94196 507325
rect 93876 500325 93918 500561
rect 94154 500325 94196 500561
rect 93876 493561 94196 500325
rect 93876 493325 93918 493561
rect 94154 493325 94196 493561
rect 93876 486561 94196 493325
rect 93876 486325 93918 486561
rect 94154 486325 94196 486561
rect 93876 479561 94196 486325
rect 93876 479325 93918 479561
rect 94154 479325 94196 479561
rect 93876 472561 94196 479325
rect 93876 472325 93918 472561
rect 94154 472325 94196 472561
rect 93876 465561 94196 472325
rect 93876 465325 93918 465561
rect 94154 465325 94196 465561
rect 93876 458561 94196 465325
rect 93876 458325 93918 458561
rect 94154 458325 94196 458561
rect 93876 451561 94196 458325
rect 93876 451325 93918 451561
rect 94154 451325 94196 451561
rect 93876 444561 94196 451325
rect 93876 444325 93918 444561
rect 94154 444325 94196 444561
rect 93876 437561 94196 444325
rect 93876 437325 93918 437561
rect 94154 437325 94196 437561
rect 93876 430561 94196 437325
rect 93876 430325 93918 430561
rect 94154 430325 94196 430561
rect 93876 423561 94196 430325
rect 93876 423325 93918 423561
rect 94154 423325 94196 423561
rect 93876 416561 94196 423325
rect 93876 416325 93918 416561
rect 94154 416325 94196 416561
rect 93876 409561 94196 416325
rect 93876 409325 93918 409561
rect 94154 409325 94196 409561
rect 93876 402561 94196 409325
rect 93876 402325 93918 402561
rect 94154 402325 94196 402561
rect 93876 395561 94196 402325
rect 93876 395325 93918 395561
rect 94154 395325 94196 395561
rect 93876 388561 94196 395325
rect 93876 388325 93918 388561
rect 94154 388325 94196 388561
rect 93876 381561 94196 388325
rect 93876 381325 93918 381561
rect 94154 381325 94196 381561
rect 93876 374561 94196 381325
rect 93876 374325 93918 374561
rect 94154 374325 94196 374561
rect 93876 367561 94196 374325
rect 93876 367325 93918 367561
rect 94154 367325 94196 367561
rect 93876 360561 94196 367325
rect 93876 360325 93918 360561
rect 94154 360325 94196 360561
rect 93876 353561 94196 360325
rect 93876 353325 93918 353561
rect 94154 353325 94196 353561
rect 93876 346561 94196 353325
rect 93876 346325 93918 346561
rect 94154 346325 94196 346561
rect 93876 339561 94196 346325
rect 93876 339325 93918 339561
rect 94154 339325 94196 339561
rect 93876 332561 94196 339325
rect 93876 332325 93918 332561
rect 94154 332325 94196 332561
rect 93876 325561 94196 332325
rect 93876 325325 93918 325561
rect 94154 325325 94196 325561
rect 93876 318561 94196 325325
rect 93876 318325 93918 318561
rect 94154 318325 94196 318561
rect 93876 311561 94196 318325
rect 93876 311325 93918 311561
rect 94154 311325 94196 311561
rect 93876 304561 94196 311325
rect 93876 304325 93918 304561
rect 94154 304325 94196 304561
rect 93876 297561 94196 304325
rect 93876 297325 93918 297561
rect 94154 297325 94196 297561
rect 93876 290561 94196 297325
rect 93876 290325 93918 290561
rect 94154 290325 94196 290561
rect 93876 283561 94196 290325
rect 93876 283325 93918 283561
rect 94154 283325 94196 283561
rect 93876 276561 94196 283325
rect 93876 276325 93918 276561
rect 94154 276325 94196 276561
rect 93876 269561 94196 276325
rect 93876 269325 93918 269561
rect 94154 269325 94196 269561
rect 93876 262561 94196 269325
rect 93876 262325 93918 262561
rect 94154 262325 94196 262561
rect 93876 255561 94196 262325
rect 93876 255325 93918 255561
rect 94154 255325 94196 255561
rect 93876 248561 94196 255325
rect 93876 248325 93918 248561
rect 94154 248325 94196 248561
rect 93876 241561 94196 248325
rect 93876 241325 93918 241561
rect 94154 241325 94196 241561
rect 93876 234561 94196 241325
rect 93876 234325 93918 234561
rect 94154 234325 94196 234561
rect 93876 227561 94196 234325
rect 93876 227325 93918 227561
rect 94154 227325 94196 227561
rect 93876 220561 94196 227325
rect 93876 220325 93918 220561
rect 94154 220325 94196 220561
rect 93876 213561 94196 220325
rect 93876 213325 93918 213561
rect 94154 213325 94196 213561
rect 93876 206561 94196 213325
rect 93876 206325 93918 206561
rect 94154 206325 94196 206561
rect 93876 199561 94196 206325
rect 93876 199325 93918 199561
rect 94154 199325 94196 199561
rect 93876 192561 94196 199325
rect 93876 192325 93918 192561
rect 94154 192325 94196 192561
rect 93876 185561 94196 192325
rect 93876 185325 93918 185561
rect 94154 185325 94196 185561
rect 93876 178561 94196 185325
rect 93876 178325 93918 178561
rect 94154 178325 94196 178561
rect 93876 171561 94196 178325
rect 93876 171325 93918 171561
rect 94154 171325 94196 171561
rect 93876 164561 94196 171325
rect 93876 164325 93918 164561
rect 94154 164325 94196 164561
rect 93876 157561 94196 164325
rect 93876 157325 93918 157561
rect 94154 157325 94196 157561
rect 93876 150561 94196 157325
rect 93876 150325 93918 150561
rect 94154 150325 94196 150561
rect 93876 143561 94196 150325
rect 93876 143325 93918 143561
rect 94154 143325 94196 143561
rect 93876 136561 94196 143325
rect 93876 136325 93918 136561
rect 94154 136325 94196 136561
rect 93876 129561 94196 136325
rect 93876 129325 93918 129561
rect 94154 129325 94196 129561
rect 93876 122561 94196 129325
rect 93876 122325 93918 122561
rect 94154 122325 94196 122561
rect 93876 115561 94196 122325
rect 93876 115325 93918 115561
rect 94154 115325 94196 115561
rect 93876 108561 94196 115325
rect 93876 108325 93918 108561
rect 94154 108325 94196 108561
rect 93876 101561 94196 108325
rect 93876 101325 93918 101561
rect 94154 101325 94196 101561
rect 93876 94561 94196 101325
rect 93876 94325 93918 94561
rect 94154 94325 94196 94561
rect 93876 87561 94196 94325
rect 93876 87325 93918 87561
rect 94154 87325 94196 87561
rect 93876 80561 94196 87325
rect 93876 80325 93918 80561
rect 94154 80325 94196 80561
rect 93876 73561 94196 80325
rect 93876 73325 93918 73561
rect 94154 73325 94196 73561
rect 93876 66561 94196 73325
rect 93876 66325 93918 66561
rect 94154 66325 94196 66561
rect 93876 59561 94196 66325
rect 93876 59325 93918 59561
rect 94154 59325 94196 59561
rect 93876 52561 94196 59325
rect 93876 52325 93918 52561
rect 94154 52325 94196 52561
rect 93876 45561 94196 52325
rect 93876 45325 93918 45561
rect 94154 45325 94196 45561
rect 93876 38561 94196 45325
rect 93876 38325 93918 38561
rect 94154 38325 94196 38561
rect 93876 31561 94196 38325
rect 93876 31325 93918 31561
rect 94154 31325 94196 31561
rect 93876 24561 94196 31325
rect 93876 24325 93918 24561
rect 94154 24325 94196 24561
rect 93876 17561 94196 24325
rect 93876 17325 93918 17561
rect 94154 17325 94196 17561
rect 93876 10561 94196 17325
rect 93876 10325 93918 10561
rect 94154 10325 94196 10561
rect 93876 3561 94196 10325
rect 93876 3325 93918 3561
rect 94154 3325 94196 3561
rect 93876 -1706 94196 3325
rect 93876 -1942 93918 -1706
rect 94154 -1942 94196 -1706
rect 93876 -2026 94196 -1942
rect 93876 -2262 93918 -2026
rect 94154 -2262 94196 -2026
rect 93876 -2294 94196 -2262
rect 99144 705238 99464 706230
rect 99144 705002 99186 705238
rect 99422 705002 99464 705238
rect 99144 704918 99464 705002
rect 99144 704682 99186 704918
rect 99422 704682 99464 704918
rect 99144 695494 99464 704682
rect 99144 695258 99186 695494
rect 99422 695258 99464 695494
rect 99144 688494 99464 695258
rect 99144 688258 99186 688494
rect 99422 688258 99464 688494
rect 99144 681494 99464 688258
rect 99144 681258 99186 681494
rect 99422 681258 99464 681494
rect 99144 674494 99464 681258
rect 99144 674258 99186 674494
rect 99422 674258 99464 674494
rect 99144 667494 99464 674258
rect 99144 667258 99186 667494
rect 99422 667258 99464 667494
rect 99144 660494 99464 667258
rect 99144 660258 99186 660494
rect 99422 660258 99464 660494
rect 99144 653494 99464 660258
rect 99144 653258 99186 653494
rect 99422 653258 99464 653494
rect 99144 646494 99464 653258
rect 99144 646258 99186 646494
rect 99422 646258 99464 646494
rect 99144 639494 99464 646258
rect 99144 639258 99186 639494
rect 99422 639258 99464 639494
rect 99144 632494 99464 639258
rect 99144 632258 99186 632494
rect 99422 632258 99464 632494
rect 99144 625494 99464 632258
rect 99144 625258 99186 625494
rect 99422 625258 99464 625494
rect 99144 618494 99464 625258
rect 99144 618258 99186 618494
rect 99422 618258 99464 618494
rect 99144 611494 99464 618258
rect 99144 611258 99186 611494
rect 99422 611258 99464 611494
rect 99144 604494 99464 611258
rect 99144 604258 99186 604494
rect 99422 604258 99464 604494
rect 99144 597494 99464 604258
rect 99144 597258 99186 597494
rect 99422 597258 99464 597494
rect 99144 590494 99464 597258
rect 99144 590258 99186 590494
rect 99422 590258 99464 590494
rect 99144 583494 99464 590258
rect 99144 583258 99186 583494
rect 99422 583258 99464 583494
rect 99144 576494 99464 583258
rect 99144 576258 99186 576494
rect 99422 576258 99464 576494
rect 99144 569494 99464 576258
rect 99144 569258 99186 569494
rect 99422 569258 99464 569494
rect 99144 562494 99464 569258
rect 99144 562258 99186 562494
rect 99422 562258 99464 562494
rect 99144 555494 99464 562258
rect 99144 555258 99186 555494
rect 99422 555258 99464 555494
rect 99144 548494 99464 555258
rect 99144 548258 99186 548494
rect 99422 548258 99464 548494
rect 99144 541494 99464 548258
rect 99144 541258 99186 541494
rect 99422 541258 99464 541494
rect 99144 534494 99464 541258
rect 99144 534258 99186 534494
rect 99422 534258 99464 534494
rect 99144 527494 99464 534258
rect 99144 527258 99186 527494
rect 99422 527258 99464 527494
rect 99144 520494 99464 527258
rect 99144 520258 99186 520494
rect 99422 520258 99464 520494
rect 99144 513494 99464 520258
rect 99144 513258 99186 513494
rect 99422 513258 99464 513494
rect 99144 506494 99464 513258
rect 99144 506258 99186 506494
rect 99422 506258 99464 506494
rect 99144 499494 99464 506258
rect 99144 499258 99186 499494
rect 99422 499258 99464 499494
rect 99144 492494 99464 499258
rect 99144 492258 99186 492494
rect 99422 492258 99464 492494
rect 99144 485494 99464 492258
rect 99144 485258 99186 485494
rect 99422 485258 99464 485494
rect 99144 478494 99464 485258
rect 99144 478258 99186 478494
rect 99422 478258 99464 478494
rect 99144 471494 99464 478258
rect 99144 471258 99186 471494
rect 99422 471258 99464 471494
rect 99144 464494 99464 471258
rect 99144 464258 99186 464494
rect 99422 464258 99464 464494
rect 99144 457494 99464 464258
rect 99144 457258 99186 457494
rect 99422 457258 99464 457494
rect 99144 450494 99464 457258
rect 99144 450258 99186 450494
rect 99422 450258 99464 450494
rect 99144 443494 99464 450258
rect 99144 443258 99186 443494
rect 99422 443258 99464 443494
rect 99144 436494 99464 443258
rect 99144 436258 99186 436494
rect 99422 436258 99464 436494
rect 99144 429494 99464 436258
rect 99144 429258 99186 429494
rect 99422 429258 99464 429494
rect 99144 422494 99464 429258
rect 99144 422258 99186 422494
rect 99422 422258 99464 422494
rect 99144 415494 99464 422258
rect 99144 415258 99186 415494
rect 99422 415258 99464 415494
rect 99144 408494 99464 415258
rect 99144 408258 99186 408494
rect 99422 408258 99464 408494
rect 99144 401494 99464 408258
rect 99144 401258 99186 401494
rect 99422 401258 99464 401494
rect 99144 394494 99464 401258
rect 99144 394258 99186 394494
rect 99422 394258 99464 394494
rect 99144 387494 99464 394258
rect 99144 387258 99186 387494
rect 99422 387258 99464 387494
rect 99144 380494 99464 387258
rect 99144 380258 99186 380494
rect 99422 380258 99464 380494
rect 99144 373494 99464 380258
rect 99144 373258 99186 373494
rect 99422 373258 99464 373494
rect 99144 366494 99464 373258
rect 99144 366258 99186 366494
rect 99422 366258 99464 366494
rect 99144 359494 99464 366258
rect 99144 359258 99186 359494
rect 99422 359258 99464 359494
rect 99144 352494 99464 359258
rect 99144 352258 99186 352494
rect 99422 352258 99464 352494
rect 99144 345494 99464 352258
rect 99144 345258 99186 345494
rect 99422 345258 99464 345494
rect 99144 338494 99464 345258
rect 99144 338258 99186 338494
rect 99422 338258 99464 338494
rect 99144 331494 99464 338258
rect 99144 331258 99186 331494
rect 99422 331258 99464 331494
rect 99144 324494 99464 331258
rect 99144 324258 99186 324494
rect 99422 324258 99464 324494
rect 99144 317494 99464 324258
rect 99144 317258 99186 317494
rect 99422 317258 99464 317494
rect 99144 310494 99464 317258
rect 99144 310258 99186 310494
rect 99422 310258 99464 310494
rect 99144 303494 99464 310258
rect 99144 303258 99186 303494
rect 99422 303258 99464 303494
rect 99144 296494 99464 303258
rect 99144 296258 99186 296494
rect 99422 296258 99464 296494
rect 99144 289494 99464 296258
rect 99144 289258 99186 289494
rect 99422 289258 99464 289494
rect 99144 282494 99464 289258
rect 99144 282258 99186 282494
rect 99422 282258 99464 282494
rect 99144 275494 99464 282258
rect 99144 275258 99186 275494
rect 99422 275258 99464 275494
rect 99144 268494 99464 275258
rect 99144 268258 99186 268494
rect 99422 268258 99464 268494
rect 99144 261494 99464 268258
rect 99144 261258 99186 261494
rect 99422 261258 99464 261494
rect 99144 254494 99464 261258
rect 99144 254258 99186 254494
rect 99422 254258 99464 254494
rect 99144 247494 99464 254258
rect 99144 247258 99186 247494
rect 99422 247258 99464 247494
rect 99144 240494 99464 247258
rect 99144 240258 99186 240494
rect 99422 240258 99464 240494
rect 99144 233494 99464 240258
rect 99144 233258 99186 233494
rect 99422 233258 99464 233494
rect 99144 226494 99464 233258
rect 99144 226258 99186 226494
rect 99422 226258 99464 226494
rect 99144 219494 99464 226258
rect 99144 219258 99186 219494
rect 99422 219258 99464 219494
rect 99144 212494 99464 219258
rect 99144 212258 99186 212494
rect 99422 212258 99464 212494
rect 99144 205494 99464 212258
rect 99144 205258 99186 205494
rect 99422 205258 99464 205494
rect 99144 198494 99464 205258
rect 99144 198258 99186 198494
rect 99422 198258 99464 198494
rect 99144 191494 99464 198258
rect 99144 191258 99186 191494
rect 99422 191258 99464 191494
rect 99144 184494 99464 191258
rect 99144 184258 99186 184494
rect 99422 184258 99464 184494
rect 99144 177494 99464 184258
rect 99144 177258 99186 177494
rect 99422 177258 99464 177494
rect 99144 170494 99464 177258
rect 99144 170258 99186 170494
rect 99422 170258 99464 170494
rect 99144 163494 99464 170258
rect 99144 163258 99186 163494
rect 99422 163258 99464 163494
rect 99144 156494 99464 163258
rect 99144 156258 99186 156494
rect 99422 156258 99464 156494
rect 99144 149494 99464 156258
rect 99144 149258 99186 149494
rect 99422 149258 99464 149494
rect 99144 142494 99464 149258
rect 99144 142258 99186 142494
rect 99422 142258 99464 142494
rect 99144 135494 99464 142258
rect 99144 135258 99186 135494
rect 99422 135258 99464 135494
rect 99144 128494 99464 135258
rect 99144 128258 99186 128494
rect 99422 128258 99464 128494
rect 99144 121494 99464 128258
rect 99144 121258 99186 121494
rect 99422 121258 99464 121494
rect 99144 114494 99464 121258
rect 99144 114258 99186 114494
rect 99422 114258 99464 114494
rect 99144 107494 99464 114258
rect 99144 107258 99186 107494
rect 99422 107258 99464 107494
rect 99144 100494 99464 107258
rect 99144 100258 99186 100494
rect 99422 100258 99464 100494
rect 99144 93494 99464 100258
rect 99144 93258 99186 93494
rect 99422 93258 99464 93494
rect 99144 86494 99464 93258
rect 99144 86258 99186 86494
rect 99422 86258 99464 86494
rect 99144 79494 99464 86258
rect 99144 79258 99186 79494
rect 99422 79258 99464 79494
rect 99144 72494 99464 79258
rect 99144 72258 99186 72494
rect 99422 72258 99464 72494
rect 99144 65494 99464 72258
rect 99144 65258 99186 65494
rect 99422 65258 99464 65494
rect 99144 58494 99464 65258
rect 99144 58258 99186 58494
rect 99422 58258 99464 58494
rect 99144 51494 99464 58258
rect 99144 51258 99186 51494
rect 99422 51258 99464 51494
rect 99144 44494 99464 51258
rect 99144 44258 99186 44494
rect 99422 44258 99464 44494
rect 99144 37494 99464 44258
rect 99144 37258 99186 37494
rect 99422 37258 99464 37494
rect 99144 30494 99464 37258
rect 99144 30258 99186 30494
rect 99422 30258 99464 30494
rect 99144 23494 99464 30258
rect 99144 23258 99186 23494
rect 99422 23258 99464 23494
rect 99144 16494 99464 23258
rect 99144 16258 99186 16494
rect 99422 16258 99464 16494
rect 99144 9494 99464 16258
rect 99144 9258 99186 9494
rect 99422 9258 99464 9494
rect 99144 2494 99464 9258
rect 99144 2258 99186 2494
rect 99422 2258 99464 2494
rect 99144 -746 99464 2258
rect 99144 -982 99186 -746
rect 99422 -982 99464 -746
rect 99144 -1066 99464 -982
rect 99144 -1302 99186 -1066
rect 99422 -1302 99464 -1066
rect 99144 -2294 99464 -1302
rect 100876 706198 101196 706230
rect 100876 705962 100918 706198
rect 101154 705962 101196 706198
rect 100876 705878 101196 705962
rect 100876 705642 100918 705878
rect 101154 705642 101196 705878
rect 100876 696561 101196 705642
rect 100876 696325 100918 696561
rect 101154 696325 101196 696561
rect 100876 689561 101196 696325
rect 100876 689325 100918 689561
rect 101154 689325 101196 689561
rect 100876 682561 101196 689325
rect 100876 682325 100918 682561
rect 101154 682325 101196 682561
rect 100876 675561 101196 682325
rect 100876 675325 100918 675561
rect 101154 675325 101196 675561
rect 100876 668561 101196 675325
rect 100876 668325 100918 668561
rect 101154 668325 101196 668561
rect 100876 661561 101196 668325
rect 100876 661325 100918 661561
rect 101154 661325 101196 661561
rect 100876 654561 101196 661325
rect 100876 654325 100918 654561
rect 101154 654325 101196 654561
rect 100876 647561 101196 654325
rect 100876 647325 100918 647561
rect 101154 647325 101196 647561
rect 100876 640561 101196 647325
rect 100876 640325 100918 640561
rect 101154 640325 101196 640561
rect 100876 633561 101196 640325
rect 100876 633325 100918 633561
rect 101154 633325 101196 633561
rect 100876 626561 101196 633325
rect 100876 626325 100918 626561
rect 101154 626325 101196 626561
rect 100876 619561 101196 626325
rect 100876 619325 100918 619561
rect 101154 619325 101196 619561
rect 100876 612561 101196 619325
rect 100876 612325 100918 612561
rect 101154 612325 101196 612561
rect 100876 605561 101196 612325
rect 100876 605325 100918 605561
rect 101154 605325 101196 605561
rect 100876 598561 101196 605325
rect 100876 598325 100918 598561
rect 101154 598325 101196 598561
rect 100876 591561 101196 598325
rect 100876 591325 100918 591561
rect 101154 591325 101196 591561
rect 100876 584561 101196 591325
rect 100876 584325 100918 584561
rect 101154 584325 101196 584561
rect 100876 577561 101196 584325
rect 100876 577325 100918 577561
rect 101154 577325 101196 577561
rect 100876 570561 101196 577325
rect 100876 570325 100918 570561
rect 101154 570325 101196 570561
rect 100876 563561 101196 570325
rect 100876 563325 100918 563561
rect 101154 563325 101196 563561
rect 100876 556561 101196 563325
rect 100876 556325 100918 556561
rect 101154 556325 101196 556561
rect 100876 549561 101196 556325
rect 100876 549325 100918 549561
rect 101154 549325 101196 549561
rect 100876 542561 101196 549325
rect 100876 542325 100918 542561
rect 101154 542325 101196 542561
rect 100876 535561 101196 542325
rect 100876 535325 100918 535561
rect 101154 535325 101196 535561
rect 100876 528561 101196 535325
rect 100876 528325 100918 528561
rect 101154 528325 101196 528561
rect 100876 521561 101196 528325
rect 100876 521325 100918 521561
rect 101154 521325 101196 521561
rect 100876 514561 101196 521325
rect 100876 514325 100918 514561
rect 101154 514325 101196 514561
rect 100876 507561 101196 514325
rect 100876 507325 100918 507561
rect 101154 507325 101196 507561
rect 100876 500561 101196 507325
rect 100876 500325 100918 500561
rect 101154 500325 101196 500561
rect 100876 493561 101196 500325
rect 100876 493325 100918 493561
rect 101154 493325 101196 493561
rect 100876 486561 101196 493325
rect 100876 486325 100918 486561
rect 101154 486325 101196 486561
rect 100876 479561 101196 486325
rect 100876 479325 100918 479561
rect 101154 479325 101196 479561
rect 100876 472561 101196 479325
rect 100876 472325 100918 472561
rect 101154 472325 101196 472561
rect 100876 465561 101196 472325
rect 100876 465325 100918 465561
rect 101154 465325 101196 465561
rect 100876 458561 101196 465325
rect 100876 458325 100918 458561
rect 101154 458325 101196 458561
rect 100876 451561 101196 458325
rect 100876 451325 100918 451561
rect 101154 451325 101196 451561
rect 100876 444561 101196 451325
rect 100876 444325 100918 444561
rect 101154 444325 101196 444561
rect 100876 437561 101196 444325
rect 100876 437325 100918 437561
rect 101154 437325 101196 437561
rect 100876 430561 101196 437325
rect 100876 430325 100918 430561
rect 101154 430325 101196 430561
rect 100876 423561 101196 430325
rect 100876 423325 100918 423561
rect 101154 423325 101196 423561
rect 100876 416561 101196 423325
rect 100876 416325 100918 416561
rect 101154 416325 101196 416561
rect 100876 409561 101196 416325
rect 100876 409325 100918 409561
rect 101154 409325 101196 409561
rect 100876 402561 101196 409325
rect 100876 402325 100918 402561
rect 101154 402325 101196 402561
rect 100876 395561 101196 402325
rect 100876 395325 100918 395561
rect 101154 395325 101196 395561
rect 100876 388561 101196 395325
rect 100876 388325 100918 388561
rect 101154 388325 101196 388561
rect 100876 381561 101196 388325
rect 100876 381325 100918 381561
rect 101154 381325 101196 381561
rect 100876 374561 101196 381325
rect 100876 374325 100918 374561
rect 101154 374325 101196 374561
rect 100876 367561 101196 374325
rect 100876 367325 100918 367561
rect 101154 367325 101196 367561
rect 100876 360561 101196 367325
rect 100876 360325 100918 360561
rect 101154 360325 101196 360561
rect 100876 353561 101196 360325
rect 100876 353325 100918 353561
rect 101154 353325 101196 353561
rect 100876 346561 101196 353325
rect 100876 346325 100918 346561
rect 101154 346325 101196 346561
rect 100876 339561 101196 346325
rect 100876 339325 100918 339561
rect 101154 339325 101196 339561
rect 100876 332561 101196 339325
rect 100876 332325 100918 332561
rect 101154 332325 101196 332561
rect 100876 325561 101196 332325
rect 100876 325325 100918 325561
rect 101154 325325 101196 325561
rect 100876 318561 101196 325325
rect 100876 318325 100918 318561
rect 101154 318325 101196 318561
rect 100876 311561 101196 318325
rect 100876 311325 100918 311561
rect 101154 311325 101196 311561
rect 100876 304561 101196 311325
rect 100876 304325 100918 304561
rect 101154 304325 101196 304561
rect 100876 297561 101196 304325
rect 100876 297325 100918 297561
rect 101154 297325 101196 297561
rect 100876 290561 101196 297325
rect 100876 290325 100918 290561
rect 101154 290325 101196 290561
rect 100876 283561 101196 290325
rect 100876 283325 100918 283561
rect 101154 283325 101196 283561
rect 100876 276561 101196 283325
rect 100876 276325 100918 276561
rect 101154 276325 101196 276561
rect 100876 269561 101196 276325
rect 100876 269325 100918 269561
rect 101154 269325 101196 269561
rect 100876 262561 101196 269325
rect 100876 262325 100918 262561
rect 101154 262325 101196 262561
rect 100876 255561 101196 262325
rect 100876 255325 100918 255561
rect 101154 255325 101196 255561
rect 100876 248561 101196 255325
rect 100876 248325 100918 248561
rect 101154 248325 101196 248561
rect 100876 241561 101196 248325
rect 100876 241325 100918 241561
rect 101154 241325 101196 241561
rect 100876 234561 101196 241325
rect 100876 234325 100918 234561
rect 101154 234325 101196 234561
rect 100876 227561 101196 234325
rect 100876 227325 100918 227561
rect 101154 227325 101196 227561
rect 100876 220561 101196 227325
rect 100876 220325 100918 220561
rect 101154 220325 101196 220561
rect 100876 213561 101196 220325
rect 100876 213325 100918 213561
rect 101154 213325 101196 213561
rect 100876 206561 101196 213325
rect 100876 206325 100918 206561
rect 101154 206325 101196 206561
rect 100876 199561 101196 206325
rect 100876 199325 100918 199561
rect 101154 199325 101196 199561
rect 100876 192561 101196 199325
rect 100876 192325 100918 192561
rect 101154 192325 101196 192561
rect 100876 185561 101196 192325
rect 100876 185325 100918 185561
rect 101154 185325 101196 185561
rect 100876 178561 101196 185325
rect 100876 178325 100918 178561
rect 101154 178325 101196 178561
rect 100876 171561 101196 178325
rect 100876 171325 100918 171561
rect 101154 171325 101196 171561
rect 100876 164561 101196 171325
rect 100876 164325 100918 164561
rect 101154 164325 101196 164561
rect 100876 157561 101196 164325
rect 100876 157325 100918 157561
rect 101154 157325 101196 157561
rect 100876 150561 101196 157325
rect 100876 150325 100918 150561
rect 101154 150325 101196 150561
rect 100876 143561 101196 150325
rect 100876 143325 100918 143561
rect 101154 143325 101196 143561
rect 100876 136561 101196 143325
rect 100876 136325 100918 136561
rect 101154 136325 101196 136561
rect 100876 129561 101196 136325
rect 100876 129325 100918 129561
rect 101154 129325 101196 129561
rect 100876 122561 101196 129325
rect 100876 122325 100918 122561
rect 101154 122325 101196 122561
rect 100876 115561 101196 122325
rect 100876 115325 100918 115561
rect 101154 115325 101196 115561
rect 100876 108561 101196 115325
rect 100876 108325 100918 108561
rect 101154 108325 101196 108561
rect 100876 101561 101196 108325
rect 100876 101325 100918 101561
rect 101154 101325 101196 101561
rect 100876 94561 101196 101325
rect 100876 94325 100918 94561
rect 101154 94325 101196 94561
rect 100876 87561 101196 94325
rect 100876 87325 100918 87561
rect 101154 87325 101196 87561
rect 100876 80561 101196 87325
rect 100876 80325 100918 80561
rect 101154 80325 101196 80561
rect 100876 73561 101196 80325
rect 100876 73325 100918 73561
rect 101154 73325 101196 73561
rect 100876 66561 101196 73325
rect 100876 66325 100918 66561
rect 101154 66325 101196 66561
rect 100876 59561 101196 66325
rect 100876 59325 100918 59561
rect 101154 59325 101196 59561
rect 100876 52561 101196 59325
rect 100876 52325 100918 52561
rect 101154 52325 101196 52561
rect 100876 45561 101196 52325
rect 100876 45325 100918 45561
rect 101154 45325 101196 45561
rect 100876 38561 101196 45325
rect 100876 38325 100918 38561
rect 101154 38325 101196 38561
rect 100876 31561 101196 38325
rect 100876 31325 100918 31561
rect 101154 31325 101196 31561
rect 100876 24561 101196 31325
rect 100876 24325 100918 24561
rect 101154 24325 101196 24561
rect 100876 17561 101196 24325
rect 100876 17325 100918 17561
rect 101154 17325 101196 17561
rect 100876 10561 101196 17325
rect 100876 10325 100918 10561
rect 101154 10325 101196 10561
rect 100876 3561 101196 10325
rect 100876 3325 100918 3561
rect 101154 3325 101196 3561
rect 100876 -1706 101196 3325
rect 100876 -1942 100918 -1706
rect 101154 -1942 101196 -1706
rect 100876 -2026 101196 -1942
rect 100876 -2262 100918 -2026
rect 101154 -2262 101196 -2026
rect 100876 -2294 101196 -2262
rect 106144 705238 106464 706230
rect 106144 705002 106186 705238
rect 106422 705002 106464 705238
rect 106144 704918 106464 705002
rect 106144 704682 106186 704918
rect 106422 704682 106464 704918
rect 106144 695494 106464 704682
rect 106144 695258 106186 695494
rect 106422 695258 106464 695494
rect 106144 688494 106464 695258
rect 106144 688258 106186 688494
rect 106422 688258 106464 688494
rect 106144 681494 106464 688258
rect 106144 681258 106186 681494
rect 106422 681258 106464 681494
rect 106144 674494 106464 681258
rect 106144 674258 106186 674494
rect 106422 674258 106464 674494
rect 106144 667494 106464 674258
rect 106144 667258 106186 667494
rect 106422 667258 106464 667494
rect 106144 660494 106464 667258
rect 106144 660258 106186 660494
rect 106422 660258 106464 660494
rect 106144 653494 106464 660258
rect 106144 653258 106186 653494
rect 106422 653258 106464 653494
rect 106144 646494 106464 653258
rect 106144 646258 106186 646494
rect 106422 646258 106464 646494
rect 106144 639494 106464 646258
rect 106144 639258 106186 639494
rect 106422 639258 106464 639494
rect 106144 632494 106464 639258
rect 106144 632258 106186 632494
rect 106422 632258 106464 632494
rect 106144 625494 106464 632258
rect 106144 625258 106186 625494
rect 106422 625258 106464 625494
rect 106144 618494 106464 625258
rect 106144 618258 106186 618494
rect 106422 618258 106464 618494
rect 106144 611494 106464 618258
rect 106144 611258 106186 611494
rect 106422 611258 106464 611494
rect 106144 604494 106464 611258
rect 106144 604258 106186 604494
rect 106422 604258 106464 604494
rect 106144 597494 106464 604258
rect 106144 597258 106186 597494
rect 106422 597258 106464 597494
rect 106144 590494 106464 597258
rect 106144 590258 106186 590494
rect 106422 590258 106464 590494
rect 106144 583494 106464 590258
rect 106144 583258 106186 583494
rect 106422 583258 106464 583494
rect 106144 576494 106464 583258
rect 106144 576258 106186 576494
rect 106422 576258 106464 576494
rect 106144 569494 106464 576258
rect 106144 569258 106186 569494
rect 106422 569258 106464 569494
rect 106144 562494 106464 569258
rect 106144 562258 106186 562494
rect 106422 562258 106464 562494
rect 106144 555494 106464 562258
rect 106144 555258 106186 555494
rect 106422 555258 106464 555494
rect 106144 548494 106464 555258
rect 106144 548258 106186 548494
rect 106422 548258 106464 548494
rect 106144 541494 106464 548258
rect 106144 541258 106186 541494
rect 106422 541258 106464 541494
rect 106144 534494 106464 541258
rect 106144 534258 106186 534494
rect 106422 534258 106464 534494
rect 106144 527494 106464 534258
rect 106144 527258 106186 527494
rect 106422 527258 106464 527494
rect 106144 520494 106464 527258
rect 106144 520258 106186 520494
rect 106422 520258 106464 520494
rect 106144 513494 106464 520258
rect 106144 513258 106186 513494
rect 106422 513258 106464 513494
rect 106144 506494 106464 513258
rect 106144 506258 106186 506494
rect 106422 506258 106464 506494
rect 106144 499494 106464 506258
rect 106144 499258 106186 499494
rect 106422 499258 106464 499494
rect 106144 492494 106464 499258
rect 106144 492258 106186 492494
rect 106422 492258 106464 492494
rect 106144 485494 106464 492258
rect 106144 485258 106186 485494
rect 106422 485258 106464 485494
rect 106144 478494 106464 485258
rect 106144 478258 106186 478494
rect 106422 478258 106464 478494
rect 106144 471494 106464 478258
rect 106144 471258 106186 471494
rect 106422 471258 106464 471494
rect 106144 464494 106464 471258
rect 106144 464258 106186 464494
rect 106422 464258 106464 464494
rect 106144 457494 106464 464258
rect 106144 457258 106186 457494
rect 106422 457258 106464 457494
rect 106144 450494 106464 457258
rect 106144 450258 106186 450494
rect 106422 450258 106464 450494
rect 106144 443494 106464 450258
rect 106144 443258 106186 443494
rect 106422 443258 106464 443494
rect 106144 436494 106464 443258
rect 106144 436258 106186 436494
rect 106422 436258 106464 436494
rect 106144 429494 106464 436258
rect 106144 429258 106186 429494
rect 106422 429258 106464 429494
rect 106144 422494 106464 429258
rect 106144 422258 106186 422494
rect 106422 422258 106464 422494
rect 106144 415494 106464 422258
rect 106144 415258 106186 415494
rect 106422 415258 106464 415494
rect 106144 408494 106464 415258
rect 106144 408258 106186 408494
rect 106422 408258 106464 408494
rect 106144 401494 106464 408258
rect 106144 401258 106186 401494
rect 106422 401258 106464 401494
rect 106144 394494 106464 401258
rect 106144 394258 106186 394494
rect 106422 394258 106464 394494
rect 106144 387494 106464 394258
rect 106144 387258 106186 387494
rect 106422 387258 106464 387494
rect 106144 380494 106464 387258
rect 106144 380258 106186 380494
rect 106422 380258 106464 380494
rect 106144 373494 106464 380258
rect 106144 373258 106186 373494
rect 106422 373258 106464 373494
rect 106144 366494 106464 373258
rect 106144 366258 106186 366494
rect 106422 366258 106464 366494
rect 106144 359494 106464 366258
rect 106144 359258 106186 359494
rect 106422 359258 106464 359494
rect 106144 352494 106464 359258
rect 106144 352258 106186 352494
rect 106422 352258 106464 352494
rect 106144 345494 106464 352258
rect 106144 345258 106186 345494
rect 106422 345258 106464 345494
rect 106144 338494 106464 345258
rect 106144 338258 106186 338494
rect 106422 338258 106464 338494
rect 106144 331494 106464 338258
rect 106144 331258 106186 331494
rect 106422 331258 106464 331494
rect 106144 324494 106464 331258
rect 106144 324258 106186 324494
rect 106422 324258 106464 324494
rect 106144 317494 106464 324258
rect 106144 317258 106186 317494
rect 106422 317258 106464 317494
rect 106144 310494 106464 317258
rect 106144 310258 106186 310494
rect 106422 310258 106464 310494
rect 106144 303494 106464 310258
rect 106144 303258 106186 303494
rect 106422 303258 106464 303494
rect 106144 296494 106464 303258
rect 106144 296258 106186 296494
rect 106422 296258 106464 296494
rect 106144 289494 106464 296258
rect 106144 289258 106186 289494
rect 106422 289258 106464 289494
rect 106144 282494 106464 289258
rect 106144 282258 106186 282494
rect 106422 282258 106464 282494
rect 106144 275494 106464 282258
rect 106144 275258 106186 275494
rect 106422 275258 106464 275494
rect 106144 268494 106464 275258
rect 106144 268258 106186 268494
rect 106422 268258 106464 268494
rect 106144 261494 106464 268258
rect 106144 261258 106186 261494
rect 106422 261258 106464 261494
rect 106144 254494 106464 261258
rect 106144 254258 106186 254494
rect 106422 254258 106464 254494
rect 106144 247494 106464 254258
rect 106144 247258 106186 247494
rect 106422 247258 106464 247494
rect 106144 240494 106464 247258
rect 106144 240258 106186 240494
rect 106422 240258 106464 240494
rect 106144 233494 106464 240258
rect 106144 233258 106186 233494
rect 106422 233258 106464 233494
rect 106144 226494 106464 233258
rect 106144 226258 106186 226494
rect 106422 226258 106464 226494
rect 106144 219494 106464 226258
rect 106144 219258 106186 219494
rect 106422 219258 106464 219494
rect 106144 212494 106464 219258
rect 106144 212258 106186 212494
rect 106422 212258 106464 212494
rect 106144 205494 106464 212258
rect 106144 205258 106186 205494
rect 106422 205258 106464 205494
rect 106144 198494 106464 205258
rect 106144 198258 106186 198494
rect 106422 198258 106464 198494
rect 106144 191494 106464 198258
rect 106144 191258 106186 191494
rect 106422 191258 106464 191494
rect 106144 184494 106464 191258
rect 106144 184258 106186 184494
rect 106422 184258 106464 184494
rect 106144 177494 106464 184258
rect 106144 177258 106186 177494
rect 106422 177258 106464 177494
rect 106144 170494 106464 177258
rect 106144 170258 106186 170494
rect 106422 170258 106464 170494
rect 106144 163494 106464 170258
rect 106144 163258 106186 163494
rect 106422 163258 106464 163494
rect 106144 156494 106464 163258
rect 106144 156258 106186 156494
rect 106422 156258 106464 156494
rect 106144 149494 106464 156258
rect 106144 149258 106186 149494
rect 106422 149258 106464 149494
rect 106144 142494 106464 149258
rect 106144 142258 106186 142494
rect 106422 142258 106464 142494
rect 106144 135494 106464 142258
rect 106144 135258 106186 135494
rect 106422 135258 106464 135494
rect 106144 128494 106464 135258
rect 106144 128258 106186 128494
rect 106422 128258 106464 128494
rect 106144 121494 106464 128258
rect 106144 121258 106186 121494
rect 106422 121258 106464 121494
rect 106144 114494 106464 121258
rect 106144 114258 106186 114494
rect 106422 114258 106464 114494
rect 106144 107494 106464 114258
rect 106144 107258 106186 107494
rect 106422 107258 106464 107494
rect 106144 100494 106464 107258
rect 106144 100258 106186 100494
rect 106422 100258 106464 100494
rect 106144 93494 106464 100258
rect 106144 93258 106186 93494
rect 106422 93258 106464 93494
rect 106144 86494 106464 93258
rect 106144 86258 106186 86494
rect 106422 86258 106464 86494
rect 106144 79494 106464 86258
rect 106144 79258 106186 79494
rect 106422 79258 106464 79494
rect 106144 72494 106464 79258
rect 106144 72258 106186 72494
rect 106422 72258 106464 72494
rect 106144 65494 106464 72258
rect 106144 65258 106186 65494
rect 106422 65258 106464 65494
rect 106144 58494 106464 65258
rect 106144 58258 106186 58494
rect 106422 58258 106464 58494
rect 106144 51494 106464 58258
rect 106144 51258 106186 51494
rect 106422 51258 106464 51494
rect 106144 44494 106464 51258
rect 106144 44258 106186 44494
rect 106422 44258 106464 44494
rect 106144 37494 106464 44258
rect 106144 37258 106186 37494
rect 106422 37258 106464 37494
rect 106144 30494 106464 37258
rect 106144 30258 106186 30494
rect 106422 30258 106464 30494
rect 106144 23494 106464 30258
rect 106144 23258 106186 23494
rect 106422 23258 106464 23494
rect 106144 16494 106464 23258
rect 106144 16258 106186 16494
rect 106422 16258 106464 16494
rect 106144 9494 106464 16258
rect 106144 9258 106186 9494
rect 106422 9258 106464 9494
rect 106144 2494 106464 9258
rect 106144 2258 106186 2494
rect 106422 2258 106464 2494
rect 106144 -746 106464 2258
rect 106144 -982 106186 -746
rect 106422 -982 106464 -746
rect 106144 -1066 106464 -982
rect 106144 -1302 106186 -1066
rect 106422 -1302 106464 -1066
rect 106144 -2294 106464 -1302
rect 107876 706198 108196 706230
rect 107876 705962 107918 706198
rect 108154 705962 108196 706198
rect 107876 705878 108196 705962
rect 107876 705642 107918 705878
rect 108154 705642 108196 705878
rect 107876 696561 108196 705642
rect 107876 696325 107918 696561
rect 108154 696325 108196 696561
rect 107876 689561 108196 696325
rect 107876 689325 107918 689561
rect 108154 689325 108196 689561
rect 107876 682561 108196 689325
rect 107876 682325 107918 682561
rect 108154 682325 108196 682561
rect 107876 675561 108196 682325
rect 107876 675325 107918 675561
rect 108154 675325 108196 675561
rect 107876 668561 108196 675325
rect 107876 668325 107918 668561
rect 108154 668325 108196 668561
rect 107876 661561 108196 668325
rect 107876 661325 107918 661561
rect 108154 661325 108196 661561
rect 107876 654561 108196 661325
rect 107876 654325 107918 654561
rect 108154 654325 108196 654561
rect 107876 647561 108196 654325
rect 107876 647325 107918 647561
rect 108154 647325 108196 647561
rect 107876 640561 108196 647325
rect 107876 640325 107918 640561
rect 108154 640325 108196 640561
rect 107876 633561 108196 640325
rect 107876 633325 107918 633561
rect 108154 633325 108196 633561
rect 107876 626561 108196 633325
rect 107876 626325 107918 626561
rect 108154 626325 108196 626561
rect 107876 619561 108196 626325
rect 107876 619325 107918 619561
rect 108154 619325 108196 619561
rect 107876 612561 108196 619325
rect 107876 612325 107918 612561
rect 108154 612325 108196 612561
rect 107876 605561 108196 612325
rect 107876 605325 107918 605561
rect 108154 605325 108196 605561
rect 107876 598561 108196 605325
rect 107876 598325 107918 598561
rect 108154 598325 108196 598561
rect 107876 591561 108196 598325
rect 107876 591325 107918 591561
rect 108154 591325 108196 591561
rect 107876 584561 108196 591325
rect 107876 584325 107918 584561
rect 108154 584325 108196 584561
rect 107876 577561 108196 584325
rect 107876 577325 107918 577561
rect 108154 577325 108196 577561
rect 107876 570561 108196 577325
rect 107876 570325 107918 570561
rect 108154 570325 108196 570561
rect 107876 563561 108196 570325
rect 107876 563325 107918 563561
rect 108154 563325 108196 563561
rect 107876 556561 108196 563325
rect 107876 556325 107918 556561
rect 108154 556325 108196 556561
rect 107876 549561 108196 556325
rect 107876 549325 107918 549561
rect 108154 549325 108196 549561
rect 107876 542561 108196 549325
rect 107876 542325 107918 542561
rect 108154 542325 108196 542561
rect 107876 535561 108196 542325
rect 107876 535325 107918 535561
rect 108154 535325 108196 535561
rect 107876 528561 108196 535325
rect 107876 528325 107918 528561
rect 108154 528325 108196 528561
rect 107876 521561 108196 528325
rect 107876 521325 107918 521561
rect 108154 521325 108196 521561
rect 107876 514561 108196 521325
rect 107876 514325 107918 514561
rect 108154 514325 108196 514561
rect 107876 507561 108196 514325
rect 107876 507325 107918 507561
rect 108154 507325 108196 507561
rect 107876 500561 108196 507325
rect 107876 500325 107918 500561
rect 108154 500325 108196 500561
rect 107876 493561 108196 500325
rect 107876 493325 107918 493561
rect 108154 493325 108196 493561
rect 107876 486561 108196 493325
rect 107876 486325 107918 486561
rect 108154 486325 108196 486561
rect 107876 479561 108196 486325
rect 107876 479325 107918 479561
rect 108154 479325 108196 479561
rect 107876 472561 108196 479325
rect 107876 472325 107918 472561
rect 108154 472325 108196 472561
rect 107876 465561 108196 472325
rect 107876 465325 107918 465561
rect 108154 465325 108196 465561
rect 107876 458561 108196 465325
rect 107876 458325 107918 458561
rect 108154 458325 108196 458561
rect 107876 451561 108196 458325
rect 107876 451325 107918 451561
rect 108154 451325 108196 451561
rect 107876 444561 108196 451325
rect 107876 444325 107918 444561
rect 108154 444325 108196 444561
rect 107876 437561 108196 444325
rect 107876 437325 107918 437561
rect 108154 437325 108196 437561
rect 107876 430561 108196 437325
rect 107876 430325 107918 430561
rect 108154 430325 108196 430561
rect 107876 423561 108196 430325
rect 107876 423325 107918 423561
rect 108154 423325 108196 423561
rect 107876 416561 108196 423325
rect 107876 416325 107918 416561
rect 108154 416325 108196 416561
rect 107876 409561 108196 416325
rect 107876 409325 107918 409561
rect 108154 409325 108196 409561
rect 107876 402561 108196 409325
rect 107876 402325 107918 402561
rect 108154 402325 108196 402561
rect 107876 395561 108196 402325
rect 107876 395325 107918 395561
rect 108154 395325 108196 395561
rect 107876 388561 108196 395325
rect 107876 388325 107918 388561
rect 108154 388325 108196 388561
rect 107876 381561 108196 388325
rect 107876 381325 107918 381561
rect 108154 381325 108196 381561
rect 107876 374561 108196 381325
rect 107876 374325 107918 374561
rect 108154 374325 108196 374561
rect 107876 367561 108196 374325
rect 107876 367325 107918 367561
rect 108154 367325 108196 367561
rect 107876 360561 108196 367325
rect 107876 360325 107918 360561
rect 108154 360325 108196 360561
rect 107876 353561 108196 360325
rect 107876 353325 107918 353561
rect 108154 353325 108196 353561
rect 107876 346561 108196 353325
rect 107876 346325 107918 346561
rect 108154 346325 108196 346561
rect 107876 339561 108196 346325
rect 107876 339325 107918 339561
rect 108154 339325 108196 339561
rect 107876 332561 108196 339325
rect 107876 332325 107918 332561
rect 108154 332325 108196 332561
rect 107876 325561 108196 332325
rect 107876 325325 107918 325561
rect 108154 325325 108196 325561
rect 107876 318561 108196 325325
rect 107876 318325 107918 318561
rect 108154 318325 108196 318561
rect 107876 311561 108196 318325
rect 107876 311325 107918 311561
rect 108154 311325 108196 311561
rect 107876 304561 108196 311325
rect 107876 304325 107918 304561
rect 108154 304325 108196 304561
rect 107876 297561 108196 304325
rect 107876 297325 107918 297561
rect 108154 297325 108196 297561
rect 107876 290561 108196 297325
rect 107876 290325 107918 290561
rect 108154 290325 108196 290561
rect 107876 283561 108196 290325
rect 107876 283325 107918 283561
rect 108154 283325 108196 283561
rect 107876 276561 108196 283325
rect 107876 276325 107918 276561
rect 108154 276325 108196 276561
rect 107876 269561 108196 276325
rect 107876 269325 107918 269561
rect 108154 269325 108196 269561
rect 107876 262561 108196 269325
rect 107876 262325 107918 262561
rect 108154 262325 108196 262561
rect 107876 255561 108196 262325
rect 107876 255325 107918 255561
rect 108154 255325 108196 255561
rect 107876 248561 108196 255325
rect 107876 248325 107918 248561
rect 108154 248325 108196 248561
rect 107876 241561 108196 248325
rect 107876 241325 107918 241561
rect 108154 241325 108196 241561
rect 107876 234561 108196 241325
rect 107876 234325 107918 234561
rect 108154 234325 108196 234561
rect 107876 227561 108196 234325
rect 107876 227325 107918 227561
rect 108154 227325 108196 227561
rect 107876 220561 108196 227325
rect 107876 220325 107918 220561
rect 108154 220325 108196 220561
rect 107876 213561 108196 220325
rect 107876 213325 107918 213561
rect 108154 213325 108196 213561
rect 107876 206561 108196 213325
rect 107876 206325 107918 206561
rect 108154 206325 108196 206561
rect 107876 199561 108196 206325
rect 107876 199325 107918 199561
rect 108154 199325 108196 199561
rect 107876 192561 108196 199325
rect 107876 192325 107918 192561
rect 108154 192325 108196 192561
rect 107876 185561 108196 192325
rect 107876 185325 107918 185561
rect 108154 185325 108196 185561
rect 107876 178561 108196 185325
rect 107876 178325 107918 178561
rect 108154 178325 108196 178561
rect 107876 171561 108196 178325
rect 107876 171325 107918 171561
rect 108154 171325 108196 171561
rect 107876 164561 108196 171325
rect 107876 164325 107918 164561
rect 108154 164325 108196 164561
rect 107876 157561 108196 164325
rect 107876 157325 107918 157561
rect 108154 157325 108196 157561
rect 107876 150561 108196 157325
rect 107876 150325 107918 150561
rect 108154 150325 108196 150561
rect 107876 143561 108196 150325
rect 107876 143325 107918 143561
rect 108154 143325 108196 143561
rect 107876 136561 108196 143325
rect 107876 136325 107918 136561
rect 108154 136325 108196 136561
rect 107876 129561 108196 136325
rect 107876 129325 107918 129561
rect 108154 129325 108196 129561
rect 107876 122561 108196 129325
rect 107876 122325 107918 122561
rect 108154 122325 108196 122561
rect 107876 115561 108196 122325
rect 107876 115325 107918 115561
rect 108154 115325 108196 115561
rect 107876 108561 108196 115325
rect 107876 108325 107918 108561
rect 108154 108325 108196 108561
rect 107876 101561 108196 108325
rect 107876 101325 107918 101561
rect 108154 101325 108196 101561
rect 107876 94561 108196 101325
rect 107876 94325 107918 94561
rect 108154 94325 108196 94561
rect 107876 87561 108196 94325
rect 107876 87325 107918 87561
rect 108154 87325 108196 87561
rect 107876 80561 108196 87325
rect 107876 80325 107918 80561
rect 108154 80325 108196 80561
rect 107876 73561 108196 80325
rect 107876 73325 107918 73561
rect 108154 73325 108196 73561
rect 107876 66561 108196 73325
rect 107876 66325 107918 66561
rect 108154 66325 108196 66561
rect 107876 59561 108196 66325
rect 107876 59325 107918 59561
rect 108154 59325 108196 59561
rect 107876 52561 108196 59325
rect 107876 52325 107918 52561
rect 108154 52325 108196 52561
rect 107876 45561 108196 52325
rect 107876 45325 107918 45561
rect 108154 45325 108196 45561
rect 107876 38561 108196 45325
rect 107876 38325 107918 38561
rect 108154 38325 108196 38561
rect 107876 31561 108196 38325
rect 107876 31325 107918 31561
rect 108154 31325 108196 31561
rect 107876 24561 108196 31325
rect 107876 24325 107918 24561
rect 108154 24325 108196 24561
rect 107876 17561 108196 24325
rect 107876 17325 107918 17561
rect 108154 17325 108196 17561
rect 107876 10561 108196 17325
rect 107876 10325 107918 10561
rect 108154 10325 108196 10561
rect 107876 3561 108196 10325
rect 107876 3325 107918 3561
rect 108154 3325 108196 3561
rect 107876 -1706 108196 3325
rect 107876 -1942 107918 -1706
rect 108154 -1942 108196 -1706
rect 107876 -2026 108196 -1942
rect 107876 -2262 107918 -2026
rect 108154 -2262 108196 -2026
rect 107876 -2294 108196 -2262
rect 113144 705238 113464 706230
rect 113144 705002 113186 705238
rect 113422 705002 113464 705238
rect 113144 704918 113464 705002
rect 113144 704682 113186 704918
rect 113422 704682 113464 704918
rect 113144 695494 113464 704682
rect 113144 695258 113186 695494
rect 113422 695258 113464 695494
rect 113144 688494 113464 695258
rect 113144 688258 113186 688494
rect 113422 688258 113464 688494
rect 113144 681494 113464 688258
rect 113144 681258 113186 681494
rect 113422 681258 113464 681494
rect 113144 674494 113464 681258
rect 113144 674258 113186 674494
rect 113422 674258 113464 674494
rect 113144 667494 113464 674258
rect 113144 667258 113186 667494
rect 113422 667258 113464 667494
rect 113144 660494 113464 667258
rect 113144 660258 113186 660494
rect 113422 660258 113464 660494
rect 113144 653494 113464 660258
rect 113144 653258 113186 653494
rect 113422 653258 113464 653494
rect 113144 646494 113464 653258
rect 113144 646258 113186 646494
rect 113422 646258 113464 646494
rect 113144 639494 113464 646258
rect 113144 639258 113186 639494
rect 113422 639258 113464 639494
rect 113144 632494 113464 639258
rect 113144 632258 113186 632494
rect 113422 632258 113464 632494
rect 113144 625494 113464 632258
rect 113144 625258 113186 625494
rect 113422 625258 113464 625494
rect 113144 618494 113464 625258
rect 113144 618258 113186 618494
rect 113422 618258 113464 618494
rect 113144 611494 113464 618258
rect 113144 611258 113186 611494
rect 113422 611258 113464 611494
rect 113144 604494 113464 611258
rect 113144 604258 113186 604494
rect 113422 604258 113464 604494
rect 113144 597494 113464 604258
rect 113144 597258 113186 597494
rect 113422 597258 113464 597494
rect 113144 590494 113464 597258
rect 113144 590258 113186 590494
rect 113422 590258 113464 590494
rect 113144 583494 113464 590258
rect 113144 583258 113186 583494
rect 113422 583258 113464 583494
rect 113144 576494 113464 583258
rect 113144 576258 113186 576494
rect 113422 576258 113464 576494
rect 113144 569494 113464 576258
rect 113144 569258 113186 569494
rect 113422 569258 113464 569494
rect 113144 562494 113464 569258
rect 113144 562258 113186 562494
rect 113422 562258 113464 562494
rect 113144 555494 113464 562258
rect 113144 555258 113186 555494
rect 113422 555258 113464 555494
rect 113144 548494 113464 555258
rect 113144 548258 113186 548494
rect 113422 548258 113464 548494
rect 113144 541494 113464 548258
rect 113144 541258 113186 541494
rect 113422 541258 113464 541494
rect 113144 534494 113464 541258
rect 113144 534258 113186 534494
rect 113422 534258 113464 534494
rect 113144 527494 113464 534258
rect 113144 527258 113186 527494
rect 113422 527258 113464 527494
rect 113144 520494 113464 527258
rect 113144 520258 113186 520494
rect 113422 520258 113464 520494
rect 113144 513494 113464 520258
rect 113144 513258 113186 513494
rect 113422 513258 113464 513494
rect 113144 506494 113464 513258
rect 113144 506258 113186 506494
rect 113422 506258 113464 506494
rect 113144 499494 113464 506258
rect 113144 499258 113186 499494
rect 113422 499258 113464 499494
rect 113144 492494 113464 499258
rect 113144 492258 113186 492494
rect 113422 492258 113464 492494
rect 113144 485494 113464 492258
rect 113144 485258 113186 485494
rect 113422 485258 113464 485494
rect 113144 478494 113464 485258
rect 113144 478258 113186 478494
rect 113422 478258 113464 478494
rect 113144 471494 113464 478258
rect 113144 471258 113186 471494
rect 113422 471258 113464 471494
rect 113144 464494 113464 471258
rect 113144 464258 113186 464494
rect 113422 464258 113464 464494
rect 113144 457494 113464 464258
rect 113144 457258 113186 457494
rect 113422 457258 113464 457494
rect 113144 450494 113464 457258
rect 113144 450258 113186 450494
rect 113422 450258 113464 450494
rect 113144 443494 113464 450258
rect 113144 443258 113186 443494
rect 113422 443258 113464 443494
rect 113144 436494 113464 443258
rect 113144 436258 113186 436494
rect 113422 436258 113464 436494
rect 113144 429494 113464 436258
rect 113144 429258 113186 429494
rect 113422 429258 113464 429494
rect 113144 422494 113464 429258
rect 113144 422258 113186 422494
rect 113422 422258 113464 422494
rect 113144 415494 113464 422258
rect 113144 415258 113186 415494
rect 113422 415258 113464 415494
rect 113144 408494 113464 415258
rect 113144 408258 113186 408494
rect 113422 408258 113464 408494
rect 113144 401494 113464 408258
rect 113144 401258 113186 401494
rect 113422 401258 113464 401494
rect 113144 394494 113464 401258
rect 113144 394258 113186 394494
rect 113422 394258 113464 394494
rect 113144 387494 113464 394258
rect 113144 387258 113186 387494
rect 113422 387258 113464 387494
rect 113144 380494 113464 387258
rect 113144 380258 113186 380494
rect 113422 380258 113464 380494
rect 113144 373494 113464 380258
rect 113144 373258 113186 373494
rect 113422 373258 113464 373494
rect 113144 366494 113464 373258
rect 113144 366258 113186 366494
rect 113422 366258 113464 366494
rect 113144 359494 113464 366258
rect 113144 359258 113186 359494
rect 113422 359258 113464 359494
rect 113144 352494 113464 359258
rect 113144 352258 113186 352494
rect 113422 352258 113464 352494
rect 113144 345494 113464 352258
rect 113144 345258 113186 345494
rect 113422 345258 113464 345494
rect 113144 338494 113464 345258
rect 113144 338258 113186 338494
rect 113422 338258 113464 338494
rect 113144 331494 113464 338258
rect 113144 331258 113186 331494
rect 113422 331258 113464 331494
rect 113144 324494 113464 331258
rect 113144 324258 113186 324494
rect 113422 324258 113464 324494
rect 113144 317494 113464 324258
rect 113144 317258 113186 317494
rect 113422 317258 113464 317494
rect 113144 310494 113464 317258
rect 113144 310258 113186 310494
rect 113422 310258 113464 310494
rect 113144 303494 113464 310258
rect 113144 303258 113186 303494
rect 113422 303258 113464 303494
rect 113144 296494 113464 303258
rect 113144 296258 113186 296494
rect 113422 296258 113464 296494
rect 113144 289494 113464 296258
rect 113144 289258 113186 289494
rect 113422 289258 113464 289494
rect 113144 282494 113464 289258
rect 113144 282258 113186 282494
rect 113422 282258 113464 282494
rect 113144 275494 113464 282258
rect 113144 275258 113186 275494
rect 113422 275258 113464 275494
rect 113144 268494 113464 275258
rect 113144 268258 113186 268494
rect 113422 268258 113464 268494
rect 113144 261494 113464 268258
rect 113144 261258 113186 261494
rect 113422 261258 113464 261494
rect 113144 254494 113464 261258
rect 113144 254258 113186 254494
rect 113422 254258 113464 254494
rect 113144 247494 113464 254258
rect 113144 247258 113186 247494
rect 113422 247258 113464 247494
rect 113144 240494 113464 247258
rect 113144 240258 113186 240494
rect 113422 240258 113464 240494
rect 113144 233494 113464 240258
rect 113144 233258 113186 233494
rect 113422 233258 113464 233494
rect 113144 226494 113464 233258
rect 113144 226258 113186 226494
rect 113422 226258 113464 226494
rect 113144 219494 113464 226258
rect 113144 219258 113186 219494
rect 113422 219258 113464 219494
rect 113144 212494 113464 219258
rect 113144 212258 113186 212494
rect 113422 212258 113464 212494
rect 113144 205494 113464 212258
rect 113144 205258 113186 205494
rect 113422 205258 113464 205494
rect 113144 198494 113464 205258
rect 113144 198258 113186 198494
rect 113422 198258 113464 198494
rect 113144 191494 113464 198258
rect 113144 191258 113186 191494
rect 113422 191258 113464 191494
rect 113144 184494 113464 191258
rect 113144 184258 113186 184494
rect 113422 184258 113464 184494
rect 113144 177494 113464 184258
rect 113144 177258 113186 177494
rect 113422 177258 113464 177494
rect 113144 170494 113464 177258
rect 113144 170258 113186 170494
rect 113422 170258 113464 170494
rect 113144 163494 113464 170258
rect 113144 163258 113186 163494
rect 113422 163258 113464 163494
rect 113144 156494 113464 163258
rect 113144 156258 113186 156494
rect 113422 156258 113464 156494
rect 113144 149494 113464 156258
rect 113144 149258 113186 149494
rect 113422 149258 113464 149494
rect 113144 142494 113464 149258
rect 113144 142258 113186 142494
rect 113422 142258 113464 142494
rect 113144 135494 113464 142258
rect 113144 135258 113186 135494
rect 113422 135258 113464 135494
rect 113144 128494 113464 135258
rect 113144 128258 113186 128494
rect 113422 128258 113464 128494
rect 113144 121494 113464 128258
rect 113144 121258 113186 121494
rect 113422 121258 113464 121494
rect 113144 114494 113464 121258
rect 113144 114258 113186 114494
rect 113422 114258 113464 114494
rect 113144 107494 113464 114258
rect 113144 107258 113186 107494
rect 113422 107258 113464 107494
rect 113144 100494 113464 107258
rect 113144 100258 113186 100494
rect 113422 100258 113464 100494
rect 113144 93494 113464 100258
rect 113144 93258 113186 93494
rect 113422 93258 113464 93494
rect 113144 86494 113464 93258
rect 113144 86258 113186 86494
rect 113422 86258 113464 86494
rect 113144 79494 113464 86258
rect 113144 79258 113186 79494
rect 113422 79258 113464 79494
rect 113144 72494 113464 79258
rect 113144 72258 113186 72494
rect 113422 72258 113464 72494
rect 113144 65494 113464 72258
rect 113144 65258 113186 65494
rect 113422 65258 113464 65494
rect 113144 58494 113464 65258
rect 113144 58258 113186 58494
rect 113422 58258 113464 58494
rect 113144 51494 113464 58258
rect 113144 51258 113186 51494
rect 113422 51258 113464 51494
rect 113144 44494 113464 51258
rect 113144 44258 113186 44494
rect 113422 44258 113464 44494
rect 113144 37494 113464 44258
rect 113144 37258 113186 37494
rect 113422 37258 113464 37494
rect 113144 30494 113464 37258
rect 113144 30258 113186 30494
rect 113422 30258 113464 30494
rect 113144 23494 113464 30258
rect 113144 23258 113186 23494
rect 113422 23258 113464 23494
rect 113144 16494 113464 23258
rect 113144 16258 113186 16494
rect 113422 16258 113464 16494
rect 113144 9494 113464 16258
rect 113144 9258 113186 9494
rect 113422 9258 113464 9494
rect 113144 2494 113464 9258
rect 113144 2258 113186 2494
rect 113422 2258 113464 2494
rect 113144 -746 113464 2258
rect 113144 -982 113186 -746
rect 113422 -982 113464 -746
rect 113144 -1066 113464 -982
rect 113144 -1302 113186 -1066
rect 113422 -1302 113464 -1066
rect 113144 -2294 113464 -1302
rect 114876 706198 115196 706230
rect 114876 705962 114918 706198
rect 115154 705962 115196 706198
rect 114876 705878 115196 705962
rect 114876 705642 114918 705878
rect 115154 705642 115196 705878
rect 114876 696561 115196 705642
rect 114876 696325 114918 696561
rect 115154 696325 115196 696561
rect 114876 689561 115196 696325
rect 114876 689325 114918 689561
rect 115154 689325 115196 689561
rect 114876 682561 115196 689325
rect 114876 682325 114918 682561
rect 115154 682325 115196 682561
rect 114876 675561 115196 682325
rect 114876 675325 114918 675561
rect 115154 675325 115196 675561
rect 114876 668561 115196 675325
rect 114876 668325 114918 668561
rect 115154 668325 115196 668561
rect 114876 661561 115196 668325
rect 114876 661325 114918 661561
rect 115154 661325 115196 661561
rect 114876 654561 115196 661325
rect 114876 654325 114918 654561
rect 115154 654325 115196 654561
rect 114876 647561 115196 654325
rect 114876 647325 114918 647561
rect 115154 647325 115196 647561
rect 114876 640561 115196 647325
rect 114876 640325 114918 640561
rect 115154 640325 115196 640561
rect 114876 633561 115196 640325
rect 114876 633325 114918 633561
rect 115154 633325 115196 633561
rect 114876 626561 115196 633325
rect 114876 626325 114918 626561
rect 115154 626325 115196 626561
rect 114876 619561 115196 626325
rect 114876 619325 114918 619561
rect 115154 619325 115196 619561
rect 114876 612561 115196 619325
rect 114876 612325 114918 612561
rect 115154 612325 115196 612561
rect 114876 605561 115196 612325
rect 114876 605325 114918 605561
rect 115154 605325 115196 605561
rect 114876 598561 115196 605325
rect 114876 598325 114918 598561
rect 115154 598325 115196 598561
rect 114876 591561 115196 598325
rect 114876 591325 114918 591561
rect 115154 591325 115196 591561
rect 114876 584561 115196 591325
rect 114876 584325 114918 584561
rect 115154 584325 115196 584561
rect 114876 577561 115196 584325
rect 114876 577325 114918 577561
rect 115154 577325 115196 577561
rect 114876 570561 115196 577325
rect 114876 570325 114918 570561
rect 115154 570325 115196 570561
rect 114876 563561 115196 570325
rect 114876 563325 114918 563561
rect 115154 563325 115196 563561
rect 114876 556561 115196 563325
rect 114876 556325 114918 556561
rect 115154 556325 115196 556561
rect 114876 549561 115196 556325
rect 114876 549325 114918 549561
rect 115154 549325 115196 549561
rect 114876 542561 115196 549325
rect 114876 542325 114918 542561
rect 115154 542325 115196 542561
rect 114876 535561 115196 542325
rect 114876 535325 114918 535561
rect 115154 535325 115196 535561
rect 114876 528561 115196 535325
rect 114876 528325 114918 528561
rect 115154 528325 115196 528561
rect 114876 521561 115196 528325
rect 114876 521325 114918 521561
rect 115154 521325 115196 521561
rect 114876 514561 115196 521325
rect 114876 514325 114918 514561
rect 115154 514325 115196 514561
rect 114876 507561 115196 514325
rect 114876 507325 114918 507561
rect 115154 507325 115196 507561
rect 114876 500561 115196 507325
rect 114876 500325 114918 500561
rect 115154 500325 115196 500561
rect 114876 493561 115196 500325
rect 114876 493325 114918 493561
rect 115154 493325 115196 493561
rect 114876 486561 115196 493325
rect 114876 486325 114918 486561
rect 115154 486325 115196 486561
rect 114876 479561 115196 486325
rect 114876 479325 114918 479561
rect 115154 479325 115196 479561
rect 114876 472561 115196 479325
rect 114876 472325 114918 472561
rect 115154 472325 115196 472561
rect 114876 465561 115196 472325
rect 114876 465325 114918 465561
rect 115154 465325 115196 465561
rect 114876 458561 115196 465325
rect 114876 458325 114918 458561
rect 115154 458325 115196 458561
rect 114876 451561 115196 458325
rect 114876 451325 114918 451561
rect 115154 451325 115196 451561
rect 114876 444561 115196 451325
rect 114876 444325 114918 444561
rect 115154 444325 115196 444561
rect 114876 437561 115196 444325
rect 114876 437325 114918 437561
rect 115154 437325 115196 437561
rect 114876 430561 115196 437325
rect 114876 430325 114918 430561
rect 115154 430325 115196 430561
rect 114876 423561 115196 430325
rect 114876 423325 114918 423561
rect 115154 423325 115196 423561
rect 114876 416561 115196 423325
rect 114876 416325 114918 416561
rect 115154 416325 115196 416561
rect 114876 409561 115196 416325
rect 114876 409325 114918 409561
rect 115154 409325 115196 409561
rect 114876 402561 115196 409325
rect 114876 402325 114918 402561
rect 115154 402325 115196 402561
rect 114876 395561 115196 402325
rect 114876 395325 114918 395561
rect 115154 395325 115196 395561
rect 114876 388561 115196 395325
rect 114876 388325 114918 388561
rect 115154 388325 115196 388561
rect 114876 381561 115196 388325
rect 114876 381325 114918 381561
rect 115154 381325 115196 381561
rect 114876 374561 115196 381325
rect 114876 374325 114918 374561
rect 115154 374325 115196 374561
rect 114876 367561 115196 374325
rect 114876 367325 114918 367561
rect 115154 367325 115196 367561
rect 114876 360561 115196 367325
rect 114876 360325 114918 360561
rect 115154 360325 115196 360561
rect 114876 353561 115196 360325
rect 114876 353325 114918 353561
rect 115154 353325 115196 353561
rect 114876 346561 115196 353325
rect 114876 346325 114918 346561
rect 115154 346325 115196 346561
rect 114876 339561 115196 346325
rect 114876 339325 114918 339561
rect 115154 339325 115196 339561
rect 114876 332561 115196 339325
rect 114876 332325 114918 332561
rect 115154 332325 115196 332561
rect 114876 325561 115196 332325
rect 114876 325325 114918 325561
rect 115154 325325 115196 325561
rect 114876 318561 115196 325325
rect 114876 318325 114918 318561
rect 115154 318325 115196 318561
rect 114876 311561 115196 318325
rect 114876 311325 114918 311561
rect 115154 311325 115196 311561
rect 114876 304561 115196 311325
rect 114876 304325 114918 304561
rect 115154 304325 115196 304561
rect 114876 297561 115196 304325
rect 114876 297325 114918 297561
rect 115154 297325 115196 297561
rect 114876 290561 115196 297325
rect 114876 290325 114918 290561
rect 115154 290325 115196 290561
rect 114876 283561 115196 290325
rect 114876 283325 114918 283561
rect 115154 283325 115196 283561
rect 114876 276561 115196 283325
rect 114876 276325 114918 276561
rect 115154 276325 115196 276561
rect 114876 269561 115196 276325
rect 114876 269325 114918 269561
rect 115154 269325 115196 269561
rect 114876 262561 115196 269325
rect 114876 262325 114918 262561
rect 115154 262325 115196 262561
rect 114876 255561 115196 262325
rect 114876 255325 114918 255561
rect 115154 255325 115196 255561
rect 114876 248561 115196 255325
rect 114876 248325 114918 248561
rect 115154 248325 115196 248561
rect 114876 241561 115196 248325
rect 114876 241325 114918 241561
rect 115154 241325 115196 241561
rect 114876 234561 115196 241325
rect 114876 234325 114918 234561
rect 115154 234325 115196 234561
rect 114876 227561 115196 234325
rect 114876 227325 114918 227561
rect 115154 227325 115196 227561
rect 114876 220561 115196 227325
rect 114876 220325 114918 220561
rect 115154 220325 115196 220561
rect 114876 213561 115196 220325
rect 114876 213325 114918 213561
rect 115154 213325 115196 213561
rect 114876 206561 115196 213325
rect 114876 206325 114918 206561
rect 115154 206325 115196 206561
rect 114876 199561 115196 206325
rect 114876 199325 114918 199561
rect 115154 199325 115196 199561
rect 114876 192561 115196 199325
rect 114876 192325 114918 192561
rect 115154 192325 115196 192561
rect 114876 185561 115196 192325
rect 114876 185325 114918 185561
rect 115154 185325 115196 185561
rect 114876 178561 115196 185325
rect 114876 178325 114918 178561
rect 115154 178325 115196 178561
rect 114876 171561 115196 178325
rect 114876 171325 114918 171561
rect 115154 171325 115196 171561
rect 114876 164561 115196 171325
rect 114876 164325 114918 164561
rect 115154 164325 115196 164561
rect 114876 157561 115196 164325
rect 114876 157325 114918 157561
rect 115154 157325 115196 157561
rect 114876 150561 115196 157325
rect 114876 150325 114918 150561
rect 115154 150325 115196 150561
rect 114876 143561 115196 150325
rect 114876 143325 114918 143561
rect 115154 143325 115196 143561
rect 114876 136561 115196 143325
rect 114876 136325 114918 136561
rect 115154 136325 115196 136561
rect 114876 129561 115196 136325
rect 114876 129325 114918 129561
rect 115154 129325 115196 129561
rect 114876 122561 115196 129325
rect 114876 122325 114918 122561
rect 115154 122325 115196 122561
rect 114876 115561 115196 122325
rect 114876 115325 114918 115561
rect 115154 115325 115196 115561
rect 114876 108561 115196 115325
rect 114876 108325 114918 108561
rect 115154 108325 115196 108561
rect 114876 101561 115196 108325
rect 114876 101325 114918 101561
rect 115154 101325 115196 101561
rect 114876 94561 115196 101325
rect 114876 94325 114918 94561
rect 115154 94325 115196 94561
rect 114876 87561 115196 94325
rect 114876 87325 114918 87561
rect 115154 87325 115196 87561
rect 114876 80561 115196 87325
rect 114876 80325 114918 80561
rect 115154 80325 115196 80561
rect 114876 73561 115196 80325
rect 114876 73325 114918 73561
rect 115154 73325 115196 73561
rect 114876 66561 115196 73325
rect 114876 66325 114918 66561
rect 115154 66325 115196 66561
rect 114876 59561 115196 66325
rect 114876 59325 114918 59561
rect 115154 59325 115196 59561
rect 114876 52561 115196 59325
rect 114876 52325 114918 52561
rect 115154 52325 115196 52561
rect 114876 45561 115196 52325
rect 114876 45325 114918 45561
rect 115154 45325 115196 45561
rect 114876 38561 115196 45325
rect 114876 38325 114918 38561
rect 115154 38325 115196 38561
rect 114876 31561 115196 38325
rect 114876 31325 114918 31561
rect 115154 31325 115196 31561
rect 114876 24561 115196 31325
rect 114876 24325 114918 24561
rect 115154 24325 115196 24561
rect 114876 17561 115196 24325
rect 114876 17325 114918 17561
rect 115154 17325 115196 17561
rect 114876 10561 115196 17325
rect 114876 10325 114918 10561
rect 115154 10325 115196 10561
rect 114876 3561 115196 10325
rect 114876 3325 114918 3561
rect 115154 3325 115196 3561
rect 114876 -1706 115196 3325
rect 114876 -1942 114918 -1706
rect 115154 -1942 115196 -1706
rect 114876 -2026 115196 -1942
rect 114876 -2262 114918 -2026
rect 115154 -2262 115196 -2026
rect 114876 -2294 115196 -2262
rect 120144 705238 120464 706230
rect 120144 705002 120186 705238
rect 120422 705002 120464 705238
rect 120144 704918 120464 705002
rect 120144 704682 120186 704918
rect 120422 704682 120464 704918
rect 120144 695494 120464 704682
rect 120144 695258 120186 695494
rect 120422 695258 120464 695494
rect 120144 688494 120464 695258
rect 120144 688258 120186 688494
rect 120422 688258 120464 688494
rect 120144 681494 120464 688258
rect 120144 681258 120186 681494
rect 120422 681258 120464 681494
rect 120144 674494 120464 681258
rect 120144 674258 120186 674494
rect 120422 674258 120464 674494
rect 120144 667494 120464 674258
rect 120144 667258 120186 667494
rect 120422 667258 120464 667494
rect 120144 660494 120464 667258
rect 120144 660258 120186 660494
rect 120422 660258 120464 660494
rect 120144 653494 120464 660258
rect 120144 653258 120186 653494
rect 120422 653258 120464 653494
rect 120144 646494 120464 653258
rect 120144 646258 120186 646494
rect 120422 646258 120464 646494
rect 120144 639494 120464 646258
rect 120144 639258 120186 639494
rect 120422 639258 120464 639494
rect 120144 632494 120464 639258
rect 120144 632258 120186 632494
rect 120422 632258 120464 632494
rect 120144 625494 120464 632258
rect 120144 625258 120186 625494
rect 120422 625258 120464 625494
rect 120144 618494 120464 625258
rect 120144 618258 120186 618494
rect 120422 618258 120464 618494
rect 120144 611494 120464 618258
rect 120144 611258 120186 611494
rect 120422 611258 120464 611494
rect 120144 604494 120464 611258
rect 120144 604258 120186 604494
rect 120422 604258 120464 604494
rect 120144 597494 120464 604258
rect 120144 597258 120186 597494
rect 120422 597258 120464 597494
rect 120144 590494 120464 597258
rect 120144 590258 120186 590494
rect 120422 590258 120464 590494
rect 120144 583494 120464 590258
rect 120144 583258 120186 583494
rect 120422 583258 120464 583494
rect 120144 576494 120464 583258
rect 120144 576258 120186 576494
rect 120422 576258 120464 576494
rect 120144 569494 120464 576258
rect 120144 569258 120186 569494
rect 120422 569258 120464 569494
rect 120144 562494 120464 569258
rect 120144 562258 120186 562494
rect 120422 562258 120464 562494
rect 120144 555494 120464 562258
rect 120144 555258 120186 555494
rect 120422 555258 120464 555494
rect 120144 548494 120464 555258
rect 120144 548258 120186 548494
rect 120422 548258 120464 548494
rect 120144 541494 120464 548258
rect 120144 541258 120186 541494
rect 120422 541258 120464 541494
rect 120144 534494 120464 541258
rect 120144 534258 120186 534494
rect 120422 534258 120464 534494
rect 120144 527494 120464 534258
rect 120144 527258 120186 527494
rect 120422 527258 120464 527494
rect 120144 520494 120464 527258
rect 120144 520258 120186 520494
rect 120422 520258 120464 520494
rect 120144 513494 120464 520258
rect 120144 513258 120186 513494
rect 120422 513258 120464 513494
rect 120144 506494 120464 513258
rect 120144 506258 120186 506494
rect 120422 506258 120464 506494
rect 120144 499494 120464 506258
rect 120144 499258 120186 499494
rect 120422 499258 120464 499494
rect 120144 492494 120464 499258
rect 120144 492258 120186 492494
rect 120422 492258 120464 492494
rect 120144 485494 120464 492258
rect 120144 485258 120186 485494
rect 120422 485258 120464 485494
rect 120144 478494 120464 485258
rect 120144 478258 120186 478494
rect 120422 478258 120464 478494
rect 120144 471494 120464 478258
rect 120144 471258 120186 471494
rect 120422 471258 120464 471494
rect 120144 464494 120464 471258
rect 120144 464258 120186 464494
rect 120422 464258 120464 464494
rect 120144 457494 120464 464258
rect 120144 457258 120186 457494
rect 120422 457258 120464 457494
rect 120144 450494 120464 457258
rect 120144 450258 120186 450494
rect 120422 450258 120464 450494
rect 120144 443494 120464 450258
rect 120144 443258 120186 443494
rect 120422 443258 120464 443494
rect 120144 436494 120464 443258
rect 120144 436258 120186 436494
rect 120422 436258 120464 436494
rect 120144 429494 120464 436258
rect 120144 429258 120186 429494
rect 120422 429258 120464 429494
rect 120144 422494 120464 429258
rect 120144 422258 120186 422494
rect 120422 422258 120464 422494
rect 120144 415494 120464 422258
rect 120144 415258 120186 415494
rect 120422 415258 120464 415494
rect 120144 408494 120464 415258
rect 120144 408258 120186 408494
rect 120422 408258 120464 408494
rect 120144 401494 120464 408258
rect 120144 401258 120186 401494
rect 120422 401258 120464 401494
rect 120144 394494 120464 401258
rect 120144 394258 120186 394494
rect 120422 394258 120464 394494
rect 120144 387494 120464 394258
rect 120144 387258 120186 387494
rect 120422 387258 120464 387494
rect 120144 380494 120464 387258
rect 120144 380258 120186 380494
rect 120422 380258 120464 380494
rect 120144 373494 120464 380258
rect 120144 373258 120186 373494
rect 120422 373258 120464 373494
rect 120144 366494 120464 373258
rect 120144 366258 120186 366494
rect 120422 366258 120464 366494
rect 120144 359494 120464 366258
rect 120144 359258 120186 359494
rect 120422 359258 120464 359494
rect 120144 352494 120464 359258
rect 120144 352258 120186 352494
rect 120422 352258 120464 352494
rect 120144 345494 120464 352258
rect 120144 345258 120186 345494
rect 120422 345258 120464 345494
rect 120144 338494 120464 345258
rect 120144 338258 120186 338494
rect 120422 338258 120464 338494
rect 120144 331494 120464 338258
rect 120144 331258 120186 331494
rect 120422 331258 120464 331494
rect 120144 324494 120464 331258
rect 120144 324258 120186 324494
rect 120422 324258 120464 324494
rect 120144 317494 120464 324258
rect 120144 317258 120186 317494
rect 120422 317258 120464 317494
rect 120144 310494 120464 317258
rect 120144 310258 120186 310494
rect 120422 310258 120464 310494
rect 120144 303494 120464 310258
rect 120144 303258 120186 303494
rect 120422 303258 120464 303494
rect 120144 296494 120464 303258
rect 120144 296258 120186 296494
rect 120422 296258 120464 296494
rect 120144 289494 120464 296258
rect 120144 289258 120186 289494
rect 120422 289258 120464 289494
rect 120144 282494 120464 289258
rect 120144 282258 120186 282494
rect 120422 282258 120464 282494
rect 120144 275494 120464 282258
rect 120144 275258 120186 275494
rect 120422 275258 120464 275494
rect 120144 268494 120464 275258
rect 120144 268258 120186 268494
rect 120422 268258 120464 268494
rect 120144 261494 120464 268258
rect 120144 261258 120186 261494
rect 120422 261258 120464 261494
rect 120144 254494 120464 261258
rect 120144 254258 120186 254494
rect 120422 254258 120464 254494
rect 120144 247494 120464 254258
rect 120144 247258 120186 247494
rect 120422 247258 120464 247494
rect 120144 240494 120464 247258
rect 120144 240258 120186 240494
rect 120422 240258 120464 240494
rect 120144 233494 120464 240258
rect 120144 233258 120186 233494
rect 120422 233258 120464 233494
rect 120144 226494 120464 233258
rect 120144 226258 120186 226494
rect 120422 226258 120464 226494
rect 120144 219494 120464 226258
rect 120144 219258 120186 219494
rect 120422 219258 120464 219494
rect 120144 212494 120464 219258
rect 120144 212258 120186 212494
rect 120422 212258 120464 212494
rect 120144 205494 120464 212258
rect 120144 205258 120186 205494
rect 120422 205258 120464 205494
rect 120144 198494 120464 205258
rect 120144 198258 120186 198494
rect 120422 198258 120464 198494
rect 120144 191494 120464 198258
rect 120144 191258 120186 191494
rect 120422 191258 120464 191494
rect 120144 184494 120464 191258
rect 120144 184258 120186 184494
rect 120422 184258 120464 184494
rect 120144 177494 120464 184258
rect 120144 177258 120186 177494
rect 120422 177258 120464 177494
rect 120144 170494 120464 177258
rect 120144 170258 120186 170494
rect 120422 170258 120464 170494
rect 120144 163494 120464 170258
rect 120144 163258 120186 163494
rect 120422 163258 120464 163494
rect 120144 156494 120464 163258
rect 120144 156258 120186 156494
rect 120422 156258 120464 156494
rect 120144 149494 120464 156258
rect 120144 149258 120186 149494
rect 120422 149258 120464 149494
rect 120144 142494 120464 149258
rect 120144 142258 120186 142494
rect 120422 142258 120464 142494
rect 120144 135494 120464 142258
rect 120144 135258 120186 135494
rect 120422 135258 120464 135494
rect 120144 128494 120464 135258
rect 120144 128258 120186 128494
rect 120422 128258 120464 128494
rect 120144 121494 120464 128258
rect 120144 121258 120186 121494
rect 120422 121258 120464 121494
rect 120144 114494 120464 121258
rect 120144 114258 120186 114494
rect 120422 114258 120464 114494
rect 120144 107494 120464 114258
rect 120144 107258 120186 107494
rect 120422 107258 120464 107494
rect 120144 100494 120464 107258
rect 120144 100258 120186 100494
rect 120422 100258 120464 100494
rect 120144 93494 120464 100258
rect 120144 93258 120186 93494
rect 120422 93258 120464 93494
rect 120144 86494 120464 93258
rect 120144 86258 120186 86494
rect 120422 86258 120464 86494
rect 120144 79494 120464 86258
rect 120144 79258 120186 79494
rect 120422 79258 120464 79494
rect 120144 72494 120464 79258
rect 120144 72258 120186 72494
rect 120422 72258 120464 72494
rect 120144 65494 120464 72258
rect 120144 65258 120186 65494
rect 120422 65258 120464 65494
rect 120144 58494 120464 65258
rect 120144 58258 120186 58494
rect 120422 58258 120464 58494
rect 120144 51494 120464 58258
rect 120144 51258 120186 51494
rect 120422 51258 120464 51494
rect 120144 44494 120464 51258
rect 120144 44258 120186 44494
rect 120422 44258 120464 44494
rect 120144 37494 120464 44258
rect 120144 37258 120186 37494
rect 120422 37258 120464 37494
rect 120144 30494 120464 37258
rect 120144 30258 120186 30494
rect 120422 30258 120464 30494
rect 120144 23494 120464 30258
rect 120144 23258 120186 23494
rect 120422 23258 120464 23494
rect 120144 16494 120464 23258
rect 120144 16258 120186 16494
rect 120422 16258 120464 16494
rect 120144 9494 120464 16258
rect 120144 9258 120186 9494
rect 120422 9258 120464 9494
rect 120144 2494 120464 9258
rect 120144 2258 120186 2494
rect 120422 2258 120464 2494
rect 120144 -746 120464 2258
rect 120144 -982 120186 -746
rect 120422 -982 120464 -746
rect 120144 -1066 120464 -982
rect 120144 -1302 120186 -1066
rect 120422 -1302 120464 -1066
rect 120144 -2294 120464 -1302
rect 121876 706198 122196 706230
rect 121876 705962 121918 706198
rect 122154 705962 122196 706198
rect 121876 705878 122196 705962
rect 121876 705642 121918 705878
rect 122154 705642 122196 705878
rect 121876 696561 122196 705642
rect 121876 696325 121918 696561
rect 122154 696325 122196 696561
rect 121876 689561 122196 696325
rect 121876 689325 121918 689561
rect 122154 689325 122196 689561
rect 121876 682561 122196 689325
rect 121876 682325 121918 682561
rect 122154 682325 122196 682561
rect 121876 675561 122196 682325
rect 121876 675325 121918 675561
rect 122154 675325 122196 675561
rect 121876 668561 122196 675325
rect 121876 668325 121918 668561
rect 122154 668325 122196 668561
rect 121876 661561 122196 668325
rect 121876 661325 121918 661561
rect 122154 661325 122196 661561
rect 121876 654561 122196 661325
rect 121876 654325 121918 654561
rect 122154 654325 122196 654561
rect 121876 647561 122196 654325
rect 121876 647325 121918 647561
rect 122154 647325 122196 647561
rect 121876 640561 122196 647325
rect 121876 640325 121918 640561
rect 122154 640325 122196 640561
rect 121876 633561 122196 640325
rect 121876 633325 121918 633561
rect 122154 633325 122196 633561
rect 121876 626561 122196 633325
rect 121876 626325 121918 626561
rect 122154 626325 122196 626561
rect 121876 619561 122196 626325
rect 121876 619325 121918 619561
rect 122154 619325 122196 619561
rect 121876 612561 122196 619325
rect 121876 612325 121918 612561
rect 122154 612325 122196 612561
rect 121876 605561 122196 612325
rect 121876 605325 121918 605561
rect 122154 605325 122196 605561
rect 121876 598561 122196 605325
rect 121876 598325 121918 598561
rect 122154 598325 122196 598561
rect 121876 591561 122196 598325
rect 121876 591325 121918 591561
rect 122154 591325 122196 591561
rect 121876 584561 122196 591325
rect 121876 584325 121918 584561
rect 122154 584325 122196 584561
rect 121876 577561 122196 584325
rect 121876 577325 121918 577561
rect 122154 577325 122196 577561
rect 121876 570561 122196 577325
rect 121876 570325 121918 570561
rect 122154 570325 122196 570561
rect 121876 563561 122196 570325
rect 121876 563325 121918 563561
rect 122154 563325 122196 563561
rect 121876 556561 122196 563325
rect 121876 556325 121918 556561
rect 122154 556325 122196 556561
rect 121876 549561 122196 556325
rect 121876 549325 121918 549561
rect 122154 549325 122196 549561
rect 121876 542561 122196 549325
rect 121876 542325 121918 542561
rect 122154 542325 122196 542561
rect 121876 535561 122196 542325
rect 121876 535325 121918 535561
rect 122154 535325 122196 535561
rect 121876 528561 122196 535325
rect 121876 528325 121918 528561
rect 122154 528325 122196 528561
rect 121876 521561 122196 528325
rect 121876 521325 121918 521561
rect 122154 521325 122196 521561
rect 121876 514561 122196 521325
rect 121876 514325 121918 514561
rect 122154 514325 122196 514561
rect 121876 507561 122196 514325
rect 121876 507325 121918 507561
rect 122154 507325 122196 507561
rect 121876 500561 122196 507325
rect 121876 500325 121918 500561
rect 122154 500325 122196 500561
rect 121876 493561 122196 500325
rect 121876 493325 121918 493561
rect 122154 493325 122196 493561
rect 121876 486561 122196 493325
rect 121876 486325 121918 486561
rect 122154 486325 122196 486561
rect 121876 479561 122196 486325
rect 121876 479325 121918 479561
rect 122154 479325 122196 479561
rect 121876 472561 122196 479325
rect 121876 472325 121918 472561
rect 122154 472325 122196 472561
rect 121876 465561 122196 472325
rect 121876 465325 121918 465561
rect 122154 465325 122196 465561
rect 121876 458561 122196 465325
rect 121876 458325 121918 458561
rect 122154 458325 122196 458561
rect 121876 451561 122196 458325
rect 121876 451325 121918 451561
rect 122154 451325 122196 451561
rect 121876 444561 122196 451325
rect 121876 444325 121918 444561
rect 122154 444325 122196 444561
rect 121876 437561 122196 444325
rect 121876 437325 121918 437561
rect 122154 437325 122196 437561
rect 121876 430561 122196 437325
rect 121876 430325 121918 430561
rect 122154 430325 122196 430561
rect 121876 423561 122196 430325
rect 121876 423325 121918 423561
rect 122154 423325 122196 423561
rect 121876 416561 122196 423325
rect 121876 416325 121918 416561
rect 122154 416325 122196 416561
rect 121876 409561 122196 416325
rect 121876 409325 121918 409561
rect 122154 409325 122196 409561
rect 121876 402561 122196 409325
rect 121876 402325 121918 402561
rect 122154 402325 122196 402561
rect 121876 395561 122196 402325
rect 121876 395325 121918 395561
rect 122154 395325 122196 395561
rect 121876 388561 122196 395325
rect 121876 388325 121918 388561
rect 122154 388325 122196 388561
rect 121876 381561 122196 388325
rect 121876 381325 121918 381561
rect 122154 381325 122196 381561
rect 121876 374561 122196 381325
rect 121876 374325 121918 374561
rect 122154 374325 122196 374561
rect 121876 367561 122196 374325
rect 121876 367325 121918 367561
rect 122154 367325 122196 367561
rect 121876 360561 122196 367325
rect 121876 360325 121918 360561
rect 122154 360325 122196 360561
rect 121876 353561 122196 360325
rect 121876 353325 121918 353561
rect 122154 353325 122196 353561
rect 121876 346561 122196 353325
rect 121876 346325 121918 346561
rect 122154 346325 122196 346561
rect 121876 339561 122196 346325
rect 121876 339325 121918 339561
rect 122154 339325 122196 339561
rect 121876 332561 122196 339325
rect 121876 332325 121918 332561
rect 122154 332325 122196 332561
rect 121876 325561 122196 332325
rect 121876 325325 121918 325561
rect 122154 325325 122196 325561
rect 121876 318561 122196 325325
rect 121876 318325 121918 318561
rect 122154 318325 122196 318561
rect 121876 311561 122196 318325
rect 121876 311325 121918 311561
rect 122154 311325 122196 311561
rect 121876 304561 122196 311325
rect 121876 304325 121918 304561
rect 122154 304325 122196 304561
rect 121876 297561 122196 304325
rect 121876 297325 121918 297561
rect 122154 297325 122196 297561
rect 121876 290561 122196 297325
rect 121876 290325 121918 290561
rect 122154 290325 122196 290561
rect 121876 283561 122196 290325
rect 121876 283325 121918 283561
rect 122154 283325 122196 283561
rect 121876 276561 122196 283325
rect 121876 276325 121918 276561
rect 122154 276325 122196 276561
rect 121876 269561 122196 276325
rect 121876 269325 121918 269561
rect 122154 269325 122196 269561
rect 121876 262561 122196 269325
rect 121876 262325 121918 262561
rect 122154 262325 122196 262561
rect 121876 255561 122196 262325
rect 121876 255325 121918 255561
rect 122154 255325 122196 255561
rect 121876 248561 122196 255325
rect 121876 248325 121918 248561
rect 122154 248325 122196 248561
rect 121876 241561 122196 248325
rect 121876 241325 121918 241561
rect 122154 241325 122196 241561
rect 121876 234561 122196 241325
rect 121876 234325 121918 234561
rect 122154 234325 122196 234561
rect 121876 227561 122196 234325
rect 121876 227325 121918 227561
rect 122154 227325 122196 227561
rect 121876 220561 122196 227325
rect 121876 220325 121918 220561
rect 122154 220325 122196 220561
rect 121876 213561 122196 220325
rect 121876 213325 121918 213561
rect 122154 213325 122196 213561
rect 121876 206561 122196 213325
rect 121876 206325 121918 206561
rect 122154 206325 122196 206561
rect 121876 199561 122196 206325
rect 121876 199325 121918 199561
rect 122154 199325 122196 199561
rect 121876 192561 122196 199325
rect 121876 192325 121918 192561
rect 122154 192325 122196 192561
rect 121876 185561 122196 192325
rect 121876 185325 121918 185561
rect 122154 185325 122196 185561
rect 121876 178561 122196 185325
rect 121876 178325 121918 178561
rect 122154 178325 122196 178561
rect 121876 171561 122196 178325
rect 121876 171325 121918 171561
rect 122154 171325 122196 171561
rect 121876 164561 122196 171325
rect 121876 164325 121918 164561
rect 122154 164325 122196 164561
rect 121876 157561 122196 164325
rect 121876 157325 121918 157561
rect 122154 157325 122196 157561
rect 121876 150561 122196 157325
rect 121876 150325 121918 150561
rect 122154 150325 122196 150561
rect 121876 143561 122196 150325
rect 121876 143325 121918 143561
rect 122154 143325 122196 143561
rect 121876 136561 122196 143325
rect 121876 136325 121918 136561
rect 122154 136325 122196 136561
rect 121876 129561 122196 136325
rect 121876 129325 121918 129561
rect 122154 129325 122196 129561
rect 121876 122561 122196 129325
rect 121876 122325 121918 122561
rect 122154 122325 122196 122561
rect 121876 115561 122196 122325
rect 121876 115325 121918 115561
rect 122154 115325 122196 115561
rect 121876 108561 122196 115325
rect 121876 108325 121918 108561
rect 122154 108325 122196 108561
rect 121876 101561 122196 108325
rect 121876 101325 121918 101561
rect 122154 101325 122196 101561
rect 121876 94561 122196 101325
rect 121876 94325 121918 94561
rect 122154 94325 122196 94561
rect 121876 87561 122196 94325
rect 121876 87325 121918 87561
rect 122154 87325 122196 87561
rect 121876 80561 122196 87325
rect 121876 80325 121918 80561
rect 122154 80325 122196 80561
rect 121876 73561 122196 80325
rect 121876 73325 121918 73561
rect 122154 73325 122196 73561
rect 121876 66561 122196 73325
rect 121876 66325 121918 66561
rect 122154 66325 122196 66561
rect 121876 59561 122196 66325
rect 121876 59325 121918 59561
rect 122154 59325 122196 59561
rect 121876 52561 122196 59325
rect 121876 52325 121918 52561
rect 122154 52325 122196 52561
rect 121876 45561 122196 52325
rect 121876 45325 121918 45561
rect 122154 45325 122196 45561
rect 121876 38561 122196 45325
rect 121876 38325 121918 38561
rect 122154 38325 122196 38561
rect 121876 31561 122196 38325
rect 121876 31325 121918 31561
rect 122154 31325 122196 31561
rect 121876 24561 122196 31325
rect 121876 24325 121918 24561
rect 122154 24325 122196 24561
rect 121876 17561 122196 24325
rect 121876 17325 121918 17561
rect 122154 17325 122196 17561
rect 121876 10561 122196 17325
rect 121876 10325 121918 10561
rect 122154 10325 122196 10561
rect 121876 3561 122196 10325
rect 121876 3325 121918 3561
rect 122154 3325 122196 3561
rect 121876 -1706 122196 3325
rect 121876 -1942 121918 -1706
rect 122154 -1942 122196 -1706
rect 121876 -2026 122196 -1942
rect 121876 -2262 121918 -2026
rect 122154 -2262 122196 -2026
rect 121876 -2294 122196 -2262
rect 127144 705238 127464 706230
rect 127144 705002 127186 705238
rect 127422 705002 127464 705238
rect 127144 704918 127464 705002
rect 127144 704682 127186 704918
rect 127422 704682 127464 704918
rect 127144 695494 127464 704682
rect 127144 695258 127186 695494
rect 127422 695258 127464 695494
rect 127144 688494 127464 695258
rect 127144 688258 127186 688494
rect 127422 688258 127464 688494
rect 127144 681494 127464 688258
rect 127144 681258 127186 681494
rect 127422 681258 127464 681494
rect 127144 674494 127464 681258
rect 127144 674258 127186 674494
rect 127422 674258 127464 674494
rect 127144 667494 127464 674258
rect 127144 667258 127186 667494
rect 127422 667258 127464 667494
rect 127144 660494 127464 667258
rect 127144 660258 127186 660494
rect 127422 660258 127464 660494
rect 127144 653494 127464 660258
rect 127144 653258 127186 653494
rect 127422 653258 127464 653494
rect 127144 646494 127464 653258
rect 127144 646258 127186 646494
rect 127422 646258 127464 646494
rect 127144 639494 127464 646258
rect 127144 639258 127186 639494
rect 127422 639258 127464 639494
rect 127144 632494 127464 639258
rect 127144 632258 127186 632494
rect 127422 632258 127464 632494
rect 127144 625494 127464 632258
rect 127144 625258 127186 625494
rect 127422 625258 127464 625494
rect 127144 618494 127464 625258
rect 127144 618258 127186 618494
rect 127422 618258 127464 618494
rect 127144 611494 127464 618258
rect 127144 611258 127186 611494
rect 127422 611258 127464 611494
rect 127144 604494 127464 611258
rect 127144 604258 127186 604494
rect 127422 604258 127464 604494
rect 127144 597494 127464 604258
rect 127144 597258 127186 597494
rect 127422 597258 127464 597494
rect 127144 590494 127464 597258
rect 127144 590258 127186 590494
rect 127422 590258 127464 590494
rect 127144 583494 127464 590258
rect 127144 583258 127186 583494
rect 127422 583258 127464 583494
rect 127144 576494 127464 583258
rect 127144 576258 127186 576494
rect 127422 576258 127464 576494
rect 127144 569494 127464 576258
rect 127144 569258 127186 569494
rect 127422 569258 127464 569494
rect 127144 562494 127464 569258
rect 127144 562258 127186 562494
rect 127422 562258 127464 562494
rect 127144 555494 127464 562258
rect 127144 555258 127186 555494
rect 127422 555258 127464 555494
rect 127144 548494 127464 555258
rect 127144 548258 127186 548494
rect 127422 548258 127464 548494
rect 127144 541494 127464 548258
rect 127144 541258 127186 541494
rect 127422 541258 127464 541494
rect 127144 534494 127464 541258
rect 127144 534258 127186 534494
rect 127422 534258 127464 534494
rect 127144 527494 127464 534258
rect 127144 527258 127186 527494
rect 127422 527258 127464 527494
rect 127144 520494 127464 527258
rect 127144 520258 127186 520494
rect 127422 520258 127464 520494
rect 127144 513494 127464 520258
rect 127144 513258 127186 513494
rect 127422 513258 127464 513494
rect 127144 506494 127464 513258
rect 127144 506258 127186 506494
rect 127422 506258 127464 506494
rect 127144 499494 127464 506258
rect 127144 499258 127186 499494
rect 127422 499258 127464 499494
rect 127144 492494 127464 499258
rect 127144 492258 127186 492494
rect 127422 492258 127464 492494
rect 127144 485494 127464 492258
rect 127144 485258 127186 485494
rect 127422 485258 127464 485494
rect 127144 478494 127464 485258
rect 127144 478258 127186 478494
rect 127422 478258 127464 478494
rect 127144 471494 127464 478258
rect 127144 471258 127186 471494
rect 127422 471258 127464 471494
rect 127144 464494 127464 471258
rect 127144 464258 127186 464494
rect 127422 464258 127464 464494
rect 127144 457494 127464 464258
rect 127144 457258 127186 457494
rect 127422 457258 127464 457494
rect 127144 450494 127464 457258
rect 127144 450258 127186 450494
rect 127422 450258 127464 450494
rect 127144 443494 127464 450258
rect 127144 443258 127186 443494
rect 127422 443258 127464 443494
rect 127144 436494 127464 443258
rect 127144 436258 127186 436494
rect 127422 436258 127464 436494
rect 127144 429494 127464 436258
rect 127144 429258 127186 429494
rect 127422 429258 127464 429494
rect 127144 422494 127464 429258
rect 127144 422258 127186 422494
rect 127422 422258 127464 422494
rect 127144 415494 127464 422258
rect 127144 415258 127186 415494
rect 127422 415258 127464 415494
rect 127144 408494 127464 415258
rect 127144 408258 127186 408494
rect 127422 408258 127464 408494
rect 127144 401494 127464 408258
rect 127144 401258 127186 401494
rect 127422 401258 127464 401494
rect 127144 394494 127464 401258
rect 127144 394258 127186 394494
rect 127422 394258 127464 394494
rect 127144 387494 127464 394258
rect 127144 387258 127186 387494
rect 127422 387258 127464 387494
rect 127144 380494 127464 387258
rect 127144 380258 127186 380494
rect 127422 380258 127464 380494
rect 127144 373494 127464 380258
rect 127144 373258 127186 373494
rect 127422 373258 127464 373494
rect 127144 366494 127464 373258
rect 127144 366258 127186 366494
rect 127422 366258 127464 366494
rect 127144 359494 127464 366258
rect 127144 359258 127186 359494
rect 127422 359258 127464 359494
rect 127144 352494 127464 359258
rect 127144 352258 127186 352494
rect 127422 352258 127464 352494
rect 127144 345494 127464 352258
rect 127144 345258 127186 345494
rect 127422 345258 127464 345494
rect 127144 338494 127464 345258
rect 127144 338258 127186 338494
rect 127422 338258 127464 338494
rect 127144 331494 127464 338258
rect 127144 331258 127186 331494
rect 127422 331258 127464 331494
rect 127144 324494 127464 331258
rect 127144 324258 127186 324494
rect 127422 324258 127464 324494
rect 127144 317494 127464 324258
rect 127144 317258 127186 317494
rect 127422 317258 127464 317494
rect 127144 310494 127464 317258
rect 127144 310258 127186 310494
rect 127422 310258 127464 310494
rect 127144 303494 127464 310258
rect 127144 303258 127186 303494
rect 127422 303258 127464 303494
rect 127144 296494 127464 303258
rect 127144 296258 127186 296494
rect 127422 296258 127464 296494
rect 127144 289494 127464 296258
rect 127144 289258 127186 289494
rect 127422 289258 127464 289494
rect 127144 282494 127464 289258
rect 127144 282258 127186 282494
rect 127422 282258 127464 282494
rect 127144 275494 127464 282258
rect 127144 275258 127186 275494
rect 127422 275258 127464 275494
rect 127144 268494 127464 275258
rect 127144 268258 127186 268494
rect 127422 268258 127464 268494
rect 127144 261494 127464 268258
rect 127144 261258 127186 261494
rect 127422 261258 127464 261494
rect 127144 254494 127464 261258
rect 127144 254258 127186 254494
rect 127422 254258 127464 254494
rect 127144 247494 127464 254258
rect 127144 247258 127186 247494
rect 127422 247258 127464 247494
rect 127144 240494 127464 247258
rect 127144 240258 127186 240494
rect 127422 240258 127464 240494
rect 127144 233494 127464 240258
rect 127144 233258 127186 233494
rect 127422 233258 127464 233494
rect 127144 226494 127464 233258
rect 127144 226258 127186 226494
rect 127422 226258 127464 226494
rect 127144 219494 127464 226258
rect 127144 219258 127186 219494
rect 127422 219258 127464 219494
rect 127144 212494 127464 219258
rect 127144 212258 127186 212494
rect 127422 212258 127464 212494
rect 127144 205494 127464 212258
rect 127144 205258 127186 205494
rect 127422 205258 127464 205494
rect 127144 198494 127464 205258
rect 127144 198258 127186 198494
rect 127422 198258 127464 198494
rect 127144 191494 127464 198258
rect 127144 191258 127186 191494
rect 127422 191258 127464 191494
rect 127144 184494 127464 191258
rect 127144 184258 127186 184494
rect 127422 184258 127464 184494
rect 127144 177494 127464 184258
rect 127144 177258 127186 177494
rect 127422 177258 127464 177494
rect 127144 170494 127464 177258
rect 127144 170258 127186 170494
rect 127422 170258 127464 170494
rect 127144 163494 127464 170258
rect 127144 163258 127186 163494
rect 127422 163258 127464 163494
rect 127144 156494 127464 163258
rect 127144 156258 127186 156494
rect 127422 156258 127464 156494
rect 127144 149494 127464 156258
rect 127144 149258 127186 149494
rect 127422 149258 127464 149494
rect 127144 142494 127464 149258
rect 127144 142258 127186 142494
rect 127422 142258 127464 142494
rect 127144 135494 127464 142258
rect 127144 135258 127186 135494
rect 127422 135258 127464 135494
rect 127144 128494 127464 135258
rect 127144 128258 127186 128494
rect 127422 128258 127464 128494
rect 127144 121494 127464 128258
rect 127144 121258 127186 121494
rect 127422 121258 127464 121494
rect 127144 114494 127464 121258
rect 127144 114258 127186 114494
rect 127422 114258 127464 114494
rect 127144 107494 127464 114258
rect 127144 107258 127186 107494
rect 127422 107258 127464 107494
rect 127144 100494 127464 107258
rect 127144 100258 127186 100494
rect 127422 100258 127464 100494
rect 127144 93494 127464 100258
rect 127144 93258 127186 93494
rect 127422 93258 127464 93494
rect 127144 86494 127464 93258
rect 127144 86258 127186 86494
rect 127422 86258 127464 86494
rect 127144 79494 127464 86258
rect 127144 79258 127186 79494
rect 127422 79258 127464 79494
rect 127144 72494 127464 79258
rect 127144 72258 127186 72494
rect 127422 72258 127464 72494
rect 127144 65494 127464 72258
rect 127144 65258 127186 65494
rect 127422 65258 127464 65494
rect 127144 58494 127464 65258
rect 127144 58258 127186 58494
rect 127422 58258 127464 58494
rect 127144 51494 127464 58258
rect 127144 51258 127186 51494
rect 127422 51258 127464 51494
rect 127144 44494 127464 51258
rect 127144 44258 127186 44494
rect 127422 44258 127464 44494
rect 127144 37494 127464 44258
rect 127144 37258 127186 37494
rect 127422 37258 127464 37494
rect 127144 30494 127464 37258
rect 127144 30258 127186 30494
rect 127422 30258 127464 30494
rect 127144 23494 127464 30258
rect 127144 23258 127186 23494
rect 127422 23258 127464 23494
rect 127144 16494 127464 23258
rect 127144 16258 127186 16494
rect 127422 16258 127464 16494
rect 127144 9494 127464 16258
rect 127144 9258 127186 9494
rect 127422 9258 127464 9494
rect 127144 2494 127464 9258
rect 127144 2258 127186 2494
rect 127422 2258 127464 2494
rect 127144 -746 127464 2258
rect 127144 -982 127186 -746
rect 127422 -982 127464 -746
rect 127144 -1066 127464 -982
rect 127144 -1302 127186 -1066
rect 127422 -1302 127464 -1066
rect 127144 -2294 127464 -1302
rect 128876 706198 129196 706230
rect 128876 705962 128918 706198
rect 129154 705962 129196 706198
rect 128876 705878 129196 705962
rect 128876 705642 128918 705878
rect 129154 705642 129196 705878
rect 128876 696561 129196 705642
rect 128876 696325 128918 696561
rect 129154 696325 129196 696561
rect 128876 689561 129196 696325
rect 128876 689325 128918 689561
rect 129154 689325 129196 689561
rect 128876 682561 129196 689325
rect 128876 682325 128918 682561
rect 129154 682325 129196 682561
rect 128876 675561 129196 682325
rect 128876 675325 128918 675561
rect 129154 675325 129196 675561
rect 128876 668561 129196 675325
rect 128876 668325 128918 668561
rect 129154 668325 129196 668561
rect 128876 661561 129196 668325
rect 128876 661325 128918 661561
rect 129154 661325 129196 661561
rect 128876 654561 129196 661325
rect 128876 654325 128918 654561
rect 129154 654325 129196 654561
rect 128876 647561 129196 654325
rect 128876 647325 128918 647561
rect 129154 647325 129196 647561
rect 128876 640561 129196 647325
rect 128876 640325 128918 640561
rect 129154 640325 129196 640561
rect 128876 633561 129196 640325
rect 128876 633325 128918 633561
rect 129154 633325 129196 633561
rect 128876 626561 129196 633325
rect 128876 626325 128918 626561
rect 129154 626325 129196 626561
rect 128876 619561 129196 626325
rect 128876 619325 128918 619561
rect 129154 619325 129196 619561
rect 128876 612561 129196 619325
rect 128876 612325 128918 612561
rect 129154 612325 129196 612561
rect 128876 605561 129196 612325
rect 128876 605325 128918 605561
rect 129154 605325 129196 605561
rect 128876 598561 129196 605325
rect 128876 598325 128918 598561
rect 129154 598325 129196 598561
rect 128876 591561 129196 598325
rect 128876 591325 128918 591561
rect 129154 591325 129196 591561
rect 128876 584561 129196 591325
rect 128876 584325 128918 584561
rect 129154 584325 129196 584561
rect 128876 577561 129196 584325
rect 128876 577325 128918 577561
rect 129154 577325 129196 577561
rect 128876 570561 129196 577325
rect 128876 570325 128918 570561
rect 129154 570325 129196 570561
rect 128876 563561 129196 570325
rect 128876 563325 128918 563561
rect 129154 563325 129196 563561
rect 128876 556561 129196 563325
rect 128876 556325 128918 556561
rect 129154 556325 129196 556561
rect 128876 549561 129196 556325
rect 128876 549325 128918 549561
rect 129154 549325 129196 549561
rect 128876 542561 129196 549325
rect 128876 542325 128918 542561
rect 129154 542325 129196 542561
rect 128876 535561 129196 542325
rect 128876 535325 128918 535561
rect 129154 535325 129196 535561
rect 128876 528561 129196 535325
rect 128876 528325 128918 528561
rect 129154 528325 129196 528561
rect 128876 521561 129196 528325
rect 128876 521325 128918 521561
rect 129154 521325 129196 521561
rect 128876 514561 129196 521325
rect 128876 514325 128918 514561
rect 129154 514325 129196 514561
rect 128876 507561 129196 514325
rect 128876 507325 128918 507561
rect 129154 507325 129196 507561
rect 128876 500561 129196 507325
rect 128876 500325 128918 500561
rect 129154 500325 129196 500561
rect 128876 493561 129196 500325
rect 128876 493325 128918 493561
rect 129154 493325 129196 493561
rect 128876 486561 129196 493325
rect 128876 486325 128918 486561
rect 129154 486325 129196 486561
rect 128876 479561 129196 486325
rect 128876 479325 128918 479561
rect 129154 479325 129196 479561
rect 128876 472561 129196 479325
rect 128876 472325 128918 472561
rect 129154 472325 129196 472561
rect 128876 465561 129196 472325
rect 128876 465325 128918 465561
rect 129154 465325 129196 465561
rect 128876 458561 129196 465325
rect 128876 458325 128918 458561
rect 129154 458325 129196 458561
rect 128876 451561 129196 458325
rect 128876 451325 128918 451561
rect 129154 451325 129196 451561
rect 128876 444561 129196 451325
rect 128876 444325 128918 444561
rect 129154 444325 129196 444561
rect 128876 437561 129196 444325
rect 128876 437325 128918 437561
rect 129154 437325 129196 437561
rect 128876 430561 129196 437325
rect 128876 430325 128918 430561
rect 129154 430325 129196 430561
rect 128876 423561 129196 430325
rect 128876 423325 128918 423561
rect 129154 423325 129196 423561
rect 128876 416561 129196 423325
rect 128876 416325 128918 416561
rect 129154 416325 129196 416561
rect 128876 409561 129196 416325
rect 128876 409325 128918 409561
rect 129154 409325 129196 409561
rect 128876 402561 129196 409325
rect 128876 402325 128918 402561
rect 129154 402325 129196 402561
rect 128876 395561 129196 402325
rect 128876 395325 128918 395561
rect 129154 395325 129196 395561
rect 128876 388561 129196 395325
rect 128876 388325 128918 388561
rect 129154 388325 129196 388561
rect 128876 381561 129196 388325
rect 128876 381325 128918 381561
rect 129154 381325 129196 381561
rect 128876 374561 129196 381325
rect 128876 374325 128918 374561
rect 129154 374325 129196 374561
rect 128876 367561 129196 374325
rect 128876 367325 128918 367561
rect 129154 367325 129196 367561
rect 128876 360561 129196 367325
rect 128876 360325 128918 360561
rect 129154 360325 129196 360561
rect 128876 353561 129196 360325
rect 128876 353325 128918 353561
rect 129154 353325 129196 353561
rect 128876 346561 129196 353325
rect 128876 346325 128918 346561
rect 129154 346325 129196 346561
rect 128876 339561 129196 346325
rect 128876 339325 128918 339561
rect 129154 339325 129196 339561
rect 128876 332561 129196 339325
rect 128876 332325 128918 332561
rect 129154 332325 129196 332561
rect 128876 325561 129196 332325
rect 128876 325325 128918 325561
rect 129154 325325 129196 325561
rect 128876 318561 129196 325325
rect 128876 318325 128918 318561
rect 129154 318325 129196 318561
rect 128876 311561 129196 318325
rect 128876 311325 128918 311561
rect 129154 311325 129196 311561
rect 128876 304561 129196 311325
rect 128876 304325 128918 304561
rect 129154 304325 129196 304561
rect 128876 297561 129196 304325
rect 128876 297325 128918 297561
rect 129154 297325 129196 297561
rect 128876 290561 129196 297325
rect 128876 290325 128918 290561
rect 129154 290325 129196 290561
rect 128876 283561 129196 290325
rect 128876 283325 128918 283561
rect 129154 283325 129196 283561
rect 128876 276561 129196 283325
rect 128876 276325 128918 276561
rect 129154 276325 129196 276561
rect 128876 269561 129196 276325
rect 128876 269325 128918 269561
rect 129154 269325 129196 269561
rect 128876 262561 129196 269325
rect 128876 262325 128918 262561
rect 129154 262325 129196 262561
rect 128876 255561 129196 262325
rect 128876 255325 128918 255561
rect 129154 255325 129196 255561
rect 128876 248561 129196 255325
rect 128876 248325 128918 248561
rect 129154 248325 129196 248561
rect 128876 241561 129196 248325
rect 128876 241325 128918 241561
rect 129154 241325 129196 241561
rect 128876 234561 129196 241325
rect 128876 234325 128918 234561
rect 129154 234325 129196 234561
rect 128876 227561 129196 234325
rect 128876 227325 128918 227561
rect 129154 227325 129196 227561
rect 128876 220561 129196 227325
rect 128876 220325 128918 220561
rect 129154 220325 129196 220561
rect 128876 213561 129196 220325
rect 128876 213325 128918 213561
rect 129154 213325 129196 213561
rect 128876 206561 129196 213325
rect 128876 206325 128918 206561
rect 129154 206325 129196 206561
rect 128876 199561 129196 206325
rect 128876 199325 128918 199561
rect 129154 199325 129196 199561
rect 128876 192561 129196 199325
rect 128876 192325 128918 192561
rect 129154 192325 129196 192561
rect 128876 185561 129196 192325
rect 128876 185325 128918 185561
rect 129154 185325 129196 185561
rect 128876 178561 129196 185325
rect 128876 178325 128918 178561
rect 129154 178325 129196 178561
rect 128876 171561 129196 178325
rect 128876 171325 128918 171561
rect 129154 171325 129196 171561
rect 128876 164561 129196 171325
rect 128876 164325 128918 164561
rect 129154 164325 129196 164561
rect 128876 157561 129196 164325
rect 128876 157325 128918 157561
rect 129154 157325 129196 157561
rect 128876 150561 129196 157325
rect 128876 150325 128918 150561
rect 129154 150325 129196 150561
rect 128876 143561 129196 150325
rect 128876 143325 128918 143561
rect 129154 143325 129196 143561
rect 128876 136561 129196 143325
rect 128876 136325 128918 136561
rect 129154 136325 129196 136561
rect 128876 129561 129196 136325
rect 128876 129325 128918 129561
rect 129154 129325 129196 129561
rect 128876 122561 129196 129325
rect 128876 122325 128918 122561
rect 129154 122325 129196 122561
rect 128876 115561 129196 122325
rect 128876 115325 128918 115561
rect 129154 115325 129196 115561
rect 128876 108561 129196 115325
rect 128876 108325 128918 108561
rect 129154 108325 129196 108561
rect 128876 101561 129196 108325
rect 128876 101325 128918 101561
rect 129154 101325 129196 101561
rect 128876 94561 129196 101325
rect 128876 94325 128918 94561
rect 129154 94325 129196 94561
rect 128876 87561 129196 94325
rect 128876 87325 128918 87561
rect 129154 87325 129196 87561
rect 128876 80561 129196 87325
rect 128876 80325 128918 80561
rect 129154 80325 129196 80561
rect 128876 73561 129196 80325
rect 128876 73325 128918 73561
rect 129154 73325 129196 73561
rect 128876 66561 129196 73325
rect 128876 66325 128918 66561
rect 129154 66325 129196 66561
rect 128876 59561 129196 66325
rect 128876 59325 128918 59561
rect 129154 59325 129196 59561
rect 128876 52561 129196 59325
rect 128876 52325 128918 52561
rect 129154 52325 129196 52561
rect 128876 45561 129196 52325
rect 128876 45325 128918 45561
rect 129154 45325 129196 45561
rect 128876 38561 129196 45325
rect 128876 38325 128918 38561
rect 129154 38325 129196 38561
rect 128876 31561 129196 38325
rect 128876 31325 128918 31561
rect 129154 31325 129196 31561
rect 128876 24561 129196 31325
rect 128876 24325 128918 24561
rect 129154 24325 129196 24561
rect 128876 17561 129196 24325
rect 128876 17325 128918 17561
rect 129154 17325 129196 17561
rect 128876 10561 129196 17325
rect 128876 10325 128918 10561
rect 129154 10325 129196 10561
rect 128876 3561 129196 10325
rect 128876 3325 128918 3561
rect 129154 3325 129196 3561
rect 128876 -1706 129196 3325
rect 128876 -1942 128918 -1706
rect 129154 -1942 129196 -1706
rect 128876 -2026 129196 -1942
rect 128876 -2262 128918 -2026
rect 129154 -2262 129196 -2026
rect 128876 -2294 129196 -2262
rect 134144 705238 134464 706230
rect 134144 705002 134186 705238
rect 134422 705002 134464 705238
rect 134144 704918 134464 705002
rect 134144 704682 134186 704918
rect 134422 704682 134464 704918
rect 134144 695494 134464 704682
rect 134144 695258 134186 695494
rect 134422 695258 134464 695494
rect 134144 688494 134464 695258
rect 134144 688258 134186 688494
rect 134422 688258 134464 688494
rect 134144 681494 134464 688258
rect 134144 681258 134186 681494
rect 134422 681258 134464 681494
rect 134144 674494 134464 681258
rect 134144 674258 134186 674494
rect 134422 674258 134464 674494
rect 134144 667494 134464 674258
rect 134144 667258 134186 667494
rect 134422 667258 134464 667494
rect 134144 660494 134464 667258
rect 134144 660258 134186 660494
rect 134422 660258 134464 660494
rect 134144 653494 134464 660258
rect 134144 653258 134186 653494
rect 134422 653258 134464 653494
rect 134144 646494 134464 653258
rect 134144 646258 134186 646494
rect 134422 646258 134464 646494
rect 134144 639494 134464 646258
rect 134144 639258 134186 639494
rect 134422 639258 134464 639494
rect 134144 632494 134464 639258
rect 134144 632258 134186 632494
rect 134422 632258 134464 632494
rect 134144 625494 134464 632258
rect 134144 625258 134186 625494
rect 134422 625258 134464 625494
rect 134144 618494 134464 625258
rect 134144 618258 134186 618494
rect 134422 618258 134464 618494
rect 134144 611494 134464 618258
rect 134144 611258 134186 611494
rect 134422 611258 134464 611494
rect 134144 604494 134464 611258
rect 134144 604258 134186 604494
rect 134422 604258 134464 604494
rect 134144 597494 134464 604258
rect 134144 597258 134186 597494
rect 134422 597258 134464 597494
rect 134144 590494 134464 597258
rect 134144 590258 134186 590494
rect 134422 590258 134464 590494
rect 134144 583494 134464 590258
rect 134144 583258 134186 583494
rect 134422 583258 134464 583494
rect 134144 576494 134464 583258
rect 134144 576258 134186 576494
rect 134422 576258 134464 576494
rect 134144 569494 134464 576258
rect 134144 569258 134186 569494
rect 134422 569258 134464 569494
rect 134144 562494 134464 569258
rect 134144 562258 134186 562494
rect 134422 562258 134464 562494
rect 134144 555494 134464 562258
rect 134144 555258 134186 555494
rect 134422 555258 134464 555494
rect 134144 548494 134464 555258
rect 134144 548258 134186 548494
rect 134422 548258 134464 548494
rect 134144 541494 134464 548258
rect 134144 541258 134186 541494
rect 134422 541258 134464 541494
rect 134144 534494 134464 541258
rect 134144 534258 134186 534494
rect 134422 534258 134464 534494
rect 134144 527494 134464 534258
rect 134144 527258 134186 527494
rect 134422 527258 134464 527494
rect 134144 520494 134464 527258
rect 134144 520258 134186 520494
rect 134422 520258 134464 520494
rect 134144 513494 134464 520258
rect 134144 513258 134186 513494
rect 134422 513258 134464 513494
rect 134144 506494 134464 513258
rect 134144 506258 134186 506494
rect 134422 506258 134464 506494
rect 134144 499494 134464 506258
rect 134144 499258 134186 499494
rect 134422 499258 134464 499494
rect 134144 492494 134464 499258
rect 134144 492258 134186 492494
rect 134422 492258 134464 492494
rect 134144 485494 134464 492258
rect 134144 485258 134186 485494
rect 134422 485258 134464 485494
rect 134144 478494 134464 485258
rect 134144 478258 134186 478494
rect 134422 478258 134464 478494
rect 134144 471494 134464 478258
rect 134144 471258 134186 471494
rect 134422 471258 134464 471494
rect 134144 464494 134464 471258
rect 134144 464258 134186 464494
rect 134422 464258 134464 464494
rect 134144 457494 134464 464258
rect 134144 457258 134186 457494
rect 134422 457258 134464 457494
rect 134144 450494 134464 457258
rect 134144 450258 134186 450494
rect 134422 450258 134464 450494
rect 134144 443494 134464 450258
rect 134144 443258 134186 443494
rect 134422 443258 134464 443494
rect 134144 436494 134464 443258
rect 134144 436258 134186 436494
rect 134422 436258 134464 436494
rect 134144 429494 134464 436258
rect 134144 429258 134186 429494
rect 134422 429258 134464 429494
rect 134144 422494 134464 429258
rect 134144 422258 134186 422494
rect 134422 422258 134464 422494
rect 134144 415494 134464 422258
rect 134144 415258 134186 415494
rect 134422 415258 134464 415494
rect 134144 408494 134464 415258
rect 134144 408258 134186 408494
rect 134422 408258 134464 408494
rect 134144 401494 134464 408258
rect 134144 401258 134186 401494
rect 134422 401258 134464 401494
rect 134144 394494 134464 401258
rect 134144 394258 134186 394494
rect 134422 394258 134464 394494
rect 134144 387494 134464 394258
rect 134144 387258 134186 387494
rect 134422 387258 134464 387494
rect 134144 380494 134464 387258
rect 134144 380258 134186 380494
rect 134422 380258 134464 380494
rect 134144 373494 134464 380258
rect 134144 373258 134186 373494
rect 134422 373258 134464 373494
rect 134144 366494 134464 373258
rect 134144 366258 134186 366494
rect 134422 366258 134464 366494
rect 134144 359494 134464 366258
rect 134144 359258 134186 359494
rect 134422 359258 134464 359494
rect 134144 352494 134464 359258
rect 134144 352258 134186 352494
rect 134422 352258 134464 352494
rect 134144 345494 134464 352258
rect 134144 345258 134186 345494
rect 134422 345258 134464 345494
rect 134144 338494 134464 345258
rect 134144 338258 134186 338494
rect 134422 338258 134464 338494
rect 134144 331494 134464 338258
rect 134144 331258 134186 331494
rect 134422 331258 134464 331494
rect 134144 324494 134464 331258
rect 134144 324258 134186 324494
rect 134422 324258 134464 324494
rect 134144 317494 134464 324258
rect 134144 317258 134186 317494
rect 134422 317258 134464 317494
rect 134144 310494 134464 317258
rect 134144 310258 134186 310494
rect 134422 310258 134464 310494
rect 134144 303494 134464 310258
rect 134144 303258 134186 303494
rect 134422 303258 134464 303494
rect 134144 296494 134464 303258
rect 134144 296258 134186 296494
rect 134422 296258 134464 296494
rect 134144 289494 134464 296258
rect 134144 289258 134186 289494
rect 134422 289258 134464 289494
rect 134144 282494 134464 289258
rect 134144 282258 134186 282494
rect 134422 282258 134464 282494
rect 134144 275494 134464 282258
rect 134144 275258 134186 275494
rect 134422 275258 134464 275494
rect 134144 268494 134464 275258
rect 134144 268258 134186 268494
rect 134422 268258 134464 268494
rect 134144 261494 134464 268258
rect 134144 261258 134186 261494
rect 134422 261258 134464 261494
rect 134144 254494 134464 261258
rect 134144 254258 134186 254494
rect 134422 254258 134464 254494
rect 134144 247494 134464 254258
rect 134144 247258 134186 247494
rect 134422 247258 134464 247494
rect 134144 240494 134464 247258
rect 134144 240258 134186 240494
rect 134422 240258 134464 240494
rect 134144 233494 134464 240258
rect 134144 233258 134186 233494
rect 134422 233258 134464 233494
rect 134144 226494 134464 233258
rect 134144 226258 134186 226494
rect 134422 226258 134464 226494
rect 134144 219494 134464 226258
rect 134144 219258 134186 219494
rect 134422 219258 134464 219494
rect 134144 212494 134464 219258
rect 134144 212258 134186 212494
rect 134422 212258 134464 212494
rect 134144 205494 134464 212258
rect 134144 205258 134186 205494
rect 134422 205258 134464 205494
rect 134144 198494 134464 205258
rect 134144 198258 134186 198494
rect 134422 198258 134464 198494
rect 134144 191494 134464 198258
rect 134144 191258 134186 191494
rect 134422 191258 134464 191494
rect 134144 184494 134464 191258
rect 134144 184258 134186 184494
rect 134422 184258 134464 184494
rect 134144 177494 134464 184258
rect 134144 177258 134186 177494
rect 134422 177258 134464 177494
rect 134144 170494 134464 177258
rect 134144 170258 134186 170494
rect 134422 170258 134464 170494
rect 134144 163494 134464 170258
rect 134144 163258 134186 163494
rect 134422 163258 134464 163494
rect 134144 156494 134464 163258
rect 134144 156258 134186 156494
rect 134422 156258 134464 156494
rect 134144 149494 134464 156258
rect 134144 149258 134186 149494
rect 134422 149258 134464 149494
rect 134144 142494 134464 149258
rect 134144 142258 134186 142494
rect 134422 142258 134464 142494
rect 134144 135494 134464 142258
rect 134144 135258 134186 135494
rect 134422 135258 134464 135494
rect 134144 128494 134464 135258
rect 134144 128258 134186 128494
rect 134422 128258 134464 128494
rect 134144 121494 134464 128258
rect 134144 121258 134186 121494
rect 134422 121258 134464 121494
rect 134144 114494 134464 121258
rect 134144 114258 134186 114494
rect 134422 114258 134464 114494
rect 134144 107494 134464 114258
rect 134144 107258 134186 107494
rect 134422 107258 134464 107494
rect 134144 100494 134464 107258
rect 134144 100258 134186 100494
rect 134422 100258 134464 100494
rect 134144 93494 134464 100258
rect 134144 93258 134186 93494
rect 134422 93258 134464 93494
rect 134144 86494 134464 93258
rect 134144 86258 134186 86494
rect 134422 86258 134464 86494
rect 134144 79494 134464 86258
rect 134144 79258 134186 79494
rect 134422 79258 134464 79494
rect 134144 72494 134464 79258
rect 134144 72258 134186 72494
rect 134422 72258 134464 72494
rect 134144 65494 134464 72258
rect 134144 65258 134186 65494
rect 134422 65258 134464 65494
rect 134144 58494 134464 65258
rect 134144 58258 134186 58494
rect 134422 58258 134464 58494
rect 134144 51494 134464 58258
rect 134144 51258 134186 51494
rect 134422 51258 134464 51494
rect 134144 44494 134464 51258
rect 134144 44258 134186 44494
rect 134422 44258 134464 44494
rect 134144 37494 134464 44258
rect 134144 37258 134186 37494
rect 134422 37258 134464 37494
rect 134144 30494 134464 37258
rect 134144 30258 134186 30494
rect 134422 30258 134464 30494
rect 134144 23494 134464 30258
rect 134144 23258 134186 23494
rect 134422 23258 134464 23494
rect 134144 16494 134464 23258
rect 134144 16258 134186 16494
rect 134422 16258 134464 16494
rect 134144 9494 134464 16258
rect 134144 9258 134186 9494
rect 134422 9258 134464 9494
rect 134144 2494 134464 9258
rect 134144 2258 134186 2494
rect 134422 2258 134464 2494
rect 134144 -746 134464 2258
rect 134144 -982 134186 -746
rect 134422 -982 134464 -746
rect 134144 -1066 134464 -982
rect 134144 -1302 134186 -1066
rect 134422 -1302 134464 -1066
rect 134144 -2294 134464 -1302
rect 135876 706198 136196 706230
rect 135876 705962 135918 706198
rect 136154 705962 136196 706198
rect 135876 705878 136196 705962
rect 135876 705642 135918 705878
rect 136154 705642 136196 705878
rect 135876 696561 136196 705642
rect 135876 696325 135918 696561
rect 136154 696325 136196 696561
rect 135876 689561 136196 696325
rect 135876 689325 135918 689561
rect 136154 689325 136196 689561
rect 135876 682561 136196 689325
rect 135876 682325 135918 682561
rect 136154 682325 136196 682561
rect 135876 675561 136196 682325
rect 135876 675325 135918 675561
rect 136154 675325 136196 675561
rect 135876 668561 136196 675325
rect 135876 668325 135918 668561
rect 136154 668325 136196 668561
rect 135876 661561 136196 668325
rect 135876 661325 135918 661561
rect 136154 661325 136196 661561
rect 135876 654561 136196 661325
rect 135876 654325 135918 654561
rect 136154 654325 136196 654561
rect 135876 647561 136196 654325
rect 135876 647325 135918 647561
rect 136154 647325 136196 647561
rect 135876 640561 136196 647325
rect 135876 640325 135918 640561
rect 136154 640325 136196 640561
rect 135876 633561 136196 640325
rect 135876 633325 135918 633561
rect 136154 633325 136196 633561
rect 135876 626561 136196 633325
rect 135876 626325 135918 626561
rect 136154 626325 136196 626561
rect 135876 619561 136196 626325
rect 135876 619325 135918 619561
rect 136154 619325 136196 619561
rect 135876 612561 136196 619325
rect 135876 612325 135918 612561
rect 136154 612325 136196 612561
rect 135876 605561 136196 612325
rect 135876 605325 135918 605561
rect 136154 605325 136196 605561
rect 135876 598561 136196 605325
rect 135876 598325 135918 598561
rect 136154 598325 136196 598561
rect 135876 591561 136196 598325
rect 135876 591325 135918 591561
rect 136154 591325 136196 591561
rect 135876 584561 136196 591325
rect 135876 584325 135918 584561
rect 136154 584325 136196 584561
rect 135876 577561 136196 584325
rect 135876 577325 135918 577561
rect 136154 577325 136196 577561
rect 135876 570561 136196 577325
rect 135876 570325 135918 570561
rect 136154 570325 136196 570561
rect 135876 563561 136196 570325
rect 135876 563325 135918 563561
rect 136154 563325 136196 563561
rect 135876 556561 136196 563325
rect 135876 556325 135918 556561
rect 136154 556325 136196 556561
rect 135876 549561 136196 556325
rect 135876 549325 135918 549561
rect 136154 549325 136196 549561
rect 135876 542561 136196 549325
rect 135876 542325 135918 542561
rect 136154 542325 136196 542561
rect 135876 535561 136196 542325
rect 135876 535325 135918 535561
rect 136154 535325 136196 535561
rect 135876 528561 136196 535325
rect 135876 528325 135918 528561
rect 136154 528325 136196 528561
rect 135876 521561 136196 528325
rect 135876 521325 135918 521561
rect 136154 521325 136196 521561
rect 135876 514561 136196 521325
rect 135876 514325 135918 514561
rect 136154 514325 136196 514561
rect 135876 507561 136196 514325
rect 135876 507325 135918 507561
rect 136154 507325 136196 507561
rect 135876 500561 136196 507325
rect 135876 500325 135918 500561
rect 136154 500325 136196 500561
rect 135876 493561 136196 500325
rect 135876 493325 135918 493561
rect 136154 493325 136196 493561
rect 135876 486561 136196 493325
rect 135876 486325 135918 486561
rect 136154 486325 136196 486561
rect 135876 479561 136196 486325
rect 135876 479325 135918 479561
rect 136154 479325 136196 479561
rect 135876 472561 136196 479325
rect 135876 472325 135918 472561
rect 136154 472325 136196 472561
rect 135876 465561 136196 472325
rect 135876 465325 135918 465561
rect 136154 465325 136196 465561
rect 135876 458561 136196 465325
rect 135876 458325 135918 458561
rect 136154 458325 136196 458561
rect 135876 451561 136196 458325
rect 135876 451325 135918 451561
rect 136154 451325 136196 451561
rect 135876 444561 136196 451325
rect 135876 444325 135918 444561
rect 136154 444325 136196 444561
rect 135876 437561 136196 444325
rect 135876 437325 135918 437561
rect 136154 437325 136196 437561
rect 135876 430561 136196 437325
rect 135876 430325 135918 430561
rect 136154 430325 136196 430561
rect 135876 423561 136196 430325
rect 135876 423325 135918 423561
rect 136154 423325 136196 423561
rect 135876 416561 136196 423325
rect 135876 416325 135918 416561
rect 136154 416325 136196 416561
rect 135876 409561 136196 416325
rect 135876 409325 135918 409561
rect 136154 409325 136196 409561
rect 135876 402561 136196 409325
rect 135876 402325 135918 402561
rect 136154 402325 136196 402561
rect 135876 395561 136196 402325
rect 135876 395325 135918 395561
rect 136154 395325 136196 395561
rect 135876 388561 136196 395325
rect 135876 388325 135918 388561
rect 136154 388325 136196 388561
rect 135876 381561 136196 388325
rect 135876 381325 135918 381561
rect 136154 381325 136196 381561
rect 135876 374561 136196 381325
rect 135876 374325 135918 374561
rect 136154 374325 136196 374561
rect 135876 367561 136196 374325
rect 135876 367325 135918 367561
rect 136154 367325 136196 367561
rect 135876 360561 136196 367325
rect 135876 360325 135918 360561
rect 136154 360325 136196 360561
rect 135876 353561 136196 360325
rect 135876 353325 135918 353561
rect 136154 353325 136196 353561
rect 135876 346561 136196 353325
rect 135876 346325 135918 346561
rect 136154 346325 136196 346561
rect 135876 339561 136196 346325
rect 135876 339325 135918 339561
rect 136154 339325 136196 339561
rect 135876 332561 136196 339325
rect 135876 332325 135918 332561
rect 136154 332325 136196 332561
rect 135876 325561 136196 332325
rect 135876 325325 135918 325561
rect 136154 325325 136196 325561
rect 135876 318561 136196 325325
rect 135876 318325 135918 318561
rect 136154 318325 136196 318561
rect 135876 311561 136196 318325
rect 135876 311325 135918 311561
rect 136154 311325 136196 311561
rect 135876 304561 136196 311325
rect 135876 304325 135918 304561
rect 136154 304325 136196 304561
rect 135876 297561 136196 304325
rect 135876 297325 135918 297561
rect 136154 297325 136196 297561
rect 135876 290561 136196 297325
rect 135876 290325 135918 290561
rect 136154 290325 136196 290561
rect 135876 283561 136196 290325
rect 135876 283325 135918 283561
rect 136154 283325 136196 283561
rect 135876 276561 136196 283325
rect 135876 276325 135918 276561
rect 136154 276325 136196 276561
rect 135876 269561 136196 276325
rect 135876 269325 135918 269561
rect 136154 269325 136196 269561
rect 135876 262561 136196 269325
rect 135876 262325 135918 262561
rect 136154 262325 136196 262561
rect 135876 255561 136196 262325
rect 135876 255325 135918 255561
rect 136154 255325 136196 255561
rect 135876 248561 136196 255325
rect 135876 248325 135918 248561
rect 136154 248325 136196 248561
rect 135876 241561 136196 248325
rect 135876 241325 135918 241561
rect 136154 241325 136196 241561
rect 135876 234561 136196 241325
rect 135876 234325 135918 234561
rect 136154 234325 136196 234561
rect 135876 227561 136196 234325
rect 135876 227325 135918 227561
rect 136154 227325 136196 227561
rect 135876 220561 136196 227325
rect 135876 220325 135918 220561
rect 136154 220325 136196 220561
rect 135876 213561 136196 220325
rect 135876 213325 135918 213561
rect 136154 213325 136196 213561
rect 135876 206561 136196 213325
rect 135876 206325 135918 206561
rect 136154 206325 136196 206561
rect 135876 199561 136196 206325
rect 135876 199325 135918 199561
rect 136154 199325 136196 199561
rect 135876 192561 136196 199325
rect 135876 192325 135918 192561
rect 136154 192325 136196 192561
rect 135876 185561 136196 192325
rect 135876 185325 135918 185561
rect 136154 185325 136196 185561
rect 135876 178561 136196 185325
rect 135876 178325 135918 178561
rect 136154 178325 136196 178561
rect 135876 171561 136196 178325
rect 135876 171325 135918 171561
rect 136154 171325 136196 171561
rect 135876 164561 136196 171325
rect 135876 164325 135918 164561
rect 136154 164325 136196 164561
rect 135876 157561 136196 164325
rect 135876 157325 135918 157561
rect 136154 157325 136196 157561
rect 135876 150561 136196 157325
rect 135876 150325 135918 150561
rect 136154 150325 136196 150561
rect 135876 143561 136196 150325
rect 135876 143325 135918 143561
rect 136154 143325 136196 143561
rect 135876 136561 136196 143325
rect 135876 136325 135918 136561
rect 136154 136325 136196 136561
rect 135876 129561 136196 136325
rect 135876 129325 135918 129561
rect 136154 129325 136196 129561
rect 135876 122561 136196 129325
rect 135876 122325 135918 122561
rect 136154 122325 136196 122561
rect 135876 115561 136196 122325
rect 135876 115325 135918 115561
rect 136154 115325 136196 115561
rect 135876 108561 136196 115325
rect 135876 108325 135918 108561
rect 136154 108325 136196 108561
rect 135876 101561 136196 108325
rect 135876 101325 135918 101561
rect 136154 101325 136196 101561
rect 135876 94561 136196 101325
rect 135876 94325 135918 94561
rect 136154 94325 136196 94561
rect 135876 87561 136196 94325
rect 135876 87325 135918 87561
rect 136154 87325 136196 87561
rect 135876 80561 136196 87325
rect 135876 80325 135918 80561
rect 136154 80325 136196 80561
rect 135876 73561 136196 80325
rect 135876 73325 135918 73561
rect 136154 73325 136196 73561
rect 135876 66561 136196 73325
rect 135876 66325 135918 66561
rect 136154 66325 136196 66561
rect 135876 59561 136196 66325
rect 135876 59325 135918 59561
rect 136154 59325 136196 59561
rect 135876 52561 136196 59325
rect 135876 52325 135918 52561
rect 136154 52325 136196 52561
rect 135876 45561 136196 52325
rect 135876 45325 135918 45561
rect 136154 45325 136196 45561
rect 135876 38561 136196 45325
rect 135876 38325 135918 38561
rect 136154 38325 136196 38561
rect 135876 31561 136196 38325
rect 135876 31325 135918 31561
rect 136154 31325 136196 31561
rect 135876 24561 136196 31325
rect 135876 24325 135918 24561
rect 136154 24325 136196 24561
rect 135876 17561 136196 24325
rect 135876 17325 135918 17561
rect 136154 17325 136196 17561
rect 135876 10561 136196 17325
rect 135876 10325 135918 10561
rect 136154 10325 136196 10561
rect 135876 3561 136196 10325
rect 135876 3325 135918 3561
rect 136154 3325 136196 3561
rect 135876 -1706 136196 3325
rect 135876 -1942 135918 -1706
rect 136154 -1942 136196 -1706
rect 135876 -2026 136196 -1942
rect 135876 -2262 135918 -2026
rect 136154 -2262 136196 -2026
rect 135876 -2294 136196 -2262
rect 141144 705238 141464 706230
rect 141144 705002 141186 705238
rect 141422 705002 141464 705238
rect 141144 704918 141464 705002
rect 141144 704682 141186 704918
rect 141422 704682 141464 704918
rect 141144 695494 141464 704682
rect 141144 695258 141186 695494
rect 141422 695258 141464 695494
rect 141144 688494 141464 695258
rect 141144 688258 141186 688494
rect 141422 688258 141464 688494
rect 141144 681494 141464 688258
rect 141144 681258 141186 681494
rect 141422 681258 141464 681494
rect 141144 674494 141464 681258
rect 141144 674258 141186 674494
rect 141422 674258 141464 674494
rect 141144 667494 141464 674258
rect 141144 667258 141186 667494
rect 141422 667258 141464 667494
rect 141144 660494 141464 667258
rect 141144 660258 141186 660494
rect 141422 660258 141464 660494
rect 141144 653494 141464 660258
rect 141144 653258 141186 653494
rect 141422 653258 141464 653494
rect 141144 646494 141464 653258
rect 141144 646258 141186 646494
rect 141422 646258 141464 646494
rect 141144 639494 141464 646258
rect 141144 639258 141186 639494
rect 141422 639258 141464 639494
rect 141144 632494 141464 639258
rect 141144 632258 141186 632494
rect 141422 632258 141464 632494
rect 141144 625494 141464 632258
rect 141144 625258 141186 625494
rect 141422 625258 141464 625494
rect 141144 618494 141464 625258
rect 141144 618258 141186 618494
rect 141422 618258 141464 618494
rect 141144 611494 141464 618258
rect 141144 611258 141186 611494
rect 141422 611258 141464 611494
rect 141144 604494 141464 611258
rect 141144 604258 141186 604494
rect 141422 604258 141464 604494
rect 141144 597494 141464 604258
rect 141144 597258 141186 597494
rect 141422 597258 141464 597494
rect 141144 590494 141464 597258
rect 141144 590258 141186 590494
rect 141422 590258 141464 590494
rect 141144 583494 141464 590258
rect 141144 583258 141186 583494
rect 141422 583258 141464 583494
rect 141144 576494 141464 583258
rect 141144 576258 141186 576494
rect 141422 576258 141464 576494
rect 141144 569494 141464 576258
rect 141144 569258 141186 569494
rect 141422 569258 141464 569494
rect 141144 562494 141464 569258
rect 141144 562258 141186 562494
rect 141422 562258 141464 562494
rect 141144 555494 141464 562258
rect 141144 555258 141186 555494
rect 141422 555258 141464 555494
rect 141144 548494 141464 555258
rect 141144 548258 141186 548494
rect 141422 548258 141464 548494
rect 141144 541494 141464 548258
rect 141144 541258 141186 541494
rect 141422 541258 141464 541494
rect 141144 534494 141464 541258
rect 141144 534258 141186 534494
rect 141422 534258 141464 534494
rect 141144 527494 141464 534258
rect 141144 527258 141186 527494
rect 141422 527258 141464 527494
rect 141144 520494 141464 527258
rect 141144 520258 141186 520494
rect 141422 520258 141464 520494
rect 141144 513494 141464 520258
rect 141144 513258 141186 513494
rect 141422 513258 141464 513494
rect 141144 506494 141464 513258
rect 141144 506258 141186 506494
rect 141422 506258 141464 506494
rect 141144 499494 141464 506258
rect 141144 499258 141186 499494
rect 141422 499258 141464 499494
rect 141144 492494 141464 499258
rect 141144 492258 141186 492494
rect 141422 492258 141464 492494
rect 141144 485494 141464 492258
rect 141144 485258 141186 485494
rect 141422 485258 141464 485494
rect 141144 478494 141464 485258
rect 141144 478258 141186 478494
rect 141422 478258 141464 478494
rect 141144 471494 141464 478258
rect 141144 471258 141186 471494
rect 141422 471258 141464 471494
rect 141144 464494 141464 471258
rect 141144 464258 141186 464494
rect 141422 464258 141464 464494
rect 141144 457494 141464 464258
rect 141144 457258 141186 457494
rect 141422 457258 141464 457494
rect 141144 450494 141464 457258
rect 141144 450258 141186 450494
rect 141422 450258 141464 450494
rect 141144 443494 141464 450258
rect 141144 443258 141186 443494
rect 141422 443258 141464 443494
rect 141144 436494 141464 443258
rect 141144 436258 141186 436494
rect 141422 436258 141464 436494
rect 141144 429494 141464 436258
rect 141144 429258 141186 429494
rect 141422 429258 141464 429494
rect 141144 422494 141464 429258
rect 141144 422258 141186 422494
rect 141422 422258 141464 422494
rect 141144 415494 141464 422258
rect 141144 415258 141186 415494
rect 141422 415258 141464 415494
rect 141144 408494 141464 415258
rect 141144 408258 141186 408494
rect 141422 408258 141464 408494
rect 141144 401494 141464 408258
rect 141144 401258 141186 401494
rect 141422 401258 141464 401494
rect 141144 394494 141464 401258
rect 141144 394258 141186 394494
rect 141422 394258 141464 394494
rect 141144 387494 141464 394258
rect 141144 387258 141186 387494
rect 141422 387258 141464 387494
rect 141144 380494 141464 387258
rect 141144 380258 141186 380494
rect 141422 380258 141464 380494
rect 141144 373494 141464 380258
rect 141144 373258 141186 373494
rect 141422 373258 141464 373494
rect 141144 366494 141464 373258
rect 141144 366258 141186 366494
rect 141422 366258 141464 366494
rect 141144 359494 141464 366258
rect 141144 359258 141186 359494
rect 141422 359258 141464 359494
rect 141144 352494 141464 359258
rect 141144 352258 141186 352494
rect 141422 352258 141464 352494
rect 141144 345494 141464 352258
rect 141144 345258 141186 345494
rect 141422 345258 141464 345494
rect 141144 338494 141464 345258
rect 141144 338258 141186 338494
rect 141422 338258 141464 338494
rect 141144 331494 141464 338258
rect 141144 331258 141186 331494
rect 141422 331258 141464 331494
rect 141144 324494 141464 331258
rect 141144 324258 141186 324494
rect 141422 324258 141464 324494
rect 141144 317494 141464 324258
rect 141144 317258 141186 317494
rect 141422 317258 141464 317494
rect 141144 310494 141464 317258
rect 141144 310258 141186 310494
rect 141422 310258 141464 310494
rect 141144 303494 141464 310258
rect 141144 303258 141186 303494
rect 141422 303258 141464 303494
rect 141144 296494 141464 303258
rect 141144 296258 141186 296494
rect 141422 296258 141464 296494
rect 141144 289494 141464 296258
rect 141144 289258 141186 289494
rect 141422 289258 141464 289494
rect 141144 282494 141464 289258
rect 141144 282258 141186 282494
rect 141422 282258 141464 282494
rect 141144 275494 141464 282258
rect 141144 275258 141186 275494
rect 141422 275258 141464 275494
rect 141144 268494 141464 275258
rect 141144 268258 141186 268494
rect 141422 268258 141464 268494
rect 141144 261494 141464 268258
rect 141144 261258 141186 261494
rect 141422 261258 141464 261494
rect 141144 254494 141464 261258
rect 141144 254258 141186 254494
rect 141422 254258 141464 254494
rect 141144 247494 141464 254258
rect 141144 247258 141186 247494
rect 141422 247258 141464 247494
rect 141144 240494 141464 247258
rect 141144 240258 141186 240494
rect 141422 240258 141464 240494
rect 141144 233494 141464 240258
rect 141144 233258 141186 233494
rect 141422 233258 141464 233494
rect 141144 226494 141464 233258
rect 141144 226258 141186 226494
rect 141422 226258 141464 226494
rect 141144 219494 141464 226258
rect 141144 219258 141186 219494
rect 141422 219258 141464 219494
rect 141144 212494 141464 219258
rect 141144 212258 141186 212494
rect 141422 212258 141464 212494
rect 141144 205494 141464 212258
rect 141144 205258 141186 205494
rect 141422 205258 141464 205494
rect 141144 198494 141464 205258
rect 141144 198258 141186 198494
rect 141422 198258 141464 198494
rect 141144 191494 141464 198258
rect 141144 191258 141186 191494
rect 141422 191258 141464 191494
rect 141144 184494 141464 191258
rect 141144 184258 141186 184494
rect 141422 184258 141464 184494
rect 141144 177494 141464 184258
rect 141144 177258 141186 177494
rect 141422 177258 141464 177494
rect 141144 170494 141464 177258
rect 141144 170258 141186 170494
rect 141422 170258 141464 170494
rect 141144 163494 141464 170258
rect 141144 163258 141186 163494
rect 141422 163258 141464 163494
rect 141144 156494 141464 163258
rect 141144 156258 141186 156494
rect 141422 156258 141464 156494
rect 141144 149494 141464 156258
rect 141144 149258 141186 149494
rect 141422 149258 141464 149494
rect 141144 142494 141464 149258
rect 141144 142258 141186 142494
rect 141422 142258 141464 142494
rect 141144 135494 141464 142258
rect 141144 135258 141186 135494
rect 141422 135258 141464 135494
rect 141144 128494 141464 135258
rect 141144 128258 141186 128494
rect 141422 128258 141464 128494
rect 141144 121494 141464 128258
rect 141144 121258 141186 121494
rect 141422 121258 141464 121494
rect 141144 114494 141464 121258
rect 141144 114258 141186 114494
rect 141422 114258 141464 114494
rect 141144 107494 141464 114258
rect 141144 107258 141186 107494
rect 141422 107258 141464 107494
rect 141144 100494 141464 107258
rect 141144 100258 141186 100494
rect 141422 100258 141464 100494
rect 141144 93494 141464 100258
rect 141144 93258 141186 93494
rect 141422 93258 141464 93494
rect 141144 86494 141464 93258
rect 141144 86258 141186 86494
rect 141422 86258 141464 86494
rect 141144 79494 141464 86258
rect 141144 79258 141186 79494
rect 141422 79258 141464 79494
rect 141144 72494 141464 79258
rect 141144 72258 141186 72494
rect 141422 72258 141464 72494
rect 141144 65494 141464 72258
rect 141144 65258 141186 65494
rect 141422 65258 141464 65494
rect 141144 58494 141464 65258
rect 141144 58258 141186 58494
rect 141422 58258 141464 58494
rect 141144 51494 141464 58258
rect 141144 51258 141186 51494
rect 141422 51258 141464 51494
rect 141144 44494 141464 51258
rect 141144 44258 141186 44494
rect 141422 44258 141464 44494
rect 141144 37494 141464 44258
rect 141144 37258 141186 37494
rect 141422 37258 141464 37494
rect 141144 30494 141464 37258
rect 141144 30258 141186 30494
rect 141422 30258 141464 30494
rect 141144 23494 141464 30258
rect 141144 23258 141186 23494
rect 141422 23258 141464 23494
rect 141144 16494 141464 23258
rect 141144 16258 141186 16494
rect 141422 16258 141464 16494
rect 141144 9494 141464 16258
rect 141144 9258 141186 9494
rect 141422 9258 141464 9494
rect 141144 2494 141464 9258
rect 141144 2258 141186 2494
rect 141422 2258 141464 2494
rect 141144 -746 141464 2258
rect 141144 -982 141186 -746
rect 141422 -982 141464 -746
rect 141144 -1066 141464 -982
rect 141144 -1302 141186 -1066
rect 141422 -1302 141464 -1066
rect 141144 -2294 141464 -1302
rect 142876 706198 143196 706230
rect 142876 705962 142918 706198
rect 143154 705962 143196 706198
rect 142876 705878 143196 705962
rect 142876 705642 142918 705878
rect 143154 705642 143196 705878
rect 142876 696561 143196 705642
rect 142876 696325 142918 696561
rect 143154 696325 143196 696561
rect 142876 689561 143196 696325
rect 142876 689325 142918 689561
rect 143154 689325 143196 689561
rect 142876 682561 143196 689325
rect 142876 682325 142918 682561
rect 143154 682325 143196 682561
rect 142876 675561 143196 682325
rect 142876 675325 142918 675561
rect 143154 675325 143196 675561
rect 142876 668561 143196 675325
rect 142876 668325 142918 668561
rect 143154 668325 143196 668561
rect 142876 661561 143196 668325
rect 142876 661325 142918 661561
rect 143154 661325 143196 661561
rect 142876 654561 143196 661325
rect 142876 654325 142918 654561
rect 143154 654325 143196 654561
rect 142876 647561 143196 654325
rect 142876 647325 142918 647561
rect 143154 647325 143196 647561
rect 142876 640561 143196 647325
rect 142876 640325 142918 640561
rect 143154 640325 143196 640561
rect 142876 633561 143196 640325
rect 142876 633325 142918 633561
rect 143154 633325 143196 633561
rect 142876 626561 143196 633325
rect 142876 626325 142918 626561
rect 143154 626325 143196 626561
rect 142876 619561 143196 626325
rect 142876 619325 142918 619561
rect 143154 619325 143196 619561
rect 142876 612561 143196 619325
rect 142876 612325 142918 612561
rect 143154 612325 143196 612561
rect 142876 605561 143196 612325
rect 142876 605325 142918 605561
rect 143154 605325 143196 605561
rect 142876 598561 143196 605325
rect 142876 598325 142918 598561
rect 143154 598325 143196 598561
rect 142876 591561 143196 598325
rect 142876 591325 142918 591561
rect 143154 591325 143196 591561
rect 142876 584561 143196 591325
rect 142876 584325 142918 584561
rect 143154 584325 143196 584561
rect 142876 577561 143196 584325
rect 142876 577325 142918 577561
rect 143154 577325 143196 577561
rect 142876 570561 143196 577325
rect 142876 570325 142918 570561
rect 143154 570325 143196 570561
rect 142876 563561 143196 570325
rect 142876 563325 142918 563561
rect 143154 563325 143196 563561
rect 142876 556561 143196 563325
rect 142876 556325 142918 556561
rect 143154 556325 143196 556561
rect 142876 549561 143196 556325
rect 142876 549325 142918 549561
rect 143154 549325 143196 549561
rect 142876 542561 143196 549325
rect 142876 542325 142918 542561
rect 143154 542325 143196 542561
rect 142876 535561 143196 542325
rect 142876 535325 142918 535561
rect 143154 535325 143196 535561
rect 142876 528561 143196 535325
rect 142876 528325 142918 528561
rect 143154 528325 143196 528561
rect 142876 521561 143196 528325
rect 142876 521325 142918 521561
rect 143154 521325 143196 521561
rect 142876 514561 143196 521325
rect 142876 514325 142918 514561
rect 143154 514325 143196 514561
rect 142876 507561 143196 514325
rect 142876 507325 142918 507561
rect 143154 507325 143196 507561
rect 142876 500561 143196 507325
rect 142876 500325 142918 500561
rect 143154 500325 143196 500561
rect 142876 493561 143196 500325
rect 142876 493325 142918 493561
rect 143154 493325 143196 493561
rect 142876 486561 143196 493325
rect 142876 486325 142918 486561
rect 143154 486325 143196 486561
rect 142876 479561 143196 486325
rect 142876 479325 142918 479561
rect 143154 479325 143196 479561
rect 142876 472561 143196 479325
rect 142876 472325 142918 472561
rect 143154 472325 143196 472561
rect 142876 465561 143196 472325
rect 142876 465325 142918 465561
rect 143154 465325 143196 465561
rect 142876 458561 143196 465325
rect 142876 458325 142918 458561
rect 143154 458325 143196 458561
rect 142876 451561 143196 458325
rect 142876 451325 142918 451561
rect 143154 451325 143196 451561
rect 142876 444561 143196 451325
rect 142876 444325 142918 444561
rect 143154 444325 143196 444561
rect 142876 437561 143196 444325
rect 142876 437325 142918 437561
rect 143154 437325 143196 437561
rect 142876 430561 143196 437325
rect 142876 430325 142918 430561
rect 143154 430325 143196 430561
rect 142876 423561 143196 430325
rect 142876 423325 142918 423561
rect 143154 423325 143196 423561
rect 142876 416561 143196 423325
rect 142876 416325 142918 416561
rect 143154 416325 143196 416561
rect 142876 409561 143196 416325
rect 142876 409325 142918 409561
rect 143154 409325 143196 409561
rect 142876 402561 143196 409325
rect 142876 402325 142918 402561
rect 143154 402325 143196 402561
rect 142876 395561 143196 402325
rect 142876 395325 142918 395561
rect 143154 395325 143196 395561
rect 142876 388561 143196 395325
rect 142876 388325 142918 388561
rect 143154 388325 143196 388561
rect 142876 381561 143196 388325
rect 142876 381325 142918 381561
rect 143154 381325 143196 381561
rect 142876 374561 143196 381325
rect 142876 374325 142918 374561
rect 143154 374325 143196 374561
rect 142876 367561 143196 374325
rect 142876 367325 142918 367561
rect 143154 367325 143196 367561
rect 142876 360561 143196 367325
rect 142876 360325 142918 360561
rect 143154 360325 143196 360561
rect 142876 353561 143196 360325
rect 142876 353325 142918 353561
rect 143154 353325 143196 353561
rect 142876 346561 143196 353325
rect 142876 346325 142918 346561
rect 143154 346325 143196 346561
rect 142876 339561 143196 346325
rect 142876 339325 142918 339561
rect 143154 339325 143196 339561
rect 142876 332561 143196 339325
rect 142876 332325 142918 332561
rect 143154 332325 143196 332561
rect 142876 325561 143196 332325
rect 142876 325325 142918 325561
rect 143154 325325 143196 325561
rect 142876 318561 143196 325325
rect 142876 318325 142918 318561
rect 143154 318325 143196 318561
rect 142876 311561 143196 318325
rect 142876 311325 142918 311561
rect 143154 311325 143196 311561
rect 142876 304561 143196 311325
rect 142876 304325 142918 304561
rect 143154 304325 143196 304561
rect 142876 297561 143196 304325
rect 142876 297325 142918 297561
rect 143154 297325 143196 297561
rect 142876 290561 143196 297325
rect 142876 290325 142918 290561
rect 143154 290325 143196 290561
rect 142876 283561 143196 290325
rect 142876 283325 142918 283561
rect 143154 283325 143196 283561
rect 142876 276561 143196 283325
rect 142876 276325 142918 276561
rect 143154 276325 143196 276561
rect 142876 269561 143196 276325
rect 142876 269325 142918 269561
rect 143154 269325 143196 269561
rect 142876 262561 143196 269325
rect 142876 262325 142918 262561
rect 143154 262325 143196 262561
rect 142876 255561 143196 262325
rect 142876 255325 142918 255561
rect 143154 255325 143196 255561
rect 142876 248561 143196 255325
rect 142876 248325 142918 248561
rect 143154 248325 143196 248561
rect 142876 241561 143196 248325
rect 142876 241325 142918 241561
rect 143154 241325 143196 241561
rect 142876 234561 143196 241325
rect 142876 234325 142918 234561
rect 143154 234325 143196 234561
rect 142876 227561 143196 234325
rect 142876 227325 142918 227561
rect 143154 227325 143196 227561
rect 142876 220561 143196 227325
rect 142876 220325 142918 220561
rect 143154 220325 143196 220561
rect 142876 213561 143196 220325
rect 142876 213325 142918 213561
rect 143154 213325 143196 213561
rect 142876 206561 143196 213325
rect 142876 206325 142918 206561
rect 143154 206325 143196 206561
rect 142876 199561 143196 206325
rect 142876 199325 142918 199561
rect 143154 199325 143196 199561
rect 142876 192561 143196 199325
rect 142876 192325 142918 192561
rect 143154 192325 143196 192561
rect 142876 185561 143196 192325
rect 142876 185325 142918 185561
rect 143154 185325 143196 185561
rect 142876 178561 143196 185325
rect 142876 178325 142918 178561
rect 143154 178325 143196 178561
rect 142876 171561 143196 178325
rect 142876 171325 142918 171561
rect 143154 171325 143196 171561
rect 142876 164561 143196 171325
rect 142876 164325 142918 164561
rect 143154 164325 143196 164561
rect 142876 157561 143196 164325
rect 142876 157325 142918 157561
rect 143154 157325 143196 157561
rect 142876 150561 143196 157325
rect 142876 150325 142918 150561
rect 143154 150325 143196 150561
rect 142876 143561 143196 150325
rect 142876 143325 142918 143561
rect 143154 143325 143196 143561
rect 142876 136561 143196 143325
rect 142876 136325 142918 136561
rect 143154 136325 143196 136561
rect 142876 129561 143196 136325
rect 142876 129325 142918 129561
rect 143154 129325 143196 129561
rect 142876 122561 143196 129325
rect 142876 122325 142918 122561
rect 143154 122325 143196 122561
rect 142876 115561 143196 122325
rect 142876 115325 142918 115561
rect 143154 115325 143196 115561
rect 142876 108561 143196 115325
rect 142876 108325 142918 108561
rect 143154 108325 143196 108561
rect 142876 101561 143196 108325
rect 142876 101325 142918 101561
rect 143154 101325 143196 101561
rect 142876 94561 143196 101325
rect 142876 94325 142918 94561
rect 143154 94325 143196 94561
rect 142876 87561 143196 94325
rect 142876 87325 142918 87561
rect 143154 87325 143196 87561
rect 142876 80561 143196 87325
rect 142876 80325 142918 80561
rect 143154 80325 143196 80561
rect 142876 73561 143196 80325
rect 142876 73325 142918 73561
rect 143154 73325 143196 73561
rect 142876 66561 143196 73325
rect 142876 66325 142918 66561
rect 143154 66325 143196 66561
rect 142876 59561 143196 66325
rect 142876 59325 142918 59561
rect 143154 59325 143196 59561
rect 142876 52561 143196 59325
rect 142876 52325 142918 52561
rect 143154 52325 143196 52561
rect 142876 45561 143196 52325
rect 142876 45325 142918 45561
rect 143154 45325 143196 45561
rect 142876 38561 143196 45325
rect 142876 38325 142918 38561
rect 143154 38325 143196 38561
rect 142876 31561 143196 38325
rect 142876 31325 142918 31561
rect 143154 31325 143196 31561
rect 142876 24561 143196 31325
rect 142876 24325 142918 24561
rect 143154 24325 143196 24561
rect 142876 17561 143196 24325
rect 142876 17325 142918 17561
rect 143154 17325 143196 17561
rect 142876 10561 143196 17325
rect 142876 10325 142918 10561
rect 143154 10325 143196 10561
rect 142876 3561 143196 10325
rect 142876 3325 142918 3561
rect 143154 3325 143196 3561
rect 142876 -1706 143196 3325
rect 142876 -1942 142918 -1706
rect 143154 -1942 143196 -1706
rect 142876 -2026 143196 -1942
rect 142876 -2262 142918 -2026
rect 143154 -2262 143196 -2026
rect 142876 -2294 143196 -2262
rect 148144 705238 148464 706230
rect 148144 705002 148186 705238
rect 148422 705002 148464 705238
rect 148144 704918 148464 705002
rect 148144 704682 148186 704918
rect 148422 704682 148464 704918
rect 148144 695494 148464 704682
rect 148144 695258 148186 695494
rect 148422 695258 148464 695494
rect 148144 688494 148464 695258
rect 148144 688258 148186 688494
rect 148422 688258 148464 688494
rect 148144 681494 148464 688258
rect 148144 681258 148186 681494
rect 148422 681258 148464 681494
rect 148144 674494 148464 681258
rect 148144 674258 148186 674494
rect 148422 674258 148464 674494
rect 148144 667494 148464 674258
rect 148144 667258 148186 667494
rect 148422 667258 148464 667494
rect 148144 660494 148464 667258
rect 148144 660258 148186 660494
rect 148422 660258 148464 660494
rect 148144 653494 148464 660258
rect 148144 653258 148186 653494
rect 148422 653258 148464 653494
rect 148144 646494 148464 653258
rect 148144 646258 148186 646494
rect 148422 646258 148464 646494
rect 148144 639494 148464 646258
rect 148144 639258 148186 639494
rect 148422 639258 148464 639494
rect 148144 632494 148464 639258
rect 148144 632258 148186 632494
rect 148422 632258 148464 632494
rect 148144 625494 148464 632258
rect 148144 625258 148186 625494
rect 148422 625258 148464 625494
rect 148144 618494 148464 625258
rect 148144 618258 148186 618494
rect 148422 618258 148464 618494
rect 148144 611494 148464 618258
rect 148144 611258 148186 611494
rect 148422 611258 148464 611494
rect 148144 604494 148464 611258
rect 148144 604258 148186 604494
rect 148422 604258 148464 604494
rect 148144 597494 148464 604258
rect 148144 597258 148186 597494
rect 148422 597258 148464 597494
rect 148144 590494 148464 597258
rect 148144 590258 148186 590494
rect 148422 590258 148464 590494
rect 148144 583494 148464 590258
rect 148144 583258 148186 583494
rect 148422 583258 148464 583494
rect 148144 576494 148464 583258
rect 148144 576258 148186 576494
rect 148422 576258 148464 576494
rect 148144 569494 148464 576258
rect 148144 569258 148186 569494
rect 148422 569258 148464 569494
rect 148144 562494 148464 569258
rect 148144 562258 148186 562494
rect 148422 562258 148464 562494
rect 148144 555494 148464 562258
rect 148144 555258 148186 555494
rect 148422 555258 148464 555494
rect 148144 548494 148464 555258
rect 148144 548258 148186 548494
rect 148422 548258 148464 548494
rect 148144 541494 148464 548258
rect 148144 541258 148186 541494
rect 148422 541258 148464 541494
rect 148144 534494 148464 541258
rect 148144 534258 148186 534494
rect 148422 534258 148464 534494
rect 148144 527494 148464 534258
rect 148144 527258 148186 527494
rect 148422 527258 148464 527494
rect 148144 520494 148464 527258
rect 148144 520258 148186 520494
rect 148422 520258 148464 520494
rect 148144 513494 148464 520258
rect 148144 513258 148186 513494
rect 148422 513258 148464 513494
rect 148144 506494 148464 513258
rect 148144 506258 148186 506494
rect 148422 506258 148464 506494
rect 148144 499494 148464 506258
rect 148144 499258 148186 499494
rect 148422 499258 148464 499494
rect 148144 492494 148464 499258
rect 148144 492258 148186 492494
rect 148422 492258 148464 492494
rect 148144 485494 148464 492258
rect 148144 485258 148186 485494
rect 148422 485258 148464 485494
rect 148144 478494 148464 485258
rect 148144 478258 148186 478494
rect 148422 478258 148464 478494
rect 148144 471494 148464 478258
rect 148144 471258 148186 471494
rect 148422 471258 148464 471494
rect 148144 464494 148464 471258
rect 148144 464258 148186 464494
rect 148422 464258 148464 464494
rect 148144 457494 148464 464258
rect 148144 457258 148186 457494
rect 148422 457258 148464 457494
rect 148144 450494 148464 457258
rect 148144 450258 148186 450494
rect 148422 450258 148464 450494
rect 148144 443494 148464 450258
rect 148144 443258 148186 443494
rect 148422 443258 148464 443494
rect 148144 436494 148464 443258
rect 148144 436258 148186 436494
rect 148422 436258 148464 436494
rect 148144 429494 148464 436258
rect 148144 429258 148186 429494
rect 148422 429258 148464 429494
rect 148144 422494 148464 429258
rect 148144 422258 148186 422494
rect 148422 422258 148464 422494
rect 148144 415494 148464 422258
rect 148144 415258 148186 415494
rect 148422 415258 148464 415494
rect 148144 408494 148464 415258
rect 148144 408258 148186 408494
rect 148422 408258 148464 408494
rect 148144 401494 148464 408258
rect 148144 401258 148186 401494
rect 148422 401258 148464 401494
rect 148144 394494 148464 401258
rect 148144 394258 148186 394494
rect 148422 394258 148464 394494
rect 148144 387494 148464 394258
rect 148144 387258 148186 387494
rect 148422 387258 148464 387494
rect 148144 380494 148464 387258
rect 148144 380258 148186 380494
rect 148422 380258 148464 380494
rect 148144 373494 148464 380258
rect 148144 373258 148186 373494
rect 148422 373258 148464 373494
rect 148144 366494 148464 373258
rect 148144 366258 148186 366494
rect 148422 366258 148464 366494
rect 148144 359494 148464 366258
rect 148144 359258 148186 359494
rect 148422 359258 148464 359494
rect 148144 352494 148464 359258
rect 148144 352258 148186 352494
rect 148422 352258 148464 352494
rect 148144 345494 148464 352258
rect 148144 345258 148186 345494
rect 148422 345258 148464 345494
rect 148144 338494 148464 345258
rect 148144 338258 148186 338494
rect 148422 338258 148464 338494
rect 148144 331494 148464 338258
rect 148144 331258 148186 331494
rect 148422 331258 148464 331494
rect 148144 324494 148464 331258
rect 148144 324258 148186 324494
rect 148422 324258 148464 324494
rect 148144 317494 148464 324258
rect 148144 317258 148186 317494
rect 148422 317258 148464 317494
rect 148144 310494 148464 317258
rect 148144 310258 148186 310494
rect 148422 310258 148464 310494
rect 148144 303494 148464 310258
rect 148144 303258 148186 303494
rect 148422 303258 148464 303494
rect 148144 296494 148464 303258
rect 148144 296258 148186 296494
rect 148422 296258 148464 296494
rect 148144 289494 148464 296258
rect 148144 289258 148186 289494
rect 148422 289258 148464 289494
rect 148144 282494 148464 289258
rect 148144 282258 148186 282494
rect 148422 282258 148464 282494
rect 148144 275494 148464 282258
rect 148144 275258 148186 275494
rect 148422 275258 148464 275494
rect 148144 268494 148464 275258
rect 148144 268258 148186 268494
rect 148422 268258 148464 268494
rect 148144 261494 148464 268258
rect 148144 261258 148186 261494
rect 148422 261258 148464 261494
rect 148144 254494 148464 261258
rect 148144 254258 148186 254494
rect 148422 254258 148464 254494
rect 148144 247494 148464 254258
rect 148144 247258 148186 247494
rect 148422 247258 148464 247494
rect 148144 240494 148464 247258
rect 148144 240258 148186 240494
rect 148422 240258 148464 240494
rect 148144 233494 148464 240258
rect 148144 233258 148186 233494
rect 148422 233258 148464 233494
rect 148144 226494 148464 233258
rect 148144 226258 148186 226494
rect 148422 226258 148464 226494
rect 148144 219494 148464 226258
rect 148144 219258 148186 219494
rect 148422 219258 148464 219494
rect 148144 212494 148464 219258
rect 148144 212258 148186 212494
rect 148422 212258 148464 212494
rect 148144 205494 148464 212258
rect 148144 205258 148186 205494
rect 148422 205258 148464 205494
rect 148144 198494 148464 205258
rect 148144 198258 148186 198494
rect 148422 198258 148464 198494
rect 148144 191494 148464 198258
rect 148144 191258 148186 191494
rect 148422 191258 148464 191494
rect 148144 184494 148464 191258
rect 148144 184258 148186 184494
rect 148422 184258 148464 184494
rect 148144 177494 148464 184258
rect 148144 177258 148186 177494
rect 148422 177258 148464 177494
rect 148144 170494 148464 177258
rect 148144 170258 148186 170494
rect 148422 170258 148464 170494
rect 148144 163494 148464 170258
rect 148144 163258 148186 163494
rect 148422 163258 148464 163494
rect 148144 156494 148464 163258
rect 148144 156258 148186 156494
rect 148422 156258 148464 156494
rect 148144 149494 148464 156258
rect 148144 149258 148186 149494
rect 148422 149258 148464 149494
rect 148144 142494 148464 149258
rect 148144 142258 148186 142494
rect 148422 142258 148464 142494
rect 148144 135494 148464 142258
rect 148144 135258 148186 135494
rect 148422 135258 148464 135494
rect 148144 128494 148464 135258
rect 148144 128258 148186 128494
rect 148422 128258 148464 128494
rect 148144 121494 148464 128258
rect 148144 121258 148186 121494
rect 148422 121258 148464 121494
rect 148144 114494 148464 121258
rect 148144 114258 148186 114494
rect 148422 114258 148464 114494
rect 148144 107494 148464 114258
rect 148144 107258 148186 107494
rect 148422 107258 148464 107494
rect 148144 100494 148464 107258
rect 148144 100258 148186 100494
rect 148422 100258 148464 100494
rect 148144 93494 148464 100258
rect 148144 93258 148186 93494
rect 148422 93258 148464 93494
rect 148144 86494 148464 93258
rect 148144 86258 148186 86494
rect 148422 86258 148464 86494
rect 148144 79494 148464 86258
rect 148144 79258 148186 79494
rect 148422 79258 148464 79494
rect 148144 72494 148464 79258
rect 148144 72258 148186 72494
rect 148422 72258 148464 72494
rect 148144 65494 148464 72258
rect 148144 65258 148186 65494
rect 148422 65258 148464 65494
rect 148144 58494 148464 65258
rect 148144 58258 148186 58494
rect 148422 58258 148464 58494
rect 148144 51494 148464 58258
rect 148144 51258 148186 51494
rect 148422 51258 148464 51494
rect 148144 44494 148464 51258
rect 148144 44258 148186 44494
rect 148422 44258 148464 44494
rect 148144 37494 148464 44258
rect 148144 37258 148186 37494
rect 148422 37258 148464 37494
rect 148144 30494 148464 37258
rect 148144 30258 148186 30494
rect 148422 30258 148464 30494
rect 148144 23494 148464 30258
rect 148144 23258 148186 23494
rect 148422 23258 148464 23494
rect 148144 16494 148464 23258
rect 148144 16258 148186 16494
rect 148422 16258 148464 16494
rect 148144 9494 148464 16258
rect 148144 9258 148186 9494
rect 148422 9258 148464 9494
rect 148144 2494 148464 9258
rect 148144 2258 148186 2494
rect 148422 2258 148464 2494
rect 148144 -746 148464 2258
rect 148144 -982 148186 -746
rect 148422 -982 148464 -746
rect 148144 -1066 148464 -982
rect 148144 -1302 148186 -1066
rect 148422 -1302 148464 -1066
rect 148144 -2294 148464 -1302
rect 149876 706198 150196 706230
rect 149876 705962 149918 706198
rect 150154 705962 150196 706198
rect 149876 705878 150196 705962
rect 149876 705642 149918 705878
rect 150154 705642 150196 705878
rect 149876 696561 150196 705642
rect 149876 696325 149918 696561
rect 150154 696325 150196 696561
rect 149876 689561 150196 696325
rect 149876 689325 149918 689561
rect 150154 689325 150196 689561
rect 149876 682561 150196 689325
rect 149876 682325 149918 682561
rect 150154 682325 150196 682561
rect 149876 675561 150196 682325
rect 149876 675325 149918 675561
rect 150154 675325 150196 675561
rect 149876 668561 150196 675325
rect 149876 668325 149918 668561
rect 150154 668325 150196 668561
rect 149876 661561 150196 668325
rect 149876 661325 149918 661561
rect 150154 661325 150196 661561
rect 149876 654561 150196 661325
rect 149876 654325 149918 654561
rect 150154 654325 150196 654561
rect 149876 647561 150196 654325
rect 149876 647325 149918 647561
rect 150154 647325 150196 647561
rect 149876 640561 150196 647325
rect 149876 640325 149918 640561
rect 150154 640325 150196 640561
rect 149876 633561 150196 640325
rect 149876 633325 149918 633561
rect 150154 633325 150196 633561
rect 149876 626561 150196 633325
rect 149876 626325 149918 626561
rect 150154 626325 150196 626561
rect 149876 619561 150196 626325
rect 149876 619325 149918 619561
rect 150154 619325 150196 619561
rect 149876 612561 150196 619325
rect 149876 612325 149918 612561
rect 150154 612325 150196 612561
rect 149876 605561 150196 612325
rect 149876 605325 149918 605561
rect 150154 605325 150196 605561
rect 149876 598561 150196 605325
rect 149876 598325 149918 598561
rect 150154 598325 150196 598561
rect 149876 591561 150196 598325
rect 149876 591325 149918 591561
rect 150154 591325 150196 591561
rect 149876 584561 150196 591325
rect 149876 584325 149918 584561
rect 150154 584325 150196 584561
rect 149876 577561 150196 584325
rect 149876 577325 149918 577561
rect 150154 577325 150196 577561
rect 149876 570561 150196 577325
rect 149876 570325 149918 570561
rect 150154 570325 150196 570561
rect 149876 563561 150196 570325
rect 149876 563325 149918 563561
rect 150154 563325 150196 563561
rect 149876 556561 150196 563325
rect 149876 556325 149918 556561
rect 150154 556325 150196 556561
rect 149876 549561 150196 556325
rect 149876 549325 149918 549561
rect 150154 549325 150196 549561
rect 149876 542561 150196 549325
rect 149876 542325 149918 542561
rect 150154 542325 150196 542561
rect 149876 535561 150196 542325
rect 149876 535325 149918 535561
rect 150154 535325 150196 535561
rect 149876 528561 150196 535325
rect 149876 528325 149918 528561
rect 150154 528325 150196 528561
rect 149876 521561 150196 528325
rect 149876 521325 149918 521561
rect 150154 521325 150196 521561
rect 149876 514561 150196 521325
rect 149876 514325 149918 514561
rect 150154 514325 150196 514561
rect 149876 507561 150196 514325
rect 149876 507325 149918 507561
rect 150154 507325 150196 507561
rect 149876 500561 150196 507325
rect 149876 500325 149918 500561
rect 150154 500325 150196 500561
rect 149876 493561 150196 500325
rect 149876 493325 149918 493561
rect 150154 493325 150196 493561
rect 149876 486561 150196 493325
rect 149876 486325 149918 486561
rect 150154 486325 150196 486561
rect 149876 479561 150196 486325
rect 149876 479325 149918 479561
rect 150154 479325 150196 479561
rect 149876 472561 150196 479325
rect 149876 472325 149918 472561
rect 150154 472325 150196 472561
rect 149876 465561 150196 472325
rect 149876 465325 149918 465561
rect 150154 465325 150196 465561
rect 149876 458561 150196 465325
rect 149876 458325 149918 458561
rect 150154 458325 150196 458561
rect 149876 451561 150196 458325
rect 149876 451325 149918 451561
rect 150154 451325 150196 451561
rect 149876 444561 150196 451325
rect 149876 444325 149918 444561
rect 150154 444325 150196 444561
rect 149876 437561 150196 444325
rect 149876 437325 149918 437561
rect 150154 437325 150196 437561
rect 149876 430561 150196 437325
rect 149876 430325 149918 430561
rect 150154 430325 150196 430561
rect 149876 423561 150196 430325
rect 149876 423325 149918 423561
rect 150154 423325 150196 423561
rect 149876 416561 150196 423325
rect 149876 416325 149918 416561
rect 150154 416325 150196 416561
rect 149876 409561 150196 416325
rect 149876 409325 149918 409561
rect 150154 409325 150196 409561
rect 149876 402561 150196 409325
rect 149876 402325 149918 402561
rect 150154 402325 150196 402561
rect 149876 395561 150196 402325
rect 149876 395325 149918 395561
rect 150154 395325 150196 395561
rect 149876 388561 150196 395325
rect 149876 388325 149918 388561
rect 150154 388325 150196 388561
rect 149876 381561 150196 388325
rect 149876 381325 149918 381561
rect 150154 381325 150196 381561
rect 149876 374561 150196 381325
rect 149876 374325 149918 374561
rect 150154 374325 150196 374561
rect 149876 367561 150196 374325
rect 149876 367325 149918 367561
rect 150154 367325 150196 367561
rect 149876 360561 150196 367325
rect 149876 360325 149918 360561
rect 150154 360325 150196 360561
rect 149876 353561 150196 360325
rect 149876 353325 149918 353561
rect 150154 353325 150196 353561
rect 149876 346561 150196 353325
rect 149876 346325 149918 346561
rect 150154 346325 150196 346561
rect 149876 339561 150196 346325
rect 149876 339325 149918 339561
rect 150154 339325 150196 339561
rect 149876 332561 150196 339325
rect 149876 332325 149918 332561
rect 150154 332325 150196 332561
rect 149876 325561 150196 332325
rect 149876 325325 149918 325561
rect 150154 325325 150196 325561
rect 149876 318561 150196 325325
rect 149876 318325 149918 318561
rect 150154 318325 150196 318561
rect 149876 311561 150196 318325
rect 149876 311325 149918 311561
rect 150154 311325 150196 311561
rect 149876 304561 150196 311325
rect 149876 304325 149918 304561
rect 150154 304325 150196 304561
rect 149876 297561 150196 304325
rect 149876 297325 149918 297561
rect 150154 297325 150196 297561
rect 149876 290561 150196 297325
rect 149876 290325 149918 290561
rect 150154 290325 150196 290561
rect 149876 283561 150196 290325
rect 149876 283325 149918 283561
rect 150154 283325 150196 283561
rect 149876 276561 150196 283325
rect 149876 276325 149918 276561
rect 150154 276325 150196 276561
rect 149876 269561 150196 276325
rect 149876 269325 149918 269561
rect 150154 269325 150196 269561
rect 149876 262561 150196 269325
rect 149876 262325 149918 262561
rect 150154 262325 150196 262561
rect 149876 255561 150196 262325
rect 149876 255325 149918 255561
rect 150154 255325 150196 255561
rect 149876 248561 150196 255325
rect 149876 248325 149918 248561
rect 150154 248325 150196 248561
rect 149876 241561 150196 248325
rect 149876 241325 149918 241561
rect 150154 241325 150196 241561
rect 149876 234561 150196 241325
rect 149876 234325 149918 234561
rect 150154 234325 150196 234561
rect 149876 227561 150196 234325
rect 149876 227325 149918 227561
rect 150154 227325 150196 227561
rect 149876 220561 150196 227325
rect 149876 220325 149918 220561
rect 150154 220325 150196 220561
rect 149876 213561 150196 220325
rect 149876 213325 149918 213561
rect 150154 213325 150196 213561
rect 149876 206561 150196 213325
rect 149876 206325 149918 206561
rect 150154 206325 150196 206561
rect 149876 199561 150196 206325
rect 149876 199325 149918 199561
rect 150154 199325 150196 199561
rect 149876 192561 150196 199325
rect 149876 192325 149918 192561
rect 150154 192325 150196 192561
rect 149876 185561 150196 192325
rect 149876 185325 149918 185561
rect 150154 185325 150196 185561
rect 149876 178561 150196 185325
rect 149876 178325 149918 178561
rect 150154 178325 150196 178561
rect 149876 171561 150196 178325
rect 149876 171325 149918 171561
rect 150154 171325 150196 171561
rect 149876 164561 150196 171325
rect 149876 164325 149918 164561
rect 150154 164325 150196 164561
rect 149876 157561 150196 164325
rect 149876 157325 149918 157561
rect 150154 157325 150196 157561
rect 149876 150561 150196 157325
rect 149876 150325 149918 150561
rect 150154 150325 150196 150561
rect 149876 143561 150196 150325
rect 149876 143325 149918 143561
rect 150154 143325 150196 143561
rect 149876 136561 150196 143325
rect 149876 136325 149918 136561
rect 150154 136325 150196 136561
rect 149876 129561 150196 136325
rect 149876 129325 149918 129561
rect 150154 129325 150196 129561
rect 149876 122561 150196 129325
rect 149876 122325 149918 122561
rect 150154 122325 150196 122561
rect 149876 115561 150196 122325
rect 149876 115325 149918 115561
rect 150154 115325 150196 115561
rect 149876 108561 150196 115325
rect 149876 108325 149918 108561
rect 150154 108325 150196 108561
rect 149876 101561 150196 108325
rect 149876 101325 149918 101561
rect 150154 101325 150196 101561
rect 149876 94561 150196 101325
rect 149876 94325 149918 94561
rect 150154 94325 150196 94561
rect 149876 87561 150196 94325
rect 149876 87325 149918 87561
rect 150154 87325 150196 87561
rect 149876 80561 150196 87325
rect 149876 80325 149918 80561
rect 150154 80325 150196 80561
rect 149876 73561 150196 80325
rect 149876 73325 149918 73561
rect 150154 73325 150196 73561
rect 149876 66561 150196 73325
rect 149876 66325 149918 66561
rect 150154 66325 150196 66561
rect 149876 59561 150196 66325
rect 149876 59325 149918 59561
rect 150154 59325 150196 59561
rect 149876 52561 150196 59325
rect 149876 52325 149918 52561
rect 150154 52325 150196 52561
rect 149876 45561 150196 52325
rect 149876 45325 149918 45561
rect 150154 45325 150196 45561
rect 149876 38561 150196 45325
rect 149876 38325 149918 38561
rect 150154 38325 150196 38561
rect 149876 31561 150196 38325
rect 149876 31325 149918 31561
rect 150154 31325 150196 31561
rect 149876 24561 150196 31325
rect 149876 24325 149918 24561
rect 150154 24325 150196 24561
rect 149876 17561 150196 24325
rect 149876 17325 149918 17561
rect 150154 17325 150196 17561
rect 149876 10561 150196 17325
rect 149876 10325 149918 10561
rect 150154 10325 150196 10561
rect 149876 3561 150196 10325
rect 149876 3325 149918 3561
rect 150154 3325 150196 3561
rect 149876 -1706 150196 3325
rect 149876 -1942 149918 -1706
rect 150154 -1942 150196 -1706
rect 149876 -2026 150196 -1942
rect 149876 -2262 149918 -2026
rect 150154 -2262 150196 -2026
rect 149876 -2294 150196 -2262
rect 155144 705238 155464 706230
rect 155144 705002 155186 705238
rect 155422 705002 155464 705238
rect 155144 704918 155464 705002
rect 155144 704682 155186 704918
rect 155422 704682 155464 704918
rect 155144 695494 155464 704682
rect 155144 695258 155186 695494
rect 155422 695258 155464 695494
rect 155144 688494 155464 695258
rect 155144 688258 155186 688494
rect 155422 688258 155464 688494
rect 155144 681494 155464 688258
rect 155144 681258 155186 681494
rect 155422 681258 155464 681494
rect 155144 674494 155464 681258
rect 155144 674258 155186 674494
rect 155422 674258 155464 674494
rect 155144 667494 155464 674258
rect 155144 667258 155186 667494
rect 155422 667258 155464 667494
rect 155144 660494 155464 667258
rect 155144 660258 155186 660494
rect 155422 660258 155464 660494
rect 155144 653494 155464 660258
rect 155144 653258 155186 653494
rect 155422 653258 155464 653494
rect 155144 646494 155464 653258
rect 155144 646258 155186 646494
rect 155422 646258 155464 646494
rect 155144 639494 155464 646258
rect 155144 639258 155186 639494
rect 155422 639258 155464 639494
rect 155144 632494 155464 639258
rect 155144 632258 155186 632494
rect 155422 632258 155464 632494
rect 155144 625494 155464 632258
rect 155144 625258 155186 625494
rect 155422 625258 155464 625494
rect 155144 618494 155464 625258
rect 155144 618258 155186 618494
rect 155422 618258 155464 618494
rect 155144 611494 155464 618258
rect 155144 611258 155186 611494
rect 155422 611258 155464 611494
rect 155144 604494 155464 611258
rect 155144 604258 155186 604494
rect 155422 604258 155464 604494
rect 155144 597494 155464 604258
rect 155144 597258 155186 597494
rect 155422 597258 155464 597494
rect 155144 590494 155464 597258
rect 155144 590258 155186 590494
rect 155422 590258 155464 590494
rect 155144 583494 155464 590258
rect 155144 583258 155186 583494
rect 155422 583258 155464 583494
rect 155144 576494 155464 583258
rect 155144 576258 155186 576494
rect 155422 576258 155464 576494
rect 155144 569494 155464 576258
rect 155144 569258 155186 569494
rect 155422 569258 155464 569494
rect 155144 562494 155464 569258
rect 155144 562258 155186 562494
rect 155422 562258 155464 562494
rect 155144 555494 155464 562258
rect 155144 555258 155186 555494
rect 155422 555258 155464 555494
rect 155144 548494 155464 555258
rect 155144 548258 155186 548494
rect 155422 548258 155464 548494
rect 155144 541494 155464 548258
rect 155144 541258 155186 541494
rect 155422 541258 155464 541494
rect 155144 534494 155464 541258
rect 155144 534258 155186 534494
rect 155422 534258 155464 534494
rect 155144 527494 155464 534258
rect 155144 527258 155186 527494
rect 155422 527258 155464 527494
rect 155144 520494 155464 527258
rect 155144 520258 155186 520494
rect 155422 520258 155464 520494
rect 155144 513494 155464 520258
rect 155144 513258 155186 513494
rect 155422 513258 155464 513494
rect 155144 506494 155464 513258
rect 155144 506258 155186 506494
rect 155422 506258 155464 506494
rect 155144 499494 155464 506258
rect 155144 499258 155186 499494
rect 155422 499258 155464 499494
rect 155144 492494 155464 499258
rect 155144 492258 155186 492494
rect 155422 492258 155464 492494
rect 155144 485494 155464 492258
rect 155144 485258 155186 485494
rect 155422 485258 155464 485494
rect 155144 478494 155464 485258
rect 155144 478258 155186 478494
rect 155422 478258 155464 478494
rect 155144 471494 155464 478258
rect 155144 471258 155186 471494
rect 155422 471258 155464 471494
rect 155144 464494 155464 471258
rect 155144 464258 155186 464494
rect 155422 464258 155464 464494
rect 155144 457494 155464 464258
rect 155144 457258 155186 457494
rect 155422 457258 155464 457494
rect 155144 450494 155464 457258
rect 155144 450258 155186 450494
rect 155422 450258 155464 450494
rect 155144 443494 155464 450258
rect 155144 443258 155186 443494
rect 155422 443258 155464 443494
rect 155144 436494 155464 443258
rect 155144 436258 155186 436494
rect 155422 436258 155464 436494
rect 155144 429494 155464 436258
rect 155144 429258 155186 429494
rect 155422 429258 155464 429494
rect 155144 422494 155464 429258
rect 155144 422258 155186 422494
rect 155422 422258 155464 422494
rect 155144 415494 155464 422258
rect 155144 415258 155186 415494
rect 155422 415258 155464 415494
rect 155144 408494 155464 415258
rect 155144 408258 155186 408494
rect 155422 408258 155464 408494
rect 155144 401494 155464 408258
rect 155144 401258 155186 401494
rect 155422 401258 155464 401494
rect 155144 394494 155464 401258
rect 155144 394258 155186 394494
rect 155422 394258 155464 394494
rect 155144 387494 155464 394258
rect 155144 387258 155186 387494
rect 155422 387258 155464 387494
rect 155144 380494 155464 387258
rect 155144 380258 155186 380494
rect 155422 380258 155464 380494
rect 155144 373494 155464 380258
rect 155144 373258 155186 373494
rect 155422 373258 155464 373494
rect 155144 366494 155464 373258
rect 155144 366258 155186 366494
rect 155422 366258 155464 366494
rect 155144 359494 155464 366258
rect 155144 359258 155186 359494
rect 155422 359258 155464 359494
rect 155144 352494 155464 359258
rect 155144 352258 155186 352494
rect 155422 352258 155464 352494
rect 155144 345494 155464 352258
rect 155144 345258 155186 345494
rect 155422 345258 155464 345494
rect 155144 338494 155464 345258
rect 155144 338258 155186 338494
rect 155422 338258 155464 338494
rect 155144 331494 155464 338258
rect 155144 331258 155186 331494
rect 155422 331258 155464 331494
rect 155144 324494 155464 331258
rect 155144 324258 155186 324494
rect 155422 324258 155464 324494
rect 155144 317494 155464 324258
rect 155144 317258 155186 317494
rect 155422 317258 155464 317494
rect 155144 310494 155464 317258
rect 155144 310258 155186 310494
rect 155422 310258 155464 310494
rect 155144 303494 155464 310258
rect 155144 303258 155186 303494
rect 155422 303258 155464 303494
rect 155144 296494 155464 303258
rect 155144 296258 155186 296494
rect 155422 296258 155464 296494
rect 155144 289494 155464 296258
rect 155144 289258 155186 289494
rect 155422 289258 155464 289494
rect 155144 282494 155464 289258
rect 155144 282258 155186 282494
rect 155422 282258 155464 282494
rect 155144 275494 155464 282258
rect 155144 275258 155186 275494
rect 155422 275258 155464 275494
rect 155144 268494 155464 275258
rect 155144 268258 155186 268494
rect 155422 268258 155464 268494
rect 155144 261494 155464 268258
rect 155144 261258 155186 261494
rect 155422 261258 155464 261494
rect 155144 254494 155464 261258
rect 155144 254258 155186 254494
rect 155422 254258 155464 254494
rect 155144 247494 155464 254258
rect 155144 247258 155186 247494
rect 155422 247258 155464 247494
rect 155144 240494 155464 247258
rect 155144 240258 155186 240494
rect 155422 240258 155464 240494
rect 155144 233494 155464 240258
rect 155144 233258 155186 233494
rect 155422 233258 155464 233494
rect 155144 226494 155464 233258
rect 155144 226258 155186 226494
rect 155422 226258 155464 226494
rect 155144 219494 155464 226258
rect 155144 219258 155186 219494
rect 155422 219258 155464 219494
rect 155144 212494 155464 219258
rect 155144 212258 155186 212494
rect 155422 212258 155464 212494
rect 155144 205494 155464 212258
rect 155144 205258 155186 205494
rect 155422 205258 155464 205494
rect 155144 198494 155464 205258
rect 155144 198258 155186 198494
rect 155422 198258 155464 198494
rect 155144 191494 155464 198258
rect 155144 191258 155186 191494
rect 155422 191258 155464 191494
rect 155144 184494 155464 191258
rect 155144 184258 155186 184494
rect 155422 184258 155464 184494
rect 155144 177494 155464 184258
rect 155144 177258 155186 177494
rect 155422 177258 155464 177494
rect 155144 170494 155464 177258
rect 155144 170258 155186 170494
rect 155422 170258 155464 170494
rect 155144 163494 155464 170258
rect 155144 163258 155186 163494
rect 155422 163258 155464 163494
rect 155144 156494 155464 163258
rect 155144 156258 155186 156494
rect 155422 156258 155464 156494
rect 155144 149494 155464 156258
rect 155144 149258 155186 149494
rect 155422 149258 155464 149494
rect 155144 142494 155464 149258
rect 155144 142258 155186 142494
rect 155422 142258 155464 142494
rect 155144 135494 155464 142258
rect 155144 135258 155186 135494
rect 155422 135258 155464 135494
rect 155144 128494 155464 135258
rect 155144 128258 155186 128494
rect 155422 128258 155464 128494
rect 155144 121494 155464 128258
rect 155144 121258 155186 121494
rect 155422 121258 155464 121494
rect 155144 114494 155464 121258
rect 155144 114258 155186 114494
rect 155422 114258 155464 114494
rect 155144 107494 155464 114258
rect 155144 107258 155186 107494
rect 155422 107258 155464 107494
rect 155144 100494 155464 107258
rect 155144 100258 155186 100494
rect 155422 100258 155464 100494
rect 155144 93494 155464 100258
rect 155144 93258 155186 93494
rect 155422 93258 155464 93494
rect 155144 86494 155464 93258
rect 155144 86258 155186 86494
rect 155422 86258 155464 86494
rect 155144 79494 155464 86258
rect 155144 79258 155186 79494
rect 155422 79258 155464 79494
rect 155144 72494 155464 79258
rect 155144 72258 155186 72494
rect 155422 72258 155464 72494
rect 155144 65494 155464 72258
rect 155144 65258 155186 65494
rect 155422 65258 155464 65494
rect 155144 58494 155464 65258
rect 155144 58258 155186 58494
rect 155422 58258 155464 58494
rect 155144 51494 155464 58258
rect 155144 51258 155186 51494
rect 155422 51258 155464 51494
rect 155144 44494 155464 51258
rect 155144 44258 155186 44494
rect 155422 44258 155464 44494
rect 155144 37494 155464 44258
rect 155144 37258 155186 37494
rect 155422 37258 155464 37494
rect 155144 30494 155464 37258
rect 155144 30258 155186 30494
rect 155422 30258 155464 30494
rect 155144 23494 155464 30258
rect 155144 23258 155186 23494
rect 155422 23258 155464 23494
rect 155144 16494 155464 23258
rect 155144 16258 155186 16494
rect 155422 16258 155464 16494
rect 155144 9494 155464 16258
rect 155144 9258 155186 9494
rect 155422 9258 155464 9494
rect 155144 2494 155464 9258
rect 155144 2258 155186 2494
rect 155422 2258 155464 2494
rect 155144 -746 155464 2258
rect 155144 -982 155186 -746
rect 155422 -982 155464 -746
rect 155144 -1066 155464 -982
rect 155144 -1302 155186 -1066
rect 155422 -1302 155464 -1066
rect 155144 -2294 155464 -1302
rect 156876 706198 157196 706230
rect 156876 705962 156918 706198
rect 157154 705962 157196 706198
rect 156876 705878 157196 705962
rect 156876 705642 156918 705878
rect 157154 705642 157196 705878
rect 156876 696561 157196 705642
rect 156876 696325 156918 696561
rect 157154 696325 157196 696561
rect 156876 689561 157196 696325
rect 156876 689325 156918 689561
rect 157154 689325 157196 689561
rect 156876 682561 157196 689325
rect 156876 682325 156918 682561
rect 157154 682325 157196 682561
rect 156876 675561 157196 682325
rect 156876 675325 156918 675561
rect 157154 675325 157196 675561
rect 156876 668561 157196 675325
rect 156876 668325 156918 668561
rect 157154 668325 157196 668561
rect 156876 661561 157196 668325
rect 156876 661325 156918 661561
rect 157154 661325 157196 661561
rect 156876 654561 157196 661325
rect 156876 654325 156918 654561
rect 157154 654325 157196 654561
rect 156876 647561 157196 654325
rect 156876 647325 156918 647561
rect 157154 647325 157196 647561
rect 156876 640561 157196 647325
rect 156876 640325 156918 640561
rect 157154 640325 157196 640561
rect 156876 633561 157196 640325
rect 156876 633325 156918 633561
rect 157154 633325 157196 633561
rect 156876 626561 157196 633325
rect 156876 626325 156918 626561
rect 157154 626325 157196 626561
rect 156876 619561 157196 626325
rect 156876 619325 156918 619561
rect 157154 619325 157196 619561
rect 156876 612561 157196 619325
rect 156876 612325 156918 612561
rect 157154 612325 157196 612561
rect 156876 605561 157196 612325
rect 156876 605325 156918 605561
rect 157154 605325 157196 605561
rect 156876 598561 157196 605325
rect 156876 598325 156918 598561
rect 157154 598325 157196 598561
rect 156876 591561 157196 598325
rect 156876 591325 156918 591561
rect 157154 591325 157196 591561
rect 156876 584561 157196 591325
rect 156876 584325 156918 584561
rect 157154 584325 157196 584561
rect 156876 577561 157196 584325
rect 156876 577325 156918 577561
rect 157154 577325 157196 577561
rect 156876 570561 157196 577325
rect 156876 570325 156918 570561
rect 157154 570325 157196 570561
rect 156876 563561 157196 570325
rect 156876 563325 156918 563561
rect 157154 563325 157196 563561
rect 156876 556561 157196 563325
rect 156876 556325 156918 556561
rect 157154 556325 157196 556561
rect 156876 549561 157196 556325
rect 156876 549325 156918 549561
rect 157154 549325 157196 549561
rect 156876 542561 157196 549325
rect 156876 542325 156918 542561
rect 157154 542325 157196 542561
rect 156876 535561 157196 542325
rect 156876 535325 156918 535561
rect 157154 535325 157196 535561
rect 156876 528561 157196 535325
rect 156876 528325 156918 528561
rect 157154 528325 157196 528561
rect 156876 521561 157196 528325
rect 156876 521325 156918 521561
rect 157154 521325 157196 521561
rect 156876 514561 157196 521325
rect 156876 514325 156918 514561
rect 157154 514325 157196 514561
rect 156876 507561 157196 514325
rect 156876 507325 156918 507561
rect 157154 507325 157196 507561
rect 156876 500561 157196 507325
rect 156876 500325 156918 500561
rect 157154 500325 157196 500561
rect 156876 493561 157196 500325
rect 156876 493325 156918 493561
rect 157154 493325 157196 493561
rect 156876 486561 157196 493325
rect 156876 486325 156918 486561
rect 157154 486325 157196 486561
rect 156876 479561 157196 486325
rect 156876 479325 156918 479561
rect 157154 479325 157196 479561
rect 156876 472561 157196 479325
rect 156876 472325 156918 472561
rect 157154 472325 157196 472561
rect 156876 465561 157196 472325
rect 156876 465325 156918 465561
rect 157154 465325 157196 465561
rect 156876 458561 157196 465325
rect 156876 458325 156918 458561
rect 157154 458325 157196 458561
rect 156876 451561 157196 458325
rect 156876 451325 156918 451561
rect 157154 451325 157196 451561
rect 156876 444561 157196 451325
rect 156876 444325 156918 444561
rect 157154 444325 157196 444561
rect 156876 437561 157196 444325
rect 156876 437325 156918 437561
rect 157154 437325 157196 437561
rect 156876 430561 157196 437325
rect 156876 430325 156918 430561
rect 157154 430325 157196 430561
rect 156876 423561 157196 430325
rect 156876 423325 156918 423561
rect 157154 423325 157196 423561
rect 156876 416561 157196 423325
rect 156876 416325 156918 416561
rect 157154 416325 157196 416561
rect 156876 409561 157196 416325
rect 156876 409325 156918 409561
rect 157154 409325 157196 409561
rect 156876 402561 157196 409325
rect 156876 402325 156918 402561
rect 157154 402325 157196 402561
rect 156876 395561 157196 402325
rect 156876 395325 156918 395561
rect 157154 395325 157196 395561
rect 156876 388561 157196 395325
rect 156876 388325 156918 388561
rect 157154 388325 157196 388561
rect 156876 381561 157196 388325
rect 156876 381325 156918 381561
rect 157154 381325 157196 381561
rect 156876 374561 157196 381325
rect 156876 374325 156918 374561
rect 157154 374325 157196 374561
rect 156876 367561 157196 374325
rect 156876 367325 156918 367561
rect 157154 367325 157196 367561
rect 156876 360561 157196 367325
rect 156876 360325 156918 360561
rect 157154 360325 157196 360561
rect 156876 353561 157196 360325
rect 156876 353325 156918 353561
rect 157154 353325 157196 353561
rect 156876 346561 157196 353325
rect 156876 346325 156918 346561
rect 157154 346325 157196 346561
rect 156876 339561 157196 346325
rect 156876 339325 156918 339561
rect 157154 339325 157196 339561
rect 156876 332561 157196 339325
rect 156876 332325 156918 332561
rect 157154 332325 157196 332561
rect 156876 325561 157196 332325
rect 156876 325325 156918 325561
rect 157154 325325 157196 325561
rect 156876 318561 157196 325325
rect 156876 318325 156918 318561
rect 157154 318325 157196 318561
rect 156876 311561 157196 318325
rect 156876 311325 156918 311561
rect 157154 311325 157196 311561
rect 156876 304561 157196 311325
rect 156876 304325 156918 304561
rect 157154 304325 157196 304561
rect 156876 297561 157196 304325
rect 156876 297325 156918 297561
rect 157154 297325 157196 297561
rect 156876 290561 157196 297325
rect 156876 290325 156918 290561
rect 157154 290325 157196 290561
rect 156876 283561 157196 290325
rect 156876 283325 156918 283561
rect 157154 283325 157196 283561
rect 156876 276561 157196 283325
rect 156876 276325 156918 276561
rect 157154 276325 157196 276561
rect 156876 269561 157196 276325
rect 156876 269325 156918 269561
rect 157154 269325 157196 269561
rect 156876 262561 157196 269325
rect 156876 262325 156918 262561
rect 157154 262325 157196 262561
rect 156876 255561 157196 262325
rect 156876 255325 156918 255561
rect 157154 255325 157196 255561
rect 156876 248561 157196 255325
rect 156876 248325 156918 248561
rect 157154 248325 157196 248561
rect 156876 241561 157196 248325
rect 156876 241325 156918 241561
rect 157154 241325 157196 241561
rect 156876 234561 157196 241325
rect 156876 234325 156918 234561
rect 157154 234325 157196 234561
rect 156876 227561 157196 234325
rect 156876 227325 156918 227561
rect 157154 227325 157196 227561
rect 156876 220561 157196 227325
rect 156876 220325 156918 220561
rect 157154 220325 157196 220561
rect 156876 213561 157196 220325
rect 156876 213325 156918 213561
rect 157154 213325 157196 213561
rect 156876 206561 157196 213325
rect 156876 206325 156918 206561
rect 157154 206325 157196 206561
rect 156876 199561 157196 206325
rect 156876 199325 156918 199561
rect 157154 199325 157196 199561
rect 156876 192561 157196 199325
rect 156876 192325 156918 192561
rect 157154 192325 157196 192561
rect 156876 185561 157196 192325
rect 156876 185325 156918 185561
rect 157154 185325 157196 185561
rect 156876 178561 157196 185325
rect 156876 178325 156918 178561
rect 157154 178325 157196 178561
rect 156876 171561 157196 178325
rect 156876 171325 156918 171561
rect 157154 171325 157196 171561
rect 156876 164561 157196 171325
rect 156876 164325 156918 164561
rect 157154 164325 157196 164561
rect 156876 157561 157196 164325
rect 156876 157325 156918 157561
rect 157154 157325 157196 157561
rect 156876 150561 157196 157325
rect 156876 150325 156918 150561
rect 157154 150325 157196 150561
rect 156876 143561 157196 150325
rect 156876 143325 156918 143561
rect 157154 143325 157196 143561
rect 156876 136561 157196 143325
rect 156876 136325 156918 136561
rect 157154 136325 157196 136561
rect 156876 129561 157196 136325
rect 156876 129325 156918 129561
rect 157154 129325 157196 129561
rect 156876 122561 157196 129325
rect 156876 122325 156918 122561
rect 157154 122325 157196 122561
rect 156876 115561 157196 122325
rect 156876 115325 156918 115561
rect 157154 115325 157196 115561
rect 156876 108561 157196 115325
rect 156876 108325 156918 108561
rect 157154 108325 157196 108561
rect 156876 101561 157196 108325
rect 156876 101325 156918 101561
rect 157154 101325 157196 101561
rect 156876 94561 157196 101325
rect 156876 94325 156918 94561
rect 157154 94325 157196 94561
rect 156876 87561 157196 94325
rect 156876 87325 156918 87561
rect 157154 87325 157196 87561
rect 156876 80561 157196 87325
rect 156876 80325 156918 80561
rect 157154 80325 157196 80561
rect 156876 73561 157196 80325
rect 156876 73325 156918 73561
rect 157154 73325 157196 73561
rect 156876 66561 157196 73325
rect 156876 66325 156918 66561
rect 157154 66325 157196 66561
rect 156876 59561 157196 66325
rect 156876 59325 156918 59561
rect 157154 59325 157196 59561
rect 156876 52561 157196 59325
rect 156876 52325 156918 52561
rect 157154 52325 157196 52561
rect 156876 45561 157196 52325
rect 156876 45325 156918 45561
rect 157154 45325 157196 45561
rect 156876 38561 157196 45325
rect 156876 38325 156918 38561
rect 157154 38325 157196 38561
rect 156876 31561 157196 38325
rect 156876 31325 156918 31561
rect 157154 31325 157196 31561
rect 156876 24561 157196 31325
rect 156876 24325 156918 24561
rect 157154 24325 157196 24561
rect 156876 17561 157196 24325
rect 156876 17325 156918 17561
rect 157154 17325 157196 17561
rect 156876 10561 157196 17325
rect 156876 10325 156918 10561
rect 157154 10325 157196 10561
rect 156876 3561 157196 10325
rect 156876 3325 156918 3561
rect 157154 3325 157196 3561
rect 156876 -1706 157196 3325
rect 156876 -1942 156918 -1706
rect 157154 -1942 157196 -1706
rect 156876 -2026 157196 -1942
rect 156876 -2262 156918 -2026
rect 157154 -2262 157196 -2026
rect 156876 -2294 157196 -2262
rect 162144 705238 162464 706230
rect 162144 705002 162186 705238
rect 162422 705002 162464 705238
rect 162144 704918 162464 705002
rect 162144 704682 162186 704918
rect 162422 704682 162464 704918
rect 162144 695494 162464 704682
rect 162144 695258 162186 695494
rect 162422 695258 162464 695494
rect 162144 688494 162464 695258
rect 162144 688258 162186 688494
rect 162422 688258 162464 688494
rect 162144 681494 162464 688258
rect 162144 681258 162186 681494
rect 162422 681258 162464 681494
rect 162144 674494 162464 681258
rect 162144 674258 162186 674494
rect 162422 674258 162464 674494
rect 162144 667494 162464 674258
rect 162144 667258 162186 667494
rect 162422 667258 162464 667494
rect 162144 660494 162464 667258
rect 162144 660258 162186 660494
rect 162422 660258 162464 660494
rect 162144 653494 162464 660258
rect 162144 653258 162186 653494
rect 162422 653258 162464 653494
rect 162144 646494 162464 653258
rect 162144 646258 162186 646494
rect 162422 646258 162464 646494
rect 162144 639494 162464 646258
rect 162144 639258 162186 639494
rect 162422 639258 162464 639494
rect 162144 632494 162464 639258
rect 162144 632258 162186 632494
rect 162422 632258 162464 632494
rect 162144 625494 162464 632258
rect 162144 625258 162186 625494
rect 162422 625258 162464 625494
rect 162144 618494 162464 625258
rect 162144 618258 162186 618494
rect 162422 618258 162464 618494
rect 162144 611494 162464 618258
rect 162144 611258 162186 611494
rect 162422 611258 162464 611494
rect 162144 604494 162464 611258
rect 162144 604258 162186 604494
rect 162422 604258 162464 604494
rect 162144 597494 162464 604258
rect 162144 597258 162186 597494
rect 162422 597258 162464 597494
rect 162144 590494 162464 597258
rect 162144 590258 162186 590494
rect 162422 590258 162464 590494
rect 162144 583494 162464 590258
rect 162144 583258 162186 583494
rect 162422 583258 162464 583494
rect 162144 576494 162464 583258
rect 162144 576258 162186 576494
rect 162422 576258 162464 576494
rect 162144 569494 162464 576258
rect 162144 569258 162186 569494
rect 162422 569258 162464 569494
rect 162144 562494 162464 569258
rect 162144 562258 162186 562494
rect 162422 562258 162464 562494
rect 162144 555494 162464 562258
rect 162144 555258 162186 555494
rect 162422 555258 162464 555494
rect 162144 548494 162464 555258
rect 162144 548258 162186 548494
rect 162422 548258 162464 548494
rect 162144 541494 162464 548258
rect 162144 541258 162186 541494
rect 162422 541258 162464 541494
rect 162144 534494 162464 541258
rect 162144 534258 162186 534494
rect 162422 534258 162464 534494
rect 162144 527494 162464 534258
rect 162144 527258 162186 527494
rect 162422 527258 162464 527494
rect 162144 520494 162464 527258
rect 162144 520258 162186 520494
rect 162422 520258 162464 520494
rect 162144 513494 162464 520258
rect 162144 513258 162186 513494
rect 162422 513258 162464 513494
rect 162144 506494 162464 513258
rect 162144 506258 162186 506494
rect 162422 506258 162464 506494
rect 162144 499494 162464 506258
rect 162144 499258 162186 499494
rect 162422 499258 162464 499494
rect 162144 492494 162464 499258
rect 162144 492258 162186 492494
rect 162422 492258 162464 492494
rect 162144 485494 162464 492258
rect 162144 485258 162186 485494
rect 162422 485258 162464 485494
rect 162144 478494 162464 485258
rect 162144 478258 162186 478494
rect 162422 478258 162464 478494
rect 162144 471494 162464 478258
rect 162144 471258 162186 471494
rect 162422 471258 162464 471494
rect 162144 464494 162464 471258
rect 162144 464258 162186 464494
rect 162422 464258 162464 464494
rect 162144 457494 162464 464258
rect 162144 457258 162186 457494
rect 162422 457258 162464 457494
rect 162144 450494 162464 457258
rect 162144 450258 162186 450494
rect 162422 450258 162464 450494
rect 162144 443494 162464 450258
rect 162144 443258 162186 443494
rect 162422 443258 162464 443494
rect 162144 436494 162464 443258
rect 162144 436258 162186 436494
rect 162422 436258 162464 436494
rect 162144 429494 162464 436258
rect 162144 429258 162186 429494
rect 162422 429258 162464 429494
rect 162144 422494 162464 429258
rect 162144 422258 162186 422494
rect 162422 422258 162464 422494
rect 162144 415494 162464 422258
rect 162144 415258 162186 415494
rect 162422 415258 162464 415494
rect 162144 408494 162464 415258
rect 162144 408258 162186 408494
rect 162422 408258 162464 408494
rect 162144 401494 162464 408258
rect 162144 401258 162186 401494
rect 162422 401258 162464 401494
rect 162144 394494 162464 401258
rect 162144 394258 162186 394494
rect 162422 394258 162464 394494
rect 162144 387494 162464 394258
rect 162144 387258 162186 387494
rect 162422 387258 162464 387494
rect 162144 380494 162464 387258
rect 162144 380258 162186 380494
rect 162422 380258 162464 380494
rect 162144 373494 162464 380258
rect 162144 373258 162186 373494
rect 162422 373258 162464 373494
rect 162144 366494 162464 373258
rect 162144 366258 162186 366494
rect 162422 366258 162464 366494
rect 162144 359494 162464 366258
rect 162144 359258 162186 359494
rect 162422 359258 162464 359494
rect 162144 352494 162464 359258
rect 162144 352258 162186 352494
rect 162422 352258 162464 352494
rect 162144 345494 162464 352258
rect 162144 345258 162186 345494
rect 162422 345258 162464 345494
rect 162144 338494 162464 345258
rect 162144 338258 162186 338494
rect 162422 338258 162464 338494
rect 162144 331494 162464 338258
rect 162144 331258 162186 331494
rect 162422 331258 162464 331494
rect 162144 324494 162464 331258
rect 162144 324258 162186 324494
rect 162422 324258 162464 324494
rect 162144 317494 162464 324258
rect 162144 317258 162186 317494
rect 162422 317258 162464 317494
rect 162144 310494 162464 317258
rect 162144 310258 162186 310494
rect 162422 310258 162464 310494
rect 162144 303494 162464 310258
rect 162144 303258 162186 303494
rect 162422 303258 162464 303494
rect 162144 296494 162464 303258
rect 162144 296258 162186 296494
rect 162422 296258 162464 296494
rect 162144 289494 162464 296258
rect 162144 289258 162186 289494
rect 162422 289258 162464 289494
rect 162144 282494 162464 289258
rect 162144 282258 162186 282494
rect 162422 282258 162464 282494
rect 162144 275494 162464 282258
rect 162144 275258 162186 275494
rect 162422 275258 162464 275494
rect 162144 268494 162464 275258
rect 162144 268258 162186 268494
rect 162422 268258 162464 268494
rect 162144 261494 162464 268258
rect 162144 261258 162186 261494
rect 162422 261258 162464 261494
rect 162144 254494 162464 261258
rect 162144 254258 162186 254494
rect 162422 254258 162464 254494
rect 162144 247494 162464 254258
rect 162144 247258 162186 247494
rect 162422 247258 162464 247494
rect 162144 240494 162464 247258
rect 162144 240258 162186 240494
rect 162422 240258 162464 240494
rect 162144 233494 162464 240258
rect 162144 233258 162186 233494
rect 162422 233258 162464 233494
rect 162144 226494 162464 233258
rect 162144 226258 162186 226494
rect 162422 226258 162464 226494
rect 162144 219494 162464 226258
rect 162144 219258 162186 219494
rect 162422 219258 162464 219494
rect 162144 212494 162464 219258
rect 162144 212258 162186 212494
rect 162422 212258 162464 212494
rect 162144 205494 162464 212258
rect 162144 205258 162186 205494
rect 162422 205258 162464 205494
rect 162144 198494 162464 205258
rect 162144 198258 162186 198494
rect 162422 198258 162464 198494
rect 162144 191494 162464 198258
rect 162144 191258 162186 191494
rect 162422 191258 162464 191494
rect 162144 184494 162464 191258
rect 162144 184258 162186 184494
rect 162422 184258 162464 184494
rect 162144 177494 162464 184258
rect 162144 177258 162186 177494
rect 162422 177258 162464 177494
rect 162144 170494 162464 177258
rect 162144 170258 162186 170494
rect 162422 170258 162464 170494
rect 162144 163494 162464 170258
rect 162144 163258 162186 163494
rect 162422 163258 162464 163494
rect 162144 156494 162464 163258
rect 162144 156258 162186 156494
rect 162422 156258 162464 156494
rect 162144 149494 162464 156258
rect 162144 149258 162186 149494
rect 162422 149258 162464 149494
rect 162144 142494 162464 149258
rect 162144 142258 162186 142494
rect 162422 142258 162464 142494
rect 162144 135494 162464 142258
rect 162144 135258 162186 135494
rect 162422 135258 162464 135494
rect 162144 128494 162464 135258
rect 162144 128258 162186 128494
rect 162422 128258 162464 128494
rect 162144 121494 162464 128258
rect 162144 121258 162186 121494
rect 162422 121258 162464 121494
rect 162144 114494 162464 121258
rect 162144 114258 162186 114494
rect 162422 114258 162464 114494
rect 162144 107494 162464 114258
rect 162144 107258 162186 107494
rect 162422 107258 162464 107494
rect 162144 100494 162464 107258
rect 162144 100258 162186 100494
rect 162422 100258 162464 100494
rect 162144 93494 162464 100258
rect 162144 93258 162186 93494
rect 162422 93258 162464 93494
rect 162144 86494 162464 93258
rect 162144 86258 162186 86494
rect 162422 86258 162464 86494
rect 162144 79494 162464 86258
rect 162144 79258 162186 79494
rect 162422 79258 162464 79494
rect 162144 72494 162464 79258
rect 162144 72258 162186 72494
rect 162422 72258 162464 72494
rect 162144 65494 162464 72258
rect 162144 65258 162186 65494
rect 162422 65258 162464 65494
rect 162144 58494 162464 65258
rect 162144 58258 162186 58494
rect 162422 58258 162464 58494
rect 162144 51494 162464 58258
rect 162144 51258 162186 51494
rect 162422 51258 162464 51494
rect 162144 44494 162464 51258
rect 162144 44258 162186 44494
rect 162422 44258 162464 44494
rect 162144 37494 162464 44258
rect 162144 37258 162186 37494
rect 162422 37258 162464 37494
rect 162144 30494 162464 37258
rect 162144 30258 162186 30494
rect 162422 30258 162464 30494
rect 162144 23494 162464 30258
rect 162144 23258 162186 23494
rect 162422 23258 162464 23494
rect 162144 16494 162464 23258
rect 162144 16258 162186 16494
rect 162422 16258 162464 16494
rect 162144 9494 162464 16258
rect 162144 9258 162186 9494
rect 162422 9258 162464 9494
rect 162144 2494 162464 9258
rect 162144 2258 162186 2494
rect 162422 2258 162464 2494
rect 162144 -746 162464 2258
rect 162144 -982 162186 -746
rect 162422 -982 162464 -746
rect 162144 -1066 162464 -982
rect 162144 -1302 162186 -1066
rect 162422 -1302 162464 -1066
rect 162144 -2294 162464 -1302
rect 163876 706198 164196 706230
rect 163876 705962 163918 706198
rect 164154 705962 164196 706198
rect 163876 705878 164196 705962
rect 163876 705642 163918 705878
rect 164154 705642 164196 705878
rect 163876 696561 164196 705642
rect 163876 696325 163918 696561
rect 164154 696325 164196 696561
rect 163876 689561 164196 696325
rect 163876 689325 163918 689561
rect 164154 689325 164196 689561
rect 163876 682561 164196 689325
rect 163876 682325 163918 682561
rect 164154 682325 164196 682561
rect 163876 675561 164196 682325
rect 163876 675325 163918 675561
rect 164154 675325 164196 675561
rect 163876 668561 164196 675325
rect 163876 668325 163918 668561
rect 164154 668325 164196 668561
rect 163876 661561 164196 668325
rect 163876 661325 163918 661561
rect 164154 661325 164196 661561
rect 163876 654561 164196 661325
rect 163876 654325 163918 654561
rect 164154 654325 164196 654561
rect 163876 647561 164196 654325
rect 163876 647325 163918 647561
rect 164154 647325 164196 647561
rect 163876 640561 164196 647325
rect 163876 640325 163918 640561
rect 164154 640325 164196 640561
rect 163876 633561 164196 640325
rect 163876 633325 163918 633561
rect 164154 633325 164196 633561
rect 163876 626561 164196 633325
rect 163876 626325 163918 626561
rect 164154 626325 164196 626561
rect 163876 619561 164196 626325
rect 163876 619325 163918 619561
rect 164154 619325 164196 619561
rect 163876 612561 164196 619325
rect 163876 612325 163918 612561
rect 164154 612325 164196 612561
rect 163876 605561 164196 612325
rect 163876 605325 163918 605561
rect 164154 605325 164196 605561
rect 163876 598561 164196 605325
rect 163876 598325 163918 598561
rect 164154 598325 164196 598561
rect 163876 591561 164196 598325
rect 163876 591325 163918 591561
rect 164154 591325 164196 591561
rect 163876 584561 164196 591325
rect 163876 584325 163918 584561
rect 164154 584325 164196 584561
rect 163876 577561 164196 584325
rect 163876 577325 163918 577561
rect 164154 577325 164196 577561
rect 163876 570561 164196 577325
rect 163876 570325 163918 570561
rect 164154 570325 164196 570561
rect 163876 563561 164196 570325
rect 163876 563325 163918 563561
rect 164154 563325 164196 563561
rect 163876 556561 164196 563325
rect 163876 556325 163918 556561
rect 164154 556325 164196 556561
rect 163876 549561 164196 556325
rect 163876 549325 163918 549561
rect 164154 549325 164196 549561
rect 163876 542561 164196 549325
rect 163876 542325 163918 542561
rect 164154 542325 164196 542561
rect 163876 535561 164196 542325
rect 163876 535325 163918 535561
rect 164154 535325 164196 535561
rect 163876 528561 164196 535325
rect 163876 528325 163918 528561
rect 164154 528325 164196 528561
rect 163876 521561 164196 528325
rect 163876 521325 163918 521561
rect 164154 521325 164196 521561
rect 163876 514561 164196 521325
rect 163876 514325 163918 514561
rect 164154 514325 164196 514561
rect 163876 507561 164196 514325
rect 163876 507325 163918 507561
rect 164154 507325 164196 507561
rect 163876 500561 164196 507325
rect 163876 500325 163918 500561
rect 164154 500325 164196 500561
rect 163876 493561 164196 500325
rect 163876 493325 163918 493561
rect 164154 493325 164196 493561
rect 163876 486561 164196 493325
rect 163876 486325 163918 486561
rect 164154 486325 164196 486561
rect 163876 479561 164196 486325
rect 163876 479325 163918 479561
rect 164154 479325 164196 479561
rect 163876 472561 164196 479325
rect 163876 472325 163918 472561
rect 164154 472325 164196 472561
rect 163876 465561 164196 472325
rect 163876 465325 163918 465561
rect 164154 465325 164196 465561
rect 163876 458561 164196 465325
rect 163876 458325 163918 458561
rect 164154 458325 164196 458561
rect 163876 451561 164196 458325
rect 163876 451325 163918 451561
rect 164154 451325 164196 451561
rect 163876 444561 164196 451325
rect 163876 444325 163918 444561
rect 164154 444325 164196 444561
rect 163876 437561 164196 444325
rect 163876 437325 163918 437561
rect 164154 437325 164196 437561
rect 163876 430561 164196 437325
rect 163876 430325 163918 430561
rect 164154 430325 164196 430561
rect 163876 423561 164196 430325
rect 163876 423325 163918 423561
rect 164154 423325 164196 423561
rect 163876 416561 164196 423325
rect 163876 416325 163918 416561
rect 164154 416325 164196 416561
rect 163876 409561 164196 416325
rect 163876 409325 163918 409561
rect 164154 409325 164196 409561
rect 163876 402561 164196 409325
rect 163876 402325 163918 402561
rect 164154 402325 164196 402561
rect 163876 395561 164196 402325
rect 163876 395325 163918 395561
rect 164154 395325 164196 395561
rect 163876 388561 164196 395325
rect 163876 388325 163918 388561
rect 164154 388325 164196 388561
rect 163876 381561 164196 388325
rect 163876 381325 163918 381561
rect 164154 381325 164196 381561
rect 163876 374561 164196 381325
rect 163876 374325 163918 374561
rect 164154 374325 164196 374561
rect 163876 367561 164196 374325
rect 163876 367325 163918 367561
rect 164154 367325 164196 367561
rect 163876 360561 164196 367325
rect 163876 360325 163918 360561
rect 164154 360325 164196 360561
rect 163876 353561 164196 360325
rect 163876 353325 163918 353561
rect 164154 353325 164196 353561
rect 163876 346561 164196 353325
rect 163876 346325 163918 346561
rect 164154 346325 164196 346561
rect 163876 339561 164196 346325
rect 163876 339325 163918 339561
rect 164154 339325 164196 339561
rect 163876 332561 164196 339325
rect 163876 332325 163918 332561
rect 164154 332325 164196 332561
rect 163876 325561 164196 332325
rect 163876 325325 163918 325561
rect 164154 325325 164196 325561
rect 163876 318561 164196 325325
rect 163876 318325 163918 318561
rect 164154 318325 164196 318561
rect 163876 311561 164196 318325
rect 163876 311325 163918 311561
rect 164154 311325 164196 311561
rect 163876 304561 164196 311325
rect 163876 304325 163918 304561
rect 164154 304325 164196 304561
rect 163876 297561 164196 304325
rect 163876 297325 163918 297561
rect 164154 297325 164196 297561
rect 163876 290561 164196 297325
rect 163876 290325 163918 290561
rect 164154 290325 164196 290561
rect 163876 283561 164196 290325
rect 163876 283325 163918 283561
rect 164154 283325 164196 283561
rect 163876 276561 164196 283325
rect 163876 276325 163918 276561
rect 164154 276325 164196 276561
rect 163876 269561 164196 276325
rect 163876 269325 163918 269561
rect 164154 269325 164196 269561
rect 163876 262561 164196 269325
rect 163876 262325 163918 262561
rect 164154 262325 164196 262561
rect 163876 255561 164196 262325
rect 163876 255325 163918 255561
rect 164154 255325 164196 255561
rect 163876 248561 164196 255325
rect 163876 248325 163918 248561
rect 164154 248325 164196 248561
rect 163876 241561 164196 248325
rect 163876 241325 163918 241561
rect 164154 241325 164196 241561
rect 163876 234561 164196 241325
rect 163876 234325 163918 234561
rect 164154 234325 164196 234561
rect 163876 227561 164196 234325
rect 163876 227325 163918 227561
rect 164154 227325 164196 227561
rect 163876 220561 164196 227325
rect 163876 220325 163918 220561
rect 164154 220325 164196 220561
rect 163876 213561 164196 220325
rect 163876 213325 163918 213561
rect 164154 213325 164196 213561
rect 163876 206561 164196 213325
rect 163876 206325 163918 206561
rect 164154 206325 164196 206561
rect 163876 199561 164196 206325
rect 163876 199325 163918 199561
rect 164154 199325 164196 199561
rect 163876 192561 164196 199325
rect 163876 192325 163918 192561
rect 164154 192325 164196 192561
rect 163876 185561 164196 192325
rect 163876 185325 163918 185561
rect 164154 185325 164196 185561
rect 163876 178561 164196 185325
rect 163876 178325 163918 178561
rect 164154 178325 164196 178561
rect 163876 171561 164196 178325
rect 163876 171325 163918 171561
rect 164154 171325 164196 171561
rect 163876 164561 164196 171325
rect 163876 164325 163918 164561
rect 164154 164325 164196 164561
rect 163876 157561 164196 164325
rect 163876 157325 163918 157561
rect 164154 157325 164196 157561
rect 163876 150561 164196 157325
rect 163876 150325 163918 150561
rect 164154 150325 164196 150561
rect 163876 143561 164196 150325
rect 163876 143325 163918 143561
rect 164154 143325 164196 143561
rect 163876 136561 164196 143325
rect 163876 136325 163918 136561
rect 164154 136325 164196 136561
rect 163876 129561 164196 136325
rect 163876 129325 163918 129561
rect 164154 129325 164196 129561
rect 163876 122561 164196 129325
rect 163876 122325 163918 122561
rect 164154 122325 164196 122561
rect 163876 115561 164196 122325
rect 163876 115325 163918 115561
rect 164154 115325 164196 115561
rect 163876 108561 164196 115325
rect 163876 108325 163918 108561
rect 164154 108325 164196 108561
rect 163876 101561 164196 108325
rect 163876 101325 163918 101561
rect 164154 101325 164196 101561
rect 163876 94561 164196 101325
rect 163876 94325 163918 94561
rect 164154 94325 164196 94561
rect 163876 87561 164196 94325
rect 163876 87325 163918 87561
rect 164154 87325 164196 87561
rect 163876 80561 164196 87325
rect 163876 80325 163918 80561
rect 164154 80325 164196 80561
rect 163876 73561 164196 80325
rect 163876 73325 163918 73561
rect 164154 73325 164196 73561
rect 163876 66561 164196 73325
rect 163876 66325 163918 66561
rect 164154 66325 164196 66561
rect 163876 59561 164196 66325
rect 163876 59325 163918 59561
rect 164154 59325 164196 59561
rect 163876 52561 164196 59325
rect 163876 52325 163918 52561
rect 164154 52325 164196 52561
rect 163876 45561 164196 52325
rect 163876 45325 163918 45561
rect 164154 45325 164196 45561
rect 163876 38561 164196 45325
rect 163876 38325 163918 38561
rect 164154 38325 164196 38561
rect 163876 31561 164196 38325
rect 163876 31325 163918 31561
rect 164154 31325 164196 31561
rect 163876 24561 164196 31325
rect 163876 24325 163918 24561
rect 164154 24325 164196 24561
rect 163876 17561 164196 24325
rect 163876 17325 163918 17561
rect 164154 17325 164196 17561
rect 163876 10561 164196 17325
rect 163876 10325 163918 10561
rect 164154 10325 164196 10561
rect 163876 3561 164196 10325
rect 163876 3325 163918 3561
rect 164154 3325 164196 3561
rect 163876 -1706 164196 3325
rect 163876 -1942 163918 -1706
rect 164154 -1942 164196 -1706
rect 163876 -2026 164196 -1942
rect 163876 -2262 163918 -2026
rect 164154 -2262 164196 -2026
rect 163876 -2294 164196 -2262
rect 169144 705238 169464 706230
rect 169144 705002 169186 705238
rect 169422 705002 169464 705238
rect 169144 704918 169464 705002
rect 169144 704682 169186 704918
rect 169422 704682 169464 704918
rect 169144 695494 169464 704682
rect 169144 695258 169186 695494
rect 169422 695258 169464 695494
rect 169144 688494 169464 695258
rect 169144 688258 169186 688494
rect 169422 688258 169464 688494
rect 169144 681494 169464 688258
rect 169144 681258 169186 681494
rect 169422 681258 169464 681494
rect 169144 674494 169464 681258
rect 169144 674258 169186 674494
rect 169422 674258 169464 674494
rect 169144 667494 169464 674258
rect 169144 667258 169186 667494
rect 169422 667258 169464 667494
rect 169144 660494 169464 667258
rect 169144 660258 169186 660494
rect 169422 660258 169464 660494
rect 169144 653494 169464 660258
rect 169144 653258 169186 653494
rect 169422 653258 169464 653494
rect 169144 646494 169464 653258
rect 169144 646258 169186 646494
rect 169422 646258 169464 646494
rect 169144 639494 169464 646258
rect 169144 639258 169186 639494
rect 169422 639258 169464 639494
rect 169144 632494 169464 639258
rect 169144 632258 169186 632494
rect 169422 632258 169464 632494
rect 169144 625494 169464 632258
rect 169144 625258 169186 625494
rect 169422 625258 169464 625494
rect 169144 618494 169464 625258
rect 169144 618258 169186 618494
rect 169422 618258 169464 618494
rect 169144 611494 169464 618258
rect 169144 611258 169186 611494
rect 169422 611258 169464 611494
rect 169144 604494 169464 611258
rect 169144 604258 169186 604494
rect 169422 604258 169464 604494
rect 169144 597494 169464 604258
rect 169144 597258 169186 597494
rect 169422 597258 169464 597494
rect 169144 590494 169464 597258
rect 169144 590258 169186 590494
rect 169422 590258 169464 590494
rect 169144 583494 169464 590258
rect 169144 583258 169186 583494
rect 169422 583258 169464 583494
rect 169144 576494 169464 583258
rect 169144 576258 169186 576494
rect 169422 576258 169464 576494
rect 169144 569494 169464 576258
rect 169144 569258 169186 569494
rect 169422 569258 169464 569494
rect 169144 562494 169464 569258
rect 169144 562258 169186 562494
rect 169422 562258 169464 562494
rect 169144 555494 169464 562258
rect 169144 555258 169186 555494
rect 169422 555258 169464 555494
rect 169144 548494 169464 555258
rect 169144 548258 169186 548494
rect 169422 548258 169464 548494
rect 169144 541494 169464 548258
rect 169144 541258 169186 541494
rect 169422 541258 169464 541494
rect 169144 534494 169464 541258
rect 169144 534258 169186 534494
rect 169422 534258 169464 534494
rect 169144 527494 169464 534258
rect 169144 527258 169186 527494
rect 169422 527258 169464 527494
rect 169144 520494 169464 527258
rect 169144 520258 169186 520494
rect 169422 520258 169464 520494
rect 169144 513494 169464 520258
rect 169144 513258 169186 513494
rect 169422 513258 169464 513494
rect 169144 506494 169464 513258
rect 169144 506258 169186 506494
rect 169422 506258 169464 506494
rect 169144 499494 169464 506258
rect 169144 499258 169186 499494
rect 169422 499258 169464 499494
rect 169144 492494 169464 499258
rect 169144 492258 169186 492494
rect 169422 492258 169464 492494
rect 169144 485494 169464 492258
rect 169144 485258 169186 485494
rect 169422 485258 169464 485494
rect 169144 478494 169464 485258
rect 169144 478258 169186 478494
rect 169422 478258 169464 478494
rect 169144 471494 169464 478258
rect 169144 471258 169186 471494
rect 169422 471258 169464 471494
rect 169144 464494 169464 471258
rect 169144 464258 169186 464494
rect 169422 464258 169464 464494
rect 169144 457494 169464 464258
rect 169144 457258 169186 457494
rect 169422 457258 169464 457494
rect 169144 450494 169464 457258
rect 169144 450258 169186 450494
rect 169422 450258 169464 450494
rect 169144 443494 169464 450258
rect 169144 443258 169186 443494
rect 169422 443258 169464 443494
rect 169144 436494 169464 443258
rect 169144 436258 169186 436494
rect 169422 436258 169464 436494
rect 169144 429494 169464 436258
rect 169144 429258 169186 429494
rect 169422 429258 169464 429494
rect 169144 422494 169464 429258
rect 169144 422258 169186 422494
rect 169422 422258 169464 422494
rect 169144 415494 169464 422258
rect 169144 415258 169186 415494
rect 169422 415258 169464 415494
rect 169144 408494 169464 415258
rect 169144 408258 169186 408494
rect 169422 408258 169464 408494
rect 169144 401494 169464 408258
rect 169144 401258 169186 401494
rect 169422 401258 169464 401494
rect 169144 394494 169464 401258
rect 169144 394258 169186 394494
rect 169422 394258 169464 394494
rect 169144 387494 169464 394258
rect 169144 387258 169186 387494
rect 169422 387258 169464 387494
rect 169144 380494 169464 387258
rect 169144 380258 169186 380494
rect 169422 380258 169464 380494
rect 169144 373494 169464 380258
rect 169144 373258 169186 373494
rect 169422 373258 169464 373494
rect 169144 366494 169464 373258
rect 169144 366258 169186 366494
rect 169422 366258 169464 366494
rect 169144 359494 169464 366258
rect 169144 359258 169186 359494
rect 169422 359258 169464 359494
rect 169144 352494 169464 359258
rect 169144 352258 169186 352494
rect 169422 352258 169464 352494
rect 169144 345494 169464 352258
rect 169144 345258 169186 345494
rect 169422 345258 169464 345494
rect 169144 338494 169464 345258
rect 169144 338258 169186 338494
rect 169422 338258 169464 338494
rect 169144 331494 169464 338258
rect 169144 331258 169186 331494
rect 169422 331258 169464 331494
rect 169144 324494 169464 331258
rect 169144 324258 169186 324494
rect 169422 324258 169464 324494
rect 169144 317494 169464 324258
rect 169144 317258 169186 317494
rect 169422 317258 169464 317494
rect 169144 310494 169464 317258
rect 169144 310258 169186 310494
rect 169422 310258 169464 310494
rect 169144 303494 169464 310258
rect 169144 303258 169186 303494
rect 169422 303258 169464 303494
rect 169144 296494 169464 303258
rect 169144 296258 169186 296494
rect 169422 296258 169464 296494
rect 169144 289494 169464 296258
rect 169144 289258 169186 289494
rect 169422 289258 169464 289494
rect 169144 282494 169464 289258
rect 169144 282258 169186 282494
rect 169422 282258 169464 282494
rect 169144 275494 169464 282258
rect 169144 275258 169186 275494
rect 169422 275258 169464 275494
rect 169144 268494 169464 275258
rect 169144 268258 169186 268494
rect 169422 268258 169464 268494
rect 169144 261494 169464 268258
rect 169144 261258 169186 261494
rect 169422 261258 169464 261494
rect 169144 254494 169464 261258
rect 169144 254258 169186 254494
rect 169422 254258 169464 254494
rect 169144 247494 169464 254258
rect 169144 247258 169186 247494
rect 169422 247258 169464 247494
rect 169144 240494 169464 247258
rect 169144 240258 169186 240494
rect 169422 240258 169464 240494
rect 169144 233494 169464 240258
rect 169144 233258 169186 233494
rect 169422 233258 169464 233494
rect 169144 226494 169464 233258
rect 169144 226258 169186 226494
rect 169422 226258 169464 226494
rect 169144 219494 169464 226258
rect 169144 219258 169186 219494
rect 169422 219258 169464 219494
rect 169144 212494 169464 219258
rect 169144 212258 169186 212494
rect 169422 212258 169464 212494
rect 169144 205494 169464 212258
rect 169144 205258 169186 205494
rect 169422 205258 169464 205494
rect 169144 198494 169464 205258
rect 169144 198258 169186 198494
rect 169422 198258 169464 198494
rect 169144 191494 169464 198258
rect 169144 191258 169186 191494
rect 169422 191258 169464 191494
rect 169144 184494 169464 191258
rect 169144 184258 169186 184494
rect 169422 184258 169464 184494
rect 169144 177494 169464 184258
rect 169144 177258 169186 177494
rect 169422 177258 169464 177494
rect 169144 170494 169464 177258
rect 169144 170258 169186 170494
rect 169422 170258 169464 170494
rect 169144 163494 169464 170258
rect 169144 163258 169186 163494
rect 169422 163258 169464 163494
rect 169144 156494 169464 163258
rect 169144 156258 169186 156494
rect 169422 156258 169464 156494
rect 169144 149494 169464 156258
rect 169144 149258 169186 149494
rect 169422 149258 169464 149494
rect 169144 142494 169464 149258
rect 169144 142258 169186 142494
rect 169422 142258 169464 142494
rect 169144 135494 169464 142258
rect 169144 135258 169186 135494
rect 169422 135258 169464 135494
rect 169144 128494 169464 135258
rect 169144 128258 169186 128494
rect 169422 128258 169464 128494
rect 169144 121494 169464 128258
rect 169144 121258 169186 121494
rect 169422 121258 169464 121494
rect 169144 114494 169464 121258
rect 169144 114258 169186 114494
rect 169422 114258 169464 114494
rect 169144 107494 169464 114258
rect 169144 107258 169186 107494
rect 169422 107258 169464 107494
rect 169144 100494 169464 107258
rect 169144 100258 169186 100494
rect 169422 100258 169464 100494
rect 169144 93494 169464 100258
rect 169144 93258 169186 93494
rect 169422 93258 169464 93494
rect 169144 86494 169464 93258
rect 169144 86258 169186 86494
rect 169422 86258 169464 86494
rect 169144 79494 169464 86258
rect 169144 79258 169186 79494
rect 169422 79258 169464 79494
rect 169144 72494 169464 79258
rect 169144 72258 169186 72494
rect 169422 72258 169464 72494
rect 169144 65494 169464 72258
rect 169144 65258 169186 65494
rect 169422 65258 169464 65494
rect 169144 58494 169464 65258
rect 169144 58258 169186 58494
rect 169422 58258 169464 58494
rect 169144 51494 169464 58258
rect 169144 51258 169186 51494
rect 169422 51258 169464 51494
rect 169144 44494 169464 51258
rect 169144 44258 169186 44494
rect 169422 44258 169464 44494
rect 169144 37494 169464 44258
rect 169144 37258 169186 37494
rect 169422 37258 169464 37494
rect 169144 30494 169464 37258
rect 169144 30258 169186 30494
rect 169422 30258 169464 30494
rect 169144 23494 169464 30258
rect 169144 23258 169186 23494
rect 169422 23258 169464 23494
rect 169144 16494 169464 23258
rect 169144 16258 169186 16494
rect 169422 16258 169464 16494
rect 169144 9494 169464 16258
rect 169144 9258 169186 9494
rect 169422 9258 169464 9494
rect 169144 2494 169464 9258
rect 169144 2258 169186 2494
rect 169422 2258 169464 2494
rect 169144 -746 169464 2258
rect 169144 -982 169186 -746
rect 169422 -982 169464 -746
rect 169144 -1066 169464 -982
rect 169144 -1302 169186 -1066
rect 169422 -1302 169464 -1066
rect 169144 -2294 169464 -1302
rect 170876 706198 171196 706230
rect 170876 705962 170918 706198
rect 171154 705962 171196 706198
rect 170876 705878 171196 705962
rect 170876 705642 170918 705878
rect 171154 705642 171196 705878
rect 170876 696561 171196 705642
rect 170876 696325 170918 696561
rect 171154 696325 171196 696561
rect 170876 689561 171196 696325
rect 170876 689325 170918 689561
rect 171154 689325 171196 689561
rect 170876 682561 171196 689325
rect 170876 682325 170918 682561
rect 171154 682325 171196 682561
rect 170876 675561 171196 682325
rect 170876 675325 170918 675561
rect 171154 675325 171196 675561
rect 170876 668561 171196 675325
rect 170876 668325 170918 668561
rect 171154 668325 171196 668561
rect 170876 661561 171196 668325
rect 170876 661325 170918 661561
rect 171154 661325 171196 661561
rect 170876 654561 171196 661325
rect 170876 654325 170918 654561
rect 171154 654325 171196 654561
rect 170876 647561 171196 654325
rect 170876 647325 170918 647561
rect 171154 647325 171196 647561
rect 170876 640561 171196 647325
rect 170876 640325 170918 640561
rect 171154 640325 171196 640561
rect 170876 633561 171196 640325
rect 170876 633325 170918 633561
rect 171154 633325 171196 633561
rect 170876 626561 171196 633325
rect 170876 626325 170918 626561
rect 171154 626325 171196 626561
rect 170876 619561 171196 626325
rect 170876 619325 170918 619561
rect 171154 619325 171196 619561
rect 170876 612561 171196 619325
rect 170876 612325 170918 612561
rect 171154 612325 171196 612561
rect 170876 605561 171196 612325
rect 170876 605325 170918 605561
rect 171154 605325 171196 605561
rect 170876 598561 171196 605325
rect 170876 598325 170918 598561
rect 171154 598325 171196 598561
rect 170876 591561 171196 598325
rect 170876 591325 170918 591561
rect 171154 591325 171196 591561
rect 170876 584561 171196 591325
rect 170876 584325 170918 584561
rect 171154 584325 171196 584561
rect 170876 577561 171196 584325
rect 170876 577325 170918 577561
rect 171154 577325 171196 577561
rect 170876 570561 171196 577325
rect 170876 570325 170918 570561
rect 171154 570325 171196 570561
rect 170876 563561 171196 570325
rect 170876 563325 170918 563561
rect 171154 563325 171196 563561
rect 170876 556561 171196 563325
rect 170876 556325 170918 556561
rect 171154 556325 171196 556561
rect 170876 549561 171196 556325
rect 170876 549325 170918 549561
rect 171154 549325 171196 549561
rect 170876 542561 171196 549325
rect 170876 542325 170918 542561
rect 171154 542325 171196 542561
rect 170876 535561 171196 542325
rect 170876 535325 170918 535561
rect 171154 535325 171196 535561
rect 170876 528561 171196 535325
rect 170876 528325 170918 528561
rect 171154 528325 171196 528561
rect 170876 521561 171196 528325
rect 170876 521325 170918 521561
rect 171154 521325 171196 521561
rect 170876 514561 171196 521325
rect 170876 514325 170918 514561
rect 171154 514325 171196 514561
rect 170876 507561 171196 514325
rect 170876 507325 170918 507561
rect 171154 507325 171196 507561
rect 170876 500561 171196 507325
rect 170876 500325 170918 500561
rect 171154 500325 171196 500561
rect 170876 493561 171196 500325
rect 170876 493325 170918 493561
rect 171154 493325 171196 493561
rect 170876 486561 171196 493325
rect 170876 486325 170918 486561
rect 171154 486325 171196 486561
rect 170876 479561 171196 486325
rect 170876 479325 170918 479561
rect 171154 479325 171196 479561
rect 170876 472561 171196 479325
rect 170876 472325 170918 472561
rect 171154 472325 171196 472561
rect 170876 465561 171196 472325
rect 170876 465325 170918 465561
rect 171154 465325 171196 465561
rect 170876 458561 171196 465325
rect 170876 458325 170918 458561
rect 171154 458325 171196 458561
rect 170876 451561 171196 458325
rect 170876 451325 170918 451561
rect 171154 451325 171196 451561
rect 170876 444561 171196 451325
rect 170876 444325 170918 444561
rect 171154 444325 171196 444561
rect 170876 437561 171196 444325
rect 170876 437325 170918 437561
rect 171154 437325 171196 437561
rect 170876 430561 171196 437325
rect 170876 430325 170918 430561
rect 171154 430325 171196 430561
rect 170876 423561 171196 430325
rect 170876 423325 170918 423561
rect 171154 423325 171196 423561
rect 170876 416561 171196 423325
rect 170876 416325 170918 416561
rect 171154 416325 171196 416561
rect 170876 409561 171196 416325
rect 170876 409325 170918 409561
rect 171154 409325 171196 409561
rect 170876 402561 171196 409325
rect 170876 402325 170918 402561
rect 171154 402325 171196 402561
rect 170876 395561 171196 402325
rect 170876 395325 170918 395561
rect 171154 395325 171196 395561
rect 170876 388561 171196 395325
rect 170876 388325 170918 388561
rect 171154 388325 171196 388561
rect 170876 381561 171196 388325
rect 170876 381325 170918 381561
rect 171154 381325 171196 381561
rect 170876 374561 171196 381325
rect 170876 374325 170918 374561
rect 171154 374325 171196 374561
rect 170876 367561 171196 374325
rect 170876 367325 170918 367561
rect 171154 367325 171196 367561
rect 170876 360561 171196 367325
rect 170876 360325 170918 360561
rect 171154 360325 171196 360561
rect 170876 353561 171196 360325
rect 170876 353325 170918 353561
rect 171154 353325 171196 353561
rect 170876 346561 171196 353325
rect 170876 346325 170918 346561
rect 171154 346325 171196 346561
rect 170876 339561 171196 346325
rect 170876 339325 170918 339561
rect 171154 339325 171196 339561
rect 170876 332561 171196 339325
rect 170876 332325 170918 332561
rect 171154 332325 171196 332561
rect 170876 325561 171196 332325
rect 170876 325325 170918 325561
rect 171154 325325 171196 325561
rect 170876 318561 171196 325325
rect 170876 318325 170918 318561
rect 171154 318325 171196 318561
rect 170876 311561 171196 318325
rect 170876 311325 170918 311561
rect 171154 311325 171196 311561
rect 170876 304561 171196 311325
rect 170876 304325 170918 304561
rect 171154 304325 171196 304561
rect 170876 297561 171196 304325
rect 170876 297325 170918 297561
rect 171154 297325 171196 297561
rect 170876 290561 171196 297325
rect 170876 290325 170918 290561
rect 171154 290325 171196 290561
rect 170876 283561 171196 290325
rect 170876 283325 170918 283561
rect 171154 283325 171196 283561
rect 170876 276561 171196 283325
rect 170876 276325 170918 276561
rect 171154 276325 171196 276561
rect 170876 269561 171196 276325
rect 170876 269325 170918 269561
rect 171154 269325 171196 269561
rect 170876 262561 171196 269325
rect 170876 262325 170918 262561
rect 171154 262325 171196 262561
rect 170876 255561 171196 262325
rect 170876 255325 170918 255561
rect 171154 255325 171196 255561
rect 170876 248561 171196 255325
rect 170876 248325 170918 248561
rect 171154 248325 171196 248561
rect 170876 241561 171196 248325
rect 170876 241325 170918 241561
rect 171154 241325 171196 241561
rect 170876 234561 171196 241325
rect 170876 234325 170918 234561
rect 171154 234325 171196 234561
rect 170876 227561 171196 234325
rect 170876 227325 170918 227561
rect 171154 227325 171196 227561
rect 170876 220561 171196 227325
rect 170876 220325 170918 220561
rect 171154 220325 171196 220561
rect 170876 213561 171196 220325
rect 170876 213325 170918 213561
rect 171154 213325 171196 213561
rect 170876 206561 171196 213325
rect 170876 206325 170918 206561
rect 171154 206325 171196 206561
rect 170876 199561 171196 206325
rect 170876 199325 170918 199561
rect 171154 199325 171196 199561
rect 170876 192561 171196 199325
rect 170876 192325 170918 192561
rect 171154 192325 171196 192561
rect 170876 185561 171196 192325
rect 170876 185325 170918 185561
rect 171154 185325 171196 185561
rect 170876 178561 171196 185325
rect 170876 178325 170918 178561
rect 171154 178325 171196 178561
rect 170876 171561 171196 178325
rect 170876 171325 170918 171561
rect 171154 171325 171196 171561
rect 170876 164561 171196 171325
rect 170876 164325 170918 164561
rect 171154 164325 171196 164561
rect 170876 157561 171196 164325
rect 170876 157325 170918 157561
rect 171154 157325 171196 157561
rect 170876 150561 171196 157325
rect 170876 150325 170918 150561
rect 171154 150325 171196 150561
rect 170876 143561 171196 150325
rect 170876 143325 170918 143561
rect 171154 143325 171196 143561
rect 170876 136561 171196 143325
rect 170876 136325 170918 136561
rect 171154 136325 171196 136561
rect 170876 129561 171196 136325
rect 170876 129325 170918 129561
rect 171154 129325 171196 129561
rect 170876 122561 171196 129325
rect 170876 122325 170918 122561
rect 171154 122325 171196 122561
rect 170876 115561 171196 122325
rect 170876 115325 170918 115561
rect 171154 115325 171196 115561
rect 170876 108561 171196 115325
rect 170876 108325 170918 108561
rect 171154 108325 171196 108561
rect 170876 101561 171196 108325
rect 170876 101325 170918 101561
rect 171154 101325 171196 101561
rect 170876 94561 171196 101325
rect 170876 94325 170918 94561
rect 171154 94325 171196 94561
rect 170876 87561 171196 94325
rect 170876 87325 170918 87561
rect 171154 87325 171196 87561
rect 170876 80561 171196 87325
rect 170876 80325 170918 80561
rect 171154 80325 171196 80561
rect 170876 73561 171196 80325
rect 170876 73325 170918 73561
rect 171154 73325 171196 73561
rect 170876 66561 171196 73325
rect 170876 66325 170918 66561
rect 171154 66325 171196 66561
rect 170876 59561 171196 66325
rect 170876 59325 170918 59561
rect 171154 59325 171196 59561
rect 170876 52561 171196 59325
rect 170876 52325 170918 52561
rect 171154 52325 171196 52561
rect 170876 45561 171196 52325
rect 170876 45325 170918 45561
rect 171154 45325 171196 45561
rect 170876 38561 171196 45325
rect 170876 38325 170918 38561
rect 171154 38325 171196 38561
rect 170876 31561 171196 38325
rect 170876 31325 170918 31561
rect 171154 31325 171196 31561
rect 170876 24561 171196 31325
rect 170876 24325 170918 24561
rect 171154 24325 171196 24561
rect 170876 17561 171196 24325
rect 170876 17325 170918 17561
rect 171154 17325 171196 17561
rect 170876 10561 171196 17325
rect 170876 10325 170918 10561
rect 171154 10325 171196 10561
rect 170876 3561 171196 10325
rect 170876 3325 170918 3561
rect 171154 3325 171196 3561
rect 170876 -1706 171196 3325
rect 170876 -1942 170918 -1706
rect 171154 -1942 171196 -1706
rect 170876 -2026 171196 -1942
rect 170876 -2262 170918 -2026
rect 171154 -2262 171196 -2026
rect 170876 -2294 171196 -2262
rect 176144 705238 176464 706230
rect 176144 705002 176186 705238
rect 176422 705002 176464 705238
rect 176144 704918 176464 705002
rect 176144 704682 176186 704918
rect 176422 704682 176464 704918
rect 176144 695494 176464 704682
rect 176144 695258 176186 695494
rect 176422 695258 176464 695494
rect 176144 688494 176464 695258
rect 176144 688258 176186 688494
rect 176422 688258 176464 688494
rect 176144 681494 176464 688258
rect 176144 681258 176186 681494
rect 176422 681258 176464 681494
rect 176144 674494 176464 681258
rect 176144 674258 176186 674494
rect 176422 674258 176464 674494
rect 176144 667494 176464 674258
rect 176144 667258 176186 667494
rect 176422 667258 176464 667494
rect 176144 660494 176464 667258
rect 176144 660258 176186 660494
rect 176422 660258 176464 660494
rect 176144 653494 176464 660258
rect 176144 653258 176186 653494
rect 176422 653258 176464 653494
rect 176144 646494 176464 653258
rect 176144 646258 176186 646494
rect 176422 646258 176464 646494
rect 176144 639494 176464 646258
rect 176144 639258 176186 639494
rect 176422 639258 176464 639494
rect 176144 632494 176464 639258
rect 176144 632258 176186 632494
rect 176422 632258 176464 632494
rect 176144 625494 176464 632258
rect 176144 625258 176186 625494
rect 176422 625258 176464 625494
rect 176144 618494 176464 625258
rect 176144 618258 176186 618494
rect 176422 618258 176464 618494
rect 176144 611494 176464 618258
rect 176144 611258 176186 611494
rect 176422 611258 176464 611494
rect 176144 604494 176464 611258
rect 176144 604258 176186 604494
rect 176422 604258 176464 604494
rect 176144 597494 176464 604258
rect 176144 597258 176186 597494
rect 176422 597258 176464 597494
rect 176144 590494 176464 597258
rect 176144 590258 176186 590494
rect 176422 590258 176464 590494
rect 176144 583494 176464 590258
rect 176144 583258 176186 583494
rect 176422 583258 176464 583494
rect 176144 576494 176464 583258
rect 176144 576258 176186 576494
rect 176422 576258 176464 576494
rect 176144 569494 176464 576258
rect 176144 569258 176186 569494
rect 176422 569258 176464 569494
rect 176144 562494 176464 569258
rect 176144 562258 176186 562494
rect 176422 562258 176464 562494
rect 176144 555494 176464 562258
rect 176144 555258 176186 555494
rect 176422 555258 176464 555494
rect 176144 548494 176464 555258
rect 176144 548258 176186 548494
rect 176422 548258 176464 548494
rect 176144 541494 176464 548258
rect 176144 541258 176186 541494
rect 176422 541258 176464 541494
rect 176144 534494 176464 541258
rect 176144 534258 176186 534494
rect 176422 534258 176464 534494
rect 176144 527494 176464 534258
rect 176144 527258 176186 527494
rect 176422 527258 176464 527494
rect 176144 520494 176464 527258
rect 176144 520258 176186 520494
rect 176422 520258 176464 520494
rect 176144 513494 176464 520258
rect 176144 513258 176186 513494
rect 176422 513258 176464 513494
rect 176144 506494 176464 513258
rect 176144 506258 176186 506494
rect 176422 506258 176464 506494
rect 176144 499494 176464 506258
rect 176144 499258 176186 499494
rect 176422 499258 176464 499494
rect 176144 492494 176464 499258
rect 176144 492258 176186 492494
rect 176422 492258 176464 492494
rect 176144 485494 176464 492258
rect 176144 485258 176186 485494
rect 176422 485258 176464 485494
rect 176144 478494 176464 485258
rect 176144 478258 176186 478494
rect 176422 478258 176464 478494
rect 176144 471494 176464 478258
rect 176144 471258 176186 471494
rect 176422 471258 176464 471494
rect 176144 464494 176464 471258
rect 176144 464258 176186 464494
rect 176422 464258 176464 464494
rect 176144 457494 176464 464258
rect 176144 457258 176186 457494
rect 176422 457258 176464 457494
rect 176144 450494 176464 457258
rect 176144 450258 176186 450494
rect 176422 450258 176464 450494
rect 176144 443494 176464 450258
rect 176144 443258 176186 443494
rect 176422 443258 176464 443494
rect 176144 436494 176464 443258
rect 176144 436258 176186 436494
rect 176422 436258 176464 436494
rect 176144 429494 176464 436258
rect 176144 429258 176186 429494
rect 176422 429258 176464 429494
rect 176144 422494 176464 429258
rect 176144 422258 176186 422494
rect 176422 422258 176464 422494
rect 176144 415494 176464 422258
rect 176144 415258 176186 415494
rect 176422 415258 176464 415494
rect 176144 408494 176464 415258
rect 176144 408258 176186 408494
rect 176422 408258 176464 408494
rect 176144 401494 176464 408258
rect 176144 401258 176186 401494
rect 176422 401258 176464 401494
rect 176144 394494 176464 401258
rect 176144 394258 176186 394494
rect 176422 394258 176464 394494
rect 176144 387494 176464 394258
rect 176144 387258 176186 387494
rect 176422 387258 176464 387494
rect 176144 380494 176464 387258
rect 176144 380258 176186 380494
rect 176422 380258 176464 380494
rect 176144 373494 176464 380258
rect 176144 373258 176186 373494
rect 176422 373258 176464 373494
rect 176144 366494 176464 373258
rect 176144 366258 176186 366494
rect 176422 366258 176464 366494
rect 176144 359494 176464 366258
rect 176144 359258 176186 359494
rect 176422 359258 176464 359494
rect 176144 352494 176464 359258
rect 176144 352258 176186 352494
rect 176422 352258 176464 352494
rect 176144 345494 176464 352258
rect 176144 345258 176186 345494
rect 176422 345258 176464 345494
rect 176144 338494 176464 345258
rect 176144 338258 176186 338494
rect 176422 338258 176464 338494
rect 176144 331494 176464 338258
rect 176144 331258 176186 331494
rect 176422 331258 176464 331494
rect 176144 324494 176464 331258
rect 176144 324258 176186 324494
rect 176422 324258 176464 324494
rect 176144 317494 176464 324258
rect 176144 317258 176186 317494
rect 176422 317258 176464 317494
rect 176144 310494 176464 317258
rect 176144 310258 176186 310494
rect 176422 310258 176464 310494
rect 176144 303494 176464 310258
rect 176144 303258 176186 303494
rect 176422 303258 176464 303494
rect 176144 296494 176464 303258
rect 176144 296258 176186 296494
rect 176422 296258 176464 296494
rect 176144 289494 176464 296258
rect 176144 289258 176186 289494
rect 176422 289258 176464 289494
rect 176144 282494 176464 289258
rect 176144 282258 176186 282494
rect 176422 282258 176464 282494
rect 176144 275494 176464 282258
rect 176144 275258 176186 275494
rect 176422 275258 176464 275494
rect 176144 268494 176464 275258
rect 176144 268258 176186 268494
rect 176422 268258 176464 268494
rect 176144 261494 176464 268258
rect 176144 261258 176186 261494
rect 176422 261258 176464 261494
rect 176144 254494 176464 261258
rect 176144 254258 176186 254494
rect 176422 254258 176464 254494
rect 176144 247494 176464 254258
rect 176144 247258 176186 247494
rect 176422 247258 176464 247494
rect 176144 240494 176464 247258
rect 176144 240258 176186 240494
rect 176422 240258 176464 240494
rect 176144 233494 176464 240258
rect 176144 233258 176186 233494
rect 176422 233258 176464 233494
rect 176144 226494 176464 233258
rect 176144 226258 176186 226494
rect 176422 226258 176464 226494
rect 176144 219494 176464 226258
rect 176144 219258 176186 219494
rect 176422 219258 176464 219494
rect 176144 212494 176464 219258
rect 176144 212258 176186 212494
rect 176422 212258 176464 212494
rect 176144 205494 176464 212258
rect 176144 205258 176186 205494
rect 176422 205258 176464 205494
rect 176144 198494 176464 205258
rect 176144 198258 176186 198494
rect 176422 198258 176464 198494
rect 176144 191494 176464 198258
rect 176144 191258 176186 191494
rect 176422 191258 176464 191494
rect 176144 184494 176464 191258
rect 176144 184258 176186 184494
rect 176422 184258 176464 184494
rect 176144 177494 176464 184258
rect 176144 177258 176186 177494
rect 176422 177258 176464 177494
rect 176144 170494 176464 177258
rect 176144 170258 176186 170494
rect 176422 170258 176464 170494
rect 176144 163494 176464 170258
rect 176144 163258 176186 163494
rect 176422 163258 176464 163494
rect 176144 156494 176464 163258
rect 176144 156258 176186 156494
rect 176422 156258 176464 156494
rect 176144 149494 176464 156258
rect 176144 149258 176186 149494
rect 176422 149258 176464 149494
rect 176144 142494 176464 149258
rect 176144 142258 176186 142494
rect 176422 142258 176464 142494
rect 176144 135494 176464 142258
rect 176144 135258 176186 135494
rect 176422 135258 176464 135494
rect 176144 128494 176464 135258
rect 176144 128258 176186 128494
rect 176422 128258 176464 128494
rect 176144 121494 176464 128258
rect 176144 121258 176186 121494
rect 176422 121258 176464 121494
rect 176144 114494 176464 121258
rect 176144 114258 176186 114494
rect 176422 114258 176464 114494
rect 176144 107494 176464 114258
rect 176144 107258 176186 107494
rect 176422 107258 176464 107494
rect 176144 100494 176464 107258
rect 176144 100258 176186 100494
rect 176422 100258 176464 100494
rect 176144 93494 176464 100258
rect 176144 93258 176186 93494
rect 176422 93258 176464 93494
rect 176144 86494 176464 93258
rect 176144 86258 176186 86494
rect 176422 86258 176464 86494
rect 176144 79494 176464 86258
rect 176144 79258 176186 79494
rect 176422 79258 176464 79494
rect 176144 72494 176464 79258
rect 176144 72258 176186 72494
rect 176422 72258 176464 72494
rect 176144 65494 176464 72258
rect 176144 65258 176186 65494
rect 176422 65258 176464 65494
rect 176144 58494 176464 65258
rect 176144 58258 176186 58494
rect 176422 58258 176464 58494
rect 176144 51494 176464 58258
rect 176144 51258 176186 51494
rect 176422 51258 176464 51494
rect 176144 44494 176464 51258
rect 176144 44258 176186 44494
rect 176422 44258 176464 44494
rect 176144 37494 176464 44258
rect 176144 37258 176186 37494
rect 176422 37258 176464 37494
rect 176144 30494 176464 37258
rect 176144 30258 176186 30494
rect 176422 30258 176464 30494
rect 176144 23494 176464 30258
rect 176144 23258 176186 23494
rect 176422 23258 176464 23494
rect 176144 16494 176464 23258
rect 176144 16258 176186 16494
rect 176422 16258 176464 16494
rect 176144 9494 176464 16258
rect 176144 9258 176186 9494
rect 176422 9258 176464 9494
rect 176144 2494 176464 9258
rect 176144 2258 176186 2494
rect 176422 2258 176464 2494
rect 176144 -746 176464 2258
rect 176144 -982 176186 -746
rect 176422 -982 176464 -746
rect 176144 -1066 176464 -982
rect 176144 -1302 176186 -1066
rect 176422 -1302 176464 -1066
rect 176144 -2294 176464 -1302
rect 177876 706198 178196 706230
rect 177876 705962 177918 706198
rect 178154 705962 178196 706198
rect 177876 705878 178196 705962
rect 177876 705642 177918 705878
rect 178154 705642 178196 705878
rect 177876 696561 178196 705642
rect 177876 696325 177918 696561
rect 178154 696325 178196 696561
rect 177876 689561 178196 696325
rect 177876 689325 177918 689561
rect 178154 689325 178196 689561
rect 177876 682561 178196 689325
rect 177876 682325 177918 682561
rect 178154 682325 178196 682561
rect 177876 675561 178196 682325
rect 177876 675325 177918 675561
rect 178154 675325 178196 675561
rect 177876 668561 178196 675325
rect 177876 668325 177918 668561
rect 178154 668325 178196 668561
rect 177876 661561 178196 668325
rect 177876 661325 177918 661561
rect 178154 661325 178196 661561
rect 177876 654561 178196 661325
rect 177876 654325 177918 654561
rect 178154 654325 178196 654561
rect 177876 647561 178196 654325
rect 177876 647325 177918 647561
rect 178154 647325 178196 647561
rect 177876 640561 178196 647325
rect 177876 640325 177918 640561
rect 178154 640325 178196 640561
rect 177876 633561 178196 640325
rect 177876 633325 177918 633561
rect 178154 633325 178196 633561
rect 177876 626561 178196 633325
rect 177876 626325 177918 626561
rect 178154 626325 178196 626561
rect 177876 619561 178196 626325
rect 177876 619325 177918 619561
rect 178154 619325 178196 619561
rect 177876 612561 178196 619325
rect 177876 612325 177918 612561
rect 178154 612325 178196 612561
rect 177876 605561 178196 612325
rect 177876 605325 177918 605561
rect 178154 605325 178196 605561
rect 177876 598561 178196 605325
rect 177876 598325 177918 598561
rect 178154 598325 178196 598561
rect 177876 591561 178196 598325
rect 177876 591325 177918 591561
rect 178154 591325 178196 591561
rect 177876 584561 178196 591325
rect 177876 584325 177918 584561
rect 178154 584325 178196 584561
rect 177876 577561 178196 584325
rect 177876 577325 177918 577561
rect 178154 577325 178196 577561
rect 177876 570561 178196 577325
rect 177876 570325 177918 570561
rect 178154 570325 178196 570561
rect 177876 563561 178196 570325
rect 177876 563325 177918 563561
rect 178154 563325 178196 563561
rect 177876 556561 178196 563325
rect 177876 556325 177918 556561
rect 178154 556325 178196 556561
rect 177876 549561 178196 556325
rect 177876 549325 177918 549561
rect 178154 549325 178196 549561
rect 177876 542561 178196 549325
rect 177876 542325 177918 542561
rect 178154 542325 178196 542561
rect 177876 535561 178196 542325
rect 177876 535325 177918 535561
rect 178154 535325 178196 535561
rect 177876 528561 178196 535325
rect 177876 528325 177918 528561
rect 178154 528325 178196 528561
rect 177876 521561 178196 528325
rect 177876 521325 177918 521561
rect 178154 521325 178196 521561
rect 177876 514561 178196 521325
rect 177876 514325 177918 514561
rect 178154 514325 178196 514561
rect 177876 507561 178196 514325
rect 177876 507325 177918 507561
rect 178154 507325 178196 507561
rect 177876 500561 178196 507325
rect 177876 500325 177918 500561
rect 178154 500325 178196 500561
rect 177876 493561 178196 500325
rect 177876 493325 177918 493561
rect 178154 493325 178196 493561
rect 177876 486561 178196 493325
rect 177876 486325 177918 486561
rect 178154 486325 178196 486561
rect 177876 479561 178196 486325
rect 177876 479325 177918 479561
rect 178154 479325 178196 479561
rect 177876 472561 178196 479325
rect 177876 472325 177918 472561
rect 178154 472325 178196 472561
rect 177876 465561 178196 472325
rect 177876 465325 177918 465561
rect 178154 465325 178196 465561
rect 177876 458561 178196 465325
rect 177876 458325 177918 458561
rect 178154 458325 178196 458561
rect 177876 451561 178196 458325
rect 177876 451325 177918 451561
rect 178154 451325 178196 451561
rect 177876 444561 178196 451325
rect 177876 444325 177918 444561
rect 178154 444325 178196 444561
rect 177876 437561 178196 444325
rect 177876 437325 177918 437561
rect 178154 437325 178196 437561
rect 177876 430561 178196 437325
rect 177876 430325 177918 430561
rect 178154 430325 178196 430561
rect 177876 423561 178196 430325
rect 177876 423325 177918 423561
rect 178154 423325 178196 423561
rect 177876 416561 178196 423325
rect 177876 416325 177918 416561
rect 178154 416325 178196 416561
rect 177876 409561 178196 416325
rect 177876 409325 177918 409561
rect 178154 409325 178196 409561
rect 177876 402561 178196 409325
rect 177876 402325 177918 402561
rect 178154 402325 178196 402561
rect 177876 395561 178196 402325
rect 177876 395325 177918 395561
rect 178154 395325 178196 395561
rect 177876 388561 178196 395325
rect 177876 388325 177918 388561
rect 178154 388325 178196 388561
rect 177876 381561 178196 388325
rect 177876 381325 177918 381561
rect 178154 381325 178196 381561
rect 177876 374561 178196 381325
rect 177876 374325 177918 374561
rect 178154 374325 178196 374561
rect 177876 367561 178196 374325
rect 177876 367325 177918 367561
rect 178154 367325 178196 367561
rect 177876 360561 178196 367325
rect 177876 360325 177918 360561
rect 178154 360325 178196 360561
rect 177876 353561 178196 360325
rect 177876 353325 177918 353561
rect 178154 353325 178196 353561
rect 177876 346561 178196 353325
rect 177876 346325 177918 346561
rect 178154 346325 178196 346561
rect 177876 339561 178196 346325
rect 177876 339325 177918 339561
rect 178154 339325 178196 339561
rect 177876 332561 178196 339325
rect 177876 332325 177918 332561
rect 178154 332325 178196 332561
rect 177876 325561 178196 332325
rect 177876 325325 177918 325561
rect 178154 325325 178196 325561
rect 177876 318561 178196 325325
rect 177876 318325 177918 318561
rect 178154 318325 178196 318561
rect 177876 311561 178196 318325
rect 177876 311325 177918 311561
rect 178154 311325 178196 311561
rect 177876 304561 178196 311325
rect 177876 304325 177918 304561
rect 178154 304325 178196 304561
rect 177876 297561 178196 304325
rect 177876 297325 177918 297561
rect 178154 297325 178196 297561
rect 177876 290561 178196 297325
rect 177876 290325 177918 290561
rect 178154 290325 178196 290561
rect 177876 283561 178196 290325
rect 177876 283325 177918 283561
rect 178154 283325 178196 283561
rect 177876 276561 178196 283325
rect 177876 276325 177918 276561
rect 178154 276325 178196 276561
rect 177876 269561 178196 276325
rect 177876 269325 177918 269561
rect 178154 269325 178196 269561
rect 177876 262561 178196 269325
rect 177876 262325 177918 262561
rect 178154 262325 178196 262561
rect 177876 255561 178196 262325
rect 177876 255325 177918 255561
rect 178154 255325 178196 255561
rect 177876 248561 178196 255325
rect 177876 248325 177918 248561
rect 178154 248325 178196 248561
rect 177876 241561 178196 248325
rect 177876 241325 177918 241561
rect 178154 241325 178196 241561
rect 177876 234561 178196 241325
rect 177876 234325 177918 234561
rect 178154 234325 178196 234561
rect 177876 227561 178196 234325
rect 177876 227325 177918 227561
rect 178154 227325 178196 227561
rect 177876 220561 178196 227325
rect 177876 220325 177918 220561
rect 178154 220325 178196 220561
rect 177876 213561 178196 220325
rect 177876 213325 177918 213561
rect 178154 213325 178196 213561
rect 177876 206561 178196 213325
rect 177876 206325 177918 206561
rect 178154 206325 178196 206561
rect 177876 199561 178196 206325
rect 177876 199325 177918 199561
rect 178154 199325 178196 199561
rect 177876 192561 178196 199325
rect 177876 192325 177918 192561
rect 178154 192325 178196 192561
rect 177876 185561 178196 192325
rect 177876 185325 177918 185561
rect 178154 185325 178196 185561
rect 177876 178561 178196 185325
rect 177876 178325 177918 178561
rect 178154 178325 178196 178561
rect 177876 171561 178196 178325
rect 177876 171325 177918 171561
rect 178154 171325 178196 171561
rect 177876 164561 178196 171325
rect 177876 164325 177918 164561
rect 178154 164325 178196 164561
rect 177876 157561 178196 164325
rect 177876 157325 177918 157561
rect 178154 157325 178196 157561
rect 177876 150561 178196 157325
rect 177876 150325 177918 150561
rect 178154 150325 178196 150561
rect 177876 143561 178196 150325
rect 177876 143325 177918 143561
rect 178154 143325 178196 143561
rect 177876 136561 178196 143325
rect 177876 136325 177918 136561
rect 178154 136325 178196 136561
rect 177876 129561 178196 136325
rect 177876 129325 177918 129561
rect 178154 129325 178196 129561
rect 177876 122561 178196 129325
rect 177876 122325 177918 122561
rect 178154 122325 178196 122561
rect 177876 115561 178196 122325
rect 177876 115325 177918 115561
rect 178154 115325 178196 115561
rect 177876 108561 178196 115325
rect 177876 108325 177918 108561
rect 178154 108325 178196 108561
rect 177876 101561 178196 108325
rect 177876 101325 177918 101561
rect 178154 101325 178196 101561
rect 177876 94561 178196 101325
rect 177876 94325 177918 94561
rect 178154 94325 178196 94561
rect 177876 87561 178196 94325
rect 177876 87325 177918 87561
rect 178154 87325 178196 87561
rect 177876 80561 178196 87325
rect 177876 80325 177918 80561
rect 178154 80325 178196 80561
rect 177876 73561 178196 80325
rect 177876 73325 177918 73561
rect 178154 73325 178196 73561
rect 177876 66561 178196 73325
rect 177876 66325 177918 66561
rect 178154 66325 178196 66561
rect 177876 59561 178196 66325
rect 177876 59325 177918 59561
rect 178154 59325 178196 59561
rect 177876 52561 178196 59325
rect 177876 52325 177918 52561
rect 178154 52325 178196 52561
rect 177876 45561 178196 52325
rect 177876 45325 177918 45561
rect 178154 45325 178196 45561
rect 177876 38561 178196 45325
rect 177876 38325 177918 38561
rect 178154 38325 178196 38561
rect 177876 31561 178196 38325
rect 177876 31325 177918 31561
rect 178154 31325 178196 31561
rect 177876 24561 178196 31325
rect 177876 24325 177918 24561
rect 178154 24325 178196 24561
rect 177876 17561 178196 24325
rect 177876 17325 177918 17561
rect 178154 17325 178196 17561
rect 177876 10561 178196 17325
rect 177876 10325 177918 10561
rect 178154 10325 178196 10561
rect 177876 3561 178196 10325
rect 177876 3325 177918 3561
rect 178154 3325 178196 3561
rect 177876 -1706 178196 3325
rect 177876 -1942 177918 -1706
rect 178154 -1942 178196 -1706
rect 177876 -2026 178196 -1942
rect 177876 -2262 177918 -2026
rect 178154 -2262 178196 -2026
rect 177876 -2294 178196 -2262
rect 183144 705238 183464 706230
rect 183144 705002 183186 705238
rect 183422 705002 183464 705238
rect 183144 704918 183464 705002
rect 183144 704682 183186 704918
rect 183422 704682 183464 704918
rect 183144 695494 183464 704682
rect 183144 695258 183186 695494
rect 183422 695258 183464 695494
rect 183144 688494 183464 695258
rect 183144 688258 183186 688494
rect 183422 688258 183464 688494
rect 183144 681494 183464 688258
rect 183144 681258 183186 681494
rect 183422 681258 183464 681494
rect 183144 674494 183464 681258
rect 183144 674258 183186 674494
rect 183422 674258 183464 674494
rect 183144 667494 183464 674258
rect 183144 667258 183186 667494
rect 183422 667258 183464 667494
rect 183144 660494 183464 667258
rect 183144 660258 183186 660494
rect 183422 660258 183464 660494
rect 183144 653494 183464 660258
rect 183144 653258 183186 653494
rect 183422 653258 183464 653494
rect 183144 646494 183464 653258
rect 183144 646258 183186 646494
rect 183422 646258 183464 646494
rect 183144 639494 183464 646258
rect 183144 639258 183186 639494
rect 183422 639258 183464 639494
rect 183144 632494 183464 639258
rect 183144 632258 183186 632494
rect 183422 632258 183464 632494
rect 183144 625494 183464 632258
rect 183144 625258 183186 625494
rect 183422 625258 183464 625494
rect 183144 618494 183464 625258
rect 183144 618258 183186 618494
rect 183422 618258 183464 618494
rect 183144 611494 183464 618258
rect 183144 611258 183186 611494
rect 183422 611258 183464 611494
rect 183144 604494 183464 611258
rect 183144 604258 183186 604494
rect 183422 604258 183464 604494
rect 183144 597494 183464 604258
rect 183144 597258 183186 597494
rect 183422 597258 183464 597494
rect 183144 590494 183464 597258
rect 183144 590258 183186 590494
rect 183422 590258 183464 590494
rect 183144 583494 183464 590258
rect 183144 583258 183186 583494
rect 183422 583258 183464 583494
rect 183144 576494 183464 583258
rect 183144 576258 183186 576494
rect 183422 576258 183464 576494
rect 183144 569494 183464 576258
rect 183144 569258 183186 569494
rect 183422 569258 183464 569494
rect 183144 562494 183464 569258
rect 183144 562258 183186 562494
rect 183422 562258 183464 562494
rect 183144 555494 183464 562258
rect 183144 555258 183186 555494
rect 183422 555258 183464 555494
rect 183144 548494 183464 555258
rect 183144 548258 183186 548494
rect 183422 548258 183464 548494
rect 183144 541494 183464 548258
rect 183144 541258 183186 541494
rect 183422 541258 183464 541494
rect 183144 534494 183464 541258
rect 183144 534258 183186 534494
rect 183422 534258 183464 534494
rect 183144 527494 183464 534258
rect 183144 527258 183186 527494
rect 183422 527258 183464 527494
rect 183144 520494 183464 527258
rect 183144 520258 183186 520494
rect 183422 520258 183464 520494
rect 183144 513494 183464 520258
rect 183144 513258 183186 513494
rect 183422 513258 183464 513494
rect 183144 506494 183464 513258
rect 183144 506258 183186 506494
rect 183422 506258 183464 506494
rect 183144 499494 183464 506258
rect 183144 499258 183186 499494
rect 183422 499258 183464 499494
rect 183144 492494 183464 499258
rect 183144 492258 183186 492494
rect 183422 492258 183464 492494
rect 183144 485494 183464 492258
rect 183144 485258 183186 485494
rect 183422 485258 183464 485494
rect 183144 478494 183464 485258
rect 183144 478258 183186 478494
rect 183422 478258 183464 478494
rect 183144 471494 183464 478258
rect 183144 471258 183186 471494
rect 183422 471258 183464 471494
rect 183144 464494 183464 471258
rect 183144 464258 183186 464494
rect 183422 464258 183464 464494
rect 183144 457494 183464 464258
rect 183144 457258 183186 457494
rect 183422 457258 183464 457494
rect 183144 450494 183464 457258
rect 183144 450258 183186 450494
rect 183422 450258 183464 450494
rect 183144 443494 183464 450258
rect 183144 443258 183186 443494
rect 183422 443258 183464 443494
rect 183144 436494 183464 443258
rect 183144 436258 183186 436494
rect 183422 436258 183464 436494
rect 183144 429494 183464 436258
rect 183144 429258 183186 429494
rect 183422 429258 183464 429494
rect 183144 422494 183464 429258
rect 183144 422258 183186 422494
rect 183422 422258 183464 422494
rect 183144 415494 183464 422258
rect 183144 415258 183186 415494
rect 183422 415258 183464 415494
rect 183144 408494 183464 415258
rect 183144 408258 183186 408494
rect 183422 408258 183464 408494
rect 183144 401494 183464 408258
rect 183144 401258 183186 401494
rect 183422 401258 183464 401494
rect 183144 394494 183464 401258
rect 183144 394258 183186 394494
rect 183422 394258 183464 394494
rect 183144 387494 183464 394258
rect 183144 387258 183186 387494
rect 183422 387258 183464 387494
rect 183144 380494 183464 387258
rect 183144 380258 183186 380494
rect 183422 380258 183464 380494
rect 183144 373494 183464 380258
rect 183144 373258 183186 373494
rect 183422 373258 183464 373494
rect 183144 366494 183464 373258
rect 183144 366258 183186 366494
rect 183422 366258 183464 366494
rect 183144 359494 183464 366258
rect 183144 359258 183186 359494
rect 183422 359258 183464 359494
rect 183144 352494 183464 359258
rect 183144 352258 183186 352494
rect 183422 352258 183464 352494
rect 183144 345494 183464 352258
rect 183144 345258 183186 345494
rect 183422 345258 183464 345494
rect 183144 338494 183464 345258
rect 183144 338258 183186 338494
rect 183422 338258 183464 338494
rect 183144 331494 183464 338258
rect 183144 331258 183186 331494
rect 183422 331258 183464 331494
rect 183144 324494 183464 331258
rect 183144 324258 183186 324494
rect 183422 324258 183464 324494
rect 183144 317494 183464 324258
rect 183144 317258 183186 317494
rect 183422 317258 183464 317494
rect 183144 310494 183464 317258
rect 183144 310258 183186 310494
rect 183422 310258 183464 310494
rect 183144 303494 183464 310258
rect 183144 303258 183186 303494
rect 183422 303258 183464 303494
rect 183144 296494 183464 303258
rect 183144 296258 183186 296494
rect 183422 296258 183464 296494
rect 183144 289494 183464 296258
rect 183144 289258 183186 289494
rect 183422 289258 183464 289494
rect 183144 282494 183464 289258
rect 183144 282258 183186 282494
rect 183422 282258 183464 282494
rect 183144 275494 183464 282258
rect 183144 275258 183186 275494
rect 183422 275258 183464 275494
rect 183144 268494 183464 275258
rect 183144 268258 183186 268494
rect 183422 268258 183464 268494
rect 183144 261494 183464 268258
rect 183144 261258 183186 261494
rect 183422 261258 183464 261494
rect 183144 254494 183464 261258
rect 183144 254258 183186 254494
rect 183422 254258 183464 254494
rect 183144 247494 183464 254258
rect 183144 247258 183186 247494
rect 183422 247258 183464 247494
rect 183144 240494 183464 247258
rect 183144 240258 183186 240494
rect 183422 240258 183464 240494
rect 183144 233494 183464 240258
rect 183144 233258 183186 233494
rect 183422 233258 183464 233494
rect 183144 226494 183464 233258
rect 183144 226258 183186 226494
rect 183422 226258 183464 226494
rect 183144 219494 183464 226258
rect 183144 219258 183186 219494
rect 183422 219258 183464 219494
rect 183144 212494 183464 219258
rect 183144 212258 183186 212494
rect 183422 212258 183464 212494
rect 183144 205494 183464 212258
rect 183144 205258 183186 205494
rect 183422 205258 183464 205494
rect 183144 198494 183464 205258
rect 183144 198258 183186 198494
rect 183422 198258 183464 198494
rect 183144 191494 183464 198258
rect 183144 191258 183186 191494
rect 183422 191258 183464 191494
rect 183144 184494 183464 191258
rect 183144 184258 183186 184494
rect 183422 184258 183464 184494
rect 183144 177494 183464 184258
rect 183144 177258 183186 177494
rect 183422 177258 183464 177494
rect 183144 170494 183464 177258
rect 183144 170258 183186 170494
rect 183422 170258 183464 170494
rect 183144 163494 183464 170258
rect 183144 163258 183186 163494
rect 183422 163258 183464 163494
rect 183144 156494 183464 163258
rect 183144 156258 183186 156494
rect 183422 156258 183464 156494
rect 183144 149494 183464 156258
rect 183144 149258 183186 149494
rect 183422 149258 183464 149494
rect 183144 142494 183464 149258
rect 183144 142258 183186 142494
rect 183422 142258 183464 142494
rect 183144 135494 183464 142258
rect 183144 135258 183186 135494
rect 183422 135258 183464 135494
rect 183144 128494 183464 135258
rect 183144 128258 183186 128494
rect 183422 128258 183464 128494
rect 183144 121494 183464 128258
rect 183144 121258 183186 121494
rect 183422 121258 183464 121494
rect 183144 114494 183464 121258
rect 183144 114258 183186 114494
rect 183422 114258 183464 114494
rect 183144 107494 183464 114258
rect 183144 107258 183186 107494
rect 183422 107258 183464 107494
rect 183144 100494 183464 107258
rect 183144 100258 183186 100494
rect 183422 100258 183464 100494
rect 183144 93494 183464 100258
rect 183144 93258 183186 93494
rect 183422 93258 183464 93494
rect 183144 86494 183464 93258
rect 183144 86258 183186 86494
rect 183422 86258 183464 86494
rect 183144 79494 183464 86258
rect 183144 79258 183186 79494
rect 183422 79258 183464 79494
rect 183144 72494 183464 79258
rect 183144 72258 183186 72494
rect 183422 72258 183464 72494
rect 183144 65494 183464 72258
rect 183144 65258 183186 65494
rect 183422 65258 183464 65494
rect 183144 58494 183464 65258
rect 183144 58258 183186 58494
rect 183422 58258 183464 58494
rect 183144 51494 183464 58258
rect 183144 51258 183186 51494
rect 183422 51258 183464 51494
rect 183144 44494 183464 51258
rect 183144 44258 183186 44494
rect 183422 44258 183464 44494
rect 183144 37494 183464 44258
rect 183144 37258 183186 37494
rect 183422 37258 183464 37494
rect 183144 30494 183464 37258
rect 183144 30258 183186 30494
rect 183422 30258 183464 30494
rect 183144 23494 183464 30258
rect 183144 23258 183186 23494
rect 183422 23258 183464 23494
rect 183144 16494 183464 23258
rect 183144 16258 183186 16494
rect 183422 16258 183464 16494
rect 183144 9494 183464 16258
rect 183144 9258 183186 9494
rect 183422 9258 183464 9494
rect 183144 2494 183464 9258
rect 183144 2258 183186 2494
rect 183422 2258 183464 2494
rect 183144 -746 183464 2258
rect 183144 -982 183186 -746
rect 183422 -982 183464 -746
rect 183144 -1066 183464 -982
rect 183144 -1302 183186 -1066
rect 183422 -1302 183464 -1066
rect 183144 -2294 183464 -1302
rect 184876 706198 185196 706230
rect 184876 705962 184918 706198
rect 185154 705962 185196 706198
rect 184876 705878 185196 705962
rect 184876 705642 184918 705878
rect 185154 705642 185196 705878
rect 184876 696561 185196 705642
rect 184876 696325 184918 696561
rect 185154 696325 185196 696561
rect 184876 689561 185196 696325
rect 184876 689325 184918 689561
rect 185154 689325 185196 689561
rect 184876 682561 185196 689325
rect 184876 682325 184918 682561
rect 185154 682325 185196 682561
rect 184876 675561 185196 682325
rect 184876 675325 184918 675561
rect 185154 675325 185196 675561
rect 184876 668561 185196 675325
rect 184876 668325 184918 668561
rect 185154 668325 185196 668561
rect 184876 661561 185196 668325
rect 184876 661325 184918 661561
rect 185154 661325 185196 661561
rect 184876 654561 185196 661325
rect 184876 654325 184918 654561
rect 185154 654325 185196 654561
rect 184876 647561 185196 654325
rect 184876 647325 184918 647561
rect 185154 647325 185196 647561
rect 184876 640561 185196 647325
rect 184876 640325 184918 640561
rect 185154 640325 185196 640561
rect 184876 633561 185196 640325
rect 184876 633325 184918 633561
rect 185154 633325 185196 633561
rect 184876 626561 185196 633325
rect 184876 626325 184918 626561
rect 185154 626325 185196 626561
rect 184876 619561 185196 626325
rect 184876 619325 184918 619561
rect 185154 619325 185196 619561
rect 184876 612561 185196 619325
rect 184876 612325 184918 612561
rect 185154 612325 185196 612561
rect 184876 605561 185196 612325
rect 184876 605325 184918 605561
rect 185154 605325 185196 605561
rect 184876 598561 185196 605325
rect 184876 598325 184918 598561
rect 185154 598325 185196 598561
rect 184876 591561 185196 598325
rect 184876 591325 184918 591561
rect 185154 591325 185196 591561
rect 184876 584561 185196 591325
rect 184876 584325 184918 584561
rect 185154 584325 185196 584561
rect 184876 577561 185196 584325
rect 184876 577325 184918 577561
rect 185154 577325 185196 577561
rect 184876 570561 185196 577325
rect 184876 570325 184918 570561
rect 185154 570325 185196 570561
rect 184876 563561 185196 570325
rect 184876 563325 184918 563561
rect 185154 563325 185196 563561
rect 184876 556561 185196 563325
rect 184876 556325 184918 556561
rect 185154 556325 185196 556561
rect 184876 549561 185196 556325
rect 184876 549325 184918 549561
rect 185154 549325 185196 549561
rect 184876 542561 185196 549325
rect 184876 542325 184918 542561
rect 185154 542325 185196 542561
rect 184876 535561 185196 542325
rect 184876 535325 184918 535561
rect 185154 535325 185196 535561
rect 184876 528561 185196 535325
rect 184876 528325 184918 528561
rect 185154 528325 185196 528561
rect 184876 521561 185196 528325
rect 184876 521325 184918 521561
rect 185154 521325 185196 521561
rect 184876 514561 185196 521325
rect 184876 514325 184918 514561
rect 185154 514325 185196 514561
rect 184876 507561 185196 514325
rect 184876 507325 184918 507561
rect 185154 507325 185196 507561
rect 184876 500561 185196 507325
rect 184876 500325 184918 500561
rect 185154 500325 185196 500561
rect 184876 493561 185196 500325
rect 184876 493325 184918 493561
rect 185154 493325 185196 493561
rect 184876 486561 185196 493325
rect 184876 486325 184918 486561
rect 185154 486325 185196 486561
rect 184876 479561 185196 486325
rect 184876 479325 184918 479561
rect 185154 479325 185196 479561
rect 184876 472561 185196 479325
rect 184876 472325 184918 472561
rect 185154 472325 185196 472561
rect 184876 465561 185196 472325
rect 184876 465325 184918 465561
rect 185154 465325 185196 465561
rect 184876 458561 185196 465325
rect 184876 458325 184918 458561
rect 185154 458325 185196 458561
rect 184876 451561 185196 458325
rect 184876 451325 184918 451561
rect 185154 451325 185196 451561
rect 184876 444561 185196 451325
rect 184876 444325 184918 444561
rect 185154 444325 185196 444561
rect 184876 437561 185196 444325
rect 184876 437325 184918 437561
rect 185154 437325 185196 437561
rect 184876 430561 185196 437325
rect 184876 430325 184918 430561
rect 185154 430325 185196 430561
rect 184876 423561 185196 430325
rect 184876 423325 184918 423561
rect 185154 423325 185196 423561
rect 184876 416561 185196 423325
rect 184876 416325 184918 416561
rect 185154 416325 185196 416561
rect 184876 409561 185196 416325
rect 184876 409325 184918 409561
rect 185154 409325 185196 409561
rect 184876 402561 185196 409325
rect 184876 402325 184918 402561
rect 185154 402325 185196 402561
rect 184876 395561 185196 402325
rect 184876 395325 184918 395561
rect 185154 395325 185196 395561
rect 184876 388561 185196 395325
rect 184876 388325 184918 388561
rect 185154 388325 185196 388561
rect 184876 381561 185196 388325
rect 184876 381325 184918 381561
rect 185154 381325 185196 381561
rect 184876 374561 185196 381325
rect 184876 374325 184918 374561
rect 185154 374325 185196 374561
rect 184876 367561 185196 374325
rect 184876 367325 184918 367561
rect 185154 367325 185196 367561
rect 184876 360561 185196 367325
rect 184876 360325 184918 360561
rect 185154 360325 185196 360561
rect 184876 353561 185196 360325
rect 184876 353325 184918 353561
rect 185154 353325 185196 353561
rect 184876 346561 185196 353325
rect 184876 346325 184918 346561
rect 185154 346325 185196 346561
rect 184876 339561 185196 346325
rect 184876 339325 184918 339561
rect 185154 339325 185196 339561
rect 184876 332561 185196 339325
rect 184876 332325 184918 332561
rect 185154 332325 185196 332561
rect 184876 325561 185196 332325
rect 184876 325325 184918 325561
rect 185154 325325 185196 325561
rect 184876 318561 185196 325325
rect 184876 318325 184918 318561
rect 185154 318325 185196 318561
rect 184876 311561 185196 318325
rect 184876 311325 184918 311561
rect 185154 311325 185196 311561
rect 184876 304561 185196 311325
rect 184876 304325 184918 304561
rect 185154 304325 185196 304561
rect 184876 297561 185196 304325
rect 184876 297325 184918 297561
rect 185154 297325 185196 297561
rect 184876 290561 185196 297325
rect 184876 290325 184918 290561
rect 185154 290325 185196 290561
rect 184876 283561 185196 290325
rect 184876 283325 184918 283561
rect 185154 283325 185196 283561
rect 184876 276561 185196 283325
rect 184876 276325 184918 276561
rect 185154 276325 185196 276561
rect 184876 269561 185196 276325
rect 184876 269325 184918 269561
rect 185154 269325 185196 269561
rect 184876 262561 185196 269325
rect 184876 262325 184918 262561
rect 185154 262325 185196 262561
rect 184876 255561 185196 262325
rect 184876 255325 184918 255561
rect 185154 255325 185196 255561
rect 184876 248561 185196 255325
rect 184876 248325 184918 248561
rect 185154 248325 185196 248561
rect 184876 241561 185196 248325
rect 184876 241325 184918 241561
rect 185154 241325 185196 241561
rect 184876 234561 185196 241325
rect 184876 234325 184918 234561
rect 185154 234325 185196 234561
rect 184876 227561 185196 234325
rect 184876 227325 184918 227561
rect 185154 227325 185196 227561
rect 184876 220561 185196 227325
rect 184876 220325 184918 220561
rect 185154 220325 185196 220561
rect 184876 213561 185196 220325
rect 184876 213325 184918 213561
rect 185154 213325 185196 213561
rect 184876 206561 185196 213325
rect 184876 206325 184918 206561
rect 185154 206325 185196 206561
rect 184876 199561 185196 206325
rect 184876 199325 184918 199561
rect 185154 199325 185196 199561
rect 184876 192561 185196 199325
rect 184876 192325 184918 192561
rect 185154 192325 185196 192561
rect 184876 185561 185196 192325
rect 184876 185325 184918 185561
rect 185154 185325 185196 185561
rect 184876 178561 185196 185325
rect 184876 178325 184918 178561
rect 185154 178325 185196 178561
rect 184876 171561 185196 178325
rect 184876 171325 184918 171561
rect 185154 171325 185196 171561
rect 184876 164561 185196 171325
rect 184876 164325 184918 164561
rect 185154 164325 185196 164561
rect 184876 157561 185196 164325
rect 184876 157325 184918 157561
rect 185154 157325 185196 157561
rect 184876 150561 185196 157325
rect 184876 150325 184918 150561
rect 185154 150325 185196 150561
rect 184876 143561 185196 150325
rect 184876 143325 184918 143561
rect 185154 143325 185196 143561
rect 184876 136561 185196 143325
rect 184876 136325 184918 136561
rect 185154 136325 185196 136561
rect 184876 129561 185196 136325
rect 184876 129325 184918 129561
rect 185154 129325 185196 129561
rect 184876 122561 185196 129325
rect 184876 122325 184918 122561
rect 185154 122325 185196 122561
rect 184876 115561 185196 122325
rect 184876 115325 184918 115561
rect 185154 115325 185196 115561
rect 184876 108561 185196 115325
rect 184876 108325 184918 108561
rect 185154 108325 185196 108561
rect 184876 101561 185196 108325
rect 184876 101325 184918 101561
rect 185154 101325 185196 101561
rect 184876 94561 185196 101325
rect 184876 94325 184918 94561
rect 185154 94325 185196 94561
rect 184876 87561 185196 94325
rect 184876 87325 184918 87561
rect 185154 87325 185196 87561
rect 184876 80561 185196 87325
rect 184876 80325 184918 80561
rect 185154 80325 185196 80561
rect 184876 73561 185196 80325
rect 184876 73325 184918 73561
rect 185154 73325 185196 73561
rect 184876 66561 185196 73325
rect 184876 66325 184918 66561
rect 185154 66325 185196 66561
rect 184876 59561 185196 66325
rect 184876 59325 184918 59561
rect 185154 59325 185196 59561
rect 184876 52561 185196 59325
rect 184876 52325 184918 52561
rect 185154 52325 185196 52561
rect 184876 45561 185196 52325
rect 184876 45325 184918 45561
rect 185154 45325 185196 45561
rect 184876 38561 185196 45325
rect 184876 38325 184918 38561
rect 185154 38325 185196 38561
rect 184876 31561 185196 38325
rect 184876 31325 184918 31561
rect 185154 31325 185196 31561
rect 184876 24561 185196 31325
rect 184876 24325 184918 24561
rect 185154 24325 185196 24561
rect 184876 17561 185196 24325
rect 184876 17325 184918 17561
rect 185154 17325 185196 17561
rect 184876 10561 185196 17325
rect 184876 10325 184918 10561
rect 185154 10325 185196 10561
rect 184876 3561 185196 10325
rect 184876 3325 184918 3561
rect 185154 3325 185196 3561
rect 184876 -1706 185196 3325
rect 184876 -1942 184918 -1706
rect 185154 -1942 185196 -1706
rect 184876 -2026 185196 -1942
rect 184876 -2262 184918 -2026
rect 185154 -2262 185196 -2026
rect 184876 -2294 185196 -2262
rect 190144 705238 190464 706230
rect 190144 705002 190186 705238
rect 190422 705002 190464 705238
rect 190144 704918 190464 705002
rect 190144 704682 190186 704918
rect 190422 704682 190464 704918
rect 190144 695494 190464 704682
rect 190144 695258 190186 695494
rect 190422 695258 190464 695494
rect 190144 688494 190464 695258
rect 190144 688258 190186 688494
rect 190422 688258 190464 688494
rect 190144 681494 190464 688258
rect 190144 681258 190186 681494
rect 190422 681258 190464 681494
rect 190144 674494 190464 681258
rect 190144 674258 190186 674494
rect 190422 674258 190464 674494
rect 190144 667494 190464 674258
rect 190144 667258 190186 667494
rect 190422 667258 190464 667494
rect 190144 660494 190464 667258
rect 190144 660258 190186 660494
rect 190422 660258 190464 660494
rect 190144 653494 190464 660258
rect 190144 653258 190186 653494
rect 190422 653258 190464 653494
rect 190144 646494 190464 653258
rect 190144 646258 190186 646494
rect 190422 646258 190464 646494
rect 190144 639494 190464 646258
rect 190144 639258 190186 639494
rect 190422 639258 190464 639494
rect 190144 632494 190464 639258
rect 190144 632258 190186 632494
rect 190422 632258 190464 632494
rect 190144 625494 190464 632258
rect 190144 625258 190186 625494
rect 190422 625258 190464 625494
rect 190144 618494 190464 625258
rect 190144 618258 190186 618494
rect 190422 618258 190464 618494
rect 190144 611494 190464 618258
rect 190144 611258 190186 611494
rect 190422 611258 190464 611494
rect 190144 604494 190464 611258
rect 190144 604258 190186 604494
rect 190422 604258 190464 604494
rect 190144 597494 190464 604258
rect 190144 597258 190186 597494
rect 190422 597258 190464 597494
rect 190144 590494 190464 597258
rect 190144 590258 190186 590494
rect 190422 590258 190464 590494
rect 190144 583494 190464 590258
rect 190144 583258 190186 583494
rect 190422 583258 190464 583494
rect 190144 576494 190464 583258
rect 190144 576258 190186 576494
rect 190422 576258 190464 576494
rect 190144 569494 190464 576258
rect 190144 569258 190186 569494
rect 190422 569258 190464 569494
rect 190144 562494 190464 569258
rect 190144 562258 190186 562494
rect 190422 562258 190464 562494
rect 190144 555494 190464 562258
rect 190144 555258 190186 555494
rect 190422 555258 190464 555494
rect 190144 548494 190464 555258
rect 190144 548258 190186 548494
rect 190422 548258 190464 548494
rect 190144 541494 190464 548258
rect 190144 541258 190186 541494
rect 190422 541258 190464 541494
rect 190144 534494 190464 541258
rect 190144 534258 190186 534494
rect 190422 534258 190464 534494
rect 190144 527494 190464 534258
rect 190144 527258 190186 527494
rect 190422 527258 190464 527494
rect 190144 520494 190464 527258
rect 190144 520258 190186 520494
rect 190422 520258 190464 520494
rect 190144 513494 190464 520258
rect 190144 513258 190186 513494
rect 190422 513258 190464 513494
rect 190144 506494 190464 513258
rect 190144 506258 190186 506494
rect 190422 506258 190464 506494
rect 190144 499494 190464 506258
rect 190144 499258 190186 499494
rect 190422 499258 190464 499494
rect 190144 492494 190464 499258
rect 190144 492258 190186 492494
rect 190422 492258 190464 492494
rect 190144 485494 190464 492258
rect 190144 485258 190186 485494
rect 190422 485258 190464 485494
rect 190144 478494 190464 485258
rect 190144 478258 190186 478494
rect 190422 478258 190464 478494
rect 190144 471494 190464 478258
rect 190144 471258 190186 471494
rect 190422 471258 190464 471494
rect 190144 464494 190464 471258
rect 190144 464258 190186 464494
rect 190422 464258 190464 464494
rect 190144 457494 190464 464258
rect 190144 457258 190186 457494
rect 190422 457258 190464 457494
rect 190144 450494 190464 457258
rect 190144 450258 190186 450494
rect 190422 450258 190464 450494
rect 190144 443494 190464 450258
rect 190144 443258 190186 443494
rect 190422 443258 190464 443494
rect 190144 436494 190464 443258
rect 190144 436258 190186 436494
rect 190422 436258 190464 436494
rect 190144 429494 190464 436258
rect 190144 429258 190186 429494
rect 190422 429258 190464 429494
rect 190144 422494 190464 429258
rect 190144 422258 190186 422494
rect 190422 422258 190464 422494
rect 190144 415494 190464 422258
rect 190144 415258 190186 415494
rect 190422 415258 190464 415494
rect 190144 408494 190464 415258
rect 190144 408258 190186 408494
rect 190422 408258 190464 408494
rect 190144 401494 190464 408258
rect 190144 401258 190186 401494
rect 190422 401258 190464 401494
rect 190144 394494 190464 401258
rect 190144 394258 190186 394494
rect 190422 394258 190464 394494
rect 190144 387494 190464 394258
rect 190144 387258 190186 387494
rect 190422 387258 190464 387494
rect 190144 380494 190464 387258
rect 190144 380258 190186 380494
rect 190422 380258 190464 380494
rect 190144 373494 190464 380258
rect 190144 373258 190186 373494
rect 190422 373258 190464 373494
rect 190144 366494 190464 373258
rect 190144 366258 190186 366494
rect 190422 366258 190464 366494
rect 190144 359494 190464 366258
rect 190144 359258 190186 359494
rect 190422 359258 190464 359494
rect 190144 352494 190464 359258
rect 190144 352258 190186 352494
rect 190422 352258 190464 352494
rect 190144 345494 190464 352258
rect 190144 345258 190186 345494
rect 190422 345258 190464 345494
rect 190144 338494 190464 345258
rect 190144 338258 190186 338494
rect 190422 338258 190464 338494
rect 190144 331494 190464 338258
rect 190144 331258 190186 331494
rect 190422 331258 190464 331494
rect 190144 324494 190464 331258
rect 190144 324258 190186 324494
rect 190422 324258 190464 324494
rect 190144 317494 190464 324258
rect 190144 317258 190186 317494
rect 190422 317258 190464 317494
rect 190144 310494 190464 317258
rect 190144 310258 190186 310494
rect 190422 310258 190464 310494
rect 190144 303494 190464 310258
rect 190144 303258 190186 303494
rect 190422 303258 190464 303494
rect 190144 296494 190464 303258
rect 190144 296258 190186 296494
rect 190422 296258 190464 296494
rect 190144 289494 190464 296258
rect 190144 289258 190186 289494
rect 190422 289258 190464 289494
rect 190144 282494 190464 289258
rect 190144 282258 190186 282494
rect 190422 282258 190464 282494
rect 190144 275494 190464 282258
rect 190144 275258 190186 275494
rect 190422 275258 190464 275494
rect 190144 268494 190464 275258
rect 190144 268258 190186 268494
rect 190422 268258 190464 268494
rect 190144 261494 190464 268258
rect 190144 261258 190186 261494
rect 190422 261258 190464 261494
rect 190144 254494 190464 261258
rect 190144 254258 190186 254494
rect 190422 254258 190464 254494
rect 190144 247494 190464 254258
rect 190144 247258 190186 247494
rect 190422 247258 190464 247494
rect 190144 240494 190464 247258
rect 190144 240258 190186 240494
rect 190422 240258 190464 240494
rect 190144 233494 190464 240258
rect 190144 233258 190186 233494
rect 190422 233258 190464 233494
rect 190144 226494 190464 233258
rect 190144 226258 190186 226494
rect 190422 226258 190464 226494
rect 190144 219494 190464 226258
rect 190144 219258 190186 219494
rect 190422 219258 190464 219494
rect 190144 212494 190464 219258
rect 190144 212258 190186 212494
rect 190422 212258 190464 212494
rect 190144 205494 190464 212258
rect 190144 205258 190186 205494
rect 190422 205258 190464 205494
rect 190144 198494 190464 205258
rect 190144 198258 190186 198494
rect 190422 198258 190464 198494
rect 190144 191494 190464 198258
rect 190144 191258 190186 191494
rect 190422 191258 190464 191494
rect 190144 184494 190464 191258
rect 190144 184258 190186 184494
rect 190422 184258 190464 184494
rect 190144 177494 190464 184258
rect 190144 177258 190186 177494
rect 190422 177258 190464 177494
rect 190144 170494 190464 177258
rect 190144 170258 190186 170494
rect 190422 170258 190464 170494
rect 190144 163494 190464 170258
rect 190144 163258 190186 163494
rect 190422 163258 190464 163494
rect 190144 156494 190464 163258
rect 190144 156258 190186 156494
rect 190422 156258 190464 156494
rect 190144 149494 190464 156258
rect 190144 149258 190186 149494
rect 190422 149258 190464 149494
rect 190144 142494 190464 149258
rect 190144 142258 190186 142494
rect 190422 142258 190464 142494
rect 190144 135494 190464 142258
rect 190144 135258 190186 135494
rect 190422 135258 190464 135494
rect 190144 128494 190464 135258
rect 190144 128258 190186 128494
rect 190422 128258 190464 128494
rect 190144 121494 190464 128258
rect 190144 121258 190186 121494
rect 190422 121258 190464 121494
rect 190144 114494 190464 121258
rect 190144 114258 190186 114494
rect 190422 114258 190464 114494
rect 190144 107494 190464 114258
rect 190144 107258 190186 107494
rect 190422 107258 190464 107494
rect 190144 100494 190464 107258
rect 190144 100258 190186 100494
rect 190422 100258 190464 100494
rect 190144 93494 190464 100258
rect 190144 93258 190186 93494
rect 190422 93258 190464 93494
rect 190144 86494 190464 93258
rect 190144 86258 190186 86494
rect 190422 86258 190464 86494
rect 190144 79494 190464 86258
rect 190144 79258 190186 79494
rect 190422 79258 190464 79494
rect 190144 72494 190464 79258
rect 190144 72258 190186 72494
rect 190422 72258 190464 72494
rect 190144 65494 190464 72258
rect 190144 65258 190186 65494
rect 190422 65258 190464 65494
rect 190144 58494 190464 65258
rect 190144 58258 190186 58494
rect 190422 58258 190464 58494
rect 190144 51494 190464 58258
rect 190144 51258 190186 51494
rect 190422 51258 190464 51494
rect 190144 44494 190464 51258
rect 190144 44258 190186 44494
rect 190422 44258 190464 44494
rect 190144 37494 190464 44258
rect 190144 37258 190186 37494
rect 190422 37258 190464 37494
rect 190144 30494 190464 37258
rect 190144 30258 190186 30494
rect 190422 30258 190464 30494
rect 190144 23494 190464 30258
rect 190144 23258 190186 23494
rect 190422 23258 190464 23494
rect 190144 16494 190464 23258
rect 190144 16258 190186 16494
rect 190422 16258 190464 16494
rect 190144 9494 190464 16258
rect 190144 9258 190186 9494
rect 190422 9258 190464 9494
rect 190144 2494 190464 9258
rect 190144 2258 190186 2494
rect 190422 2258 190464 2494
rect 190144 -746 190464 2258
rect 190144 -982 190186 -746
rect 190422 -982 190464 -746
rect 190144 -1066 190464 -982
rect 190144 -1302 190186 -1066
rect 190422 -1302 190464 -1066
rect 190144 -2294 190464 -1302
rect 191876 706198 192196 706230
rect 191876 705962 191918 706198
rect 192154 705962 192196 706198
rect 191876 705878 192196 705962
rect 191876 705642 191918 705878
rect 192154 705642 192196 705878
rect 191876 696561 192196 705642
rect 191876 696325 191918 696561
rect 192154 696325 192196 696561
rect 191876 689561 192196 696325
rect 191876 689325 191918 689561
rect 192154 689325 192196 689561
rect 191876 682561 192196 689325
rect 191876 682325 191918 682561
rect 192154 682325 192196 682561
rect 191876 675561 192196 682325
rect 191876 675325 191918 675561
rect 192154 675325 192196 675561
rect 191876 668561 192196 675325
rect 191876 668325 191918 668561
rect 192154 668325 192196 668561
rect 191876 661561 192196 668325
rect 191876 661325 191918 661561
rect 192154 661325 192196 661561
rect 191876 654561 192196 661325
rect 191876 654325 191918 654561
rect 192154 654325 192196 654561
rect 191876 647561 192196 654325
rect 191876 647325 191918 647561
rect 192154 647325 192196 647561
rect 191876 640561 192196 647325
rect 191876 640325 191918 640561
rect 192154 640325 192196 640561
rect 191876 633561 192196 640325
rect 191876 633325 191918 633561
rect 192154 633325 192196 633561
rect 191876 626561 192196 633325
rect 191876 626325 191918 626561
rect 192154 626325 192196 626561
rect 191876 619561 192196 626325
rect 191876 619325 191918 619561
rect 192154 619325 192196 619561
rect 191876 612561 192196 619325
rect 191876 612325 191918 612561
rect 192154 612325 192196 612561
rect 191876 605561 192196 612325
rect 191876 605325 191918 605561
rect 192154 605325 192196 605561
rect 191876 598561 192196 605325
rect 191876 598325 191918 598561
rect 192154 598325 192196 598561
rect 191876 591561 192196 598325
rect 191876 591325 191918 591561
rect 192154 591325 192196 591561
rect 191876 584561 192196 591325
rect 191876 584325 191918 584561
rect 192154 584325 192196 584561
rect 191876 577561 192196 584325
rect 191876 577325 191918 577561
rect 192154 577325 192196 577561
rect 191876 570561 192196 577325
rect 191876 570325 191918 570561
rect 192154 570325 192196 570561
rect 191876 563561 192196 570325
rect 191876 563325 191918 563561
rect 192154 563325 192196 563561
rect 191876 556561 192196 563325
rect 191876 556325 191918 556561
rect 192154 556325 192196 556561
rect 191876 549561 192196 556325
rect 191876 549325 191918 549561
rect 192154 549325 192196 549561
rect 191876 542561 192196 549325
rect 191876 542325 191918 542561
rect 192154 542325 192196 542561
rect 191876 535561 192196 542325
rect 191876 535325 191918 535561
rect 192154 535325 192196 535561
rect 191876 528561 192196 535325
rect 191876 528325 191918 528561
rect 192154 528325 192196 528561
rect 191876 521561 192196 528325
rect 191876 521325 191918 521561
rect 192154 521325 192196 521561
rect 191876 514561 192196 521325
rect 191876 514325 191918 514561
rect 192154 514325 192196 514561
rect 191876 507561 192196 514325
rect 191876 507325 191918 507561
rect 192154 507325 192196 507561
rect 191876 500561 192196 507325
rect 191876 500325 191918 500561
rect 192154 500325 192196 500561
rect 191876 493561 192196 500325
rect 191876 493325 191918 493561
rect 192154 493325 192196 493561
rect 191876 486561 192196 493325
rect 191876 486325 191918 486561
rect 192154 486325 192196 486561
rect 191876 479561 192196 486325
rect 191876 479325 191918 479561
rect 192154 479325 192196 479561
rect 191876 472561 192196 479325
rect 191876 472325 191918 472561
rect 192154 472325 192196 472561
rect 191876 465561 192196 472325
rect 191876 465325 191918 465561
rect 192154 465325 192196 465561
rect 191876 458561 192196 465325
rect 191876 458325 191918 458561
rect 192154 458325 192196 458561
rect 191876 451561 192196 458325
rect 191876 451325 191918 451561
rect 192154 451325 192196 451561
rect 191876 444561 192196 451325
rect 191876 444325 191918 444561
rect 192154 444325 192196 444561
rect 191876 437561 192196 444325
rect 191876 437325 191918 437561
rect 192154 437325 192196 437561
rect 191876 430561 192196 437325
rect 191876 430325 191918 430561
rect 192154 430325 192196 430561
rect 191876 423561 192196 430325
rect 191876 423325 191918 423561
rect 192154 423325 192196 423561
rect 191876 416561 192196 423325
rect 191876 416325 191918 416561
rect 192154 416325 192196 416561
rect 191876 409561 192196 416325
rect 191876 409325 191918 409561
rect 192154 409325 192196 409561
rect 191876 402561 192196 409325
rect 191876 402325 191918 402561
rect 192154 402325 192196 402561
rect 191876 395561 192196 402325
rect 191876 395325 191918 395561
rect 192154 395325 192196 395561
rect 191876 388561 192196 395325
rect 191876 388325 191918 388561
rect 192154 388325 192196 388561
rect 191876 381561 192196 388325
rect 191876 381325 191918 381561
rect 192154 381325 192196 381561
rect 191876 374561 192196 381325
rect 191876 374325 191918 374561
rect 192154 374325 192196 374561
rect 191876 367561 192196 374325
rect 191876 367325 191918 367561
rect 192154 367325 192196 367561
rect 191876 360561 192196 367325
rect 191876 360325 191918 360561
rect 192154 360325 192196 360561
rect 191876 353561 192196 360325
rect 191876 353325 191918 353561
rect 192154 353325 192196 353561
rect 191876 346561 192196 353325
rect 191876 346325 191918 346561
rect 192154 346325 192196 346561
rect 191876 339561 192196 346325
rect 191876 339325 191918 339561
rect 192154 339325 192196 339561
rect 191876 332561 192196 339325
rect 191876 332325 191918 332561
rect 192154 332325 192196 332561
rect 191876 325561 192196 332325
rect 191876 325325 191918 325561
rect 192154 325325 192196 325561
rect 191876 318561 192196 325325
rect 191876 318325 191918 318561
rect 192154 318325 192196 318561
rect 191876 311561 192196 318325
rect 191876 311325 191918 311561
rect 192154 311325 192196 311561
rect 191876 304561 192196 311325
rect 191876 304325 191918 304561
rect 192154 304325 192196 304561
rect 191876 297561 192196 304325
rect 191876 297325 191918 297561
rect 192154 297325 192196 297561
rect 191876 290561 192196 297325
rect 191876 290325 191918 290561
rect 192154 290325 192196 290561
rect 191876 283561 192196 290325
rect 191876 283325 191918 283561
rect 192154 283325 192196 283561
rect 191876 276561 192196 283325
rect 191876 276325 191918 276561
rect 192154 276325 192196 276561
rect 191876 269561 192196 276325
rect 191876 269325 191918 269561
rect 192154 269325 192196 269561
rect 191876 262561 192196 269325
rect 191876 262325 191918 262561
rect 192154 262325 192196 262561
rect 191876 255561 192196 262325
rect 191876 255325 191918 255561
rect 192154 255325 192196 255561
rect 191876 248561 192196 255325
rect 191876 248325 191918 248561
rect 192154 248325 192196 248561
rect 191876 241561 192196 248325
rect 191876 241325 191918 241561
rect 192154 241325 192196 241561
rect 191876 234561 192196 241325
rect 191876 234325 191918 234561
rect 192154 234325 192196 234561
rect 191876 227561 192196 234325
rect 191876 227325 191918 227561
rect 192154 227325 192196 227561
rect 191876 220561 192196 227325
rect 191876 220325 191918 220561
rect 192154 220325 192196 220561
rect 191876 213561 192196 220325
rect 191876 213325 191918 213561
rect 192154 213325 192196 213561
rect 191876 206561 192196 213325
rect 191876 206325 191918 206561
rect 192154 206325 192196 206561
rect 191876 199561 192196 206325
rect 191876 199325 191918 199561
rect 192154 199325 192196 199561
rect 191876 192561 192196 199325
rect 191876 192325 191918 192561
rect 192154 192325 192196 192561
rect 191876 185561 192196 192325
rect 191876 185325 191918 185561
rect 192154 185325 192196 185561
rect 191876 178561 192196 185325
rect 191876 178325 191918 178561
rect 192154 178325 192196 178561
rect 191876 171561 192196 178325
rect 191876 171325 191918 171561
rect 192154 171325 192196 171561
rect 191876 164561 192196 171325
rect 191876 164325 191918 164561
rect 192154 164325 192196 164561
rect 191876 157561 192196 164325
rect 191876 157325 191918 157561
rect 192154 157325 192196 157561
rect 191876 150561 192196 157325
rect 191876 150325 191918 150561
rect 192154 150325 192196 150561
rect 191876 143561 192196 150325
rect 191876 143325 191918 143561
rect 192154 143325 192196 143561
rect 191876 136561 192196 143325
rect 191876 136325 191918 136561
rect 192154 136325 192196 136561
rect 191876 129561 192196 136325
rect 191876 129325 191918 129561
rect 192154 129325 192196 129561
rect 191876 122561 192196 129325
rect 191876 122325 191918 122561
rect 192154 122325 192196 122561
rect 191876 115561 192196 122325
rect 191876 115325 191918 115561
rect 192154 115325 192196 115561
rect 191876 108561 192196 115325
rect 191876 108325 191918 108561
rect 192154 108325 192196 108561
rect 191876 101561 192196 108325
rect 191876 101325 191918 101561
rect 192154 101325 192196 101561
rect 191876 94561 192196 101325
rect 191876 94325 191918 94561
rect 192154 94325 192196 94561
rect 191876 87561 192196 94325
rect 191876 87325 191918 87561
rect 192154 87325 192196 87561
rect 191876 80561 192196 87325
rect 191876 80325 191918 80561
rect 192154 80325 192196 80561
rect 191876 73561 192196 80325
rect 191876 73325 191918 73561
rect 192154 73325 192196 73561
rect 191876 66561 192196 73325
rect 191876 66325 191918 66561
rect 192154 66325 192196 66561
rect 191876 59561 192196 66325
rect 191876 59325 191918 59561
rect 192154 59325 192196 59561
rect 191876 52561 192196 59325
rect 191876 52325 191918 52561
rect 192154 52325 192196 52561
rect 191876 45561 192196 52325
rect 191876 45325 191918 45561
rect 192154 45325 192196 45561
rect 191876 38561 192196 45325
rect 191876 38325 191918 38561
rect 192154 38325 192196 38561
rect 191876 31561 192196 38325
rect 191876 31325 191918 31561
rect 192154 31325 192196 31561
rect 191876 24561 192196 31325
rect 191876 24325 191918 24561
rect 192154 24325 192196 24561
rect 191876 17561 192196 24325
rect 191876 17325 191918 17561
rect 192154 17325 192196 17561
rect 191876 10561 192196 17325
rect 191876 10325 191918 10561
rect 192154 10325 192196 10561
rect 191876 3561 192196 10325
rect 191876 3325 191918 3561
rect 192154 3325 192196 3561
rect 191876 -1706 192196 3325
rect 191876 -1942 191918 -1706
rect 192154 -1942 192196 -1706
rect 191876 -2026 192196 -1942
rect 191876 -2262 191918 -2026
rect 192154 -2262 192196 -2026
rect 191876 -2294 192196 -2262
rect 197144 705238 197464 706230
rect 197144 705002 197186 705238
rect 197422 705002 197464 705238
rect 197144 704918 197464 705002
rect 197144 704682 197186 704918
rect 197422 704682 197464 704918
rect 197144 695494 197464 704682
rect 197144 695258 197186 695494
rect 197422 695258 197464 695494
rect 197144 688494 197464 695258
rect 197144 688258 197186 688494
rect 197422 688258 197464 688494
rect 197144 681494 197464 688258
rect 197144 681258 197186 681494
rect 197422 681258 197464 681494
rect 197144 674494 197464 681258
rect 197144 674258 197186 674494
rect 197422 674258 197464 674494
rect 197144 667494 197464 674258
rect 197144 667258 197186 667494
rect 197422 667258 197464 667494
rect 197144 660494 197464 667258
rect 197144 660258 197186 660494
rect 197422 660258 197464 660494
rect 197144 653494 197464 660258
rect 197144 653258 197186 653494
rect 197422 653258 197464 653494
rect 197144 646494 197464 653258
rect 197144 646258 197186 646494
rect 197422 646258 197464 646494
rect 197144 639494 197464 646258
rect 197144 639258 197186 639494
rect 197422 639258 197464 639494
rect 197144 632494 197464 639258
rect 197144 632258 197186 632494
rect 197422 632258 197464 632494
rect 197144 625494 197464 632258
rect 197144 625258 197186 625494
rect 197422 625258 197464 625494
rect 197144 618494 197464 625258
rect 197144 618258 197186 618494
rect 197422 618258 197464 618494
rect 197144 611494 197464 618258
rect 197144 611258 197186 611494
rect 197422 611258 197464 611494
rect 197144 604494 197464 611258
rect 197144 604258 197186 604494
rect 197422 604258 197464 604494
rect 197144 597494 197464 604258
rect 197144 597258 197186 597494
rect 197422 597258 197464 597494
rect 197144 590494 197464 597258
rect 197144 590258 197186 590494
rect 197422 590258 197464 590494
rect 197144 583494 197464 590258
rect 197144 583258 197186 583494
rect 197422 583258 197464 583494
rect 197144 576494 197464 583258
rect 197144 576258 197186 576494
rect 197422 576258 197464 576494
rect 197144 569494 197464 576258
rect 197144 569258 197186 569494
rect 197422 569258 197464 569494
rect 197144 562494 197464 569258
rect 197144 562258 197186 562494
rect 197422 562258 197464 562494
rect 197144 555494 197464 562258
rect 197144 555258 197186 555494
rect 197422 555258 197464 555494
rect 197144 548494 197464 555258
rect 197144 548258 197186 548494
rect 197422 548258 197464 548494
rect 197144 541494 197464 548258
rect 197144 541258 197186 541494
rect 197422 541258 197464 541494
rect 197144 534494 197464 541258
rect 197144 534258 197186 534494
rect 197422 534258 197464 534494
rect 197144 527494 197464 534258
rect 197144 527258 197186 527494
rect 197422 527258 197464 527494
rect 197144 520494 197464 527258
rect 197144 520258 197186 520494
rect 197422 520258 197464 520494
rect 197144 513494 197464 520258
rect 197144 513258 197186 513494
rect 197422 513258 197464 513494
rect 197144 506494 197464 513258
rect 197144 506258 197186 506494
rect 197422 506258 197464 506494
rect 197144 499494 197464 506258
rect 197144 499258 197186 499494
rect 197422 499258 197464 499494
rect 197144 492494 197464 499258
rect 197144 492258 197186 492494
rect 197422 492258 197464 492494
rect 197144 485494 197464 492258
rect 197144 485258 197186 485494
rect 197422 485258 197464 485494
rect 197144 478494 197464 485258
rect 197144 478258 197186 478494
rect 197422 478258 197464 478494
rect 197144 471494 197464 478258
rect 197144 471258 197186 471494
rect 197422 471258 197464 471494
rect 197144 464494 197464 471258
rect 197144 464258 197186 464494
rect 197422 464258 197464 464494
rect 197144 457494 197464 464258
rect 197144 457258 197186 457494
rect 197422 457258 197464 457494
rect 197144 450494 197464 457258
rect 197144 450258 197186 450494
rect 197422 450258 197464 450494
rect 197144 443494 197464 450258
rect 197144 443258 197186 443494
rect 197422 443258 197464 443494
rect 197144 436494 197464 443258
rect 197144 436258 197186 436494
rect 197422 436258 197464 436494
rect 197144 429494 197464 436258
rect 197144 429258 197186 429494
rect 197422 429258 197464 429494
rect 197144 422494 197464 429258
rect 197144 422258 197186 422494
rect 197422 422258 197464 422494
rect 197144 415494 197464 422258
rect 197144 415258 197186 415494
rect 197422 415258 197464 415494
rect 197144 408494 197464 415258
rect 197144 408258 197186 408494
rect 197422 408258 197464 408494
rect 197144 401494 197464 408258
rect 197144 401258 197186 401494
rect 197422 401258 197464 401494
rect 197144 394494 197464 401258
rect 197144 394258 197186 394494
rect 197422 394258 197464 394494
rect 197144 387494 197464 394258
rect 197144 387258 197186 387494
rect 197422 387258 197464 387494
rect 197144 380494 197464 387258
rect 197144 380258 197186 380494
rect 197422 380258 197464 380494
rect 197144 373494 197464 380258
rect 197144 373258 197186 373494
rect 197422 373258 197464 373494
rect 197144 366494 197464 373258
rect 197144 366258 197186 366494
rect 197422 366258 197464 366494
rect 197144 359494 197464 366258
rect 197144 359258 197186 359494
rect 197422 359258 197464 359494
rect 197144 352494 197464 359258
rect 197144 352258 197186 352494
rect 197422 352258 197464 352494
rect 197144 345494 197464 352258
rect 197144 345258 197186 345494
rect 197422 345258 197464 345494
rect 197144 338494 197464 345258
rect 197144 338258 197186 338494
rect 197422 338258 197464 338494
rect 197144 331494 197464 338258
rect 197144 331258 197186 331494
rect 197422 331258 197464 331494
rect 197144 324494 197464 331258
rect 197144 324258 197186 324494
rect 197422 324258 197464 324494
rect 197144 317494 197464 324258
rect 197144 317258 197186 317494
rect 197422 317258 197464 317494
rect 197144 310494 197464 317258
rect 197144 310258 197186 310494
rect 197422 310258 197464 310494
rect 197144 303494 197464 310258
rect 197144 303258 197186 303494
rect 197422 303258 197464 303494
rect 197144 296494 197464 303258
rect 197144 296258 197186 296494
rect 197422 296258 197464 296494
rect 197144 289494 197464 296258
rect 197144 289258 197186 289494
rect 197422 289258 197464 289494
rect 197144 282494 197464 289258
rect 197144 282258 197186 282494
rect 197422 282258 197464 282494
rect 197144 275494 197464 282258
rect 197144 275258 197186 275494
rect 197422 275258 197464 275494
rect 197144 268494 197464 275258
rect 197144 268258 197186 268494
rect 197422 268258 197464 268494
rect 197144 261494 197464 268258
rect 197144 261258 197186 261494
rect 197422 261258 197464 261494
rect 197144 254494 197464 261258
rect 197144 254258 197186 254494
rect 197422 254258 197464 254494
rect 197144 247494 197464 254258
rect 197144 247258 197186 247494
rect 197422 247258 197464 247494
rect 197144 240494 197464 247258
rect 197144 240258 197186 240494
rect 197422 240258 197464 240494
rect 197144 233494 197464 240258
rect 197144 233258 197186 233494
rect 197422 233258 197464 233494
rect 197144 226494 197464 233258
rect 197144 226258 197186 226494
rect 197422 226258 197464 226494
rect 197144 219494 197464 226258
rect 197144 219258 197186 219494
rect 197422 219258 197464 219494
rect 197144 212494 197464 219258
rect 197144 212258 197186 212494
rect 197422 212258 197464 212494
rect 197144 205494 197464 212258
rect 197144 205258 197186 205494
rect 197422 205258 197464 205494
rect 197144 198494 197464 205258
rect 197144 198258 197186 198494
rect 197422 198258 197464 198494
rect 197144 191494 197464 198258
rect 197144 191258 197186 191494
rect 197422 191258 197464 191494
rect 197144 184494 197464 191258
rect 197144 184258 197186 184494
rect 197422 184258 197464 184494
rect 197144 177494 197464 184258
rect 197144 177258 197186 177494
rect 197422 177258 197464 177494
rect 197144 170494 197464 177258
rect 197144 170258 197186 170494
rect 197422 170258 197464 170494
rect 197144 163494 197464 170258
rect 197144 163258 197186 163494
rect 197422 163258 197464 163494
rect 197144 156494 197464 163258
rect 197144 156258 197186 156494
rect 197422 156258 197464 156494
rect 197144 149494 197464 156258
rect 197144 149258 197186 149494
rect 197422 149258 197464 149494
rect 197144 142494 197464 149258
rect 197144 142258 197186 142494
rect 197422 142258 197464 142494
rect 197144 135494 197464 142258
rect 197144 135258 197186 135494
rect 197422 135258 197464 135494
rect 197144 128494 197464 135258
rect 197144 128258 197186 128494
rect 197422 128258 197464 128494
rect 197144 121494 197464 128258
rect 197144 121258 197186 121494
rect 197422 121258 197464 121494
rect 197144 114494 197464 121258
rect 197144 114258 197186 114494
rect 197422 114258 197464 114494
rect 197144 107494 197464 114258
rect 197144 107258 197186 107494
rect 197422 107258 197464 107494
rect 197144 100494 197464 107258
rect 197144 100258 197186 100494
rect 197422 100258 197464 100494
rect 197144 93494 197464 100258
rect 197144 93258 197186 93494
rect 197422 93258 197464 93494
rect 197144 86494 197464 93258
rect 197144 86258 197186 86494
rect 197422 86258 197464 86494
rect 197144 79494 197464 86258
rect 197144 79258 197186 79494
rect 197422 79258 197464 79494
rect 197144 72494 197464 79258
rect 197144 72258 197186 72494
rect 197422 72258 197464 72494
rect 197144 65494 197464 72258
rect 197144 65258 197186 65494
rect 197422 65258 197464 65494
rect 197144 58494 197464 65258
rect 197144 58258 197186 58494
rect 197422 58258 197464 58494
rect 197144 51494 197464 58258
rect 197144 51258 197186 51494
rect 197422 51258 197464 51494
rect 197144 44494 197464 51258
rect 197144 44258 197186 44494
rect 197422 44258 197464 44494
rect 197144 37494 197464 44258
rect 197144 37258 197186 37494
rect 197422 37258 197464 37494
rect 197144 30494 197464 37258
rect 197144 30258 197186 30494
rect 197422 30258 197464 30494
rect 197144 23494 197464 30258
rect 197144 23258 197186 23494
rect 197422 23258 197464 23494
rect 197144 16494 197464 23258
rect 197144 16258 197186 16494
rect 197422 16258 197464 16494
rect 197144 9494 197464 16258
rect 197144 9258 197186 9494
rect 197422 9258 197464 9494
rect 197144 2494 197464 9258
rect 197144 2258 197186 2494
rect 197422 2258 197464 2494
rect 197144 -746 197464 2258
rect 197144 -982 197186 -746
rect 197422 -982 197464 -746
rect 197144 -1066 197464 -982
rect 197144 -1302 197186 -1066
rect 197422 -1302 197464 -1066
rect 197144 -2294 197464 -1302
rect 198876 706198 199196 706230
rect 198876 705962 198918 706198
rect 199154 705962 199196 706198
rect 198876 705878 199196 705962
rect 198876 705642 198918 705878
rect 199154 705642 199196 705878
rect 198876 696561 199196 705642
rect 198876 696325 198918 696561
rect 199154 696325 199196 696561
rect 198876 689561 199196 696325
rect 198876 689325 198918 689561
rect 199154 689325 199196 689561
rect 198876 682561 199196 689325
rect 198876 682325 198918 682561
rect 199154 682325 199196 682561
rect 198876 675561 199196 682325
rect 198876 675325 198918 675561
rect 199154 675325 199196 675561
rect 198876 668561 199196 675325
rect 198876 668325 198918 668561
rect 199154 668325 199196 668561
rect 198876 661561 199196 668325
rect 198876 661325 198918 661561
rect 199154 661325 199196 661561
rect 198876 654561 199196 661325
rect 198876 654325 198918 654561
rect 199154 654325 199196 654561
rect 198876 647561 199196 654325
rect 198876 647325 198918 647561
rect 199154 647325 199196 647561
rect 198876 640561 199196 647325
rect 198876 640325 198918 640561
rect 199154 640325 199196 640561
rect 198876 633561 199196 640325
rect 198876 633325 198918 633561
rect 199154 633325 199196 633561
rect 198876 626561 199196 633325
rect 198876 626325 198918 626561
rect 199154 626325 199196 626561
rect 198876 619561 199196 626325
rect 198876 619325 198918 619561
rect 199154 619325 199196 619561
rect 198876 612561 199196 619325
rect 198876 612325 198918 612561
rect 199154 612325 199196 612561
rect 198876 605561 199196 612325
rect 198876 605325 198918 605561
rect 199154 605325 199196 605561
rect 198876 598561 199196 605325
rect 198876 598325 198918 598561
rect 199154 598325 199196 598561
rect 198876 591561 199196 598325
rect 198876 591325 198918 591561
rect 199154 591325 199196 591561
rect 198876 584561 199196 591325
rect 198876 584325 198918 584561
rect 199154 584325 199196 584561
rect 198876 577561 199196 584325
rect 198876 577325 198918 577561
rect 199154 577325 199196 577561
rect 198876 570561 199196 577325
rect 198876 570325 198918 570561
rect 199154 570325 199196 570561
rect 198876 563561 199196 570325
rect 198876 563325 198918 563561
rect 199154 563325 199196 563561
rect 198876 556561 199196 563325
rect 198876 556325 198918 556561
rect 199154 556325 199196 556561
rect 198876 549561 199196 556325
rect 198876 549325 198918 549561
rect 199154 549325 199196 549561
rect 198876 542561 199196 549325
rect 198876 542325 198918 542561
rect 199154 542325 199196 542561
rect 198876 535561 199196 542325
rect 198876 535325 198918 535561
rect 199154 535325 199196 535561
rect 198876 528561 199196 535325
rect 198876 528325 198918 528561
rect 199154 528325 199196 528561
rect 198876 521561 199196 528325
rect 198876 521325 198918 521561
rect 199154 521325 199196 521561
rect 198876 514561 199196 521325
rect 198876 514325 198918 514561
rect 199154 514325 199196 514561
rect 198876 507561 199196 514325
rect 198876 507325 198918 507561
rect 199154 507325 199196 507561
rect 198876 500561 199196 507325
rect 198876 500325 198918 500561
rect 199154 500325 199196 500561
rect 198876 493561 199196 500325
rect 198876 493325 198918 493561
rect 199154 493325 199196 493561
rect 198876 486561 199196 493325
rect 198876 486325 198918 486561
rect 199154 486325 199196 486561
rect 198876 479561 199196 486325
rect 198876 479325 198918 479561
rect 199154 479325 199196 479561
rect 198876 472561 199196 479325
rect 198876 472325 198918 472561
rect 199154 472325 199196 472561
rect 198876 465561 199196 472325
rect 198876 465325 198918 465561
rect 199154 465325 199196 465561
rect 198876 458561 199196 465325
rect 198876 458325 198918 458561
rect 199154 458325 199196 458561
rect 198876 451561 199196 458325
rect 198876 451325 198918 451561
rect 199154 451325 199196 451561
rect 198876 444561 199196 451325
rect 198876 444325 198918 444561
rect 199154 444325 199196 444561
rect 198876 437561 199196 444325
rect 198876 437325 198918 437561
rect 199154 437325 199196 437561
rect 198876 430561 199196 437325
rect 198876 430325 198918 430561
rect 199154 430325 199196 430561
rect 198876 423561 199196 430325
rect 198876 423325 198918 423561
rect 199154 423325 199196 423561
rect 198876 416561 199196 423325
rect 198876 416325 198918 416561
rect 199154 416325 199196 416561
rect 198876 409561 199196 416325
rect 198876 409325 198918 409561
rect 199154 409325 199196 409561
rect 198876 402561 199196 409325
rect 198876 402325 198918 402561
rect 199154 402325 199196 402561
rect 198876 395561 199196 402325
rect 198876 395325 198918 395561
rect 199154 395325 199196 395561
rect 198876 388561 199196 395325
rect 198876 388325 198918 388561
rect 199154 388325 199196 388561
rect 198876 381561 199196 388325
rect 198876 381325 198918 381561
rect 199154 381325 199196 381561
rect 198876 374561 199196 381325
rect 198876 374325 198918 374561
rect 199154 374325 199196 374561
rect 198876 367561 199196 374325
rect 198876 367325 198918 367561
rect 199154 367325 199196 367561
rect 198876 360561 199196 367325
rect 198876 360325 198918 360561
rect 199154 360325 199196 360561
rect 198876 353561 199196 360325
rect 198876 353325 198918 353561
rect 199154 353325 199196 353561
rect 198876 346561 199196 353325
rect 198876 346325 198918 346561
rect 199154 346325 199196 346561
rect 198876 339561 199196 346325
rect 198876 339325 198918 339561
rect 199154 339325 199196 339561
rect 198876 332561 199196 339325
rect 198876 332325 198918 332561
rect 199154 332325 199196 332561
rect 198876 325561 199196 332325
rect 198876 325325 198918 325561
rect 199154 325325 199196 325561
rect 198876 318561 199196 325325
rect 198876 318325 198918 318561
rect 199154 318325 199196 318561
rect 198876 311561 199196 318325
rect 198876 311325 198918 311561
rect 199154 311325 199196 311561
rect 198876 304561 199196 311325
rect 198876 304325 198918 304561
rect 199154 304325 199196 304561
rect 198876 297561 199196 304325
rect 198876 297325 198918 297561
rect 199154 297325 199196 297561
rect 198876 290561 199196 297325
rect 198876 290325 198918 290561
rect 199154 290325 199196 290561
rect 198876 283561 199196 290325
rect 198876 283325 198918 283561
rect 199154 283325 199196 283561
rect 198876 276561 199196 283325
rect 198876 276325 198918 276561
rect 199154 276325 199196 276561
rect 198876 269561 199196 276325
rect 198876 269325 198918 269561
rect 199154 269325 199196 269561
rect 198876 262561 199196 269325
rect 198876 262325 198918 262561
rect 199154 262325 199196 262561
rect 198876 255561 199196 262325
rect 198876 255325 198918 255561
rect 199154 255325 199196 255561
rect 198876 248561 199196 255325
rect 198876 248325 198918 248561
rect 199154 248325 199196 248561
rect 198876 241561 199196 248325
rect 198876 241325 198918 241561
rect 199154 241325 199196 241561
rect 198876 234561 199196 241325
rect 198876 234325 198918 234561
rect 199154 234325 199196 234561
rect 198876 227561 199196 234325
rect 198876 227325 198918 227561
rect 199154 227325 199196 227561
rect 198876 220561 199196 227325
rect 198876 220325 198918 220561
rect 199154 220325 199196 220561
rect 198876 213561 199196 220325
rect 198876 213325 198918 213561
rect 199154 213325 199196 213561
rect 198876 206561 199196 213325
rect 198876 206325 198918 206561
rect 199154 206325 199196 206561
rect 198876 199561 199196 206325
rect 198876 199325 198918 199561
rect 199154 199325 199196 199561
rect 198876 192561 199196 199325
rect 198876 192325 198918 192561
rect 199154 192325 199196 192561
rect 198876 185561 199196 192325
rect 198876 185325 198918 185561
rect 199154 185325 199196 185561
rect 198876 178561 199196 185325
rect 198876 178325 198918 178561
rect 199154 178325 199196 178561
rect 198876 171561 199196 178325
rect 198876 171325 198918 171561
rect 199154 171325 199196 171561
rect 198876 164561 199196 171325
rect 198876 164325 198918 164561
rect 199154 164325 199196 164561
rect 198876 157561 199196 164325
rect 198876 157325 198918 157561
rect 199154 157325 199196 157561
rect 198876 150561 199196 157325
rect 198876 150325 198918 150561
rect 199154 150325 199196 150561
rect 198876 143561 199196 150325
rect 198876 143325 198918 143561
rect 199154 143325 199196 143561
rect 198876 136561 199196 143325
rect 198876 136325 198918 136561
rect 199154 136325 199196 136561
rect 198876 129561 199196 136325
rect 198876 129325 198918 129561
rect 199154 129325 199196 129561
rect 198876 122561 199196 129325
rect 198876 122325 198918 122561
rect 199154 122325 199196 122561
rect 198876 115561 199196 122325
rect 198876 115325 198918 115561
rect 199154 115325 199196 115561
rect 198876 108561 199196 115325
rect 198876 108325 198918 108561
rect 199154 108325 199196 108561
rect 198876 101561 199196 108325
rect 198876 101325 198918 101561
rect 199154 101325 199196 101561
rect 198876 94561 199196 101325
rect 198876 94325 198918 94561
rect 199154 94325 199196 94561
rect 198876 87561 199196 94325
rect 198876 87325 198918 87561
rect 199154 87325 199196 87561
rect 198876 80561 199196 87325
rect 198876 80325 198918 80561
rect 199154 80325 199196 80561
rect 198876 73561 199196 80325
rect 198876 73325 198918 73561
rect 199154 73325 199196 73561
rect 198876 66561 199196 73325
rect 198876 66325 198918 66561
rect 199154 66325 199196 66561
rect 198876 59561 199196 66325
rect 198876 59325 198918 59561
rect 199154 59325 199196 59561
rect 198876 52561 199196 59325
rect 198876 52325 198918 52561
rect 199154 52325 199196 52561
rect 198876 45561 199196 52325
rect 198876 45325 198918 45561
rect 199154 45325 199196 45561
rect 198876 38561 199196 45325
rect 198876 38325 198918 38561
rect 199154 38325 199196 38561
rect 198876 31561 199196 38325
rect 198876 31325 198918 31561
rect 199154 31325 199196 31561
rect 198876 24561 199196 31325
rect 198876 24325 198918 24561
rect 199154 24325 199196 24561
rect 198876 17561 199196 24325
rect 198876 17325 198918 17561
rect 199154 17325 199196 17561
rect 198876 10561 199196 17325
rect 198876 10325 198918 10561
rect 199154 10325 199196 10561
rect 198876 3561 199196 10325
rect 198876 3325 198918 3561
rect 199154 3325 199196 3561
rect 198876 -1706 199196 3325
rect 198876 -1942 198918 -1706
rect 199154 -1942 199196 -1706
rect 198876 -2026 199196 -1942
rect 198876 -2262 198918 -2026
rect 199154 -2262 199196 -2026
rect 198876 -2294 199196 -2262
rect 204144 705238 204464 706230
rect 204144 705002 204186 705238
rect 204422 705002 204464 705238
rect 204144 704918 204464 705002
rect 204144 704682 204186 704918
rect 204422 704682 204464 704918
rect 204144 695494 204464 704682
rect 204144 695258 204186 695494
rect 204422 695258 204464 695494
rect 204144 688494 204464 695258
rect 204144 688258 204186 688494
rect 204422 688258 204464 688494
rect 204144 681494 204464 688258
rect 204144 681258 204186 681494
rect 204422 681258 204464 681494
rect 204144 674494 204464 681258
rect 204144 674258 204186 674494
rect 204422 674258 204464 674494
rect 204144 667494 204464 674258
rect 204144 667258 204186 667494
rect 204422 667258 204464 667494
rect 204144 660494 204464 667258
rect 204144 660258 204186 660494
rect 204422 660258 204464 660494
rect 204144 653494 204464 660258
rect 204144 653258 204186 653494
rect 204422 653258 204464 653494
rect 204144 646494 204464 653258
rect 204144 646258 204186 646494
rect 204422 646258 204464 646494
rect 204144 639494 204464 646258
rect 204144 639258 204186 639494
rect 204422 639258 204464 639494
rect 204144 632494 204464 639258
rect 204144 632258 204186 632494
rect 204422 632258 204464 632494
rect 204144 625494 204464 632258
rect 204144 625258 204186 625494
rect 204422 625258 204464 625494
rect 204144 618494 204464 625258
rect 204144 618258 204186 618494
rect 204422 618258 204464 618494
rect 204144 611494 204464 618258
rect 204144 611258 204186 611494
rect 204422 611258 204464 611494
rect 204144 604494 204464 611258
rect 204144 604258 204186 604494
rect 204422 604258 204464 604494
rect 204144 597494 204464 604258
rect 204144 597258 204186 597494
rect 204422 597258 204464 597494
rect 204144 590494 204464 597258
rect 204144 590258 204186 590494
rect 204422 590258 204464 590494
rect 204144 583494 204464 590258
rect 204144 583258 204186 583494
rect 204422 583258 204464 583494
rect 204144 576494 204464 583258
rect 204144 576258 204186 576494
rect 204422 576258 204464 576494
rect 204144 569494 204464 576258
rect 204144 569258 204186 569494
rect 204422 569258 204464 569494
rect 204144 562494 204464 569258
rect 204144 562258 204186 562494
rect 204422 562258 204464 562494
rect 204144 555494 204464 562258
rect 204144 555258 204186 555494
rect 204422 555258 204464 555494
rect 204144 548494 204464 555258
rect 204144 548258 204186 548494
rect 204422 548258 204464 548494
rect 204144 541494 204464 548258
rect 204144 541258 204186 541494
rect 204422 541258 204464 541494
rect 204144 534494 204464 541258
rect 204144 534258 204186 534494
rect 204422 534258 204464 534494
rect 204144 527494 204464 534258
rect 204144 527258 204186 527494
rect 204422 527258 204464 527494
rect 204144 520494 204464 527258
rect 204144 520258 204186 520494
rect 204422 520258 204464 520494
rect 204144 513494 204464 520258
rect 204144 513258 204186 513494
rect 204422 513258 204464 513494
rect 204144 506494 204464 513258
rect 204144 506258 204186 506494
rect 204422 506258 204464 506494
rect 204144 499494 204464 506258
rect 204144 499258 204186 499494
rect 204422 499258 204464 499494
rect 204144 492494 204464 499258
rect 204144 492258 204186 492494
rect 204422 492258 204464 492494
rect 204144 485494 204464 492258
rect 204144 485258 204186 485494
rect 204422 485258 204464 485494
rect 204144 478494 204464 485258
rect 204144 478258 204186 478494
rect 204422 478258 204464 478494
rect 204144 471494 204464 478258
rect 204144 471258 204186 471494
rect 204422 471258 204464 471494
rect 204144 464494 204464 471258
rect 204144 464258 204186 464494
rect 204422 464258 204464 464494
rect 204144 457494 204464 464258
rect 204144 457258 204186 457494
rect 204422 457258 204464 457494
rect 204144 450494 204464 457258
rect 204144 450258 204186 450494
rect 204422 450258 204464 450494
rect 204144 443494 204464 450258
rect 204144 443258 204186 443494
rect 204422 443258 204464 443494
rect 204144 436494 204464 443258
rect 204144 436258 204186 436494
rect 204422 436258 204464 436494
rect 204144 429494 204464 436258
rect 204144 429258 204186 429494
rect 204422 429258 204464 429494
rect 204144 422494 204464 429258
rect 204144 422258 204186 422494
rect 204422 422258 204464 422494
rect 204144 415494 204464 422258
rect 204144 415258 204186 415494
rect 204422 415258 204464 415494
rect 204144 408494 204464 415258
rect 204144 408258 204186 408494
rect 204422 408258 204464 408494
rect 204144 401494 204464 408258
rect 204144 401258 204186 401494
rect 204422 401258 204464 401494
rect 204144 394494 204464 401258
rect 204144 394258 204186 394494
rect 204422 394258 204464 394494
rect 204144 387494 204464 394258
rect 204144 387258 204186 387494
rect 204422 387258 204464 387494
rect 204144 380494 204464 387258
rect 204144 380258 204186 380494
rect 204422 380258 204464 380494
rect 204144 373494 204464 380258
rect 204144 373258 204186 373494
rect 204422 373258 204464 373494
rect 204144 366494 204464 373258
rect 204144 366258 204186 366494
rect 204422 366258 204464 366494
rect 204144 359494 204464 366258
rect 204144 359258 204186 359494
rect 204422 359258 204464 359494
rect 204144 352494 204464 359258
rect 204144 352258 204186 352494
rect 204422 352258 204464 352494
rect 204144 345494 204464 352258
rect 204144 345258 204186 345494
rect 204422 345258 204464 345494
rect 204144 338494 204464 345258
rect 204144 338258 204186 338494
rect 204422 338258 204464 338494
rect 204144 331494 204464 338258
rect 204144 331258 204186 331494
rect 204422 331258 204464 331494
rect 204144 324494 204464 331258
rect 204144 324258 204186 324494
rect 204422 324258 204464 324494
rect 204144 317494 204464 324258
rect 204144 317258 204186 317494
rect 204422 317258 204464 317494
rect 204144 310494 204464 317258
rect 204144 310258 204186 310494
rect 204422 310258 204464 310494
rect 204144 303494 204464 310258
rect 204144 303258 204186 303494
rect 204422 303258 204464 303494
rect 204144 296494 204464 303258
rect 204144 296258 204186 296494
rect 204422 296258 204464 296494
rect 204144 289494 204464 296258
rect 204144 289258 204186 289494
rect 204422 289258 204464 289494
rect 204144 282494 204464 289258
rect 204144 282258 204186 282494
rect 204422 282258 204464 282494
rect 204144 275494 204464 282258
rect 204144 275258 204186 275494
rect 204422 275258 204464 275494
rect 204144 268494 204464 275258
rect 204144 268258 204186 268494
rect 204422 268258 204464 268494
rect 204144 261494 204464 268258
rect 204144 261258 204186 261494
rect 204422 261258 204464 261494
rect 204144 254494 204464 261258
rect 204144 254258 204186 254494
rect 204422 254258 204464 254494
rect 204144 247494 204464 254258
rect 204144 247258 204186 247494
rect 204422 247258 204464 247494
rect 204144 240494 204464 247258
rect 204144 240258 204186 240494
rect 204422 240258 204464 240494
rect 204144 233494 204464 240258
rect 204144 233258 204186 233494
rect 204422 233258 204464 233494
rect 204144 226494 204464 233258
rect 204144 226258 204186 226494
rect 204422 226258 204464 226494
rect 204144 219494 204464 226258
rect 204144 219258 204186 219494
rect 204422 219258 204464 219494
rect 204144 212494 204464 219258
rect 204144 212258 204186 212494
rect 204422 212258 204464 212494
rect 204144 205494 204464 212258
rect 204144 205258 204186 205494
rect 204422 205258 204464 205494
rect 204144 198494 204464 205258
rect 204144 198258 204186 198494
rect 204422 198258 204464 198494
rect 204144 191494 204464 198258
rect 204144 191258 204186 191494
rect 204422 191258 204464 191494
rect 204144 184494 204464 191258
rect 204144 184258 204186 184494
rect 204422 184258 204464 184494
rect 204144 177494 204464 184258
rect 204144 177258 204186 177494
rect 204422 177258 204464 177494
rect 204144 170494 204464 177258
rect 204144 170258 204186 170494
rect 204422 170258 204464 170494
rect 204144 163494 204464 170258
rect 204144 163258 204186 163494
rect 204422 163258 204464 163494
rect 204144 156494 204464 163258
rect 204144 156258 204186 156494
rect 204422 156258 204464 156494
rect 204144 149494 204464 156258
rect 204144 149258 204186 149494
rect 204422 149258 204464 149494
rect 204144 142494 204464 149258
rect 204144 142258 204186 142494
rect 204422 142258 204464 142494
rect 204144 135494 204464 142258
rect 204144 135258 204186 135494
rect 204422 135258 204464 135494
rect 204144 128494 204464 135258
rect 204144 128258 204186 128494
rect 204422 128258 204464 128494
rect 204144 121494 204464 128258
rect 204144 121258 204186 121494
rect 204422 121258 204464 121494
rect 204144 114494 204464 121258
rect 204144 114258 204186 114494
rect 204422 114258 204464 114494
rect 204144 107494 204464 114258
rect 204144 107258 204186 107494
rect 204422 107258 204464 107494
rect 204144 100494 204464 107258
rect 204144 100258 204186 100494
rect 204422 100258 204464 100494
rect 204144 93494 204464 100258
rect 204144 93258 204186 93494
rect 204422 93258 204464 93494
rect 204144 86494 204464 93258
rect 204144 86258 204186 86494
rect 204422 86258 204464 86494
rect 204144 79494 204464 86258
rect 204144 79258 204186 79494
rect 204422 79258 204464 79494
rect 204144 72494 204464 79258
rect 204144 72258 204186 72494
rect 204422 72258 204464 72494
rect 204144 65494 204464 72258
rect 204144 65258 204186 65494
rect 204422 65258 204464 65494
rect 204144 58494 204464 65258
rect 204144 58258 204186 58494
rect 204422 58258 204464 58494
rect 204144 51494 204464 58258
rect 204144 51258 204186 51494
rect 204422 51258 204464 51494
rect 204144 44494 204464 51258
rect 204144 44258 204186 44494
rect 204422 44258 204464 44494
rect 204144 37494 204464 44258
rect 204144 37258 204186 37494
rect 204422 37258 204464 37494
rect 204144 30494 204464 37258
rect 204144 30258 204186 30494
rect 204422 30258 204464 30494
rect 204144 23494 204464 30258
rect 204144 23258 204186 23494
rect 204422 23258 204464 23494
rect 204144 16494 204464 23258
rect 204144 16258 204186 16494
rect 204422 16258 204464 16494
rect 204144 9494 204464 16258
rect 204144 9258 204186 9494
rect 204422 9258 204464 9494
rect 204144 2494 204464 9258
rect 204144 2258 204186 2494
rect 204422 2258 204464 2494
rect 204144 -746 204464 2258
rect 204144 -982 204186 -746
rect 204422 -982 204464 -746
rect 204144 -1066 204464 -982
rect 204144 -1302 204186 -1066
rect 204422 -1302 204464 -1066
rect 204144 -2294 204464 -1302
rect 205876 706198 206196 706230
rect 205876 705962 205918 706198
rect 206154 705962 206196 706198
rect 205876 705878 206196 705962
rect 205876 705642 205918 705878
rect 206154 705642 206196 705878
rect 205876 696561 206196 705642
rect 205876 696325 205918 696561
rect 206154 696325 206196 696561
rect 205876 689561 206196 696325
rect 205876 689325 205918 689561
rect 206154 689325 206196 689561
rect 205876 682561 206196 689325
rect 205876 682325 205918 682561
rect 206154 682325 206196 682561
rect 205876 675561 206196 682325
rect 205876 675325 205918 675561
rect 206154 675325 206196 675561
rect 205876 668561 206196 675325
rect 205876 668325 205918 668561
rect 206154 668325 206196 668561
rect 205876 661561 206196 668325
rect 205876 661325 205918 661561
rect 206154 661325 206196 661561
rect 205876 654561 206196 661325
rect 205876 654325 205918 654561
rect 206154 654325 206196 654561
rect 205876 647561 206196 654325
rect 205876 647325 205918 647561
rect 206154 647325 206196 647561
rect 205876 640561 206196 647325
rect 205876 640325 205918 640561
rect 206154 640325 206196 640561
rect 205876 633561 206196 640325
rect 205876 633325 205918 633561
rect 206154 633325 206196 633561
rect 205876 626561 206196 633325
rect 205876 626325 205918 626561
rect 206154 626325 206196 626561
rect 205876 619561 206196 626325
rect 205876 619325 205918 619561
rect 206154 619325 206196 619561
rect 205876 612561 206196 619325
rect 205876 612325 205918 612561
rect 206154 612325 206196 612561
rect 205876 605561 206196 612325
rect 205876 605325 205918 605561
rect 206154 605325 206196 605561
rect 205876 598561 206196 605325
rect 205876 598325 205918 598561
rect 206154 598325 206196 598561
rect 205876 591561 206196 598325
rect 205876 591325 205918 591561
rect 206154 591325 206196 591561
rect 205876 584561 206196 591325
rect 205876 584325 205918 584561
rect 206154 584325 206196 584561
rect 205876 577561 206196 584325
rect 205876 577325 205918 577561
rect 206154 577325 206196 577561
rect 205876 570561 206196 577325
rect 205876 570325 205918 570561
rect 206154 570325 206196 570561
rect 205876 563561 206196 570325
rect 205876 563325 205918 563561
rect 206154 563325 206196 563561
rect 205876 556561 206196 563325
rect 205876 556325 205918 556561
rect 206154 556325 206196 556561
rect 205876 549561 206196 556325
rect 205876 549325 205918 549561
rect 206154 549325 206196 549561
rect 205876 542561 206196 549325
rect 205876 542325 205918 542561
rect 206154 542325 206196 542561
rect 205876 535561 206196 542325
rect 205876 535325 205918 535561
rect 206154 535325 206196 535561
rect 205876 528561 206196 535325
rect 205876 528325 205918 528561
rect 206154 528325 206196 528561
rect 205876 521561 206196 528325
rect 205876 521325 205918 521561
rect 206154 521325 206196 521561
rect 205876 514561 206196 521325
rect 205876 514325 205918 514561
rect 206154 514325 206196 514561
rect 205876 507561 206196 514325
rect 205876 507325 205918 507561
rect 206154 507325 206196 507561
rect 205876 500561 206196 507325
rect 205876 500325 205918 500561
rect 206154 500325 206196 500561
rect 205876 493561 206196 500325
rect 205876 493325 205918 493561
rect 206154 493325 206196 493561
rect 205876 486561 206196 493325
rect 205876 486325 205918 486561
rect 206154 486325 206196 486561
rect 205876 479561 206196 486325
rect 205876 479325 205918 479561
rect 206154 479325 206196 479561
rect 205876 472561 206196 479325
rect 205876 472325 205918 472561
rect 206154 472325 206196 472561
rect 205876 465561 206196 472325
rect 205876 465325 205918 465561
rect 206154 465325 206196 465561
rect 205876 458561 206196 465325
rect 205876 458325 205918 458561
rect 206154 458325 206196 458561
rect 205876 451561 206196 458325
rect 205876 451325 205918 451561
rect 206154 451325 206196 451561
rect 205876 444561 206196 451325
rect 205876 444325 205918 444561
rect 206154 444325 206196 444561
rect 205876 437561 206196 444325
rect 205876 437325 205918 437561
rect 206154 437325 206196 437561
rect 205876 430561 206196 437325
rect 205876 430325 205918 430561
rect 206154 430325 206196 430561
rect 205876 423561 206196 430325
rect 205876 423325 205918 423561
rect 206154 423325 206196 423561
rect 205876 416561 206196 423325
rect 205876 416325 205918 416561
rect 206154 416325 206196 416561
rect 205876 409561 206196 416325
rect 205876 409325 205918 409561
rect 206154 409325 206196 409561
rect 205876 402561 206196 409325
rect 205876 402325 205918 402561
rect 206154 402325 206196 402561
rect 205876 395561 206196 402325
rect 205876 395325 205918 395561
rect 206154 395325 206196 395561
rect 205876 388561 206196 395325
rect 205876 388325 205918 388561
rect 206154 388325 206196 388561
rect 205876 381561 206196 388325
rect 205876 381325 205918 381561
rect 206154 381325 206196 381561
rect 205876 374561 206196 381325
rect 205876 374325 205918 374561
rect 206154 374325 206196 374561
rect 205876 367561 206196 374325
rect 205876 367325 205918 367561
rect 206154 367325 206196 367561
rect 205876 360561 206196 367325
rect 205876 360325 205918 360561
rect 206154 360325 206196 360561
rect 205876 353561 206196 360325
rect 205876 353325 205918 353561
rect 206154 353325 206196 353561
rect 205876 346561 206196 353325
rect 205876 346325 205918 346561
rect 206154 346325 206196 346561
rect 205876 339561 206196 346325
rect 205876 339325 205918 339561
rect 206154 339325 206196 339561
rect 205876 332561 206196 339325
rect 205876 332325 205918 332561
rect 206154 332325 206196 332561
rect 205876 325561 206196 332325
rect 205876 325325 205918 325561
rect 206154 325325 206196 325561
rect 205876 318561 206196 325325
rect 205876 318325 205918 318561
rect 206154 318325 206196 318561
rect 205876 311561 206196 318325
rect 205876 311325 205918 311561
rect 206154 311325 206196 311561
rect 205876 304561 206196 311325
rect 205876 304325 205918 304561
rect 206154 304325 206196 304561
rect 205876 297561 206196 304325
rect 205876 297325 205918 297561
rect 206154 297325 206196 297561
rect 205876 290561 206196 297325
rect 205876 290325 205918 290561
rect 206154 290325 206196 290561
rect 205876 283561 206196 290325
rect 205876 283325 205918 283561
rect 206154 283325 206196 283561
rect 205876 276561 206196 283325
rect 205876 276325 205918 276561
rect 206154 276325 206196 276561
rect 205876 269561 206196 276325
rect 205876 269325 205918 269561
rect 206154 269325 206196 269561
rect 205876 262561 206196 269325
rect 205876 262325 205918 262561
rect 206154 262325 206196 262561
rect 205876 255561 206196 262325
rect 205876 255325 205918 255561
rect 206154 255325 206196 255561
rect 205876 248561 206196 255325
rect 205876 248325 205918 248561
rect 206154 248325 206196 248561
rect 205876 241561 206196 248325
rect 205876 241325 205918 241561
rect 206154 241325 206196 241561
rect 205876 234561 206196 241325
rect 205876 234325 205918 234561
rect 206154 234325 206196 234561
rect 205876 227561 206196 234325
rect 205876 227325 205918 227561
rect 206154 227325 206196 227561
rect 205876 220561 206196 227325
rect 205876 220325 205918 220561
rect 206154 220325 206196 220561
rect 205876 213561 206196 220325
rect 205876 213325 205918 213561
rect 206154 213325 206196 213561
rect 205876 206561 206196 213325
rect 205876 206325 205918 206561
rect 206154 206325 206196 206561
rect 205876 199561 206196 206325
rect 205876 199325 205918 199561
rect 206154 199325 206196 199561
rect 205876 192561 206196 199325
rect 205876 192325 205918 192561
rect 206154 192325 206196 192561
rect 205876 185561 206196 192325
rect 205876 185325 205918 185561
rect 206154 185325 206196 185561
rect 205876 178561 206196 185325
rect 205876 178325 205918 178561
rect 206154 178325 206196 178561
rect 205876 171561 206196 178325
rect 205876 171325 205918 171561
rect 206154 171325 206196 171561
rect 205876 164561 206196 171325
rect 205876 164325 205918 164561
rect 206154 164325 206196 164561
rect 205876 157561 206196 164325
rect 205876 157325 205918 157561
rect 206154 157325 206196 157561
rect 205876 150561 206196 157325
rect 205876 150325 205918 150561
rect 206154 150325 206196 150561
rect 205876 143561 206196 150325
rect 205876 143325 205918 143561
rect 206154 143325 206196 143561
rect 205876 136561 206196 143325
rect 205876 136325 205918 136561
rect 206154 136325 206196 136561
rect 205876 129561 206196 136325
rect 205876 129325 205918 129561
rect 206154 129325 206196 129561
rect 205876 122561 206196 129325
rect 205876 122325 205918 122561
rect 206154 122325 206196 122561
rect 205876 115561 206196 122325
rect 205876 115325 205918 115561
rect 206154 115325 206196 115561
rect 205876 108561 206196 115325
rect 205876 108325 205918 108561
rect 206154 108325 206196 108561
rect 205876 101561 206196 108325
rect 205876 101325 205918 101561
rect 206154 101325 206196 101561
rect 205876 94561 206196 101325
rect 205876 94325 205918 94561
rect 206154 94325 206196 94561
rect 205876 87561 206196 94325
rect 205876 87325 205918 87561
rect 206154 87325 206196 87561
rect 205876 80561 206196 87325
rect 205876 80325 205918 80561
rect 206154 80325 206196 80561
rect 205876 73561 206196 80325
rect 205876 73325 205918 73561
rect 206154 73325 206196 73561
rect 205876 66561 206196 73325
rect 205876 66325 205918 66561
rect 206154 66325 206196 66561
rect 205876 59561 206196 66325
rect 205876 59325 205918 59561
rect 206154 59325 206196 59561
rect 205876 52561 206196 59325
rect 205876 52325 205918 52561
rect 206154 52325 206196 52561
rect 205876 45561 206196 52325
rect 205876 45325 205918 45561
rect 206154 45325 206196 45561
rect 205876 38561 206196 45325
rect 205876 38325 205918 38561
rect 206154 38325 206196 38561
rect 205876 31561 206196 38325
rect 205876 31325 205918 31561
rect 206154 31325 206196 31561
rect 205876 24561 206196 31325
rect 205876 24325 205918 24561
rect 206154 24325 206196 24561
rect 205876 17561 206196 24325
rect 205876 17325 205918 17561
rect 206154 17325 206196 17561
rect 205876 10561 206196 17325
rect 205876 10325 205918 10561
rect 206154 10325 206196 10561
rect 205876 3561 206196 10325
rect 205876 3325 205918 3561
rect 206154 3325 206196 3561
rect 205876 -1706 206196 3325
rect 205876 -1942 205918 -1706
rect 206154 -1942 206196 -1706
rect 205876 -2026 206196 -1942
rect 205876 -2262 205918 -2026
rect 206154 -2262 206196 -2026
rect 205876 -2294 206196 -2262
rect 211144 705238 211464 706230
rect 211144 705002 211186 705238
rect 211422 705002 211464 705238
rect 211144 704918 211464 705002
rect 211144 704682 211186 704918
rect 211422 704682 211464 704918
rect 211144 695494 211464 704682
rect 211144 695258 211186 695494
rect 211422 695258 211464 695494
rect 211144 688494 211464 695258
rect 211144 688258 211186 688494
rect 211422 688258 211464 688494
rect 211144 681494 211464 688258
rect 211144 681258 211186 681494
rect 211422 681258 211464 681494
rect 211144 674494 211464 681258
rect 211144 674258 211186 674494
rect 211422 674258 211464 674494
rect 211144 667494 211464 674258
rect 211144 667258 211186 667494
rect 211422 667258 211464 667494
rect 211144 660494 211464 667258
rect 211144 660258 211186 660494
rect 211422 660258 211464 660494
rect 211144 653494 211464 660258
rect 211144 653258 211186 653494
rect 211422 653258 211464 653494
rect 211144 646494 211464 653258
rect 211144 646258 211186 646494
rect 211422 646258 211464 646494
rect 211144 639494 211464 646258
rect 211144 639258 211186 639494
rect 211422 639258 211464 639494
rect 211144 632494 211464 639258
rect 211144 632258 211186 632494
rect 211422 632258 211464 632494
rect 211144 625494 211464 632258
rect 211144 625258 211186 625494
rect 211422 625258 211464 625494
rect 211144 618494 211464 625258
rect 211144 618258 211186 618494
rect 211422 618258 211464 618494
rect 211144 611494 211464 618258
rect 211144 611258 211186 611494
rect 211422 611258 211464 611494
rect 211144 604494 211464 611258
rect 211144 604258 211186 604494
rect 211422 604258 211464 604494
rect 211144 597494 211464 604258
rect 211144 597258 211186 597494
rect 211422 597258 211464 597494
rect 211144 590494 211464 597258
rect 211144 590258 211186 590494
rect 211422 590258 211464 590494
rect 211144 583494 211464 590258
rect 211144 583258 211186 583494
rect 211422 583258 211464 583494
rect 211144 576494 211464 583258
rect 211144 576258 211186 576494
rect 211422 576258 211464 576494
rect 211144 569494 211464 576258
rect 211144 569258 211186 569494
rect 211422 569258 211464 569494
rect 211144 562494 211464 569258
rect 211144 562258 211186 562494
rect 211422 562258 211464 562494
rect 211144 555494 211464 562258
rect 211144 555258 211186 555494
rect 211422 555258 211464 555494
rect 211144 548494 211464 555258
rect 211144 548258 211186 548494
rect 211422 548258 211464 548494
rect 211144 541494 211464 548258
rect 211144 541258 211186 541494
rect 211422 541258 211464 541494
rect 211144 534494 211464 541258
rect 211144 534258 211186 534494
rect 211422 534258 211464 534494
rect 211144 527494 211464 534258
rect 211144 527258 211186 527494
rect 211422 527258 211464 527494
rect 211144 520494 211464 527258
rect 211144 520258 211186 520494
rect 211422 520258 211464 520494
rect 211144 513494 211464 520258
rect 211144 513258 211186 513494
rect 211422 513258 211464 513494
rect 211144 506494 211464 513258
rect 211144 506258 211186 506494
rect 211422 506258 211464 506494
rect 211144 499494 211464 506258
rect 211144 499258 211186 499494
rect 211422 499258 211464 499494
rect 211144 492494 211464 499258
rect 211144 492258 211186 492494
rect 211422 492258 211464 492494
rect 211144 485494 211464 492258
rect 211144 485258 211186 485494
rect 211422 485258 211464 485494
rect 211144 478494 211464 485258
rect 211144 478258 211186 478494
rect 211422 478258 211464 478494
rect 211144 471494 211464 478258
rect 211144 471258 211186 471494
rect 211422 471258 211464 471494
rect 211144 464494 211464 471258
rect 211144 464258 211186 464494
rect 211422 464258 211464 464494
rect 211144 457494 211464 464258
rect 211144 457258 211186 457494
rect 211422 457258 211464 457494
rect 211144 450494 211464 457258
rect 211144 450258 211186 450494
rect 211422 450258 211464 450494
rect 211144 443494 211464 450258
rect 211144 443258 211186 443494
rect 211422 443258 211464 443494
rect 211144 436494 211464 443258
rect 211144 436258 211186 436494
rect 211422 436258 211464 436494
rect 211144 429494 211464 436258
rect 211144 429258 211186 429494
rect 211422 429258 211464 429494
rect 211144 422494 211464 429258
rect 211144 422258 211186 422494
rect 211422 422258 211464 422494
rect 211144 415494 211464 422258
rect 211144 415258 211186 415494
rect 211422 415258 211464 415494
rect 211144 408494 211464 415258
rect 211144 408258 211186 408494
rect 211422 408258 211464 408494
rect 211144 401494 211464 408258
rect 211144 401258 211186 401494
rect 211422 401258 211464 401494
rect 211144 394494 211464 401258
rect 211144 394258 211186 394494
rect 211422 394258 211464 394494
rect 211144 387494 211464 394258
rect 211144 387258 211186 387494
rect 211422 387258 211464 387494
rect 211144 380494 211464 387258
rect 211144 380258 211186 380494
rect 211422 380258 211464 380494
rect 211144 373494 211464 380258
rect 211144 373258 211186 373494
rect 211422 373258 211464 373494
rect 211144 366494 211464 373258
rect 211144 366258 211186 366494
rect 211422 366258 211464 366494
rect 211144 359494 211464 366258
rect 211144 359258 211186 359494
rect 211422 359258 211464 359494
rect 211144 352494 211464 359258
rect 211144 352258 211186 352494
rect 211422 352258 211464 352494
rect 211144 345494 211464 352258
rect 211144 345258 211186 345494
rect 211422 345258 211464 345494
rect 211144 338494 211464 345258
rect 211144 338258 211186 338494
rect 211422 338258 211464 338494
rect 211144 331494 211464 338258
rect 211144 331258 211186 331494
rect 211422 331258 211464 331494
rect 211144 324494 211464 331258
rect 211144 324258 211186 324494
rect 211422 324258 211464 324494
rect 211144 317494 211464 324258
rect 211144 317258 211186 317494
rect 211422 317258 211464 317494
rect 211144 310494 211464 317258
rect 211144 310258 211186 310494
rect 211422 310258 211464 310494
rect 211144 303494 211464 310258
rect 211144 303258 211186 303494
rect 211422 303258 211464 303494
rect 211144 296494 211464 303258
rect 211144 296258 211186 296494
rect 211422 296258 211464 296494
rect 211144 289494 211464 296258
rect 211144 289258 211186 289494
rect 211422 289258 211464 289494
rect 211144 282494 211464 289258
rect 211144 282258 211186 282494
rect 211422 282258 211464 282494
rect 211144 275494 211464 282258
rect 211144 275258 211186 275494
rect 211422 275258 211464 275494
rect 211144 268494 211464 275258
rect 211144 268258 211186 268494
rect 211422 268258 211464 268494
rect 211144 261494 211464 268258
rect 211144 261258 211186 261494
rect 211422 261258 211464 261494
rect 211144 254494 211464 261258
rect 211144 254258 211186 254494
rect 211422 254258 211464 254494
rect 211144 247494 211464 254258
rect 211144 247258 211186 247494
rect 211422 247258 211464 247494
rect 211144 240494 211464 247258
rect 211144 240258 211186 240494
rect 211422 240258 211464 240494
rect 211144 233494 211464 240258
rect 211144 233258 211186 233494
rect 211422 233258 211464 233494
rect 211144 226494 211464 233258
rect 211144 226258 211186 226494
rect 211422 226258 211464 226494
rect 211144 219494 211464 226258
rect 211144 219258 211186 219494
rect 211422 219258 211464 219494
rect 211144 212494 211464 219258
rect 211144 212258 211186 212494
rect 211422 212258 211464 212494
rect 211144 205494 211464 212258
rect 211144 205258 211186 205494
rect 211422 205258 211464 205494
rect 211144 198494 211464 205258
rect 211144 198258 211186 198494
rect 211422 198258 211464 198494
rect 211144 191494 211464 198258
rect 211144 191258 211186 191494
rect 211422 191258 211464 191494
rect 211144 184494 211464 191258
rect 211144 184258 211186 184494
rect 211422 184258 211464 184494
rect 211144 177494 211464 184258
rect 211144 177258 211186 177494
rect 211422 177258 211464 177494
rect 211144 170494 211464 177258
rect 211144 170258 211186 170494
rect 211422 170258 211464 170494
rect 211144 163494 211464 170258
rect 211144 163258 211186 163494
rect 211422 163258 211464 163494
rect 211144 156494 211464 163258
rect 211144 156258 211186 156494
rect 211422 156258 211464 156494
rect 211144 149494 211464 156258
rect 211144 149258 211186 149494
rect 211422 149258 211464 149494
rect 211144 142494 211464 149258
rect 211144 142258 211186 142494
rect 211422 142258 211464 142494
rect 211144 135494 211464 142258
rect 211144 135258 211186 135494
rect 211422 135258 211464 135494
rect 211144 128494 211464 135258
rect 211144 128258 211186 128494
rect 211422 128258 211464 128494
rect 211144 121494 211464 128258
rect 211144 121258 211186 121494
rect 211422 121258 211464 121494
rect 211144 114494 211464 121258
rect 211144 114258 211186 114494
rect 211422 114258 211464 114494
rect 211144 107494 211464 114258
rect 211144 107258 211186 107494
rect 211422 107258 211464 107494
rect 211144 100494 211464 107258
rect 211144 100258 211186 100494
rect 211422 100258 211464 100494
rect 211144 93494 211464 100258
rect 211144 93258 211186 93494
rect 211422 93258 211464 93494
rect 211144 86494 211464 93258
rect 211144 86258 211186 86494
rect 211422 86258 211464 86494
rect 211144 79494 211464 86258
rect 211144 79258 211186 79494
rect 211422 79258 211464 79494
rect 211144 72494 211464 79258
rect 211144 72258 211186 72494
rect 211422 72258 211464 72494
rect 211144 65494 211464 72258
rect 211144 65258 211186 65494
rect 211422 65258 211464 65494
rect 211144 58494 211464 65258
rect 211144 58258 211186 58494
rect 211422 58258 211464 58494
rect 211144 51494 211464 58258
rect 211144 51258 211186 51494
rect 211422 51258 211464 51494
rect 211144 44494 211464 51258
rect 211144 44258 211186 44494
rect 211422 44258 211464 44494
rect 211144 37494 211464 44258
rect 211144 37258 211186 37494
rect 211422 37258 211464 37494
rect 211144 30494 211464 37258
rect 211144 30258 211186 30494
rect 211422 30258 211464 30494
rect 211144 23494 211464 30258
rect 211144 23258 211186 23494
rect 211422 23258 211464 23494
rect 211144 16494 211464 23258
rect 211144 16258 211186 16494
rect 211422 16258 211464 16494
rect 211144 9494 211464 16258
rect 211144 9258 211186 9494
rect 211422 9258 211464 9494
rect 211144 2494 211464 9258
rect 211144 2258 211186 2494
rect 211422 2258 211464 2494
rect 211144 -746 211464 2258
rect 211144 -982 211186 -746
rect 211422 -982 211464 -746
rect 211144 -1066 211464 -982
rect 211144 -1302 211186 -1066
rect 211422 -1302 211464 -1066
rect 211144 -2294 211464 -1302
rect 212876 706198 213196 706230
rect 212876 705962 212918 706198
rect 213154 705962 213196 706198
rect 212876 705878 213196 705962
rect 212876 705642 212918 705878
rect 213154 705642 213196 705878
rect 212876 696561 213196 705642
rect 212876 696325 212918 696561
rect 213154 696325 213196 696561
rect 212876 689561 213196 696325
rect 212876 689325 212918 689561
rect 213154 689325 213196 689561
rect 212876 682561 213196 689325
rect 212876 682325 212918 682561
rect 213154 682325 213196 682561
rect 212876 675561 213196 682325
rect 212876 675325 212918 675561
rect 213154 675325 213196 675561
rect 212876 668561 213196 675325
rect 212876 668325 212918 668561
rect 213154 668325 213196 668561
rect 212876 661561 213196 668325
rect 212876 661325 212918 661561
rect 213154 661325 213196 661561
rect 212876 654561 213196 661325
rect 212876 654325 212918 654561
rect 213154 654325 213196 654561
rect 212876 647561 213196 654325
rect 212876 647325 212918 647561
rect 213154 647325 213196 647561
rect 212876 640561 213196 647325
rect 212876 640325 212918 640561
rect 213154 640325 213196 640561
rect 212876 633561 213196 640325
rect 212876 633325 212918 633561
rect 213154 633325 213196 633561
rect 212876 626561 213196 633325
rect 212876 626325 212918 626561
rect 213154 626325 213196 626561
rect 212876 619561 213196 626325
rect 212876 619325 212918 619561
rect 213154 619325 213196 619561
rect 212876 612561 213196 619325
rect 212876 612325 212918 612561
rect 213154 612325 213196 612561
rect 212876 605561 213196 612325
rect 212876 605325 212918 605561
rect 213154 605325 213196 605561
rect 212876 598561 213196 605325
rect 212876 598325 212918 598561
rect 213154 598325 213196 598561
rect 212876 591561 213196 598325
rect 212876 591325 212918 591561
rect 213154 591325 213196 591561
rect 212876 584561 213196 591325
rect 212876 584325 212918 584561
rect 213154 584325 213196 584561
rect 212876 577561 213196 584325
rect 212876 577325 212918 577561
rect 213154 577325 213196 577561
rect 212876 570561 213196 577325
rect 212876 570325 212918 570561
rect 213154 570325 213196 570561
rect 212876 563561 213196 570325
rect 212876 563325 212918 563561
rect 213154 563325 213196 563561
rect 212876 556561 213196 563325
rect 212876 556325 212918 556561
rect 213154 556325 213196 556561
rect 212876 549561 213196 556325
rect 212876 549325 212918 549561
rect 213154 549325 213196 549561
rect 212876 542561 213196 549325
rect 212876 542325 212918 542561
rect 213154 542325 213196 542561
rect 212876 535561 213196 542325
rect 212876 535325 212918 535561
rect 213154 535325 213196 535561
rect 212876 528561 213196 535325
rect 212876 528325 212918 528561
rect 213154 528325 213196 528561
rect 212876 521561 213196 528325
rect 212876 521325 212918 521561
rect 213154 521325 213196 521561
rect 212876 514561 213196 521325
rect 212876 514325 212918 514561
rect 213154 514325 213196 514561
rect 212876 507561 213196 514325
rect 212876 507325 212918 507561
rect 213154 507325 213196 507561
rect 212876 500561 213196 507325
rect 212876 500325 212918 500561
rect 213154 500325 213196 500561
rect 212876 493561 213196 500325
rect 212876 493325 212918 493561
rect 213154 493325 213196 493561
rect 212876 486561 213196 493325
rect 212876 486325 212918 486561
rect 213154 486325 213196 486561
rect 212876 479561 213196 486325
rect 212876 479325 212918 479561
rect 213154 479325 213196 479561
rect 212876 472561 213196 479325
rect 212876 472325 212918 472561
rect 213154 472325 213196 472561
rect 212876 465561 213196 472325
rect 212876 465325 212918 465561
rect 213154 465325 213196 465561
rect 212876 458561 213196 465325
rect 212876 458325 212918 458561
rect 213154 458325 213196 458561
rect 212876 451561 213196 458325
rect 212876 451325 212918 451561
rect 213154 451325 213196 451561
rect 212876 444561 213196 451325
rect 212876 444325 212918 444561
rect 213154 444325 213196 444561
rect 212876 437561 213196 444325
rect 212876 437325 212918 437561
rect 213154 437325 213196 437561
rect 212876 430561 213196 437325
rect 212876 430325 212918 430561
rect 213154 430325 213196 430561
rect 212876 423561 213196 430325
rect 212876 423325 212918 423561
rect 213154 423325 213196 423561
rect 212876 416561 213196 423325
rect 212876 416325 212918 416561
rect 213154 416325 213196 416561
rect 212876 409561 213196 416325
rect 212876 409325 212918 409561
rect 213154 409325 213196 409561
rect 212876 402561 213196 409325
rect 212876 402325 212918 402561
rect 213154 402325 213196 402561
rect 212876 395561 213196 402325
rect 212876 395325 212918 395561
rect 213154 395325 213196 395561
rect 212876 388561 213196 395325
rect 212876 388325 212918 388561
rect 213154 388325 213196 388561
rect 212876 381561 213196 388325
rect 212876 381325 212918 381561
rect 213154 381325 213196 381561
rect 212876 374561 213196 381325
rect 212876 374325 212918 374561
rect 213154 374325 213196 374561
rect 212876 367561 213196 374325
rect 212876 367325 212918 367561
rect 213154 367325 213196 367561
rect 212876 360561 213196 367325
rect 212876 360325 212918 360561
rect 213154 360325 213196 360561
rect 212876 353561 213196 360325
rect 212876 353325 212918 353561
rect 213154 353325 213196 353561
rect 212876 346561 213196 353325
rect 212876 346325 212918 346561
rect 213154 346325 213196 346561
rect 212876 339561 213196 346325
rect 212876 339325 212918 339561
rect 213154 339325 213196 339561
rect 212876 332561 213196 339325
rect 212876 332325 212918 332561
rect 213154 332325 213196 332561
rect 212876 325561 213196 332325
rect 212876 325325 212918 325561
rect 213154 325325 213196 325561
rect 212876 318561 213196 325325
rect 212876 318325 212918 318561
rect 213154 318325 213196 318561
rect 212876 311561 213196 318325
rect 212876 311325 212918 311561
rect 213154 311325 213196 311561
rect 212876 304561 213196 311325
rect 212876 304325 212918 304561
rect 213154 304325 213196 304561
rect 212876 297561 213196 304325
rect 212876 297325 212918 297561
rect 213154 297325 213196 297561
rect 212876 290561 213196 297325
rect 212876 290325 212918 290561
rect 213154 290325 213196 290561
rect 212876 283561 213196 290325
rect 212876 283325 212918 283561
rect 213154 283325 213196 283561
rect 212876 276561 213196 283325
rect 212876 276325 212918 276561
rect 213154 276325 213196 276561
rect 212876 269561 213196 276325
rect 212876 269325 212918 269561
rect 213154 269325 213196 269561
rect 212876 262561 213196 269325
rect 212876 262325 212918 262561
rect 213154 262325 213196 262561
rect 212876 255561 213196 262325
rect 212876 255325 212918 255561
rect 213154 255325 213196 255561
rect 212876 248561 213196 255325
rect 212876 248325 212918 248561
rect 213154 248325 213196 248561
rect 212876 241561 213196 248325
rect 212876 241325 212918 241561
rect 213154 241325 213196 241561
rect 212876 234561 213196 241325
rect 212876 234325 212918 234561
rect 213154 234325 213196 234561
rect 212876 227561 213196 234325
rect 212876 227325 212918 227561
rect 213154 227325 213196 227561
rect 212876 220561 213196 227325
rect 212876 220325 212918 220561
rect 213154 220325 213196 220561
rect 212876 213561 213196 220325
rect 212876 213325 212918 213561
rect 213154 213325 213196 213561
rect 212876 206561 213196 213325
rect 212876 206325 212918 206561
rect 213154 206325 213196 206561
rect 212876 199561 213196 206325
rect 212876 199325 212918 199561
rect 213154 199325 213196 199561
rect 212876 192561 213196 199325
rect 212876 192325 212918 192561
rect 213154 192325 213196 192561
rect 212876 185561 213196 192325
rect 212876 185325 212918 185561
rect 213154 185325 213196 185561
rect 212876 178561 213196 185325
rect 212876 178325 212918 178561
rect 213154 178325 213196 178561
rect 212876 171561 213196 178325
rect 212876 171325 212918 171561
rect 213154 171325 213196 171561
rect 212876 164561 213196 171325
rect 212876 164325 212918 164561
rect 213154 164325 213196 164561
rect 212876 157561 213196 164325
rect 212876 157325 212918 157561
rect 213154 157325 213196 157561
rect 212876 150561 213196 157325
rect 212876 150325 212918 150561
rect 213154 150325 213196 150561
rect 212876 143561 213196 150325
rect 212876 143325 212918 143561
rect 213154 143325 213196 143561
rect 212876 136561 213196 143325
rect 212876 136325 212918 136561
rect 213154 136325 213196 136561
rect 212876 129561 213196 136325
rect 212876 129325 212918 129561
rect 213154 129325 213196 129561
rect 212876 122561 213196 129325
rect 212876 122325 212918 122561
rect 213154 122325 213196 122561
rect 212876 115561 213196 122325
rect 212876 115325 212918 115561
rect 213154 115325 213196 115561
rect 212876 108561 213196 115325
rect 212876 108325 212918 108561
rect 213154 108325 213196 108561
rect 212876 101561 213196 108325
rect 212876 101325 212918 101561
rect 213154 101325 213196 101561
rect 212876 94561 213196 101325
rect 212876 94325 212918 94561
rect 213154 94325 213196 94561
rect 212876 87561 213196 94325
rect 212876 87325 212918 87561
rect 213154 87325 213196 87561
rect 212876 80561 213196 87325
rect 212876 80325 212918 80561
rect 213154 80325 213196 80561
rect 212876 73561 213196 80325
rect 212876 73325 212918 73561
rect 213154 73325 213196 73561
rect 212876 66561 213196 73325
rect 212876 66325 212918 66561
rect 213154 66325 213196 66561
rect 212876 59561 213196 66325
rect 212876 59325 212918 59561
rect 213154 59325 213196 59561
rect 212876 52561 213196 59325
rect 212876 52325 212918 52561
rect 213154 52325 213196 52561
rect 212876 45561 213196 52325
rect 212876 45325 212918 45561
rect 213154 45325 213196 45561
rect 212876 38561 213196 45325
rect 212876 38325 212918 38561
rect 213154 38325 213196 38561
rect 212876 31561 213196 38325
rect 212876 31325 212918 31561
rect 213154 31325 213196 31561
rect 212876 24561 213196 31325
rect 212876 24325 212918 24561
rect 213154 24325 213196 24561
rect 212876 17561 213196 24325
rect 212876 17325 212918 17561
rect 213154 17325 213196 17561
rect 212876 10561 213196 17325
rect 212876 10325 212918 10561
rect 213154 10325 213196 10561
rect 212876 3561 213196 10325
rect 212876 3325 212918 3561
rect 213154 3325 213196 3561
rect 212876 -1706 213196 3325
rect 212876 -1942 212918 -1706
rect 213154 -1942 213196 -1706
rect 212876 -2026 213196 -1942
rect 212876 -2262 212918 -2026
rect 213154 -2262 213196 -2026
rect 212876 -2294 213196 -2262
rect 218144 705238 218464 706230
rect 218144 705002 218186 705238
rect 218422 705002 218464 705238
rect 218144 704918 218464 705002
rect 218144 704682 218186 704918
rect 218422 704682 218464 704918
rect 218144 695494 218464 704682
rect 218144 695258 218186 695494
rect 218422 695258 218464 695494
rect 218144 688494 218464 695258
rect 218144 688258 218186 688494
rect 218422 688258 218464 688494
rect 218144 681494 218464 688258
rect 218144 681258 218186 681494
rect 218422 681258 218464 681494
rect 218144 674494 218464 681258
rect 218144 674258 218186 674494
rect 218422 674258 218464 674494
rect 218144 667494 218464 674258
rect 218144 667258 218186 667494
rect 218422 667258 218464 667494
rect 218144 660494 218464 667258
rect 218144 660258 218186 660494
rect 218422 660258 218464 660494
rect 218144 653494 218464 660258
rect 218144 653258 218186 653494
rect 218422 653258 218464 653494
rect 218144 646494 218464 653258
rect 218144 646258 218186 646494
rect 218422 646258 218464 646494
rect 218144 639494 218464 646258
rect 218144 639258 218186 639494
rect 218422 639258 218464 639494
rect 218144 632494 218464 639258
rect 218144 632258 218186 632494
rect 218422 632258 218464 632494
rect 218144 625494 218464 632258
rect 218144 625258 218186 625494
rect 218422 625258 218464 625494
rect 218144 618494 218464 625258
rect 218144 618258 218186 618494
rect 218422 618258 218464 618494
rect 218144 611494 218464 618258
rect 218144 611258 218186 611494
rect 218422 611258 218464 611494
rect 218144 604494 218464 611258
rect 218144 604258 218186 604494
rect 218422 604258 218464 604494
rect 218144 597494 218464 604258
rect 218144 597258 218186 597494
rect 218422 597258 218464 597494
rect 218144 590494 218464 597258
rect 218144 590258 218186 590494
rect 218422 590258 218464 590494
rect 218144 583494 218464 590258
rect 218144 583258 218186 583494
rect 218422 583258 218464 583494
rect 218144 576494 218464 583258
rect 218144 576258 218186 576494
rect 218422 576258 218464 576494
rect 218144 569494 218464 576258
rect 218144 569258 218186 569494
rect 218422 569258 218464 569494
rect 218144 562494 218464 569258
rect 218144 562258 218186 562494
rect 218422 562258 218464 562494
rect 218144 555494 218464 562258
rect 218144 555258 218186 555494
rect 218422 555258 218464 555494
rect 218144 548494 218464 555258
rect 218144 548258 218186 548494
rect 218422 548258 218464 548494
rect 218144 541494 218464 548258
rect 218144 541258 218186 541494
rect 218422 541258 218464 541494
rect 218144 534494 218464 541258
rect 218144 534258 218186 534494
rect 218422 534258 218464 534494
rect 218144 527494 218464 534258
rect 218144 527258 218186 527494
rect 218422 527258 218464 527494
rect 218144 520494 218464 527258
rect 218144 520258 218186 520494
rect 218422 520258 218464 520494
rect 218144 513494 218464 520258
rect 218144 513258 218186 513494
rect 218422 513258 218464 513494
rect 218144 506494 218464 513258
rect 218144 506258 218186 506494
rect 218422 506258 218464 506494
rect 218144 499494 218464 506258
rect 218144 499258 218186 499494
rect 218422 499258 218464 499494
rect 218144 492494 218464 499258
rect 218144 492258 218186 492494
rect 218422 492258 218464 492494
rect 218144 485494 218464 492258
rect 218144 485258 218186 485494
rect 218422 485258 218464 485494
rect 218144 478494 218464 485258
rect 218144 478258 218186 478494
rect 218422 478258 218464 478494
rect 218144 471494 218464 478258
rect 218144 471258 218186 471494
rect 218422 471258 218464 471494
rect 218144 464494 218464 471258
rect 218144 464258 218186 464494
rect 218422 464258 218464 464494
rect 218144 457494 218464 464258
rect 218144 457258 218186 457494
rect 218422 457258 218464 457494
rect 218144 450494 218464 457258
rect 218144 450258 218186 450494
rect 218422 450258 218464 450494
rect 218144 443494 218464 450258
rect 218144 443258 218186 443494
rect 218422 443258 218464 443494
rect 218144 436494 218464 443258
rect 218144 436258 218186 436494
rect 218422 436258 218464 436494
rect 218144 429494 218464 436258
rect 218144 429258 218186 429494
rect 218422 429258 218464 429494
rect 218144 422494 218464 429258
rect 218144 422258 218186 422494
rect 218422 422258 218464 422494
rect 218144 415494 218464 422258
rect 218144 415258 218186 415494
rect 218422 415258 218464 415494
rect 218144 408494 218464 415258
rect 218144 408258 218186 408494
rect 218422 408258 218464 408494
rect 218144 401494 218464 408258
rect 218144 401258 218186 401494
rect 218422 401258 218464 401494
rect 218144 394494 218464 401258
rect 218144 394258 218186 394494
rect 218422 394258 218464 394494
rect 218144 387494 218464 394258
rect 218144 387258 218186 387494
rect 218422 387258 218464 387494
rect 218144 380494 218464 387258
rect 218144 380258 218186 380494
rect 218422 380258 218464 380494
rect 218144 373494 218464 380258
rect 218144 373258 218186 373494
rect 218422 373258 218464 373494
rect 218144 366494 218464 373258
rect 218144 366258 218186 366494
rect 218422 366258 218464 366494
rect 218144 359494 218464 366258
rect 218144 359258 218186 359494
rect 218422 359258 218464 359494
rect 218144 352494 218464 359258
rect 218144 352258 218186 352494
rect 218422 352258 218464 352494
rect 218144 345494 218464 352258
rect 218144 345258 218186 345494
rect 218422 345258 218464 345494
rect 218144 338494 218464 345258
rect 218144 338258 218186 338494
rect 218422 338258 218464 338494
rect 218144 331494 218464 338258
rect 218144 331258 218186 331494
rect 218422 331258 218464 331494
rect 218144 324494 218464 331258
rect 218144 324258 218186 324494
rect 218422 324258 218464 324494
rect 218144 317494 218464 324258
rect 218144 317258 218186 317494
rect 218422 317258 218464 317494
rect 218144 310494 218464 317258
rect 218144 310258 218186 310494
rect 218422 310258 218464 310494
rect 218144 303494 218464 310258
rect 218144 303258 218186 303494
rect 218422 303258 218464 303494
rect 218144 296494 218464 303258
rect 218144 296258 218186 296494
rect 218422 296258 218464 296494
rect 218144 289494 218464 296258
rect 218144 289258 218186 289494
rect 218422 289258 218464 289494
rect 218144 282494 218464 289258
rect 218144 282258 218186 282494
rect 218422 282258 218464 282494
rect 218144 275494 218464 282258
rect 218144 275258 218186 275494
rect 218422 275258 218464 275494
rect 218144 268494 218464 275258
rect 218144 268258 218186 268494
rect 218422 268258 218464 268494
rect 218144 261494 218464 268258
rect 218144 261258 218186 261494
rect 218422 261258 218464 261494
rect 218144 254494 218464 261258
rect 218144 254258 218186 254494
rect 218422 254258 218464 254494
rect 218144 247494 218464 254258
rect 218144 247258 218186 247494
rect 218422 247258 218464 247494
rect 218144 240494 218464 247258
rect 218144 240258 218186 240494
rect 218422 240258 218464 240494
rect 218144 233494 218464 240258
rect 218144 233258 218186 233494
rect 218422 233258 218464 233494
rect 218144 226494 218464 233258
rect 218144 226258 218186 226494
rect 218422 226258 218464 226494
rect 218144 219494 218464 226258
rect 218144 219258 218186 219494
rect 218422 219258 218464 219494
rect 218144 212494 218464 219258
rect 218144 212258 218186 212494
rect 218422 212258 218464 212494
rect 218144 205494 218464 212258
rect 218144 205258 218186 205494
rect 218422 205258 218464 205494
rect 218144 198494 218464 205258
rect 218144 198258 218186 198494
rect 218422 198258 218464 198494
rect 218144 191494 218464 198258
rect 218144 191258 218186 191494
rect 218422 191258 218464 191494
rect 218144 184494 218464 191258
rect 218144 184258 218186 184494
rect 218422 184258 218464 184494
rect 218144 177494 218464 184258
rect 218144 177258 218186 177494
rect 218422 177258 218464 177494
rect 218144 170494 218464 177258
rect 218144 170258 218186 170494
rect 218422 170258 218464 170494
rect 218144 163494 218464 170258
rect 218144 163258 218186 163494
rect 218422 163258 218464 163494
rect 218144 156494 218464 163258
rect 218144 156258 218186 156494
rect 218422 156258 218464 156494
rect 218144 149494 218464 156258
rect 218144 149258 218186 149494
rect 218422 149258 218464 149494
rect 218144 142494 218464 149258
rect 218144 142258 218186 142494
rect 218422 142258 218464 142494
rect 218144 135494 218464 142258
rect 218144 135258 218186 135494
rect 218422 135258 218464 135494
rect 218144 128494 218464 135258
rect 218144 128258 218186 128494
rect 218422 128258 218464 128494
rect 218144 121494 218464 128258
rect 218144 121258 218186 121494
rect 218422 121258 218464 121494
rect 218144 114494 218464 121258
rect 218144 114258 218186 114494
rect 218422 114258 218464 114494
rect 218144 107494 218464 114258
rect 218144 107258 218186 107494
rect 218422 107258 218464 107494
rect 218144 100494 218464 107258
rect 218144 100258 218186 100494
rect 218422 100258 218464 100494
rect 218144 93494 218464 100258
rect 218144 93258 218186 93494
rect 218422 93258 218464 93494
rect 218144 86494 218464 93258
rect 218144 86258 218186 86494
rect 218422 86258 218464 86494
rect 218144 79494 218464 86258
rect 218144 79258 218186 79494
rect 218422 79258 218464 79494
rect 218144 72494 218464 79258
rect 218144 72258 218186 72494
rect 218422 72258 218464 72494
rect 218144 65494 218464 72258
rect 218144 65258 218186 65494
rect 218422 65258 218464 65494
rect 218144 58494 218464 65258
rect 218144 58258 218186 58494
rect 218422 58258 218464 58494
rect 218144 51494 218464 58258
rect 218144 51258 218186 51494
rect 218422 51258 218464 51494
rect 218144 44494 218464 51258
rect 218144 44258 218186 44494
rect 218422 44258 218464 44494
rect 218144 37494 218464 44258
rect 218144 37258 218186 37494
rect 218422 37258 218464 37494
rect 218144 30494 218464 37258
rect 218144 30258 218186 30494
rect 218422 30258 218464 30494
rect 218144 23494 218464 30258
rect 218144 23258 218186 23494
rect 218422 23258 218464 23494
rect 218144 16494 218464 23258
rect 218144 16258 218186 16494
rect 218422 16258 218464 16494
rect 218144 9494 218464 16258
rect 218144 9258 218186 9494
rect 218422 9258 218464 9494
rect 218144 2494 218464 9258
rect 218144 2258 218186 2494
rect 218422 2258 218464 2494
rect 218144 -746 218464 2258
rect 218144 -982 218186 -746
rect 218422 -982 218464 -746
rect 218144 -1066 218464 -982
rect 218144 -1302 218186 -1066
rect 218422 -1302 218464 -1066
rect 218144 -2294 218464 -1302
rect 219876 706198 220196 706230
rect 219876 705962 219918 706198
rect 220154 705962 220196 706198
rect 219876 705878 220196 705962
rect 219876 705642 219918 705878
rect 220154 705642 220196 705878
rect 219876 696561 220196 705642
rect 219876 696325 219918 696561
rect 220154 696325 220196 696561
rect 219876 689561 220196 696325
rect 219876 689325 219918 689561
rect 220154 689325 220196 689561
rect 219876 682561 220196 689325
rect 219876 682325 219918 682561
rect 220154 682325 220196 682561
rect 219876 675561 220196 682325
rect 219876 675325 219918 675561
rect 220154 675325 220196 675561
rect 219876 668561 220196 675325
rect 219876 668325 219918 668561
rect 220154 668325 220196 668561
rect 219876 661561 220196 668325
rect 219876 661325 219918 661561
rect 220154 661325 220196 661561
rect 219876 654561 220196 661325
rect 219876 654325 219918 654561
rect 220154 654325 220196 654561
rect 219876 647561 220196 654325
rect 219876 647325 219918 647561
rect 220154 647325 220196 647561
rect 219876 640561 220196 647325
rect 219876 640325 219918 640561
rect 220154 640325 220196 640561
rect 219876 633561 220196 640325
rect 219876 633325 219918 633561
rect 220154 633325 220196 633561
rect 219876 626561 220196 633325
rect 219876 626325 219918 626561
rect 220154 626325 220196 626561
rect 219876 619561 220196 626325
rect 219876 619325 219918 619561
rect 220154 619325 220196 619561
rect 219876 612561 220196 619325
rect 219876 612325 219918 612561
rect 220154 612325 220196 612561
rect 219876 605561 220196 612325
rect 219876 605325 219918 605561
rect 220154 605325 220196 605561
rect 219876 598561 220196 605325
rect 219876 598325 219918 598561
rect 220154 598325 220196 598561
rect 219876 591561 220196 598325
rect 219876 591325 219918 591561
rect 220154 591325 220196 591561
rect 219876 584561 220196 591325
rect 219876 584325 219918 584561
rect 220154 584325 220196 584561
rect 219876 577561 220196 584325
rect 219876 577325 219918 577561
rect 220154 577325 220196 577561
rect 219876 570561 220196 577325
rect 219876 570325 219918 570561
rect 220154 570325 220196 570561
rect 219876 563561 220196 570325
rect 219876 563325 219918 563561
rect 220154 563325 220196 563561
rect 219876 556561 220196 563325
rect 219876 556325 219918 556561
rect 220154 556325 220196 556561
rect 219876 549561 220196 556325
rect 219876 549325 219918 549561
rect 220154 549325 220196 549561
rect 219876 542561 220196 549325
rect 219876 542325 219918 542561
rect 220154 542325 220196 542561
rect 219876 535561 220196 542325
rect 219876 535325 219918 535561
rect 220154 535325 220196 535561
rect 219876 528561 220196 535325
rect 219876 528325 219918 528561
rect 220154 528325 220196 528561
rect 219876 521561 220196 528325
rect 219876 521325 219918 521561
rect 220154 521325 220196 521561
rect 219876 514561 220196 521325
rect 219876 514325 219918 514561
rect 220154 514325 220196 514561
rect 219876 507561 220196 514325
rect 219876 507325 219918 507561
rect 220154 507325 220196 507561
rect 219876 500561 220196 507325
rect 219876 500325 219918 500561
rect 220154 500325 220196 500561
rect 219876 493561 220196 500325
rect 219876 493325 219918 493561
rect 220154 493325 220196 493561
rect 219876 486561 220196 493325
rect 219876 486325 219918 486561
rect 220154 486325 220196 486561
rect 219876 479561 220196 486325
rect 219876 479325 219918 479561
rect 220154 479325 220196 479561
rect 219876 472561 220196 479325
rect 219876 472325 219918 472561
rect 220154 472325 220196 472561
rect 219876 465561 220196 472325
rect 219876 465325 219918 465561
rect 220154 465325 220196 465561
rect 219876 458561 220196 465325
rect 219876 458325 219918 458561
rect 220154 458325 220196 458561
rect 219876 451561 220196 458325
rect 219876 451325 219918 451561
rect 220154 451325 220196 451561
rect 219876 444561 220196 451325
rect 219876 444325 219918 444561
rect 220154 444325 220196 444561
rect 219876 437561 220196 444325
rect 219876 437325 219918 437561
rect 220154 437325 220196 437561
rect 219876 430561 220196 437325
rect 219876 430325 219918 430561
rect 220154 430325 220196 430561
rect 219876 423561 220196 430325
rect 219876 423325 219918 423561
rect 220154 423325 220196 423561
rect 219876 416561 220196 423325
rect 219876 416325 219918 416561
rect 220154 416325 220196 416561
rect 219876 409561 220196 416325
rect 219876 409325 219918 409561
rect 220154 409325 220196 409561
rect 219876 402561 220196 409325
rect 219876 402325 219918 402561
rect 220154 402325 220196 402561
rect 219876 395561 220196 402325
rect 219876 395325 219918 395561
rect 220154 395325 220196 395561
rect 219876 388561 220196 395325
rect 219876 388325 219918 388561
rect 220154 388325 220196 388561
rect 219876 381561 220196 388325
rect 219876 381325 219918 381561
rect 220154 381325 220196 381561
rect 219876 374561 220196 381325
rect 219876 374325 219918 374561
rect 220154 374325 220196 374561
rect 219876 367561 220196 374325
rect 219876 367325 219918 367561
rect 220154 367325 220196 367561
rect 219876 360561 220196 367325
rect 219876 360325 219918 360561
rect 220154 360325 220196 360561
rect 219876 353561 220196 360325
rect 219876 353325 219918 353561
rect 220154 353325 220196 353561
rect 219876 346561 220196 353325
rect 219876 346325 219918 346561
rect 220154 346325 220196 346561
rect 219876 339561 220196 346325
rect 219876 339325 219918 339561
rect 220154 339325 220196 339561
rect 219876 332561 220196 339325
rect 219876 332325 219918 332561
rect 220154 332325 220196 332561
rect 219876 325561 220196 332325
rect 219876 325325 219918 325561
rect 220154 325325 220196 325561
rect 219876 318561 220196 325325
rect 219876 318325 219918 318561
rect 220154 318325 220196 318561
rect 219876 311561 220196 318325
rect 219876 311325 219918 311561
rect 220154 311325 220196 311561
rect 219876 304561 220196 311325
rect 219876 304325 219918 304561
rect 220154 304325 220196 304561
rect 219876 297561 220196 304325
rect 219876 297325 219918 297561
rect 220154 297325 220196 297561
rect 219876 290561 220196 297325
rect 219876 290325 219918 290561
rect 220154 290325 220196 290561
rect 219876 283561 220196 290325
rect 219876 283325 219918 283561
rect 220154 283325 220196 283561
rect 219876 276561 220196 283325
rect 219876 276325 219918 276561
rect 220154 276325 220196 276561
rect 219876 269561 220196 276325
rect 219876 269325 219918 269561
rect 220154 269325 220196 269561
rect 219876 262561 220196 269325
rect 219876 262325 219918 262561
rect 220154 262325 220196 262561
rect 219876 255561 220196 262325
rect 219876 255325 219918 255561
rect 220154 255325 220196 255561
rect 219876 248561 220196 255325
rect 219876 248325 219918 248561
rect 220154 248325 220196 248561
rect 219876 241561 220196 248325
rect 219876 241325 219918 241561
rect 220154 241325 220196 241561
rect 219876 234561 220196 241325
rect 219876 234325 219918 234561
rect 220154 234325 220196 234561
rect 219876 227561 220196 234325
rect 219876 227325 219918 227561
rect 220154 227325 220196 227561
rect 219876 220561 220196 227325
rect 219876 220325 219918 220561
rect 220154 220325 220196 220561
rect 219876 213561 220196 220325
rect 219876 213325 219918 213561
rect 220154 213325 220196 213561
rect 219876 206561 220196 213325
rect 219876 206325 219918 206561
rect 220154 206325 220196 206561
rect 219876 199561 220196 206325
rect 219876 199325 219918 199561
rect 220154 199325 220196 199561
rect 219876 192561 220196 199325
rect 219876 192325 219918 192561
rect 220154 192325 220196 192561
rect 219876 185561 220196 192325
rect 219876 185325 219918 185561
rect 220154 185325 220196 185561
rect 219876 178561 220196 185325
rect 219876 178325 219918 178561
rect 220154 178325 220196 178561
rect 219876 171561 220196 178325
rect 219876 171325 219918 171561
rect 220154 171325 220196 171561
rect 219876 164561 220196 171325
rect 219876 164325 219918 164561
rect 220154 164325 220196 164561
rect 219876 157561 220196 164325
rect 219876 157325 219918 157561
rect 220154 157325 220196 157561
rect 219876 150561 220196 157325
rect 219876 150325 219918 150561
rect 220154 150325 220196 150561
rect 219876 143561 220196 150325
rect 219876 143325 219918 143561
rect 220154 143325 220196 143561
rect 219876 136561 220196 143325
rect 219876 136325 219918 136561
rect 220154 136325 220196 136561
rect 219876 129561 220196 136325
rect 219876 129325 219918 129561
rect 220154 129325 220196 129561
rect 219876 122561 220196 129325
rect 219876 122325 219918 122561
rect 220154 122325 220196 122561
rect 219876 115561 220196 122325
rect 219876 115325 219918 115561
rect 220154 115325 220196 115561
rect 219876 108561 220196 115325
rect 219876 108325 219918 108561
rect 220154 108325 220196 108561
rect 219876 101561 220196 108325
rect 219876 101325 219918 101561
rect 220154 101325 220196 101561
rect 219876 94561 220196 101325
rect 219876 94325 219918 94561
rect 220154 94325 220196 94561
rect 219876 87561 220196 94325
rect 219876 87325 219918 87561
rect 220154 87325 220196 87561
rect 219876 80561 220196 87325
rect 219876 80325 219918 80561
rect 220154 80325 220196 80561
rect 219876 73561 220196 80325
rect 219876 73325 219918 73561
rect 220154 73325 220196 73561
rect 219876 66561 220196 73325
rect 219876 66325 219918 66561
rect 220154 66325 220196 66561
rect 219876 59561 220196 66325
rect 219876 59325 219918 59561
rect 220154 59325 220196 59561
rect 219876 52561 220196 59325
rect 219876 52325 219918 52561
rect 220154 52325 220196 52561
rect 219876 45561 220196 52325
rect 219876 45325 219918 45561
rect 220154 45325 220196 45561
rect 219876 38561 220196 45325
rect 219876 38325 219918 38561
rect 220154 38325 220196 38561
rect 219876 31561 220196 38325
rect 219876 31325 219918 31561
rect 220154 31325 220196 31561
rect 219876 24561 220196 31325
rect 219876 24325 219918 24561
rect 220154 24325 220196 24561
rect 219876 17561 220196 24325
rect 219876 17325 219918 17561
rect 220154 17325 220196 17561
rect 219876 10561 220196 17325
rect 219876 10325 219918 10561
rect 220154 10325 220196 10561
rect 219876 3561 220196 10325
rect 219876 3325 219918 3561
rect 220154 3325 220196 3561
rect 219876 -1706 220196 3325
rect 219876 -1942 219918 -1706
rect 220154 -1942 220196 -1706
rect 219876 -2026 220196 -1942
rect 219876 -2262 219918 -2026
rect 220154 -2262 220196 -2026
rect 219876 -2294 220196 -2262
rect 225144 705238 225464 706230
rect 225144 705002 225186 705238
rect 225422 705002 225464 705238
rect 225144 704918 225464 705002
rect 225144 704682 225186 704918
rect 225422 704682 225464 704918
rect 225144 695494 225464 704682
rect 225144 695258 225186 695494
rect 225422 695258 225464 695494
rect 225144 688494 225464 695258
rect 225144 688258 225186 688494
rect 225422 688258 225464 688494
rect 225144 681494 225464 688258
rect 225144 681258 225186 681494
rect 225422 681258 225464 681494
rect 225144 674494 225464 681258
rect 225144 674258 225186 674494
rect 225422 674258 225464 674494
rect 225144 667494 225464 674258
rect 225144 667258 225186 667494
rect 225422 667258 225464 667494
rect 225144 660494 225464 667258
rect 225144 660258 225186 660494
rect 225422 660258 225464 660494
rect 225144 653494 225464 660258
rect 225144 653258 225186 653494
rect 225422 653258 225464 653494
rect 225144 646494 225464 653258
rect 225144 646258 225186 646494
rect 225422 646258 225464 646494
rect 225144 639494 225464 646258
rect 225144 639258 225186 639494
rect 225422 639258 225464 639494
rect 225144 632494 225464 639258
rect 225144 632258 225186 632494
rect 225422 632258 225464 632494
rect 225144 625494 225464 632258
rect 225144 625258 225186 625494
rect 225422 625258 225464 625494
rect 225144 618494 225464 625258
rect 225144 618258 225186 618494
rect 225422 618258 225464 618494
rect 225144 611494 225464 618258
rect 225144 611258 225186 611494
rect 225422 611258 225464 611494
rect 225144 604494 225464 611258
rect 225144 604258 225186 604494
rect 225422 604258 225464 604494
rect 225144 597494 225464 604258
rect 225144 597258 225186 597494
rect 225422 597258 225464 597494
rect 225144 590494 225464 597258
rect 225144 590258 225186 590494
rect 225422 590258 225464 590494
rect 225144 583494 225464 590258
rect 225144 583258 225186 583494
rect 225422 583258 225464 583494
rect 225144 576494 225464 583258
rect 225144 576258 225186 576494
rect 225422 576258 225464 576494
rect 225144 569494 225464 576258
rect 225144 569258 225186 569494
rect 225422 569258 225464 569494
rect 225144 562494 225464 569258
rect 225144 562258 225186 562494
rect 225422 562258 225464 562494
rect 225144 555494 225464 562258
rect 225144 555258 225186 555494
rect 225422 555258 225464 555494
rect 225144 548494 225464 555258
rect 225144 548258 225186 548494
rect 225422 548258 225464 548494
rect 225144 541494 225464 548258
rect 225144 541258 225186 541494
rect 225422 541258 225464 541494
rect 225144 534494 225464 541258
rect 225144 534258 225186 534494
rect 225422 534258 225464 534494
rect 225144 527494 225464 534258
rect 225144 527258 225186 527494
rect 225422 527258 225464 527494
rect 225144 520494 225464 527258
rect 225144 520258 225186 520494
rect 225422 520258 225464 520494
rect 225144 513494 225464 520258
rect 225144 513258 225186 513494
rect 225422 513258 225464 513494
rect 225144 506494 225464 513258
rect 225144 506258 225186 506494
rect 225422 506258 225464 506494
rect 225144 499494 225464 506258
rect 225144 499258 225186 499494
rect 225422 499258 225464 499494
rect 225144 492494 225464 499258
rect 225144 492258 225186 492494
rect 225422 492258 225464 492494
rect 225144 485494 225464 492258
rect 225144 485258 225186 485494
rect 225422 485258 225464 485494
rect 225144 478494 225464 485258
rect 225144 478258 225186 478494
rect 225422 478258 225464 478494
rect 225144 471494 225464 478258
rect 225144 471258 225186 471494
rect 225422 471258 225464 471494
rect 225144 464494 225464 471258
rect 225144 464258 225186 464494
rect 225422 464258 225464 464494
rect 225144 457494 225464 464258
rect 225144 457258 225186 457494
rect 225422 457258 225464 457494
rect 225144 450494 225464 457258
rect 225144 450258 225186 450494
rect 225422 450258 225464 450494
rect 225144 443494 225464 450258
rect 225144 443258 225186 443494
rect 225422 443258 225464 443494
rect 225144 436494 225464 443258
rect 225144 436258 225186 436494
rect 225422 436258 225464 436494
rect 225144 429494 225464 436258
rect 225144 429258 225186 429494
rect 225422 429258 225464 429494
rect 225144 422494 225464 429258
rect 225144 422258 225186 422494
rect 225422 422258 225464 422494
rect 225144 415494 225464 422258
rect 225144 415258 225186 415494
rect 225422 415258 225464 415494
rect 225144 408494 225464 415258
rect 225144 408258 225186 408494
rect 225422 408258 225464 408494
rect 225144 401494 225464 408258
rect 225144 401258 225186 401494
rect 225422 401258 225464 401494
rect 225144 394494 225464 401258
rect 225144 394258 225186 394494
rect 225422 394258 225464 394494
rect 225144 387494 225464 394258
rect 225144 387258 225186 387494
rect 225422 387258 225464 387494
rect 225144 380494 225464 387258
rect 225144 380258 225186 380494
rect 225422 380258 225464 380494
rect 225144 373494 225464 380258
rect 225144 373258 225186 373494
rect 225422 373258 225464 373494
rect 225144 366494 225464 373258
rect 225144 366258 225186 366494
rect 225422 366258 225464 366494
rect 225144 359494 225464 366258
rect 225144 359258 225186 359494
rect 225422 359258 225464 359494
rect 225144 352494 225464 359258
rect 225144 352258 225186 352494
rect 225422 352258 225464 352494
rect 225144 345494 225464 352258
rect 225144 345258 225186 345494
rect 225422 345258 225464 345494
rect 225144 338494 225464 345258
rect 225144 338258 225186 338494
rect 225422 338258 225464 338494
rect 225144 331494 225464 338258
rect 225144 331258 225186 331494
rect 225422 331258 225464 331494
rect 225144 324494 225464 331258
rect 225144 324258 225186 324494
rect 225422 324258 225464 324494
rect 225144 317494 225464 324258
rect 225144 317258 225186 317494
rect 225422 317258 225464 317494
rect 225144 310494 225464 317258
rect 225144 310258 225186 310494
rect 225422 310258 225464 310494
rect 225144 303494 225464 310258
rect 225144 303258 225186 303494
rect 225422 303258 225464 303494
rect 225144 296494 225464 303258
rect 225144 296258 225186 296494
rect 225422 296258 225464 296494
rect 225144 289494 225464 296258
rect 225144 289258 225186 289494
rect 225422 289258 225464 289494
rect 225144 282494 225464 289258
rect 225144 282258 225186 282494
rect 225422 282258 225464 282494
rect 225144 275494 225464 282258
rect 225144 275258 225186 275494
rect 225422 275258 225464 275494
rect 225144 268494 225464 275258
rect 225144 268258 225186 268494
rect 225422 268258 225464 268494
rect 225144 261494 225464 268258
rect 225144 261258 225186 261494
rect 225422 261258 225464 261494
rect 225144 254494 225464 261258
rect 225144 254258 225186 254494
rect 225422 254258 225464 254494
rect 225144 247494 225464 254258
rect 225144 247258 225186 247494
rect 225422 247258 225464 247494
rect 225144 240494 225464 247258
rect 225144 240258 225186 240494
rect 225422 240258 225464 240494
rect 225144 233494 225464 240258
rect 225144 233258 225186 233494
rect 225422 233258 225464 233494
rect 225144 226494 225464 233258
rect 225144 226258 225186 226494
rect 225422 226258 225464 226494
rect 225144 219494 225464 226258
rect 225144 219258 225186 219494
rect 225422 219258 225464 219494
rect 225144 212494 225464 219258
rect 225144 212258 225186 212494
rect 225422 212258 225464 212494
rect 225144 205494 225464 212258
rect 225144 205258 225186 205494
rect 225422 205258 225464 205494
rect 225144 198494 225464 205258
rect 225144 198258 225186 198494
rect 225422 198258 225464 198494
rect 225144 191494 225464 198258
rect 225144 191258 225186 191494
rect 225422 191258 225464 191494
rect 225144 184494 225464 191258
rect 225144 184258 225186 184494
rect 225422 184258 225464 184494
rect 225144 177494 225464 184258
rect 225144 177258 225186 177494
rect 225422 177258 225464 177494
rect 225144 170494 225464 177258
rect 225144 170258 225186 170494
rect 225422 170258 225464 170494
rect 225144 163494 225464 170258
rect 225144 163258 225186 163494
rect 225422 163258 225464 163494
rect 225144 156494 225464 163258
rect 225144 156258 225186 156494
rect 225422 156258 225464 156494
rect 225144 149494 225464 156258
rect 225144 149258 225186 149494
rect 225422 149258 225464 149494
rect 225144 142494 225464 149258
rect 225144 142258 225186 142494
rect 225422 142258 225464 142494
rect 225144 135494 225464 142258
rect 225144 135258 225186 135494
rect 225422 135258 225464 135494
rect 225144 128494 225464 135258
rect 225144 128258 225186 128494
rect 225422 128258 225464 128494
rect 225144 121494 225464 128258
rect 225144 121258 225186 121494
rect 225422 121258 225464 121494
rect 225144 114494 225464 121258
rect 225144 114258 225186 114494
rect 225422 114258 225464 114494
rect 225144 107494 225464 114258
rect 225144 107258 225186 107494
rect 225422 107258 225464 107494
rect 225144 100494 225464 107258
rect 225144 100258 225186 100494
rect 225422 100258 225464 100494
rect 225144 93494 225464 100258
rect 225144 93258 225186 93494
rect 225422 93258 225464 93494
rect 225144 86494 225464 93258
rect 225144 86258 225186 86494
rect 225422 86258 225464 86494
rect 225144 79494 225464 86258
rect 225144 79258 225186 79494
rect 225422 79258 225464 79494
rect 225144 72494 225464 79258
rect 225144 72258 225186 72494
rect 225422 72258 225464 72494
rect 225144 65494 225464 72258
rect 225144 65258 225186 65494
rect 225422 65258 225464 65494
rect 225144 58494 225464 65258
rect 225144 58258 225186 58494
rect 225422 58258 225464 58494
rect 225144 51494 225464 58258
rect 225144 51258 225186 51494
rect 225422 51258 225464 51494
rect 225144 44494 225464 51258
rect 225144 44258 225186 44494
rect 225422 44258 225464 44494
rect 225144 37494 225464 44258
rect 225144 37258 225186 37494
rect 225422 37258 225464 37494
rect 225144 30494 225464 37258
rect 225144 30258 225186 30494
rect 225422 30258 225464 30494
rect 225144 23494 225464 30258
rect 225144 23258 225186 23494
rect 225422 23258 225464 23494
rect 225144 16494 225464 23258
rect 225144 16258 225186 16494
rect 225422 16258 225464 16494
rect 225144 9494 225464 16258
rect 225144 9258 225186 9494
rect 225422 9258 225464 9494
rect 225144 2494 225464 9258
rect 225144 2258 225186 2494
rect 225422 2258 225464 2494
rect 225144 -746 225464 2258
rect 225144 -982 225186 -746
rect 225422 -982 225464 -746
rect 225144 -1066 225464 -982
rect 225144 -1302 225186 -1066
rect 225422 -1302 225464 -1066
rect 225144 -2294 225464 -1302
rect 226876 706198 227196 706230
rect 226876 705962 226918 706198
rect 227154 705962 227196 706198
rect 226876 705878 227196 705962
rect 226876 705642 226918 705878
rect 227154 705642 227196 705878
rect 226876 696561 227196 705642
rect 226876 696325 226918 696561
rect 227154 696325 227196 696561
rect 226876 689561 227196 696325
rect 226876 689325 226918 689561
rect 227154 689325 227196 689561
rect 226876 682561 227196 689325
rect 226876 682325 226918 682561
rect 227154 682325 227196 682561
rect 226876 675561 227196 682325
rect 226876 675325 226918 675561
rect 227154 675325 227196 675561
rect 226876 668561 227196 675325
rect 226876 668325 226918 668561
rect 227154 668325 227196 668561
rect 226876 661561 227196 668325
rect 226876 661325 226918 661561
rect 227154 661325 227196 661561
rect 226876 654561 227196 661325
rect 226876 654325 226918 654561
rect 227154 654325 227196 654561
rect 226876 647561 227196 654325
rect 226876 647325 226918 647561
rect 227154 647325 227196 647561
rect 226876 640561 227196 647325
rect 226876 640325 226918 640561
rect 227154 640325 227196 640561
rect 226876 633561 227196 640325
rect 226876 633325 226918 633561
rect 227154 633325 227196 633561
rect 226876 626561 227196 633325
rect 226876 626325 226918 626561
rect 227154 626325 227196 626561
rect 226876 619561 227196 626325
rect 226876 619325 226918 619561
rect 227154 619325 227196 619561
rect 226876 612561 227196 619325
rect 226876 612325 226918 612561
rect 227154 612325 227196 612561
rect 226876 605561 227196 612325
rect 226876 605325 226918 605561
rect 227154 605325 227196 605561
rect 226876 598561 227196 605325
rect 226876 598325 226918 598561
rect 227154 598325 227196 598561
rect 226876 591561 227196 598325
rect 226876 591325 226918 591561
rect 227154 591325 227196 591561
rect 226876 584561 227196 591325
rect 226876 584325 226918 584561
rect 227154 584325 227196 584561
rect 226876 577561 227196 584325
rect 226876 577325 226918 577561
rect 227154 577325 227196 577561
rect 226876 570561 227196 577325
rect 226876 570325 226918 570561
rect 227154 570325 227196 570561
rect 226876 563561 227196 570325
rect 226876 563325 226918 563561
rect 227154 563325 227196 563561
rect 226876 556561 227196 563325
rect 226876 556325 226918 556561
rect 227154 556325 227196 556561
rect 226876 549561 227196 556325
rect 226876 549325 226918 549561
rect 227154 549325 227196 549561
rect 226876 542561 227196 549325
rect 226876 542325 226918 542561
rect 227154 542325 227196 542561
rect 226876 535561 227196 542325
rect 226876 535325 226918 535561
rect 227154 535325 227196 535561
rect 226876 528561 227196 535325
rect 226876 528325 226918 528561
rect 227154 528325 227196 528561
rect 226876 521561 227196 528325
rect 226876 521325 226918 521561
rect 227154 521325 227196 521561
rect 226876 514561 227196 521325
rect 226876 514325 226918 514561
rect 227154 514325 227196 514561
rect 226876 507561 227196 514325
rect 226876 507325 226918 507561
rect 227154 507325 227196 507561
rect 226876 500561 227196 507325
rect 226876 500325 226918 500561
rect 227154 500325 227196 500561
rect 226876 493561 227196 500325
rect 226876 493325 226918 493561
rect 227154 493325 227196 493561
rect 226876 486561 227196 493325
rect 226876 486325 226918 486561
rect 227154 486325 227196 486561
rect 226876 479561 227196 486325
rect 226876 479325 226918 479561
rect 227154 479325 227196 479561
rect 226876 472561 227196 479325
rect 226876 472325 226918 472561
rect 227154 472325 227196 472561
rect 226876 465561 227196 472325
rect 226876 465325 226918 465561
rect 227154 465325 227196 465561
rect 226876 458561 227196 465325
rect 226876 458325 226918 458561
rect 227154 458325 227196 458561
rect 226876 451561 227196 458325
rect 226876 451325 226918 451561
rect 227154 451325 227196 451561
rect 226876 444561 227196 451325
rect 226876 444325 226918 444561
rect 227154 444325 227196 444561
rect 226876 437561 227196 444325
rect 226876 437325 226918 437561
rect 227154 437325 227196 437561
rect 226876 430561 227196 437325
rect 226876 430325 226918 430561
rect 227154 430325 227196 430561
rect 226876 423561 227196 430325
rect 226876 423325 226918 423561
rect 227154 423325 227196 423561
rect 226876 416561 227196 423325
rect 226876 416325 226918 416561
rect 227154 416325 227196 416561
rect 226876 409561 227196 416325
rect 226876 409325 226918 409561
rect 227154 409325 227196 409561
rect 226876 402561 227196 409325
rect 226876 402325 226918 402561
rect 227154 402325 227196 402561
rect 226876 395561 227196 402325
rect 226876 395325 226918 395561
rect 227154 395325 227196 395561
rect 226876 388561 227196 395325
rect 226876 388325 226918 388561
rect 227154 388325 227196 388561
rect 226876 381561 227196 388325
rect 226876 381325 226918 381561
rect 227154 381325 227196 381561
rect 226876 374561 227196 381325
rect 226876 374325 226918 374561
rect 227154 374325 227196 374561
rect 226876 367561 227196 374325
rect 226876 367325 226918 367561
rect 227154 367325 227196 367561
rect 226876 360561 227196 367325
rect 226876 360325 226918 360561
rect 227154 360325 227196 360561
rect 226876 353561 227196 360325
rect 226876 353325 226918 353561
rect 227154 353325 227196 353561
rect 226876 346561 227196 353325
rect 226876 346325 226918 346561
rect 227154 346325 227196 346561
rect 226876 339561 227196 346325
rect 226876 339325 226918 339561
rect 227154 339325 227196 339561
rect 226876 332561 227196 339325
rect 226876 332325 226918 332561
rect 227154 332325 227196 332561
rect 226876 325561 227196 332325
rect 226876 325325 226918 325561
rect 227154 325325 227196 325561
rect 226876 318561 227196 325325
rect 226876 318325 226918 318561
rect 227154 318325 227196 318561
rect 226876 311561 227196 318325
rect 226876 311325 226918 311561
rect 227154 311325 227196 311561
rect 226876 304561 227196 311325
rect 226876 304325 226918 304561
rect 227154 304325 227196 304561
rect 226876 297561 227196 304325
rect 226876 297325 226918 297561
rect 227154 297325 227196 297561
rect 226876 290561 227196 297325
rect 226876 290325 226918 290561
rect 227154 290325 227196 290561
rect 226876 283561 227196 290325
rect 226876 283325 226918 283561
rect 227154 283325 227196 283561
rect 226876 276561 227196 283325
rect 226876 276325 226918 276561
rect 227154 276325 227196 276561
rect 226876 269561 227196 276325
rect 226876 269325 226918 269561
rect 227154 269325 227196 269561
rect 226876 262561 227196 269325
rect 226876 262325 226918 262561
rect 227154 262325 227196 262561
rect 226876 255561 227196 262325
rect 226876 255325 226918 255561
rect 227154 255325 227196 255561
rect 226876 248561 227196 255325
rect 226876 248325 226918 248561
rect 227154 248325 227196 248561
rect 226876 241561 227196 248325
rect 226876 241325 226918 241561
rect 227154 241325 227196 241561
rect 226876 234561 227196 241325
rect 226876 234325 226918 234561
rect 227154 234325 227196 234561
rect 226876 227561 227196 234325
rect 226876 227325 226918 227561
rect 227154 227325 227196 227561
rect 226876 220561 227196 227325
rect 226876 220325 226918 220561
rect 227154 220325 227196 220561
rect 226876 213561 227196 220325
rect 226876 213325 226918 213561
rect 227154 213325 227196 213561
rect 226876 206561 227196 213325
rect 226876 206325 226918 206561
rect 227154 206325 227196 206561
rect 226876 199561 227196 206325
rect 226876 199325 226918 199561
rect 227154 199325 227196 199561
rect 226876 192561 227196 199325
rect 226876 192325 226918 192561
rect 227154 192325 227196 192561
rect 226876 185561 227196 192325
rect 226876 185325 226918 185561
rect 227154 185325 227196 185561
rect 226876 178561 227196 185325
rect 226876 178325 226918 178561
rect 227154 178325 227196 178561
rect 226876 171561 227196 178325
rect 226876 171325 226918 171561
rect 227154 171325 227196 171561
rect 226876 164561 227196 171325
rect 226876 164325 226918 164561
rect 227154 164325 227196 164561
rect 226876 157561 227196 164325
rect 226876 157325 226918 157561
rect 227154 157325 227196 157561
rect 226876 150561 227196 157325
rect 226876 150325 226918 150561
rect 227154 150325 227196 150561
rect 226876 143561 227196 150325
rect 226876 143325 226918 143561
rect 227154 143325 227196 143561
rect 226876 136561 227196 143325
rect 226876 136325 226918 136561
rect 227154 136325 227196 136561
rect 226876 129561 227196 136325
rect 226876 129325 226918 129561
rect 227154 129325 227196 129561
rect 226876 122561 227196 129325
rect 226876 122325 226918 122561
rect 227154 122325 227196 122561
rect 226876 115561 227196 122325
rect 226876 115325 226918 115561
rect 227154 115325 227196 115561
rect 226876 108561 227196 115325
rect 226876 108325 226918 108561
rect 227154 108325 227196 108561
rect 226876 101561 227196 108325
rect 226876 101325 226918 101561
rect 227154 101325 227196 101561
rect 226876 94561 227196 101325
rect 226876 94325 226918 94561
rect 227154 94325 227196 94561
rect 226876 87561 227196 94325
rect 226876 87325 226918 87561
rect 227154 87325 227196 87561
rect 226876 80561 227196 87325
rect 226876 80325 226918 80561
rect 227154 80325 227196 80561
rect 226876 73561 227196 80325
rect 226876 73325 226918 73561
rect 227154 73325 227196 73561
rect 226876 66561 227196 73325
rect 226876 66325 226918 66561
rect 227154 66325 227196 66561
rect 226876 59561 227196 66325
rect 226876 59325 226918 59561
rect 227154 59325 227196 59561
rect 226876 52561 227196 59325
rect 226876 52325 226918 52561
rect 227154 52325 227196 52561
rect 226876 45561 227196 52325
rect 226876 45325 226918 45561
rect 227154 45325 227196 45561
rect 226876 38561 227196 45325
rect 226876 38325 226918 38561
rect 227154 38325 227196 38561
rect 226876 31561 227196 38325
rect 226876 31325 226918 31561
rect 227154 31325 227196 31561
rect 226876 24561 227196 31325
rect 226876 24325 226918 24561
rect 227154 24325 227196 24561
rect 226876 17561 227196 24325
rect 226876 17325 226918 17561
rect 227154 17325 227196 17561
rect 226876 10561 227196 17325
rect 226876 10325 226918 10561
rect 227154 10325 227196 10561
rect 226876 3561 227196 10325
rect 226876 3325 226918 3561
rect 227154 3325 227196 3561
rect 226876 -1706 227196 3325
rect 226876 -1942 226918 -1706
rect 227154 -1942 227196 -1706
rect 226876 -2026 227196 -1942
rect 226876 -2262 226918 -2026
rect 227154 -2262 227196 -2026
rect 226876 -2294 227196 -2262
rect 232144 705238 232464 706230
rect 232144 705002 232186 705238
rect 232422 705002 232464 705238
rect 232144 704918 232464 705002
rect 232144 704682 232186 704918
rect 232422 704682 232464 704918
rect 232144 695494 232464 704682
rect 232144 695258 232186 695494
rect 232422 695258 232464 695494
rect 232144 688494 232464 695258
rect 232144 688258 232186 688494
rect 232422 688258 232464 688494
rect 232144 681494 232464 688258
rect 232144 681258 232186 681494
rect 232422 681258 232464 681494
rect 232144 674494 232464 681258
rect 232144 674258 232186 674494
rect 232422 674258 232464 674494
rect 232144 667494 232464 674258
rect 232144 667258 232186 667494
rect 232422 667258 232464 667494
rect 232144 660494 232464 667258
rect 232144 660258 232186 660494
rect 232422 660258 232464 660494
rect 232144 653494 232464 660258
rect 232144 653258 232186 653494
rect 232422 653258 232464 653494
rect 232144 646494 232464 653258
rect 232144 646258 232186 646494
rect 232422 646258 232464 646494
rect 232144 639494 232464 646258
rect 232144 639258 232186 639494
rect 232422 639258 232464 639494
rect 232144 632494 232464 639258
rect 232144 632258 232186 632494
rect 232422 632258 232464 632494
rect 232144 625494 232464 632258
rect 232144 625258 232186 625494
rect 232422 625258 232464 625494
rect 232144 618494 232464 625258
rect 232144 618258 232186 618494
rect 232422 618258 232464 618494
rect 232144 611494 232464 618258
rect 232144 611258 232186 611494
rect 232422 611258 232464 611494
rect 232144 604494 232464 611258
rect 232144 604258 232186 604494
rect 232422 604258 232464 604494
rect 232144 597494 232464 604258
rect 232144 597258 232186 597494
rect 232422 597258 232464 597494
rect 232144 590494 232464 597258
rect 232144 590258 232186 590494
rect 232422 590258 232464 590494
rect 232144 583494 232464 590258
rect 232144 583258 232186 583494
rect 232422 583258 232464 583494
rect 232144 576494 232464 583258
rect 232144 576258 232186 576494
rect 232422 576258 232464 576494
rect 232144 569494 232464 576258
rect 232144 569258 232186 569494
rect 232422 569258 232464 569494
rect 232144 562494 232464 569258
rect 232144 562258 232186 562494
rect 232422 562258 232464 562494
rect 232144 555494 232464 562258
rect 232144 555258 232186 555494
rect 232422 555258 232464 555494
rect 232144 548494 232464 555258
rect 232144 548258 232186 548494
rect 232422 548258 232464 548494
rect 232144 541494 232464 548258
rect 232144 541258 232186 541494
rect 232422 541258 232464 541494
rect 232144 534494 232464 541258
rect 232144 534258 232186 534494
rect 232422 534258 232464 534494
rect 232144 527494 232464 534258
rect 232144 527258 232186 527494
rect 232422 527258 232464 527494
rect 232144 520494 232464 527258
rect 232144 520258 232186 520494
rect 232422 520258 232464 520494
rect 232144 513494 232464 520258
rect 232144 513258 232186 513494
rect 232422 513258 232464 513494
rect 232144 506494 232464 513258
rect 232144 506258 232186 506494
rect 232422 506258 232464 506494
rect 232144 499494 232464 506258
rect 232144 499258 232186 499494
rect 232422 499258 232464 499494
rect 232144 492494 232464 499258
rect 232144 492258 232186 492494
rect 232422 492258 232464 492494
rect 232144 485494 232464 492258
rect 232144 485258 232186 485494
rect 232422 485258 232464 485494
rect 232144 478494 232464 485258
rect 232144 478258 232186 478494
rect 232422 478258 232464 478494
rect 232144 471494 232464 478258
rect 232144 471258 232186 471494
rect 232422 471258 232464 471494
rect 232144 464494 232464 471258
rect 232144 464258 232186 464494
rect 232422 464258 232464 464494
rect 232144 457494 232464 464258
rect 232144 457258 232186 457494
rect 232422 457258 232464 457494
rect 232144 450494 232464 457258
rect 232144 450258 232186 450494
rect 232422 450258 232464 450494
rect 232144 443494 232464 450258
rect 232144 443258 232186 443494
rect 232422 443258 232464 443494
rect 232144 436494 232464 443258
rect 232144 436258 232186 436494
rect 232422 436258 232464 436494
rect 232144 429494 232464 436258
rect 232144 429258 232186 429494
rect 232422 429258 232464 429494
rect 232144 422494 232464 429258
rect 232144 422258 232186 422494
rect 232422 422258 232464 422494
rect 232144 415494 232464 422258
rect 232144 415258 232186 415494
rect 232422 415258 232464 415494
rect 232144 408494 232464 415258
rect 232144 408258 232186 408494
rect 232422 408258 232464 408494
rect 232144 401494 232464 408258
rect 232144 401258 232186 401494
rect 232422 401258 232464 401494
rect 232144 394494 232464 401258
rect 232144 394258 232186 394494
rect 232422 394258 232464 394494
rect 232144 387494 232464 394258
rect 232144 387258 232186 387494
rect 232422 387258 232464 387494
rect 232144 380494 232464 387258
rect 232144 380258 232186 380494
rect 232422 380258 232464 380494
rect 232144 373494 232464 380258
rect 232144 373258 232186 373494
rect 232422 373258 232464 373494
rect 232144 366494 232464 373258
rect 232144 366258 232186 366494
rect 232422 366258 232464 366494
rect 232144 359494 232464 366258
rect 232144 359258 232186 359494
rect 232422 359258 232464 359494
rect 232144 352494 232464 359258
rect 232144 352258 232186 352494
rect 232422 352258 232464 352494
rect 232144 345494 232464 352258
rect 232144 345258 232186 345494
rect 232422 345258 232464 345494
rect 232144 338494 232464 345258
rect 232144 338258 232186 338494
rect 232422 338258 232464 338494
rect 232144 331494 232464 338258
rect 232144 331258 232186 331494
rect 232422 331258 232464 331494
rect 232144 324494 232464 331258
rect 232144 324258 232186 324494
rect 232422 324258 232464 324494
rect 232144 317494 232464 324258
rect 232144 317258 232186 317494
rect 232422 317258 232464 317494
rect 232144 310494 232464 317258
rect 232144 310258 232186 310494
rect 232422 310258 232464 310494
rect 232144 303494 232464 310258
rect 232144 303258 232186 303494
rect 232422 303258 232464 303494
rect 232144 296494 232464 303258
rect 232144 296258 232186 296494
rect 232422 296258 232464 296494
rect 232144 289494 232464 296258
rect 232144 289258 232186 289494
rect 232422 289258 232464 289494
rect 232144 282494 232464 289258
rect 232144 282258 232186 282494
rect 232422 282258 232464 282494
rect 232144 275494 232464 282258
rect 232144 275258 232186 275494
rect 232422 275258 232464 275494
rect 232144 268494 232464 275258
rect 232144 268258 232186 268494
rect 232422 268258 232464 268494
rect 232144 261494 232464 268258
rect 232144 261258 232186 261494
rect 232422 261258 232464 261494
rect 232144 254494 232464 261258
rect 232144 254258 232186 254494
rect 232422 254258 232464 254494
rect 232144 247494 232464 254258
rect 232144 247258 232186 247494
rect 232422 247258 232464 247494
rect 232144 240494 232464 247258
rect 232144 240258 232186 240494
rect 232422 240258 232464 240494
rect 232144 233494 232464 240258
rect 232144 233258 232186 233494
rect 232422 233258 232464 233494
rect 232144 226494 232464 233258
rect 232144 226258 232186 226494
rect 232422 226258 232464 226494
rect 232144 219494 232464 226258
rect 232144 219258 232186 219494
rect 232422 219258 232464 219494
rect 232144 212494 232464 219258
rect 232144 212258 232186 212494
rect 232422 212258 232464 212494
rect 232144 205494 232464 212258
rect 232144 205258 232186 205494
rect 232422 205258 232464 205494
rect 232144 198494 232464 205258
rect 232144 198258 232186 198494
rect 232422 198258 232464 198494
rect 232144 191494 232464 198258
rect 232144 191258 232186 191494
rect 232422 191258 232464 191494
rect 232144 184494 232464 191258
rect 232144 184258 232186 184494
rect 232422 184258 232464 184494
rect 232144 177494 232464 184258
rect 232144 177258 232186 177494
rect 232422 177258 232464 177494
rect 232144 170494 232464 177258
rect 232144 170258 232186 170494
rect 232422 170258 232464 170494
rect 232144 163494 232464 170258
rect 232144 163258 232186 163494
rect 232422 163258 232464 163494
rect 232144 156494 232464 163258
rect 232144 156258 232186 156494
rect 232422 156258 232464 156494
rect 232144 149494 232464 156258
rect 232144 149258 232186 149494
rect 232422 149258 232464 149494
rect 232144 142494 232464 149258
rect 232144 142258 232186 142494
rect 232422 142258 232464 142494
rect 232144 135494 232464 142258
rect 232144 135258 232186 135494
rect 232422 135258 232464 135494
rect 232144 128494 232464 135258
rect 232144 128258 232186 128494
rect 232422 128258 232464 128494
rect 232144 121494 232464 128258
rect 232144 121258 232186 121494
rect 232422 121258 232464 121494
rect 232144 114494 232464 121258
rect 232144 114258 232186 114494
rect 232422 114258 232464 114494
rect 232144 107494 232464 114258
rect 232144 107258 232186 107494
rect 232422 107258 232464 107494
rect 232144 100494 232464 107258
rect 232144 100258 232186 100494
rect 232422 100258 232464 100494
rect 232144 93494 232464 100258
rect 232144 93258 232186 93494
rect 232422 93258 232464 93494
rect 232144 86494 232464 93258
rect 232144 86258 232186 86494
rect 232422 86258 232464 86494
rect 232144 79494 232464 86258
rect 232144 79258 232186 79494
rect 232422 79258 232464 79494
rect 232144 72494 232464 79258
rect 232144 72258 232186 72494
rect 232422 72258 232464 72494
rect 232144 65494 232464 72258
rect 232144 65258 232186 65494
rect 232422 65258 232464 65494
rect 232144 58494 232464 65258
rect 232144 58258 232186 58494
rect 232422 58258 232464 58494
rect 232144 51494 232464 58258
rect 232144 51258 232186 51494
rect 232422 51258 232464 51494
rect 232144 44494 232464 51258
rect 232144 44258 232186 44494
rect 232422 44258 232464 44494
rect 232144 37494 232464 44258
rect 232144 37258 232186 37494
rect 232422 37258 232464 37494
rect 232144 30494 232464 37258
rect 232144 30258 232186 30494
rect 232422 30258 232464 30494
rect 232144 23494 232464 30258
rect 232144 23258 232186 23494
rect 232422 23258 232464 23494
rect 232144 16494 232464 23258
rect 232144 16258 232186 16494
rect 232422 16258 232464 16494
rect 232144 9494 232464 16258
rect 232144 9258 232186 9494
rect 232422 9258 232464 9494
rect 232144 2494 232464 9258
rect 232144 2258 232186 2494
rect 232422 2258 232464 2494
rect 232144 -746 232464 2258
rect 232144 -982 232186 -746
rect 232422 -982 232464 -746
rect 232144 -1066 232464 -982
rect 232144 -1302 232186 -1066
rect 232422 -1302 232464 -1066
rect 232144 -2294 232464 -1302
rect 233876 706198 234196 706230
rect 233876 705962 233918 706198
rect 234154 705962 234196 706198
rect 233876 705878 234196 705962
rect 233876 705642 233918 705878
rect 234154 705642 234196 705878
rect 233876 696561 234196 705642
rect 233876 696325 233918 696561
rect 234154 696325 234196 696561
rect 233876 689561 234196 696325
rect 233876 689325 233918 689561
rect 234154 689325 234196 689561
rect 233876 682561 234196 689325
rect 233876 682325 233918 682561
rect 234154 682325 234196 682561
rect 233876 675561 234196 682325
rect 233876 675325 233918 675561
rect 234154 675325 234196 675561
rect 233876 668561 234196 675325
rect 233876 668325 233918 668561
rect 234154 668325 234196 668561
rect 233876 661561 234196 668325
rect 233876 661325 233918 661561
rect 234154 661325 234196 661561
rect 233876 654561 234196 661325
rect 233876 654325 233918 654561
rect 234154 654325 234196 654561
rect 233876 647561 234196 654325
rect 233876 647325 233918 647561
rect 234154 647325 234196 647561
rect 233876 640561 234196 647325
rect 233876 640325 233918 640561
rect 234154 640325 234196 640561
rect 233876 633561 234196 640325
rect 233876 633325 233918 633561
rect 234154 633325 234196 633561
rect 233876 626561 234196 633325
rect 233876 626325 233918 626561
rect 234154 626325 234196 626561
rect 233876 619561 234196 626325
rect 233876 619325 233918 619561
rect 234154 619325 234196 619561
rect 233876 612561 234196 619325
rect 233876 612325 233918 612561
rect 234154 612325 234196 612561
rect 233876 605561 234196 612325
rect 233876 605325 233918 605561
rect 234154 605325 234196 605561
rect 233876 598561 234196 605325
rect 233876 598325 233918 598561
rect 234154 598325 234196 598561
rect 233876 591561 234196 598325
rect 233876 591325 233918 591561
rect 234154 591325 234196 591561
rect 233876 584561 234196 591325
rect 233876 584325 233918 584561
rect 234154 584325 234196 584561
rect 233876 577561 234196 584325
rect 233876 577325 233918 577561
rect 234154 577325 234196 577561
rect 233876 570561 234196 577325
rect 233876 570325 233918 570561
rect 234154 570325 234196 570561
rect 233876 563561 234196 570325
rect 233876 563325 233918 563561
rect 234154 563325 234196 563561
rect 233876 556561 234196 563325
rect 233876 556325 233918 556561
rect 234154 556325 234196 556561
rect 233876 549561 234196 556325
rect 233876 549325 233918 549561
rect 234154 549325 234196 549561
rect 233876 542561 234196 549325
rect 233876 542325 233918 542561
rect 234154 542325 234196 542561
rect 233876 535561 234196 542325
rect 233876 535325 233918 535561
rect 234154 535325 234196 535561
rect 233876 528561 234196 535325
rect 233876 528325 233918 528561
rect 234154 528325 234196 528561
rect 233876 521561 234196 528325
rect 233876 521325 233918 521561
rect 234154 521325 234196 521561
rect 233876 514561 234196 521325
rect 233876 514325 233918 514561
rect 234154 514325 234196 514561
rect 233876 507561 234196 514325
rect 233876 507325 233918 507561
rect 234154 507325 234196 507561
rect 233876 500561 234196 507325
rect 233876 500325 233918 500561
rect 234154 500325 234196 500561
rect 233876 493561 234196 500325
rect 233876 493325 233918 493561
rect 234154 493325 234196 493561
rect 233876 486561 234196 493325
rect 233876 486325 233918 486561
rect 234154 486325 234196 486561
rect 233876 479561 234196 486325
rect 233876 479325 233918 479561
rect 234154 479325 234196 479561
rect 233876 472561 234196 479325
rect 233876 472325 233918 472561
rect 234154 472325 234196 472561
rect 233876 465561 234196 472325
rect 233876 465325 233918 465561
rect 234154 465325 234196 465561
rect 233876 458561 234196 465325
rect 233876 458325 233918 458561
rect 234154 458325 234196 458561
rect 233876 451561 234196 458325
rect 233876 451325 233918 451561
rect 234154 451325 234196 451561
rect 233876 444561 234196 451325
rect 233876 444325 233918 444561
rect 234154 444325 234196 444561
rect 233876 437561 234196 444325
rect 233876 437325 233918 437561
rect 234154 437325 234196 437561
rect 233876 430561 234196 437325
rect 233876 430325 233918 430561
rect 234154 430325 234196 430561
rect 233876 423561 234196 430325
rect 233876 423325 233918 423561
rect 234154 423325 234196 423561
rect 233876 416561 234196 423325
rect 233876 416325 233918 416561
rect 234154 416325 234196 416561
rect 233876 409561 234196 416325
rect 233876 409325 233918 409561
rect 234154 409325 234196 409561
rect 233876 402561 234196 409325
rect 233876 402325 233918 402561
rect 234154 402325 234196 402561
rect 233876 395561 234196 402325
rect 233876 395325 233918 395561
rect 234154 395325 234196 395561
rect 233876 388561 234196 395325
rect 233876 388325 233918 388561
rect 234154 388325 234196 388561
rect 233876 381561 234196 388325
rect 233876 381325 233918 381561
rect 234154 381325 234196 381561
rect 233876 374561 234196 381325
rect 233876 374325 233918 374561
rect 234154 374325 234196 374561
rect 233876 367561 234196 374325
rect 233876 367325 233918 367561
rect 234154 367325 234196 367561
rect 233876 360561 234196 367325
rect 233876 360325 233918 360561
rect 234154 360325 234196 360561
rect 233876 353561 234196 360325
rect 233876 353325 233918 353561
rect 234154 353325 234196 353561
rect 233876 346561 234196 353325
rect 233876 346325 233918 346561
rect 234154 346325 234196 346561
rect 233876 339561 234196 346325
rect 233876 339325 233918 339561
rect 234154 339325 234196 339561
rect 233876 332561 234196 339325
rect 233876 332325 233918 332561
rect 234154 332325 234196 332561
rect 233876 325561 234196 332325
rect 233876 325325 233918 325561
rect 234154 325325 234196 325561
rect 233876 318561 234196 325325
rect 233876 318325 233918 318561
rect 234154 318325 234196 318561
rect 233876 311561 234196 318325
rect 233876 311325 233918 311561
rect 234154 311325 234196 311561
rect 233876 304561 234196 311325
rect 233876 304325 233918 304561
rect 234154 304325 234196 304561
rect 233876 297561 234196 304325
rect 233876 297325 233918 297561
rect 234154 297325 234196 297561
rect 233876 290561 234196 297325
rect 233876 290325 233918 290561
rect 234154 290325 234196 290561
rect 233876 283561 234196 290325
rect 233876 283325 233918 283561
rect 234154 283325 234196 283561
rect 233876 276561 234196 283325
rect 233876 276325 233918 276561
rect 234154 276325 234196 276561
rect 233876 269561 234196 276325
rect 233876 269325 233918 269561
rect 234154 269325 234196 269561
rect 233876 262561 234196 269325
rect 233876 262325 233918 262561
rect 234154 262325 234196 262561
rect 233876 255561 234196 262325
rect 233876 255325 233918 255561
rect 234154 255325 234196 255561
rect 233876 248561 234196 255325
rect 233876 248325 233918 248561
rect 234154 248325 234196 248561
rect 233876 241561 234196 248325
rect 233876 241325 233918 241561
rect 234154 241325 234196 241561
rect 233876 234561 234196 241325
rect 233876 234325 233918 234561
rect 234154 234325 234196 234561
rect 233876 227561 234196 234325
rect 233876 227325 233918 227561
rect 234154 227325 234196 227561
rect 233876 220561 234196 227325
rect 233876 220325 233918 220561
rect 234154 220325 234196 220561
rect 233876 213561 234196 220325
rect 233876 213325 233918 213561
rect 234154 213325 234196 213561
rect 233876 206561 234196 213325
rect 233876 206325 233918 206561
rect 234154 206325 234196 206561
rect 233876 199561 234196 206325
rect 233876 199325 233918 199561
rect 234154 199325 234196 199561
rect 233876 192561 234196 199325
rect 233876 192325 233918 192561
rect 234154 192325 234196 192561
rect 233876 185561 234196 192325
rect 233876 185325 233918 185561
rect 234154 185325 234196 185561
rect 233876 178561 234196 185325
rect 233876 178325 233918 178561
rect 234154 178325 234196 178561
rect 233876 171561 234196 178325
rect 233876 171325 233918 171561
rect 234154 171325 234196 171561
rect 233876 164561 234196 171325
rect 233876 164325 233918 164561
rect 234154 164325 234196 164561
rect 233876 157561 234196 164325
rect 233876 157325 233918 157561
rect 234154 157325 234196 157561
rect 233876 150561 234196 157325
rect 233876 150325 233918 150561
rect 234154 150325 234196 150561
rect 233876 143561 234196 150325
rect 233876 143325 233918 143561
rect 234154 143325 234196 143561
rect 233876 136561 234196 143325
rect 233876 136325 233918 136561
rect 234154 136325 234196 136561
rect 233876 129561 234196 136325
rect 233876 129325 233918 129561
rect 234154 129325 234196 129561
rect 233876 122561 234196 129325
rect 233876 122325 233918 122561
rect 234154 122325 234196 122561
rect 233876 115561 234196 122325
rect 233876 115325 233918 115561
rect 234154 115325 234196 115561
rect 233876 108561 234196 115325
rect 233876 108325 233918 108561
rect 234154 108325 234196 108561
rect 233876 101561 234196 108325
rect 233876 101325 233918 101561
rect 234154 101325 234196 101561
rect 233876 94561 234196 101325
rect 233876 94325 233918 94561
rect 234154 94325 234196 94561
rect 233876 87561 234196 94325
rect 233876 87325 233918 87561
rect 234154 87325 234196 87561
rect 233876 80561 234196 87325
rect 233876 80325 233918 80561
rect 234154 80325 234196 80561
rect 233876 73561 234196 80325
rect 233876 73325 233918 73561
rect 234154 73325 234196 73561
rect 233876 66561 234196 73325
rect 233876 66325 233918 66561
rect 234154 66325 234196 66561
rect 233876 59561 234196 66325
rect 233876 59325 233918 59561
rect 234154 59325 234196 59561
rect 233876 52561 234196 59325
rect 233876 52325 233918 52561
rect 234154 52325 234196 52561
rect 233876 45561 234196 52325
rect 233876 45325 233918 45561
rect 234154 45325 234196 45561
rect 233876 38561 234196 45325
rect 233876 38325 233918 38561
rect 234154 38325 234196 38561
rect 233876 31561 234196 38325
rect 233876 31325 233918 31561
rect 234154 31325 234196 31561
rect 233876 24561 234196 31325
rect 233876 24325 233918 24561
rect 234154 24325 234196 24561
rect 233876 17561 234196 24325
rect 233876 17325 233918 17561
rect 234154 17325 234196 17561
rect 233876 10561 234196 17325
rect 233876 10325 233918 10561
rect 234154 10325 234196 10561
rect 233876 3561 234196 10325
rect 233876 3325 233918 3561
rect 234154 3325 234196 3561
rect 233876 -1706 234196 3325
rect 233876 -1942 233918 -1706
rect 234154 -1942 234196 -1706
rect 233876 -2026 234196 -1942
rect 233876 -2262 233918 -2026
rect 234154 -2262 234196 -2026
rect 233876 -2294 234196 -2262
rect 239144 705238 239464 706230
rect 239144 705002 239186 705238
rect 239422 705002 239464 705238
rect 239144 704918 239464 705002
rect 239144 704682 239186 704918
rect 239422 704682 239464 704918
rect 239144 695494 239464 704682
rect 239144 695258 239186 695494
rect 239422 695258 239464 695494
rect 239144 688494 239464 695258
rect 239144 688258 239186 688494
rect 239422 688258 239464 688494
rect 239144 681494 239464 688258
rect 239144 681258 239186 681494
rect 239422 681258 239464 681494
rect 239144 674494 239464 681258
rect 239144 674258 239186 674494
rect 239422 674258 239464 674494
rect 239144 667494 239464 674258
rect 239144 667258 239186 667494
rect 239422 667258 239464 667494
rect 239144 660494 239464 667258
rect 239144 660258 239186 660494
rect 239422 660258 239464 660494
rect 239144 653494 239464 660258
rect 239144 653258 239186 653494
rect 239422 653258 239464 653494
rect 239144 646494 239464 653258
rect 239144 646258 239186 646494
rect 239422 646258 239464 646494
rect 239144 639494 239464 646258
rect 239144 639258 239186 639494
rect 239422 639258 239464 639494
rect 239144 632494 239464 639258
rect 239144 632258 239186 632494
rect 239422 632258 239464 632494
rect 239144 625494 239464 632258
rect 239144 625258 239186 625494
rect 239422 625258 239464 625494
rect 239144 618494 239464 625258
rect 239144 618258 239186 618494
rect 239422 618258 239464 618494
rect 239144 611494 239464 618258
rect 239144 611258 239186 611494
rect 239422 611258 239464 611494
rect 239144 604494 239464 611258
rect 239144 604258 239186 604494
rect 239422 604258 239464 604494
rect 239144 597494 239464 604258
rect 239144 597258 239186 597494
rect 239422 597258 239464 597494
rect 239144 590494 239464 597258
rect 239144 590258 239186 590494
rect 239422 590258 239464 590494
rect 239144 583494 239464 590258
rect 239144 583258 239186 583494
rect 239422 583258 239464 583494
rect 239144 576494 239464 583258
rect 239144 576258 239186 576494
rect 239422 576258 239464 576494
rect 239144 569494 239464 576258
rect 239144 569258 239186 569494
rect 239422 569258 239464 569494
rect 239144 562494 239464 569258
rect 239144 562258 239186 562494
rect 239422 562258 239464 562494
rect 239144 555494 239464 562258
rect 239144 555258 239186 555494
rect 239422 555258 239464 555494
rect 239144 548494 239464 555258
rect 239144 548258 239186 548494
rect 239422 548258 239464 548494
rect 239144 541494 239464 548258
rect 239144 541258 239186 541494
rect 239422 541258 239464 541494
rect 239144 534494 239464 541258
rect 239144 534258 239186 534494
rect 239422 534258 239464 534494
rect 239144 527494 239464 534258
rect 239144 527258 239186 527494
rect 239422 527258 239464 527494
rect 239144 520494 239464 527258
rect 239144 520258 239186 520494
rect 239422 520258 239464 520494
rect 239144 513494 239464 520258
rect 239144 513258 239186 513494
rect 239422 513258 239464 513494
rect 239144 506494 239464 513258
rect 239144 506258 239186 506494
rect 239422 506258 239464 506494
rect 239144 499494 239464 506258
rect 239144 499258 239186 499494
rect 239422 499258 239464 499494
rect 239144 492494 239464 499258
rect 239144 492258 239186 492494
rect 239422 492258 239464 492494
rect 239144 485494 239464 492258
rect 239144 485258 239186 485494
rect 239422 485258 239464 485494
rect 239144 478494 239464 485258
rect 239144 478258 239186 478494
rect 239422 478258 239464 478494
rect 239144 471494 239464 478258
rect 239144 471258 239186 471494
rect 239422 471258 239464 471494
rect 239144 464494 239464 471258
rect 239144 464258 239186 464494
rect 239422 464258 239464 464494
rect 239144 457494 239464 464258
rect 239144 457258 239186 457494
rect 239422 457258 239464 457494
rect 239144 450494 239464 457258
rect 239144 450258 239186 450494
rect 239422 450258 239464 450494
rect 239144 443494 239464 450258
rect 239144 443258 239186 443494
rect 239422 443258 239464 443494
rect 239144 436494 239464 443258
rect 239144 436258 239186 436494
rect 239422 436258 239464 436494
rect 239144 429494 239464 436258
rect 239144 429258 239186 429494
rect 239422 429258 239464 429494
rect 239144 422494 239464 429258
rect 239144 422258 239186 422494
rect 239422 422258 239464 422494
rect 239144 415494 239464 422258
rect 239144 415258 239186 415494
rect 239422 415258 239464 415494
rect 239144 408494 239464 415258
rect 239144 408258 239186 408494
rect 239422 408258 239464 408494
rect 239144 401494 239464 408258
rect 239144 401258 239186 401494
rect 239422 401258 239464 401494
rect 239144 394494 239464 401258
rect 239144 394258 239186 394494
rect 239422 394258 239464 394494
rect 239144 387494 239464 394258
rect 239144 387258 239186 387494
rect 239422 387258 239464 387494
rect 239144 380494 239464 387258
rect 239144 380258 239186 380494
rect 239422 380258 239464 380494
rect 239144 373494 239464 380258
rect 239144 373258 239186 373494
rect 239422 373258 239464 373494
rect 239144 366494 239464 373258
rect 239144 366258 239186 366494
rect 239422 366258 239464 366494
rect 239144 359494 239464 366258
rect 239144 359258 239186 359494
rect 239422 359258 239464 359494
rect 239144 352494 239464 359258
rect 239144 352258 239186 352494
rect 239422 352258 239464 352494
rect 239144 345494 239464 352258
rect 239144 345258 239186 345494
rect 239422 345258 239464 345494
rect 239144 338494 239464 345258
rect 239144 338258 239186 338494
rect 239422 338258 239464 338494
rect 239144 331494 239464 338258
rect 239144 331258 239186 331494
rect 239422 331258 239464 331494
rect 239144 324494 239464 331258
rect 239144 324258 239186 324494
rect 239422 324258 239464 324494
rect 239144 317494 239464 324258
rect 239144 317258 239186 317494
rect 239422 317258 239464 317494
rect 239144 310494 239464 317258
rect 239144 310258 239186 310494
rect 239422 310258 239464 310494
rect 239144 303494 239464 310258
rect 239144 303258 239186 303494
rect 239422 303258 239464 303494
rect 239144 296494 239464 303258
rect 239144 296258 239186 296494
rect 239422 296258 239464 296494
rect 239144 289494 239464 296258
rect 239144 289258 239186 289494
rect 239422 289258 239464 289494
rect 239144 282494 239464 289258
rect 239144 282258 239186 282494
rect 239422 282258 239464 282494
rect 239144 275494 239464 282258
rect 239144 275258 239186 275494
rect 239422 275258 239464 275494
rect 239144 268494 239464 275258
rect 239144 268258 239186 268494
rect 239422 268258 239464 268494
rect 239144 261494 239464 268258
rect 239144 261258 239186 261494
rect 239422 261258 239464 261494
rect 239144 254494 239464 261258
rect 239144 254258 239186 254494
rect 239422 254258 239464 254494
rect 239144 247494 239464 254258
rect 239144 247258 239186 247494
rect 239422 247258 239464 247494
rect 239144 240494 239464 247258
rect 239144 240258 239186 240494
rect 239422 240258 239464 240494
rect 239144 233494 239464 240258
rect 239144 233258 239186 233494
rect 239422 233258 239464 233494
rect 239144 226494 239464 233258
rect 239144 226258 239186 226494
rect 239422 226258 239464 226494
rect 239144 219494 239464 226258
rect 239144 219258 239186 219494
rect 239422 219258 239464 219494
rect 239144 212494 239464 219258
rect 239144 212258 239186 212494
rect 239422 212258 239464 212494
rect 239144 205494 239464 212258
rect 239144 205258 239186 205494
rect 239422 205258 239464 205494
rect 239144 198494 239464 205258
rect 239144 198258 239186 198494
rect 239422 198258 239464 198494
rect 239144 191494 239464 198258
rect 239144 191258 239186 191494
rect 239422 191258 239464 191494
rect 239144 184494 239464 191258
rect 239144 184258 239186 184494
rect 239422 184258 239464 184494
rect 239144 177494 239464 184258
rect 239144 177258 239186 177494
rect 239422 177258 239464 177494
rect 239144 170494 239464 177258
rect 239144 170258 239186 170494
rect 239422 170258 239464 170494
rect 239144 163494 239464 170258
rect 239144 163258 239186 163494
rect 239422 163258 239464 163494
rect 239144 156494 239464 163258
rect 239144 156258 239186 156494
rect 239422 156258 239464 156494
rect 239144 149494 239464 156258
rect 239144 149258 239186 149494
rect 239422 149258 239464 149494
rect 239144 142494 239464 149258
rect 239144 142258 239186 142494
rect 239422 142258 239464 142494
rect 239144 135494 239464 142258
rect 239144 135258 239186 135494
rect 239422 135258 239464 135494
rect 239144 128494 239464 135258
rect 239144 128258 239186 128494
rect 239422 128258 239464 128494
rect 239144 121494 239464 128258
rect 239144 121258 239186 121494
rect 239422 121258 239464 121494
rect 239144 114494 239464 121258
rect 239144 114258 239186 114494
rect 239422 114258 239464 114494
rect 239144 107494 239464 114258
rect 239144 107258 239186 107494
rect 239422 107258 239464 107494
rect 239144 100494 239464 107258
rect 239144 100258 239186 100494
rect 239422 100258 239464 100494
rect 239144 93494 239464 100258
rect 239144 93258 239186 93494
rect 239422 93258 239464 93494
rect 239144 86494 239464 93258
rect 239144 86258 239186 86494
rect 239422 86258 239464 86494
rect 239144 79494 239464 86258
rect 239144 79258 239186 79494
rect 239422 79258 239464 79494
rect 239144 72494 239464 79258
rect 239144 72258 239186 72494
rect 239422 72258 239464 72494
rect 239144 65494 239464 72258
rect 239144 65258 239186 65494
rect 239422 65258 239464 65494
rect 239144 58494 239464 65258
rect 239144 58258 239186 58494
rect 239422 58258 239464 58494
rect 239144 51494 239464 58258
rect 239144 51258 239186 51494
rect 239422 51258 239464 51494
rect 239144 44494 239464 51258
rect 239144 44258 239186 44494
rect 239422 44258 239464 44494
rect 239144 37494 239464 44258
rect 239144 37258 239186 37494
rect 239422 37258 239464 37494
rect 239144 30494 239464 37258
rect 239144 30258 239186 30494
rect 239422 30258 239464 30494
rect 239144 23494 239464 30258
rect 239144 23258 239186 23494
rect 239422 23258 239464 23494
rect 239144 16494 239464 23258
rect 239144 16258 239186 16494
rect 239422 16258 239464 16494
rect 239144 9494 239464 16258
rect 239144 9258 239186 9494
rect 239422 9258 239464 9494
rect 239144 2494 239464 9258
rect 239144 2258 239186 2494
rect 239422 2258 239464 2494
rect 239144 -746 239464 2258
rect 239144 -982 239186 -746
rect 239422 -982 239464 -746
rect 239144 -1066 239464 -982
rect 239144 -1302 239186 -1066
rect 239422 -1302 239464 -1066
rect 239144 -2294 239464 -1302
rect 240876 706198 241196 706230
rect 240876 705962 240918 706198
rect 241154 705962 241196 706198
rect 240876 705878 241196 705962
rect 240876 705642 240918 705878
rect 241154 705642 241196 705878
rect 240876 696561 241196 705642
rect 240876 696325 240918 696561
rect 241154 696325 241196 696561
rect 240876 689561 241196 696325
rect 240876 689325 240918 689561
rect 241154 689325 241196 689561
rect 240876 682561 241196 689325
rect 240876 682325 240918 682561
rect 241154 682325 241196 682561
rect 240876 675561 241196 682325
rect 240876 675325 240918 675561
rect 241154 675325 241196 675561
rect 240876 668561 241196 675325
rect 240876 668325 240918 668561
rect 241154 668325 241196 668561
rect 240876 661561 241196 668325
rect 240876 661325 240918 661561
rect 241154 661325 241196 661561
rect 240876 654561 241196 661325
rect 240876 654325 240918 654561
rect 241154 654325 241196 654561
rect 240876 647561 241196 654325
rect 240876 647325 240918 647561
rect 241154 647325 241196 647561
rect 240876 640561 241196 647325
rect 240876 640325 240918 640561
rect 241154 640325 241196 640561
rect 240876 633561 241196 640325
rect 240876 633325 240918 633561
rect 241154 633325 241196 633561
rect 240876 626561 241196 633325
rect 240876 626325 240918 626561
rect 241154 626325 241196 626561
rect 240876 619561 241196 626325
rect 240876 619325 240918 619561
rect 241154 619325 241196 619561
rect 240876 612561 241196 619325
rect 240876 612325 240918 612561
rect 241154 612325 241196 612561
rect 240876 605561 241196 612325
rect 240876 605325 240918 605561
rect 241154 605325 241196 605561
rect 240876 598561 241196 605325
rect 240876 598325 240918 598561
rect 241154 598325 241196 598561
rect 240876 591561 241196 598325
rect 240876 591325 240918 591561
rect 241154 591325 241196 591561
rect 240876 584561 241196 591325
rect 240876 584325 240918 584561
rect 241154 584325 241196 584561
rect 240876 577561 241196 584325
rect 240876 577325 240918 577561
rect 241154 577325 241196 577561
rect 240876 570561 241196 577325
rect 240876 570325 240918 570561
rect 241154 570325 241196 570561
rect 240876 563561 241196 570325
rect 240876 563325 240918 563561
rect 241154 563325 241196 563561
rect 240876 556561 241196 563325
rect 240876 556325 240918 556561
rect 241154 556325 241196 556561
rect 240876 549561 241196 556325
rect 240876 549325 240918 549561
rect 241154 549325 241196 549561
rect 240876 542561 241196 549325
rect 240876 542325 240918 542561
rect 241154 542325 241196 542561
rect 240876 535561 241196 542325
rect 240876 535325 240918 535561
rect 241154 535325 241196 535561
rect 240876 528561 241196 535325
rect 240876 528325 240918 528561
rect 241154 528325 241196 528561
rect 240876 521561 241196 528325
rect 240876 521325 240918 521561
rect 241154 521325 241196 521561
rect 240876 514561 241196 521325
rect 240876 514325 240918 514561
rect 241154 514325 241196 514561
rect 240876 507561 241196 514325
rect 240876 507325 240918 507561
rect 241154 507325 241196 507561
rect 240876 500561 241196 507325
rect 240876 500325 240918 500561
rect 241154 500325 241196 500561
rect 240876 493561 241196 500325
rect 240876 493325 240918 493561
rect 241154 493325 241196 493561
rect 240876 486561 241196 493325
rect 240876 486325 240918 486561
rect 241154 486325 241196 486561
rect 240876 479561 241196 486325
rect 240876 479325 240918 479561
rect 241154 479325 241196 479561
rect 240876 472561 241196 479325
rect 240876 472325 240918 472561
rect 241154 472325 241196 472561
rect 240876 465561 241196 472325
rect 240876 465325 240918 465561
rect 241154 465325 241196 465561
rect 240876 458561 241196 465325
rect 240876 458325 240918 458561
rect 241154 458325 241196 458561
rect 240876 451561 241196 458325
rect 240876 451325 240918 451561
rect 241154 451325 241196 451561
rect 240876 444561 241196 451325
rect 240876 444325 240918 444561
rect 241154 444325 241196 444561
rect 240876 437561 241196 444325
rect 240876 437325 240918 437561
rect 241154 437325 241196 437561
rect 240876 430561 241196 437325
rect 240876 430325 240918 430561
rect 241154 430325 241196 430561
rect 240876 423561 241196 430325
rect 240876 423325 240918 423561
rect 241154 423325 241196 423561
rect 240876 416561 241196 423325
rect 240876 416325 240918 416561
rect 241154 416325 241196 416561
rect 240876 409561 241196 416325
rect 240876 409325 240918 409561
rect 241154 409325 241196 409561
rect 240876 402561 241196 409325
rect 240876 402325 240918 402561
rect 241154 402325 241196 402561
rect 240876 395561 241196 402325
rect 240876 395325 240918 395561
rect 241154 395325 241196 395561
rect 240876 388561 241196 395325
rect 240876 388325 240918 388561
rect 241154 388325 241196 388561
rect 240876 381561 241196 388325
rect 240876 381325 240918 381561
rect 241154 381325 241196 381561
rect 240876 374561 241196 381325
rect 240876 374325 240918 374561
rect 241154 374325 241196 374561
rect 240876 367561 241196 374325
rect 240876 367325 240918 367561
rect 241154 367325 241196 367561
rect 240876 360561 241196 367325
rect 240876 360325 240918 360561
rect 241154 360325 241196 360561
rect 240876 353561 241196 360325
rect 240876 353325 240918 353561
rect 241154 353325 241196 353561
rect 240876 346561 241196 353325
rect 240876 346325 240918 346561
rect 241154 346325 241196 346561
rect 240876 339561 241196 346325
rect 240876 339325 240918 339561
rect 241154 339325 241196 339561
rect 240876 332561 241196 339325
rect 240876 332325 240918 332561
rect 241154 332325 241196 332561
rect 240876 325561 241196 332325
rect 240876 325325 240918 325561
rect 241154 325325 241196 325561
rect 240876 318561 241196 325325
rect 240876 318325 240918 318561
rect 241154 318325 241196 318561
rect 240876 311561 241196 318325
rect 240876 311325 240918 311561
rect 241154 311325 241196 311561
rect 240876 304561 241196 311325
rect 240876 304325 240918 304561
rect 241154 304325 241196 304561
rect 240876 297561 241196 304325
rect 240876 297325 240918 297561
rect 241154 297325 241196 297561
rect 240876 290561 241196 297325
rect 240876 290325 240918 290561
rect 241154 290325 241196 290561
rect 240876 283561 241196 290325
rect 240876 283325 240918 283561
rect 241154 283325 241196 283561
rect 240876 276561 241196 283325
rect 240876 276325 240918 276561
rect 241154 276325 241196 276561
rect 240876 269561 241196 276325
rect 240876 269325 240918 269561
rect 241154 269325 241196 269561
rect 240876 262561 241196 269325
rect 240876 262325 240918 262561
rect 241154 262325 241196 262561
rect 240876 255561 241196 262325
rect 240876 255325 240918 255561
rect 241154 255325 241196 255561
rect 240876 248561 241196 255325
rect 240876 248325 240918 248561
rect 241154 248325 241196 248561
rect 240876 241561 241196 248325
rect 240876 241325 240918 241561
rect 241154 241325 241196 241561
rect 240876 234561 241196 241325
rect 240876 234325 240918 234561
rect 241154 234325 241196 234561
rect 240876 227561 241196 234325
rect 240876 227325 240918 227561
rect 241154 227325 241196 227561
rect 240876 220561 241196 227325
rect 240876 220325 240918 220561
rect 241154 220325 241196 220561
rect 240876 213561 241196 220325
rect 240876 213325 240918 213561
rect 241154 213325 241196 213561
rect 240876 206561 241196 213325
rect 240876 206325 240918 206561
rect 241154 206325 241196 206561
rect 240876 199561 241196 206325
rect 240876 199325 240918 199561
rect 241154 199325 241196 199561
rect 240876 192561 241196 199325
rect 240876 192325 240918 192561
rect 241154 192325 241196 192561
rect 240876 185561 241196 192325
rect 240876 185325 240918 185561
rect 241154 185325 241196 185561
rect 240876 178561 241196 185325
rect 240876 178325 240918 178561
rect 241154 178325 241196 178561
rect 240876 171561 241196 178325
rect 240876 171325 240918 171561
rect 241154 171325 241196 171561
rect 240876 164561 241196 171325
rect 240876 164325 240918 164561
rect 241154 164325 241196 164561
rect 240876 157561 241196 164325
rect 240876 157325 240918 157561
rect 241154 157325 241196 157561
rect 240876 150561 241196 157325
rect 240876 150325 240918 150561
rect 241154 150325 241196 150561
rect 240876 143561 241196 150325
rect 240876 143325 240918 143561
rect 241154 143325 241196 143561
rect 240876 136561 241196 143325
rect 240876 136325 240918 136561
rect 241154 136325 241196 136561
rect 240876 129561 241196 136325
rect 240876 129325 240918 129561
rect 241154 129325 241196 129561
rect 240876 122561 241196 129325
rect 240876 122325 240918 122561
rect 241154 122325 241196 122561
rect 240876 115561 241196 122325
rect 240876 115325 240918 115561
rect 241154 115325 241196 115561
rect 240876 108561 241196 115325
rect 240876 108325 240918 108561
rect 241154 108325 241196 108561
rect 240876 101561 241196 108325
rect 240876 101325 240918 101561
rect 241154 101325 241196 101561
rect 240876 94561 241196 101325
rect 240876 94325 240918 94561
rect 241154 94325 241196 94561
rect 240876 87561 241196 94325
rect 240876 87325 240918 87561
rect 241154 87325 241196 87561
rect 240876 80561 241196 87325
rect 240876 80325 240918 80561
rect 241154 80325 241196 80561
rect 240876 73561 241196 80325
rect 240876 73325 240918 73561
rect 241154 73325 241196 73561
rect 240876 66561 241196 73325
rect 240876 66325 240918 66561
rect 241154 66325 241196 66561
rect 240876 59561 241196 66325
rect 240876 59325 240918 59561
rect 241154 59325 241196 59561
rect 240876 52561 241196 59325
rect 240876 52325 240918 52561
rect 241154 52325 241196 52561
rect 240876 45561 241196 52325
rect 240876 45325 240918 45561
rect 241154 45325 241196 45561
rect 240876 38561 241196 45325
rect 240876 38325 240918 38561
rect 241154 38325 241196 38561
rect 240876 31561 241196 38325
rect 240876 31325 240918 31561
rect 241154 31325 241196 31561
rect 240876 24561 241196 31325
rect 240876 24325 240918 24561
rect 241154 24325 241196 24561
rect 240876 17561 241196 24325
rect 240876 17325 240918 17561
rect 241154 17325 241196 17561
rect 240876 10561 241196 17325
rect 240876 10325 240918 10561
rect 241154 10325 241196 10561
rect 240876 3561 241196 10325
rect 240876 3325 240918 3561
rect 241154 3325 241196 3561
rect 240876 -1706 241196 3325
rect 240876 -1942 240918 -1706
rect 241154 -1942 241196 -1706
rect 240876 -2026 241196 -1942
rect 240876 -2262 240918 -2026
rect 241154 -2262 241196 -2026
rect 240876 -2294 241196 -2262
rect 246144 705238 246464 706230
rect 246144 705002 246186 705238
rect 246422 705002 246464 705238
rect 246144 704918 246464 705002
rect 246144 704682 246186 704918
rect 246422 704682 246464 704918
rect 246144 695494 246464 704682
rect 246144 695258 246186 695494
rect 246422 695258 246464 695494
rect 246144 688494 246464 695258
rect 246144 688258 246186 688494
rect 246422 688258 246464 688494
rect 246144 681494 246464 688258
rect 246144 681258 246186 681494
rect 246422 681258 246464 681494
rect 246144 674494 246464 681258
rect 246144 674258 246186 674494
rect 246422 674258 246464 674494
rect 246144 667494 246464 674258
rect 246144 667258 246186 667494
rect 246422 667258 246464 667494
rect 246144 660494 246464 667258
rect 246144 660258 246186 660494
rect 246422 660258 246464 660494
rect 246144 653494 246464 660258
rect 246144 653258 246186 653494
rect 246422 653258 246464 653494
rect 246144 646494 246464 653258
rect 246144 646258 246186 646494
rect 246422 646258 246464 646494
rect 246144 639494 246464 646258
rect 246144 639258 246186 639494
rect 246422 639258 246464 639494
rect 246144 632494 246464 639258
rect 246144 632258 246186 632494
rect 246422 632258 246464 632494
rect 246144 625494 246464 632258
rect 246144 625258 246186 625494
rect 246422 625258 246464 625494
rect 246144 618494 246464 625258
rect 246144 618258 246186 618494
rect 246422 618258 246464 618494
rect 246144 611494 246464 618258
rect 246144 611258 246186 611494
rect 246422 611258 246464 611494
rect 246144 604494 246464 611258
rect 246144 604258 246186 604494
rect 246422 604258 246464 604494
rect 246144 597494 246464 604258
rect 246144 597258 246186 597494
rect 246422 597258 246464 597494
rect 246144 590494 246464 597258
rect 246144 590258 246186 590494
rect 246422 590258 246464 590494
rect 246144 583494 246464 590258
rect 246144 583258 246186 583494
rect 246422 583258 246464 583494
rect 246144 576494 246464 583258
rect 246144 576258 246186 576494
rect 246422 576258 246464 576494
rect 246144 569494 246464 576258
rect 246144 569258 246186 569494
rect 246422 569258 246464 569494
rect 246144 562494 246464 569258
rect 246144 562258 246186 562494
rect 246422 562258 246464 562494
rect 246144 555494 246464 562258
rect 246144 555258 246186 555494
rect 246422 555258 246464 555494
rect 246144 548494 246464 555258
rect 246144 548258 246186 548494
rect 246422 548258 246464 548494
rect 246144 541494 246464 548258
rect 246144 541258 246186 541494
rect 246422 541258 246464 541494
rect 246144 534494 246464 541258
rect 246144 534258 246186 534494
rect 246422 534258 246464 534494
rect 246144 527494 246464 534258
rect 246144 527258 246186 527494
rect 246422 527258 246464 527494
rect 246144 520494 246464 527258
rect 246144 520258 246186 520494
rect 246422 520258 246464 520494
rect 246144 513494 246464 520258
rect 246144 513258 246186 513494
rect 246422 513258 246464 513494
rect 246144 506494 246464 513258
rect 246144 506258 246186 506494
rect 246422 506258 246464 506494
rect 246144 499494 246464 506258
rect 246144 499258 246186 499494
rect 246422 499258 246464 499494
rect 246144 492494 246464 499258
rect 246144 492258 246186 492494
rect 246422 492258 246464 492494
rect 246144 485494 246464 492258
rect 246144 485258 246186 485494
rect 246422 485258 246464 485494
rect 246144 478494 246464 485258
rect 246144 478258 246186 478494
rect 246422 478258 246464 478494
rect 246144 471494 246464 478258
rect 246144 471258 246186 471494
rect 246422 471258 246464 471494
rect 246144 464494 246464 471258
rect 246144 464258 246186 464494
rect 246422 464258 246464 464494
rect 246144 457494 246464 464258
rect 246144 457258 246186 457494
rect 246422 457258 246464 457494
rect 246144 450494 246464 457258
rect 246144 450258 246186 450494
rect 246422 450258 246464 450494
rect 246144 443494 246464 450258
rect 246144 443258 246186 443494
rect 246422 443258 246464 443494
rect 246144 436494 246464 443258
rect 246144 436258 246186 436494
rect 246422 436258 246464 436494
rect 246144 429494 246464 436258
rect 246144 429258 246186 429494
rect 246422 429258 246464 429494
rect 246144 422494 246464 429258
rect 246144 422258 246186 422494
rect 246422 422258 246464 422494
rect 246144 415494 246464 422258
rect 246144 415258 246186 415494
rect 246422 415258 246464 415494
rect 246144 408494 246464 415258
rect 246144 408258 246186 408494
rect 246422 408258 246464 408494
rect 246144 401494 246464 408258
rect 246144 401258 246186 401494
rect 246422 401258 246464 401494
rect 246144 394494 246464 401258
rect 246144 394258 246186 394494
rect 246422 394258 246464 394494
rect 246144 387494 246464 394258
rect 246144 387258 246186 387494
rect 246422 387258 246464 387494
rect 246144 380494 246464 387258
rect 246144 380258 246186 380494
rect 246422 380258 246464 380494
rect 246144 373494 246464 380258
rect 246144 373258 246186 373494
rect 246422 373258 246464 373494
rect 246144 366494 246464 373258
rect 246144 366258 246186 366494
rect 246422 366258 246464 366494
rect 246144 359494 246464 366258
rect 246144 359258 246186 359494
rect 246422 359258 246464 359494
rect 246144 352494 246464 359258
rect 246144 352258 246186 352494
rect 246422 352258 246464 352494
rect 246144 345494 246464 352258
rect 246144 345258 246186 345494
rect 246422 345258 246464 345494
rect 246144 338494 246464 345258
rect 246144 338258 246186 338494
rect 246422 338258 246464 338494
rect 246144 331494 246464 338258
rect 246144 331258 246186 331494
rect 246422 331258 246464 331494
rect 246144 324494 246464 331258
rect 246144 324258 246186 324494
rect 246422 324258 246464 324494
rect 246144 317494 246464 324258
rect 246144 317258 246186 317494
rect 246422 317258 246464 317494
rect 246144 310494 246464 317258
rect 246144 310258 246186 310494
rect 246422 310258 246464 310494
rect 246144 303494 246464 310258
rect 246144 303258 246186 303494
rect 246422 303258 246464 303494
rect 246144 296494 246464 303258
rect 246144 296258 246186 296494
rect 246422 296258 246464 296494
rect 246144 289494 246464 296258
rect 246144 289258 246186 289494
rect 246422 289258 246464 289494
rect 246144 282494 246464 289258
rect 246144 282258 246186 282494
rect 246422 282258 246464 282494
rect 246144 275494 246464 282258
rect 246144 275258 246186 275494
rect 246422 275258 246464 275494
rect 246144 268494 246464 275258
rect 246144 268258 246186 268494
rect 246422 268258 246464 268494
rect 246144 261494 246464 268258
rect 246144 261258 246186 261494
rect 246422 261258 246464 261494
rect 246144 254494 246464 261258
rect 246144 254258 246186 254494
rect 246422 254258 246464 254494
rect 246144 247494 246464 254258
rect 246144 247258 246186 247494
rect 246422 247258 246464 247494
rect 246144 240494 246464 247258
rect 246144 240258 246186 240494
rect 246422 240258 246464 240494
rect 246144 233494 246464 240258
rect 246144 233258 246186 233494
rect 246422 233258 246464 233494
rect 246144 226494 246464 233258
rect 246144 226258 246186 226494
rect 246422 226258 246464 226494
rect 246144 219494 246464 226258
rect 246144 219258 246186 219494
rect 246422 219258 246464 219494
rect 246144 212494 246464 219258
rect 246144 212258 246186 212494
rect 246422 212258 246464 212494
rect 246144 205494 246464 212258
rect 246144 205258 246186 205494
rect 246422 205258 246464 205494
rect 246144 198494 246464 205258
rect 246144 198258 246186 198494
rect 246422 198258 246464 198494
rect 246144 191494 246464 198258
rect 246144 191258 246186 191494
rect 246422 191258 246464 191494
rect 246144 184494 246464 191258
rect 246144 184258 246186 184494
rect 246422 184258 246464 184494
rect 246144 177494 246464 184258
rect 246144 177258 246186 177494
rect 246422 177258 246464 177494
rect 246144 170494 246464 177258
rect 246144 170258 246186 170494
rect 246422 170258 246464 170494
rect 246144 163494 246464 170258
rect 246144 163258 246186 163494
rect 246422 163258 246464 163494
rect 246144 156494 246464 163258
rect 246144 156258 246186 156494
rect 246422 156258 246464 156494
rect 246144 149494 246464 156258
rect 246144 149258 246186 149494
rect 246422 149258 246464 149494
rect 246144 142494 246464 149258
rect 246144 142258 246186 142494
rect 246422 142258 246464 142494
rect 246144 135494 246464 142258
rect 246144 135258 246186 135494
rect 246422 135258 246464 135494
rect 246144 128494 246464 135258
rect 246144 128258 246186 128494
rect 246422 128258 246464 128494
rect 246144 121494 246464 128258
rect 246144 121258 246186 121494
rect 246422 121258 246464 121494
rect 246144 114494 246464 121258
rect 246144 114258 246186 114494
rect 246422 114258 246464 114494
rect 246144 107494 246464 114258
rect 246144 107258 246186 107494
rect 246422 107258 246464 107494
rect 246144 100494 246464 107258
rect 246144 100258 246186 100494
rect 246422 100258 246464 100494
rect 246144 93494 246464 100258
rect 246144 93258 246186 93494
rect 246422 93258 246464 93494
rect 246144 86494 246464 93258
rect 246144 86258 246186 86494
rect 246422 86258 246464 86494
rect 246144 79494 246464 86258
rect 246144 79258 246186 79494
rect 246422 79258 246464 79494
rect 246144 72494 246464 79258
rect 246144 72258 246186 72494
rect 246422 72258 246464 72494
rect 246144 65494 246464 72258
rect 246144 65258 246186 65494
rect 246422 65258 246464 65494
rect 246144 58494 246464 65258
rect 246144 58258 246186 58494
rect 246422 58258 246464 58494
rect 246144 51494 246464 58258
rect 246144 51258 246186 51494
rect 246422 51258 246464 51494
rect 246144 44494 246464 51258
rect 246144 44258 246186 44494
rect 246422 44258 246464 44494
rect 246144 37494 246464 44258
rect 246144 37258 246186 37494
rect 246422 37258 246464 37494
rect 246144 30494 246464 37258
rect 246144 30258 246186 30494
rect 246422 30258 246464 30494
rect 246144 23494 246464 30258
rect 246144 23258 246186 23494
rect 246422 23258 246464 23494
rect 246144 16494 246464 23258
rect 246144 16258 246186 16494
rect 246422 16258 246464 16494
rect 246144 9494 246464 16258
rect 246144 9258 246186 9494
rect 246422 9258 246464 9494
rect 246144 2494 246464 9258
rect 246144 2258 246186 2494
rect 246422 2258 246464 2494
rect 246144 -746 246464 2258
rect 246144 -982 246186 -746
rect 246422 -982 246464 -746
rect 246144 -1066 246464 -982
rect 246144 -1302 246186 -1066
rect 246422 -1302 246464 -1066
rect 246144 -2294 246464 -1302
rect 247876 706198 248196 706230
rect 247876 705962 247918 706198
rect 248154 705962 248196 706198
rect 247876 705878 248196 705962
rect 247876 705642 247918 705878
rect 248154 705642 248196 705878
rect 247876 696561 248196 705642
rect 247876 696325 247918 696561
rect 248154 696325 248196 696561
rect 247876 689561 248196 696325
rect 247876 689325 247918 689561
rect 248154 689325 248196 689561
rect 247876 682561 248196 689325
rect 247876 682325 247918 682561
rect 248154 682325 248196 682561
rect 247876 675561 248196 682325
rect 247876 675325 247918 675561
rect 248154 675325 248196 675561
rect 247876 668561 248196 675325
rect 247876 668325 247918 668561
rect 248154 668325 248196 668561
rect 247876 661561 248196 668325
rect 247876 661325 247918 661561
rect 248154 661325 248196 661561
rect 247876 654561 248196 661325
rect 247876 654325 247918 654561
rect 248154 654325 248196 654561
rect 247876 647561 248196 654325
rect 247876 647325 247918 647561
rect 248154 647325 248196 647561
rect 247876 640561 248196 647325
rect 247876 640325 247918 640561
rect 248154 640325 248196 640561
rect 247876 633561 248196 640325
rect 247876 633325 247918 633561
rect 248154 633325 248196 633561
rect 247876 626561 248196 633325
rect 247876 626325 247918 626561
rect 248154 626325 248196 626561
rect 247876 619561 248196 626325
rect 247876 619325 247918 619561
rect 248154 619325 248196 619561
rect 247876 612561 248196 619325
rect 247876 612325 247918 612561
rect 248154 612325 248196 612561
rect 247876 605561 248196 612325
rect 247876 605325 247918 605561
rect 248154 605325 248196 605561
rect 247876 598561 248196 605325
rect 247876 598325 247918 598561
rect 248154 598325 248196 598561
rect 247876 591561 248196 598325
rect 247876 591325 247918 591561
rect 248154 591325 248196 591561
rect 247876 584561 248196 591325
rect 247876 584325 247918 584561
rect 248154 584325 248196 584561
rect 247876 577561 248196 584325
rect 247876 577325 247918 577561
rect 248154 577325 248196 577561
rect 247876 570561 248196 577325
rect 247876 570325 247918 570561
rect 248154 570325 248196 570561
rect 247876 563561 248196 570325
rect 247876 563325 247918 563561
rect 248154 563325 248196 563561
rect 247876 556561 248196 563325
rect 247876 556325 247918 556561
rect 248154 556325 248196 556561
rect 247876 549561 248196 556325
rect 247876 549325 247918 549561
rect 248154 549325 248196 549561
rect 247876 542561 248196 549325
rect 247876 542325 247918 542561
rect 248154 542325 248196 542561
rect 247876 535561 248196 542325
rect 247876 535325 247918 535561
rect 248154 535325 248196 535561
rect 247876 528561 248196 535325
rect 247876 528325 247918 528561
rect 248154 528325 248196 528561
rect 247876 521561 248196 528325
rect 247876 521325 247918 521561
rect 248154 521325 248196 521561
rect 247876 514561 248196 521325
rect 247876 514325 247918 514561
rect 248154 514325 248196 514561
rect 247876 507561 248196 514325
rect 247876 507325 247918 507561
rect 248154 507325 248196 507561
rect 247876 500561 248196 507325
rect 247876 500325 247918 500561
rect 248154 500325 248196 500561
rect 247876 493561 248196 500325
rect 247876 493325 247918 493561
rect 248154 493325 248196 493561
rect 247876 486561 248196 493325
rect 247876 486325 247918 486561
rect 248154 486325 248196 486561
rect 247876 479561 248196 486325
rect 247876 479325 247918 479561
rect 248154 479325 248196 479561
rect 247876 472561 248196 479325
rect 247876 472325 247918 472561
rect 248154 472325 248196 472561
rect 247876 465561 248196 472325
rect 247876 465325 247918 465561
rect 248154 465325 248196 465561
rect 247876 458561 248196 465325
rect 247876 458325 247918 458561
rect 248154 458325 248196 458561
rect 247876 451561 248196 458325
rect 247876 451325 247918 451561
rect 248154 451325 248196 451561
rect 247876 444561 248196 451325
rect 247876 444325 247918 444561
rect 248154 444325 248196 444561
rect 247876 437561 248196 444325
rect 247876 437325 247918 437561
rect 248154 437325 248196 437561
rect 247876 430561 248196 437325
rect 247876 430325 247918 430561
rect 248154 430325 248196 430561
rect 247876 423561 248196 430325
rect 247876 423325 247918 423561
rect 248154 423325 248196 423561
rect 247876 416561 248196 423325
rect 247876 416325 247918 416561
rect 248154 416325 248196 416561
rect 247876 409561 248196 416325
rect 247876 409325 247918 409561
rect 248154 409325 248196 409561
rect 247876 402561 248196 409325
rect 247876 402325 247918 402561
rect 248154 402325 248196 402561
rect 247876 395561 248196 402325
rect 247876 395325 247918 395561
rect 248154 395325 248196 395561
rect 247876 388561 248196 395325
rect 247876 388325 247918 388561
rect 248154 388325 248196 388561
rect 247876 381561 248196 388325
rect 247876 381325 247918 381561
rect 248154 381325 248196 381561
rect 247876 374561 248196 381325
rect 247876 374325 247918 374561
rect 248154 374325 248196 374561
rect 247876 367561 248196 374325
rect 247876 367325 247918 367561
rect 248154 367325 248196 367561
rect 247876 360561 248196 367325
rect 247876 360325 247918 360561
rect 248154 360325 248196 360561
rect 247876 353561 248196 360325
rect 247876 353325 247918 353561
rect 248154 353325 248196 353561
rect 247876 346561 248196 353325
rect 247876 346325 247918 346561
rect 248154 346325 248196 346561
rect 247876 339561 248196 346325
rect 247876 339325 247918 339561
rect 248154 339325 248196 339561
rect 247876 332561 248196 339325
rect 247876 332325 247918 332561
rect 248154 332325 248196 332561
rect 247876 325561 248196 332325
rect 247876 325325 247918 325561
rect 248154 325325 248196 325561
rect 247876 318561 248196 325325
rect 247876 318325 247918 318561
rect 248154 318325 248196 318561
rect 247876 311561 248196 318325
rect 247876 311325 247918 311561
rect 248154 311325 248196 311561
rect 247876 304561 248196 311325
rect 247876 304325 247918 304561
rect 248154 304325 248196 304561
rect 247876 297561 248196 304325
rect 247876 297325 247918 297561
rect 248154 297325 248196 297561
rect 247876 290561 248196 297325
rect 247876 290325 247918 290561
rect 248154 290325 248196 290561
rect 247876 283561 248196 290325
rect 247876 283325 247918 283561
rect 248154 283325 248196 283561
rect 247876 276561 248196 283325
rect 247876 276325 247918 276561
rect 248154 276325 248196 276561
rect 247876 269561 248196 276325
rect 247876 269325 247918 269561
rect 248154 269325 248196 269561
rect 247876 262561 248196 269325
rect 247876 262325 247918 262561
rect 248154 262325 248196 262561
rect 247876 255561 248196 262325
rect 247876 255325 247918 255561
rect 248154 255325 248196 255561
rect 247876 248561 248196 255325
rect 247876 248325 247918 248561
rect 248154 248325 248196 248561
rect 247876 241561 248196 248325
rect 247876 241325 247918 241561
rect 248154 241325 248196 241561
rect 247876 234561 248196 241325
rect 247876 234325 247918 234561
rect 248154 234325 248196 234561
rect 247876 227561 248196 234325
rect 247876 227325 247918 227561
rect 248154 227325 248196 227561
rect 247876 220561 248196 227325
rect 247876 220325 247918 220561
rect 248154 220325 248196 220561
rect 247876 213561 248196 220325
rect 247876 213325 247918 213561
rect 248154 213325 248196 213561
rect 247876 206561 248196 213325
rect 247876 206325 247918 206561
rect 248154 206325 248196 206561
rect 247876 199561 248196 206325
rect 247876 199325 247918 199561
rect 248154 199325 248196 199561
rect 247876 192561 248196 199325
rect 247876 192325 247918 192561
rect 248154 192325 248196 192561
rect 247876 185561 248196 192325
rect 247876 185325 247918 185561
rect 248154 185325 248196 185561
rect 247876 178561 248196 185325
rect 247876 178325 247918 178561
rect 248154 178325 248196 178561
rect 247876 171561 248196 178325
rect 247876 171325 247918 171561
rect 248154 171325 248196 171561
rect 247876 164561 248196 171325
rect 247876 164325 247918 164561
rect 248154 164325 248196 164561
rect 247876 157561 248196 164325
rect 247876 157325 247918 157561
rect 248154 157325 248196 157561
rect 247876 150561 248196 157325
rect 247876 150325 247918 150561
rect 248154 150325 248196 150561
rect 247876 143561 248196 150325
rect 247876 143325 247918 143561
rect 248154 143325 248196 143561
rect 247876 136561 248196 143325
rect 247876 136325 247918 136561
rect 248154 136325 248196 136561
rect 247876 129561 248196 136325
rect 247876 129325 247918 129561
rect 248154 129325 248196 129561
rect 247876 122561 248196 129325
rect 247876 122325 247918 122561
rect 248154 122325 248196 122561
rect 247876 115561 248196 122325
rect 247876 115325 247918 115561
rect 248154 115325 248196 115561
rect 247876 108561 248196 115325
rect 247876 108325 247918 108561
rect 248154 108325 248196 108561
rect 247876 101561 248196 108325
rect 247876 101325 247918 101561
rect 248154 101325 248196 101561
rect 247876 94561 248196 101325
rect 247876 94325 247918 94561
rect 248154 94325 248196 94561
rect 247876 87561 248196 94325
rect 247876 87325 247918 87561
rect 248154 87325 248196 87561
rect 247876 80561 248196 87325
rect 247876 80325 247918 80561
rect 248154 80325 248196 80561
rect 247876 73561 248196 80325
rect 247876 73325 247918 73561
rect 248154 73325 248196 73561
rect 247876 66561 248196 73325
rect 247876 66325 247918 66561
rect 248154 66325 248196 66561
rect 247876 59561 248196 66325
rect 247876 59325 247918 59561
rect 248154 59325 248196 59561
rect 247876 52561 248196 59325
rect 247876 52325 247918 52561
rect 248154 52325 248196 52561
rect 247876 45561 248196 52325
rect 247876 45325 247918 45561
rect 248154 45325 248196 45561
rect 247876 38561 248196 45325
rect 247876 38325 247918 38561
rect 248154 38325 248196 38561
rect 247876 31561 248196 38325
rect 247876 31325 247918 31561
rect 248154 31325 248196 31561
rect 247876 24561 248196 31325
rect 247876 24325 247918 24561
rect 248154 24325 248196 24561
rect 247876 17561 248196 24325
rect 247876 17325 247918 17561
rect 248154 17325 248196 17561
rect 247876 10561 248196 17325
rect 247876 10325 247918 10561
rect 248154 10325 248196 10561
rect 247876 3561 248196 10325
rect 247876 3325 247918 3561
rect 248154 3325 248196 3561
rect 247876 -1706 248196 3325
rect 247876 -1942 247918 -1706
rect 248154 -1942 248196 -1706
rect 247876 -2026 248196 -1942
rect 247876 -2262 247918 -2026
rect 248154 -2262 248196 -2026
rect 247876 -2294 248196 -2262
rect 253144 705238 253464 706230
rect 253144 705002 253186 705238
rect 253422 705002 253464 705238
rect 253144 704918 253464 705002
rect 253144 704682 253186 704918
rect 253422 704682 253464 704918
rect 253144 695494 253464 704682
rect 253144 695258 253186 695494
rect 253422 695258 253464 695494
rect 253144 688494 253464 695258
rect 253144 688258 253186 688494
rect 253422 688258 253464 688494
rect 253144 681494 253464 688258
rect 253144 681258 253186 681494
rect 253422 681258 253464 681494
rect 253144 674494 253464 681258
rect 253144 674258 253186 674494
rect 253422 674258 253464 674494
rect 253144 667494 253464 674258
rect 253144 667258 253186 667494
rect 253422 667258 253464 667494
rect 253144 660494 253464 667258
rect 253144 660258 253186 660494
rect 253422 660258 253464 660494
rect 253144 653494 253464 660258
rect 253144 653258 253186 653494
rect 253422 653258 253464 653494
rect 253144 646494 253464 653258
rect 253144 646258 253186 646494
rect 253422 646258 253464 646494
rect 253144 639494 253464 646258
rect 253144 639258 253186 639494
rect 253422 639258 253464 639494
rect 253144 632494 253464 639258
rect 253144 632258 253186 632494
rect 253422 632258 253464 632494
rect 253144 625494 253464 632258
rect 253144 625258 253186 625494
rect 253422 625258 253464 625494
rect 253144 618494 253464 625258
rect 253144 618258 253186 618494
rect 253422 618258 253464 618494
rect 253144 611494 253464 618258
rect 253144 611258 253186 611494
rect 253422 611258 253464 611494
rect 253144 604494 253464 611258
rect 253144 604258 253186 604494
rect 253422 604258 253464 604494
rect 253144 597494 253464 604258
rect 253144 597258 253186 597494
rect 253422 597258 253464 597494
rect 253144 590494 253464 597258
rect 253144 590258 253186 590494
rect 253422 590258 253464 590494
rect 253144 583494 253464 590258
rect 253144 583258 253186 583494
rect 253422 583258 253464 583494
rect 253144 576494 253464 583258
rect 253144 576258 253186 576494
rect 253422 576258 253464 576494
rect 253144 569494 253464 576258
rect 253144 569258 253186 569494
rect 253422 569258 253464 569494
rect 253144 562494 253464 569258
rect 253144 562258 253186 562494
rect 253422 562258 253464 562494
rect 253144 555494 253464 562258
rect 253144 555258 253186 555494
rect 253422 555258 253464 555494
rect 253144 548494 253464 555258
rect 253144 548258 253186 548494
rect 253422 548258 253464 548494
rect 253144 541494 253464 548258
rect 253144 541258 253186 541494
rect 253422 541258 253464 541494
rect 253144 534494 253464 541258
rect 253144 534258 253186 534494
rect 253422 534258 253464 534494
rect 253144 527494 253464 534258
rect 253144 527258 253186 527494
rect 253422 527258 253464 527494
rect 253144 520494 253464 527258
rect 253144 520258 253186 520494
rect 253422 520258 253464 520494
rect 253144 513494 253464 520258
rect 253144 513258 253186 513494
rect 253422 513258 253464 513494
rect 253144 506494 253464 513258
rect 253144 506258 253186 506494
rect 253422 506258 253464 506494
rect 253144 499494 253464 506258
rect 253144 499258 253186 499494
rect 253422 499258 253464 499494
rect 253144 492494 253464 499258
rect 253144 492258 253186 492494
rect 253422 492258 253464 492494
rect 253144 485494 253464 492258
rect 253144 485258 253186 485494
rect 253422 485258 253464 485494
rect 253144 478494 253464 485258
rect 253144 478258 253186 478494
rect 253422 478258 253464 478494
rect 253144 471494 253464 478258
rect 253144 471258 253186 471494
rect 253422 471258 253464 471494
rect 253144 464494 253464 471258
rect 253144 464258 253186 464494
rect 253422 464258 253464 464494
rect 253144 457494 253464 464258
rect 253144 457258 253186 457494
rect 253422 457258 253464 457494
rect 253144 450494 253464 457258
rect 253144 450258 253186 450494
rect 253422 450258 253464 450494
rect 253144 443494 253464 450258
rect 253144 443258 253186 443494
rect 253422 443258 253464 443494
rect 253144 436494 253464 443258
rect 253144 436258 253186 436494
rect 253422 436258 253464 436494
rect 253144 429494 253464 436258
rect 253144 429258 253186 429494
rect 253422 429258 253464 429494
rect 253144 422494 253464 429258
rect 253144 422258 253186 422494
rect 253422 422258 253464 422494
rect 253144 415494 253464 422258
rect 253144 415258 253186 415494
rect 253422 415258 253464 415494
rect 253144 408494 253464 415258
rect 253144 408258 253186 408494
rect 253422 408258 253464 408494
rect 253144 401494 253464 408258
rect 253144 401258 253186 401494
rect 253422 401258 253464 401494
rect 253144 394494 253464 401258
rect 253144 394258 253186 394494
rect 253422 394258 253464 394494
rect 253144 387494 253464 394258
rect 253144 387258 253186 387494
rect 253422 387258 253464 387494
rect 253144 380494 253464 387258
rect 253144 380258 253186 380494
rect 253422 380258 253464 380494
rect 253144 373494 253464 380258
rect 253144 373258 253186 373494
rect 253422 373258 253464 373494
rect 253144 366494 253464 373258
rect 253144 366258 253186 366494
rect 253422 366258 253464 366494
rect 253144 359494 253464 366258
rect 253144 359258 253186 359494
rect 253422 359258 253464 359494
rect 253144 352494 253464 359258
rect 253144 352258 253186 352494
rect 253422 352258 253464 352494
rect 253144 345494 253464 352258
rect 253144 345258 253186 345494
rect 253422 345258 253464 345494
rect 253144 338494 253464 345258
rect 253144 338258 253186 338494
rect 253422 338258 253464 338494
rect 253144 331494 253464 338258
rect 253144 331258 253186 331494
rect 253422 331258 253464 331494
rect 253144 324494 253464 331258
rect 253144 324258 253186 324494
rect 253422 324258 253464 324494
rect 253144 317494 253464 324258
rect 253144 317258 253186 317494
rect 253422 317258 253464 317494
rect 253144 310494 253464 317258
rect 253144 310258 253186 310494
rect 253422 310258 253464 310494
rect 253144 303494 253464 310258
rect 253144 303258 253186 303494
rect 253422 303258 253464 303494
rect 253144 296494 253464 303258
rect 253144 296258 253186 296494
rect 253422 296258 253464 296494
rect 253144 289494 253464 296258
rect 253144 289258 253186 289494
rect 253422 289258 253464 289494
rect 253144 282494 253464 289258
rect 253144 282258 253186 282494
rect 253422 282258 253464 282494
rect 253144 275494 253464 282258
rect 253144 275258 253186 275494
rect 253422 275258 253464 275494
rect 253144 268494 253464 275258
rect 253144 268258 253186 268494
rect 253422 268258 253464 268494
rect 253144 261494 253464 268258
rect 253144 261258 253186 261494
rect 253422 261258 253464 261494
rect 253144 254494 253464 261258
rect 253144 254258 253186 254494
rect 253422 254258 253464 254494
rect 253144 247494 253464 254258
rect 253144 247258 253186 247494
rect 253422 247258 253464 247494
rect 253144 240494 253464 247258
rect 253144 240258 253186 240494
rect 253422 240258 253464 240494
rect 253144 233494 253464 240258
rect 253144 233258 253186 233494
rect 253422 233258 253464 233494
rect 253144 226494 253464 233258
rect 253144 226258 253186 226494
rect 253422 226258 253464 226494
rect 253144 219494 253464 226258
rect 253144 219258 253186 219494
rect 253422 219258 253464 219494
rect 253144 212494 253464 219258
rect 253144 212258 253186 212494
rect 253422 212258 253464 212494
rect 253144 205494 253464 212258
rect 253144 205258 253186 205494
rect 253422 205258 253464 205494
rect 253144 198494 253464 205258
rect 253144 198258 253186 198494
rect 253422 198258 253464 198494
rect 253144 191494 253464 198258
rect 253144 191258 253186 191494
rect 253422 191258 253464 191494
rect 253144 184494 253464 191258
rect 253144 184258 253186 184494
rect 253422 184258 253464 184494
rect 253144 177494 253464 184258
rect 253144 177258 253186 177494
rect 253422 177258 253464 177494
rect 253144 170494 253464 177258
rect 253144 170258 253186 170494
rect 253422 170258 253464 170494
rect 253144 163494 253464 170258
rect 253144 163258 253186 163494
rect 253422 163258 253464 163494
rect 253144 156494 253464 163258
rect 253144 156258 253186 156494
rect 253422 156258 253464 156494
rect 253144 149494 253464 156258
rect 253144 149258 253186 149494
rect 253422 149258 253464 149494
rect 253144 142494 253464 149258
rect 253144 142258 253186 142494
rect 253422 142258 253464 142494
rect 253144 135494 253464 142258
rect 253144 135258 253186 135494
rect 253422 135258 253464 135494
rect 253144 128494 253464 135258
rect 253144 128258 253186 128494
rect 253422 128258 253464 128494
rect 253144 121494 253464 128258
rect 253144 121258 253186 121494
rect 253422 121258 253464 121494
rect 253144 114494 253464 121258
rect 253144 114258 253186 114494
rect 253422 114258 253464 114494
rect 253144 107494 253464 114258
rect 253144 107258 253186 107494
rect 253422 107258 253464 107494
rect 253144 100494 253464 107258
rect 253144 100258 253186 100494
rect 253422 100258 253464 100494
rect 253144 93494 253464 100258
rect 253144 93258 253186 93494
rect 253422 93258 253464 93494
rect 253144 86494 253464 93258
rect 253144 86258 253186 86494
rect 253422 86258 253464 86494
rect 253144 79494 253464 86258
rect 253144 79258 253186 79494
rect 253422 79258 253464 79494
rect 253144 72494 253464 79258
rect 253144 72258 253186 72494
rect 253422 72258 253464 72494
rect 253144 65494 253464 72258
rect 253144 65258 253186 65494
rect 253422 65258 253464 65494
rect 253144 58494 253464 65258
rect 253144 58258 253186 58494
rect 253422 58258 253464 58494
rect 253144 51494 253464 58258
rect 253144 51258 253186 51494
rect 253422 51258 253464 51494
rect 253144 44494 253464 51258
rect 253144 44258 253186 44494
rect 253422 44258 253464 44494
rect 253144 37494 253464 44258
rect 253144 37258 253186 37494
rect 253422 37258 253464 37494
rect 253144 30494 253464 37258
rect 253144 30258 253186 30494
rect 253422 30258 253464 30494
rect 253144 23494 253464 30258
rect 253144 23258 253186 23494
rect 253422 23258 253464 23494
rect 253144 16494 253464 23258
rect 253144 16258 253186 16494
rect 253422 16258 253464 16494
rect 253144 9494 253464 16258
rect 253144 9258 253186 9494
rect 253422 9258 253464 9494
rect 253144 2494 253464 9258
rect 253144 2258 253186 2494
rect 253422 2258 253464 2494
rect 253144 -746 253464 2258
rect 253144 -982 253186 -746
rect 253422 -982 253464 -746
rect 253144 -1066 253464 -982
rect 253144 -1302 253186 -1066
rect 253422 -1302 253464 -1066
rect 253144 -2294 253464 -1302
rect 254876 706198 255196 706230
rect 254876 705962 254918 706198
rect 255154 705962 255196 706198
rect 254876 705878 255196 705962
rect 254876 705642 254918 705878
rect 255154 705642 255196 705878
rect 254876 696561 255196 705642
rect 254876 696325 254918 696561
rect 255154 696325 255196 696561
rect 254876 689561 255196 696325
rect 254876 689325 254918 689561
rect 255154 689325 255196 689561
rect 254876 682561 255196 689325
rect 254876 682325 254918 682561
rect 255154 682325 255196 682561
rect 254876 675561 255196 682325
rect 254876 675325 254918 675561
rect 255154 675325 255196 675561
rect 254876 668561 255196 675325
rect 254876 668325 254918 668561
rect 255154 668325 255196 668561
rect 254876 661561 255196 668325
rect 254876 661325 254918 661561
rect 255154 661325 255196 661561
rect 254876 654561 255196 661325
rect 254876 654325 254918 654561
rect 255154 654325 255196 654561
rect 254876 647561 255196 654325
rect 254876 647325 254918 647561
rect 255154 647325 255196 647561
rect 254876 640561 255196 647325
rect 254876 640325 254918 640561
rect 255154 640325 255196 640561
rect 254876 633561 255196 640325
rect 254876 633325 254918 633561
rect 255154 633325 255196 633561
rect 254876 626561 255196 633325
rect 254876 626325 254918 626561
rect 255154 626325 255196 626561
rect 254876 619561 255196 626325
rect 254876 619325 254918 619561
rect 255154 619325 255196 619561
rect 254876 612561 255196 619325
rect 254876 612325 254918 612561
rect 255154 612325 255196 612561
rect 254876 605561 255196 612325
rect 254876 605325 254918 605561
rect 255154 605325 255196 605561
rect 254876 598561 255196 605325
rect 254876 598325 254918 598561
rect 255154 598325 255196 598561
rect 254876 591561 255196 598325
rect 254876 591325 254918 591561
rect 255154 591325 255196 591561
rect 254876 584561 255196 591325
rect 254876 584325 254918 584561
rect 255154 584325 255196 584561
rect 254876 577561 255196 584325
rect 254876 577325 254918 577561
rect 255154 577325 255196 577561
rect 254876 570561 255196 577325
rect 254876 570325 254918 570561
rect 255154 570325 255196 570561
rect 254876 563561 255196 570325
rect 254876 563325 254918 563561
rect 255154 563325 255196 563561
rect 254876 556561 255196 563325
rect 254876 556325 254918 556561
rect 255154 556325 255196 556561
rect 254876 549561 255196 556325
rect 254876 549325 254918 549561
rect 255154 549325 255196 549561
rect 254876 542561 255196 549325
rect 254876 542325 254918 542561
rect 255154 542325 255196 542561
rect 254876 535561 255196 542325
rect 254876 535325 254918 535561
rect 255154 535325 255196 535561
rect 254876 528561 255196 535325
rect 254876 528325 254918 528561
rect 255154 528325 255196 528561
rect 254876 521561 255196 528325
rect 254876 521325 254918 521561
rect 255154 521325 255196 521561
rect 254876 514561 255196 521325
rect 254876 514325 254918 514561
rect 255154 514325 255196 514561
rect 254876 507561 255196 514325
rect 254876 507325 254918 507561
rect 255154 507325 255196 507561
rect 254876 500561 255196 507325
rect 254876 500325 254918 500561
rect 255154 500325 255196 500561
rect 254876 493561 255196 500325
rect 254876 493325 254918 493561
rect 255154 493325 255196 493561
rect 254876 486561 255196 493325
rect 254876 486325 254918 486561
rect 255154 486325 255196 486561
rect 254876 479561 255196 486325
rect 254876 479325 254918 479561
rect 255154 479325 255196 479561
rect 254876 472561 255196 479325
rect 254876 472325 254918 472561
rect 255154 472325 255196 472561
rect 254876 465561 255196 472325
rect 254876 465325 254918 465561
rect 255154 465325 255196 465561
rect 254876 458561 255196 465325
rect 254876 458325 254918 458561
rect 255154 458325 255196 458561
rect 254876 451561 255196 458325
rect 254876 451325 254918 451561
rect 255154 451325 255196 451561
rect 254876 444561 255196 451325
rect 254876 444325 254918 444561
rect 255154 444325 255196 444561
rect 254876 437561 255196 444325
rect 254876 437325 254918 437561
rect 255154 437325 255196 437561
rect 254876 430561 255196 437325
rect 254876 430325 254918 430561
rect 255154 430325 255196 430561
rect 254876 423561 255196 430325
rect 254876 423325 254918 423561
rect 255154 423325 255196 423561
rect 254876 416561 255196 423325
rect 254876 416325 254918 416561
rect 255154 416325 255196 416561
rect 254876 409561 255196 416325
rect 254876 409325 254918 409561
rect 255154 409325 255196 409561
rect 254876 402561 255196 409325
rect 254876 402325 254918 402561
rect 255154 402325 255196 402561
rect 254876 395561 255196 402325
rect 254876 395325 254918 395561
rect 255154 395325 255196 395561
rect 254876 388561 255196 395325
rect 254876 388325 254918 388561
rect 255154 388325 255196 388561
rect 254876 381561 255196 388325
rect 254876 381325 254918 381561
rect 255154 381325 255196 381561
rect 254876 374561 255196 381325
rect 254876 374325 254918 374561
rect 255154 374325 255196 374561
rect 254876 367561 255196 374325
rect 254876 367325 254918 367561
rect 255154 367325 255196 367561
rect 254876 360561 255196 367325
rect 254876 360325 254918 360561
rect 255154 360325 255196 360561
rect 254876 353561 255196 360325
rect 254876 353325 254918 353561
rect 255154 353325 255196 353561
rect 254876 346561 255196 353325
rect 254876 346325 254918 346561
rect 255154 346325 255196 346561
rect 254876 339561 255196 346325
rect 254876 339325 254918 339561
rect 255154 339325 255196 339561
rect 254876 332561 255196 339325
rect 254876 332325 254918 332561
rect 255154 332325 255196 332561
rect 254876 325561 255196 332325
rect 254876 325325 254918 325561
rect 255154 325325 255196 325561
rect 254876 318561 255196 325325
rect 254876 318325 254918 318561
rect 255154 318325 255196 318561
rect 254876 311561 255196 318325
rect 254876 311325 254918 311561
rect 255154 311325 255196 311561
rect 254876 304561 255196 311325
rect 254876 304325 254918 304561
rect 255154 304325 255196 304561
rect 254876 297561 255196 304325
rect 254876 297325 254918 297561
rect 255154 297325 255196 297561
rect 254876 290561 255196 297325
rect 254876 290325 254918 290561
rect 255154 290325 255196 290561
rect 254876 283561 255196 290325
rect 254876 283325 254918 283561
rect 255154 283325 255196 283561
rect 254876 276561 255196 283325
rect 254876 276325 254918 276561
rect 255154 276325 255196 276561
rect 254876 269561 255196 276325
rect 254876 269325 254918 269561
rect 255154 269325 255196 269561
rect 254876 262561 255196 269325
rect 254876 262325 254918 262561
rect 255154 262325 255196 262561
rect 254876 255561 255196 262325
rect 254876 255325 254918 255561
rect 255154 255325 255196 255561
rect 254876 248561 255196 255325
rect 254876 248325 254918 248561
rect 255154 248325 255196 248561
rect 254876 241561 255196 248325
rect 254876 241325 254918 241561
rect 255154 241325 255196 241561
rect 254876 234561 255196 241325
rect 254876 234325 254918 234561
rect 255154 234325 255196 234561
rect 254876 227561 255196 234325
rect 254876 227325 254918 227561
rect 255154 227325 255196 227561
rect 254876 220561 255196 227325
rect 254876 220325 254918 220561
rect 255154 220325 255196 220561
rect 254876 213561 255196 220325
rect 254876 213325 254918 213561
rect 255154 213325 255196 213561
rect 254876 206561 255196 213325
rect 254876 206325 254918 206561
rect 255154 206325 255196 206561
rect 254876 199561 255196 206325
rect 254876 199325 254918 199561
rect 255154 199325 255196 199561
rect 254876 192561 255196 199325
rect 254876 192325 254918 192561
rect 255154 192325 255196 192561
rect 254876 185561 255196 192325
rect 254876 185325 254918 185561
rect 255154 185325 255196 185561
rect 254876 178561 255196 185325
rect 254876 178325 254918 178561
rect 255154 178325 255196 178561
rect 254876 171561 255196 178325
rect 254876 171325 254918 171561
rect 255154 171325 255196 171561
rect 254876 164561 255196 171325
rect 254876 164325 254918 164561
rect 255154 164325 255196 164561
rect 254876 157561 255196 164325
rect 254876 157325 254918 157561
rect 255154 157325 255196 157561
rect 254876 150561 255196 157325
rect 254876 150325 254918 150561
rect 255154 150325 255196 150561
rect 254876 143561 255196 150325
rect 254876 143325 254918 143561
rect 255154 143325 255196 143561
rect 254876 136561 255196 143325
rect 254876 136325 254918 136561
rect 255154 136325 255196 136561
rect 254876 129561 255196 136325
rect 254876 129325 254918 129561
rect 255154 129325 255196 129561
rect 254876 122561 255196 129325
rect 254876 122325 254918 122561
rect 255154 122325 255196 122561
rect 254876 115561 255196 122325
rect 254876 115325 254918 115561
rect 255154 115325 255196 115561
rect 254876 108561 255196 115325
rect 254876 108325 254918 108561
rect 255154 108325 255196 108561
rect 254876 101561 255196 108325
rect 254876 101325 254918 101561
rect 255154 101325 255196 101561
rect 254876 94561 255196 101325
rect 254876 94325 254918 94561
rect 255154 94325 255196 94561
rect 254876 87561 255196 94325
rect 254876 87325 254918 87561
rect 255154 87325 255196 87561
rect 254876 80561 255196 87325
rect 254876 80325 254918 80561
rect 255154 80325 255196 80561
rect 254876 73561 255196 80325
rect 254876 73325 254918 73561
rect 255154 73325 255196 73561
rect 254876 66561 255196 73325
rect 254876 66325 254918 66561
rect 255154 66325 255196 66561
rect 254876 59561 255196 66325
rect 254876 59325 254918 59561
rect 255154 59325 255196 59561
rect 254876 52561 255196 59325
rect 254876 52325 254918 52561
rect 255154 52325 255196 52561
rect 254876 45561 255196 52325
rect 254876 45325 254918 45561
rect 255154 45325 255196 45561
rect 254876 38561 255196 45325
rect 254876 38325 254918 38561
rect 255154 38325 255196 38561
rect 254876 31561 255196 38325
rect 254876 31325 254918 31561
rect 255154 31325 255196 31561
rect 254876 24561 255196 31325
rect 254876 24325 254918 24561
rect 255154 24325 255196 24561
rect 254876 17561 255196 24325
rect 254876 17325 254918 17561
rect 255154 17325 255196 17561
rect 254876 10561 255196 17325
rect 254876 10325 254918 10561
rect 255154 10325 255196 10561
rect 254876 3561 255196 10325
rect 254876 3325 254918 3561
rect 255154 3325 255196 3561
rect 254876 -1706 255196 3325
rect 254876 -1942 254918 -1706
rect 255154 -1942 255196 -1706
rect 254876 -2026 255196 -1942
rect 254876 -2262 254918 -2026
rect 255154 -2262 255196 -2026
rect 254876 -2294 255196 -2262
rect 260144 705238 260464 706230
rect 260144 705002 260186 705238
rect 260422 705002 260464 705238
rect 260144 704918 260464 705002
rect 260144 704682 260186 704918
rect 260422 704682 260464 704918
rect 260144 695494 260464 704682
rect 260144 695258 260186 695494
rect 260422 695258 260464 695494
rect 260144 688494 260464 695258
rect 260144 688258 260186 688494
rect 260422 688258 260464 688494
rect 260144 681494 260464 688258
rect 260144 681258 260186 681494
rect 260422 681258 260464 681494
rect 260144 674494 260464 681258
rect 260144 674258 260186 674494
rect 260422 674258 260464 674494
rect 260144 667494 260464 674258
rect 260144 667258 260186 667494
rect 260422 667258 260464 667494
rect 260144 660494 260464 667258
rect 260144 660258 260186 660494
rect 260422 660258 260464 660494
rect 260144 653494 260464 660258
rect 260144 653258 260186 653494
rect 260422 653258 260464 653494
rect 260144 646494 260464 653258
rect 260144 646258 260186 646494
rect 260422 646258 260464 646494
rect 260144 639494 260464 646258
rect 260144 639258 260186 639494
rect 260422 639258 260464 639494
rect 260144 632494 260464 639258
rect 260144 632258 260186 632494
rect 260422 632258 260464 632494
rect 260144 625494 260464 632258
rect 260144 625258 260186 625494
rect 260422 625258 260464 625494
rect 260144 618494 260464 625258
rect 260144 618258 260186 618494
rect 260422 618258 260464 618494
rect 260144 611494 260464 618258
rect 260144 611258 260186 611494
rect 260422 611258 260464 611494
rect 260144 604494 260464 611258
rect 260144 604258 260186 604494
rect 260422 604258 260464 604494
rect 260144 597494 260464 604258
rect 260144 597258 260186 597494
rect 260422 597258 260464 597494
rect 260144 590494 260464 597258
rect 260144 590258 260186 590494
rect 260422 590258 260464 590494
rect 260144 583494 260464 590258
rect 260144 583258 260186 583494
rect 260422 583258 260464 583494
rect 260144 576494 260464 583258
rect 260144 576258 260186 576494
rect 260422 576258 260464 576494
rect 260144 569494 260464 576258
rect 260144 569258 260186 569494
rect 260422 569258 260464 569494
rect 260144 562494 260464 569258
rect 260144 562258 260186 562494
rect 260422 562258 260464 562494
rect 260144 555494 260464 562258
rect 260144 555258 260186 555494
rect 260422 555258 260464 555494
rect 260144 548494 260464 555258
rect 260144 548258 260186 548494
rect 260422 548258 260464 548494
rect 260144 541494 260464 548258
rect 260144 541258 260186 541494
rect 260422 541258 260464 541494
rect 260144 534494 260464 541258
rect 260144 534258 260186 534494
rect 260422 534258 260464 534494
rect 260144 527494 260464 534258
rect 260144 527258 260186 527494
rect 260422 527258 260464 527494
rect 260144 520494 260464 527258
rect 260144 520258 260186 520494
rect 260422 520258 260464 520494
rect 260144 513494 260464 520258
rect 260144 513258 260186 513494
rect 260422 513258 260464 513494
rect 260144 506494 260464 513258
rect 260144 506258 260186 506494
rect 260422 506258 260464 506494
rect 260144 499494 260464 506258
rect 260144 499258 260186 499494
rect 260422 499258 260464 499494
rect 260144 492494 260464 499258
rect 260144 492258 260186 492494
rect 260422 492258 260464 492494
rect 260144 485494 260464 492258
rect 260144 485258 260186 485494
rect 260422 485258 260464 485494
rect 260144 478494 260464 485258
rect 260144 478258 260186 478494
rect 260422 478258 260464 478494
rect 260144 471494 260464 478258
rect 260144 471258 260186 471494
rect 260422 471258 260464 471494
rect 260144 464494 260464 471258
rect 260144 464258 260186 464494
rect 260422 464258 260464 464494
rect 260144 457494 260464 464258
rect 260144 457258 260186 457494
rect 260422 457258 260464 457494
rect 260144 450494 260464 457258
rect 260144 450258 260186 450494
rect 260422 450258 260464 450494
rect 260144 443494 260464 450258
rect 260144 443258 260186 443494
rect 260422 443258 260464 443494
rect 260144 436494 260464 443258
rect 260144 436258 260186 436494
rect 260422 436258 260464 436494
rect 260144 429494 260464 436258
rect 260144 429258 260186 429494
rect 260422 429258 260464 429494
rect 260144 422494 260464 429258
rect 260144 422258 260186 422494
rect 260422 422258 260464 422494
rect 260144 415494 260464 422258
rect 260144 415258 260186 415494
rect 260422 415258 260464 415494
rect 260144 408494 260464 415258
rect 260144 408258 260186 408494
rect 260422 408258 260464 408494
rect 260144 401494 260464 408258
rect 260144 401258 260186 401494
rect 260422 401258 260464 401494
rect 260144 394494 260464 401258
rect 260144 394258 260186 394494
rect 260422 394258 260464 394494
rect 260144 387494 260464 394258
rect 260144 387258 260186 387494
rect 260422 387258 260464 387494
rect 260144 380494 260464 387258
rect 260144 380258 260186 380494
rect 260422 380258 260464 380494
rect 260144 373494 260464 380258
rect 260144 373258 260186 373494
rect 260422 373258 260464 373494
rect 260144 366494 260464 373258
rect 260144 366258 260186 366494
rect 260422 366258 260464 366494
rect 260144 359494 260464 366258
rect 260144 359258 260186 359494
rect 260422 359258 260464 359494
rect 260144 352494 260464 359258
rect 260144 352258 260186 352494
rect 260422 352258 260464 352494
rect 260144 345494 260464 352258
rect 260144 345258 260186 345494
rect 260422 345258 260464 345494
rect 260144 338494 260464 345258
rect 260144 338258 260186 338494
rect 260422 338258 260464 338494
rect 260144 331494 260464 338258
rect 260144 331258 260186 331494
rect 260422 331258 260464 331494
rect 260144 324494 260464 331258
rect 260144 324258 260186 324494
rect 260422 324258 260464 324494
rect 260144 317494 260464 324258
rect 260144 317258 260186 317494
rect 260422 317258 260464 317494
rect 260144 310494 260464 317258
rect 260144 310258 260186 310494
rect 260422 310258 260464 310494
rect 260144 303494 260464 310258
rect 260144 303258 260186 303494
rect 260422 303258 260464 303494
rect 260144 296494 260464 303258
rect 260144 296258 260186 296494
rect 260422 296258 260464 296494
rect 260144 289494 260464 296258
rect 260144 289258 260186 289494
rect 260422 289258 260464 289494
rect 260144 282494 260464 289258
rect 260144 282258 260186 282494
rect 260422 282258 260464 282494
rect 260144 275494 260464 282258
rect 260144 275258 260186 275494
rect 260422 275258 260464 275494
rect 260144 268494 260464 275258
rect 260144 268258 260186 268494
rect 260422 268258 260464 268494
rect 260144 261494 260464 268258
rect 260144 261258 260186 261494
rect 260422 261258 260464 261494
rect 260144 254494 260464 261258
rect 260144 254258 260186 254494
rect 260422 254258 260464 254494
rect 260144 247494 260464 254258
rect 260144 247258 260186 247494
rect 260422 247258 260464 247494
rect 260144 240494 260464 247258
rect 260144 240258 260186 240494
rect 260422 240258 260464 240494
rect 260144 233494 260464 240258
rect 260144 233258 260186 233494
rect 260422 233258 260464 233494
rect 260144 226494 260464 233258
rect 260144 226258 260186 226494
rect 260422 226258 260464 226494
rect 260144 219494 260464 226258
rect 260144 219258 260186 219494
rect 260422 219258 260464 219494
rect 260144 212494 260464 219258
rect 260144 212258 260186 212494
rect 260422 212258 260464 212494
rect 260144 205494 260464 212258
rect 260144 205258 260186 205494
rect 260422 205258 260464 205494
rect 260144 198494 260464 205258
rect 260144 198258 260186 198494
rect 260422 198258 260464 198494
rect 260144 191494 260464 198258
rect 260144 191258 260186 191494
rect 260422 191258 260464 191494
rect 260144 184494 260464 191258
rect 260144 184258 260186 184494
rect 260422 184258 260464 184494
rect 260144 177494 260464 184258
rect 260144 177258 260186 177494
rect 260422 177258 260464 177494
rect 260144 170494 260464 177258
rect 260144 170258 260186 170494
rect 260422 170258 260464 170494
rect 260144 163494 260464 170258
rect 260144 163258 260186 163494
rect 260422 163258 260464 163494
rect 260144 156494 260464 163258
rect 260144 156258 260186 156494
rect 260422 156258 260464 156494
rect 260144 149494 260464 156258
rect 260144 149258 260186 149494
rect 260422 149258 260464 149494
rect 260144 142494 260464 149258
rect 260144 142258 260186 142494
rect 260422 142258 260464 142494
rect 260144 135494 260464 142258
rect 260144 135258 260186 135494
rect 260422 135258 260464 135494
rect 260144 128494 260464 135258
rect 260144 128258 260186 128494
rect 260422 128258 260464 128494
rect 260144 121494 260464 128258
rect 260144 121258 260186 121494
rect 260422 121258 260464 121494
rect 260144 114494 260464 121258
rect 260144 114258 260186 114494
rect 260422 114258 260464 114494
rect 260144 107494 260464 114258
rect 260144 107258 260186 107494
rect 260422 107258 260464 107494
rect 260144 100494 260464 107258
rect 260144 100258 260186 100494
rect 260422 100258 260464 100494
rect 260144 93494 260464 100258
rect 260144 93258 260186 93494
rect 260422 93258 260464 93494
rect 260144 86494 260464 93258
rect 260144 86258 260186 86494
rect 260422 86258 260464 86494
rect 260144 79494 260464 86258
rect 260144 79258 260186 79494
rect 260422 79258 260464 79494
rect 260144 72494 260464 79258
rect 260144 72258 260186 72494
rect 260422 72258 260464 72494
rect 260144 65494 260464 72258
rect 260144 65258 260186 65494
rect 260422 65258 260464 65494
rect 260144 58494 260464 65258
rect 260144 58258 260186 58494
rect 260422 58258 260464 58494
rect 260144 51494 260464 58258
rect 260144 51258 260186 51494
rect 260422 51258 260464 51494
rect 260144 44494 260464 51258
rect 260144 44258 260186 44494
rect 260422 44258 260464 44494
rect 260144 37494 260464 44258
rect 260144 37258 260186 37494
rect 260422 37258 260464 37494
rect 260144 30494 260464 37258
rect 260144 30258 260186 30494
rect 260422 30258 260464 30494
rect 260144 23494 260464 30258
rect 260144 23258 260186 23494
rect 260422 23258 260464 23494
rect 260144 16494 260464 23258
rect 260144 16258 260186 16494
rect 260422 16258 260464 16494
rect 260144 9494 260464 16258
rect 260144 9258 260186 9494
rect 260422 9258 260464 9494
rect 260144 2494 260464 9258
rect 260144 2258 260186 2494
rect 260422 2258 260464 2494
rect 260144 -746 260464 2258
rect 260144 -982 260186 -746
rect 260422 -982 260464 -746
rect 260144 -1066 260464 -982
rect 260144 -1302 260186 -1066
rect 260422 -1302 260464 -1066
rect 260144 -2294 260464 -1302
rect 261876 706198 262196 706230
rect 261876 705962 261918 706198
rect 262154 705962 262196 706198
rect 261876 705878 262196 705962
rect 261876 705642 261918 705878
rect 262154 705642 262196 705878
rect 261876 696561 262196 705642
rect 261876 696325 261918 696561
rect 262154 696325 262196 696561
rect 261876 689561 262196 696325
rect 261876 689325 261918 689561
rect 262154 689325 262196 689561
rect 261876 682561 262196 689325
rect 261876 682325 261918 682561
rect 262154 682325 262196 682561
rect 261876 675561 262196 682325
rect 261876 675325 261918 675561
rect 262154 675325 262196 675561
rect 261876 668561 262196 675325
rect 261876 668325 261918 668561
rect 262154 668325 262196 668561
rect 261876 661561 262196 668325
rect 261876 661325 261918 661561
rect 262154 661325 262196 661561
rect 261876 654561 262196 661325
rect 261876 654325 261918 654561
rect 262154 654325 262196 654561
rect 261876 647561 262196 654325
rect 261876 647325 261918 647561
rect 262154 647325 262196 647561
rect 261876 640561 262196 647325
rect 261876 640325 261918 640561
rect 262154 640325 262196 640561
rect 261876 633561 262196 640325
rect 261876 633325 261918 633561
rect 262154 633325 262196 633561
rect 261876 626561 262196 633325
rect 261876 626325 261918 626561
rect 262154 626325 262196 626561
rect 261876 619561 262196 626325
rect 261876 619325 261918 619561
rect 262154 619325 262196 619561
rect 261876 612561 262196 619325
rect 261876 612325 261918 612561
rect 262154 612325 262196 612561
rect 261876 605561 262196 612325
rect 261876 605325 261918 605561
rect 262154 605325 262196 605561
rect 261876 598561 262196 605325
rect 261876 598325 261918 598561
rect 262154 598325 262196 598561
rect 261876 591561 262196 598325
rect 261876 591325 261918 591561
rect 262154 591325 262196 591561
rect 261876 584561 262196 591325
rect 261876 584325 261918 584561
rect 262154 584325 262196 584561
rect 261876 577561 262196 584325
rect 261876 577325 261918 577561
rect 262154 577325 262196 577561
rect 261876 570561 262196 577325
rect 261876 570325 261918 570561
rect 262154 570325 262196 570561
rect 261876 563561 262196 570325
rect 261876 563325 261918 563561
rect 262154 563325 262196 563561
rect 261876 556561 262196 563325
rect 261876 556325 261918 556561
rect 262154 556325 262196 556561
rect 261876 549561 262196 556325
rect 261876 549325 261918 549561
rect 262154 549325 262196 549561
rect 261876 542561 262196 549325
rect 261876 542325 261918 542561
rect 262154 542325 262196 542561
rect 261876 535561 262196 542325
rect 261876 535325 261918 535561
rect 262154 535325 262196 535561
rect 261876 528561 262196 535325
rect 261876 528325 261918 528561
rect 262154 528325 262196 528561
rect 261876 521561 262196 528325
rect 261876 521325 261918 521561
rect 262154 521325 262196 521561
rect 261876 514561 262196 521325
rect 261876 514325 261918 514561
rect 262154 514325 262196 514561
rect 261876 507561 262196 514325
rect 261876 507325 261918 507561
rect 262154 507325 262196 507561
rect 261876 500561 262196 507325
rect 261876 500325 261918 500561
rect 262154 500325 262196 500561
rect 261876 493561 262196 500325
rect 261876 493325 261918 493561
rect 262154 493325 262196 493561
rect 261876 486561 262196 493325
rect 261876 486325 261918 486561
rect 262154 486325 262196 486561
rect 261876 479561 262196 486325
rect 261876 479325 261918 479561
rect 262154 479325 262196 479561
rect 261876 472561 262196 479325
rect 261876 472325 261918 472561
rect 262154 472325 262196 472561
rect 261876 465561 262196 472325
rect 261876 465325 261918 465561
rect 262154 465325 262196 465561
rect 261876 458561 262196 465325
rect 261876 458325 261918 458561
rect 262154 458325 262196 458561
rect 261876 451561 262196 458325
rect 261876 451325 261918 451561
rect 262154 451325 262196 451561
rect 261876 444561 262196 451325
rect 261876 444325 261918 444561
rect 262154 444325 262196 444561
rect 261876 437561 262196 444325
rect 261876 437325 261918 437561
rect 262154 437325 262196 437561
rect 261876 430561 262196 437325
rect 261876 430325 261918 430561
rect 262154 430325 262196 430561
rect 261876 423561 262196 430325
rect 261876 423325 261918 423561
rect 262154 423325 262196 423561
rect 261876 416561 262196 423325
rect 261876 416325 261918 416561
rect 262154 416325 262196 416561
rect 261876 409561 262196 416325
rect 261876 409325 261918 409561
rect 262154 409325 262196 409561
rect 261876 402561 262196 409325
rect 261876 402325 261918 402561
rect 262154 402325 262196 402561
rect 261876 395561 262196 402325
rect 261876 395325 261918 395561
rect 262154 395325 262196 395561
rect 261876 388561 262196 395325
rect 261876 388325 261918 388561
rect 262154 388325 262196 388561
rect 261876 381561 262196 388325
rect 261876 381325 261918 381561
rect 262154 381325 262196 381561
rect 261876 374561 262196 381325
rect 261876 374325 261918 374561
rect 262154 374325 262196 374561
rect 261876 367561 262196 374325
rect 261876 367325 261918 367561
rect 262154 367325 262196 367561
rect 261876 360561 262196 367325
rect 261876 360325 261918 360561
rect 262154 360325 262196 360561
rect 261876 353561 262196 360325
rect 261876 353325 261918 353561
rect 262154 353325 262196 353561
rect 261876 346561 262196 353325
rect 261876 346325 261918 346561
rect 262154 346325 262196 346561
rect 261876 339561 262196 346325
rect 261876 339325 261918 339561
rect 262154 339325 262196 339561
rect 261876 332561 262196 339325
rect 261876 332325 261918 332561
rect 262154 332325 262196 332561
rect 261876 325561 262196 332325
rect 261876 325325 261918 325561
rect 262154 325325 262196 325561
rect 261876 318561 262196 325325
rect 261876 318325 261918 318561
rect 262154 318325 262196 318561
rect 261876 311561 262196 318325
rect 261876 311325 261918 311561
rect 262154 311325 262196 311561
rect 261876 304561 262196 311325
rect 261876 304325 261918 304561
rect 262154 304325 262196 304561
rect 261876 297561 262196 304325
rect 261876 297325 261918 297561
rect 262154 297325 262196 297561
rect 261876 290561 262196 297325
rect 261876 290325 261918 290561
rect 262154 290325 262196 290561
rect 261876 283561 262196 290325
rect 261876 283325 261918 283561
rect 262154 283325 262196 283561
rect 261876 276561 262196 283325
rect 261876 276325 261918 276561
rect 262154 276325 262196 276561
rect 261876 269561 262196 276325
rect 261876 269325 261918 269561
rect 262154 269325 262196 269561
rect 261876 262561 262196 269325
rect 261876 262325 261918 262561
rect 262154 262325 262196 262561
rect 261876 255561 262196 262325
rect 261876 255325 261918 255561
rect 262154 255325 262196 255561
rect 261876 248561 262196 255325
rect 261876 248325 261918 248561
rect 262154 248325 262196 248561
rect 261876 241561 262196 248325
rect 261876 241325 261918 241561
rect 262154 241325 262196 241561
rect 261876 234561 262196 241325
rect 261876 234325 261918 234561
rect 262154 234325 262196 234561
rect 261876 227561 262196 234325
rect 261876 227325 261918 227561
rect 262154 227325 262196 227561
rect 261876 220561 262196 227325
rect 261876 220325 261918 220561
rect 262154 220325 262196 220561
rect 261876 213561 262196 220325
rect 261876 213325 261918 213561
rect 262154 213325 262196 213561
rect 261876 206561 262196 213325
rect 261876 206325 261918 206561
rect 262154 206325 262196 206561
rect 261876 199561 262196 206325
rect 261876 199325 261918 199561
rect 262154 199325 262196 199561
rect 261876 192561 262196 199325
rect 261876 192325 261918 192561
rect 262154 192325 262196 192561
rect 261876 185561 262196 192325
rect 261876 185325 261918 185561
rect 262154 185325 262196 185561
rect 261876 178561 262196 185325
rect 261876 178325 261918 178561
rect 262154 178325 262196 178561
rect 261876 171561 262196 178325
rect 261876 171325 261918 171561
rect 262154 171325 262196 171561
rect 261876 164561 262196 171325
rect 261876 164325 261918 164561
rect 262154 164325 262196 164561
rect 261876 157561 262196 164325
rect 261876 157325 261918 157561
rect 262154 157325 262196 157561
rect 261876 150561 262196 157325
rect 261876 150325 261918 150561
rect 262154 150325 262196 150561
rect 261876 143561 262196 150325
rect 261876 143325 261918 143561
rect 262154 143325 262196 143561
rect 261876 136561 262196 143325
rect 261876 136325 261918 136561
rect 262154 136325 262196 136561
rect 261876 129561 262196 136325
rect 261876 129325 261918 129561
rect 262154 129325 262196 129561
rect 261876 122561 262196 129325
rect 261876 122325 261918 122561
rect 262154 122325 262196 122561
rect 261876 115561 262196 122325
rect 261876 115325 261918 115561
rect 262154 115325 262196 115561
rect 261876 108561 262196 115325
rect 261876 108325 261918 108561
rect 262154 108325 262196 108561
rect 261876 101561 262196 108325
rect 261876 101325 261918 101561
rect 262154 101325 262196 101561
rect 261876 94561 262196 101325
rect 261876 94325 261918 94561
rect 262154 94325 262196 94561
rect 261876 87561 262196 94325
rect 261876 87325 261918 87561
rect 262154 87325 262196 87561
rect 261876 80561 262196 87325
rect 261876 80325 261918 80561
rect 262154 80325 262196 80561
rect 261876 73561 262196 80325
rect 261876 73325 261918 73561
rect 262154 73325 262196 73561
rect 261876 66561 262196 73325
rect 261876 66325 261918 66561
rect 262154 66325 262196 66561
rect 261876 59561 262196 66325
rect 261876 59325 261918 59561
rect 262154 59325 262196 59561
rect 261876 52561 262196 59325
rect 261876 52325 261918 52561
rect 262154 52325 262196 52561
rect 261876 45561 262196 52325
rect 261876 45325 261918 45561
rect 262154 45325 262196 45561
rect 261876 38561 262196 45325
rect 261876 38325 261918 38561
rect 262154 38325 262196 38561
rect 261876 31561 262196 38325
rect 261876 31325 261918 31561
rect 262154 31325 262196 31561
rect 261876 24561 262196 31325
rect 261876 24325 261918 24561
rect 262154 24325 262196 24561
rect 261876 17561 262196 24325
rect 261876 17325 261918 17561
rect 262154 17325 262196 17561
rect 261876 10561 262196 17325
rect 261876 10325 261918 10561
rect 262154 10325 262196 10561
rect 261876 3561 262196 10325
rect 261876 3325 261918 3561
rect 262154 3325 262196 3561
rect 261876 -1706 262196 3325
rect 261876 -1942 261918 -1706
rect 262154 -1942 262196 -1706
rect 261876 -2026 262196 -1942
rect 261876 -2262 261918 -2026
rect 262154 -2262 262196 -2026
rect 261876 -2294 262196 -2262
rect 267144 705238 267464 706230
rect 267144 705002 267186 705238
rect 267422 705002 267464 705238
rect 267144 704918 267464 705002
rect 267144 704682 267186 704918
rect 267422 704682 267464 704918
rect 267144 695494 267464 704682
rect 267144 695258 267186 695494
rect 267422 695258 267464 695494
rect 267144 688494 267464 695258
rect 267144 688258 267186 688494
rect 267422 688258 267464 688494
rect 267144 681494 267464 688258
rect 267144 681258 267186 681494
rect 267422 681258 267464 681494
rect 267144 674494 267464 681258
rect 267144 674258 267186 674494
rect 267422 674258 267464 674494
rect 267144 667494 267464 674258
rect 267144 667258 267186 667494
rect 267422 667258 267464 667494
rect 267144 660494 267464 667258
rect 267144 660258 267186 660494
rect 267422 660258 267464 660494
rect 267144 653494 267464 660258
rect 267144 653258 267186 653494
rect 267422 653258 267464 653494
rect 267144 646494 267464 653258
rect 267144 646258 267186 646494
rect 267422 646258 267464 646494
rect 267144 639494 267464 646258
rect 267144 639258 267186 639494
rect 267422 639258 267464 639494
rect 267144 632494 267464 639258
rect 267144 632258 267186 632494
rect 267422 632258 267464 632494
rect 267144 625494 267464 632258
rect 267144 625258 267186 625494
rect 267422 625258 267464 625494
rect 267144 618494 267464 625258
rect 267144 618258 267186 618494
rect 267422 618258 267464 618494
rect 267144 611494 267464 618258
rect 267144 611258 267186 611494
rect 267422 611258 267464 611494
rect 267144 604494 267464 611258
rect 267144 604258 267186 604494
rect 267422 604258 267464 604494
rect 267144 597494 267464 604258
rect 267144 597258 267186 597494
rect 267422 597258 267464 597494
rect 267144 590494 267464 597258
rect 267144 590258 267186 590494
rect 267422 590258 267464 590494
rect 267144 583494 267464 590258
rect 267144 583258 267186 583494
rect 267422 583258 267464 583494
rect 267144 576494 267464 583258
rect 267144 576258 267186 576494
rect 267422 576258 267464 576494
rect 267144 569494 267464 576258
rect 267144 569258 267186 569494
rect 267422 569258 267464 569494
rect 267144 562494 267464 569258
rect 267144 562258 267186 562494
rect 267422 562258 267464 562494
rect 267144 555494 267464 562258
rect 267144 555258 267186 555494
rect 267422 555258 267464 555494
rect 267144 548494 267464 555258
rect 267144 548258 267186 548494
rect 267422 548258 267464 548494
rect 267144 541494 267464 548258
rect 267144 541258 267186 541494
rect 267422 541258 267464 541494
rect 267144 534494 267464 541258
rect 267144 534258 267186 534494
rect 267422 534258 267464 534494
rect 267144 527494 267464 534258
rect 267144 527258 267186 527494
rect 267422 527258 267464 527494
rect 267144 520494 267464 527258
rect 267144 520258 267186 520494
rect 267422 520258 267464 520494
rect 267144 513494 267464 520258
rect 267144 513258 267186 513494
rect 267422 513258 267464 513494
rect 267144 506494 267464 513258
rect 267144 506258 267186 506494
rect 267422 506258 267464 506494
rect 267144 499494 267464 506258
rect 267144 499258 267186 499494
rect 267422 499258 267464 499494
rect 267144 492494 267464 499258
rect 267144 492258 267186 492494
rect 267422 492258 267464 492494
rect 267144 485494 267464 492258
rect 267144 485258 267186 485494
rect 267422 485258 267464 485494
rect 267144 478494 267464 485258
rect 267144 478258 267186 478494
rect 267422 478258 267464 478494
rect 267144 471494 267464 478258
rect 267144 471258 267186 471494
rect 267422 471258 267464 471494
rect 267144 464494 267464 471258
rect 267144 464258 267186 464494
rect 267422 464258 267464 464494
rect 267144 457494 267464 464258
rect 267144 457258 267186 457494
rect 267422 457258 267464 457494
rect 267144 450494 267464 457258
rect 267144 450258 267186 450494
rect 267422 450258 267464 450494
rect 267144 443494 267464 450258
rect 267144 443258 267186 443494
rect 267422 443258 267464 443494
rect 267144 436494 267464 443258
rect 267144 436258 267186 436494
rect 267422 436258 267464 436494
rect 267144 429494 267464 436258
rect 267144 429258 267186 429494
rect 267422 429258 267464 429494
rect 267144 422494 267464 429258
rect 267144 422258 267186 422494
rect 267422 422258 267464 422494
rect 267144 415494 267464 422258
rect 267144 415258 267186 415494
rect 267422 415258 267464 415494
rect 267144 408494 267464 415258
rect 267144 408258 267186 408494
rect 267422 408258 267464 408494
rect 267144 401494 267464 408258
rect 267144 401258 267186 401494
rect 267422 401258 267464 401494
rect 267144 394494 267464 401258
rect 267144 394258 267186 394494
rect 267422 394258 267464 394494
rect 267144 387494 267464 394258
rect 267144 387258 267186 387494
rect 267422 387258 267464 387494
rect 267144 380494 267464 387258
rect 267144 380258 267186 380494
rect 267422 380258 267464 380494
rect 267144 373494 267464 380258
rect 267144 373258 267186 373494
rect 267422 373258 267464 373494
rect 267144 366494 267464 373258
rect 267144 366258 267186 366494
rect 267422 366258 267464 366494
rect 267144 359494 267464 366258
rect 267144 359258 267186 359494
rect 267422 359258 267464 359494
rect 267144 352494 267464 359258
rect 267144 352258 267186 352494
rect 267422 352258 267464 352494
rect 267144 345494 267464 352258
rect 267144 345258 267186 345494
rect 267422 345258 267464 345494
rect 267144 338494 267464 345258
rect 267144 338258 267186 338494
rect 267422 338258 267464 338494
rect 267144 331494 267464 338258
rect 267144 331258 267186 331494
rect 267422 331258 267464 331494
rect 267144 324494 267464 331258
rect 267144 324258 267186 324494
rect 267422 324258 267464 324494
rect 267144 317494 267464 324258
rect 267144 317258 267186 317494
rect 267422 317258 267464 317494
rect 267144 310494 267464 317258
rect 267144 310258 267186 310494
rect 267422 310258 267464 310494
rect 267144 303494 267464 310258
rect 267144 303258 267186 303494
rect 267422 303258 267464 303494
rect 267144 296494 267464 303258
rect 267144 296258 267186 296494
rect 267422 296258 267464 296494
rect 267144 289494 267464 296258
rect 267144 289258 267186 289494
rect 267422 289258 267464 289494
rect 267144 282494 267464 289258
rect 267144 282258 267186 282494
rect 267422 282258 267464 282494
rect 267144 275494 267464 282258
rect 267144 275258 267186 275494
rect 267422 275258 267464 275494
rect 267144 268494 267464 275258
rect 267144 268258 267186 268494
rect 267422 268258 267464 268494
rect 267144 261494 267464 268258
rect 267144 261258 267186 261494
rect 267422 261258 267464 261494
rect 267144 254494 267464 261258
rect 267144 254258 267186 254494
rect 267422 254258 267464 254494
rect 267144 247494 267464 254258
rect 267144 247258 267186 247494
rect 267422 247258 267464 247494
rect 267144 240494 267464 247258
rect 267144 240258 267186 240494
rect 267422 240258 267464 240494
rect 267144 233494 267464 240258
rect 267144 233258 267186 233494
rect 267422 233258 267464 233494
rect 267144 226494 267464 233258
rect 267144 226258 267186 226494
rect 267422 226258 267464 226494
rect 267144 219494 267464 226258
rect 267144 219258 267186 219494
rect 267422 219258 267464 219494
rect 267144 212494 267464 219258
rect 267144 212258 267186 212494
rect 267422 212258 267464 212494
rect 267144 205494 267464 212258
rect 267144 205258 267186 205494
rect 267422 205258 267464 205494
rect 267144 198494 267464 205258
rect 267144 198258 267186 198494
rect 267422 198258 267464 198494
rect 267144 191494 267464 198258
rect 267144 191258 267186 191494
rect 267422 191258 267464 191494
rect 267144 184494 267464 191258
rect 267144 184258 267186 184494
rect 267422 184258 267464 184494
rect 267144 177494 267464 184258
rect 267144 177258 267186 177494
rect 267422 177258 267464 177494
rect 267144 170494 267464 177258
rect 267144 170258 267186 170494
rect 267422 170258 267464 170494
rect 267144 163494 267464 170258
rect 267144 163258 267186 163494
rect 267422 163258 267464 163494
rect 267144 156494 267464 163258
rect 267144 156258 267186 156494
rect 267422 156258 267464 156494
rect 267144 149494 267464 156258
rect 267144 149258 267186 149494
rect 267422 149258 267464 149494
rect 267144 142494 267464 149258
rect 267144 142258 267186 142494
rect 267422 142258 267464 142494
rect 267144 135494 267464 142258
rect 267144 135258 267186 135494
rect 267422 135258 267464 135494
rect 267144 128494 267464 135258
rect 267144 128258 267186 128494
rect 267422 128258 267464 128494
rect 267144 121494 267464 128258
rect 267144 121258 267186 121494
rect 267422 121258 267464 121494
rect 267144 114494 267464 121258
rect 267144 114258 267186 114494
rect 267422 114258 267464 114494
rect 267144 107494 267464 114258
rect 267144 107258 267186 107494
rect 267422 107258 267464 107494
rect 267144 100494 267464 107258
rect 267144 100258 267186 100494
rect 267422 100258 267464 100494
rect 267144 93494 267464 100258
rect 267144 93258 267186 93494
rect 267422 93258 267464 93494
rect 267144 86494 267464 93258
rect 267144 86258 267186 86494
rect 267422 86258 267464 86494
rect 267144 79494 267464 86258
rect 267144 79258 267186 79494
rect 267422 79258 267464 79494
rect 267144 72494 267464 79258
rect 267144 72258 267186 72494
rect 267422 72258 267464 72494
rect 267144 65494 267464 72258
rect 267144 65258 267186 65494
rect 267422 65258 267464 65494
rect 267144 58494 267464 65258
rect 267144 58258 267186 58494
rect 267422 58258 267464 58494
rect 267144 51494 267464 58258
rect 267144 51258 267186 51494
rect 267422 51258 267464 51494
rect 267144 44494 267464 51258
rect 267144 44258 267186 44494
rect 267422 44258 267464 44494
rect 267144 37494 267464 44258
rect 267144 37258 267186 37494
rect 267422 37258 267464 37494
rect 267144 30494 267464 37258
rect 267144 30258 267186 30494
rect 267422 30258 267464 30494
rect 267144 23494 267464 30258
rect 267144 23258 267186 23494
rect 267422 23258 267464 23494
rect 267144 16494 267464 23258
rect 267144 16258 267186 16494
rect 267422 16258 267464 16494
rect 267144 9494 267464 16258
rect 267144 9258 267186 9494
rect 267422 9258 267464 9494
rect 267144 2494 267464 9258
rect 267144 2258 267186 2494
rect 267422 2258 267464 2494
rect 267144 -746 267464 2258
rect 267144 -982 267186 -746
rect 267422 -982 267464 -746
rect 267144 -1066 267464 -982
rect 267144 -1302 267186 -1066
rect 267422 -1302 267464 -1066
rect 267144 -2294 267464 -1302
rect 268876 706198 269196 706230
rect 268876 705962 268918 706198
rect 269154 705962 269196 706198
rect 268876 705878 269196 705962
rect 268876 705642 268918 705878
rect 269154 705642 269196 705878
rect 268876 696561 269196 705642
rect 268876 696325 268918 696561
rect 269154 696325 269196 696561
rect 268876 689561 269196 696325
rect 268876 689325 268918 689561
rect 269154 689325 269196 689561
rect 268876 682561 269196 689325
rect 268876 682325 268918 682561
rect 269154 682325 269196 682561
rect 268876 675561 269196 682325
rect 268876 675325 268918 675561
rect 269154 675325 269196 675561
rect 268876 668561 269196 675325
rect 268876 668325 268918 668561
rect 269154 668325 269196 668561
rect 268876 661561 269196 668325
rect 268876 661325 268918 661561
rect 269154 661325 269196 661561
rect 268876 654561 269196 661325
rect 268876 654325 268918 654561
rect 269154 654325 269196 654561
rect 268876 647561 269196 654325
rect 268876 647325 268918 647561
rect 269154 647325 269196 647561
rect 268876 640561 269196 647325
rect 268876 640325 268918 640561
rect 269154 640325 269196 640561
rect 268876 633561 269196 640325
rect 268876 633325 268918 633561
rect 269154 633325 269196 633561
rect 268876 626561 269196 633325
rect 268876 626325 268918 626561
rect 269154 626325 269196 626561
rect 268876 619561 269196 626325
rect 268876 619325 268918 619561
rect 269154 619325 269196 619561
rect 268876 612561 269196 619325
rect 268876 612325 268918 612561
rect 269154 612325 269196 612561
rect 268876 605561 269196 612325
rect 268876 605325 268918 605561
rect 269154 605325 269196 605561
rect 268876 598561 269196 605325
rect 268876 598325 268918 598561
rect 269154 598325 269196 598561
rect 268876 591561 269196 598325
rect 268876 591325 268918 591561
rect 269154 591325 269196 591561
rect 268876 584561 269196 591325
rect 268876 584325 268918 584561
rect 269154 584325 269196 584561
rect 268876 577561 269196 584325
rect 268876 577325 268918 577561
rect 269154 577325 269196 577561
rect 268876 570561 269196 577325
rect 268876 570325 268918 570561
rect 269154 570325 269196 570561
rect 268876 563561 269196 570325
rect 268876 563325 268918 563561
rect 269154 563325 269196 563561
rect 268876 556561 269196 563325
rect 268876 556325 268918 556561
rect 269154 556325 269196 556561
rect 268876 549561 269196 556325
rect 268876 549325 268918 549561
rect 269154 549325 269196 549561
rect 268876 542561 269196 549325
rect 268876 542325 268918 542561
rect 269154 542325 269196 542561
rect 268876 535561 269196 542325
rect 268876 535325 268918 535561
rect 269154 535325 269196 535561
rect 268876 528561 269196 535325
rect 268876 528325 268918 528561
rect 269154 528325 269196 528561
rect 268876 521561 269196 528325
rect 268876 521325 268918 521561
rect 269154 521325 269196 521561
rect 268876 514561 269196 521325
rect 268876 514325 268918 514561
rect 269154 514325 269196 514561
rect 268876 507561 269196 514325
rect 268876 507325 268918 507561
rect 269154 507325 269196 507561
rect 268876 500561 269196 507325
rect 268876 500325 268918 500561
rect 269154 500325 269196 500561
rect 268876 493561 269196 500325
rect 268876 493325 268918 493561
rect 269154 493325 269196 493561
rect 268876 486561 269196 493325
rect 268876 486325 268918 486561
rect 269154 486325 269196 486561
rect 268876 479561 269196 486325
rect 268876 479325 268918 479561
rect 269154 479325 269196 479561
rect 268876 472561 269196 479325
rect 268876 472325 268918 472561
rect 269154 472325 269196 472561
rect 268876 465561 269196 472325
rect 268876 465325 268918 465561
rect 269154 465325 269196 465561
rect 268876 458561 269196 465325
rect 268876 458325 268918 458561
rect 269154 458325 269196 458561
rect 268876 451561 269196 458325
rect 268876 451325 268918 451561
rect 269154 451325 269196 451561
rect 268876 444561 269196 451325
rect 268876 444325 268918 444561
rect 269154 444325 269196 444561
rect 268876 437561 269196 444325
rect 268876 437325 268918 437561
rect 269154 437325 269196 437561
rect 268876 430561 269196 437325
rect 268876 430325 268918 430561
rect 269154 430325 269196 430561
rect 268876 423561 269196 430325
rect 268876 423325 268918 423561
rect 269154 423325 269196 423561
rect 268876 416561 269196 423325
rect 268876 416325 268918 416561
rect 269154 416325 269196 416561
rect 268876 409561 269196 416325
rect 268876 409325 268918 409561
rect 269154 409325 269196 409561
rect 268876 402561 269196 409325
rect 268876 402325 268918 402561
rect 269154 402325 269196 402561
rect 268876 395561 269196 402325
rect 268876 395325 268918 395561
rect 269154 395325 269196 395561
rect 268876 388561 269196 395325
rect 268876 388325 268918 388561
rect 269154 388325 269196 388561
rect 268876 381561 269196 388325
rect 268876 381325 268918 381561
rect 269154 381325 269196 381561
rect 268876 374561 269196 381325
rect 268876 374325 268918 374561
rect 269154 374325 269196 374561
rect 268876 367561 269196 374325
rect 268876 367325 268918 367561
rect 269154 367325 269196 367561
rect 268876 360561 269196 367325
rect 268876 360325 268918 360561
rect 269154 360325 269196 360561
rect 268876 353561 269196 360325
rect 268876 353325 268918 353561
rect 269154 353325 269196 353561
rect 268876 346561 269196 353325
rect 268876 346325 268918 346561
rect 269154 346325 269196 346561
rect 268876 339561 269196 346325
rect 268876 339325 268918 339561
rect 269154 339325 269196 339561
rect 268876 332561 269196 339325
rect 268876 332325 268918 332561
rect 269154 332325 269196 332561
rect 268876 325561 269196 332325
rect 268876 325325 268918 325561
rect 269154 325325 269196 325561
rect 268876 318561 269196 325325
rect 268876 318325 268918 318561
rect 269154 318325 269196 318561
rect 268876 311561 269196 318325
rect 268876 311325 268918 311561
rect 269154 311325 269196 311561
rect 268876 304561 269196 311325
rect 268876 304325 268918 304561
rect 269154 304325 269196 304561
rect 268876 297561 269196 304325
rect 268876 297325 268918 297561
rect 269154 297325 269196 297561
rect 268876 290561 269196 297325
rect 268876 290325 268918 290561
rect 269154 290325 269196 290561
rect 268876 283561 269196 290325
rect 268876 283325 268918 283561
rect 269154 283325 269196 283561
rect 268876 276561 269196 283325
rect 268876 276325 268918 276561
rect 269154 276325 269196 276561
rect 268876 269561 269196 276325
rect 268876 269325 268918 269561
rect 269154 269325 269196 269561
rect 268876 262561 269196 269325
rect 268876 262325 268918 262561
rect 269154 262325 269196 262561
rect 268876 255561 269196 262325
rect 268876 255325 268918 255561
rect 269154 255325 269196 255561
rect 268876 248561 269196 255325
rect 268876 248325 268918 248561
rect 269154 248325 269196 248561
rect 268876 241561 269196 248325
rect 268876 241325 268918 241561
rect 269154 241325 269196 241561
rect 268876 234561 269196 241325
rect 268876 234325 268918 234561
rect 269154 234325 269196 234561
rect 268876 227561 269196 234325
rect 268876 227325 268918 227561
rect 269154 227325 269196 227561
rect 268876 220561 269196 227325
rect 268876 220325 268918 220561
rect 269154 220325 269196 220561
rect 268876 213561 269196 220325
rect 268876 213325 268918 213561
rect 269154 213325 269196 213561
rect 268876 206561 269196 213325
rect 268876 206325 268918 206561
rect 269154 206325 269196 206561
rect 268876 199561 269196 206325
rect 268876 199325 268918 199561
rect 269154 199325 269196 199561
rect 268876 192561 269196 199325
rect 268876 192325 268918 192561
rect 269154 192325 269196 192561
rect 268876 185561 269196 192325
rect 268876 185325 268918 185561
rect 269154 185325 269196 185561
rect 268876 178561 269196 185325
rect 268876 178325 268918 178561
rect 269154 178325 269196 178561
rect 268876 171561 269196 178325
rect 268876 171325 268918 171561
rect 269154 171325 269196 171561
rect 268876 164561 269196 171325
rect 268876 164325 268918 164561
rect 269154 164325 269196 164561
rect 268876 157561 269196 164325
rect 268876 157325 268918 157561
rect 269154 157325 269196 157561
rect 268876 150561 269196 157325
rect 268876 150325 268918 150561
rect 269154 150325 269196 150561
rect 268876 143561 269196 150325
rect 268876 143325 268918 143561
rect 269154 143325 269196 143561
rect 268876 136561 269196 143325
rect 268876 136325 268918 136561
rect 269154 136325 269196 136561
rect 268876 129561 269196 136325
rect 268876 129325 268918 129561
rect 269154 129325 269196 129561
rect 268876 122561 269196 129325
rect 268876 122325 268918 122561
rect 269154 122325 269196 122561
rect 268876 115561 269196 122325
rect 268876 115325 268918 115561
rect 269154 115325 269196 115561
rect 268876 108561 269196 115325
rect 268876 108325 268918 108561
rect 269154 108325 269196 108561
rect 268876 101561 269196 108325
rect 268876 101325 268918 101561
rect 269154 101325 269196 101561
rect 268876 94561 269196 101325
rect 268876 94325 268918 94561
rect 269154 94325 269196 94561
rect 268876 87561 269196 94325
rect 268876 87325 268918 87561
rect 269154 87325 269196 87561
rect 268876 80561 269196 87325
rect 268876 80325 268918 80561
rect 269154 80325 269196 80561
rect 268876 73561 269196 80325
rect 268876 73325 268918 73561
rect 269154 73325 269196 73561
rect 268876 66561 269196 73325
rect 268876 66325 268918 66561
rect 269154 66325 269196 66561
rect 268876 59561 269196 66325
rect 268876 59325 268918 59561
rect 269154 59325 269196 59561
rect 268876 52561 269196 59325
rect 268876 52325 268918 52561
rect 269154 52325 269196 52561
rect 268876 45561 269196 52325
rect 268876 45325 268918 45561
rect 269154 45325 269196 45561
rect 268876 38561 269196 45325
rect 268876 38325 268918 38561
rect 269154 38325 269196 38561
rect 268876 31561 269196 38325
rect 268876 31325 268918 31561
rect 269154 31325 269196 31561
rect 268876 24561 269196 31325
rect 268876 24325 268918 24561
rect 269154 24325 269196 24561
rect 268876 17561 269196 24325
rect 268876 17325 268918 17561
rect 269154 17325 269196 17561
rect 268876 10561 269196 17325
rect 268876 10325 268918 10561
rect 269154 10325 269196 10561
rect 268876 3561 269196 10325
rect 268876 3325 268918 3561
rect 269154 3325 269196 3561
rect 268876 -1706 269196 3325
rect 268876 -1942 268918 -1706
rect 269154 -1942 269196 -1706
rect 268876 -2026 269196 -1942
rect 268876 -2262 268918 -2026
rect 269154 -2262 269196 -2026
rect 268876 -2294 269196 -2262
rect 274144 705238 274464 706230
rect 274144 705002 274186 705238
rect 274422 705002 274464 705238
rect 274144 704918 274464 705002
rect 274144 704682 274186 704918
rect 274422 704682 274464 704918
rect 274144 695494 274464 704682
rect 274144 695258 274186 695494
rect 274422 695258 274464 695494
rect 274144 688494 274464 695258
rect 274144 688258 274186 688494
rect 274422 688258 274464 688494
rect 274144 681494 274464 688258
rect 274144 681258 274186 681494
rect 274422 681258 274464 681494
rect 274144 674494 274464 681258
rect 274144 674258 274186 674494
rect 274422 674258 274464 674494
rect 274144 667494 274464 674258
rect 274144 667258 274186 667494
rect 274422 667258 274464 667494
rect 274144 660494 274464 667258
rect 274144 660258 274186 660494
rect 274422 660258 274464 660494
rect 274144 653494 274464 660258
rect 274144 653258 274186 653494
rect 274422 653258 274464 653494
rect 274144 646494 274464 653258
rect 274144 646258 274186 646494
rect 274422 646258 274464 646494
rect 274144 639494 274464 646258
rect 274144 639258 274186 639494
rect 274422 639258 274464 639494
rect 274144 632494 274464 639258
rect 274144 632258 274186 632494
rect 274422 632258 274464 632494
rect 274144 625494 274464 632258
rect 274144 625258 274186 625494
rect 274422 625258 274464 625494
rect 274144 618494 274464 625258
rect 274144 618258 274186 618494
rect 274422 618258 274464 618494
rect 274144 611494 274464 618258
rect 274144 611258 274186 611494
rect 274422 611258 274464 611494
rect 274144 604494 274464 611258
rect 274144 604258 274186 604494
rect 274422 604258 274464 604494
rect 274144 597494 274464 604258
rect 274144 597258 274186 597494
rect 274422 597258 274464 597494
rect 274144 590494 274464 597258
rect 274144 590258 274186 590494
rect 274422 590258 274464 590494
rect 274144 583494 274464 590258
rect 274144 583258 274186 583494
rect 274422 583258 274464 583494
rect 274144 576494 274464 583258
rect 274144 576258 274186 576494
rect 274422 576258 274464 576494
rect 274144 569494 274464 576258
rect 274144 569258 274186 569494
rect 274422 569258 274464 569494
rect 274144 562494 274464 569258
rect 274144 562258 274186 562494
rect 274422 562258 274464 562494
rect 274144 555494 274464 562258
rect 274144 555258 274186 555494
rect 274422 555258 274464 555494
rect 274144 548494 274464 555258
rect 274144 548258 274186 548494
rect 274422 548258 274464 548494
rect 274144 541494 274464 548258
rect 274144 541258 274186 541494
rect 274422 541258 274464 541494
rect 274144 534494 274464 541258
rect 274144 534258 274186 534494
rect 274422 534258 274464 534494
rect 274144 527494 274464 534258
rect 274144 527258 274186 527494
rect 274422 527258 274464 527494
rect 274144 520494 274464 527258
rect 274144 520258 274186 520494
rect 274422 520258 274464 520494
rect 274144 513494 274464 520258
rect 274144 513258 274186 513494
rect 274422 513258 274464 513494
rect 274144 506494 274464 513258
rect 274144 506258 274186 506494
rect 274422 506258 274464 506494
rect 274144 499494 274464 506258
rect 274144 499258 274186 499494
rect 274422 499258 274464 499494
rect 274144 492494 274464 499258
rect 274144 492258 274186 492494
rect 274422 492258 274464 492494
rect 274144 485494 274464 492258
rect 274144 485258 274186 485494
rect 274422 485258 274464 485494
rect 274144 478494 274464 485258
rect 274144 478258 274186 478494
rect 274422 478258 274464 478494
rect 274144 471494 274464 478258
rect 274144 471258 274186 471494
rect 274422 471258 274464 471494
rect 274144 464494 274464 471258
rect 274144 464258 274186 464494
rect 274422 464258 274464 464494
rect 274144 457494 274464 464258
rect 274144 457258 274186 457494
rect 274422 457258 274464 457494
rect 274144 450494 274464 457258
rect 274144 450258 274186 450494
rect 274422 450258 274464 450494
rect 274144 443494 274464 450258
rect 274144 443258 274186 443494
rect 274422 443258 274464 443494
rect 274144 436494 274464 443258
rect 274144 436258 274186 436494
rect 274422 436258 274464 436494
rect 274144 429494 274464 436258
rect 274144 429258 274186 429494
rect 274422 429258 274464 429494
rect 274144 422494 274464 429258
rect 274144 422258 274186 422494
rect 274422 422258 274464 422494
rect 274144 415494 274464 422258
rect 274144 415258 274186 415494
rect 274422 415258 274464 415494
rect 274144 408494 274464 415258
rect 274144 408258 274186 408494
rect 274422 408258 274464 408494
rect 274144 401494 274464 408258
rect 274144 401258 274186 401494
rect 274422 401258 274464 401494
rect 274144 394494 274464 401258
rect 274144 394258 274186 394494
rect 274422 394258 274464 394494
rect 274144 387494 274464 394258
rect 274144 387258 274186 387494
rect 274422 387258 274464 387494
rect 274144 380494 274464 387258
rect 274144 380258 274186 380494
rect 274422 380258 274464 380494
rect 274144 373494 274464 380258
rect 274144 373258 274186 373494
rect 274422 373258 274464 373494
rect 274144 366494 274464 373258
rect 274144 366258 274186 366494
rect 274422 366258 274464 366494
rect 274144 359494 274464 366258
rect 274144 359258 274186 359494
rect 274422 359258 274464 359494
rect 274144 352494 274464 359258
rect 274144 352258 274186 352494
rect 274422 352258 274464 352494
rect 274144 345494 274464 352258
rect 274144 345258 274186 345494
rect 274422 345258 274464 345494
rect 274144 338494 274464 345258
rect 274144 338258 274186 338494
rect 274422 338258 274464 338494
rect 274144 331494 274464 338258
rect 274144 331258 274186 331494
rect 274422 331258 274464 331494
rect 274144 324494 274464 331258
rect 274144 324258 274186 324494
rect 274422 324258 274464 324494
rect 274144 317494 274464 324258
rect 274144 317258 274186 317494
rect 274422 317258 274464 317494
rect 274144 310494 274464 317258
rect 274144 310258 274186 310494
rect 274422 310258 274464 310494
rect 274144 303494 274464 310258
rect 274144 303258 274186 303494
rect 274422 303258 274464 303494
rect 274144 296494 274464 303258
rect 274144 296258 274186 296494
rect 274422 296258 274464 296494
rect 274144 289494 274464 296258
rect 274144 289258 274186 289494
rect 274422 289258 274464 289494
rect 274144 282494 274464 289258
rect 274144 282258 274186 282494
rect 274422 282258 274464 282494
rect 274144 275494 274464 282258
rect 274144 275258 274186 275494
rect 274422 275258 274464 275494
rect 274144 268494 274464 275258
rect 274144 268258 274186 268494
rect 274422 268258 274464 268494
rect 274144 261494 274464 268258
rect 274144 261258 274186 261494
rect 274422 261258 274464 261494
rect 274144 254494 274464 261258
rect 274144 254258 274186 254494
rect 274422 254258 274464 254494
rect 274144 247494 274464 254258
rect 274144 247258 274186 247494
rect 274422 247258 274464 247494
rect 274144 240494 274464 247258
rect 274144 240258 274186 240494
rect 274422 240258 274464 240494
rect 274144 233494 274464 240258
rect 274144 233258 274186 233494
rect 274422 233258 274464 233494
rect 274144 226494 274464 233258
rect 274144 226258 274186 226494
rect 274422 226258 274464 226494
rect 274144 219494 274464 226258
rect 274144 219258 274186 219494
rect 274422 219258 274464 219494
rect 274144 212494 274464 219258
rect 274144 212258 274186 212494
rect 274422 212258 274464 212494
rect 274144 205494 274464 212258
rect 274144 205258 274186 205494
rect 274422 205258 274464 205494
rect 274144 198494 274464 205258
rect 274144 198258 274186 198494
rect 274422 198258 274464 198494
rect 274144 191494 274464 198258
rect 274144 191258 274186 191494
rect 274422 191258 274464 191494
rect 274144 184494 274464 191258
rect 274144 184258 274186 184494
rect 274422 184258 274464 184494
rect 274144 177494 274464 184258
rect 274144 177258 274186 177494
rect 274422 177258 274464 177494
rect 274144 170494 274464 177258
rect 274144 170258 274186 170494
rect 274422 170258 274464 170494
rect 274144 163494 274464 170258
rect 274144 163258 274186 163494
rect 274422 163258 274464 163494
rect 274144 156494 274464 163258
rect 274144 156258 274186 156494
rect 274422 156258 274464 156494
rect 274144 149494 274464 156258
rect 274144 149258 274186 149494
rect 274422 149258 274464 149494
rect 274144 142494 274464 149258
rect 274144 142258 274186 142494
rect 274422 142258 274464 142494
rect 274144 135494 274464 142258
rect 274144 135258 274186 135494
rect 274422 135258 274464 135494
rect 274144 128494 274464 135258
rect 274144 128258 274186 128494
rect 274422 128258 274464 128494
rect 274144 121494 274464 128258
rect 274144 121258 274186 121494
rect 274422 121258 274464 121494
rect 274144 114494 274464 121258
rect 274144 114258 274186 114494
rect 274422 114258 274464 114494
rect 274144 107494 274464 114258
rect 274144 107258 274186 107494
rect 274422 107258 274464 107494
rect 274144 100494 274464 107258
rect 274144 100258 274186 100494
rect 274422 100258 274464 100494
rect 274144 93494 274464 100258
rect 274144 93258 274186 93494
rect 274422 93258 274464 93494
rect 274144 86494 274464 93258
rect 274144 86258 274186 86494
rect 274422 86258 274464 86494
rect 274144 79494 274464 86258
rect 274144 79258 274186 79494
rect 274422 79258 274464 79494
rect 274144 72494 274464 79258
rect 274144 72258 274186 72494
rect 274422 72258 274464 72494
rect 274144 65494 274464 72258
rect 274144 65258 274186 65494
rect 274422 65258 274464 65494
rect 274144 58494 274464 65258
rect 274144 58258 274186 58494
rect 274422 58258 274464 58494
rect 274144 51494 274464 58258
rect 274144 51258 274186 51494
rect 274422 51258 274464 51494
rect 274144 44494 274464 51258
rect 274144 44258 274186 44494
rect 274422 44258 274464 44494
rect 274144 37494 274464 44258
rect 274144 37258 274186 37494
rect 274422 37258 274464 37494
rect 274144 30494 274464 37258
rect 274144 30258 274186 30494
rect 274422 30258 274464 30494
rect 274144 23494 274464 30258
rect 274144 23258 274186 23494
rect 274422 23258 274464 23494
rect 274144 16494 274464 23258
rect 274144 16258 274186 16494
rect 274422 16258 274464 16494
rect 274144 9494 274464 16258
rect 274144 9258 274186 9494
rect 274422 9258 274464 9494
rect 274144 2494 274464 9258
rect 274144 2258 274186 2494
rect 274422 2258 274464 2494
rect 274144 -746 274464 2258
rect 274144 -982 274186 -746
rect 274422 -982 274464 -746
rect 274144 -1066 274464 -982
rect 274144 -1302 274186 -1066
rect 274422 -1302 274464 -1066
rect 274144 -2294 274464 -1302
rect 275876 706198 276196 706230
rect 275876 705962 275918 706198
rect 276154 705962 276196 706198
rect 275876 705878 276196 705962
rect 275876 705642 275918 705878
rect 276154 705642 276196 705878
rect 275876 696561 276196 705642
rect 275876 696325 275918 696561
rect 276154 696325 276196 696561
rect 275876 689561 276196 696325
rect 275876 689325 275918 689561
rect 276154 689325 276196 689561
rect 275876 682561 276196 689325
rect 275876 682325 275918 682561
rect 276154 682325 276196 682561
rect 275876 675561 276196 682325
rect 275876 675325 275918 675561
rect 276154 675325 276196 675561
rect 275876 668561 276196 675325
rect 275876 668325 275918 668561
rect 276154 668325 276196 668561
rect 275876 661561 276196 668325
rect 275876 661325 275918 661561
rect 276154 661325 276196 661561
rect 275876 654561 276196 661325
rect 275876 654325 275918 654561
rect 276154 654325 276196 654561
rect 275876 647561 276196 654325
rect 275876 647325 275918 647561
rect 276154 647325 276196 647561
rect 275876 640561 276196 647325
rect 275876 640325 275918 640561
rect 276154 640325 276196 640561
rect 275876 633561 276196 640325
rect 275876 633325 275918 633561
rect 276154 633325 276196 633561
rect 275876 626561 276196 633325
rect 275876 626325 275918 626561
rect 276154 626325 276196 626561
rect 275876 619561 276196 626325
rect 275876 619325 275918 619561
rect 276154 619325 276196 619561
rect 275876 612561 276196 619325
rect 275876 612325 275918 612561
rect 276154 612325 276196 612561
rect 275876 605561 276196 612325
rect 275876 605325 275918 605561
rect 276154 605325 276196 605561
rect 275876 598561 276196 605325
rect 275876 598325 275918 598561
rect 276154 598325 276196 598561
rect 275876 591561 276196 598325
rect 275876 591325 275918 591561
rect 276154 591325 276196 591561
rect 275876 584561 276196 591325
rect 275876 584325 275918 584561
rect 276154 584325 276196 584561
rect 275876 577561 276196 584325
rect 275876 577325 275918 577561
rect 276154 577325 276196 577561
rect 275876 570561 276196 577325
rect 275876 570325 275918 570561
rect 276154 570325 276196 570561
rect 275876 563561 276196 570325
rect 275876 563325 275918 563561
rect 276154 563325 276196 563561
rect 275876 556561 276196 563325
rect 275876 556325 275918 556561
rect 276154 556325 276196 556561
rect 275876 549561 276196 556325
rect 275876 549325 275918 549561
rect 276154 549325 276196 549561
rect 275876 542561 276196 549325
rect 275876 542325 275918 542561
rect 276154 542325 276196 542561
rect 275876 535561 276196 542325
rect 275876 535325 275918 535561
rect 276154 535325 276196 535561
rect 275876 528561 276196 535325
rect 275876 528325 275918 528561
rect 276154 528325 276196 528561
rect 275876 521561 276196 528325
rect 275876 521325 275918 521561
rect 276154 521325 276196 521561
rect 275876 514561 276196 521325
rect 275876 514325 275918 514561
rect 276154 514325 276196 514561
rect 275876 507561 276196 514325
rect 275876 507325 275918 507561
rect 276154 507325 276196 507561
rect 275876 500561 276196 507325
rect 275876 500325 275918 500561
rect 276154 500325 276196 500561
rect 275876 493561 276196 500325
rect 275876 493325 275918 493561
rect 276154 493325 276196 493561
rect 275876 486561 276196 493325
rect 275876 486325 275918 486561
rect 276154 486325 276196 486561
rect 275876 479561 276196 486325
rect 275876 479325 275918 479561
rect 276154 479325 276196 479561
rect 275876 472561 276196 479325
rect 275876 472325 275918 472561
rect 276154 472325 276196 472561
rect 275876 465561 276196 472325
rect 275876 465325 275918 465561
rect 276154 465325 276196 465561
rect 275876 458561 276196 465325
rect 275876 458325 275918 458561
rect 276154 458325 276196 458561
rect 275876 451561 276196 458325
rect 275876 451325 275918 451561
rect 276154 451325 276196 451561
rect 275876 444561 276196 451325
rect 275876 444325 275918 444561
rect 276154 444325 276196 444561
rect 275876 437561 276196 444325
rect 275876 437325 275918 437561
rect 276154 437325 276196 437561
rect 275876 430561 276196 437325
rect 275876 430325 275918 430561
rect 276154 430325 276196 430561
rect 275876 423561 276196 430325
rect 275876 423325 275918 423561
rect 276154 423325 276196 423561
rect 275876 416561 276196 423325
rect 275876 416325 275918 416561
rect 276154 416325 276196 416561
rect 275876 409561 276196 416325
rect 275876 409325 275918 409561
rect 276154 409325 276196 409561
rect 275876 402561 276196 409325
rect 275876 402325 275918 402561
rect 276154 402325 276196 402561
rect 275876 395561 276196 402325
rect 275876 395325 275918 395561
rect 276154 395325 276196 395561
rect 275876 388561 276196 395325
rect 275876 388325 275918 388561
rect 276154 388325 276196 388561
rect 275876 381561 276196 388325
rect 275876 381325 275918 381561
rect 276154 381325 276196 381561
rect 275876 374561 276196 381325
rect 275876 374325 275918 374561
rect 276154 374325 276196 374561
rect 275876 367561 276196 374325
rect 275876 367325 275918 367561
rect 276154 367325 276196 367561
rect 275876 360561 276196 367325
rect 275876 360325 275918 360561
rect 276154 360325 276196 360561
rect 275876 353561 276196 360325
rect 275876 353325 275918 353561
rect 276154 353325 276196 353561
rect 275876 346561 276196 353325
rect 275876 346325 275918 346561
rect 276154 346325 276196 346561
rect 275876 339561 276196 346325
rect 275876 339325 275918 339561
rect 276154 339325 276196 339561
rect 275876 332561 276196 339325
rect 275876 332325 275918 332561
rect 276154 332325 276196 332561
rect 275876 325561 276196 332325
rect 275876 325325 275918 325561
rect 276154 325325 276196 325561
rect 275876 318561 276196 325325
rect 275876 318325 275918 318561
rect 276154 318325 276196 318561
rect 275876 311561 276196 318325
rect 275876 311325 275918 311561
rect 276154 311325 276196 311561
rect 275876 304561 276196 311325
rect 275876 304325 275918 304561
rect 276154 304325 276196 304561
rect 275876 297561 276196 304325
rect 275876 297325 275918 297561
rect 276154 297325 276196 297561
rect 275876 290561 276196 297325
rect 275876 290325 275918 290561
rect 276154 290325 276196 290561
rect 275876 283561 276196 290325
rect 275876 283325 275918 283561
rect 276154 283325 276196 283561
rect 275876 276561 276196 283325
rect 275876 276325 275918 276561
rect 276154 276325 276196 276561
rect 275876 269561 276196 276325
rect 275876 269325 275918 269561
rect 276154 269325 276196 269561
rect 275876 262561 276196 269325
rect 275876 262325 275918 262561
rect 276154 262325 276196 262561
rect 275876 255561 276196 262325
rect 275876 255325 275918 255561
rect 276154 255325 276196 255561
rect 275876 248561 276196 255325
rect 275876 248325 275918 248561
rect 276154 248325 276196 248561
rect 275876 241561 276196 248325
rect 275876 241325 275918 241561
rect 276154 241325 276196 241561
rect 275876 234561 276196 241325
rect 275876 234325 275918 234561
rect 276154 234325 276196 234561
rect 275876 227561 276196 234325
rect 275876 227325 275918 227561
rect 276154 227325 276196 227561
rect 275876 220561 276196 227325
rect 275876 220325 275918 220561
rect 276154 220325 276196 220561
rect 275876 213561 276196 220325
rect 275876 213325 275918 213561
rect 276154 213325 276196 213561
rect 275876 206561 276196 213325
rect 275876 206325 275918 206561
rect 276154 206325 276196 206561
rect 275876 199561 276196 206325
rect 275876 199325 275918 199561
rect 276154 199325 276196 199561
rect 275876 192561 276196 199325
rect 275876 192325 275918 192561
rect 276154 192325 276196 192561
rect 275876 185561 276196 192325
rect 275876 185325 275918 185561
rect 276154 185325 276196 185561
rect 275876 178561 276196 185325
rect 275876 178325 275918 178561
rect 276154 178325 276196 178561
rect 275876 171561 276196 178325
rect 275876 171325 275918 171561
rect 276154 171325 276196 171561
rect 275876 164561 276196 171325
rect 275876 164325 275918 164561
rect 276154 164325 276196 164561
rect 275876 157561 276196 164325
rect 275876 157325 275918 157561
rect 276154 157325 276196 157561
rect 275876 150561 276196 157325
rect 275876 150325 275918 150561
rect 276154 150325 276196 150561
rect 275876 143561 276196 150325
rect 275876 143325 275918 143561
rect 276154 143325 276196 143561
rect 275876 136561 276196 143325
rect 275876 136325 275918 136561
rect 276154 136325 276196 136561
rect 275876 129561 276196 136325
rect 275876 129325 275918 129561
rect 276154 129325 276196 129561
rect 275876 122561 276196 129325
rect 275876 122325 275918 122561
rect 276154 122325 276196 122561
rect 275876 115561 276196 122325
rect 275876 115325 275918 115561
rect 276154 115325 276196 115561
rect 275876 108561 276196 115325
rect 275876 108325 275918 108561
rect 276154 108325 276196 108561
rect 275876 101561 276196 108325
rect 275876 101325 275918 101561
rect 276154 101325 276196 101561
rect 275876 94561 276196 101325
rect 275876 94325 275918 94561
rect 276154 94325 276196 94561
rect 275876 87561 276196 94325
rect 275876 87325 275918 87561
rect 276154 87325 276196 87561
rect 275876 80561 276196 87325
rect 275876 80325 275918 80561
rect 276154 80325 276196 80561
rect 275876 73561 276196 80325
rect 275876 73325 275918 73561
rect 276154 73325 276196 73561
rect 275876 66561 276196 73325
rect 275876 66325 275918 66561
rect 276154 66325 276196 66561
rect 275876 59561 276196 66325
rect 275876 59325 275918 59561
rect 276154 59325 276196 59561
rect 275876 52561 276196 59325
rect 275876 52325 275918 52561
rect 276154 52325 276196 52561
rect 275876 45561 276196 52325
rect 275876 45325 275918 45561
rect 276154 45325 276196 45561
rect 275876 38561 276196 45325
rect 275876 38325 275918 38561
rect 276154 38325 276196 38561
rect 275876 31561 276196 38325
rect 275876 31325 275918 31561
rect 276154 31325 276196 31561
rect 275876 24561 276196 31325
rect 275876 24325 275918 24561
rect 276154 24325 276196 24561
rect 275876 17561 276196 24325
rect 275876 17325 275918 17561
rect 276154 17325 276196 17561
rect 275876 10561 276196 17325
rect 275876 10325 275918 10561
rect 276154 10325 276196 10561
rect 275876 3561 276196 10325
rect 275876 3325 275918 3561
rect 276154 3325 276196 3561
rect 275876 -1706 276196 3325
rect 275876 -1942 275918 -1706
rect 276154 -1942 276196 -1706
rect 275876 -2026 276196 -1942
rect 275876 -2262 275918 -2026
rect 276154 -2262 276196 -2026
rect 275876 -2294 276196 -2262
rect 281144 705238 281464 706230
rect 281144 705002 281186 705238
rect 281422 705002 281464 705238
rect 281144 704918 281464 705002
rect 281144 704682 281186 704918
rect 281422 704682 281464 704918
rect 281144 695494 281464 704682
rect 281144 695258 281186 695494
rect 281422 695258 281464 695494
rect 281144 688494 281464 695258
rect 281144 688258 281186 688494
rect 281422 688258 281464 688494
rect 281144 681494 281464 688258
rect 281144 681258 281186 681494
rect 281422 681258 281464 681494
rect 281144 674494 281464 681258
rect 281144 674258 281186 674494
rect 281422 674258 281464 674494
rect 281144 667494 281464 674258
rect 281144 667258 281186 667494
rect 281422 667258 281464 667494
rect 281144 660494 281464 667258
rect 281144 660258 281186 660494
rect 281422 660258 281464 660494
rect 281144 653494 281464 660258
rect 281144 653258 281186 653494
rect 281422 653258 281464 653494
rect 281144 646494 281464 653258
rect 281144 646258 281186 646494
rect 281422 646258 281464 646494
rect 281144 639494 281464 646258
rect 281144 639258 281186 639494
rect 281422 639258 281464 639494
rect 281144 632494 281464 639258
rect 281144 632258 281186 632494
rect 281422 632258 281464 632494
rect 281144 625494 281464 632258
rect 281144 625258 281186 625494
rect 281422 625258 281464 625494
rect 281144 618494 281464 625258
rect 281144 618258 281186 618494
rect 281422 618258 281464 618494
rect 281144 611494 281464 618258
rect 281144 611258 281186 611494
rect 281422 611258 281464 611494
rect 281144 604494 281464 611258
rect 281144 604258 281186 604494
rect 281422 604258 281464 604494
rect 281144 597494 281464 604258
rect 281144 597258 281186 597494
rect 281422 597258 281464 597494
rect 281144 590494 281464 597258
rect 281144 590258 281186 590494
rect 281422 590258 281464 590494
rect 281144 583494 281464 590258
rect 281144 583258 281186 583494
rect 281422 583258 281464 583494
rect 281144 576494 281464 583258
rect 281144 576258 281186 576494
rect 281422 576258 281464 576494
rect 281144 569494 281464 576258
rect 281144 569258 281186 569494
rect 281422 569258 281464 569494
rect 281144 562494 281464 569258
rect 281144 562258 281186 562494
rect 281422 562258 281464 562494
rect 281144 555494 281464 562258
rect 281144 555258 281186 555494
rect 281422 555258 281464 555494
rect 281144 548494 281464 555258
rect 281144 548258 281186 548494
rect 281422 548258 281464 548494
rect 281144 541494 281464 548258
rect 281144 541258 281186 541494
rect 281422 541258 281464 541494
rect 281144 534494 281464 541258
rect 281144 534258 281186 534494
rect 281422 534258 281464 534494
rect 281144 527494 281464 534258
rect 281144 527258 281186 527494
rect 281422 527258 281464 527494
rect 281144 520494 281464 527258
rect 281144 520258 281186 520494
rect 281422 520258 281464 520494
rect 281144 513494 281464 520258
rect 281144 513258 281186 513494
rect 281422 513258 281464 513494
rect 281144 506494 281464 513258
rect 281144 506258 281186 506494
rect 281422 506258 281464 506494
rect 281144 499494 281464 506258
rect 281144 499258 281186 499494
rect 281422 499258 281464 499494
rect 281144 492494 281464 499258
rect 281144 492258 281186 492494
rect 281422 492258 281464 492494
rect 281144 485494 281464 492258
rect 281144 485258 281186 485494
rect 281422 485258 281464 485494
rect 281144 478494 281464 485258
rect 281144 478258 281186 478494
rect 281422 478258 281464 478494
rect 281144 471494 281464 478258
rect 281144 471258 281186 471494
rect 281422 471258 281464 471494
rect 281144 464494 281464 471258
rect 281144 464258 281186 464494
rect 281422 464258 281464 464494
rect 281144 457494 281464 464258
rect 281144 457258 281186 457494
rect 281422 457258 281464 457494
rect 281144 450494 281464 457258
rect 281144 450258 281186 450494
rect 281422 450258 281464 450494
rect 281144 443494 281464 450258
rect 281144 443258 281186 443494
rect 281422 443258 281464 443494
rect 281144 436494 281464 443258
rect 281144 436258 281186 436494
rect 281422 436258 281464 436494
rect 281144 429494 281464 436258
rect 281144 429258 281186 429494
rect 281422 429258 281464 429494
rect 281144 422494 281464 429258
rect 281144 422258 281186 422494
rect 281422 422258 281464 422494
rect 281144 415494 281464 422258
rect 281144 415258 281186 415494
rect 281422 415258 281464 415494
rect 281144 408494 281464 415258
rect 281144 408258 281186 408494
rect 281422 408258 281464 408494
rect 281144 401494 281464 408258
rect 281144 401258 281186 401494
rect 281422 401258 281464 401494
rect 281144 394494 281464 401258
rect 281144 394258 281186 394494
rect 281422 394258 281464 394494
rect 281144 387494 281464 394258
rect 281144 387258 281186 387494
rect 281422 387258 281464 387494
rect 281144 380494 281464 387258
rect 281144 380258 281186 380494
rect 281422 380258 281464 380494
rect 281144 373494 281464 380258
rect 281144 373258 281186 373494
rect 281422 373258 281464 373494
rect 281144 366494 281464 373258
rect 281144 366258 281186 366494
rect 281422 366258 281464 366494
rect 281144 359494 281464 366258
rect 281144 359258 281186 359494
rect 281422 359258 281464 359494
rect 281144 352494 281464 359258
rect 281144 352258 281186 352494
rect 281422 352258 281464 352494
rect 281144 345494 281464 352258
rect 281144 345258 281186 345494
rect 281422 345258 281464 345494
rect 281144 338494 281464 345258
rect 281144 338258 281186 338494
rect 281422 338258 281464 338494
rect 281144 331494 281464 338258
rect 281144 331258 281186 331494
rect 281422 331258 281464 331494
rect 281144 324494 281464 331258
rect 281144 324258 281186 324494
rect 281422 324258 281464 324494
rect 281144 317494 281464 324258
rect 281144 317258 281186 317494
rect 281422 317258 281464 317494
rect 281144 310494 281464 317258
rect 281144 310258 281186 310494
rect 281422 310258 281464 310494
rect 281144 303494 281464 310258
rect 281144 303258 281186 303494
rect 281422 303258 281464 303494
rect 281144 296494 281464 303258
rect 281144 296258 281186 296494
rect 281422 296258 281464 296494
rect 281144 289494 281464 296258
rect 281144 289258 281186 289494
rect 281422 289258 281464 289494
rect 281144 282494 281464 289258
rect 281144 282258 281186 282494
rect 281422 282258 281464 282494
rect 281144 275494 281464 282258
rect 281144 275258 281186 275494
rect 281422 275258 281464 275494
rect 281144 268494 281464 275258
rect 281144 268258 281186 268494
rect 281422 268258 281464 268494
rect 281144 261494 281464 268258
rect 281144 261258 281186 261494
rect 281422 261258 281464 261494
rect 281144 254494 281464 261258
rect 281144 254258 281186 254494
rect 281422 254258 281464 254494
rect 281144 247494 281464 254258
rect 281144 247258 281186 247494
rect 281422 247258 281464 247494
rect 281144 240494 281464 247258
rect 281144 240258 281186 240494
rect 281422 240258 281464 240494
rect 281144 233494 281464 240258
rect 281144 233258 281186 233494
rect 281422 233258 281464 233494
rect 281144 226494 281464 233258
rect 281144 226258 281186 226494
rect 281422 226258 281464 226494
rect 281144 219494 281464 226258
rect 281144 219258 281186 219494
rect 281422 219258 281464 219494
rect 281144 212494 281464 219258
rect 281144 212258 281186 212494
rect 281422 212258 281464 212494
rect 281144 205494 281464 212258
rect 281144 205258 281186 205494
rect 281422 205258 281464 205494
rect 281144 198494 281464 205258
rect 281144 198258 281186 198494
rect 281422 198258 281464 198494
rect 281144 191494 281464 198258
rect 281144 191258 281186 191494
rect 281422 191258 281464 191494
rect 281144 184494 281464 191258
rect 281144 184258 281186 184494
rect 281422 184258 281464 184494
rect 281144 177494 281464 184258
rect 281144 177258 281186 177494
rect 281422 177258 281464 177494
rect 281144 170494 281464 177258
rect 281144 170258 281186 170494
rect 281422 170258 281464 170494
rect 281144 163494 281464 170258
rect 281144 163258 281186 163494
rect 281422 163258 281464 163494
rect 281144 156494 281464 163258
rect 281144 156258 281186 156494
rect 281422 156258 281464 156494
rect 281144 149494 281464 156258
rect 281144 149258 281186 149494
rect 281422 149258 281464 149494
rect 281144 142494 281464 149258
rect 281144 142258 281186 142494
rect 281422 142258 281464 142494
rect 281144 135494 281464 142258
rect 281144 135258 281186 135494
rect 281422 135258 281464 135494
rect 281144 128494 281464 135258
rect 281144 128258 281186 128494
rect 281422 128258 281464 128494
rect 281144 121494 281464 128258
rect 281144 121258 281186 121494
rect 281422 121258 281464 121494
rect 281144 114494 281464 121258
rect 281144 114258 281186 114494
rect 281422 114258 281464 114494
rect 281144 107494 281464 114258
rect 281144 107258 281186 107494
rect 281422 107258 281464 107494
rect 281144 100494 281464 107258
rect 281144 100258 281186 100494
rect 281422 100258 281464 100494
rect 281144 93494 281464 100258
rect 281144 93258 281186 93494
rect 281422 93258 281464 93494
rect 281144 86494 281464 93258
rect 281144 86258 281186 86494
rect 281422 86258 281464 86494
rect 281144 79494 281464 86258
rect 281144 79258 281186 79494
rect 281422 79258 281464 79494
rect 281144 72494 281464 79258
rect 281144 72258 281186 72494
rect 281422 72258 281464 72494
rect 281144 65494 281464 72258
rect 281144 65258 281186 65494
rect 281422 65258 281464 65494
rect 281144 58494 281464 65258
rect 281144 58258 281186 58494
rect 281422 58258 281464 58494
rect 281144 51494 281464 58258
rect 281144 51258 281186 51494
rect 281422 51258 281464 51494
rect 281144 44494 281464 51258
rect 281144 44258 281186 44494
rect 281422 44258 281464 44494
rect 281144 37494 281464 44258
rect 281144 37258 281186 37494
rect 281422 37258 281464 37494
rect 281144 30494 281464 37258
rect 281144 30258 281186 30494
rect 281422 30258 281464 30494
rect 281144 23494 281464 30258
rect 281144 23258 281186 23494
rect 281422 23258 281464 23494
rect 281144 16494 281464 23258
rect 281144 16258 281186 16494
rect 281422 16258 281464 16494
rect 281144 9494 281464 16258
rect 281144 9258 281186 9494
rect 281422 9258 281464 9494
rect 281144 2494 281464 9258
rect 281144 2258 281186 2494
rect 281422 2258 281464 2494
rect 281144 -746 281464 2258
rect 281144 -982 281186 -746
rect 281422 -982 281464 -746
rect 281144 -1066 281464 -982
rect 281144 -1302 281186 -1066
rect 281422 -1302 281464 -1066
rect 281144 -2294 281464 -1302
rect 282876 706198 283196 706230
rect 282876 705962 282918 706198
rect 283154 705962 283196 706198
rect 282876 705878 283196 705962
rect 282876 705642 282918 705878
rect 283154 705642 283196 705878
rect 282876 696561 283196 705642
rect 282876 696325 282918 696561
rect 283154 696325 283196 696561
rect 282876 689561 283196 696325
rect 282876 689325 282918 689561
rect 283154 689325 283196 689561
rect 282876 682561 283196 689325
rect 282876 682325 282918 682561
rect 283154 682325 283196 682561
rect 282876 675561 283196 682325
rect 282876 675325 282918 675561
rect 283154 675325 283196 675561
rect 282876 668561 283196 675325
rect 282876 668325 282918 668561
rect 283154 668325 283196 668561
rect 282876 661561 283196 668325
rect 282876 661325 282918 661561
rect 283154 661325 283196 661561
rect 282876 654561 283196 661325
rect 282876 654325 282918 654561
rect 283154 654325 283196 654561
rect 282876 647561 283196 654325
rect 282876 647325 282918 647561
rect 283154 647325 283196 647561
rect 282876 640561 283196 647325
rect 282876 640325 282918 640561
rect 283154 640325 283196 640561
rect 282876 633561 283196 640325
rect 282876 633325 282918 633561
rect 283154 633325 283196 633561
rect 282876 626561 283196 633325
rect 282876 626325 282918 626561
rect 283154 626325 283196 626561
rect 282876 619561 283196 626325
rect 282876 619325 282918 619561
rect 283154 619325 283196 619561
rect 282876 612561 283196 619325
rect 282876 612325 282918 612561
rect 283154 612325 283196 612561
rect 282876 605561 283196 612325
rect 282876 605325 282918 605561
rect 283154 605325 283196 605561
rect 282876 598561 283196 605325
rect 282876 598325 282918 598561
rect 283154 598325 283196 598561
rect 282876 591561 283196 598325
rect 282876 591325 282918 591561
rect 283154 591325 283196 591561
rect 282876 584561 283196 591325
rect 282876 584325 282918 584561
rect 283154 584325 283196 584561
rect 282876 577561 283196 584325
rect 282876 577325 282918 577561
rect 283154 577325 283196 577561
rect 282876 570561 283196 577325
rect 282876 570325 282918 570561
rect 283154 570325 283196 570561
rect 282876 563561 283196 570325
rect 282876 563325 282918 563561
rect 283154 563325 283196 563561
rect 282876 556561 283196 563325
rect 282876 556325 282918 556561
rect 283154 556325 283196 556561
rect 282876 549561 283196 556325
rect 282876 549325 282918 549561
rect 283154 549325 283196 549561
rect 282876 542561 283196 549325
rect 282876 542325 282918 542561
rect 283154 542325 283196 542561
rect 282876 535561 283196 542325
rect 282876 535325 282918 535561
rect 283154 535325 283196 535561
rect 282876 528561 283196 535325
rect 282876 528325 282918 528561
rect 283154 528325 283196 528561
rect 282876 521561 283196 528325
rect 282876 521325 282918 521561
rect 283154 521325 283196 521561
rect 282876 514561 283196 521325
rect 282876 514325 282918 514561
rect 283154 514325 283196 514561
rect 282876 507561 283196 514325
rect 282876 507325 282918 507561
rect 283154 507325 283196 507561
rect 282876 500561 283196 507325
rect 282876 500325 282918 500561
rect 283154 500325 283196 500561
rect 282876 493561 283196 500325
rect 282876 493325 282918 493561
rect 283154 493325 283196 493561
rect 282876 486561 283196 493325
rect 282876 486325 282918 486561
rect 283154 486325 283196 486561
rect 282876 479561 283196 486325
rect 282876 479325 282918 479561
rect 283154 479325 283196 479561
rect 282876 472561 283196 479325
rect 282876 472325 282918 472561
rect 283154 472325 283196 472561
rect 282876 465561 283196 472325
rect 282876 465325 282918 465561
rect 283154 465325 283196 465561
rect 282876 458561 283196 465325
rect 282876 458325 282918 458561
rect 283154 458325 283196 458561
rect 282876 451561 283196 458325
rect 282876 451325 282918 451561
rect 283154 451325 283196 451561
rect 282876 444561 283196 451325
rect 282876 444325 282918 444561
rect 283154 444325 283196 444561
rect 282876 437561 283196 444325
rect 282876 437325 282918 437561
rect 283154 437325 283196 437561
rect 282876 430561 283196 437325
rect 282876 430325 282918 430561
rect 283154 430325 283196 430561
rect 282876 423561 283196 430325
rect 282876 423325 282918 423561
rect 283154 423325 283196 423561
rect 282876 416561 283196 423325
rect 282876 416325 282918 416561
rect 283154 416325 283196 416561
rect 282876 409561 283196 416325
rect 282876 409325 282918 409561
rect 283154 409325 283196 409561
rect 282876 402561 283196 409325
rect 282876 402325 282918 402561
rect 283154 402325 283196 402561
rect 282876 395561 283196 402325
rect 282876 395325 282918 395561
rect 283154 395325 283196 395561
rect 282876 388561 283196 395325
rect 282876 388325 282918 388561
rect 283154 388325 283196 388561
rect 282876 381561 283196 388325
rect 282876 381325 282918 381561
rect 283154 381325 283196 381561
rect 282876 374561 283196 381325
rect 282876 374325 282918 374561
rect 283154 374325 283196 374561
rect 282876 367561 283196 374325
rect 282876 367325 282918 367561
rect 283154 367325 283196 367561
rect 282876 360561 283196 367325
rect 282876 360325 282918 360561
rect 283154 360325 283196 360561
rect 282876 353561 283196 360325
rect 282876 353325 282918 353561
rect 283154 353325 283196 353561
rect 282876 346561 283196 353325
rect 282876 346325 282918 346561
rect 283154 346325 283196 346561
rect 282876 339561 283196 346325
rect 282876 339325 282918 339561
rect 283154 339325 283196 339561
rect 282876 332561 283196 339325
rect 282876 332325 282918 332561
rect 283154 332325 283196 332561
rect 282876 325561 283196 332325
rect 282876 325325 282918 325561
rect 283154 325325 283196 325561
rect 282876 318561 283196 325325
rect 282876 318325 282918 318561
rect 283154 318325 283196 318561
rect 282876 311561 283196 318325
rect 282876 311325 282918 311561
rect 283154 311325 283196 311561
rect 282876 304561 283196 311325
rect 282876 304325 282918 304561
rect 283154 304325 283196 304561
rect 282876 297561 283196 304325
rect 282876 297325 282918 297561
rect 283154 297325 283196 297561
rect 282876 290561 283196 297325
rect 282876 290325 282918 290561
rect 283154 290325 283196 290561
rect 282876 283561 283196 290325
rect 282876 283325 282918 283561
rect 283154 283325 283196 283561
rect 282876 276561 283196 283325
rect 282876 276325 282918 276561
rect 283154 276325 283196 276561
rect 282876 269561 283196 276325
rect 282876 269325 282918 269561
rect 283154 269325 283196 269561
rect 282876 262561 283196 269325
rect 282876 262325 282918 262561
rect 283154 262325 283196 262561
rect 282876 255561 283196 262325
rect 282876 255325 282918 255561
rect 283154 255325 283196 255561
rect 282876 248561 283196 255325
rect 282876 248325 282918 248561
rect 283154 248325 283196 248561
rect 282876 241561 283196 248325
rect 282876 241325 282918 241561
rect 283154 241325 283196 241561
rect 282876 234561 283196 241325
rect 282876 234325 282918 234561
rect 283154 234325 283196 234561
rect 282876 227561 283196 234325
rect 282876 227325 282918 227561
rect 283154 227325 283196 227561
rect 282876 220561 283196 227325
rect 282876 220325 282918 220561
rect 283154 220325 283196 220561
rect 282876 213561 283196 220325
rect 282876 213325 282918 213561
rect 283154 213325 283196 213561
rect 282876 206561 283196 213325
rect 282876 206325 282918 206561
rect 283154 206325 283196 206561
rect 282876 199561 283196 206325
rect 282876 199325 282918 199561
rect 283154 199325 283196 199561
rect 282876 192561 283196 199325
rect 282876 192325 282918 192561
rect 283154 192325 283196 192561
rect 282876 185561 283196 192325
rect 282876 185325 282918 185561
rect 283154 185325 283196 185561
rect 282876 178561 283196 185325
rect 282876 178325 282918 178561
rect 283154 178325 283196 178561
rect 282876 171561 283196 178325
rect 282876 171325 282918 171561
rect 283154 171325 283196 171561
rect 282876 164561 283196 171325
rect 282876 164325 282918 164561
rect 283154 164325 283196 164561
rect 282876 157561 283196 164325
rect 282876 157325 282918 157561
rect 283154 157325 283196 157561
rect 282876 150561 283196 157325
rect 282876 150325 282918 150561
rect 283154 150325 283196 150561
rect 282876 143561 283196 150325
rect 282876 143325 282918 143561
rect 283154 143325 283196 143561
rect 282876 136561 283196 143325
rect 282876 136325 282918 136561
rect 283154 136325 283196 136561
rect 282876 129561 283196 136325
rect 282876 129325 282918 129561
rect 283154 129325 283196 129561
rect 282876 122561 283196 129325
rect 282876 122325 282918 122561
rect 283154 122325 283196 122561
rect 282876 115561 283196 122325
rect 282876 115325 282918 115561
rect 283154 115325 283196 115561
rect 282876 108561 283196 115325
rect 282876 108325 282918 108561
rect 283154 108325 283196 108561
rect 282876 101561 283196 108325
rect 282876 101325 282918 101561
rect 283154 101325 283196 101561
rect 282876 94561 283196 101325
rect 282876 94325 282918 94561
rect 283154 94325 283196 94561
rect 282876 87561 283196 94325
rect 282876 87325 282918 87561
rect 283154 87325 283196 87561
rect 282876 80561 283196 87325
rect 282876 80325 282918 80561
rect 283154 80325 283196 80561
rect 282876 73561 283196 80325
rect 282876 73325 282918 73561
rect 283154 73325 283196 73561
rect 282876 66561 283196 73325
rect 282876 66325 282918 66561
rect 283154 66325 283196 66561
rect 282876 59561 283196 66325
rect 282876 59325 282918 59561
rect 283154 59325 283196 59561
rect 282876 52561 283196 59325
rect 282876 52325 282918 52561
rect 283154 52325 283196 52561
rect 282876 45561 283196 52325
rect 282876 45325 282918 45561
rect 283154 45325 283196 45561
rect 282876 38561 283196 45325
rect 282876 38325 282918 38561
rect 283154 38325 283196 38561
rect 282876 31561 283196 38325
rect 282876 31325 282918 31561
rect 283154 31325 283196 31561
rect 282876 24561 283196 31325
rect 282876 24325 282918 24561
rect 283154 24325 283196 24561
rect 282876 17561 283196 24325
rect 282876 17325 282918 17561
rect 283154 17325 283196 17561
rect 282876 10561 283196 17325
rect 282876 10325 282918 10561
rect 283154 10325 283196 10561
rect 282876 3561 283196 10325
rect 282876 3325 282918 3561
rect 283154 3325 283196 3561
rect 282876 -1706 283196 3325
rect 282876 -1942 282918 -1706
rect 283154 -1942 283196 -1706
rect 282876 -2026 283196 -1942
rect 282876 -2262 282918 -2026
rect 283154 -2262 283196 -2026
rect 282876 -2294 283196 -2262
rect 288144 705238 288464 706230
rect 288144 705002 288186 705238
rect 288422 705002 288464 705238
rect 288144 704918 288464 705002
rect 288144 704682 288186 704918
rect 288422 704682 288464 704918
rect 288144 695494 288464 704682
rect 288144 695258 288186 695494
rect 288422 695258 288464 695494
rect 288144 688494 288464 695258
rect 288144 688258 288186 688494
rect 288422 688258 288464 688494
rect 288144 681494 288464 688258
rect 288144 681258 288186 681494
rect 288422 681258 288464 681494
rect 288144 674494 288464 681258
rect 288144 674258 288186 674494
rect 288422 674258 288464 674494
rect 288144 667494 288464 674258
rect 288144 667258 288186 667494
rect 288422 667258 288464 667494
rect 288144 660494 288464 667258
rect 288144 660258 288186 660494
rect 288422 660258 288464 660494
rect 288144 653494 288464 660258
rect 288144 653258 288186 653494
rect 288422 653258 288464 653494
rect 288144 646494 288464 653258
rect 288144 646258 288186 646494
rect 288422 646258 288464 646494
rect 288144 639494 288464 646258
rect 288144 639258 288186 639494
rect 288422 639258 288464 639494
rect 288144 632494 288464 639258
rect 288144 632258 288186 632494
rect 288422 632258 288464 632494
rect 288144 625494 288464 632258
rect 288144 625258 288186 625494
rect 288422 625258 288464 625494
rect 288144 618494 288464 625258
rect 288144 618258 288186 618494
rect 288422 618258 288464 618494
rect 288144 611494 288464 618258
rect 288144 611258 288186 611494
rect 288422 611258 288464 611494
rect 288144 604494 288464 611258
rect 288144 604258 288186 604494
rect 288422 604258 288464 604494
rect 288144 597494 288464 604258
rect 288144 597258 288186 597494
rect 288422 597258 288464 597494
rect 288144 590494 288464 597258
rect 288144 590258 288186 590494
rect 288422 590258 288464 590494
rect 288144 583494 288464 590258
rect 288144 583258 288186 583494
rect 288422 583258 288464 583494
rect 288144 576494 288464 583258
rect 288144 576258 288186 576494
rect 288422 576258 288464 576494
rect 288144 569494 288464 576258
rect 288144 569258 288186 569494
rect 288422 569258 288464 569494
rect 288144 562494 288464 569258
rect 288144 562258 288186 562494
rect 288422 562258 288464 562494
rect 288144 555494 288464 562258
rect 288144 555258 288186 555494
rect 288422 555258 288464 555494
rect 288144 548494 288464 555258
rect 288144 548258 288186 548494
rect 288422 548258 288464 548494
rect 288144 541494 288464 548258
rect 288144 541258 288186 541494
rect 288422 541258 288464 541494
rect 288144 534494 288464 541258
rect 288144 534258 288186 534494
rect 288422 534258 288464 534494
rect 288144 527494 288464 534258
rect 288144 527258 288186 527494
rect 288422 527258 288464 527494
rect 288144 520494 288464 527258
rect 288144 520258 288186 520494
rect 288422 520258 288464 520494
rect 288144 513494 288464 520258
rect 288144 513258 288186 513494
rect 288422 513258 288464 513494
rect 288144 506494 288464 513258
rect 288144 506258 288186 506494
rect 288422 506258 288464 506494
rect 288144 499494 288464 506258
rect 288144 499258 288186 499494
rect 288422 499258 288464 499494
rect 288144 492494 288464 499258
rect 288144 492258 288186 492494
rect 288422 492258 288464 492494
rect 288144 485494 288464 492258
rect 288144 485258 288186 485494
rect 288422 485258 288464 485494
rect 288144 478494 288464 485258
rect 288144 478258 288186 478494
rect 288422 478258 288464 478494
rect 288144 471494 288464 478258
rect 288144 471258 288186 471494
rect 288422 471258 288464 471494
rect 288144 464494 288464 471258
rect 288144 464258 288186 464494
rect 288422 464258 288464 464494
rect 288144 457494 288464 464258
rect 288144 457258 288186 457494
rect 288422 457258 288464 457494
rect 288144 450494 288464 457258
rect 288144 450258 288186 450494
rect 288422 450258 288464 450494
rect 288144 443494 288464 450258
rect 288144 443258 288186 443494
rect 288422 443258 288464 443494
rect 288144 436494 288464 443258
rect 288144 436258 288186 436494
rect 288422 436258 288464 436494
rect 288144 429494 288464 436258
rect 288144 429258 288186 429494
rect 288422 429258 288464 429494
rect 288144 422494 288464 429258
rect 288144 422258 288186 422494
rect 288422 422258 288464 422494
rect 288144 415494 288464 422258
rect 288144 415258 288186 415494
rect 288422 415258 288464 415494
rect 288144 408494 288464 415258
rect 288144 408258 288186 408494
rect 288422 408258 288464 408494
rect 288144 401494 288464 408258
rect 288144 401258 288186 401494
rect 288422 401258 288464 401494
rect 288144 394494 288464 401258
rect 288144 394258 288186 394494
rect 288422 394258 288464 394494
rect 288144 387494 288464 394258
rect 288144 387258 288186 387494
rect 288422 387258 288464 387494
rect 288144 380494 288464 387258
rect 288144 380258 288186 380494
rect 288422 380258 288464 380494
rect 288144 373494 288464 380258
rect 288144 373258 288186 373494
rect 288422 373258 288464 373494
rect 288144 366494 288464 373258
rect 288144 366258 288186 366494
rect 288422 366258 288464 366494
rect 288144 359494 288464 366258
rect 288144 359258 288186 359494
rect 288422 359258 288464 359494
rect 288144 352494 288464 359258
rect 288144 352258 288186 352494
rect 288422 352258 288464 352494
rect 288144 345494 288464 352258
rect 288144 345258 288186 345494
rect 288422 345258 288464 345494
rect 288144 338494 288464 345258
rect 288144 338258 288186 338494
rect 288422 338258 288464 338494
rect 288144 331494 288464 338258
rect 288144 331258 288186 331494
rect 288422 331258 288464 331494
rect 288144 324494 288464 331258
rect 288144 324258 288186 324494
rect 288422 324258 288464 324494
rect 288144 317494 288464 324258
rect 288144 317258 288186 317494
rect 288422 317258 288464 317494
rect 288144 310494 288464 317258
rect 288144 310258 288186 310494
rect 288422 310258 288464 310494
rect 288144 303494 288464 310258
rect 288144 303258 288186 303494
rect 288422 303258 288464 303494
rect 288144 296494 288464 303258
rect 288144 296258 288186 296494
rect 288422 296258 288464 296494
rect 288144 289494 288464 296258
rect 288144 289258 288186 289494
rect 288422 289258 288464 289494
rect 288144 282494 288464 289258
rect 288144 282258 288186 282494
rect 288422 282258 288464 282494
rect 288144 275494 288464 282258
rect 288144 275258 288186 275494
rect 288422 275258 288464 275494
rect 288144 268494 288464 275258
rect 288144 268258 288186 268494
rect 288422 268258 288464 268494
rect 288144 261494 288464 268258
rect 288144 261258 288186 261494
rect 288422 261258 288464 261494
rect 288144 254494 288464 261258
rect 288144 254258 288186 254494
rect 288422 254258 288464 254494
rect 288144 247494 288464 254258
rect 288144 247258 288186 247494
rect 288422 247258 288464 247494
rect 288144 240494 288464 247258
rect 288144 240258 288186 240494
rect 288422 240258 288464 240494
rect 288144 233494 288464 240258
rect 288144 233258 288186 233494
rect 288422 233258 288464 233494
rect 288144 226494 288464 233258
rect 288144 226258 288186 226494
rect 288422 226258 288464 226494
rect 288144 219494 288464 226258
rect 288144 219258 288186 219494
rect 288422 219258 288464 219494
rect 288144 212494 288464 219258
rect 288144 212258 288186 212494
rect 288422 212258 288464 212494
rect 288144 205494 288464 212258
rect 288144 205258 288186 205494
rect 288422 205258 288464 205494
rect 288144 198494 288464 205258
rect 288144 198258 288186 198494
rect 288422 198258 288464 198494
rect 288144 191494 288464 198258
rect 288144 191258 288186 191494
rect 288422 191258 288464 191494
rect 288144 184494 288464 191258
rect 288144 184258 288186 184494
rect 288422 184258 288464 184494
rect 288144 177494 288464 184258
rect 288144 177258 288186 177494
rect 288422 177258 288464 177494
rect 288144 170494 288464 177258
rect 288144 170258 288186 170494
rect 288422 170258 288464 170494
rect 288144 163494 288464 170258
rect 288144 163258 288186 163494
rect 288422 163258 288464 163494
rect 288144 156494 288464 163258
rect 288144 156258 288186 156494
rect 288422 156258 288464 156494
rect 288144 149494 288464 156258
rect 288144 149258 288186 149494
rect 288422 149258 288464 149494
rect 288144 142494 288464 149258
rect 288144 142258 288186 142494
rect 288422 142258 288464 142494
rect 288144 135494 288464 142258
rect 288144 135258 288186 135494
rect 288422 135258 288464 135494
rect 288144 128494 288464 135258
rect 288144 128258 288186 128494
rect 288422 128258 288464 128494
rect 288144 121494 288464 128258
rect 288144 121258 288186 121494
rect 288422 121258 288464 121494
rect 288144 114494 288464 121258
rect 288144 114258 288186 114494
rect 288422 114258 288464 114494
rect 288144 107494 288464 114258
rect 288144 107258 288186 107494
rect 288422 107258 288464 107494
rect 288144 100494 288464 107258
rect 288144 100258 288186 100494
rect 288422 100258 288464 100494
rect 288144 93494 288464 100258
rect 288144 93258 288186 93494
rect 288422 93258 288464 93494
rect 288144 86494 288464 93258
rect 288144 86258 288186 86494
rect 288422 86258 288464 86494
rect 288144 79494 288464 86258
rect 288144 79258 288186 79494
rect 288422 79258 288464 79494
rect 288144 72494 288464 79258
rect 288144 72258 288186 72494
rect 288422 72258 288464 72494
rect 288144 65494 288464 72258
rect 288144 65258 288186 65494
rect 288422 65258 288464 65494
rect 288144 58494 288464 65258
rect 288144 58258 288186 58494
rect 288422 58258 288464 58494
rect 288144 51494 288464 58258
rect 288144 51258 288186 51494
rect 288422 51258 288464 51494
rect 288144 44494 288464 51258
rect 288144 44258 288186 44494
rect 288422 44258 288464 44494
rect 288144 37494 288464 44258
rect 288144 37258 288186 37494
rect 288422 37258 288464 37494
rect 288144 30494 288464 37258
rect 288144 30258 288186 30494
rect 288422 30258 288464 30494
rect 288144 23494 288464 30258
rect 288144 23258 288186 23494
rect 288422 23258 288464 23494
rect 288144 16494 288464 23258
rect 288144 16258 288186 16494
rect 288422 16258 288464 16494
rect 288144 9494 288464 16258
rect 288144 9258 288186 9494
rect 288422 9258 288464 9494
rect 288144 2494 288464 9258
rect 288144 2258 288186 2494
rect 288422 2258 288464 2494
rect 288144 -746 288464 2258
rect 288144 -982 288186 -746
rect 288422 -982 288464 -746
rect 288144 -1066 288464 -982
rect 288144 -1302 288186 -1066
rect 288422 -1302 288464 -1066
rect 288144 -2294 288464 -1302
rect 289876 706198 290196 706230
rect 289876 705962 289918 706198
rect 290154 705962 290196 706198
rect 289876 705878 290196 705962
rect 289876 705642 289918 705878
rect 290154 705642 290196 705878
rect 289876 696561 290196 705642
rect 289876 696325 289918 696561
rect 290154 696325 290196 696561
rect 289876 689561 290196 696325
rect 289876 689325 289918 689561
rect 290154 689325 290196 689561
rect 289876 682561 290196 689325
rect 289876 682325 289918 682561
rect 290154 682325 290196 682561
rect 289876 675561 290196 682325
rect 289876 675325 289918 675561
rect 290154 675325 290196 675561
rect 289876 668561 290196 675325
rect 289876 668325 289918 668561
rect 290154 668325 290196 668561
rect 289876 661561 290196 668325
rect 289876 661325 289918 661561
rect 290154 661325 290196 661561
rect 289876 654561 290196 661325
rect 289876 654325 289918 654561
rect 290154 654325 290196 654561
rect 289876 647561 290196 654325
rect 289876 647325 289918 647561
rect 290154 647325 290196 647561
rect 289876 640561 290196 647325
rect 289876 640325 289918 640561
rect 290154 640325 290196 640561
rect 289876 633561 290196 640325
rect 289876 633325 289918 633561
rect 290154 633325 290196 633561
rect 289876 626561 290196 633325
rect 289876 626325 289918 626561
rect 290154 626325 290196 626561
rect 289876 619561 290196 626325
rect 289876 619325 289918 619561
rect 290154 619325 290196 619561
rect 289876 612561 290196 619325
rect 289876 612325 289918 612561
rect 290154 612325 290196 612561
rect 289876 605561 290196 612325
rect 289876 605325 289918 605561
rect 290154 605325 290196 605561
rect 289876 598561 290196 605325
rect 289876 598325 289918 598561
rect 290154 598325 290196 598561
rect 289876 591561 290196 598325
rect 289876 591325 289918 591561
rect 290154 591325 290196 591561
rect 289876 584561 290196 591325
rect 289876 584325 289918 584561
rect 290154 584325 290196 584561
rect 289876 577561 290196 584325
rect 289876 577325 289918 577561
rect 290154 577325 290196 577561
rect 289876 570561 290196 577325
rect 289876 570325 289918 570561
rect 290154 570325 290196 570561
rect 289876 563561 290196 570325
rect 289876 563325 289918 563561
rect 290154 563325 290196 563561
rect 289876 556561 290196 563325
rect 289876 556325 289918 556561
rect 290154 556325 290196 556561
rect 289876 549561 290196 556325
rect 289876 549325 289918 549561
rect 290154 549325 290196 549561
rect 289876 542561 290196 549325
rect 289876 542325 289918 542561
rect 290154 542325 290196 542561
rect 289876 535561 290196 542325
rect 289876 535325 289918 535561
rect 290154 535325 290196 535561
rect 289876 528561 290196 535325
rect 289876 528325 289918 528561
rect 290154 528325 290196 528561
rect 289876 521561 290196 528325
rect 289876 521325 289918 521561
rect 290154 521325 290196 521561
rect 289876 514561 290196 521325
rect 289876 514325 289918 514561
rect 290154 514325 290196 514561
rect 289876 507561 290196 514325
rect 289876 507325 289918 507561
rect 290154 507325 290196 507561
rect 289876 500561 290196 507325
rect 289876 500325 289918 500561
rect 290154 500325 290196 500561
rect 289876 493561 290196 500325
rect 289876 493325 289918 493561
rect 290154 493325 290196 493561
rect 289876 486561 290196 493325
rect 289876 486325 289918 486561
rect 290154 486325 290196 486561
rect 289876 479561 290196 486325
rect 289876 479325 289918 479561
rect 290154 479325 290196 479561
rect 289876 472561 290196 479325
rect 289876 472325 289918 472561
rect 290154 472325 290196 472561
rect 289876 465561 290196 472325
rect 289876 465325 289918 465561
rect 290154 465325 290196 465561
rect 289876 458561 290196 465325
rect 289876 458325 289918 458561
rect 290154 458325 290196 458561
rect 289876 451561 290196 458325
rect 289876 451325 289918 451561
rect 290154 451325 290196 451561
rect 289876 444561 290196 451325
rect 289876 444325 289918 444561
rect 290154 444325 290196 444561
rect 289876 437561 290196 444325
rect 289876 437325 289918 437561
rect 290154 437325 290196 437561
rect 289876 430561 290196 437325
rect 289876 430325 289918 430561
rect 290154 430325 290196 430561
rect 289876 423561 290196 430325
rect 289876 423325 289918 423561
rect 290154 423325 290196 423561
rect 289876 416561 290196 423325
rect 289876 416325 289918 416561
rect 290154 416325 290196 416561
rect 289876 409561 290196 416325
rect 289876 409325 289918 409561
rect 290154 409325 290196 409561
rect 289876 402561 290196 409325
rect 289876 402325 289918 402561
rect 290154 402325 290196 402561
rect 289876 395561 290196 402325
rect 289876 395325 289918 395561
rect 290154 395325 290196 395561
rect 289876 388561 290196 395325
rect 289876 388325 289918 388561
rect 290154 388325 290196 388561
rect 289876 381561 290196 388325
rect 289876 381325 289918 381561
rect 290154 381325 290196 381561
rect 289876 374561 290196 381325
rect 289876 374325 289918 374561
rect 290154 374325 290196 374561
rect 289876 367561 290196 374325
rect 295144 705238 295464 706230
rect 295144 705002 295186 705238
rect 295422 705002 295464 705238
rect 295144 704918 295464 705002
rect 295144 704682 295186 704918
rect 295422 704682 295464 704918
rect 295144 695494 295464 704682
rect 295144 695258 295186 695494
rect 295422 695258 295464 695494
rect 295144 688494 295464 695258
rect 295144 688258 295186 688494
rect 295422 688258 295464 688494
rect 295144 681494 295464 688258
rect 295144 681258 295186 681494
rect 295422 681258 295464 681494
rect 295144 674494 295464 681258
rect 295144 674258 295186 674494
rect 295422 674258 295464 674494
rect 295144 667494 295464 674258
rect 295144 667258 295186 667494
rect 295422 667258 295464 667494
rect 295144 660494 295464 667258
rect 295144 660258 295186 660494
rect 295422 660258 295464 660494
rect 295144 653494 295464 660258
rect 295144 653258 295186 653494
rect 295422 653258 295464 653494
rect 295144 646494 295464 653258
rect 295144 646258 295186 646494
rect 295422 646258 295464 646494
rect 295144 639494 295464 646258
rect 295144 639258 295186 639494
rect 295422 639258 295464 639494
rect 295144 632494 295464 639258
rect 295144 632258 295186 632494
rect 295422 632258 295464 632494
rect 295144 625494 295464 632258
rect 295144 625258 295186 625494
rect 295422 625258 295464 625494
rect 295144 618494 295464 625258
rect 295144 618258 295186 618494
rect 295422 618258 295464 618494
rect 295144 611494 295464 618258
rect 295144 611258 295186 611494
rect 295422 611258 295464 611494
rect 295144 604494 295464 611258
rect 295144 604258 295186 604494
rect 295422 604258 295464 604494
rect 295144 597494 295464 604258
rect 295144 597258 295186 597494
rect 295422 597258 295464 597494
rect 295144 590494 295464 597258
rect 295144 590258 295186 590494
rect 295422 590258 295464 590494
rect 295144 583494 295464 590258
rect 295144 583258 295186 583494
rect 295422 583258 295464 583494
rect 295144 576494 295464 583258
rect 295144 576258 295186 576494
rect 295422 576258 295464 576494
rect 295144 569494 295464 576258
rect 295144 569258 295186 569494
rect 295422 569258 295464 569494
rect 295144 562494 295464 569258
rect 295144 562258 295186 562494
rect 295422 562258 295464 562494
rect 295144 555494 295464 562258
rect 295144 555258 295186 555494
rect 295422 555258 295464 555494
rect 295144 548494 295464 555258
rect 295144 548258 295186 548494
rect 295422 548258 295464 548494
rect 295144 541494 295464 548258
rect 295144 541258 295186 541494
rect 295422 541258 295464 541494
rect 295144 534494 295464 541258
rect 295144 534258 295186 534494
rect 295422 534258 295464 534494
rect 295144 527494 295464 534258
rect 295144 527258 295186 527494
rect 295422 527258 295464 527494
rect 295144 520494 295464 527258
rect 295144 520258 295186 520494
rect 295422 520258 295464 520494
rect 295144 513494 295464 520258
rect 295144 513258 295186 513494
rect 295422 513258 295464 513494
rect 295144 506494 295464 513258
rect 295144 506258 295186 506494
rect 295422 506258 295464 506494
rect 295144 499494 295464 506258
rect 295144 499258 295186 499494
rect 295422 499258 295464 499494
rect 295144 492494 295464 499258
rect 295144 492258 295186 492494
rect 295422 492258 295464 492494
rect 295144 490538 295464 492258
rect 295144 490474 295152 490538
rect 295216 490474 295232 490538
rect 295296 490474 295312 490538
rect 295376 490474 295392 490538
rect 295456 490474 295464 490538
rect 295144 490458 295464 490474
rect 295144 490394 295152 490458
rect 295216 490394 295232 490458
rect 295296 490394 295312 490458
rect 295376 490394 295392 490458
rect 295456 490394 295464 490458
rect 295144 490378 295464 490394
rect 295144 490314 295152 490378
rect 295216 490314 295232 490378
rect 295296 490314 295312 490378
rect 295376 490314 295392 490378
rect 295456 490314 295464 490378
rect 295144 485494 295464 490314
rect 295144 485258 295186 485494
rect 295422 485258 295464 485494
rect 295144 478494 295464 485258
rect 295144 478258 295186 478494
rect 295422 478258 295464 478494
rect 295144 471494 295464 478258
rect 295144 471258 295186 471494
rect 295422 471258 295464 471494
rect 295144 464494 295464 471258
rect 295144 464258 295186 464494
rect 295422 464258 295464 464494
rect 295144 457494 295464 464258
rect 295144 457258 295186 457494
rect 295422 457258 295464 457494
rect 295144 450494 295464 457258
rect 295144 450258 295186 450494
rect 295422 450258 295464 450494
rect 295144 443494 295464 450258
rect 295144 443258 295186 443494
rect 295422 443258 295464 443494
rect 295144 436494 295464 443258
rect 295144 436258 295186 436494
rect 295422 436258 295464 436494
rect 295144 429494 295464 436258
rect 295144 429258 295186 429494
rect 295422 429258 295464 429494
rect 295144 422494 295464 429258
rect 295144 422258 295186 422494
rect 295422 422258 295464 422494
rect 295144 415494 295464 422258
rect 295144 415258 295186 415494
rect 295422 415258 295464 415494
rect 295144 408494 295464 415258
rect 295144 408258 295186 408494
rect 295422 408258 295464 408494
rect 295144 401494 295464 408258
rect 295144 401258 295186 401494
rect 295422 401258 295464 401494
rect 295144 394494 295464 401258
rect 295144 394258 295186 394494
rect 295422 394258 295464 394494
rect 295144 388002 295464 394258
rect 295144 387938 295152 388002
rect 295216 387938 295232 388002
rect 295296 387938 295312 388002
rect 295376 387938 295392 388002
rect 295456 387938 295464 388002
rect 295144 387922 295464 387938
rect 295144 387858 295152 387922
rect 295216 387858 295232 387922
rect 295296 387858 295312 387922
rect 295376 387858 295392 387922
rect 295456 387858 295464 387922
rect 295144 387842 295464 387858
rect 295144 387778 295152 387842
rect 295216 387778 295232 387842
rect 295296 387778 295312 387842
rect 295376 387778 295392 387842
rect 295456 387778 295464 387842
rect 295144 387762 295464 387778
rect 295144 387698 295152 387762
rect 295216 387698 295232 387762
rect 295296 387698 295312 387762
rect 295376 387698 295392 387762
rect 295456 387698 295464 387762
rect 295144 387494 295464 387698
rect 295144 387258 295186 387494
rect 295422 387258 295464 387494
rect 295144 380494 295464 387258
rect 295144 380258 295186 380494
rect 295422 380258 295464 380494
rect 295144 373494 295464 380258
rect 295144 373258 295186 373494
rect 295422 373258 295464 373494
rect 295144 368640 295464 373258
rect 296876 706198 297196 706230
rect 296876 705962 296918 706198
rect 297154 705962 297196 706198
rect 296876 705878 297196 705962
rect 296876 705642 296918 705878
rect 297154 705642 297196 705878
rect 296876 696561 297196 705642
rect 296876 696325 296918 696561
rect 297154 696325 297196 696561
rect 296876 689561 297196 696325
rect 296876 689325 296918 689561
rect 297154 689325 297196 689561
rect 296876 682561 297196 689325
rect 296876 682325 296918 682561
rect 297154 682325 297196 682561
rect 296876 675561 297196 682325
rect 296876 675325 296918 675561
rect 297154 675325 297196 675561
rect 296876 668561 297196 675325
rect 296876 668325 296918 668561
rect 297154 668325 297196 668561
rect 296876 661561 297196 668325
rect 296876 661325 296918 661561
rect 297154 661325 297196 661561
rect 296876 654561 297196 661325
rect 296876 654325 296918 654561
rect 297154 654325 297196 654561
rect 296876 647561 297196 654325
rect 296876 647325 296918 647561
rect 297154 647325 297196 647561
rect 296876 640561 297196 647325
rect 296876 640325 296918 640561
rect 297154 640325 297196 640561
rect 296876 633561 297196 640325
rect 296876 633325 296918 633561
rect 297154 633325 297196 633561
rect 296876 626561 297196 633325
rect 296876 626325 296918 626561
rect 297154 626325 297196 626561
rect 296876 619561 297196 626325
rect 296876 619325 296918 619561
rect 297154 619325 297196 619561
rect 296876 612561 297196 619325
rect 296876 612325 296918 612561
rect 297154 612325 297196 612561
rect 296876 605561 297196 612325
rect 296876 605325 296918 605561
rect 297154 605325 297196 605561
rect 296876 598561 297196 605325
rect 296876 598325 296918 598561
rect 297154 598325 297196 598561
rect 296876 591561 297196 598325
rect 296876 591325 296918 591561
rect 297154 591325 297196 591561
rect 296876 584561 297196 591325
rect 296876 584325 296918 584561
rect 297154 584325 297196 584561
rect 296876 577561 297196 584325
rect 296876 577325 296918 577561
rect 297154 577325 297196 577561
rect 296876 570561 297196 577325
rect 296876 570325 296918 570561
rect 297154 570325 297196 570561
rect 296876 563561 297196 570325
rect 296876 563325 296918 563561
rect 297154 563325 297196 563561
rect 296876 556561 297196 563325
rect 296876 556325 296918 556561
rect 297154 556325 297196 556561
rect 296876 549561 297196 556325
rect 296876 549325 296918 549561
rect 297154 549325 297196 549561
rect 296876 542561 297196 549325
rect 296876 542325 296918 542561
rect 297154 542325 297196 542561
rect 296876 535561 297196 542325
rect 296876 535325 296918 535561
rect 297154 535325 297196 535561
rect 296876 528561 297196 535325
rect 296876 528325 296918 528561
rect 297154 528325 297196 528561
rect 296876 521561 297196 528325
rect 296876 521325 296918 521561
rect 297154 521325 297196 521561
rect 296876 514561 297196 521325
rect 296876 514325 296918 514561
rect 297154 514325 297196 514561
rect 296876 507561 297196 514325
rect 296876 507325 296918 507561
rect 297154 507325 297196 507561
rect 296876 500561 297196 507325
rect 296876 500325 296918 500561
rect 297154 500325 297196 500561
rect 296876 493561 297196 500325
rect 296876 493325 296918 493561
rect 297154 493325 297196 493561
rect 296876 491654 297196 493325
rect 296876 491590 296884 491654
rect 296948 491590 296964 491654
rect 297028 491590 297044 491654
rect 297108 491590 297124 491654
rect 297188 491590 297196 491654
rect 296876 491574 297196 491590
rect 296876 491510 296884 491574
rect 296948 491510 296964 491574
rect 297028 491510 297044 491574
rect 297108 491510 297124 491574
rect 297188 491510 297196 491574
rect 296876 491494 297196 491510
rect 296876 491430 296884 491494
rect 296948 491430 296964 491494
rect 297028 491430 297044 491494
rect 297108 491430 297124 491494
rect 297188 491430 297196 491494
rect 296876 491414 297196 491430
rect 296876 491350 296884 491414
rect 296948 491350 296964 491414
rect 297028 491350 297044 491414
rect 297108 491350 297124 491414
rect 297188 491350 297196 491414
rect 296876 486561 297196 491350
rect 296876 486325 296918 486561
rect 297154 486325 297196 486561
rect 296876 479561 297196 486325
rect 296876 479325 296918 479561
rect 297154 479325 297196 479561
rect 296876 473114 297196 479325
rect 296876 473050 296884 473114
rect 296948 473050 296964 473114
rect 297028 473050 297044 473114
rect 297108 473050 297124 473114
rect 297188 473050 297196 473114
rect 296876 473034 297196 473050
rect 296876 472970 296884 473034
rect 296948 472970 296964 473034
rect 297028 472970 297044 473034
rect 297108 472970 297124 473034
rect 297188 472970 297196 473034
rect 296876 472954 297196 472970
rect 296876 472890 296884 472954
rect 296948 472890 296964 472954
rect 297028 472890 297044 472954
rect 297108 472890 297124 472954
rect 297188 472890 297196 472954
rect 296876 472874 297196 472890
rect 296876 472810 296884 472874
rect 296948 472810 296964 472874
rect 297028 472810 297044 472874
rect 297108 472810 297124 472874
rect 297188 472810 297196 472874
rect 296876 472561 297196 472810
rect 296876 472325 296918 472561
rect 297154 472325 297196 472561
rect 296876 465561 297196 472325
rect 296876 465325 296918 465561
rect 297154 465325 297196 465561
rect 296876 458561 297196 465325
rect 296876 458325 296918 458561
rect 297154 458325 297196 458561
rect 296876 452058 297196 458325
rect 296876 451994 296884 452058
rect 296948 451994 296964 452058
rect 297028 451994 297044 452058
rect 297108 451994 297124 452058
rect 297188 451994 297196 452058
rect 296876 451978 297196 451994
rect 296876 451914 296884 451978
rect 296948 451914 296964 451978
rect 297028 451914 297044 451978
rect 297108 451914 297124 451978
rect 297188 451914 297196 451978
rect 296876 451898 297196 451914
rect 296876 451834 296884 451898
rect 296948 451834 296964 451898
rect 297028 451834 297044 451898
rect 297108 451834 297124 451898
rect 297188 451834 297196 451898
rect 296876 451818 297196 451834
rect 296876 451754 296884 451818
rect 296948 451754 296964 451818
rect 297028 451754 297044 451818
rect 297108 451754 297124 451818
rect 297188 451754 297196 451818
rect 296876 451738 297196 451754
rect 296876 451674 296884 451738
rect 296948 451674 296964 451738
rect 297028 451674 297044 451738
rect 297108 451674 297124 451738
rect 297188 451674 297196 451738
rect 296876 451658 297196 451674
rect 296876 451594 296884 451658
rect 296948 451594 296964 451658
rect 297028 451594 297044 451658
rect 297108 451594 297124 451658
rect 297188 451594 297196 451658
rect 296876 451578 297196 451594
rect 296876 451514 296884 451578
rect 296948 451561 296964 451578
rect 297028 451561 297044 451578
rect 297108 451561 297124 451578
rect 297188 451514 297196 451578
rect 296876 451498 296918 451514
rect 297154 451498 297196 451514
rect 296876 451434 296884 451498
rect 297188 451434 297196 451498
rect 296876 451418 296918 451434
rect 297154 451418 297196 451434
rect 296876 451354 296884 451418
rect 297188 451354 297196 451418
rect 296876 451338 296918 451354
rect 297154 451338 297196 451354
rect 296876 451274 296884 451338
rect 296948 451274 296964 451325
rect 297028 451274 297044 451325
rect 297108 451274 297124 451325
rect 297188 451274 297196 451338
rect 296876 444561 297196 451274
rect 296876 444325 296918 444561
rect 297154 444325 297196 444561
rect 296876 437561 297196 444325
rect 296876 437325 296918 437561
rect 297154 437325 297196 437561
rect 296876 430561 297196 437325
rect 296876 430325 296918 430561
rect 297154 430325 297196 430561
rect 296876 423561 297196 430325
rect 296876 423325 296918 423561
rect 297154 423325 297196 423561
rect 296876 416561 297196 423325
rect 296876 416325 296918 416561
rect 297154 416325 297196 416561
rect 296876 410084 297196 416325
rect 296876 410020 296884 410084
rect 296948 410020 296964 410084
rect 297028 410020 297044 410084
rect 297108 410020 297124 410084
rect 297188 410020 297196 410084
rect 296876 410004 297196 410020
rect 296876 409940 296884 410004
rect 296948 409940 296964 410004
rect 297028 409940 297044 410004
rect 297108 409940 297124 410004
rect 297188 409940 297196 410004
rect 296876 409924 297196 409940
rect 296876 409860 296884 409924
rect 296948 409860 296964 409924
rect 297028 409860 297044 409924
rect 297108 409860 297124 409924
rect 297188 409860 297196 409924
rect 296876 409844 297196 409860
rect 296876 409780 296884 409844
rect 296948 409780 296964 409844
rect 297028 409780 297044 409844
rect 297108 409780 297124 409844
rect 297188 409780 297196 409844
rect 296876 409561 297196 409780
rect 296876 409325 296918 409561
rect 297154 409325 297196 409561
rect 296876 402561 297196 409325
rect 296876 402325 296918 402561
rect 297154 402325 297196 402561
rect 296876 395561 297196 402325
rect 296876 395325 296918 395561
rect 297154 395325 297196 395561
rect 296876 389085 297196 395325
rect 296876 389021 296884 389085
rect 296948 389021 296964 389085
rect 297028 389021 297044 389085
rect 297108 389021 297124 389085
rect 297188 389021 297196 389085
rect 296876 389005 297196 389021
rect 296876 388941 296884 389005
rect 296948 388941 296964 389005
rect 297028 388941 297044 389005
rect 297108 388941 297124 389005
rect 297188 388941 297196 389005
rect 296876 388925 297196 388941
rect 296876 388861 296884 388925
rect 296948 388861 296964 388925
rect 297028 388861 297044 388925
rect 297108 388861 297124 388925
rect 297188 388861 297196 388925
rect 296876 388845 297196 388861
rect 296876 388781 296884 388845
rect 296948 388781 296964 388845
rect 297028 388781 297044 388845
rect 297108 388781 297124 388845
rect 297188 388781 297196 388845
rect 296876 388561 297196 388781
rect 296876 388325 296918 388561
rect 297154 388325 297196 388561
rect 296876 381561 297196 388325
rect 296876 381325 296918 381561
rect 297154 381325 297196 381561
rect 296876 374561 297196 381325
rect 296876 374325 296918 374561
rect 297154 374325 297196 374561
rect 296876 368640 297196 374325
rect 302144 705238 302464 706230
rect 302144 705002 302186 705238
rect 302422 705002 302464 705238
rect 302144 704918 302464 705002
rect 302144 704682 302186 704918
rect 302422 704682 302464 704918
rect 302144 695494 302464 704682
rect 302144 695258 302186 695494
rect 302422 695258 302464 695494
rect 302144 688494 302464 695258
rect 302144 688258 302186 688494
rect 302422 688258 302464 688494
rect 302144 681494 302464 688258
rect 302144 681258 302186 681494
rect 302422 681258 302464 681494
rect 302144 674494 302464 681258
rect 302144 674258 302186 674494
rect 302422 674258 302464 674494
rect 302144 667494 302464 674258
rect 302144 667258 302186 667494
rect 302422 667258 302464 667494
rect 302144 660494 302464 667258
rect 302144 660258 302186 660494
rect 302422 660258 302464 660494
rect 302144 653494 302464 660258
rect 302144 653258 302186 653494
rect 302422 653258 302464 653494
rect 302144 646494 302464 653258
rect 302144 646258 302186 646494
rect 302422 646258 302464 646494
rect 302144 639494 302464 646258
rect 302144 639258 302186 639494
rect 302422 639258 302464 639494
rect 302144 632494 302464 639258
rect 302144 632258 302186 632494
rect 302422 632258 302464 632494
rect 302144 625494 302464 632258
rect 302144 625258 302186 625494
rect 302422 625258 302464 625494
rect 302144 618494 302464 625258
rect 302144 618258 302186 618494
rect 302422 618258 302464 618494
rect 302144 611494 302464 618258
rect 302144 611258 302186 611494
rect 302422 611258 302464 611494
rect 302144 604494 302464 611258
rect 302144 604258 302186 604494
rect 302422 604258 302464 604494
rect 302144 597494 302464 604258
rect 302144 597258 302186 597494
rect 302422 597258 302464 597494
rect 302144 590494 302464 597258
rect 302144 590258 302186 590494
rect 302422 590258 302464 590494
rect 302144 583494 302464 590258
rect 302144 583258 302186 583494
rect 302422 583258 302464 583494
rect 302144 576494 302464 583258
rect 302144 576258 302186 576494
rect 302422 576258 302464 576494
rect 302144 569494 302464 576258
rect 302144 569258 302186 569494
rect 302422 569258 302464 569494
rect 302144 562494 302464 569258
rect 302144 562258 302186 562494
rect 302422 562258 302464 562494
rect 302144 555494 302464 562258
rect 302144 555258 302186 555494
rect 302422 555258 302464 555494
rect 302144 548494 302464 555258
rect 302144 548258 302186 548494
rect 302422 548258 302464 548494
rect 302144 541494 302464 548258
rect 302144 541258 302186 541494
rect 302422 541258 302464 541494
rect 302144 534494 302464 541258
rect 302144 534258 302186 534494
rect 302422 534258 302464 534494
rect 302144 527494 302464 534258
rect 302144 527258 302186 527494
rect 302422 527258 302464 527494
rect 302144 520494 302464 527258
rect 302144 520258 302186 520494
rect 302422 520258 302464 520494
rect 302144 513494 302464 520258
rect 302144 513258 302186 513494
rect 302422 513258 302464 513494
rect 302144 506494 302464 513258
rect 302144 506258 302186 506494
rect 302422 506258 302464 506494
rect 302144 499494 302464 506258
rect 302144 499258 302186 499494
rect 302422 499258 302464 499494
rect 302144 492494 302464 499258
rect 302144 492258 302186 492494
rect 302422 492258 302464 492494
rect 302144 485494 302464 492258
rect 302144 485258 302186 485494
rect 302422 485258 302464 485494
rect 302144 478494 302464 485258
rect 302144 478258 302186 478494
rect 302422 478258 302464 478494
rect 302144 472013 302464 478258
rect 302144 471949 302152 472013
rect 302216 471949 302232 472013
rect 302296 471949 302312 472013
rect 302376 471949 302392 472013
rect 302456 471949 302464 472013
rect 302144 471933 302464 471949
rect 302144 471869 302152 471933
rect 302216 471869 302232 471933
rect 302296 471869 302312 471933
rect 302376 471869 302392 471933
rect 302456 471869 302464 471933
rect 302144 471853 302464 471869
rect 302144 471789 302152 471853
rect 302216 471789 302232 471853
rect 302296 471789 302312 471853
rect 302376 471789 302392 471853
rect 302456 471789 302464 471853
rect 302144 471773 302464 471789
rect 302144 471709 302152 471773
rect 302216 471709 302232 471773
rect 302296 471709 302312 471773
rect 302376 471709 302392 471773
rect 302456 471709 302464 471773
rect 302144 471494 302464 471709
rect 302144 471258 302186 471494
rect 302422 471258 302464 471494
rect 302144 464494 302464 471258
rect 302144 464258 302186 464494
rect 302422 464258 302464 464494
rect 302144 457494 302464 464258
rect 302144 457258 302186 457494
rect 302422 457258 302464 457494
rect 302144 450494 302464 457258
rect 302144 450258 302186 450494
rect 302422 450258 302464 450494
rect 302144 443494 302464 450258
rect 302144 443258 302186 443494
rect 302422 443258 302464 443494
rect 302144 436494 302464 443258
rect 302144 436258 302186 436494
rect 302422 436258 302464 436494
rect 302144 429494 302464 436258
rect 302144 429258 302186 429494
rect 302422 429258 302464 429494
rect 302144 422494 302464 429258
rect 302144 422258 302186 422494
rect 302422 422258 302464 422494
rect 302144 415494 302464 422258
rect 302144 415258 302186 415494
rect 302422 415258 302464 415494
rect 302144 408998 302464 415258
rect 302144 408934 302152 408998
rect 302216 408934 302232 408998
rect 302296 408934 302312 408998
rect 302376 408934 302392 408998
rect 302456 408934 302464 408998
rect 302144 408918 302464 408934
rect 302144 408854 302152 408918
rect 302216 408854 302232 408918
rect 302296 408854 302312 408918
rect 302376 408854 302392 408918
rect 302456 408854 302464 408918
rect 302144 408838 302464 408854
rect 302144 408774 302152 408838
rect 302216 408774 302232 408838
rect 302296 408774 302312 408838
rect 302376 408774 302392 408838
rect 302456 408774 302464 408838
rect 302144 408758 302464 408774
rect 302144 408694 302152 408758
rect 302216 408694 302232 408758
rect 302296 408694 302312 408758
rect 302376 408694 302392 408758
rect 302456 408694 302464 408758
rect 302144 408494 302464 408694
rect 302144 408258 302186 408494
rect 302422 408258 302464 408494
rect 302144 401494 302464 408258
rect 302144 401258 302186 401494
rect 302422 401258 302464 401494
rect 302144 394494 302464 401258
rect 302144 394258 302186 394494
rect 302422 394258 302464 394494
rect 302144 387997 302464 394258
rect 302144 387933 302152 387997
rect 302216 387933 302232 387997
rect 302296 387933 302312 387997
rect 302376 387933 302392 387997
rect 302456 387933 302464 387997
rect 302144 387917 302464 387933
rect 302144 387853 302152 387917
rect 302216 387853 302232 387917
rect 302296 387853 302312 387917
rect 302376 387853 302392 387917
rect 302456 387853 302464 387917
rect 302144 387837 302464 387853
rect 302144 387773 302152 387837
rect 302216 387773 302232 387837
rect 302296 387773 302312 387837
rect 302376 387773 302392 387837
rect 302456 387773 302464 387837
rect 302144 387757 302464 387773
rect 302144 387693 302152 387757
rect 302216 387693 302232 387757
rect 302296 387693 302312 387757
rect 302376 387693 302392 387757
rect 302456 387693 302464 387757
rect 302144 387494 302464 387693
rect 302144 387258 302186 387494
rect 302422 387258 302464 387494
rect 302144 380494 302464 387258
rect 302144 380258 302186 380494
rect 302422 380258 302464 380494
rect 302144 373494 302464 380258
rect 302144 373258 302186 373494
rect 302422 373258 302464 373494
rect 302144 368640 302464 373258
rect 303876 706198 304196 706230
rect 303876 705962 303918 706198
rect 304154 705962 304196 706198
rect 303876 705878 304196 705962
rect 303876 705642 303918 705878
rect 304154 705642 304196 705878
rect 303876 696561 304196 705642
rect 303876 696325 303918 696561
rect 304154 696325 304196 696561
rect 303876 689561 304196 696325
rect 303876 689325 303918 689561
rect 304154 689325 304196 689561
rect 303876 682561 304196 689325
rect 303876 682325 303918 682561
rect 304154 682325 304196 682561
rect 303876 675561 304196 682325
rect 303876 675325 303918 675561
rect 304154 675325 304196 675561
rect 303876 668561 304196 675325
rect 303876 668325 303918 668561
rect 304154 668325 304196 668561
rect 303876 661561 304196 668325
rect 303876 661325 303918 661561
rect 304154 661325 304196 661561
rect 303876 654561 304196 661325
rect 303876 654325 303918 654561
rect 304154 654325 304196 654561
rect 303876 647561 304196 654325
rect 303876 647325 303918 647561
rect 304154 647325 304196 647561
rect 303876 640561 304196 647325
rect 303876 640325 303918 640561
rect 304154 640325 304196 640561
rect 303876 633561 304196 640325
rect 303876 633325 303918 633561
rect 304154 633325 304196 633561
rect 303876 626561 304196 633325
rect 303876 626325 303918 626561
rect 304154 626325 304196 626561
rect 303876 619561 304196 626325
rect 303876 619325 303918 619561
rect 304154 619325 304196 619561
rect 303876 612561 304196 619325
rect 303876 612325 303918 612561
rect 304154 612325 304196 612561
rect 303876 605561 304196 612325
rect 303876 605325 303918 605561
rect 304154 605325 304196 605561
rect 303876 598561 304196 605325
rect 303876 598325 303918 598561
rect 304154 598325 304196 598561
rect 303876 591561 304196 598325
rect 303876 591325 303918 591561
rect 304154 591325 304196 591561
rect 303876 584561 304196 591325
rect 303876 584325 303918 584561
rect 304154 584325 304196 584561
rect 303876 577561 304196 584325
rect 303876 577325 303918 577561
rect 304154 577325 304196 577561
rect 303876 570561 304196 577325
rect 303876 570325 303918 570561
rect 304154 570325 304196 570561
rect 303876 563561 304196 570325
rect 303876 563325 303918 563561
rect 304154 563325 304196 563561
rect 303876 556561 304196 563325
rect 303876 556325 303918 556561
rect 304154 556325 304196 556561
rect 303876 549561 304196 556325
rect 303876 549325 303918 549561
rect 304154 549325 304196 549561
rect 303876 542561 304196 549325
rect 303876 542325 303918 542561
rect 304154 542325 304196 542561
rect 303876 535561 304196 542325
rect 303876 535325 303918 535561
rect 304154 535325 304196 535561
rect 303876 528561 304196 535325
rect 303876 528325 303918 528561
rect 304154 528325 304196 528561
rect 303876 521561 304196 528325
rect 303876 521325 303918 521561
rect 304154 521325 304196 521561
rect 303876 514561 304196 521325
rect 303876 514325 303918 514561
rect 304154 514325 304196 514561
rect 303876 507561 304196 514325
rect 303876 507325 303918 507561
rect 304154 507325 304196 507561
rect 303876 500561 304196 507325
rect 303876 500325 303918 500561
rect 304154 500325 304196 500561
rect 303876 493561 304196 500325
rect 303876 493325 303918 493561
rect 304154 493325 304196 493561
rect 303876 491654 304196 493325
rect 303876 491590 303884 491654
rect 303948 491590 303964 491654
rect 304028 491590 304044 491654
rect 304108 491590 304124 491654
rect 304188 491590 304196 491654
rect 303876 491574 304196 491590
rect 303876 491510 303884 491574
rect 303948 491510 303964 491574
rect 304028 491510 304044 491574
rect 304108 491510 304124 491574
rect 304188 491510 304196 491574
rect 303876 491494 304196 491510
rect 303876 491430 303884 491494
rect 303948 491430 303964 491494
rect 304028 491430 304044 491494
rect 304108 491430 304124 491494
rect 304188 491430 304196 491494
rect 303876 491414 304196 491430
rect 303876 491350 303884 491414
rect 303948 491350 303964 491414
rect 304028 491350 304044 491414
rect 304108 491350 304124 491414
rect 304188 491350 304196 491414
rect 303876 489482 304196 491350
rect 303876 489418 303884 489482
rect 303948 489418 303964 489482
rect 304028 489418 304044 489482
rect 304108 489418 304124 489482
rect 304188 489418 304196 489482
rect 303876 489402 304196 489418
rect 303876 489338 303884 489402
rect 303948 489338 303964 489402
rect 304028 489338 304044 489402
rect 304108 489338 304124 489402
rect 304188 489338 304196 489402
rect 303876 489322 304196 489338
rect 303876 489258 303884 489322
rect 303948 489258 303964 489322
rect 304028 489258 304044 489322
rect 304108 489258 304124 489322
rect 304188 489258 304196 489322
rect 303876 489242 304196 489258
rect 303876 489178 303884 489242
rect 303948 489178 303964 489242
rect 304028 489178 304044 489242
rect 304108 489178 304124 489242
rect 304188 489178 304196 489242
rect 303876 486561 304196 489178
rect 303876 486325 303918 486561
rect 304154 486325 304196 486561
rect 303876 479561 304196 486325
rect 303876 479325 303918 479561
rect 304154 479325 304196 479561
rect 303876 473114 304196 479325
rect 303876 473050 303884 473114
rect 303948 473050 303964 473114
rect 304028 473050 304044 473114
rect 304108 473050 304124 473114
rect 304188 473050 304196 473114
rect 303876 473034 304196 473050
rect 303876 472970 303884 473034
rect 303948 472970 303964 473034
rect 304028 472970 304044 473034
rect 304108 472970 304124 473034
rect 304188 472970 304196 473034
rect 303876 472954 304196 472970
rect 303876 472890 303884 472954
rect 303948 472890 303964 472954
rect 304028 472890 304044 472954
rect 304108 472890 304124 472954
rect 304188 472890 304196 472954
rect 303876 472874 304196 472890
rect 303876 472810 303884 472874
rect 303948 472810 303964 472874
rect 304028 472810 304044 472874
rect 304108 472810 304124 472874
rect 304188 472810 304196 472874
rect 303876 472561 304196 472810
rect 303876 472325 303918 472561
rect 304154 472325 304196 472561
rect 303876 465561 304196 472325
rect 303876 465325 303918 465561
rect 304154 465325 304196 465561
rect 303876 458561 304196 465325
rect 303876 458325 303918 458561
rect 304154 458325 304196 458561
rect 303876 452058 304196 458325
rect 303876 451994 303884 452058
rect 303948 451994 303964 452058
rect 304028 451994 304044 452058
rect 304108 451994 304124 452058
rect 304188 451994 304196 452058
rect 303876 451978 304196 451994
rect 303876 451914 303884 451978
rect 303948 451914 303964 451978
rect 304028 451914 304044 451978
rect 304108 451914 304124 451978
rect 304188 451914 304196 451978
rect 303876 451898 304196 451914
rect 303876 451834 303884 451898
rect 303948 451834 303964 451898
rect 304028 451834 304044 451898
rect 304108 451834 304124 451898
rect 304188 451834 304196 451898
rect 303876 451818 304196 451834
rect 303876 451754 303884 451818
rect 303948 451754 303964 451818
rect 304028 451754 304044 451818
rect 304108 451754 304124 451818
rect 304188 451754 304196 451818
rect 303876 451738 304196 451754
rect 303876 451674 303884 451738
rect 303948 451674 303964 451738
rect 304028 451674 304044 451738
rect 304108 451674 304124 451738
rect 304188 451674 304196 451738
rect 303876 451658 304196 451674
rect 303876 451594 303884 451658
rect 303948 451594 303964 451658
rect 304028 451594 304044 451658
rect 304108 451594 304124 451658
rect 304188 451594 304196 451658
rect 303876 451578 304196 451594
rect 303876 451514 303884 451578
rect 303948 451561 303964 451578
rect 304028 451561 304044 451578
rect 304108 451561 304124 451578
rect 304188 451514 304196 451578
rect 303876 451498 303918 451514
rect 304154 451498 304196 451514
rect 303876 451434 303884 451498
rect 304188 451434 304196 451498
rect 303876 451418 303918 451434
rect 304154 451418 304196 451434
rect 303876 451354 303884 451418
rect 304188 451354 304196 451418
rect 303876 451338 303918 451354
rect 304154 451338 304196 451354
rect 303876 451274 303884 451338
rect 303948 451274 303964 451325
rect 304028 451274 304044 451325
rect 304108 451274 304124 451325
rect 304188 451274 304196 451338
rect 303876 444561 304196 451274
rect 303876 444325 303918 444561
rect 304154 444325 304196 444561
rect 303876 437561 304196 444325
rect 303876 437325 303918 437561
rect 304154 437325 304196 437561
rect 303876 430561 304196 437325
rect 303876 430325 303918 430561
rect 304154 430325 304196 430561
rect 303876 423561 304196 430325
rect 303876 423325 303918 423561
rect 304154 423325 304196 423561
rect 303876 416561 304196 423325
rect 303876 416325 303918 416561
rect 304154 416325 304196 416561
rect 303876 410084 304196 416325
rect 303876 410020 303884 410084
rect 303948 410020 303964 410084
rect 304028 410020 304044 410084
rect 304108 410020 304124 410084
rect 304188 410020 304196 410084
rect 303876 410004 304196 410020
rect 303876 409940 303884 410004
rect 303948 409940 303964 410004
rect 304028 409940 304044 410004
rect 304108 409940 304124 410004
rect 304188 409940 304196 410004
rect 303876 409924 304196 409940
rect 303876 409860 303884 409924
rect 303948 409860 303964 409924
rect 304028 409860 304044 409924
rect 304108 409860 304124 409924
rect 304188 409860 304196 409924
rect 303876 409844 304196 409860
rect 303876 409780 303884 409844
rect 303948 409780 303964 409844
rect 304028 409780 304044 409844
rect 304108 409780 304124 409844
rect 304188 409780 304196 409844
rect 303876 409561 304196 409780
rect 303876 409325 303918 409561
rect 304154 409325 304196 409561
rect 303876 402561 304196 409325
rect 303876 402325 303918 402561
rect 304154 402325 304196 402561
rect 303876 395561 304196 402325
rect 303876 395325 303918 395561
rect 304154 395325 304196 395561
rect 303876 389085 304196 395325
rect 303876 389021 303884 389085
rect 303948 389021 303964 389085
rect 304028 389021 304044 389085
rect 304108 389021 304124 389085
rect 304188 389021 304196 389085
rect 303876 389005 304196 389021
rect 303876 388941 303884 389005
rect 303948 388941 303964 389005
rect 304028 388941 304044 389005
rect 304108 388941 304124 389005
rect 304188 388941 304196 389005
rect 303876 388925 304196 388941
rect 303876 388861 303884 388925
rect 303948 388861 303964 388925
rect 304028 388861 304044 388925
rect 304108 388861 304124 388925
rect 304188 388861 304196 388925
rect 303876 388845 304196 388861
rect 303876 388781 303884 388845
rect 303948 388781 303964 388845
rect 304028 388781 304044 388845
rect 304108 388781 304124 388845
rect 304188 388781 304196 388845
rect 303876 388561 304196 388781
rect 303876 388325 303918 388561
rect 304154 388325 304196 388561
rect 303876 387402 304196 388325
rect 303876 387338 303960 387402
rect 304024 387338 304196 387402
rect 303876 381561 304196 387338
rect 303876 381325 303918 381561
rect 304154 381325 304196 381561
rect 303876 374561 304196 381325
rect 303876 374325 303918 374561
rect 304154 374325 304196 374561
rect 303876 368640 304196 374325
rect 309144 705238 309464 706230
rect 309144 705002 309186 705238
rect 309422 705002 309464 705238
rect 309144 704918 309464 705002
rect 309144 704682 309186 704918
rect 309422 704682 309464 704918
rect 309144 695494 309464 704682
rect 309144 695258 309186 695494
rect 309422 695258 309464 695494
rect 309144 688494 309464 695258
rect 309144 688258 309186 688494
rect 309422 688258 309464 688494
rect 309144 681494 309464 688258
rect 309144 681258 309186 681494
rect 309422 681258 309464 681494
rect 309144 674494 309464 681258
rect 309144 674258 309186 674494
rect 309422 674258 309464 674494
rect 309144 667494 309464 674258
rect 309144 667258 309186 667494
rect 309422 667258 309464 667494
rect 309144 660494 309464 667258
rect 309144 660258 309186 660494
rect 309422 660258 309464 660494
rect 309144 653494 309464 660258
rect 309144 653258 309186 653494
rect 309422 653258 309464 653494
rect 309144 646494 309464 653258
rect 309144 646258 309186 646494
rect 309422 646258 309464 646494
rect 309144 639494 309464 646258
rect 309144 639258 309186 639494
rect 309422 639258 309464 639494
rect 309144 632494 309464 639258
rect 309144 632258 309186 632494
rect 309422 632258 309464 632494
rect 309144 625494 309464 632258
rect 309144 625258 309186 625494
rect 309422 625258 309464 625494
rect 309144 618494 309464 625258
rect 309144 618258 309186 618494
rect 309422 618258 309464 618494
rect 309144 611494 309464 618258
rect 309144 611258 309186 611494
rect 309422 611258 309464 611494
rect 309144 604494 309464 611258
rect 309144 604258 309186 604494
rect 309422 604258 309464 604494
rect 309144 597494 309464 604258
rect 309144 597258 309186 597494
rect 309422 597258 309464 597494
rect 309144 590494 309464 597258
rect 309144 590258 309186 590494
rect 309422 590258 309464 590494
rect 309144 583494 309464 590258
rect 309144 583258 309186 583494
rect 309422 583258 309464 583494
rect 309144 576494 309464 583258
rect 309144 576258 309186 576494
rect 309422 576258 309464 576494
rect 309144 569494 309464 576258
rect 309144 569258 309186 569494
rect 309422 569258 309464 569494
rect 309144 562494 309464 569258
rect 309144 562258 309186 562494
rect 309422 562258 309464 562494
rect 309144 555494 309464 562258
rect 309144 555258 309186 555494
rect 309422 555258 309464 555494
rect 309144 548494 309464 555258
rect 309144 548258 309186 548494
rect 309422 548258 309464 548494
rect 309144 541494 309464 548258
rect 309144 541258 309186 541494
rect 309422 541258 309464 541494
rect 309144 534494 309464 541258
rect 309144 534258 309186 534494
rect 309422 534258 309464 534494
rect 309144 527494 309464 534258
rect 309144 527258 309186 527494
rect 309422 527258 309464 527494
rect 309144 520494 309464 527258
rect 309144 520258 309186 520494
rect 309422 520258 309464 520494
rect 309144 513494 309464 520258
rect 309144 513258 309186 513494
rect 309422 513258 309464 513494
rect 309144 506494 309464 513258
rect 309144 506258 309186 506494
rect 309422 506258 309464 506494
rect 309144 499494 309464 506258
rect 309144 499258 309186 499494
rect 309422 499258 309464 499494
rect 309144 492494 309464 499258
rect 309144 492258 309186 492494
rect 309422 492258 309464 492494
rect 309144 485494 309464 492258
rect 309144 485258 309186 485494
rect 309422 485258 309464 485494
rect 309144 478494 309464 485258
rect 309144 478258 309186 478494
rect 309422 478258 309464 478494
rect 309144 472013 309464 478258
rect 309144 471949 309152 472013
rect 309216 471949 309232 472013
rect 309296 471949 309312 472013
rect 309376 471949 309392 472013
rect 309456 471949 309464 472013
rect 309144 471933 309464 471949
rect 309144 471869 309152 471933
rect 309216 471869 309232 471933
rect 309296 471869 309312 471933
rect 309376 471869 309392 471933
rect 309456 471869 309464 471933
rect 309144 471853 309464 471869
rect 309144 471789 309152 471853
rect 309216 471789 309232 471853
rect 309296 471789 309312 471853
rect 309376 471789 309392 471853
rect 309456 471789 309464 471853
rect 309144 471773 309464 471789
rect 309144 471709 309152 471773
rect 309216 471709 309232 471773
rect 309296 471709 309312 471773
rect 309376 471709 309392 471773
rect 309456 471709 309464 471773
rect 309144 471494 309464 471709
rect 309144 471258 309186 471494
rect 309422 471258 309464 471494
rect 309144 464494 309464 471258
rect 309144 464258 309186 464494
rect 309422 464258 309464 464494
rect 309144 457494 309464 464258
rect 309144 457258 309186 457494
rect 309422 457258 309464 457494
rect 309144 450494 309464 457258
rect 309144 450258 309186 450494
rect 309422 450258 309464 450494
rect 309144 443494 309464 450258
rect 309144 443258 309186 443494
rect 309422 443258 309464 443494
rect 309144 436494 309464 443258
rect 309144 436258 309186 436494
rect 309422 436258 309464 436494
rect 309144 429998 309464 436258
rect 309144 429934 309187 429998
rect 309251 429934 309267 429998
rect 309331 429934 309347 429998
rect 309411 429934 309464 429998
rect 309144 429918 309464 429934
rect 309144 429854 309187 429918
rect 309251 429854 309267 429918
rect 309331 429854 309347 429918
rect 309411 429854 309464 429918
rect 309144 429838 309464 429854
rect 309144 429774 309187 429838
rect 309251 429774 309267 429838
rect 309331 429774 309347 429838
rect 309411 429774 309464 429838
rect 309144 429758 309464 429774
rect 309144 429694 309187 429758
rect 309251 429694 309267 429758
rect 309331 429694 309347 429758
rect 309411 429694 309464 429758
rect 309144 429494 309464 429694
rect 309144 429258 309186 429494
rect 309422 429258 309464 429494
rect 309144 422494 309464 429258
rect 309144 422258 309186 422494
rect 309422 422258 309464 422494
rect 309144 415494 309464 422258
rect 309144 415258 309186 415494
rect 309422 415258 309464 415494
rect 309144 408494 309464 415258
rect 309144 408258 309186 408494
rect 309422 408258 309464 408494
rect 309144 401494 309464 408258
rect 309144 401258 309186 401494
rect 309422 401258 309464 401494
rect 309144 394494 309464 401258
rect 309144 394258 309186 394494
rect 309422 394258 309464 394494
rect 309144 387997 309464 394258
rect 309144 387933 309152 387997
rect 309216 387933 309232 387997
rect 309296 387933 309312 387997
rect 309376 387933 309392 387997
rect 309456 387933 309464 387997
rect 309144 387917 309464 387933
rect 309144 387853 309152 387917
rect 309216 387853 309232 387917
rect 309296 387853 309312 387917
rect 309376 387853 309392 387917
rect 309456 387853 309464 387917
rect 309144 387837 309464 387853
rect 309144 387773 309152 387837
rect 309216 387773 309232 387837
rect 309296 387773 309312 387837
rect 309376 387773 309392 387837
rect 309456 387773 309464 387837
rect 309144 387757 309464 387773
rect 309144 387693 309152 387757
rect 309216 387693 309232 387757
rect 309296 387693 309312 387757
rect 309376 387693 309392 387757
rect 309456 387693 309464 387757
rect 309144 387494 309464 387693
rect 309144 387258 309186 387494
rect 309422 387258 309464 387494
rect 309144 380494 309464 387258
rect 309144 380258 309186 380494
rect 309422 380258 309464 380494
rect 309144 373494 309464 380258
rect 309144 373258 309186 373494
rect 309422 373258 309464 373494
rect 309144 368640 309464 373258
rect 310876 706198 311196 706230
rect 310876 705962 310918 706198
rect 311154 705962 311196 706198
rect 310876 705878 311196 705962
rect 310876 705642 310918 705878
rect 311154 705642 311196 705878
rect 310876 696561 311196 705642
rect 310876 696325 310918 696561
rect 311154 696325 311196 696561
rect 310876 689561 311196 696325
rect 310876 689325 310918 689561
rect 311154 689325 311196 689561
rect 310876 682561 311196 689325
rect 310876 682325 310918 682561
rect 311154 682325 311196 682561
rect 310876 675561 311196 682325
rect 310876 675325 310918 675561
rect 311154 675325 311196 675561
rect 310876 668561 311196 675325
rect 310876 668325 310918 668561
rect 311154 668325 311196 668561
rect 310876 661561 311196 668325
rect 310876 661325 310918 661561
rect 311154 661325 311196 661561
rect 310876 654561 311196 661325
rect 310876 654325 310918 654561
rect 311154 654325 311196 654561
rect 310876 647561 311196 654325
rect 310876 647325 310918 647561
rect 311154 647325 311196 647561
rect 310876 640561 311196 647325
rect 310876 640325 310918 640561
rect 311154 640325 311196 640561
rect 310876 633561 311196 640325
rect 310876 633325 310918 633561
rect 311154 633325 311196 633561
rect 310876 626561 311196 633325
rect 310876 626325 310918 626561
rect 311154 626325 311196 626561
rect 310876 619561 311196 626325
rect 310876 619325 310918 619561
rect 311154 619325 311196 619561
rect 310876 612561 311196 619325
rect 310876 612325 310918 612561
rect 311154 612325 311196 612561
rect 310876 605561 311196 612325
rect 310876 605325 310918 605561
rect 311154 605325 311196 605561
rect 310876 598561 311196 605325
rect 310876 598325 310918 598561
rect 311154 598325 311196 598561
rect 310876 591561 311196 598325
rect 310876 591325 310918 591561
rect 311154 591325 311196 591561
rect 310876 584561 311196 591325
rect 310876 584325 310918 584561
rect 311154 584325 311196 584561
rect 310876 577561 311196 584325
rect 310876 577325 310918 577561
rect 311154 577325 311196 577561
rect 310876 570561 311196 577325
rect 310876 570325 310918 570561
rect 311154 570325 311196 570561
rect 310876 563561 311196 570325
rect 310876 563325 310918 563561
rect 311154 563325 311196 563561
rect 310876 556561 311196 563325
rect 310876 556325 310918 556561
rect 311154 556325 311196 556561
rect 310876 549561 311196 556325
rect 310876 549325 310918 549561
rect 311154 549325 311196 549561
rect 310876 542561 311196 549325
rect 310876 542325 310918 542561
rect 311154 542325 311196 542561
rect 310876 535561 311196 542325
rect 310876 535325 310918 535561
rect 311154 535325 311196 535561
rect 310876 528561 311196 535325
rect 310876 528325 310918 528561
rect 311154 528325 311196 528561
rect 310876 521561 311196 528325
rect 310876 521325 310918 521561
rect 311154 521325 311196 521561
rect 310876 514561 311196 521325
rect 310876 514325 310918 514561
rect 311154 514325 311196 514561
rect 310876 507561 311196 514325
rect 310876 507325 310918 507561
rect 311154 507325 311196 507561
rect 310876 500561 311196 507325
rect 310876 500325 310918 500561
rect 311154 500325 311196 500561
rect 310876 493561 311196 500325
rect 310876 493325 310918 493561
rect 311154 493325 311196 493561
rect 310876 491654 311196 493325
rect 310876 491590 310884 491654
rect 310948 491590 310964 491654
rect 311028 491590 311044 491654
rect 311108 491590 311124 491654
rect 311188 491590 311196 491654
rect 310876 491574 311196 491590
rect 310876 491510 310884 491574
rect 310948 491510 310964 491574
rect 311028 491510 311044 491574
rect 311108 491510 311124 491574
rect 311188 491510 311196 491574
rect 310876 491494 311196 491510
rect 310876 491430 310884 491494
rect 310948 491430 310964 491494
rect 311028 491430 311044 491494
rect 311108 491430 311124 491494
rect 311188 491430 311196 491494
rect 310876 491414 311196 491430
rect 310876 491350 310884 491414
rect 310948 491350 310964 491414
rect 311028 491350 311044 491414
rect 311108 491350 311124 491414
rect 311188 491350 311196 491414
rect 310876 489482 311196 491350
rect 310876 489418 310884 489482
rect 310948 489418 310964 489482
rect 311028 489418 311044 489482
rect 311108 489418 311124 489482
rect 311188 489418 311196 489482
rect 310876 489402 311196 489418
rect 310876 489338 310884 489402
rect 310948 489338 310964 489402
rect 311028 489338 311044 489402
rect 311108 489338 311124 489402
rect 311188 489338 311196 489402
rect 310876 489322 311196 489338
rect 310876 489258 310884 489322
rect 310948 489258 310964 489322
rect 311028 489258 311044 489322
rect 311108 489258 311124 489322
rect 311188 489258 311196 489322
rect 310876 489242 311196 489258
rect 310876 489178 310884 489242
rect 310948 489178 310964 489242
rect 311028 489178 311044 489242
rect 311108 489178 311124 489242
rect 311188 489178 311196 489242
rect 310876 486561 311196 489178
rect 310876 486325 310918 486561
rect 311154 486325 311196 486561
rect 310876 479561 311196 486325
rect 310876 479325 310918 479561
rect 311154 479325 311196 479561
rect 310876 473114 311196 479325
rect 310876 473050 310884 473114
rect 310948 473050 310964 473114
rect 311028 473050 311044 473114
rect 311108 473050 311124 473114
rect 311188 473050 311196 473114
rect 310876 473034 311196 473050
rect 310876 472970 310884 473034
rect 310948 472970 310964 473034
rect 311028 472970 311044 473034
rect 311108 472970 311124 473034
rect 311188 472970 311196 473034
rect 310876 472954 311196 472970
rect 310876 472890 310884 472954
rect 310948 472890 310964 472954
rect 311028 472890 311044 472954
rect 311108 472890 311124 472954
rect 311188 472890 311196 472954
rect 310876 472874 311196 472890
rect 310876 472810 310884 472874
rect 310948 472810 310964 472874
rect 311028 472810 311044 472874
rect 311108 472810 311124 472874
rect 311188 472810 311196 472874
rect 310876 472561 311196 472810
rect 310876 472325 310918 472561
rect 311154 472325 311196 472561
rect 310876 465561 311196 472325
rect 310876 465325 310918 465561
rect 311154 465325 311196 465561
rect 310876 458561 311196 465325
rect 310876 458325 310918 458561
rect 311154 458325 311196 458561
rect 310876 452058 311196 458325
rect 310876 451994 310915 452058
rect 310979 451994 310995 452058
rect 311059 451994 311196 452058
rect 310876 451978 311196 451994
rect 310876 451914 310915 451978
rect 310979 451914 310995 451978
rect 311059 451914 311196 451978
rect 310876 451898 311196 451914
rect 310876 451834 310915 451898
rect 310979 451834 310995 451898
rect 311059 451834 311196 451898
rect 310876 451818 311196 451834
rect 310876 451754 310915 451818
rect 310979 451754 310995 451818
rect 311059 451754 311196 451818
rect 310876 451738 311196 451754
rect 310876 451674 310915 451738
rect 310979 451674 310995 451738
rect 311059 451674 311196 451738
rect 310876 451658 311196 451674
rect 310876 451594 310915 451658
rect 310979 451594 310995 451658
rect 311059 451594 311196 451658
rect 310876 451578 311196 451594
rect 310876 451514 310915 451578
rect 310979 451561 310995 451578
rect 311059 451561 311196 451578
rect 310876 451498 310918 451514
rect 310876 451434 310915 451498
rect 310876 451418 310918 451434
rect 310876 451354 310915 451418
rect 310876 451338 310918 451354
rect 310876 451274 310915 451338
rect 311154 451325 311196 451561
rect 310979 451274 310995 451325
rect 311059 451274 311196 451325
rect 310876 450181 311196 451274
rect 310876 450117 310894 450181
rect 310958 450117 310974 450181
rect 311038 450117 311054 450181
rect 311118 450117 311196 450181
rect 310876 450101 311196 450117
rect 310876 450037 310894 450101
rect 310958 450037 310974 450101
rect 311038 450037 311054 450101
rect 311118 450037 311196 450101
rect 310876 450021 311196 450037
rect 310876 449957 310894 450021
rect 310958 449957 310974 450021
rect 311038 449957 311054 450021
rect 311118 449957 311196 450021
rect 310876 449941 311196 449957
rect 310876 449877 310894 449941
rect 310958 449877 310974 449941
rect 311038 449877 311054 449941
rect 311118 449877 311196 449941
rect 310876 449861 311196 449877
rect 310876 449797 310894 449861
rect 310958 449797 310974 449861
rect 311038 449797 311054 449861
rect 311118 449797 311196 449861
rect 310876 449781 311196 449797
rect 310876 449717 310894 449781
rect 310958 449717 310974 449781
rect 311038 449717 311054 449781
rect 311118 449717 311196 449781
rect 310876 449701 311196 449717
rect 310876 449637 310894 449701
rect 310958 449637 310974 449701
rect 311038 449637 311054 449701
rect 311118 449637 311196 449701
rect 310876 444561 311196 449637
rect 310876 444325 310918 444561
rect 311154 444325 311196 444561
rect 310876 437561 311196 444325
rect 310876 437325 310918 437561
rect 311154 437325 311196 437561
rect 310876 430561 311196 437325
rect 310876 430325 310918 430561
rect 311154 430325 311196 430561
rect 310876 423561 311196 430325
rect 310876 423325 310918 423561
rect 311154 423325 311196 423561
rect 310876 416561 311196 423325
rect 310876 416325 310918 416561
rect 311154 416325 311196 416561
rect 310876 410084 311196 416325
rect 310876 410020 310884 410084
rect 310948 410020 310964 410084
rect 311028 410020 311044 410084
rect 311108 410020 311124 410084
rect 311188 410020 311196 410084
rect 310876 410004 311196 410020
rect 310876 409940 310884 410004
rect 310948 409940 310964 410004
rect 311028 409940 311044 410004
rect 311108 409940 311124 410004
rect 311188 409940 311196 410004
rect 310876 409924 311196 409940
rect 310876 409860 310884 409924
rect 310948 409860 310964 409924
rect 311028 409860 311044 409924
rect 311108 409860 311124 409924
rect 311188 409860 311196 409924
rect 310876 409844 311196 409860
rect 310876 409780 310884 409844
rect 310948 409780 310964 409844
rect 311028 409780 311044 409844
rect 311108 409780 311124 409844
rect 311188 409780 311196 409844
rect 310876 409561 311196 409780
rect 310876 409325 310918 409561
rect 311154 409325 311196 409561
rect 310876 407912 311196 409325
rect 310876 407848 310884 407912
rect 310948 407848 310964 407912
rect 311028 407848 311044 407912
rect 311108 407848 311124 407912
rect 311188 407848 311196 407912
rect 310876 407832 311196 407848
rect 310876 407768 310884 407832
rect 310948 407768 310964 407832
rect 311028 407768 311044 407832
rect 311108 407768 311124 407832
rect 311188 407768 311196 407832
rect 310876 407752 311196 407768
rect 310876 407688 310884 407752
rect 310948 407688 310964 407752
rect 311028 407688 311044 407752
rect 311108 407688 311124 407752
rect 311188 407688 311196 407752
rect 310876 407672 311196 407688
rect 310876 407608 310884 407672
rect 310948 407608 310964 407672
rect 311028 407608 311044 407672
rect 311108 407608 311124 407672
rect 311188 407608 311196 407672
rect 310876 402561 311196 407608
rect 310876 402325 310918 402561
rect 311154 402325 311196 402561
rect 310876 395561 311196 402325
rect 310876 395325 310918 395561
rect 311154 395325 311196 395561
rect 310876 389085 311196 395325
rect 310876 389021 310884 389085
rect 310948 389021 310964 389085
rect 311028 389021 311044 389085
rect 311108 389021 311124 389085
rect 311188 389021 311196 389085
rect 310876 389005 311196 389021
rect 310876 388941 310884 389005
rect 310948 388941 310964 389005
rect 311028 388941 311044 389005
rect 311108 388941 311124 389005
rect 311188 388941 311196 389005
rect 310876 388925 311196 388941
rect 310876 388861 310884 388925
rect 310948 388861 310964 388925
rect 311028 388861 311044 388925
rect 311108 388861 311124 388925
rect 311188 388861 311196 388925
rect 310876 388845 311196 388861
rect 310876 388781 310884 388845
rect 310948 388781 310964 388845
rect 311028 388781 311044 388845
rect 311108 388781 311124 388845
rect 311188 388781 311196 388845
rect 310876 388561 311196 388781
rect 310876 388325 310918 388561
rect 311154 388325 311196 388561
rect 310876 387519 311196 388325
rect 310876 387455 311040 387519
rect 311104 387455 311196 387519
rect 310876 381561 311196 387455
rect 310876 381325 310918 381561
rect 311154 381325 311196 381561
rect 310876 374561 311196 381325
rect 310876 374325 310918 374561
rect 311154 374325 311196 374561
rect 310876 368547 311196 374325
rect 316144 705238 316464 706230
rect 316144 705002 316186 705238
rect 316422 705002 316464 705238
rect 316144 704918 316464 705002
rect 316144 704682 316186 704918
rect 316422 704682 316464 704918
rect 316144 695494 316464 704682
rect 316144 695258 316186 695494
rect 316422 695258 316464 695494
rect 316144 688494 316464 695258
rect 316144 688258 316186 688494
rect 316422 688258 316464 688494
rect 316144 681494 316464 688258
rect 316144 681258 316186 681494
rect 316422 681258 316464 681494
rect 316144 674494 316464 681258
rect 316144 674258 316186 674494
rect 316422 674258 316464 674494
rect 316144 667494 316464 674258
rect 316144 667258 316186 667494
rect 316422 667258 316464 667494
rect 316144 660494 316464 667258
rect 316144 660258 316186 660494
rect 316422 660258 316464 660494
rect 316144 653494 316464 660258
rect 316144 653258 316186 653494
rect 316422 653258 316464 653494
rect 316144 646494 316464 653258
rect 316144 646258 316186 646494
rect 316422 646258 316464 646494
rect 316144 639494 316464 646258
rect 316144 639258 316186 639494
rect 316422 639258 316464 639494
rect 316144 632494 316464 639258
rect 316144 632258 316186 632494
rect 316422 632258 316464 632494
rect 316144 625494 316464 632258
rect 316144 625258 316186 625494
rect 316422 625258 316464 625494
rect 316144 618494 316464 625258
rect 316144 618258 316186 618494
rect 316422 618258 316464 618494
rect 316144 611494 316464 618258
rect 316144 611258 316186 611494
rect 316422 611258 316464 611494
rect 316144 604494 316464 611258
rect 316144 604258 316186 604494
rect 316422 604258 316464 604494
rect 316144 597494 316464 604258
rect 316144 597258 316186 597494
rect 316422 597258 316464 597494
rect 316144 590494 316464 597258
rect 316144 590258 316186 590494
rect 316422 590258 316464 590494
rect 316144 583494 316464 590258
rect 316144 583258 316186 583494
rect 316422 583258 316464 583494
rect 316144 576494 316464 583258
rect 316144 576258 316186 576494
rect 316422 576258 316464 576494
rect 316144 569494 316464 576258
rect 316144 569258 316186 569494
rect 316422 569258 316464 569494
rect 316144 562494 316464 569258
rect 316144 562258 316186 562494
rect 316422 562258 316464 562494
rect 316144 555494 316464 562258
rect 316144 555258 316186 555494
rect 316422 555258 316464 555494
rect 316144 548494 316464 555258
rect 316144 548258 316186 548494
rect 316422 548258 316464 548494
rect 316144 541494 316464 548258
rect 316144 541258 316186 541494
rect 316422 541258 316464 541494
rect 316144 534494 316464 541258
rect 316144 534258 316186 534494
rect 316422 534258 316464 534494
rect 316144 527494 316464 534258
rect 316144 527258 316186 527494
rect 316422 527258 316464 527494
rect 316144 520494 316464 527258
rect 316144 520258 316186 520494
rect 316422 520258 316464 520494
rect 316144 513494 316464 520258
rect 316144 513258 316186 513494
rect 316422 513258 316464 513494
rect 316144 506494 316464 513258
rect 316144 506258 316186 506494
rect 316422 506258 316464 506494
rect 316144 499494 316464 506258
rect 316144 499258 316186 499494
rect 316422 499258 316464 499494
rect 316144 492494 316464 499258
rect 316144 492258 316186 492494
rect 316422 492258 316464 492494
rect 316144 485494 316464 492258
rect 316144 485258 316186 485494
rect 316422 485258 316464 485494
rect 316144 478494 316464 485258
rect 316144 478258 316186 478494
rect 316422 478258 316464 478494
rect 316144 471494 316464 478258
rect 316144 471258 316186 471494
rect 316422 471258 316464 471494
rect 316144 464494 316464 471258
rect 316144 464258 316186 464494
rect 316422 464258 316464 464494
rect 316144 457494 316464 464258
rect 316144 457258 316186 457494
rect 316422 457258 316464 457494
rect 316144 450494 316464 457258
rect 316144 450258 316186 450494
rect 316422 450258 316464 450494
rect 316144 443494 316464 450258
rect 316144 443258 316186 443494
rect 316422 443258 316464 443494
rect 316144 436494 316464 443258
rect 316144 436258 316186 436494
rect 316422 436258 316464 436494
rect 316144 429494 316464 436258
rect 316144 429258 316186 429494
rect 316422 429258 316464 429494
rect 316144 422494 316464 429258
rect 316144 422258 316186 422494
rect 316422 422258 316464 422494
rect 316144 415494 316464 422258
rect 316144 415258 316186 415494
rect 316422 415258 316464 415494
rect 316144 408494 316464 415258
rect 316144 408258 316186 408494
rect 316422 408258 316464 408494
rect 316144 401494 316464 408258
rect 316144 401258 316186 401494
rect 316422 401258 316464 401494
rect 316144 394494 316464 401258
rect 316144 394258 316186 394494
rect 316422 394258 316464 394494
rect 316144 387494 316464 394258
rect 316144 387258 316186 387494
rect 316422 387258 316464 387494
rect 316144 380494 316464 387258
rect 316144 380258 316186 380494
rect 316422 380258 316464 380494
rect 316144 373494 316464 380258
rect 316144 373258 316186 373494
rect 316422 373258 316464 373494
rect 289876 367325 289918 367561
rect 290154 367325 290196 367561
rect 289876 360561 290196 367325
rect 316144 366494 316464 373258
rect 316144 366258 316186 366494
rect 316422 366258 316464 366494
rect 289876 360325 289918 360561
rect 290154 360325 290196 360561
rect 289876 353561 290196 360325
rect 289876 353325 289918 353561
rect 290154 353325 290196 353561
rect 289876 346561 290196 353325
rect 289876 346325 289918 346561
rect 290154 346325 290196 346561
rect 289876 339561 290196 346325
rect 289876 339325 289918 339561
rect 290154 339325 290196 339561
rect 289876 332561 290196 339325
rect 289876 332325 289918 332561
rect 290154 332325 290196 332561
rect 289876 325561 290196 332325
rect 289876 325325 289918 325561
rect 290154 325325 290196 325561
rect 289876 318561 290196 325325
rect 289876 318325 289918 318561
rect 290154 318325 290196 318561
rect 289876 311561 290196 318325
rect 289876 311325 289918 311561
rect 290154 311325 290196 311561
rect 289876 304561 290196 311325
rect 289876 304325 289918 304561
rect 290154 304325 290196 304561
rect 289876 297561 290196 304325
rect 289876 297325 289918 297561
rect 290154 297325 290196 297561
rect 289876 290561 290196 297325
rect 289876 290325 289918 290561
rect 290154 290325 290196 290561
rect 289876 283561 290196 290325
rect 289876 283325 289918 283561
rect 290154 283325 290196 283561
rect 289876 276561 290196 283325
rect 289876 276325 289918 276561
rect 290154 276325 290196 276561
rect 289876 269561 290196 276325
rect 289876 269325 289918 269561
rect 290154 269325 290196 269561
rect 289876 262561 290196 269325
rect 289876 262325 289918 262561
rect 290154 262325 290196 262561
rect 289876 255561 290196 262325
rect 289876 255325 289918 255561
rect 290154 255325 290196 255561
rect 289876 248561 290196 255325
rect 289876 248325 289918 248561
rect 290154 248325 290196 248561
rect 289876 241561 290196 248325
rect 289876 241325 289918 241561
rect 290154 241325 290196 241561
rect 289876 234561 290196 241325
rect 289876 234325 289918 234561
rect 290154 234325 290196 234561
rect 289876 227561 290196 234325
rect 289876 227325 289918 227561
rect 290154 227325 290196 227561
rect 289876 220561 290196 227325
rect 289876 220325 289918 220561
rect 290154 220325 290196 220561
rect 289876 213561 290196 220325
rect 289876 213325 289918 213561
rect 290154 213325 290196 213561
rect 289876 206561 290196 213325
rect 289876 206325 289918 206561
rect 290154 206325 290196 206561
rect 289876 199561 290196 206325
rect 295144 359494 295464 364236
rect 295144 359258 295186 359494
rect 295422 359258 295464 359494
rect 295144 352494 295464 359258
rect 295144 352258 295186 352494
rect 295422 352258 295464 352494
rect 295144 345494 295464 352258
rect 295144 345258 295186 345494
rect 295422 345258 295464 345494
rect 295144 338494 295464 345258
rect 295144 338258 295186 338494
rect 295422 338258 295464 338494
rect 295144 331494 295464 338258
rect 295144 331258 295186 331494
rect 295422 331258 295464 331494
rect 295144 324494 295464 331258
rect 295144 324258 295186 324494
rect 295422 324258 295464 324494
rect 295144 317494 295464 324258
rect 295144 317258 295186 317494
rect 295422 317258 295464 317494
rect 295144 310494 295464 317258
rect 295144 310258 295186 310494
rect 295422 310258 295464 310494
rect 295144 303494 295464 310258
rect 295144 303258 295186 303494
rect 295422 303258 295464 303494
rect 295144 296494 295464 303258
rect 295144 296258 295186 296494
rect 295422 296258 295464 296494
rect 295144 289494 295464 296258
rect 295144 289258 295186 289494
rect 295422 289258 295464 289494
rect 295144 282494 295464 289258
rect 295144 282258 295186 282494
rect 295422 282258 295464 282494
rect 295144 275494 295464 282258
rect 295144 275258 295186 275494
rect 295422 275258 295464 275494
rect 295144 268494 295464 275258
rect 295144 268258 295186 268494
rect 295422 268258 295464 268494
rect 295144 261494 295464 268258
rect 295144 261258 295186 261494
rect 295422 261258 295464 261494
rect 295144 254494 295464 261258
rect 295144 254258 295186 254494
rect 295422 254258 295464 254494
rect 295144 247494 295464 254258
rect 295144 247258 295186 247494
rect 295422 247258 295464 247494
rect 295144 240999 295464 247258
rect 295144 240935 295152 240999
rect 295216 240935 295232 240999
rect 295296 240935 295312 240999
rect 295376 240935 295392 240999
rect 295456 240935 295464 240999
rect 295144 240919 295464 240935
rect 295144 240855 295152 240919
rect 295216 240855 295232 240919
rect 295296 240855 295312 240919
rect 295376 240855 295392 240919
rect 295456 240855 295464 240919
rect 295144 240839 295464 240855
rect 295144 240775 295152 240839
rect 295216 240775 295232 240839
rect 295296 240775 295312 240839
rect 295376 240775 295392 240839
rect 295456 240775 295464 240839
rect 295144 240759 295464 240775
rect 295144 240695 295152 240759
rect 295216 240695 295232 240759
rect 295296 240695 295312 240759
rect 295376 240695 295392 240759
rect 295456 240695 295464 240759
rect 295144 240494 295464 240695
rect 295144 240258 295186 240494
rect 295422 240258 295464 240494
rect 295144 233494 295464 240258
rect 295144 233258 295186 233494
rect 295422 233258 295464 233494
rect 295144 226494 295464 233258
rect 295144 226258 295186 226494
rect 295422 226258 295464 226494
rect 295144 220000 295464 226258
rect 295144 219936 295152 220000
rect 295216 219936 295232 220000
rect 295296 219936 295312 220000
rect 295376 219936 295392 220000
rect 295456 219936 295464 220000
rect 295144 219920 295464 219936
rect 295144 219856 295152 219920
rect 295216 219856 295232 219920
rect 295296 219856 295312 219920
rect 295376 219856 295392 219920
rect 295456 219856 295464 219920
rect 295144 219840 295464 219856
rect 295144 219776 295152 219840
rect 295216 219776 295232 219840
rect 295296 219776 295312 219840
rect 295376 219776 295392 219840
rect 295456 219776 295464 219840
rect 295144 219760 295464 219776
rect 295144 219696 295152 219760
rect 295216 219696 295232 219760
rect 295296 219696 295312 219760
rect 295376 219696 295392 219760
rect 295456 219696 295464 219760
rect 295144 219494 295464 219696
rect 295144 219258 295186 219494
rect 295422 219258 295464 219494
rect 295144 212494 295464 219258
rect 295144 212258 295186 212494
rect 295422 212258 295464 212494
rect 295144 205494 295464 212258
rect 295144 205258 295186 205494
rect 295422 205258 295464 205494
rect 295144 200640 295464 205258
rect 296876 360561 297196 364236
rect 296876 360325 296918 360561
rect 297154 360325 297196 360561
rect 296876 353561 297196 360325
rect 296876 353325 296918 353561
rect 297154 353325 297196 353561
rect 296876 347085 297196 353325
rect 296876 347021 296884 347085
rect 296948 347021 296964 347085
rect 297028 347021 297044 347085
rect 297108 347021 297124 347085
rect 297188 347021 297196 347085
rect 296876 347005 297196 347021
rect 296876 346941 296884 347005
rect 296948 346941 296964 347005
rect 297028 346941 297044 347005
rect 297108 346941 297124 347005
rect 297188 346941 297196 347005
rect 296876 346925 297196 346941
rect 296876 346861 296884 346925
rect 296948 346861 296964 346925
rect 297028 346861 297044 346925
rect 297108 346861 297124 346925
rect 297188 346861 297196 346925
rect 296876 346845 297196 346861
rect 296876 346781 296884 346845
rect 296948 346781 296964 346845
rect 297028 346781 297044 346845
rect 297108 346781 297124 346845
rect 297188 346781 297196 346845
rect 296876 346561 297196 346781
rect 296876 346325 296918 346561
rect 297154 346325 297196 346561
rect 296876 339561 297196 346325
rect 296876 339325 296918 339561
rect 297154 339325 297196 339561
rect 296876 332561 297196 339325
rect 296876 332325 296918 332561
rect 297154 332325 297196 332561
rect 296876 326084 297196 332325
rect 296876 326020 296884 326084
rect 296948 326020 296964 326084
rect 297028 326020 297044 326084
rect 297108 326020 297124 326084
rect 297188 326020 297196 326084
rect 296876 326004 297196 326020
rect 296876 325940 296884 326004
rect 296948 325940 296964 326004
rect 297028 325940 297044 326004
rect 297108 325940 297124 326004
rect 297188 325940 297196 326004
rect 296876 325924 297196 325940
rect 296876 325860 296884 325924
rect 296948 325860 296964 325924
rect 297028 325860 297044 325924
rect 297108 325860 297124 325924
rect 297188 325860 297196 325924
rect 296876 325844 297196 325860
rect 296876 325780 296884 325844
rect 296948 325780 296964 325844
rect 297028 325780 297044 325844
rect 297108 325780 297124 325844
rect 297188 325780 297196 325844
rect 296876 325561 297196 325780
rect 296876 325325 296918 325561
rect 297154 325325 297196 325561
rect 296876 318561 297196 325325
rect 296876 318325 296918 318561
rect 297154 318325 297196 318561
rect 296876 311561 297196 318325
rect 296876 311325 296918 311561
rect 297154 311325 297196 311561
rect 296876 305114 297196 311325
rect 296876 305050 296884 305114
rect 296948 305050 296964 305114
rect 297028 305050 297044 305114
rect 297108 305050 297124 305114
rect 297188 305050 297196 305114
rect 296876 305034 297196 305050
rect 296876 304970 296884 305034
rect 296948 304970 296964 305034
rect 297028 304970 297044 305034
rect 297108 304970 297124 305034
rect 297188 304970 297196 305034
rect 296876 304954 297196 304970
rect 296876 304890 296884 304954
rect 296948 304890 296964 304954
rect 297028 304890 297044 304954
rect 297108 304890 297124 304954
rect 297188 304890 297196 304954
rect 296876 304874 297196 304890
rect 296876 304810 296884 304874
rect 296948 304810 296964 304874
rect 297028 304810 297044 304874
rect 297108 304810 297124 304874
rect 297188 304810 297196 304874
rect 296876 304561 297196 304810
rect 296876 304325 296918 304561
rect 297154 304325 297196 304561
rect 296876 297561 297196 304325
rect 296876 297325 296918 297561
rect 297154 297325 297196 297561
rect 296876 290561 297196 297325
rect 296876 290325 296918 290561
rect 297154 290325 297196 290561
rect 296876 283561 297196 290325
rect 296876 283325 296918 283561
rect 297154 283325 297196 283561
rect 296876 276561 297196 283325
rect 296876 276325 296918 276561
rect 297154 276325 297196 276561
rect 296876 269561 297196 276325
rect 296876 269325 296918 269561
rect 297154 269325 297196 269561
rect 296876 262561 297196 269325
rect 296876 262325 296918 262561
rect 297154 262325 297196 262561
rect 296876 255561 297196 262325
rect 296876 255325 296918 255561
rect 297154 255325 297196 255561
rect 296876 248561 297196 255325
rect 296876 248325 296918 248561
rect 297154 248325 297196 248561
rect 296876 242084 297196 248325
rect 296876 242020 296884 242084
rect 296948 242020 296964 242084
rect 297028 242020 297044 242084
rect 297108 242020 297124 242084
rect 297188 242020 297196 242084
rect 296876 242004 297196 242020
rect 296876 241940 296884 242004
rect 296948 241940 296964 242004
rect 297028 241940 297044 242004
rect 297108 241940 297124 242004
rect 297188 241940 297196 242004
rect 296876 241924 297196 241940
rect 296876 241860 296884 241924
rect 296948 241860 296964 241924
rect 297028 241860 297044 241924
rect 297108 241860 297124 241924
rect 297188 241860 297196 241924
rect 296876 241844 297196 241860
rect 296876 241780 296884 241844
rect 296948 241780 296964 241844
rect 297028 241780 297044 241844
rect 297108 241780 297124 241844
rect 297188 241780 297196 241844
rect 296876 241561 297196 241780
rect 296876 241325 296918 241561
rect 297154 241325 297196 241561
rect 296876 234561 297196 241325
rect 296876 234325 296918 234561
rect 297154 234325 297196 234561
rect 296876 227561 297196 234325
rect 296876 227325 296918 227561
rect 297154 227325 297196 227561
rect 296876 221085 297196 227325
rect 296876 221021 296884 221085
rect 296948 221021 296964 221085
rect 297028 221021 297044 221085
rect 297108 221021 297124 221085
rect 297188 221021 297196 221085
rect 296876 221005 297196 221021
rect 296876 220941 296884 221005
rect 296948 220941 296964 221005
rect 297028 220941 297044 221005
rect 297108 220941 297124 221005
rect 297188 220941 297196 221005
rect 296876 220925 297196 220941
rect 296876 220861 296884 220925
rect 296948 220861 296964 220925
rect 297028 220861 297044 220925
rect 297108 220861 297124 220925
rect 297188 220861 297196 220925
rect 296876 220845 297196 220861
rect 296876 220781 296884 220845
rect 296948 220781 296964 220845
rect 297028 220781 297044 220845
rect 297108 220781 297124 220845
rect 297188 220781 297196 220845
rect 296876 220561 297196 220781
rect 296876 220325 296918 220561
rect 297154 220325 297196 220561
rect 296876 213561 297196 220325
rect 296876 213325 296918 213561
rect 297154 213325 297196 213561
rect 296876 206561 297196 213325
rect 296876 206325 296918 206561
rect 297154 206325 297196 206561
rect 296876 200640 297196 206325
rect 302144 359494 302464 364236
rect 302144 359258 302186 359494
rect 302422 359258 302464 359494
rect 302144 352494 302464 359258
rect 302144 352258 302186 352494
rect 302422 352258 302464 352494
rect 302144 345983 302464 352258
rect 302144 345919 302152 345983
rect 302216 345919 302232 345983
rect 302296 345919 302312 345983
rect 302376 345919 302392 345983
rect 302456 345919 302464 345983
rect 302144 345903 302464 345919
rect 302144 345839 302152 345903
rect 302216 345839 302232 345903
rect 302296 345839 302312 345903
rect 302376 345839 302392 345903
rect 302456 345839 302464 345903
rect 302144 345823 302464 345839
rect 302144 345759 302152 345823
rect 302216 345759 302232 345823
rect 302296 345759 302312 345823
rect 302376 345759 302392 345823
rect 302456 345759 302464 345823
rect 302144 345743 302464 345759
rect 302144 345679 302152 345743
rect 302216 345679 302232 345743
rect 302296 345679 302312 345743
rect 302376 345679 302392 345743
rect 302456 345679 302464 345743
rect 302144 345494 302464 345679
rect 302144 345258 302186 345494
rect 302422 345258 302464 345494
rect 302144 338494 302464 345258
rect 302144 338258 302186 338494
rect 302422 338258 302464 338494
rect 302144 331494 302464 338258
rect 302144 331258 302186 331494
rect 302422 331258 302464 331494
rect 302144 324494 302464 331258
rect 302144 324258 302186 324494
rect 302422 324258 302464 324494
rect 302144 317494 302464 324258
rect 302144 317258 302186 317494
rect 302422 317258 302464 317494
rect 302144 310494 302464 317258
rect 302144 310258 302186 310494
rect 302422 310258 302464 310494
rect 302144 304013 302464 310258
rect 302144 303949 302152 304013
rect 302216 303949 302232 304013
rect 302296 303949 302312 304013
rect 302376 303949 302392 304013
rect 302456 303949 302464 304013
rect 302144 303933 302464 303949
rect 302144 303869 302152 303933
rect 302216 303869 302232 303933
rect 302296 303869 302312 303933
rect 302376 303869 302392 303933
rect 302456 303869 302464 303933
rect 302144 303853 302464 303869
rect 302144 303789 302152 303853
rect 302216 303789 302232 303853
rect 302296 303789 302312 303853
rect 302376 303789 302392 303853
rect 302456 303789 302464 303853
rect 302144 303773 302464 303789
rect 302144 303709 302152 303773
rect 302216 303709 302232 303773
rect 302296 303709 302312 303773
rect 302376 303709 302392 303773
rect 302456 303709 302464 303773
rect 302144 303494 302464 303709
rect 302144 303258 302186 303494
rect 302422 303258 302464 303494
rect 302144 296494 302464 303258
rect 302144 296258 302186 296494
rect 302422 296258 302464 296494
rect 302144 289494 302464 296258
rect 302144 289258 302186 289494
rect 302422 289258 302464 289494
rect 302144 282998 302464 289258
rect 302144 282934 302152 282998
rect 302216 282934 302232 282998
rect 302296 282934 302312 282998
rect 302376 282934 302392 282998
rect 302456 282934 302464 282998
rect 302144 282918 302464 282934
rect 302144 282854 302152 282918
rect 302216 282854 302232 282918
rect 302296 282854 302312 282918
rect 302376 282854 302392 282918
rect 302456 282854 302464 282918
rect 302144 282838 302464 282854
rect 302144 282774 302152 282838
rect 302216 282774 302232 282838
rect 302296 282774 302312 282838
rect 302376 282774 302392 282838
rect 302456 282774 302464 282838
rect 302144 282758 302464 282774
rect 302144 282694 302152 282758
rect 302216 282694 302232 282758
rect 302296 282694 302312 282758
rect 302376 282694 302392 282758
rect 302456 282694 302464 282758
rect 302144 282494 302464 282694
rect 302144 282258 302186 282494
rect 302422 282258 302464 282494
rect 302144 275494 302464 282258
rect 302144 275258 302186 275494
rect 302422 275258 302464 275494
rect 302144 268494 302464 275258
rect 302144 268258 302186 268494
rect 302422 268258 302464 268494
rect 302144 261998 302464 268258
rect 302144 261934 302152 261998
rect 302216 261934 302232 261998
rect 302296 261934 302312 261998
rect 302376 261934 302392 261998
rect 302456 261934 302464 261998
rect 302144 261918 302464 261934
rect 302144 261854 302152 261918
rect 302216 261854 302232 261918
rect 302296 261854 302312 261918
rect 302376 261854 302392 261918
rect 302456 261854 302464 261918
rect 302144 261838 302464 261854
rect 302144 261774 302152 261838
rect 302216 261774 302232 261838
rect 302296 261774 302312 261838
rect 302376 261774 302392 261838
rect 302456 261774 302464 261838
rect 302144 261758 302464 261774
rect 302144 261694 302152 261758
rect 302216 261694 302232 261758
rect 302296 261694 302312 261758
rect 302376 261694 302392 261758
rect 302456 261694 302464 261758
rect 302144 261494 302464 261694
rect 302144 261258 302186 261494
rect 302422 261258 302464 261494
rect 302144 254494 302464 261258
rect 302144 254258 302186 254494
rect 302422 254258 302464 254494
rect 302144 247494 302464 254258
rect 302144 247258 302186 247494
rect 302422 247258 302464 247494
rect 302144 240494 302464 247258
rect 302144 240258 302186 240494
rect 302422 240258 302464 240494
rect 302144 233494 302464 240258
rect 302144 233258 302186 233494
rect 302422 233258 302464 233494
rect 302144 226494 302464 233258
rect 302144 226258 302186 226494
rect 302422 226258 302464 226494
rect 302144 219999 302464 226258
rect 302144 219935 302152 219999
rect 302216 219935 302232 219999
rect 302296 219935 302312 219999
rect 302376 219935 302392 219999
rect 302456 219935 302464 219999
rect 302144 219919 302464 219935
rect 302144 219855 302152 219919
rect 302216 219855 302232 219919
rect 302296 219855 302312 219919
rect 302376 219855 302392 219919
rect 302456 219855 302464 219919
rect 302144 219839 302464 219855
rect 302144 219775 302152 219839
rect 302216 219775 302232 219839
rect 302296 219775 302312 219839
rect 302376 219775 302392 219839
rect 302456 219775 302464 219839
rect 302144 219759 302464 219775
rect 302144 219695 302152 219759
rect 302216 219695 302232 219759
rect 302296 219695 302312 219759
rect 302376 219695 302392 219759
rect 302456 219695 302464 219759
rect 302144 219494 302464 219695
rect 302144 219258 302186 219494
rect 302422 219258 302464 219494
rect 302144 212494 302464 219258
rect 302144 212258 302186 212494
rect 302422 212258 302464 212494
rect 302144 205494 302464 212258
rect 302144 205258 302186 205494
rect 302422 205258 302464 205494
rect 302144 200640 302464 205258
rect 303876 360561 304196 364236
rect 303876 360325 303918 360561
rect 304154 360325 304196 360561
rect 303876 353561 304196 360325
rect 303876 353325 303918 353561
rect 304154 353325 304196 353561
rect 303876 347085 304196 353325
rect 303876 347021 303884 347085
rect 303948 347021 303964 347085
rect 304028 347021 304044 347085
rect 304108 347021 304124 347085
rect 304188 347021 304196 347085
rect 303876 347005 304196 347021
rect 303876 346941 303884 347005
rect 303948 346941 303964 347005
rect 304028 346941 304044 347005
rect 304108 346941 304124 347005
rect 304188 346941 304196 347005
rect 303876 346925 304196 346941
rect 303876 346861 303884 346925
rect 303948 346861 303964 346925
rect 304028 346861 304044 346925
rect 304108 346861 304124 346925
rect 304188 346861 304196 346925
rect 303876 346845 304196 346861
rect 303876 346781 303884 346845
rect 303948 346781 303964 346845
rect 304028 346781 304044 346845
rect 304108 346781 304124 346845
rect 304188 346781 304196 346845
rect 303876 346561 304196 346781
rect 303876 346325 303918 346561
rect 304154 346325 304196 346561
rect 303876 339561 304196 346325
rect 303876 339325 303918 339561
rect 304154 339325 304196 339561
rect 303876 332561 304196 339325
rect 303876 332325 303918 332561
rect 304154 332325 304196 332561
rect 303876 326084 304196 332325
rect 303876 326020 303884 326084
rect 303948 326020 303964 326084
rect 304028 326020 304044 326084
rect 304108 326020 304124 326084
rect 304188 326020 304196 326084
rect 303876 326004 304196 326020
rect 303876 325940 303884 326004
rect 303948 325940 303964 326004
rect 304028 325940 304044 326004
rect 304108 325940 304124 326004
rect 304188 325940 304196 326004
rect 303876 325924 304196 325940
rect 303876 325860 303884 325924
rect 303948 325860 303964 325924
rect 304028 325860 304044 325924
rect 304108 325860 304124 325924
rect 304188 325860 304196 325924
rect 303876 325844 304196 325860
rect 303876 325780 303884 325844
rect 303948 325780 303964 325844
rect 304028 325780 304044 325844
rect 304108 325780 304124 325844
rect 304188 325780 304196 325844
rect 303876 325561 304196 325780
rect 303876 325325 303918 325561
rect 304154 325325 304196 325561
rect 303876 323912 304196 325325
rect 303876 323848 303884 323912
rect 303948 323848 303964 323912
rect 304028 323848 304044 323912
rect 304108 323848 304124 323912
rect 304188 323848 304196 323912
rect 303876 323832 304196 323848
rect 303876 323768 303884 323832
rect 303948 323768 303964 323832
rect 304028 323768 304044 323832
rect 304108 323768 304124 323832
rect 304188 323768 304196 323832
rect 303876 323752 304196 323768
rect 303876 323688 303884 323752
rect 303948 323688 303964 323752
rect 304028 323688 304044 323752
rect 304108 323688 304124 323752
rect 304188 323688 304196 323752
rect 303876 323672 304196 323688
rect 303876 323608 303884 323672
rect 303948 323608 303964 323672
rect 304028 323608 304044 323672
rect 304108 323608 304124 323672
rect 304188 323608 304196 323672
rect 303876 318561 304196 323608
rect 303876 318325 303918 318561
rect 304154 318325 304196 318561
rect 303876 311561 304196 318325
rect 303876 311325 303918 311561
rect 304154 311325 304196 311561
rect 303876 305114 304196 311325
rect 303876 305050 303884 305114
rect 303948 305050 303964 305114
rect 304028 305050 304044 305114
rect 304108 305050 304124 305114
rect 304188 305050 304196 305114
rect 303876 305034 304196 305050
rect 303876 304970 303884 305034
rect 303948 304970 303964 305034
rect 304028 304970 304044 305034
rect 304108 304970 304124 305034
rect 304188 304970 304196 305034
rect 303876 304954 304196 304970
rect 303876 304890 303884 304954
rect 303948 304890 303964 304954
rect 304028 304890 304044 304954
rect 304108 304890 304124 304954
rect 304188 304890 304196 304954
rect 303876 304874 304196 304890
rect 303876 304810 303884 304874
rect 303948 304810 303964 304874
rect 304028 304810 304044 304874
rect 304108 304810 304124 304874
rect 304188 304810 304196 304874
rect 303876 304561 304196 304810
rect 303876 304325 303918 304561
rect 304154 304325 304196 304561
rect 303876 297561 304196 304325
rect 303876 297325 303918 297561
rect 304154 297325 304196 297561
rect 303876 290561 304196 297325
rect 303876 290325 303918 290561
rect 304154 290325 304196 290561
rect 303876 283561 304196 290325
rect 303876 283325 303918 283561
rect 304154 283325 304196 283561
rect 303876 282237 304196 283325
rect 303876 282173 303884 282237
rect 303948 282173 303964 282237
rect 304028 282173 304044 282237
rect 304108 282173 304124 282237
rect 304188 282173 304196 282237
rect 303876 282157 304196 282173
rect 303876 282093 303884 282157
rect 303948 282093 303964 282157
rect 304028 282093 304044 282157
rect 304108 282093 304124 282157
rect 304188 282093 304196 282157
rect 303876 282077 304196 282093
rect 303876 282013 303884 282077
rect 303948 282013 303964 282077
rect 304028 282013 304044 282077
rect 304108 282013 304124 282077
rect 304188 282013 304196 282077
rect 303876 281997 304196 282013
rect 303876 281933 303884 281997
rect 303948 281933 303964 281997
rect 304028 281933 304044 281997
rect 304108 281933 304124 281997
rect 304188 281933 304196 281997
rect 303876 281917 304196 281933
rect 303876 281853 303884 281917
rect 303948 281853 303964 281917
rect 304028 281853 304044 281917
rect 304108 281853 304124 281917
rect 304188 281853 304196 281917
rect 303876 281837 304196 281853
rect 303876 281773 303884 281837
rect 303948 281773 303964 281837
rect 304028 281773 304044 281837
rect 304108 281773 304124 281837
rect 304188 281773 304196 281837
rect 303876 281757 304196 281773
rect 303876 281693 303884 281757
rect 303948 281693 303964 281757
rect 304028 281693 304044 281757
rect 304108 281693 304124 281757
rect 304188 281693 304196 281757
rect 303876 281677 304196 281693
rect 303876 281613 303884 281677
rect 303948 281613 303964 281677
rect 304028 281613 304044 281677
rect 304108 281613 304124 281677
rect 304188 281613 304196 281677
rect 303876 276561 304196 281613
rect 303876 276325 303918 276561
rect 304154 276325 304196 276561
rect 303876 269561 304196 276325
rect 303876 269325 303918 269561
rect 304154 269325 304196 269561
rect 303876 262561 304196 269325
rect 303876 262325 303918 262561
rect 304154 262325 304196 262561
rect 303876 261237 304196 262325
rect 303876 261173 303884 261237
rect 303948 261173 303964 261237
rect 304028 261173 304044 261237
rect 304108 261173 304124 261237
rect 304188 261173 304196 261237
rect 303876 261157 304196 261173
rect 303876 261093 303884 261157
rect 303948 261093 303964 261157
rect 304028 261093 304044 261157
rect 304108 261093 304124 261157
rect 304188 261093 304196 261157
rect 303876 261077 304196 261093
rect 303876 261013 303884 261077
rect 303948 261013 303964 261077
rect 304028 261013 304044 261077
rect 304108 261013 304124 261077
rect 304188 261013 304196 261077
rect 303876 260997 304196 261013
rect 303876 260933 303884 260997
rect 303948 260933 303964 260997
rect 304028 260933 304044 260997
rect 304108 260933 304124 260997
rect 304188 260933 304196 260997
rect 303876 260917 304196 260933
rect 303876 260853 303884 260917
rect 303948 260853 303964 260917
rect 304028 260853 304044 260917
rect 304108 260853 304124 260917
rect 304188 260853 304196 260917
rect 303876 260837 304196 260853
rect 303876 260773 303884 260837
rect 303948 260773 303964 260837
rect 304028 260773 304044 260837
rect 304108 260773 304124 260837
rect 304188 260773 304196 260837
rect 303876 260757 304196 260773
rect 303876 260693 303884 260757
rect 303948 260693 303964 260757
rect 304028 260693 304044 260757
rect 304108 260693 304124 260757
rect 304188 260693 304196 260757
rect 303876 260677 304196 260693
rect 303876 260613 303884 260677
rect 303948 260613 303964 260677
rect 304028 260613 304044 260677
rect 304108 260613 304124 260677
rect 304188 260613 304196 260677
rect 303876 255561 304196 260613
rect 303876 255325 303918 255561
rect 304154 255325 304196 255561
rect 303876 248561 304196 255325
rect 303876 248325 303918 248561
rect 304154 248325 304196 248561
rect 303876 242084 304196 248325
rect 303876 242020 303884 242084
rect 303948 242020 303964 242084
rect 304028 242020 304044 242084
rect 304108 242020 304124 242084
rect 304188 242020 304196 242084
rect 303876 242004 304196 242020
rect 303876 241940 303884 242004
rect 303948 241940 303964 242004
rect 304028 241940 304044 242004
rect 304108 241940 304124 242004
rect 304188 241940 304196 242004
rect 303876 241924 304196 241940
rect 303876 241860 303884 241924
rect 303948 241860 303964 241924
rect 304028 241860 304044 241924
rect 304108 241860 304124 241924
rect 304188 241860 304196 241924
rect 303876 241844 304196 241860
rect 303876 241780 303884 241844
rect 303948 241780 303964 241844
rect 304028 241780 304044 241844
rect 304108 241780 304124 241844
rect 304188 241780 304196 241844
rect 303876 241561 304196 241780
rect 303876 241325 303918 241561
rect 304154 241325 304196 241561
rect 303876 234561 304196 241325
rect 303876 234325 303918 234561
rect 304154 234325 304196 234561
rect 303876 227561 304196 234325
rect 303876 227325 303918 227561
rect 304154 227325 304196 227561
rect 303876 221085 304196 227325
rect 303876 221021 303884 221085
rect 303948 221021 303964 221085
rect 304028 221021 304044 221085
rect 304108 221021 304124 221085
rect 304188 221021 304196 221085
rect 303876 221005 304196 221021
rect 303876 220941 303884 221005
rect 303948 220941 303964 221005
rect 304028 220941 304044 221005
rect 304108 220941 304124 221005
rect 304188 220941 304196 221005
rect 303876 220925 304196 220941
rect 303876 220861 303884 220925
rect 303948 220861 303964 220925
rect 304028 220861 304044 220925
rect 304108 220861 304124 220925
rect 304188 220861 304196 220925
rect 303876 220845 304196 220861
rect 303876 220781 303884 220845
rect 303948 220781 303964 220845
rect 304028 220781 304044 220845
rect 304108 220781 304124 220845
rect 304188 220781 304196 220845
rect 303876 220561 304196 220781
rect 303876 220325 303918 220561
rect 304154 220325 304196 220561
rect 303876 219402 304196 220325
rect 303876 219338 303959 219402
rect 304023 219338 304196 219402
rect 303876 213561 304196 219338
rect 303876 213325 303918 213561
rect 304154 213325 304196 213561
rect 303876 206561 304196 213325
rect 303876 206325 303918 206561
rect 304154 206325 304196 206561
rect 303876 200640 304196 206325
rect 309144 359494 309464 364236
rect 309144 359258 309186 359494
rect 309422 359258 309464 359494
rect 309144 352494 309464 359258
rect 309144 352258 309186 352494
rect 309422 352258 309464 352494
rect 309144 345983 309464 352258
rect 309144 345919 309152 345983
rect 309216 345919 309232 345983
rect 309296 345919 309312 345983
rect 309376 345919 309392 345983
rect 309456 345919 309464 345983
rect 309144 345903 309464 345919
rect 309144 345839 309152 345903
rect 309216 345839 309232 345903
rect 309296 345839 309312 345903
rect 309376 345839 309392 345903
rect 309456 345839 309464 345903
rect 309144 345823 309464 345839
rect 309144 345759 309152 345823
rect 309216 345759 309232 345823
rect 309296 345759 309312 345823
rect 309376 345759 309392 345823
rect 309456 345759 309464 345823
rect 309144 345743 309464 345759
rect 309144 345679 309152 345743
rect 309216 345679 309232 345743
rect 309296 345679 309312 345743
rect 309376 345679 309392 345743
rect 309456 345679 309464 345743
rect 309144 345494 309464 345679
rect 309144 345258 309186 345494
rect 309422 345258 309464 345494
rect 309144 338494 309464 345258
rect 309144 338258 309186 338494
rect 309422 338258 309464 338494
rect 309144 331494 309464 338258
rect 309144 331258 309186 331494
rect 309422 331258 309464 331494
rect 309144 324494 309464 331258
rect 309144 324258 309186 324494
rect 309422 324258 309464 324494
rect 309144 317494 309464 324258
rect 309144 317258 309186 317494
rect 309422 317258 309464 317494
rect 309144 310494 309464 317258
rect 309144 310258 309186 310494
rect 309422 310258 309464 310494
rect 309144 304013 309464 310258
rect 309144 303949 309152 304013
rect 309216 303949 309232 304013
rect 309296 303949 309312 304013
rect 309376 303949 309392 304013
rect 309456 303949 309464 304013
rect 309144 303933 309464 303949
rect 309144 303869 309152 303933
rect 309216 303869 309232 303933
rect 309296 303869 309312 303933
rect 309376 303869 309392 303933
rect 309456 303869 309464 303933
rect 309144 303853 309464 303869
rect 309144 303789 309152 303853
rect 309216 303789 309232 303853
rect 309296 303789 309312 303853
rect 309376 303789 309392 303853
rect 309456 303789 309464 303853
rect 309144 303773 309464 303789
rect 309144 303709 309152 303773
rect 309216 303709 309232 303773
rect 309296 303709 309312 303773
rect 309376 303709 309392 303773
rect 309456 303709 309464 303773
rect 309144 303494 309464 303709
rect 309144 303258 309186 303494
rect 309422 303258 309464 303494
rect 309144 296494 309464 303258
rect 309144 296258 309186 296494
rect 309422 296258 309464 296494
rect 309144 289494 309464 296258
rect 309144 289258 309186 289494
rect 309422 289258 309464 289494
rect 309144 282999 309464 289258
rect 309144 282935 309152 282999
rect 309216 282935 309232 282999
rect 309296 282935 309312 282999
rect 309376 282935 309392 282999
rect 309456 282935 309464 282999
rect 309144 282919 309464 282935
rect 309144 282855 309152 282919
rect 309216 282855 309232 282919
rect 309296 282855 309312 282919
rect 309376 282855 309392 282919
rect 309456 282855 309464 282919
rect 309144 282839 309464 282855
rect 309144 282775 309152 282839
rect 309216 282775 309232 282839
rect 309296 282775 309312 282839
rect 309376 282775 309392 282839
rect 309456 282775 309464 282839
rect 309144 282759 309464 282775
rect 309144 282695 309152 282759
rect 309216 282695 309232 282759
rect 309296 282695 309312 282759
rect 309376 282695 309392 282759
rect 309456 282695 309464 282759
rect 309144 282494 309464 282695
rect 309144 282258 309186 282494
rect 309422 282258 309464 282494
rect 309144 275494 309464 282258
rect 309144 275258 309186 275494
rect 309422 275258 309464 275494
rect 309144 268494 309464 275258
rect 309144 268258 309186 268494
rect 309422 268258 309464 268494
rect 309144 261998 309464 268258
rect 309144 261934 309152 261998
rect 309216 261934 309232 261998
rect 309296 261934 309312 261998
rect 309376 261934 309392 261998
rect 309456 261934 309464 261998
rect 309144 261918 309464 261934
rect 309144 261854 309152 261918
rect 309216 261854 309232 261918
rect 309296 261854 309312 261918
rect 309376 261854 309392 261918
rect 309456 261854 309464 261918
rect 309144 261838 309464 261854
rect 309144 261774 309152 261838
rect 309216 261774 309232 261838
rect 309296 261774 309312 261838
rect 309376 261774 309392 261838
rect 309456 261774 309464 261838
rect 309144 261758 309464 261774
rect 309144 261694 309152 261758
rect 309216 261694 309232 261758
rect 309296 261694 309312 261758
rect 309376 261694 309392 261758
rect 309456 261694 309464 261758
rect 309144 261494 309464 261694
rect 309144 261258 309186 261494
rect 309422 261258 309464 261494
rect 309144 254494 309464 261258
rect 309144 254258 309186 254494
rect 309422 254258 309464 254494
rect 309144 247494 309464 254258
rect 309144 247258 309186 247494
rect 309422 247258 309464 247494
rect 309144 240973 309464 247258
rect 309144 240909 309152 240973
rect 309216 240909 309232 240973
rect 309296 240909 309312 240973
rect 309376 240909 309392 240973
rect 309456 240909 309464 240973
rect 309144 240893 309464 240909
rect 309144 240829 309152 240893
rect 309216 240829 309232 240893
rect 309296 240829 309312 240893
rect 309376 240829 309392 240893
rect 309456 240829 309464 240893
rect 309144 240813 309464 240829
rect 309144 240749 309152 240813
rect 309216 240749 309232 240813
rect 309296 240749 309312 240813
rect 309376 240749 309392 240813
rect 309456 240749 309464 240813
rect 309144 240733 309464 240749
rect 309144 240669 309152 240733
rect 309216 240669 309232 240733
rect 309296 240669 309312 240733
rect 309376 240669 309392 240733
rect 309456 240669 309464 240733
rect 309144 240494 309464 240669
rect 309144 240258 309186 240494
rect 309422 240258 309464 240494
rect 309144 233494 309464 240258
rect 309144 233258 309186 233494
rect 309422 233258 309464 233494
rect 309144 226494 309464 233258
rect 309144 226258 309186 226494
rect 309422 226258 309464 226494
rect 309144 219999 309464 226258
rect 309144 219935 309152 219999
rect 309216 219935 309232 219999
rect 309296 219935 309312 219999
rect 309376 219935 309392 219999
rect 309456 219935 309464 219999
rect 309144 219919 309464 219935
rect 309144 219855 309152 219919
rect 309216 219855 309232 219919
rect 309296 219855 309312 219919
rect 309376 219855 309392 219919
rect 309456 219855 309464 219919
rect 309144 219839 309464 219855
rect 309144 219775 309152 219839
rect 309216 219775 309232 219839
rect 309296 219775 309312 219839
rect 309376 219775 309392 219839
rect 309456 219775 309464 219839
rect 309144 219759 309464 219775
rect 309144 219695 309152 219759
rect 309216 219695 309232 219759
rect 309296 219695 309312 219759
rect 309376 219695 309392 219759
rect 309456 219695 309464 219759
rect 309144 219494 309464 219695
rect 309144 219258 309186 219494
rect 309422 219258 309464 219494
rect 309144 212494 309464 219258
rect 309144 212258 309186 212494
rect 309422 212258 309464 212494
rect 309144 205494 309464 212258
rect 309144 205258 309186 205494
rect 309422 205258 309464 205494
rect 309144 200640 309464 205258
rect 310876 360561 311196 364236
rect 310876 360325 310918 360561
rect 311154 360325 311196 360561
rect 310876 353561 311196 360325
rect 310876 353325 310918 353561
rect 311154 353325 311196 353561
rect 310876 346561 311196 353325
rect 310876 346325 310918 346561
rect 311154 346325 311196 346561
rect 310876 339561 311196 346325
rect 310876 339325 310918 339561
rect 311154 339325 311196 339561
rect 310876 332561 311196 339325
rect 310876 332325 310918 332561
rect 311154 332325 311196 332561
rect 310876 326084 311196 332325
rect 310876 326020 310884 326084
rect 310948 326020 310964 326084
rect 311028 326020 311044 326084
rect 311108 326020 311124 326084
rect 311188 326020 311196 326084
rect 310876 326004 311196 326020
rect 310876 325940 310884 326004
rect 310948 325940 310964 326004
rect 311028 325940 311044 326004
rect 311108 325940 311124 326004
rect 311188 325940 311196 326004
rect 310876 325924 311196 325940
rect 310876 325860 310884 325924
rect 310948 325860 310964 325924
rect 311028 325860 311044 325924
rect 311108 325860 311124 325924
rect 311188 325860 311196 325924
rect 310876 325844 311196 325860
rect 310876 325780 310884 325844
rect 310948 325780 310964 325844
rect 311028 325780 311044 325844
rect 311108 325780 311124 325844
rect 311188 325780 311196 325844
rect 310876 325561 311196 325780
rect 310876 325325 310918 325561
rect 311154 325325 311196 325561
rect 310876 323912 311196 325325
rect 310876 323848 310884 323912
rect 310948 323848 310964 323912
rect 311028 323848 311044 323912
rect 311108 323848 311124 323912
rect 311188 323848 311196 323912
rect 310876 323832 311196 323848
rect 310876 323768 310884 323832
rect 310948 323768 310964 323832
rect 311028 323768 311044 323832
rect 311108 323768 311124 323832
rect 311188 323768 311196 323832
rect 310876 323752 311196 323768
rect 310876 323688 310884 323752
rect 310948 323688 310964 323752
rect 311028 323688 311044 323752
rect 311108 323688 311124 323752
rect 311188 323688 311196 323752
rect 310876 323672 311196 323688
rect 310876 323608 310884 323672
rect 310948 323608 310964 323672
rect 311028 323608 311044 323672
rect 311108 323608 311124 323672
rect 311188 323608 311196 323672
rect 310876 318561 311196 323608
rect 310876 318325 310918 318561
rect 311154 318325 311196 318561
rect 310876 311561 311196 318325
rect 310876 311325 310918 311561
rect 311154 311325 311196 311561
rect 310876 305114 311196 311325
rect 310876 305050 310884 305114
rect 310948 305050 310964 305114
rect 311028 305050 311044 305114
rect 311108 305050 311124 305114
rect 311188 305050 311196 305114
rect 310876 305034 311196 305050
rect 310876 304970 310884 305034
rect 310948 304970 310964 305034
rect 311028 304970 311044 305034
rect 311108 304970 311124 305034
rect 311188 304970 311196 305034
rect 310876 304954 311196 304970
rect 310876 304890 310884 304954
rect 310948 304890 310964 304954
rect 311028 304890 311044 304954
rect 311108 304890 311124 304954
rect 311188 304890 311196 304954
rect 310876 304874 311196 304890
rect 310876 304810 310884 304874
rect 310948 304810 310964 304874
rect 311028 304810 311044 304874
rect 311108 304810 311124 304874
rect 311188 304810 311196 304874
rect 310876 304561 311196 304810
rect 310876 304325 310918 304561
rect 311154 304325 311196 304561
rect 310876 297561 311196 304325
rect 310876 297325 310918 297561
rect 311154 297325 311196 297561
rect 310876 290561 311196 297325
rect 310876 290325 310918 290561
rect 311154 290325 311196 290561
rect 310876 283561 311196 290325
rect 310876 283325 310918 283561
rect 311154 283325 311196 283561
rect 310876 282182 311196 283325
rect 310876 282118 310884 282182
rect 310948 282118 310964 282182
rect 311028 282118 311044 282182
rect 311108 282118 311124 282182
rect 311188 282118 311196 282182
rect 310876 282102 311196 282118
rect 310876 282038 310884 282102
rect 310948 282038 310964 282102
rect 311028 282038 311044 282102
rect 311108 282038 311124 282102
rect 311188 282038 311196 282102
rect 310876 282022 311196 282038
rect 310876 281958 310884 282022
rect 310948 281958 310964 282022
rect 311028 281958 311044 282022
rect 311108 281958 311124 282022
rect 311188 281958 311196 282022
rect 310876 281942 311196 281958
rect 310876 281878 310884 281942
rect 310948 281878 310964 281942
rect 311028 281878 311044 281942
rect 311108 281878 311124 281942
rect 311188 281878 311196 281942
rect 310876 281862 311196 281878
rect 310876 281798 310884 281862
rect 310948 281798 310964 281862
rect 311028 281798 311044 281862
rect 311108 281798 311124 281862
rect 311188 281798 311196 281862
rect 310876 281782 311196 281798
rect 310876 281718 310884 281782
rect 310948 281718 310964 281782
rect 311028 281718 311044 281782
rect 311108 281718 311124 281782
rect 311188 281718 311196 281782
rect 310876 281702 311196 281718
rect 310876 281638 310884 281702
rect 310948 281638 310964 281702
rect 311028 281638 311044 281702
rect 311108 281638 311124 281702
rect 311188 281638 311196 281702
rect 310876 276561 311196 281638
rect 310876 276325 310918 276561
rect 311154 276325 311196 276561
rect 310876 269561 311196 276325
rect 310876 269325 310918 269561
rect 311154 269325 311196 269561
rect 310876 262561 311196 269325
rect 310876 262325 310918 262561
rect 311154 262325 311196 262561
rect 310876 255561 311196 262325
rect 310876 255325 310918 255561
rect 311154 255325 311196 255561
rect 310876 248561 311196 255325
rect 310876 248325 310918 248561
rect 311154 248325 311196 248561
rect 310876 242084 311196 248325
rect 310876 242020 310884 242084
rect 310948 242020 310964 242084
rect 311028 242020 311044 242084
rect 311108 242020 311124 242084
rect 311188 242020 311196 242084
rect 310876 242004 311196 242020
rect 310876 241940 310884 242004
rect 310948 241940 310964 242004
rect 311028 241940 311044 242004
rect 311108 241940 311124 242004
rect 311188 241940 311196 242004
rect 310876 241924 311196 241940
rect 310876 241860 310884 241924
rect 310948 241860 310964 241924
rect 311028 241860 311044 241924
rect 311108 241860 311124 241924
rect 311188 241860 311196 241924
rect 310876 241844 311196 241860
rect 310876 241780 310884 241844
rect 310948 241780 310964 241844
rect 311028 241780 311044 241844
rect 311108 241780 311124 241844
rect 311188 241780 311196 241844
rect 310876 241561 311196 241780
rect 310876 241325 310918 241561
rect 311154 241325 311196 241561
rect 310876 239912 311196 241325
rect 310876 239848 310884 239912
rect 310948 239848 310964 239912
rect 311028 239848 311044 239912
rect 311108 239848 311124 239912
rect 311188 239848 311196 239912
rect 310876 239832 311196 239848
rect 310876 239768 310884 239832
rect 310948 239768 310964 239832
rect 311028 239768 311044 239832
rect 311108 239768 311124 239832
rect 311188 239768 311196 239832
rect 310876 239752 311196 239768
rect 310876 239688 310884 239752
rect 310948 239688 310964 239752
rect 311028 239688 311044 239752
rect 311108 239688 311124 239752
rect 311188 239688 311196 239752
rect 310876 239672 311196 239688
rect 310876 239608 310884 239672
rect 310948 239608 310964 239672
rect 311028 239608 311044 239672
rect 311108 239608 311124 239672
rect 311188 239608 311196 239672
rect 310876 234561 311196 239608
rect 310876 234325 310918 234561
rect 311154 234325 311196 234561
rect 310876 227561 311196 234325
rect 310876 227325 310918 227561
rect 311154 227325 311196 227561
rect 310876 221085 311196 227325
rect 310876 221021 310884 221085
rect 310948 221021 310964 221085
rect 311028 221021 311044 221085
rect 311108 221021 311124 221085
rect 311188 221021 311196 221085
rect 310876 221005 311196 221021
rect 310876 220941 310884 221005
rect 310948 220941 310964 221005
rect 311028 220941 311044 221005
rect 311108 220941 311124 221005
rect 311188 220941 311196 221005
rect 310876 220925 311196 220941
rect 310876 220861 310884 220925
rect 310948 220861 310964 220925
rect 311028 220861 311044 220925
rect 311108 220861 311124 220925
rect 311188 220861 311196 220925
rect 310876 220845 311196 220861
rect 310876 220781 310884 220845
rect 310948 220781 310964 220845
rect 311028 220781 311044 220845
rect 311108 220781 311124 220845
rect 311188 220781 311196 220845
rect 310876 220561 311196 220781
rect 310876 220325 310918 220561
rect 311154 220325 311196 220561
rect 310876 219519 311196 220325
rect 310876 219455 311039 219519
rect 311103 219455 311196 219519
rect 310876 213561 311196 219455
rect 310876 213325 310918 213561
rect 311154 213325 311196 213561
rect 310876 206561 311196 213325
rect 310876 206325 310918 206561
rect 311154 206325 311196 206561
rect 310876 200547 311196 206325
rect 316144 359494 316464 366258
rect 316144 359258 316186 359494
rect 316422 359258 316464 359494
rect 316144 352494 316464 359258
rect 316144 352258 316186 352494
rect 316422 352258 316464 352494
rect 316144 345494 316464 352258
rect 316144 345258 316186 345494
rect 316422 345258 316464 345494
rect 316144 338494 316464 345258
rect 316144 338258 316186 338494
rect 316422 338258 316464 338494
rect 316144 331494 316464 338258
rect 316144 331258 316186 331494
rect 316422 331258 316464 331494
rect 316144 324494 316464 331258
rect 316144 324258 316186 324494
rect 316422 324258 316464 324494
rect 316144 317494 316464 324258
rect 316144 317258 316186 317494
rect 316422 317258 316464 317494
rect 316144 310494 316464 317258
rect 316144 310258 316186 310494
rect 316422 310258 316464 310494
rect 316144 303494 316464 310258
rect 316144 303258 316186 303494
rect 316422 303258 316464 303494
rect 316144 296494 316464 303258
rect 316144 296258 316186 296494
rect 316422 296258 316464 296494
rect 316144 289494 316464 296258
rect 316144 289258 316186 289494
rect 316422 289258 316464 289494
rect 316144 282494 316464 289258
rect 316144 282258 316186 282494
rect 316422 282258 316464 282494
rect 316144 275494 316464 282258
rect 316144 275258 316186 275494
rect 316422 275258 316464 275494
rect 316144 268494 316464 275258
rect 316144 268258 316186 268494
rect 316422 268258 316464 268494
rect 316144 261494 316464 268258
rect 316144 261258 316186 261494
rect 316422 261258 316464 261494
rect 316144 254494 316464 261258
rect 316144 254258 316186 254494
rect 316422 254258 316464 254494
rect 316144 247494 316464 254258
rect 316144 247258 316186 247494
rect 316422 247258 316464 247494
rect 316144 240494 316464 247258
rect 316144 240258 316186 240494
rect 316422 240258 316464 240494
rect 316144 233494 316464 240258
rect 316144 233258 316186 233494
rect 316422 233258 316464 233494
rect 316144 226494 316464 233258
rect 316144 226258 316186 226494
rect 316422 226258 316464 226494
rect 316144 219494 316464 226258
rect 316144 219258 316186 219494
rect 316422 219258 316464 219494
rect 316144 212494 316464 219258
rect 316144 212258 316186 212494
rect 316422 212258 316464 212494
rect 316144 205494 316464 212258
rect 316144 205258 316186 205494
rect 316422 205258 316464 205494
rect 289876 199325 289918 199561
rect 290154 199325 290196 199561
rect 289876 192561 290196 199325
rect 316144 198494 316464 205258
rect 316144 198258 316186 198494
rect 316422 198258 316464 198494
rect 289876 192325 289918 192561
rect 290154 192325 290196 192561
rect 289876 185561 290196 192325
rect 289876 185325 289918 185561
rect 290154 185325 290196 185561
rect 289876 178561 290196 185325
rect 289876 178325 289918 178561
rect 290154 178325 290196 178561
rect 289876 171561 290196 178325
rect 289876 171325 289918 171561
rect 290154 171325 290196 171561
rect 289876 164561 290196 171325
rect 289876 164325 289918 164561
rect 290154 164325 290196 164561
rect 289876 157561 290196 164325
rect 289876 157325 289918 157561
rect 290154 157325 290196 157561
rect 289876 150561 290196 157325
rect 289876 150325 289918 150561
rect 290154 150325 290196 150561
rect 289876 143561 290196 150325
rect 289876 143325 289918 143561
rect 290154 143325 290196 143561
rect 289876 136561 290196 143325
rect 289876 136325 289918 136561
rect 290154 136325 290196 136561
rect 289876 129561 290196 136325
rect 289876 129325 289918 129561
rect 290154 129325 290196 129561
rect 289876 122561 290196 129325
rect 289876 122325 289918 122561
rect 290154 122325 290196 122561
rect 289876 115561 290196 122325
rect 289876 115325 289918 115561
rect 290154 115325 290196 115561
rect 289876 108561 290196 115325
rect 289876 108325 289918 108561
rect 290154 108325 290196 108561
rect 289876 101561 290196 108325
rect 289876 101325 289918 101561
rect 290154 101325 290196 101561
rect 289876 94561 290196 101325
rect 289876 94325 289918 94561
rect 290154 94325 290196 94561
rect 289876 87561 290196 94325
rect 289876 87325 289918 87561
rect 290154 87325 290196 87561
rect 289876 80561 290196 87325
rect 289876 80325 289918 80561
rect 290154 80325 290196 80561
rect 289876 73561 290196 80325
rect 289876 73325 289918 73561
rect 290154 73325 290196 73561
rect 289876 66561 290196 73325
rect 289876 66325 289918 66561
rect 290154 66325 290196 66561
rect 289876 59561 290196 66325
rect 289876 59325 289918 59561
rect 290154 59325 290196 59561
rect 289876 52561 290196 59325
rect 289876 52325 289918 52561
rect 290154 52325 290196 52561
rect 289876 45561 290196 52325
rect 289876 45325 289918 45561
rect 290154 45325 290196 45561
rect 289876 38561 290196 45325
rect 289876 38325 289918 38561
rect 290154 38325 290196 38561
rect 289876 31561 290196 38325
rect 289876 31325 289918 31561
rect 290154 31325 290196 31561
rect 289876 24561 290196 31325
rect 289876 24325 289918 24561
rect 290154 24325 290196 24561
rect 289876 17561 290196 24325
rect 289876 17325 289918 17561
rect 290154 17325 290196 17561
rect 289876 10561 290196 17325
rect 289876 10325 289918 10561
rect 290154 10325 290196 10561
rect 289876 3561 290196 10325
rect 289876 3325 289918 3561
rect 290154 3325 290196 3561
rect 289876 -1706 290196 3325
rect 289876 -1942 289918 -1706
rect 290154 -1942 290196 -1706
rect 289876 -2026 290196 -1942
rect 289876 -2262 289918 -2026
rect 290154 -2262 290196 -2026
rect 289876 -2294 290196 -2262
rect 295144 191494 295464 196236
rect 295144 191258 295186 191494
rect 295422 191258 295464 191494
rect 295144 184494 295464 191258
rect 295144 184258 295186 184494
rect 295422 184258 295464 184494
rect 295144 178199 295464 184258
rect 295144 178135 295152 178199
rect 295216 178135 295232 178199
rect 295296 178135 295312 178199
rect 295376 178135 295392 178199
rect 295456 178135 295464 178199
rect 295144 178119 295464 178135
rect 295144 178055 295152 178119
rect 295216 178055 295232 178119
rect 295296 178055 295312 178119
rect 295376 178055 295392 178119
rect 295456 178055 295464 178119
rect 295144 178039 295464 178055
rect 295144 177975 295152 178039
rect 295216 177975 295232 178039
rect 295296 177975 295312 178039
rect 295376 177975 295392 178039
rect 295456 177975 295464 178039
rect 295144 177959 295464 177975
rect 295144 177895 295152 177959
rect 295216 177895 295232 177959
rect 295296 177895 295312 177959
rect 295376 177895 295392 177959
rect 295456 177895 295464 177959
rect 295144 177494 295464 177895
rect 295144 177258 295186 177494
rect 295422 177258 295464 177494
rect 295144 170494 295464 177258
rect 295144 170258 295186 170494
rect 295422 170258 295464 170494
rect 295144 163494 295464 170258
rect 295144 163258 295186 163494
rect 295422 163258 295464 163494
rect 295144 156494 295464 163258
rect 295144 156258 295186 156494
rect 295422 156258 295464 156494
rect 295144 149494 295464 156258
rect 295144 149258 295186 149494
rect 295422 149258 295464 149494
rect 295144 142494 295464 149258
rect 295144 142258 295186 142494
rect 295422 142258 295464 142494
rect 295144 135494 295464 142258
rect 295144 135258 295186 135494
rect 295422 135258 295464 135494
rect 295144 128494 295464 135258
rect 295144 128258 295186 128494
rect 295422 128258 295464 128494
rect 295144 121494 295464 128258
rect 295144 121258 295186 121494
rect 295422 121258 295464 121494
rect 295144 114494 295464 121258
rect 295144 114258 295186 114494
rect 295422 114258 295464 114494
rect 295144 107494 295464 114258
rect 295144 107258 295186 107494
rect 295422 107258 295464 107494
rect 295144 100494 295464 107258
rect 295144 100258 295186 100494
rect 295422 100258 295464 100494
rect 295144 93494 295464 100258
rect 295144 93258 295186 93494
rect 295422 93258 295464 93494
rect 295144 86494 295464 93258
rect 295144 86258 295186 86494
rect 295422 86258 295464 86494
rect 295144 79494 295464 86258
rect 295144 79258 295186 79494
rect 295422 79258 295464 79494
rect 295144 72494 295464 79258
rect 295144 72258 295186 72494
rect 295422 72258 295464 72494
rect 295144 65494 295464 72258
rect 295144 65258 295186 65494
rect 295422 65258 295464 65494
rect 295144 58494 295464 65258
rect 295144 58258 295186 58494
rect 295422 58258 295464 58494
rect 295144 51494 295464 58258
rect 295144 51258 295186 51494
rect 295422 51258 295464 51494
rect 295144 44494 295464 51258
rect 295144 44258 295186 44494
rect 295422 44258 295464 44494
rect 295144 37494 295464 44258
rect 295144 37258 295186 37494
rect 295422 37258 295464 37494
rect 295144 30494 295464 37258
rect 295144 30258 295186 30494
rect 295422 30258 295464 30494
rect 295144 23494 295464 30258
rect 295144 23258 295186 23494
rect 295422 23258 295464 23494
rect 295144 16494 295464 23258
rect 295144 16258 295186 16494
rect 295422 16258 295464 16494
rect 295144 9494 295464 16258
rect 295144 9258 295186 9494
rect 295422 9258 295464 9494
rect 295144 2494 295464 9258
rect 295144 2258 295186 2494
rect 295422 2258 295464 2494
rect 295144 -746 295464 2258
rect 295144 -982 295186 -746
rect 295422 -982 295464 -746
rect 295144 -1066 295464 -982
rect 295144 -1302 295186 -1066
rect 295422 -1302 295464 -1066
rect 295144 -2294 295464 -1302
rect 296876 192561 297196 196236
rect 296876 192325 296918 192561
rect 297154 192325 297196 192561
rect 296876 185561 297196 192325
rect 296876 185325 296918 185561
rect 297154 185325 297196 185561
rect 296876 179285 297196 185325
rect 296876 179221 296884 179285
rect 296948 179221 296964 179285
rect 297028 179221 297044 179285
rect 297108 179221 297124 179285
rect 297188 179221 297196 179285
rect 296876 179205 297196 179221
rect 296876 179141 296884 179205
rect 296948 179141 296964 179205
rect 297028 179141 297044 179205
rect 297108 179141 297124 179205
rect 297188 179141 297196 179205
rect 296876 179125 297196 179141
rect 296876 179061 296884 179125
rect 296948 179061 296964 179125
rect 297028 179061 297044 179125
rect 297108 179061 297124 179125
rect 297188 179061 297196 179125
rect 296876 179045 297196 179061
rect 296876 178981 296884 179045
rect 296948 178981 296964 179045
rect 297028 178981 297044 179045
rect 297108 178981 297124 179045
rect 297188 178981 297196 179045
rect 296876 178561 297196 178981
rect 296876 178325 296918 178561
rect 297154 178325 297196 178561
rect 296876 171561 297196 178325
rect 296876 171325 296918 171561
rect 297154 171325 297196 171561
rect 296876 164561 297196 171325
rect 296876 164325 296918 164561
rect 297154 164325 297196 164561
rect 296876 157561 297196 164325
rect 296876 157325 296918 157561
rect 297154 157325 297196 157561
rect 296876 150561 297196 157325
rect 296876 150325 296918 150561
rect 297154 150325 297196 150561
rect 296876 143561 297196 150325
rect 296876 143325 296918 143561
rect 297154 143325 297196 143561
rect 296876 136561 297196 143325
rect 296876 136325 296918 136561
rect 297154 136325 297196 136561
rect 296876 129561 297196 136325
rect 296876 129325 296918 129561
rect 297154 129325 297196 129561
rect 296876 122561 297196 129325
rect 296876 122325 296918 122561
rect 297154 122325 297196 122561
rect 296876 115561 297196 122325
rect 296876 115325 296918 115561
rect 297154 115325 297196 115561
rect 296876 108561 297196 115325
rect 296876 108325 296918 108561
rect 297154 108325 297196 108561
rect 296876 101561 297196 108325
rect 296876 101325 296918 101561
rect 297154 101325 297196 101561
rect 296876 94561 297196 101325
rect 296876 94325 296918 94561
rect 297154 94325 297196 94561
rect 296876 87561 297196 94325
rect 296876 87325 296918 87561
rect 297154 87325 297196 87561
rect 296876 80561 297196 87325
rect 296876 80325 296918 80561
rect 297154 80325 297196 80561
rect 296876 73561 297196 80325
rect 296876 73325 296918 73561
rect 297154 73325 297196 73561
rect 296876 66561 297196 73325
rect 296876 66325 296918 66561
rect 297154 66325 297196 66561
rect 296876 59561 297196 66325
rect 296876 59325 296918 59561
rect 297154 59325 297196 59561
rect 296876 52561 297196 59325
rect 296876 52325 296918 52561
rect 297154 52325 297196 52561
rect 296876 45561 297196 52325
rect 296876 45325 296918 45561
rect 297154 45325 297196 45561
rect 296876 38561 297196 45325
rect 296876 38325 296918 38561
rect 297154 38325 297196 38561
rect 296876 31561 297196 38325
rect 296876 31325 296918 31561
rect 297154 31325 297196 31561
rect 296876 24561 297196 31325
rect 296876 24325 296918 24561
rect 297154 24325 297196 24561
rect 296876 17561 297196 24325
rect 296876 17325 296918 17561
rect 297154 17325 297196 17561
rect 296876 10561 297196 17325
rect 296876 10325 296918 10561
rect 297154 10325 297196 10561
rect 296876 3561 297196 10325
rect 296876 3325 296918 3561
rect 297154 3325 297196 3561
rect 296876 -1706 297196 3325
rect 296876 -1942 296918 -1706
rect 297154 -1942 297196 -1706
rect 296876 -2026 297196 -1942
rect 296876 -2262 296918 -2026
rect 297154 -2262 297196 -2026
rect 296876 -2294 297196 -2262
rect 302144 191494 302464 196236
rect 302144 191258 302186 191494
rect 302422 191258 302464 191494
rect 302144 184494 302464 191258
rect 302144 184258 302186 184494
rect 302422 184258 302464 184494
rect 302144 178183 302464 184258
rect 302144 178119 302152 178183
rect 302216 178119 302232 178183
rect 302296 178119 302312 178183
rect 302376 178119 302392 178183
rect 302456 178119 302464 178183
rect 302144 178103 302464 178119
rect 302144 178039 302152 178103
rect 302216 178039 302232 178103
rect 302296 178039 302312 178103
rect 302376 178039 302392 178103
rect 302456 178039 302464 178103
rect 302144 178023 302464 178039
rect 302144 177959 302152 178023
rect 302216 177959 302232 178023
rect 302296 177959 302312 178023
rect 302376 177959 302392 178023
rect 302456 177959 302464 178023
rect 302144 177943 302464 177959
rect 302144 177879 302152 177943
rect 302216 177879 302232 177943
rect 302296 177879 302312 177943
rect 302376 177879 302392 177943
rect 302456 177879 302464 177943
rect 302144 177494 302464 177879
rect 302144 177258 302186 177494
rect 302422 177258 302464 177494
rect 302144 170494 302464 177258
rect 302144 170258 302186 170494
rect 302422 170258 302464 170494
rect 302144 163494 302464 170258
rect 302144 163258 302186 163494
rect 302422 163258 302464 163494
rect 302144 156494 302464 163258
rect 302144 156258 302186 156494
rect 302422 156258 302464 156494
rect 302144 149494 302464 156258
rect 302144 149258 302186 149494
rect 302422 149258 302464 149494
rect 302144 142494 302464 149258
rect 302144 142258 302186 142494
rect 302422 142258 302464 142494
rect 302144 135494 302464 142258
rect 302144 135258 302186 135494
rect 302422 135258 302464 135494
rect 302144 128494 302464 135258
rect 302144 128258 302186 128494
rect 302422 128258 302464 128494
rect 302144 121494 302464 128258
rect 302144 121258 302186 121494
rect 302422 121258 302464 121494
rect 302144 114494 302464 121258
rect 302144 114258 302186 114494
rect 302422 114258 302464 114494
rect 302144 107494 302464 114258
rect 302144 107258 302186 107494
rect 302422 107258 302464 107494
rect 302144 100494 302464 107258
rect 302144 100258 302186 100494
rect 302422 100258 302464 100494
rect 302144 93494 302464 100258
rect 302144 93258 302186 93494
rect 302422 93258 302464 93494
rect 302144 86494 302464 93258
rect 302144 86258 302186 86494
rect 302422 86258 302464 86494
rect 302144 79494 302464 86258
rect 302144 79258 302186 79494
rect 302422 79258 302464 79494
rect 302144 72494 302464 79258
rect 302144 72258 302186 72494
rect 302422 72258 302464 72494
rect 302144 65494 302464 72258
rect 302144 65258 302186 65494
rect 302422 65258 302464 65494
rect 302144 58494 302464 65258
rect 302144 58258 302186 58494
rect 302422 58258 302464 58494
rect 302144 51494 302464 58258
rect 302144 51258 302186 51494
rect 302422 51258 302464 51494
rect 302144 44494 302464 51258
rect 302144 44258 302186 44494
rect 302422 44258 302464 44494
rect 302144 37494 302464 44258
rect 302144 37258 302186 37494
rect 302422 37258 302464 37494
rect 302144 30494 302464 37258
rect 302144 30258 302186 30494
rect 302422 30258 302464 30494
rect 302144 23494 302464 30258
rect 302144 23258 302186 23494
rect 302422 23258 302464 23494
rect 302144 16494 302464 23258
rect 302144 16258 302186 16494
rect 302422 16258 302464 16494
rect 302144 9494 302464 16258
rect 302144 9258 302186 9494
rect 302422 9258 302464 9494
rect 302144 2494 302464 9258
rect 302144 2258 302186 2494
rect 302422 2258 302464 2494
rect 302144 -746 302464 2258
rect 302144 -982 302186 -746
rect 302422 -982 302464 -746
rect 302144 -1066 302464 -982
rect 302144 -1302 302186 -1066
rect 302422 -1302 302464 -1066
rect 302144 -2294 302464 -1302
rect 303876 192561 304196 196236
rect 303876 192325 303918 192561
rect 304154 192325 304196 192561
rect 303876 185561 304196 192325
rect 303876 185325 303918 185561
rect 304154 185325 304196 185561
rect 303876 179285 304196 185325
rect 303876 179221 303884 179285
rect 303948 179221 303964 179285
rect 304028 179221 304044 179285
rect 304108 179221 304124 179285
rect 304188 179221 304196 179285
rect 303876 179205 304196 179221
rect 303876 179141 303884 179205
rect 303948 179141 303964 179205
rect 304028 179141 304044 179205
rect 304108 179141 304124 179205
rect 304188 179141 304196 179205
rect 303876 179125 304196 179141
rect 303876 179061 303884 179125
rect 303948 179061 303964 179125
rect 304028 179061 304044 179125
rect 304108 179061 304124 179125
rect 304188 179061 304196 179125
rect 303876 179045 304196 179061
rect 303876 178981 303884 179045
rect 303948 178981 303964 179045
rect 304028 178981 304044 179045
rect 304108 178981 304124 179045
rect 304188 178981 304196 179045
rect 303876 178561 304196 178981
rect 303876 178325 303918 178561
rect 304154 178325 304196 178561
rect 303876 171561 304196 178325
rect 303876 171325 303918 171561
rect 304154 171325 304196 171561
rect 303876 164561 304196 171325
rect 303876 164325 303918 164561
rect 304154 164325 304196 164561
rect 303876 157561 304196 164325
rect 303876 157325 303918 157561
rect 304154 157325 304196 157561
rect 303876 150561 304196 157325
rect 303876 150325 303918 150561
rect 304154 150325 304196 150561
rect 303876 143561 304196 150325
rect 303876 143325 303918 143561
rect 304154 143325 304196 143561
rect 303876 136561 304196 143325
rect 303876 136325 303918 136561
rect 304154 136325 304196 136561
rect 303876 129561 304196 136325
rect 303876 129325 303918 129561
rect 304154 129325 304196 129561
rect 303876 122561 304196 129325
rect 303876 122325 303918 122561
rect 304154 122325 304196 122561
rect 303876 115561 304196 122325
rect 303876 115325 303918 115561
rect 304154 115325 304196 115561
rect 303876 108561 304196 115325
rect 303876 108325 303918 108561
rect 304154 108325 304196 108561
rect 303876 101561 304196 108325
rect 303876 101325 303918 101561
rect 304154 101325 304196 101561
rect 303876 94561 304196 101325
rect 303876 94325 303918 94561
rect 304154 94325 304196 94561
rect 303876 87561 304196 94325
rect 303876 87325 303918 87561
rect 304154 87325 304196 87561
rect 303876 80561 304196 87325
rect 303876 80325 303918 80561
rect 304154 80325 304196 80561
rect 303876 73561 304196 80325
rect 303876 73325 303918 73561
rect 304154 73325 304196 73561
rect 303876 66561 304196 73325
rect 303876 66325 303918 66561
rect 304154 66325 304196 66561
rect 303876 59561 304196 66325
rect 303876 59325 303918 59561
rect 304154 59325 304196 59561
rect 303876 52561 304196 59325
rect 303876 52325 303918 52561
rect 304154 52325 304196 52561
rect 303876 45561 304196 52325
rect 303876 45325 303918 45561
rect 304154 45325 304196 45561
rect 303876 38561 304196 45325
rect 303876 38325 303918 38561
rect 304154 38325 304196 38561
rect 303876 31561 304196 38325
rect 303876 31325 303918 31561
rect 304154 31325 304196 31561
rect 303876 24561 304196 31325
rect 303876 24325 303918 24561
rect 304154 24325 304196 24561
rect 303876 17561 304196 24325
rect 303876 17325 303918 17561
rect 304154 17325 304196 17561
rect 303876 10561 304196 17325
rect 303876 10325 303918 10561
rect 304154 10325 304196 10561
rect 303876 3561 304196 10325
rect 303876 3325 303918 3561
rect 304154 3325 304196 3561
rect 303876 -1706 304196 3325
rect 303876 -1942 303918 -1706
rect 304154 -1942 304196 -1706
rect 303876 -2026 304196 -1942
rect 303876 -2262 303918 -2026
rect 304154 -2262 304196 -2026
rect 303876 -2294 304196 -2262
rect 309144 191494 309464 196236
rect 309144 191258 309186 191494
rect 309422 191258 309464 191494
rect 309144 184494 309464 191258
rect 309144 184258 309186 184494
rect 309422 184258 309464 184494
rect 309144 178183 309464 184258
rect 309144 178119 309152 178183
rect 309216 178119 309232 178183
rect 309296 178119 309312 178183
rect 309376 178119 309392 178183
rect 309456 178119 309464 178183
rect 309144 178103 309464 178119
rect 309144 178039 309152 178103
rect 309216 178039 309232 178103
rect 309296 178039 309312 178103
rect 309376 178039 309392 178103
rect 309456 178039 309464 178103
rect 309144 178023 309464 178039
rect 309144 177959 309152 178023
rect 309216 177959 309232 178023
rect 309296 177959 309312 178023
rect 309376 177959 309392 178023
rect 309456 177959 309464 178023
rect 309144 177943 309464 177959
rect 309144 177879 309152 177943
rect 309216 177879 309232 177943
rect 309296 177879 309312 177943
rect 309376 177879 309392 177943
rect 309456 177879 309464 177943
rect 309144 177494 309464 177879
rect 309144 177258 309186 177494
rect 309422 177258 309464 177494
rect 309144 170494 309464 177258
rect 309144 170258 309186 170494
rect 309422 170258 309464 170494
rect 309144 163494 309464 170258
rect 309144 163258 309186 163494
rect 309422 163258 309464 163494
rect 309144 156494 309464 163258
rect 309144 156258 309186 156494
rect 309422 156258 309464 156494
rect 309144 149494 309464 156258
rect 309144 149258 309186 149494
rect 309422 149258 309464 149494
rect 309144 142494 309464 149258
rect 309144 142258 309186 142494
rect 309422 142258 309464 142494
rect 309144 135494 309464 142258
rect 309144 135258 309186 135494
rect 309422 135258 309464 135494
rect 309144 128494 309464 135258
rect 309144 128258 309186 128494
rect 309422 128258 309464 128494
rect 309144 121494 309464 128258
rect 309144 121258 309186 121494
rect 309422 121258 309464 121494
rect 309144 114494 309464 121258
rect 309144 114258 309186 114494
rect 309422 114258 309464 114494
rect 309144 107494 309464 114258
rect 309144 107258 309186 107494
rect 309422 107258 309464 107494
rect 309144 100494 309464 107258
rect 309144 100258 309186 100494
rect 309422 100258 309464 100494
rect 309144 93494 309464 100258
rect 309144 93258 309186 93494
rect 309422 93258 309464 93494
rect 309144 86494 309464 93258
rect 309144 86258 309186 86494
rect 309422 86258 309464 86494
rect 309144 79494 309464 86258
rect 309144 79258 309186 79494
rect 309422 79258 309464 79494
rect 309144 72494 309464 79258
rect 309144 72258 309186 72494
rect 309422 72258 309464 72494
rect 309144 65494 309464 72258
rect 309144 65258 309186 65494
rect 309422 65258 309464 65494
rect 309144 58494 309464 65258
rect 309144 58258 309186 58494
rect 309422 58258 309464 58494
rect 309144 51494 309464 58258
rect 309144 51258 309186 51494
rect 309422 51258 309464 51494
rect 309144 44494 309464 51258
rect 309144 44258 309186 44494
rect 309422 44258 309464 44494
rect 309144 37494 309464 44258
rect 309144 37258 309186 37494
rect 309422 37258 309464 37494
rect 309144 30494 309464 37258
rect 309144 30258 309186 30494
rect 309422 30258 309464 30494
rect 309144 23494 309464 30258
rect 309144 23258 309186 23494
rect 309422 23258 309464 23494
rect 309144 16494 309464 23258
rect 309144 16258 309186 16494
rect 309422 16258 309464 16494
rect 309144 9494 309464 16258
rect 309144 9258 309186 9494
rect 309422 9258 309464 9494
rect 309144 2494 309464 9258
rect 309144 2258 309186 2494
rect 309422 2258 309464 2494
rect 309144 -746 309464 2258
rect 309144 -982 309186 -746
rect 309422 -982 309464 -746
rect 309144 -1066 309464 -982
rect 309144 -1302 309186 -1066
rect 309422 -1302 309464 -1066
rect 309144 -2294 309464 -1302
rect 310876 192561 311196 196236
rect 310876 192325 310918 192561
rect 311154 192325 311196 192561
rect 310876 185561 311196 192325
rect 310876 185325 310918 185561
rect 311154 185325 311196 185561
rect 310876 179285 311196 185325
rect 310876 179221 310888 179285
rect 310952 179221 311196 179285
rect 310876 179205 311196 179221
rect 310876 179141 310888 179205
rect 310952 179141 311196 179205
rect 310876 179125 311196 179141
rect 310876 179061 310888 179125
rect 310952 179061 311196 179125
rect 310876 179045 311196 179061
rect 310876 178981 310888 179045
rect 310952 178981 311196 179045
rect 310876 178561 311196 178981
rect 310876 178325 310918 178561
rect 311154 178325 311196 178561
rect 310876 171561 311196 178325
rect 310876 171325 310918 171561
rect 311154 171325 311196 171561
rect 310876 164561 311196 171325
rect 310876 164325 310918 164561
rect 311154 164325 311196 164561
rect 310876 157561 311196 164325
rect 310876 157325 310918 157561
rect 311154 157325 311196 157561
rect 310876 150561 311196 157325
rect 310876 150325 310918 150561
rect 311154 150325 311196 150561
rect 310876 143561 311196 150325
rect 310876 143325 310918 143561
rect 311154 143325 311196 143561
rect 310876 136561 311196 143325
rect 310876 136325 310918 136561
rect 311154 136325 311196 136561
rect 310876 129561 311196 136325
rect 310876 129325 310918 129561
rect 311154 129325 311196 129561
rect 310876 122561 311196 129325
rect 310876 122325 310918 122561
rect 311154 122325 311196 122561
rect 310876 115561 311196 122325
rect 310876 115325 310918 115561
rect 311154 115325 311196 115561
rect 310876 108561 311196 115325
rect 310876 108325 310918 108561
rect 311154 108325 311196 108561
rect 310876 101561 311196 108325
rect 310876 101325 310918 101561
rect 311154 101325 311196 101561
rect 310876 94561 311196 101325
rect 310876 94325 310918 94561
rect 311154 94325 311196 94561
rect 310876 87561 311196 94325
rect 310876 87325 310918 87561
rect 311154 87325 311196 87561
rect 310876 80561 311196 87325
rect 310876 80325 310918 80561
rect 311154 80325 311196 80561
rect 310876 73561 311196 80325
rect 310876 73325 310918 73561
rect 311154 73325 311196 73561
rect 310876 66561 311196 73325
rect 310876 66325 310918 66561
rect 311154 66325 311196 66561
rect 310876 59561 311196 66325
rect 310876 59325 310918 59561
rect 311154 59325 311196 59561
rect 310876 52561 311196 59325
rect 310876 52325 310918 52561
rect 311154 52325 311196 52561
rect 310876 45561 311196 52325
rect 310876 45325 310918 45561
rect 311154 45325 311196 45561
rect 310876 38561 311196 45325
rect 310876 38325 310918 38561
rect 311154 38325 311196 38561
rect 310876 31561 311196 38325
rect 310876 31325 310918 31561
rect 311154 31325 311196 31561
rect 310876 24561 311196 31325
rect 310876 24325 310918 24561
rect 311154 24325 311196 24561
rect 310876 17561 311196 24325
rect 310876 17325 310918 17561
rect 311154 17325 311196 17561
rect 310876 10561 311196 17325
rect 310876 10325 310918 10561
rect 311154 10325 311196 10561
rect 310876 3561 311196 10325
rect 310876 3325 310918 3561
rect 311154 3325 311196 3561
rect 310876 -1706 311196 3325
rect 310876 -1942 310918 -1706
rect 311154 -1942 311196 -1706
rect 310876 -2026 311196 -1942
rect 310876 -2262 310918 -2026
rect 311154 -2262 311196 -2026
rect 310876 -2294 311196 -2262
rect 316144 191494 316464 198258
rect 316144 191258 316186 191494
rect 316422 191258 316464 191494
rect 316144 184494 316464 191258
rect 316144 184258 316186 184494
rect 316422 184258 316464 184494
rect 316144 177494 316464 184258
rect 316144 177258 316186 177494
rect 316422 177258 316464 177494
rect 316144 170494 316464 177258
rect 316144 170258 316186 170494
rect 316422 170258 316464 170494
rect 316144 163494 316464 170258
rect 316144 163258 316186 163494
rect 316422 163258 316464 163494
rect 316144 156494 316464 163258
rect 316144 156258 316186 156494
rect 316422 156258 316464 156494
rect 316144 149494 316464 156258
rect 316144 149258 316186 149494
rect 316422 149258 316464 149494
rect 316144 142494 316464 149258
rect 316144 142258 316186 142494
rect 316422 142258 316464 142494
rect 316144 135494 316464 142258
rect 316144 135258 316186 135494
rect 316422 135258 316464 135494
rect 316144 128494 316464 135258
rect 316144 128258 316186 128494
rect 316422 128258 316464 128494
rect 316144 121494 316464 128258
rect 316144 121258 316186 121494
rect 316422 121258 316464 121494
rect 316144 114494 316464 121258
rect 316144 114258 316186 114494
rect 316422 114258 316464 114494
rect 316144 107494 316464 114258
rect 316144 107258 316186 107494
rect 316422 107258 316464 107494
rect 316144 100494 316464 107258
rect 316144 100258 316186 100494
rect 316422 100258 316464 100494
rect 316144 93494 316464 100258
rect 316144 93258 316186 93494
rect 316422 93258 316464 93494
rect 316144 86494 316464 93258
rect 316144 86258 316186 86494
rect 316422 86258 316464 86494
rect 316144 79494 316464 86258
rect 316144 79258 316186 79494
rect 316422 79258 316464 79494
rect 316144 72494 316464 79258
rect 316144 72258 316186 72494
rect 316422 72258 316464 72494
rect 316144 65494 316464 72258
rect 316144 65258 316186 65494
rect 316422 65258 316464 65494
rect 316144 58494 316464 65258
rect 316144 58258 316186 58494
rect 316422 58258 316464 58494
rect 316144 51494 316464 58258
rect 316144 51258 316186 51494
rect 316422 51258 316464 51494
rect 316144 44494 316464 51258
rect 316144 44258 316186 44494
rect 316422 44258 316464 44494
rect 316144 37494 316464 44258
rect 316144 37258 316186 37494
rect 316422 37258 316464 37494
rect 316144 30494 316464 37258
rect 316144 30258 316186 30494
rect 316422 30258 316464 30494
rect 316144 23494 316464 30258
rect 316144 23258 316186 23494
rect 316422 23258 316464 23494
rect 316144 16494 316464 23258
rect 316144 16258 316186 16494
rect 316422 16258 316464 16494
rect 316144 9494 316464 16258
rect 316144 9258 316186 9494
rect 316422 9258 316464 9494
rect 316144 2494 316464 9258
rect 316144 2258 316186 2494
rect 316422 2258 316464 2494
rect 316144 -746 316464 2258
rect 316144 -982 316186 -746
rect 316422 -982 316464 -746
rect 316144 -1066 316464 -982
rect 316144 -1302 316186 -1066
rect 316422 -1302 316464 -1066
rect 316144 -2294 316464 -1302
rect 317876 706198 318196 706230
rect 317876 705962 317918 706198
rect 318154 705962 318196 706198
rect 317876 705878 318196 705962
rect 317876 705642 317918 705878
rect 318154 705642 318196 705878
rect 317876 696561 318196 705642
rect 317876 696325 317918 696561
rect 318154 696325 318196 696561
rect 317876 689561 318196 696325
rect 317876 689325 317918 689561
rect 318154 689325 318196 689561
rect 317876 682561 318196 689325
rect 317876 682325 317918 682561
rect 318154 682325 318196 682561
rect 317876 675561 318196 682325
rect 317876 675325 317918 675561
rect 318154 675325 318196 675561
rect 317876 668561 318196 675325
rect 317876 668325 317918 668561
rect 318154 668325 318196 668561
rect 317876 661561 318196 668325
rect 317876 661325 317918 661561
rect 318154 661325 318196 661561
rect 317876 654561 318196 661325
rect 317876 654325 317918 654561
rect 318154 654325 318196 654561
rect 317876 647561 318196 654325
rect 317876 647325 317918 647561
rect 318154 647325 318196 647561
rect 317876 640561 318196 647325
rect 317876 640325 317918 640561
rect 318154 640325 318196 640561
rect 317876 633561 318196 640325
rect 317876 633325 317918 633561
rect 318154 633325 318196 633561
rect 317876 626561 318196 633325
rect 317876 626325 317918 626561
rect 318154 626325 318196 626561
rect 317876 619561 318196 626325
rect 317876 619325 317918 619561
rect 318154 619325 318196 619561
rect 317876 612561 318196 619325
rect 317876 612325 317918 612561
rect 318154 612325 318196 612561
rect 317876 605561 318196 612325
rect 317876 605325 317918 605561
rect 318154 605325 318196 605561
rect 317876 598561 318196 605325
rect 317876 598325 317918 598561
rect 318154 598325 318196 598561
rect 317876 591561 318196 598325
rect 317876 591325 317918 591561
rect 318154 591325 318196 591561
rect 317876 584561 318196 591325
rect 317876 584325 317918 584561
rect 318154 584325 318196 584561
rect 317876 577561 318196 584325
rect 317876 577325 317918 577561
rect 318154 577325 318196 577561
rect 317876 570561 318196 577325
rect 317876 570325 317918 570561
rect 318154 570325 318196 570561
rect 317876 563561 318196 570325
rect 317876 563325 317918 563561
rect 318154 563325 318196 563561
rect 317876 556561 318196 563325
rect 317876 556325 317918 556561
rect 318154 556325 318196 556561
rect 317876 549561 318196 556325
rect 317876 549325 317918 549561
rect 318154 549325 318196 549561
rect 317876 542561 318196 549325
rect 317876 542325 317918 542561
rect 318154 542325 318196 542561
rect 317876 535561 318196 542325
rect 317876 535325 317918 535561
rect 318154 535325 318196 535561
rect 317876 528561 318196 535325
rect 317876 528325 317918 528561
rect 318154 528325 318196 528561
rect 317876 521561 318196 528325
rect 317876 521325 317918 521561
rect 318154 521325 318196 521561
rect 317876 514561 318196 521325
rect 317876 514325 317918 514561
rect 318154 514325 318196 514561
rect 317876 507561 318196 514325
rect 317876 507325 317918 507561
rect 318154 507325 318196 507561
rect 317876 500561 318196 507325
rect 317876 500325 317918 500561
rect 318154 500325 318196 500561
rect 317876 493561 318196 500325
rect 317876 493325 317918 493561
rect 318154 493325 318196 493561
rect 317876 486561 318196 493325
rect 317876 486325 317918 486561
rect 318154 486325 318196 486561
rect 317876 479561 318196 486325
rect 317876 479325 317918 479561
rect 318154 479325 318196 479561
rect 317876 472561 318196 479325
rect 317876 472325 317918 472561
rect 318154 472325 318196 472561
rect 317876 465561 318196 472325
rect 317876 465325 317918 465561
rect 318154 465325 318196 465561
rect 317876 458561 318196 465325
rect 317876 458325 317918 458561
rect 318154 458325 318196 458561
rect 317876 451561 318196 458325
rect 317876 451325 317918 451561
rect 318154 451325 318196 451561
rect 317876 444561 318196 451325
rect 317876 444325 317918 444561
rect 318154 444325 318196 444561
rect 317876 437561 318196 444325
rect 317876 437325 317918 437561
rect 318154 437325 318196 437561
rect 317876 430561 318196 437325
rect 317876 430325 317918 430561
rect 318154 430325 318196 430561
rect 317876 423561 318196 430325
rect 317876 423325 317918 423561
rect 318154 423325 318196 423561
rect 317876 416561 318196 423325
rect 317876 416325 317918 416561
rect 318154 416325 318196 416561
rect 317876 409561 318196 416325
rect 317876 409325 317918 409561
rect 318154 409325 318196 409561
rect 317876 402561 318196 409325
rect 317876 402325 317918 402561
rect 318154 402325 318196 402561
rect 317876 395561 318196 402325
rect 317876 395325 317918 395561
rect 318154 395325 318196 395561
rect 317876 388561 318196 395325
rect 317876 388325 317918 388561
rect 318154 388325 318196 388561
rect 317876 381561 318196 388325
rect 317876 381325 317918 381561
rect 318154 381325 318196 381561
rect 317876 374561 318196 381325
rect 317876 374325 317918 374561
rect 318154 374325 318196 374561
rect 317876 367561 318196 374325
rect 317876 367325 317918 367561
rect 318154 367325 318196 367561
rect 317876 360561 318196 367325
rect 317876 360325 317918 360561
rect 318154 360325 318196 360561
rect 317876 353561 318196 360325
rect 317876 353325 317918 353561
rect 318154 353325 318196 353561
rect 317876 346561 318196 353325
rect 317876 346325 317918 346561
rect 318154 346325 318196 346561
rect 317876 339561 318196 346325
rect 317876 339325 317918 339561
rect 318154 339325 318196 339561
rect 317876 332561 318196 339325
rect 317876 332325 317918 332561
rect 318154 332325 318196 332561
rect 317876 325561 318196 332325
rect 317876 325325 317918 325561
rect 318154 325325 318196 325561
rect 317876 318561 318196 325325
rect 317876 318325 317918 318561
rect 318154 318325 318196 318561
rect 317876 311561 318196 318325
rect 317876 311325 317918 311561
rect 318154 311325 318196 311561
rect 317876 304561 318196 311325
rect 317876 304325 317918 304561
rect 318154 304325 318196 304561
rect 317876 297561 318196 304325
rect 317876 297325 317918 297561
rect 318154 297325 318196 297561
rect 317876 290561 318196 297325
rect 317876 290325 317918 290561
rect 318154 290325 318196 290561
rect 317876 283561 318196 290325
rect 317876 283325 317918 283561
rect 318154 283325 318196 283561
rect 317876 276561 318196 283325
rect 317876 276325 317918 276561
rect 318154 276325 318196 276561
rect 317876 269561 318196 276325
rect 317876 269325 317918 269561
rect 318154 269325 318196 269561
rect 317876 262561 318196 269325
rect 317876 262325 317918 262561
rect 318154 262325 318196 262561
rect 317876 255561 318196 262325
rect 317876 255325 317918 255561
rect 318154 255325 318196 255561
rect 317876 248561 318196 255325
rect 317876 248325 317918 248561
rect 318154 248325 318196 248561
rect 317876 241561 318196 248325
rect 317876 241325 317918 241561
rect 318154 241325 318196 241561
rect 317876 234561 318196 241325
rect 317876 234325 317918 234561
rect 318154 234325 318196 234561
rect 317876 227561 318196 234325
rect 317876 227325 317918 227561
rect 318154 227325 318196 227561
rect 317876 220561 318196 227325
rect 317876 220325 317918 220561
rect 318154 220325 318196 220561
rect 317876 213561 318196 220325
rect 317876 213325 317918 213561
rect 318154 213325 318196 213561
rect 317876 206561 318196 213325
rect 317876 206325 317918 206561
rect 318154 206325 318196 206561
rect 317876 199561 318196 206325
rect 317876 199325 317918 199561
rect 318154 199325 318196 199561
rect 317876 192561 318196 199325
rect 317876 192325 317918 192561
rect 318154 192325 318196 192561
rect 317876 185561 318196 192325
rect 317876 185325 317918 185561
rect 318154 185325 318196 185561
rect 317876 178561 318196 185325
rect 317876 178325 317918 178561
rect 318154 178325 318196 178561
rect 317876 171561 318196 178325
rect 317876 171325 317918 171561
rect 318154 171325 318196 171561
rect 317876 164561 318196 171325
rect 317876 164325 317918 164561
rect 318154 164325 318196 164561
rect 317876 157561 318196 164325
rect 317876 157325 317918 157561
rect 318154 157325 318196 157561
rect 317876 150561 318196 157325
rect 317876 150325 317918 150561
rect 318154 150325 318196 150561
rect 317876 143561 318196 150325
rect 317876 143325 317918 143561
rect 318154 143325 318196 143561
rect 317876 136561 318196 143325
rect 317876 136325 317918 136561
rect 318154 136325 318196 136561
rect 317876 129561 318196 136325
rect 317876 129325 317918 129561
rect 318154 129325 318196 129561
rect 317876 122561 318196 129325
rect 317876 122325 317918 122561
rect 318154 122325 318196 122561
rect 317876 115561 318196 122325
rect 317876 115325 317918 115561
rect 318154 115325 318196 115561
rect 317876 108561 318196 115325
rect 317876 108325 317918 108561
rect 318154 108325 318196 108561
rect 317876 101561 318196 108325
rect 317876 101325 317918 101561
rect 318154 101325 318196 101561
rect 317876 94561 318196 101325
rect 317876 94325 317918 94561
rect 318154 94325 318196 94561
rect 317876 87561 318196 94325
rect 317876 87325 317918 87561
rect 318154 87325 318196 87561
rect 317876 80561 318196 87325
rect 317876 80325 317918 80561
rect 318154 80325 318196 80561
rect 317876 73561 318196 80325
rect 317876 73325 317918 73561
rect 318154 73325 318196 73561
rect 317876 66561 318196 73325
rect 317876 66325 317918 66561
rect 318154 66325 318196 66561
rect 317876 59561 318196 66325
rect 317876 59325 317918 59561
rect 318154 59325 318196 59561
rect 317876 52561 318196 59325
rect 317876 52325 317918 52561
rect 318154 52325 318196 52561
rect 317876 45561 318196 52325
rect 317876 45325 317918 45561
rect 318154 45325 318196 45561
rect 317876 38561 318196 45325
rect 317876 38325 317918 38561
rect 318154 38325 318196 38561
rect 317876 31561 318196 38325
rect 317876 31325 317918 31561
rect 318154 31325 318196 31561
rect 317876 24561 318196 31325
rect 317876 24325 317918 24561
rect 318154 24325 318196 24561
rect 317876 17561 318196 24325
rect 317876 17325 317918 17561
rect 318154 17325 318196 17561
rect 317876 10561 318196 17325
rect 317876 10325 317918 10561
rect 318154 10325 318196 10561
rect 317876 3561 318196 10325
rect 317876 3325 317918 3561
rect 318154 3325 318196 3561
rect 317876 -1706 318196 3325
rect 317876 -1942 317918 -1706
rect 318154 -1942 318196 -1706
rect 317876 -2026 318196 -1942
rect 317876 -2262 317918 -2026
rect 318154 -2262 318196 -2026
rect 317876 -2294 318196 -2262
rect 323144 705238 323464 706230
rect 323144 705002 323186 705238
rect 323422 705002 323464 705238
rect 323144 704918 323464 705002
rect 323144 704682 323186 704918
rect 323422 704682 323464 704918
rect 323144 695494 323464 704682
rect 323144 695258 323186 695494
rect 323422 695258 323464 695494
rect 323144 688494 323464 695258
rect 323144 688258 323186 688494
rect 323422 688258 323464 688494
rect 323144 681494 323464 688258
rect 323144 681258 323186 681494
rect 323422 681258 323464 681494
rect 323144 674494 323464 681258
rect 323144 674258 323186 674494
rect 323422 674258 323464 674494
rect 323144 667494 323464 674258
rect 323144 667258 323186 667494
rect 323422 667258 323464 667494
rect 323144 660494 323464 667258
rect 323144 660258 323186 660494
rect 323422 660258 323464 660494
rect 323144 653494 323464 660258
rect 323144 653258 323186 653494
rect 323422 653258 323464 653494
rect 323144 646494 323464 653258
rect 323144 646258 323186 646494
rect 323422 646258 323464 646494
rect 323144 639494 323464 646258
rect 323144 639258 323186 639494
rect 323422 639258 323464 639494
rect 323144 632494 323464 639258
rect 323144 632258 323186 632494
rect 323422 632258 323464 632494
rect 323144 625494 323464 632258
rect 323144 625258 323186 625494
rect 323422 625258 323464 625494
rect 323144 618494 323464 625258
rect 323144 618258 323186 618494
rect 323422 618258 323464 618494
rect 323144 611494 323464 618258
rect 323144 611258 323186 611494
rect 323422 611258 323464 611494
rect 323144 604494 323464 611258
rect 323144 604258 323186 604494
rect 323422 604258 323464 604494
rect 323144 597494 323464 604258
rect 323144 597258 323186 597494
rect 323422 597258 323464 597494
rect 323144 590494 323464 597258
rect 323144 590258 323186 590494
rect 323422 590258 323464 590494
rect 323144 583494 323464 590258
rect 323144 583258 323186 583494
rect 323422 583258 323464 583494
rect 323144 576494 323464 583258
rect 323144 576258 323186 576494
rect 323422 576258 323464 576494
rect 323144 569494 323464 576258
rect 323144 569258 323186 569494
rect 323422 569258 323464 569494
rect 323144 562494 323464 569258
rect 323144 562258 323186 562494
rect 323422 562258 323464 562494
rect 323144 555494 323464 562258
rect 323144 555258 323186 555494
rect 323422 555258 323464 555494
rect 323144 548494 323464 555258
rect 323144 548258 323186 548494
rect 323422 548258 323464 548494
rect 323144 541494 323464 548258
rect 323144 541258 323186 541494
rect 323422 541258 323464 541494
rect 323144 534494 323464 541258
rect 323144 534258 323186 534494
rect 323422 534258 323464 534494
rect 323144 527494 323464 534258
rect 323144 527258 323186 527494
rect 323422 527258 323464 527494
rect 323144 520494 323464 527258
rect 323144 520258 323186 520494
rect 323422 520258 323464 520494
rect 323144 513494 323464 520258
rect 323144 513258 323186 513494
rect 323422 513258 323464 513494
rect 323144 506494 323464 513258
rect 323144 506258 323186 506494
rect 323422 506258 323464 506494
rect 323144 499494 323464 506258
rect 323144 499258 323186 499494
rect 323422 499258 323464 499494
rect 323144 492494 323464 499258
rect 323144 492258 323186 492494
rect 323422 492258 323464 492494
rect 323144 485494 323464 492258
rect 323144 485258 323186 485494
rect 323422 485258 323464 485494
rect 323144 478494 323464 485258
rect 323144 478258 323186 478494
rect 323422 478258 323464 478494
rect 323144 471494 323464 478258
rect 323144 471258 323186 471494
rect 323422 471258 323464 471494
rect 323144 464494 323464 471258
rect 323144 464258 323186 464494
rect 323422 464258 323464 464494
rect 323144 457494 323464 464258
rect 323144 457258 323186 457494
rect 323422 457258 323464 457494
rect 323144 450494 323464 457258
rect 323144 450258 323186 450494
rect 323422 450258 323464 450494
rect 323144 443494 323464 450258
rect 323144 443258 323186 443494
rect 323422 443258 323464 443494
rect 323144 436494 323464 443258
rect 323144 436258 323186 436494
rect 323422 436258 323464 436494
rect 323144 429494 323464 436258
rect 323144 429258 323186 429494
rect 323422 429258 323464 429494
rect 323144 422494 323464 429258
rect 323144 422258 323186 422494
rect 323422 422258 323464 422494
rect 323144 415494 323464 422258
rect 323144 415258 323186 415494
rect 323422 415258 323464 415494
rect 323144 408494 323464 415258
rect 323144 408258 323186 408494
rect 323422 408258 323464 408494
rect 323144 401494 323464 408258
rect 323144 401258 323186 401494
rect 323422 401258 323464 401494
rect 323144 394494 323464 401258
rect 323144 394258 323186 394494
rect 323422 394258 323464 394494
rect 323144 387494 323464 394258
rect 323144 387258 323186 387494
rect 323422 387258 323464 387494
rect 323144 380494 323464 387258
rect 323144 380258 323186 380494
rect 323422 380258 323464 380494
rect 323144 373494 323464 380258
rect 323144 373258 323186 373494
rect 323422 373258 323464 373494
rect 323144 366494 323464 373258
rect 323144 366258 323186 366494
rect 323422 366258 323464 366494
rect 323144 359494 323464 366258
rect 323144 359258 323186 359494
rect 323422 359258 323464 359494
rect 323144 352494 323464 359258
rect 323144 352258 323186 352494
rect 323422 352258 323464 352494
rect 323144 345494 323464 352258
rect 323144 345258 323186 345494
rect 323422 345258 323464 345494
rect 323144 338494 323464 345258
rect 323144 338258 323186 338494
rect 323422 338258 323464 338494
rect 323144 331494 323464 338258
rect 323144 331258 323186 331494
rect 323422 331258 323464 331494
rect 323144 324494 323464 331258
rect 323144 324258 323186 324494
rect 323422 324258 323464 324494
rect 323144 317494 323464 324258
rect 323144 317258 323186 317494
rect 323422 317258 323464 317494
rect 323144 310494 323464 317258
rect 323144 310258 323186 310494
rect 323422 310258 323464 310494
rect 323144 303494 323464 310258
rect 323144 303258 323186 303494
rect 323422 303258 323464 303494
rect 323144 296494 323464 303258
rect 323144 296258 323186 296494
rect 323422 296258 323464 296494
rect 323144 289494 323464 296258
rect 323144 289258 323186 289494
rect 323422 289258 323464 289494
rect 323144 282494 323464 289258
rect 323144 282258 323186 282494
rect 323422 282258 323464 282494
rect 323144 275494 323464 282258
rect 323144 275258 323186 275494
rect 323422 275258 323464 275494
rect 323144 268494 323464 275258
rect 323144 268258 323186 268494
rect 323422 268258 323464 268494
rect 323144 261494 323464 268258
rect 323144 261258 323186 261494
rect 323422 261258 323464 261494
rect 323144 254494 323464 261258
rect 323144 254258 323186 254494
rect 323422 254258 323464 254494
rect 323144 247494 323464 254258
rect 323144 247258 323186 247494
rect 323422 247258 323464 247494
rect 323144 240494 323464 247258
rect 323144 240258 323186 240494
rect 323422 240258 323464 240494
rect 323144 233494 323464 240258
rect 323144 233258 323186 233494
rect 323422 233258 323464 233494
rect 323144 226494 323464 233258
rect 323144 226258 323186 226494
rect 323422 226258 323464 226494
rect 323144 219494 323464 226258
rect 323144 219258 323186 219494
rect 323422 219258 323464 219494
rect 323144 212494 323464 219258
rect 323144 212258 323186 212494
rect 323422 212258 323464 212494
rect 323144 205494 323464 212258
rect 323144 205258 323186 205494
rect 323422 205258 323464 205494
rect 323144 198494 323464 205258
rect 323144 198258 323186 198494
rect 323422 198258 323464 198494
rect 323144 191494 323464 198258
rect 323144 191258 323186 191494
rect 323422 191258 323464 191494
rect 323144 184494 323464 191258
rect 323144 184258 323186 184494
rect 323422 184258 323464 184494
rect 323144 177494 323464 184258
rect 323144 177258 323186 177494
rect 323422 177258 323464 177494
rect 323144 170494 323464 177258
rect 323144 170258 323186 170494
rect 323422 170258 323464 170494
rect 323144 163494 323464 170258
rect 323144 163258 323186 163494
rect 323422 163258 323464 163494
rect 323144 156494 323464 163258
rect 323144 156258 323186 156494
rect 323422 156258 323464 156494
rect 323144 149494 323464 156258
rect 323144 149258 323186 149494
rect 323422 149258 323464 149494
rect 323144 142494 323464 149258
rect 323144 142258 323186 142494
rect 323422 142258 323464 142494
rect 323144 135494 323464 142258
rect 323144 135258 323186 135494
rect 323422 135258 323464 135494
rect 323144 128494 323464 135258
rect 323144 128258 323186 128494
rect 323422 128258 323464 128494
rect 323144 121494 323464 128258
rect 323144 121258 323186 121494
rect 323422 121258 323464 121494
rect 323144 114494 323464 121258
rect 323144 114258 323186 114494
rect 323422 114258 323464 114494
rect 323144 107494 323464 114258
rect 323144 107258 323186 107494
rect 323422 107258 323464 107494
rect 323144 100494 323464 107258
rect 323144 100258 323186 100494
rect 323422 100258 323464 100494
rect 323144 93494 323464 100258
rect 323144 93258 323186 93494
rect 323422 93258 323464 93494
rect 323144 86494 323464 93258
rect 323144 86258 323186 86494
rect 323422 86258 323464 86494
rect 323144 79494 323464 86258
rect 323144 79258 323186 79494
rect 323422 79258 323464 79494
rect 323144 72494 323464 79258
rect 323144 72258 323186 72494
rect 323422 72258 323464 72494
rect 323144 65494 323464 72258
rect 323144 65258 323186 65494
rect 323422 65258 323464 65494
rect 323144 58494 323464 65258
rect 323144 58258 323186 58494
rect 323422 58258 323464 58494
rect 323144 51494 323464 58258
rect 323144 51258 323186 51494
rect 323422 51258 323464 51494
rect 323144 44494 323464 51258
rect 323144 44258 323186 44494
rect 323422 44258 323464 44494
rect 323144 37494 323464 44258
rect 323144 37258 323186 37494
rect 323422 37258 323464 37494
rect 323144 30494 323464 37258
rect 323144 30258 323186 30494
rect 323422 30258 323464 30494
rect 323144 23494 323464 30258
rect 323144 23258 323186 23494
rect 323422 23258 323464 23494
rect 323144 16494 323464 23258
rect 323144 16258 323186 16494
rect 323422 16258 323464 16494
rect 323144 9494 323464 16258
rect 323144 9258 323186 9494
rect 323422 9258 323464 9494
rect 323144 2494 323464 9258
rect 323144 2258 323186 2494
rect 323422 2258 323464 2494
rect 323144 -746 323464 2258
rect 323144 -982 323186 -746
rect 323422 -982 323464 -746
rect 323144 -1066 323464 -982
rect 323144 -1302 323186 -1066
rect 323422 -1302 323464 -1066
rect 323144 -2294 323464 -1302
rect 324876 706198 325196 706230
rect 324876 705962 324918 706198
rect 325154 705962 325196 706198
rect 324876 705878 325196 705962
rect 324876 705642 324918 705878
rect 325154 705642 325196 705878
rect 324876 696561 325196 705642
rect 324876 696325 324918 696561
rect 325154 696325 325196 696561
rect 324876 689561 325196 696325
rect 324876 689325 324918 689561
rect 325154 689325 325196 689561
rect 324876 682561 325196 689325
rect 324876 682325 324918 682561
rect 325154 682325 325196 682561
rect 324876 675561 325196 682325
rect 324876 675325 324918 675561
rect 325154 675325 325196 675561
rect 324876 668561 325196 675325
rect 324876 668325 324918 668561
rect 325154 668325 325196 668561
rect 324876 661561 325196 668325
rect 324876 661325 324918 661561
rect 325154 661325 325196 661561
rect 324876 654561 325196 661325
rect 324876 654325 324918 654561
rect 325154 654325 325196 654561
rect 324876 647561 325196 654325
rect 324876 647325 324918 647561
rect 325154 647325 325196 647561
rect 324876 640561 325196 647325
rect 324876 640325 324918 640561
rect 325154 640325 325196 640561
rect 324876 633561 325196 640325
rect 324876 633325 324918 633561
rect 325154 633325 325196 633561
rect 324876 626561 325196 633325
rect 324876 626325 324918 626561
rect 325154 626325 325196 626561
rect 324876 619561 325196 626325
rect 324876 619325 324918 619561
rect 325154 619325 325196 619561
rect 324876 612561 325196 619325
rect 324876 612325 324918 612561
rect 325154 612325 325196 612561
rect 324876 605561 325196 612325
rect 324876 605325 324918 605561
rect 325154 605325 325196 605561
rect 324876 598561 325196 605325
rect 324876 598325 324918 598561
rect 325154 598325 325196 598561
rect 324876 591561 325196 598325
rect 324876 591325 324918 591561
rect 325154 591325 325196 591561
rect 324876 584561 325196 591325
rect 324876 584325 324918 584561
rect 325154 584325 325196 584561
rect 324876 577561 325196 584325
rect 324876 577325 324918 577561
rect 325154 577325 325196 577561
rect 324876 570561 325196 577325
rect 324876 570325 324918 570561
rect 325154 570325 325196 570561
rect 324876 563561 325196 570325
rect 324876 563325 324918 563561
rect 325154 563325 325196 563561
rect 324876 556561 325196 563325
rect 324876 556325 324918 556561
rect 325154 556325 325196 556561
rect 324876 549561 325196 556325
rect 324876 549325 324918 549561
rect 325154 549325 325196 549561
rect 324876 542561 325196 549325
rect 324876 542325 324918 542561
rect 325154 542325 325196 542561
rect 324876 535561 325196 542325
rect 324876 535325 324918 535561
rect 325154 535325 325196 535561
rect 324876 528561 325196 535325
rect 324876 528325 324918 528561
rect 325154 528325 325196 528561
rect 324876 521561 325196 528325
rect 324876 521325 324918 521561
rect 325154 521325 325196 521561
rect 324876 514561 325196 521325
rect 324876 514325 324918 514561
rect 325154 514325 325196 514561
rect 324876 507561 325196 514325
rect 324876 507325 324918 507561
rect 325154 507325 325196 507561
rect 324876 500561 325196 507325
rect 324876 500325 324918 500561
rect 325154 500325 325196 500561
rect 324876 493561 325196 500325
rect 324876 493325 324918 493561
rect 325154 493325 325196 493561
rect 324876 486561 325196 493325
rect 324876 486325 324918 486561
rect 325154 486325 325196 486561
rect 324876 479561 325196 486325
rect 324876 479325 324918 479561
rect 325154 479325 325196 479561
rect 324876 472561 325196 479325
rect 324876 472325 324918 472561
rect 325154 472325 325196 472561
rect 324876 465561 325196 472325
rect 324876 465325 324918 465561
rect 325154 465325 325196 465561
rect 324876 458561 325196 465325
rect 324876 458325 324918 458561
rect 325154 458325 325196 458561
rect 324876 451561 325196 458325
rect 324876 451325 324918 451561
rect 325154 451325 325196 451561
rect 324876 444561 325196 451325
rect 324876 444325 324918 444561
rect 325154 444325 325196 444561
rect 324876 437561 325196 444325
rect 324876 437325 324918 437561
rect 325154 437325 325196 437561
rect 324876 430561 325196 437325
rect 324876 430325 324918 430561
rect 325154 430325 325196 430561
rect 324876 423561 325196 430325
rect 324876 423325 324918 423561
rect 325154 423325 325196 423561
rect 324876 416561 325196 423325
rect 324876 416325 324918 416561
rect 325154 416325 325196 416561
rect 324876 409561 325196 416325
rect 324876 409325 324918 409561
rect 325154 409325 325196 409561
rect 324876 402561 325196 409325
rect 324876 402325 324918 402561
rect 325154 402325 325196 402561
rect 324876 395561 325196 402325
rect 324876 395325 324918 395561
rect 325154 395325 325196 395561
rect 324876 388561 325196 395325
rect 324876 388325 324918 388561
rect 325154 388325 325196 388561
rect 324876 381561 325196 388325
rect 324876 381325 324918 381561
rect 325154 381325 325196 381561
rect 324876 374561 325196 381325
rect 324876 374325 324918 374561
rect 325154 374325 325196 374561
rect 324876 367561 325196 374325
rect 324876 367325 324918 367561
rect 325154 367325 325196 367561
rect 324876 360561 325196 367325
rect 324876 360325 324918 360561
rect 325154 360325 325196 360561
rect 324876 353561 325196 360325
rect 324876 353325 324918 353561
rect 325154 353325 325196 353561
rect 324876 346561 325196 353325
rect 324876 346325 324918 346561
rect 325154 346325 325196 346561
rect 324876 339561 325196 346325
rect 324876 339325 324918 339561
rect 325154 339325 325196 339561
rect 324876 332561 325196 339325
rect 324876 332325 324918 332561
rect 325154 332325 325196 332561
rect 324876 325561 325196 332325
rect 324876 325325 324918 325561
rect 325154 325325 325196 325561
rect 324876 318561 325196 325325
rect 324876 318325 324918 318561
rect 325154 318325 325196 318561
rect 324876 311561 325196 318325
rect 324876 311325 324918 311561
rect 325154 311325 325196 311561
rect 324876 304561 325196 311325
rect 324876 304325 324918 304561
rect 325154 304325 325196 304561
rect 324876 297561 325196 304325
rect 324876 297325 324918 297561
rect 325154 297325 325196 297561
rect 324876 290561 325196 297325
rect 324876 290325 324918 290561
rect 325154 290325 325196 290561
rect 324876 283561 325196 290325
rect 324876 283325 324918 283561
rect 325154 283325 325196 283561
rect 324876 276561 325196 283325
rect 324876 276325 324918 276561
rect 325154 276325 325196 276561
rect 324876 269561 325196 276325
rect 324876 269325 324918 269561
rect 325154 269325 325196 269561
rect 324876 262561 325196 269325
rect 324876 262325 324918 262561
rect 325154 262325 325196 262561
rect 324876 255561 325196 262325
rect 324876 255325 324918 255561
rect 325154 255325 325196 255561
rect 324876 248561 325196 255325
rect 324876 248325 324918 248561
rect 325154 248325 325196 248561
rect 324876 241561 325196 248325
rect 324876 241325 324918 241561
rect 325154 241325 325196 241561
rect 324876 234561 325196 241325
rect 324876 234325 324918 234561
rect 325154 234325 325196 234561
rect 324876 227561 325196 234325
rect 324876 227325 324918 227561
rect 325154 227325 325196 227561
rect 324876 220561 325196 227325
rect 324876 220325 324918 220561
rect 325154 220325 325196 220561
rect 324876 213561 325196 220325
rect 324876 213325 324918 213561
rect 325154 213325 325196 213561
rect 324876 206561 325196 213325
rect 324876 206325 324918 206561
rect 325154 206325 325196 206561
rect 324876 199561 325196 206325
rect 324876 199325 324918 199561
rect 325154 199325 325196 199561
rect 324876 192561 325196 199325
rect 324876 192325 324918 192561
rect 325154 192325 325196 192561
rect 324876 185561 325196 192325
rect 324876 185325 324918 185561
rect 325154 185325 325196 185561
rect 324876 178561 325196 185325
rect 324876 178325 324918 178561
rect 325154 178325 325196 178561
rect 324876 171561 325196 178325
rect 324876 171325 324918 171561
rect 325154 171325 325196 171561
rect 324876 164561 325196 171325
rect 324876 164325 324918 164561
rect 325154 164325 325196 164561
rect 324876 157561 325196 164325
rect 324876 157325 324918 157561
rect 325154 157325 325196 157561
rect 324876 150561 325196 157325
rect 324876 150325 324918 150561
rect 325154 150325 325196 150561
rect 324876 143561 325196 150325
rect 324876 143325 324918 143561
rect 325154 143325 325196 143561
rect 324876 136561 325196 143325
rect 324876 136325 324918 136561
rect 325154 136325 325196 136561
rect 324876 129561 325196 136325
rect 324876 129325 324918 129561
rect 325154 129325 325196 129561
rect 324876 122561 325196 129325
rect 324876 122325 324918 122561
rect 325154 122325 325196 122561
rect 324876 115561 325196 122325
rect 324876 115325 324918 115561
rect 325154 115325 325196 115561
rect 324876 108561 325196 115325
rect 324876 108325 324918 108561
rect 325154 108325 325196 108561
rect 324876 101561 325196 108325
rect 324876 101325 324918 101561
rect 325154 101325 325196 101561
rect 324876 94561 325196 101325
rect 324876 94325 324918 94561
rect 325154 94325 325196 94561
rect 324876 87561 325196 94325
rect 324876 87325 324918 87561
rect 325154 87325 325196 87561
rect 324876 80561 325196 87325
rect 324876 80325 324918 80561
rect 325154 80325 325196 80561
rect 324876 73561 325196 80325
rect 324876 73325 324918 73561
rect 325154 73325 325196 73561
rect 324876 66561 325196 73325
rect 324876 66325 324918 66561
rect 325154 66325 325196 66561
rect 324876 59561 325196 66325
rect 324876 59325 324918 59561
rect 325154 59325 325196 59561
rect 324876 52561 325196 59325
rect 324876 52325 324918 52561
rect 325154 52325 325196 52561
rect 324876 45561 325196 52325
rect 324876 45325 324918 45561
rect 325154 45325 325196 45561
rect 324876 38561 325196 45325
rect 324876 38325 324918 38561
rect 325154 38325 325196 38561
rect 324876 31561 325196 38325
rect 324876 31325 324918 31561
rect 325154 31325 325196 31561
rect 324876 24561 325196 31325
rect 324876 24325 324918 24561
rect 325154 24325 325196 24561
rect 324876 17561 325196 24325
rect 324876 17325 324918 17561
rect 325154 17325 325196 17561
rect 324876 10561 325196 17325
rect 324876 10325 324918 10561
rect 325154 10325 325196 10561
rect 324876 3561 325196 10325
rect 324876 3325 324918 3561
rect 325154 3325 325196 3561
rect 324876 -1706 325196 3325
rect 324876 -1942 324918 -1706
rect 325154 -1942 325196 -1706
rect 324876 -2026 325196 -1942
rect 324876 -2262 324918 -2026
rect 325154 -2262 325196 -2026
rect 324876 -2294 325196 -2262
rect 330144 705238 330464 706230
rect 330144 705002 330186 705238
rect 330422 705002 330464 705238
rect 330144 704918 330464 705002
rect 330144 704682 330186 704918
rect 330422 704682 330464 704918
rect 330144 695494 330464 704682
rect 330144 695258 330186 695494
rect 330422 695258 330464 695494
rect 330144 688494 330464 695258
rect 330144 688258 330186 688494
rect 330422 688258 330464 688494
rect 330144 681494 330464 688258
rect 330144 681258 330186 681494
rect 330422 681258 330464 681494
rect 330144 674494 330464 681258
rect 330144 674258 330186 674494
rect 330422 674258 330464 674494
rect 330144 667494 330464 674258
rect 330144 667258 330186 667494
rect 330422 667258 330464 667494
rect 330144 660494 330464 667258
rect 330144 660258 330186 660494
rect 330422 660258 330464 660494
rect 330144 653494 330464 660258
rect 330144 653258 330186 653494
rect 330422 653258 330464 653494
rect 330144 646494 330464 653258
rect 330144 646258 330186 646494
rect 330422 646258 330464 646494
rect 330144 639494 330464 646258
rect 330144 639258 330186 639494
rect 330422 639258 330464 639494
rect 330144 632494 330464 639258
rect 330144 632258 330186 632494
rect 330422 632258 330464 632494
rect 330144 625494 330464 632258
rect 330144 625258 330186 625494
rect 330422 625258 330464 625494
rect 330144 618494 330464 625258
rect 330144 618258 330186 618494
rect 330422 618258 330464 618494
rect 330144 611494 330464 618258
rect 330144 611258 330186 611494
rect 330422 611258 330464 611494
rect 330144 604494 330464 611258
rect 330144 604258 330186 604494
rect 330422 604258 330464 604494
rect 330144 597494 330464 604258
rect 330144 597258 330186 597494
rect 330422 597258 330464 597494
rect 330144 590494 330464 597258
rect 330144 590258 330186 590494
rect 330422 590258 330464 590494
rect 330144 583494 330464 590258
rect 330144 583258 330186 583494
rect 330422 583258 330464 583494
rect 330144 576494 330464 583258
rect 330144 576258 330186 576494
rect 330422 576258 330464 576494
rect 330144 569494 330464 576258
rect 330144 569258 330186 569494
rect 330422 569258 330464 569494
rect 330144 562494 330464 569258
rect 330144 562258 330186 562494
rect 330422 562258 330464 562494
rect 330144 555494 330464 562258
rect 330144 555258 330186 555494
rect 330422 555258 330464 555494
rect 330144 548494 330464 555258
rect 330144 548258 330186 548494
rect 330422 548258 330464 548494
rect 330144 541494 330464 548258
rect 330144 541258 330186 541494
rect 330422 541258 330464 541494
rect 330144 534494 330464 541258
rect 330144 534258 330186 534494
rect 330422 534258 330464 534494
rect 330144 527494 330464 534258
rect 330144 527258 330186 527494
rect 330422 527258 330464 527494
rect 330144 520494 330464 527258
rect 330144 520258 330186 520494
rect 330422 520258 330464 520494
rect 330144 513494 330464 520258
rect 330144 513258 330186 513494
rect 330422 513258 330464 513494
rect 330144 506494 330464 513258
rect 330144 506258 330186 506494
rect 330422 506258 330464 506494
rect 330144 499494 330464 506258
rect 330144 499258 330186 499494
rect 330422 499258 330464 499494
rect 330144 492494 330464 499258
rect 330144 492258 330186 492494
rect 330422 492258 330464 492494
rect 330144 485494 330464 492258
rect 330144 485258 330186 485494
rect 330422 485258 330464 485494
rect 330144 478494 330464 485258
rect 330144 478258 330186 478494
rect 330422 478258 330464 478494
rect 330144 471494 330464 478258
rect 330144 471258 330186 471494
rect 330422 471258 330464 471494
rect 330144 464494 330464 471258
rect 330144 464258 330186 464494
rect 330422 464258 330464 464494
rect 330144 457494 330464 464258
rect 330144 457258 330186 457494
rect 330422 457258 330464 457494
rect 330144 450494 330464 457258
rect 330144 450258 330186 450494
rect 330422 450258 330464 450494
rect 330144 443494 330464 450258
rect 330144 443258 330186 443494
rect 330422 443258 330464 443494
rect 330144 436494 330464 443258
rect 330144 436258 330186 436494
rect 330422 436258 330464 436494
rect 330144 429494 330464 436258
rect 330144 429258 330186 429494
rect 330422 429258 330464 429494
rect 330144 422494 330464 429258
rect 330144 422258 330186 422494
rect 330422 422258 330464 422494
rect 330144 415494 330464 422258
rect 330144 415258 330186 415494
rect 330422 415258 330464 415494
rect 330144 408494 330464 415258
rect 330144 408258 330186 408494
rect 330422 408258 330464 408494
rect 330144 401494 330464 408258
rect 330144 401258 330186 401494
rect 330422 401258 330464 401494
rect 330144 394494 330464 401258
rect 330144 394258 330186 394494
rect 330422 394258 330464 394494
rect 330144 387494 330464 394258
rect 330144 387258 330186 387494
rect 330422 387258 330464 387494
rect 330144 380494 330464 387258
rect 330144 380258 330186 380494
rect 330422 380258 330464 380494
rect 330144 373494 330464 380258
rect 330144 373258 330186 373494
rect 330422 373258 330464 373494
rect 330144 366494 330464 373258
rect 330144 366258 330186 366494
rect 330422 366258 330464 366494
rect 330144 359494 330464 366258
rect 330144 359258 330186 359494
rect 330422 359258 330464 359494
rect 330144 352494 330464 359258
rect 330144 352258 330186 352494
rect 330422 352258 330464 352494
rect 330144 345494 330464 352258
rect 330144 345258 330186 345494
rect 330422 345258 330464 345494
rect 330144 338494 330464 345258
rect 330144 338258 330186 338494
rect 330422 338258 330464 338494
rect 330144 331494 330464 338258
rect 330144 331258 330186 331494
rect 330422 331258 330464 331494
rect 330144 324494 330464 331258
rect 330144 324258 330186 324494
rect 330422 324258 330464 324494
rect 330144 317494 330464 324258
rect 330144 317258 330186 317494
rect 330422 317258 330464 317494
rect 330144 310494 330464 317258
rect 330144 310258 330186 310494
rect 330422 310258 330464 310494
rect 330144 303494 330464 310258
rect 330144 303258 330186 303494
rect 330422 303258 330464 303494
rect 330144 296494 330464 303258
rect 330144 296258 330186 296494
rect 330422 296258 330464 296494
rect 330144 289494 330464 296258
rect 330144 289258 330186 289494
rect 330422 289258 330464 289494
rect 330144 282494 330464 289258
rect 330144 282258 330186 282494
rect 330422 282258 330464 282494
rect 330144 275494 330464 282258
rect 330144 275258 330186 275494
rect 330422 275258 330464 275494
rect 330144 268494 330464 275258
rect 330144 268258 330186 268494
rect 330422 268258 330464 268494
rect 330144 261494 330464 268258
rect 330144 261258 330186 261494
rect 330422 261258 330464 261494
rect 330144 254494 330464 261258
rect 330144 254258 330186 254494
rect 330422 254258 330464 254494
rect 330144 247494 330464 254258
rect 330144 247258 330186 247494
rect 330422 247258 330464 247494
rect 330144 240494 330464 247258
rect 330144 240258 330186 240494
rect 330422 240258 330464 240494
rect 330144 233494 330464 240258
rect 330144 233258 330186 233494
rect 330422 233258 330464 233494
rect 330144 226494 330464 233258
rect 330144 226258 330186 226494
rect 330422 226258 330464 226494
rect 330144 219494 330464 226258
rect 330144 219258 330186 219494
rect 330422 219258 330464 219494
rect 330144 212494 330464 219258
rect 330144 212258 330186 212494
rect 330422 212258 330464 212494
rect 330144 205494 330464 212258
rect 330144 205258 330186 205494
rect 330422 205258 330464 205494
rect 330144 198494 330464 205258
rect 330144 198258 330186 198494
rect 330422 198258 330464 198494
rect 330144 191494 330464 198258
rect 330144 191258 330186 191494
rect 330422 191258 330464 191494
rect 330144 184494 330464 191258
rect 330144 184258 330186 184494
rect 330422 184258 330464 184494
rect 330144 177494 330464 184258
rect 330144 177258 330186 177494
rect 330422 177258 330464 177494
rect 330144 170494 330464 177258
rect 330144 170258 330186 170494
rect 330422 170258 330464 170494
rect 330144 163494 330464 170258
rect 330144 163258 330186 163494
rect 330422 163258 330464 163494
rect 330144 156494 330464 163258
rect 330144 156258 330186 156494
rect 330422 156258 330464 156494
rect 330144 149494 330464 156258
rect 330144 149258 330186 149494
rect 330422 149258 330464 149494
rect 330144 142494 330464 149258
rect 330144 142258 330186 142494
rect 330422 142258 330464 142494
rect 330144 135494 330464 142258
rect 330144 135258 330186 135494
rect 330422 135258 330464 135494
rect 330144 128494 330464 135258
rect 330144 128258 330186 128494
rect 330422 128258 330464 128494
rect 330144 121494 330464 128258
rect 330144 121258 330186 121494
rect 330422 121258 330464 121494
rect 330144 114494 330464 121258
rect 330144 114258 330186 114494
rect 330422 114258 330464 114494
rect 330144 107494 330464 114258
rect 330144 107258 330186 107494
rect 330422 107258 330464 107494
rect 330144 100494 330464 107258
rect 330144 100258 330186 100494
rect 330422 100258 330464 100494
rect 330144 93494 330464 100258
rect 330144 93258 330186 93494
rect 330422 93258 330464 93494
rect 330144 86494 330464 93258
rect 330144 86258 330186 86494
rect 330422 86258 330464 86494
rect 330144 79494 330464 86258
rect 330144 79258 330186 79494
rect 330422 79258 330464 79494
rect 330144 72494 330464 79258
rect 330144 72258 330186 72494
rect 330422 72258 330464 72494
rect 330144 65494 330464 72258
rect 330144 65258 330186 65494
rect 330422 65258 330464 65494
rect 330144 58494 330464 65258
rect 330144 58258 330186 58494
rect 330422 58258 330464 58494
rect 330144 51494 330464 58258
rect 330144 51258 330186 51494
rect 330422 51258 330464 51494
rect 330144 44494 330464 51258
rect 330144 44258 330186 44494
rect 330422 44258 330464 44494
rect 330144 37494 330464 44258
rect 330144 37258 330186 37494
rect 330422 37258 330464 37494
rect 330144 30494 330464 37258
rect 330144 30258 330186 30494
rect 330422 30258 330464 30494
rect 330144 23494 330464 30258
rect 330144 23258 330186 23494
rect 330422 23258 330464 23494
rect 330144 16494 330464 23258
rect 330144 16258 330186 16494
rect 330422 16258 330464 16494
rect 330144 9494 330464 16258
rect 330144 9258 330186 9494
rect 330422 9258 330464 9494
rect 330144 2494 330464 9258
rect 330144 2258 330186 2494
rect 330422 2258 330464 2494
rect 330144 -746 330464 2258
rect 330144 -982 330186 -746
rect 330422 -982 330464 -746
rect 330144 -1066 330464 -982
rect 330144 -1302 330186 -1066
rect 330422 -1302 330464 -1066
rect 330144 -2294 330464 -1302
rect 331876 706198 332196 706230
rect 331876 705962 331918 706198
rect 332154 705962 332196 706198
rect 331876 705878 332196 705962
rect 331876 705642 331918 705878
rect 332154 705642 332196 705878
rect 331876 696561 332196 705642
rect 331876 696325 331918 696561
rect 332154 696325 332196 696561
rect 331876 689561 332196 696325
rect 331876 689325 331918 689561
rect 332154 689325 332196 689561
rect 331876 682561 332196 689325
rect 331876 682325 331918 682561
rect 332154 682325 332196 682561
rect 331876 675561 332196 682325
rect 331876 675325 331918 675561
rect 332154 675325 332196 675561
rect 331876 668561 332196 675325
rect 331876 668325 331918 668561
rect 332154 668325 332196 668561
rect 331876 661561 332196 668325
rect 331876 661325 331918 661561
rect 332154 661325 332196 661561
rect 331876 654561 332196 661325
rect 331876 654325 331918 654561
rect 332154 654325 332196 654561
rect 331876 647561 332196 654325
rect 331876 647325 331918 647561
rect 332154 647325 332196 647561
rect 331876 640561 332196 647325
rect 331876 640325 331918 640561
rect 332154 640325 332196 640561
rect 331876 633561 332196 640325
rect 331876 633325 331918 633561
rect 332154 633325 332196 633561
rect 331876 626561 332196 633325
rect 331876 626325 331918 626561
rect 332154 626325 332196 626561
rect 331876 619561 332196 626325
rect 331876 619325 331918 619561
rect 332154 619325 332196 619561
rect 331876 612561 332196 619325
rect 331876 612325 331918 612561
rect 332154 612325 332196 612561
rect 331876 605561 332196 612325
rect 331876 605325 331918 605561
rect 332154 605325 332196 605561
rect 331876 598561 332196 605325
rect 331876 598325 331918 598561
rect 332154 598325 332196 598561
rect 331876 591561 332196 598325
rect 331876 591325 331918 591561
rect 332154 591325 332196 591561
rect 331876 584561 332196 591325
rect 331876 584325 331918 584561
rect 332154 584325 332196 584561
rect 331876 577561 332196 584325
rect 331876 577325 331918 577561
rect 332154 577325 332196 577561
rect 331876 570561 332196 577325
rect 331876 570325 331918 570561
rect 332154 570325 332196 570561
rect 331876 563561 332196 570325
rect 331876 563325 331918 563561
rect 332154 563325 332196 563561
rect 331876 556561 332196 563325
rect 331876 556325 331918 556561
rect 332154 556325 332196 556561
rect 331876 549561 332196 556325
rect 331876 549325 331918 549561
rect 332154 549325 332196 549561
rect 331876 542561 332196 549325
rect 331876 542325 331918 542561
rect 332154 542325 332196 542561
rect 331876 535561 332196 542325
rect 331876 535325 331918 535561
rect 332154 535325 332196 535561
rect 331876 528561 332196 535325
rect 331876 528325 331918 528561
rect 332154 528325 332196 528561
rect 331876 521561 332196 528325
rect 331876 521325 331918 521561
rect 332154 521325 332196 521561
rect 331876 514561 332196 521325
rect 331876 514325 331918 514561
rect 332154 514325 332196 514561
rect 331876 507561 332196 514325
rect 331876 507325 331918 507561
rect 332154 507325 332196 507561
rect 331876 500561 332196 507325
rect 331876 500325 331918 500561
rect 332154 500325 332196 500561
rect 331876 493561 332196 500325
rect 331876 493325 331918 493561
rect 332154 493325 332196 493561
rect 331876 486561 332196 493325
rect 331876 486325 331918 486561
rect 332154 486325 332196 486561
rect 331876 479561 332196 486325
rect 331876 479325 331918 479561
rect 332154 479325 332196 479561
rect 331876 472561 332196 479325
rect 331876 472325 331918 472561
rect 332154 472325 332196 472561
rect 331876 465561 332196 472325
rect 331876 465325 331918 465561
rect 332154 465325 332196 465561
rect 331876 458561 332196 465325
rect 331876 458325 331918 458561
rect 332154 458325 332196 458561
rect 331876 451561 332196 458325
rect 331876 451325 331918 451561
rect 332154 451325 332196 451561
rect 331876 444561 332196 451325
rect 331876 444325 331918 444561
rect 332154 444325 332196 444561
rect 331876 437561 332196 444325
rect 331876 437325 331918 437561
rect 332154 437325 332196 437561
rect 331876 430561 332196 437325
rect 331876 430325 331918 430561
rect 332154 430325 332196 430561
rect 331876 423561 332196 430325
rect 331876 423325 331918 423561
rect 332154 423325 332196 423561
rect 331876 416561 332196 423325
rect 331876 416325 331918 416561
rect 332154 416325 332196 416561
rect 331876 409561 332196 416325
rect 331876 409325 331918 409561
rect 332154 409325 332196 409561
rect 331876 402561 332196 409325
rect 331876 402325 331918 402561
rect 332154 402325 332196 402561
rect 331876 395561 332196 402325
rect 331876 395325 331918 395561
rect 332154 395325 332196 395561
rect 331876 388561 332196 395325
rect 331876 388325 331918 388561
rect 332154 388325 332196 388561
rect 331876 381561 332196 388325
rect 331876 381325 331918 381561
rect 332154 381325 332196 381561
rect 331876 374561 332196 381325
rect 331876 374325 331918 374561
rect 332154 374325 332196 374561
rect 331876 367561 332196 374325
rect 331876 367325 331918 367561
rect 332154 367325 332196 367561
rect 331876 360561 332196 367325
rect 331876 360325 331918 360561
rect 332154 360325 332196 360561
rect 331876 353561 332196 360325
rect 331876 353325 331918 353561
rect 332154 353325 332196 353561
rect 331876 346561 332196 353325
rect 331876 346325 331918 346561
rect 332154 346325 332196 346561
rect 331876 339561 332196 346325
rect 331876 339325 331918 339561
rect 332154 339325 332196 339561
rect 331876 332561 332196 339325
rect 331876 332325 331918 332561
rect 332154 332325 332196 332561
rect 331876 325561 332196 332325
rect 331876 325325 331918 325561
rect 332154 325325 332196 325561
rect 331876 318561 332196 325325
rect 331876 318325 331918 318561
rect 332154 318325 332196 318561
rect 331876 311561 332196 318325
rect 331876 311325 331918 311561
rect 332154 311325 332196 311561
rect 331876 304561 332196 311325
rect 331876 304325 331918 304561
rect 332154 304325 332196 304561
rect 331876 297561 332196 304325
rect 331876 297325 331918 297561
rect 332154 297325 332196 297561
rect 331876 290561 332196 297325
rect 331876 290325 331918 290561
rect 332154 290325 332196 290561
rect 331876 283561 332196 290325
rect 331876 283325 331918 283561
rect 332154 283325 332196 283561
rect 331876 276561 332196 283325
rect 331876 276325 331918 276561
rect 332154 276325 332196 276561
rect 331876 269561 332196 276325
rect 331876 269325 331918 269561
rect 332154 269325 332196 269561
rect 331876 262561 332196 269325
rect 331876 262325 331918 262561
rect 332154 262325 332196 262561
rect 331876 255561 332196 262325
rect 331876 255325 331918 255561
rect 332154 255325 332196 255561
rect 331876 248561 332196 255325
rect 331876 248325 331918 248561
rect 332154 248325 332196 248561
rect 331876 241561 332196 248325
rect 331876 241325 331918 241561
rect 332154 241325 332196 241561
rect 331876 234561 332196 241325
rect 331876 234325 331918 234561
rect 332154 234325 332196 234561
rect 331876 227561 332196 234325
rect 331876 227325 331918 227561
rect 332154 227325 332196 227561
rect 331876 220561 332196 227325
rect 331876 220325 331918 220561
rect 332154 220325 332196 220561
rect 331876 213561 332196 220325
rect 331876 213325 331918 213561
rect 332154 213325 332196 213561
rect 331876 206561 332196 213325
rect 331876 206325 331918 206561
rect 332154 206325 332196 206561
rect 331876 199561 332196 206325
rect 331876 199325 331918 199561
rect 332154 199325 332196 199561
rect 331876 192561 332196 199325
rect 331876 192325 331918 192561
rect 332154 192325 332196 192561
rect 331876 185561 332196 192325
rect 331876 185325 331918 185561
rect 332154 185325 332196 185561
rect 331876 178561 332196 185325
rect 331876 178325 331918 178561
rect 332154 178325 332196 178561
rect 331876 171561 332196 178325
rect 331876 171325 331918 171561
rect 332154 171325 332196 171561
rect 331876 164561 332196 171325
rect 331876 164325 331918 164561
rect 332154 164325 332196 164561
rect 331876 157561 332196 164325
rect 331876 157325 331918 157561
rect 332154 157325 332196 157561
rect 331876 150561 332196 157325
rect 331876 150325 331918 150561
rect 332154 150325 332196 150561
rect 331876 143561 332196 150325
rect 331876 143325 331918 143561
rect 332154 143325 332196 143561
rect 331876 136561 332196 143325
rect 331876 136325 331918 136561
rect 332154 136325 332196 136561
rect 331876 129561 332196 136325
rect 331876 129325 331918 129561
rect 332154 129325 332196 129561
rect 331876 122561 332196 129325
rect 331876 122325 331918 122561
rect 332154 122325 332196 122561
rect 331876 115561 332196 122325
rect 331876 115325 331918 115561
rect 332154 115325 332196 115561
rect 331876 108561 332196 115325
rect 331876 108325 331918 108561
rect 332154 108325 332196 108561
rect 331876 101561 332196 108325
rect 331876 101325 331918 101561
rect 332154 101325 332196 101561
rect 331876 94561 332196 101325
rect 331876 94325 331918 94561
rect 332154 94325 332196 94561
rect 331876 87561 332196 94325
rect 331876 87325 331918 87561
rect 332154 87325 332196 87561
rect 331876 80561 332196 87325
rect 331876 80325 331918 80561
rect 332154 80325 332196 80561
rect 331876 73561 332196 80325
rect 331876 73325 331918 73561
rect 332154 73325 332196 73561
rect 331876 66561 332196 73325
rect 331876 66325 331918 66561
rect 332154 66325 332196 66561
rect 331876 59561 332196 66325
rect 331876 59325 331918 59561
rect 332154 59325 332196 59561
rect 331876 52561 332196 59325
rect 331876 52325 331918 52561
rect 332154 52325 332196 52561
rect 331876 45561 332196 52325
rect 331876 45325 331918 45561
rect 332154 45325 332196 45561
rect 331876 38561 332196 45325
rect 331876 38325 331918 38561
rect 332154 38325 332196 38561
rect 331876 31561 332196 38325
rect 331876 31325 331918 31561
rect 332154 31325 332196 31561
rect 331876 24561 332196 31325
rect 331876 24325 331918 24561
rect 332154 24325 332196 24561
rect 331876 17561 332196 24325
rect 331876 17325 331918 17561
rect 332154 17325 332196 17561
rect 331876 10561 332196 17325
rect 331876 10325 331918 10561
rect 332154 10325 332196 10561
rect 331876 3561 332196 10325
rect 331876 3325 331918 3561
rect 332154 3325 332196 3561
rect 331876 -1706 332196 3325
rect 331876 -1942 331918 -1706
rect 332154 -1942 332196 -1706
rect 331876 -2026 332196 -1942
rect 331876 -2262 331918 -2026
rect 332154 -2262 332196 -2026
rect 331876 -2294 332196 -2262
rect 337144 705238 337464 706230
rect 337144 705002 337186 705238
rect 337422 705002 337464 705238
rect 337144 704918 337464 705002
rect 337144 704682 337186 704918
rect 337422 704682 337464 704918
rect 337144 695494 337464 704682
rect 337144 695258 337186 695494
rect 337422 695258 337464 695494
rect 337144 688494 337464 695258
rect 337144 688258 337186 688494
rect 337422 688258 337464 688494
rect 337144 681494 337464 688258
rect 337144 681258 337186 681494
rect 337422 681258 337464 681494
rect 337144 674494 337464 681258
rect 337144 674258 337186 674494
rect 337422 674258 337464 674494
rect 337144 667494 337464 674258
rect 337144 667258 337186 667494
rect 337422 667258 337464 667494
rect 337144 660494 337464 667258
rect 337144 660258 337186 660494
rect 337422 660258 337464 660494
rect 337144 653494 337464 660258
rect 337144 653258 337186 653494
rect 337422 653258 337464 653494
rect 337144 646494 337464 653258
rect 337144 646258 337186 646494
rect 337422 646258 337464 646494
rect 337144 639494 337464 646258
rect 337144 639258 337186 639494
rect 337422 639258 337464 639494
rect 337144 632494 337464 639258
rect 337144 632258 337186 632494
rect 337422 632258 337464 632494
rect 337144 625494 337464 632258
rect 337144 625258 337186 625494
rect 337422 625258 337464 625494
rect 337144 618494 337464 625258
rect 337144 618258 337186 618494
rect 337422 618258 337464 618494
rect 337144 611494 337464 618258
rect 337144 611258 337186 611494
rect 337422 611258 337464 611494
rect 337144 604494 337464 611258
rect 337144 604258 337186 604494
rect 337422 604258 337464 604494
rect 337144 597494 337464 604258
rect 337144 597258 337186 597494
rect 337422 597258 337464 597494
rect 337144 590494 337464 597258
rect 337144 590258 337186 590494
rect 337422 590258 337464 590494
rect 337144 583494 337464 590258
rect 337144 583258 337186 583494
rect 337422 583258 337464 583494
rect 337144 576494 337464 583258
rect 337144 576258 337186 576494
rect 337422 576258 337464 576494
rect 337144 569494 337464 576258
rect 337144 569258 337186 569494
rect 337422 569258 337464 569494
rect 337144 562494 337464 569258
rect 337144 562258 337186 562494
rect 337422 562258 337464 562494
rect 337144 555494 337464 562258
rect 337144 555258 337186 555494
rect 337422 555258 337464 555494
rect 337144 548494 337464 555258
rect 337144 548258 337186 548494
rect 337422 548258 337464 548494
rect 337144 541494 337464 548258
rect 337144 541258 337186 541494
rect 337422 541258 337464 541494
rect 337144 534494 337464 541258
rect 337144 534258 337186 534494
rect 337422 534258 337464 534494
rect 337144 527494 337464 534258
rect 337144 527258 337186 527494
rect 337422 527258 337464 527494
rect 337144 520494 337464 527258
rect 337144 520258 337186 520494
rect 337422 520258 337464 520494
rect 337144 513494 337464 520258
rect 337144 513258 337186 513494
rect 337422 513258 337464 513494
rect 337144 506494 337464 513258
rect 337144 506258 337186 506494
rect 337422 506258 337464 506494
rect 337144 499494 337464 506258
rect 337144 499258 337186 499494
rect 337422 499258 337464 499494
rect 337144 492494 337464 499258
rect 337144 492258 337186 492494
rect 337422 492258 337464 492494
rect 337144 485494 337464 492258
rect 337144 485258 337186 485494
rect 337422 485258 337464 485494
rect 337144 478494 337464 485258
rect 337144 478258 337186 478494
rect 337422 478258 337464 478494
rect 337144 471494 337464 478258
rect 337144 471258 337186 471494
rect 337422 471258 337464 471494
rect 337144 464494 337464 471258
rect 337144 464258 337186 464494
rect 337422 464258 337464 464494
rect 337144 457494 337464 464258
rect 337144 457258 337186 457494
rect 337422 457258 337464 457494
rect 337144 450494 337464 457258
rect 337144 450258 337186 450494
rect 337422 450258 337464 450494
rect 337144 443494 337464 450258
rect 337144 443258 337186 443494
rect 337422 443258 337464 443494
rect 337144 436494 337464 443258
rect 337144 436258 337186 436494
rect 337422 436258 337464 436494
rect 337144 429494 337464 436258
rect 337144 429258 337186 429494
rect 337422 429258 337464 429494
rect 337144 422494 337464 429258
rect 337144 422258 337186 422494
rect 337422 422258 337464 422494
rect 337144 415494 337464 422258
rect 337144 415258 337186 415494
rect 337422 415258 337464 415494
rect 337144 408494 337464 415258
rect 337144 408258 337186 408494
rect 337422 408258 337464 408494
rect 337144 401494 337464 408258
rect 337144 401258 337186 401494
rect 337422 401258 337464 401494
rect 337144 394494 337464 401258
rect 337144 394258 337186 394494
rect 337422 394258 337464 394494
rect 337144 387494 337464 394258
rect 337144 387258 337186 387494
rect 337422 387258 337464 387494
rect 337144 380494 337464 387258
rect 337144 380258 337186 380494
rect 337422 380258 337464 380494
rect 337144 373494 337464 380258
rect 337144 373258 337186 373494
rect 337422 373258 337464 373494
rect 337144 366494 337464 373258
rect 337144 366258 337186 366494
rect 337422 366258 337464 366494
rect 337144 359494 337464 366258
rect 337144 359258 337186 359494
rect 337422 359258 337464 359494
rect 337144 352494 337464 359258
rect 337144 352258 337186 352494
rect 337422 352258 337464 352494
rect 337144 345494 337464 352258
rect 337144 345258 337186 345494
rect 337422 345258 337464 345494
rect 337144 338494 337464 345258
rect 337144 338258 337186 338494
rect 337422 338258 337464 338494
rect 337144 331494 337464 338258
rect 337144 331258 337186 331494
rect 337422 331258 337464 331494
rect 337144 324494 337464 331258
rect 337144 324258 337186 324494
rect 337422 324258 337464 324494
rect 337144 317494 337464 324258
rect 337144 317258 337186 317494
rect 337422 317258 337464 317494
rect 337144 310494 337464 317258
rect 337144 310258 337186 310494
rect 337422 310258 337464 310494
rect 337144 303494 337464 310258
rect 337144 303258 337186 303494
rect 337422 303258 337464 303494
rect 337144 296494 337464 303258
rect 337144 296258 337186 296494
rect 337422 296258 337464 296494
rect 337144 289494 337464 296258
rect 337144 289258 337186 289494
rect 337422 289258 337464 289494
rect 337144 282494 337464 289258
rect 337144 282258 337186 282494
rect 337422 282258 337464 282494
rect 337144 275494 337464 282258
rect 337144 275258 337186 275494
rect 337422 275258 337464 275494
rect 337144 268494 337464 275258
rect 337144 268258 337186 268494
rect 337422 268258 337464 268494
rect 337144 261494 337464 268258
rect 337144 261258 337186 261494
rect 337422 261258 337464 261494
rect 337144 254494 337464 261258
rect 337144 254258 337186 254494
rect 337422 254258 337464 254494
rect 337144 247494 337464 254258
rect 337144 247258 337186 247494
rect 337422 247258 337464 247494
rect 337144 240494 337464 247258
rect 337144 240258 337186 240494
rect 337422 240258 337464 240494
rect 337144 233494 337464 240258
rect 337144 233258 337186 233494
rect 337422 233258 337464 233494
rect 337144 226494 337464 233258
rect 337144 226258 337186 226494
rect 337422 226258 337464 226494
rect 337144 219494 337464 226258
rect 337144 219258 337186 219494
rect 337422 219258 337464 219494
rect 337144 212494 337464 219258
rect 337144 212258 337186 212494
rect 337422 212258 337464 212494
rect 337144 205494 337464 212258
rect 337144 205258 337186 205494
rect 337422 205258 337464 205494
rect 337144 198494 337464 205258
rect 337144 198258 337186 198494
rect 337422 198258 337464 198494
rect 337144 191494 337464 198258
rect 337144 191258 337186 191494
rect 337422 191258 337464 191494
rect 337144 184494 337464 191258
rect 337144 184258 337186 184494
rect 337422 184258 337464 184494
rect 337144 177494 337464 184258
rect 337144 177258 337186 177494
rect 337422 177258 337464 177494
rect 337144 170494 337464 177258
rect 337144 170258 337186 170494
rect 337422 170258 337464 170494
rect 337144 163494 337464 170258
rect 337144 163258 337186 163494
rect 337422 163258 337464 163494
rect 337144 156494 337464 163258
rect 337144 156258 337186 156494
rect 337422 156258 337464 156494
rect 337144 149494 337464 156258
rect 337144 149258 337186 149494
rect 337422 149258 337464 149494
rect 337144 142494 337464 149258
rect 337144 142258 337186 142494
rect 337422 142258 337464 142494
rect 337144 135494 337464 142258
rect 337144 135258 337186 135494
rect 337422 135258 337464 135494
rect 337144 128494 337464 135258
rect 337144 128258 337186 128494
rect 337422 128258 337464 128494
rect 337144 121494 337464 128258
rect 337144 121258 337186 121494
rect 337422 121258 337464 121494
rect 337144 114494 337464 121258
rect 337144 114258 337186 114494
rect 337422 114258 337464 114494
rect 337144 107494 337464 114258
rect 337144 107258 337186 107494
rect 337422 107258 337464 107494
rect 337144 100494 337464 107258
rect 337144 100258 337186 100494
rect 337422 100258 337464 100494
rect 337144 93494 337464 100258
rect 337144 93258 337186 93494
rect 337422 93258 337464 93494
rect 337144 86494 337464 93258
rect 337144 86258 337186 86494
rect 337422 86258 337464 86494
rect 337144 79494 337464 86258
rect 337144 79258 337186 79494
rect 337422 79258 337464 79494
rect 337144 72494 337464 79258
rect 337144 72258 337186 72494
rect 337422 72258 337464 72494
rect 337144 65494 337464 72258
rect 337144 65258 337186 65494
rect 337422 65258 337464 65494
rect 337144 58494 337464 65258
rect 337144 58258 337186 58494
rect 337422 58258 337464 58494
rect 337144 51494 337464 58258
rect 337144 51258 337186 51494
rect 337422 51258 337464 51494
rect 337144 44494 337464 51258
rect 337144 44258 337186 44494
rect 337422 44258 337464 44494
rect 337144 37494 337464 44258
rect 337144 37258 337186 37494
rect 337422 37258 337464 37494
rect 337144 30494 337464 37258
rect 337144 30258 337186 30494
rect 337422 30258 337464 30494
rect 337144 23494 337464 30258
rect 337144 23258 337186 23494
rect 337422 23258 337464 23494
rect 337144 16494 337464 23258
rect 337144 16258 337186 16494
rect 337422 16258 337464 16494
rect 337144 9494 337464 16258
rect 337144 9258 337186 9494
rect 337422 9258 337464 9494
rect 337144 2494 337464 9258
rect 337144 2258 337186 2494
rect 337422 2258 337464 2494
rect 337144 -746 337464 2258
rect 337144 -982 337186 -746
rect 337422 -982 337464 -746
rect 337144 -1066 337464 -982
rect 337144 -1302 337186 -1066
rect 337422 -1302 337464 -1066
rect 337144 -2294 337464 -1302
rect 338876 706198 339196 706230
rect 338876 705962 338918 706198
rect 339154 705962 339196 706198
rect 338876 705878 339196 705962
rect 338876 705642 338918 705878
rect 339154 705642 339196 705878
rect 338876 696561 339196 705642
rect 338876 696325 338918 696561
rect 339154 696325 339196 696561
rect 338876 689561 339196 696325
rect 338876 689325 338918 689561
rect 339154 689325 339196 689561
rect 338876 682561 339196 689325
rect 338876 682325 338918 682561
rect 339154 682325 339196 682561
rect 338876 675561 339196 682325
rect 338876 675325 338918 675561
rect 339154 675325 339196 675561
rect 338876 668561 339196 675325
rect 338876 668325 338918 668561
rect 339154 668325 339196 668561
rect 338876 661561 339196 668325
rect 338876 661325 338918 661561
rect 339154 661325 339196 661561
rect 338876 654561 339196 661325
rect 338876 654325 338918 654561
rect 339154 654325 339196 654561
rect 338876 647561 339196 654325
rect 338876 647325 338918 647561
rect 339154 647325 339196 647561
rect 338876 640561 339196 647325
rect 338876 640325 338918 640561
rect 339154 640325 339196 640561
rect 338876 633561 339196 640325
rect 338876 633325 338918 633561
rect 339154 633325 339196 633561
rect 338876 626561 339196 633325
rect 338876 626325 338918 626561
rect 339154 626325 339196 626561
rect 338876 619561 339196 626325
rect 338876 619325 338918 619561
rect 339154 619325 339196 619561
rect 338876 612561 339196 619325
rect 338876 612325 338918 612561
rect 339154 612325 339196 612561
rect 338876 605561 339196 612325
rect 338876 605325 338918 605561
rect 339154 605325 339196 605561
rect 338876 598561 339196 605325
rect 338876 598325 338918 598561
rect 339154 598325 339196 598561
rect 338876 591561 339196 598325
rect 338876 591325 338918 591561
rect 339154 591325 339196 591561
rect 338876 584561 339196 591325
rect 338876 584325 338918 584561
rect 339154 584325 339196 584561
rect 338876 577561 339196 584325
rect 338876 577325 338918 577561
rect 339154 577325 339196 577561
rect 338876 570561 339196 577325
rect 338876 570325 338918 570561
rect 339154 570325 339196 570561
rect 338876 563561 339196 570325
rect 338876 563325 338918 563561
rect 339154 563325 339196 563561
rect 338876 556561 339196 563325
rect 338876 556325 338918 556561
rect 339154 556325 339196 556561
rect 338876 549561 339196 556325
rect 338876 549325 338918 549561
rect 339154 549325 339196 549561
rect 338876 542561 339196 549325
rect 338876 542325 338918 542561
rect 339154 542325 339196 542561
rect 338876 535561 339196 542325
rect 338876 535325 338918 535561
rect 339154 535325 339196 535561
rect 338876 528561 339196 535325
rect 338876 528325 338918 528561
rect 339154 528325 339196 528561
rect 338876 521561 339196 528325
rect 338876 521325 338918 521561
rect 339154 521325 339196 521561
rect 338876 514561 339196 521325
rect 338876 514325 338918 514561
rect 339154 514325 339196 514561
rect 338876 507561 339196 514325
rect 338876 507325 338918 507561
rect 339154 507325 339196 507561
rect 338876 500561 339196 507325
rect 338876 500325 338918 500561
rect 339154 500325 339196 500561
rect 338876 493561 339196 500325
rect 338876 493325 338918 493561
rect 339154 493325 339196 493561
rect 338876 486561 339196 493325
rect 338876 486325 338918 486561
rect 339154 486325 339196 486561
rect 338876 479561 339196 486325
rect 338876 479325 338918 479561
rect 339154 479325 339196 479561
rect 338876 472561 339196 479325
rect 338876 472325 338918 472561
rect 339154 472325 339196 472561
rect 338876 465561 339196 472325
rect 338876 465325 338918 465561
rect 339154 465325 339196 465561
rect 338876 458561 339196 465325
rect 338876 458325 338918 458561
rect 339154 458325 339196 458561
rect 338876 451561 339196 458325
rect 338876 451325 338918 451561
rect 339154 451325 339196 451561
rect 338876 444561 339196 451325
rect 338876 444325 338918 444561
rect 339154 444325 339196 444561
rect 338876 437561 339196 444325
rect 338876 437325 338918 437561
rect 339154 437325 339196 437561
rect 338876 430561 339196 437325
rect 338876 430325 338918 430561
rect 339154 430325 339196 430561
rect 338876 423561 339196 430325
rect 338876 423325 338918 423561
rect 339154 423325 339196 423561
rect 338876 416561 339196 423325
rect 338876 416325 338918 416561
rect 339154 416325 339196 416561
rect 338876 409561 339196 416325
rect 338876 409325 338918 409561
rect 339154 409325 339196 409561
rect 338876 402561 339196 409325
rect 338876 402325 338918 402561
rect 339154 402325 339196 402561
rect 338876 395561 339196 402325
rect 338876 395325 338918 395561
rect 339154 395325 339196 395561
rect 338876 388561 339196 395325
rect 338876 388325 338918 388561
rect 339154 388325 339196 388561
rect 338876 381561 339196 388325
rect 338876 381325 338918 381561
rect 339154 381325 339196 381561
rect 338876 374561 339196 381325
rect 338876 374325 338918 374561
rect 339154 374325 339196 374561
rect 338876 367561 339196 374325
rect 338876 367325 338918 367561
rect 339154 367325 339196 367561
rect 338876 360561 339196 367325
rect 338876 360325 338918 360561
rect 339154 360325 339196 360561
rect 338876 353561 339196 360325
rect 338876 353325 338918 353561
rect 339154 353325 339196 353561
rect 338876 346561 339196 353325
rect 338876 346325 338918 346561
rect 339154 346325 339196 346561
rect 338876 339561 339196 346325
rect 338876 339325 338918 339561
rect 339154 339325 339196 339561
rect 338876 332561 339196 339325
rect 338876 332325 338918 332561
rect 339154 332325 339196 332561
rect 338876 325561 339196 332325
rect 338876 325325 338918 325561
rect 339154 325325 339196 325561
rect 338876 318561 339196 325325
rect 338876 318325 338918 318561
rect 339154 318325 339196 318561
rect 338876 311561 339196 318325
rect 338876 311325 338918 311561
rect 339154 311325 339196 311561
rect 338876 304561 339196 311325
rect 338876 304325 338918 304561
rect 339154 304325 339196 304561
rect 338876 297561 339196 304325
rect 338876 297325 338918 297561
rect 339154 297325 339196 297561
rect 338876 290561 339196 297325
rect 338876 290325 338918 290561
rect 339154 290325 339196 290561
rect 338876 283561 339196 290325
rect 338876 283325 338918 283561
rect 339154 283325 339196 283561
rect 338876 276561 339196 283325
rect 338876 276325 338918 276561
rect 339154 276325 339196 276561
rect 338876 269561 339196 276325
rect 338876 269325 338918 269561
rect 339154 269325 339196 269561
rect 338876 262561 339196 269325
rect 338876 262325 338918 262561
rect 339154 262325 339196 262561
rect 338876 255561 339196 262325
rect 338876 255325 338918 255561
rect 339154 255325 339196 255561
rect 338876 248561 339196 255325
rect 338876 248325 338918 248561
rect 339154 248325 339196 248561
rect 338876 241561 339196 248325
rect 338876 241325 338918 241561
rect 339154 241325 339196 241561
rect 338876 234561 339196 241325
rect 338876 234325 338918 234561
rect 339154 234325 339196 234561
rect 338876 227561 339196 234325
rect 338876 227325 338918 227561
rect 339154 227325 339196 227561
rect 338876 220561 339196 227325
rect 338876 220325 338918 220561
rect 339154 220325 339196 220561
rect 338876 213561 339196 220325
rect 338876 213325 338918 213561
rect 339154 213325 339196 213561
rect 338876 206561 339196 213325
rect 338876 206325 338918 206561
rect 339154 206325 339196 206561
rect 338876 199561 339196 206325
rect 338876 199325 338918 199561
rect 339154 199325 339196 199561
rect 338876 192561 339196 199325
rect 338876 192325 338918 192561
rect 339154 192325 339196 192561
rect 338876 185561 339196 192325
rect 338876 185325 338918 185561
rect 339154 185325 339196 185561
rect 338876 178561 339196 185325
rect 338876 178325 338918 178561
rect 339154 178325 339196 178561
rect 338876 171561 339196 178325
rect 338876 171325 338918 171561
rect 339154 171325 339196 171561
rect 338876 164561 339196 171325
rect 338876 164325 338918 164561
rect 339154 164325 339196 164561
rect 338876 157561 339196 164325
rect 338876 157325 338918 157561
rect 339154 157325 339196 157561
rect 338876 150561 339196 157325
rect 338876 150325 338918 150561
rect 339154 150325 339196 150561
rect 338876 143561 339196 150325
rect 338876 143325 338918 143561
rect 339154 143325 339196 143561
rect 338876 136561 339196 143325
rect 338876 136325 338918 136561
rect 339154 136325 339196 136561
rect 338876 129561 339196 136325
rect 338876 129325 338918 129561
rect 339154 129325 339196 129561
rect 338876 122561 339196 129325
rect 338876 122325 338918 122561
rect 339154 122325 339196 122561
rect 338876 115561 339196 122325
rect 338876 115325 338918 115561
rect 339154 115325 339196 115561
rect 338876 108561 339196 115325
rect 338876 108325 338918 108561
rect 339154 108325 339196 108561
rect 338876 101561 339196 108325
rect 338876 101325 338918 101561
rect 339154 101325 339196 101561
rect 338876 94561 339196 101325
rect 338876 94325 338918 94561
rect 339154 94325 339196 94561
rect 338876 87561 339196 94325
rect 338876 87325 338918 87561
rect 339154 87325 339196 87561
rect 338876 80561 339196 87325
rect 338876 80325 338918 80561
rect 339154 80325 339196 80561
rect 338876 73561 339196 80325
rect 338876 73325 338918 73561
rect 339154 73325 339196 73561
rect 338876 66561 339196 73325
rect 338876 66325 338918 66561
rect 339154 66325 339196 66561
rect 338876 59561 339196 66325
rect 338876 59325 338918 59561
rect 339154 59325 339196 59561
rect 338876 52561 339196 59325
rect 338876 52325 338918 52561
rect 339154 52325 339196 52561
rect 338876 45561 339196 52325
rect 338876 45325 338918 45561
rect 339154 45325 339196 45561
rect 338876 38561 339196 45325
rect 338876 38325 338918 38561
rect 339154 38325 339196 38561
rect 338876 31561 339196 38325
rect 338876 31325 338918 31561
rect 339154 31325 339196 31561
rect 338876 24561 339196 31325
rect 338876 24325 338918 24561
rect 339154 24325 339196 24561
rect 338876 17561 339196 24325
rect 338876 17325 338918 17561
rect 339154 17325 339196 17561
rect 338876 10561 339196 17325
rect 338876 10325 338918 10561
rect 339154 10325 339196 10561
rect 338876 3561 339196 10325
rect 338876 3325 338918 3561
rect 339154 3325 339196 3561
rect 338876 -1706 339196 3325
rect 338876 -1942 338918 -1706
rect 339154 -1942 339196 -1706
rect 338876 -2026 339196 -1942
rect 338876 -2262 338918 -2026
rect 339154 -2262 339196 -2026
rect 338876 -2294 339196 -2262
rect 344144 705238 344464 706230
rect 344144 705002 344186 705238
rect 344422 705002 344464 705238
rect 344144 704918 344464 705002
rect 344144 704682 344186 704918
rect 344422 704682 344464 704918
rect 344144 695494 344464 704682
rect 344144 695258 344186 695494
rect 344422 695258 344464 695494
rect 344144 688494 344464 695258
rect 344144 688258 344186 688494
rect 344422 688258 344464 688494
rect 344144 681494 344464 688258
rect 344144 681258 344186 681494
rect 344422 681258 344464 681494
rect 344144 674494 344464 681258
rect 344144 674258 344186 674494
rect 344422 674258 344464 674494
rect 344144 667494 344464 674258
rect 344144 667258 344186 667494
rect 344422 667258 344464 667494
rect 344144 660494 344464 667258
rect 344144 660258 344186 660494
rect 344422 660258 344464 660494
rect 344144 653494 344464 660258
rect 344144 653258 344186 653494
rect 344422 653258 344464 653494
rect 344144 646494 344464 653258
rect 344144 646258 344186 646494
rect 344422 646258 344464 646494
rect 344144 639494 344464 646258
rect 344144 639258 344186 639494
rect 344422 639258 344464 639494
rect 344144 632494 344464 639258
rect 344144 632258 344186 632494
rect 344422 632258 344464 632494
rect 344144 625494 344464 632258
rect 344144 625258 344186 625494
rect 344422 625258 344464 625494
rect 344144 618494 344464 625258
rect 344144 618258 344186 618494
rect 344422 618258 344464 618494
rect 344144 611494 344464 618258
rect 344144 611258 344186 611494
rect 344422 611258 344464 611494
rect 344144 604494 344464 611258
rect 344144 604258 344186 604494
rect 344422 604258 344464 604494
rect 344144 597494 344464 604258
rect 344144 597258 344186 597494
rect 344422 597258 344464 597494
rect 344144 590494 344464 597258
rect 344144 590258 344186 590494
rect 344422 590258 344464 590494
rect 344144 583494 344464 590258
rect 344144 583258 344186 583494
rect 344422 583258 344464 583494
rect 344144 576494 344464 583258
rect 344144 576258 344186 576494
rect 344422 576258 344464 576494
rect 344144 569494 344464 576258
rect 344144 569258 344186 569494
rect 344422 569258 344464 569494
rect 344144 562494 344464 569258
rect 344144 562258 344186 562494
rect 344422 562258 344464 562494
rect 344144 555494 344464 562258
rect 344144 555258 344186 555494
rect 344422 555258 344464 555494
rect 344144 548494 344464 555258
rect 344144 548258 344186 548494
rect 344422 548258 344464 548494
rect 344144 541494 344464 548258
rect 344144 541258 344186 541494
rect 344422 541258 344464 541494
rect 344144 534494 344464 541258
rect 344144 534258 344186 534494
rect 344422 534258 344464 534494
rect 344144 527494 344464 534258
rect 344144 527258 344186 527494
rect 344422 527258 344464 527494
rect 344144 520494 344464 527258
rect 344144 520258 344186 520494
rect 344422 520258 344464 520494
rect 344144 513494 344464 520258
rect 344144 513258 344186 513494
rect 344422 513258 344464 513494
rect 344144 506494 344464 513258
rect 344144 506258 344186 506494
rect 344422 506258 344464 506494
rect 344144 499494 344464 506258
rect 344144 499258 344186 499494
rect 344422 499258 344464 499494
rect 344144 492494 344464 499258
rect 344144 492258 344186 492494
rect 344422 492258 344464 492494
rect 344144 485494 344464 492258
rect 344144 485258 344186 485494
rect 344422 485258 344464 485494
rect 344144 478494 344464 485258
rect 344144 478258 344186 478494
rect 344422 478258 344464 478494
rect 344144 471494 344464 478258
rect 344144 471258 344186 471494
rect 344422 471258 344464 471494
rect 344144 464494 344464 471258
rect 344144 464258 344186 464494
rect 344422 464258 344464 464494
rect 344144 457494 344464 464258
rect 344144 457258 344186 457494
rect 344422 457258 344464 457494
rect 344144 450494 344464 457258
rect 344144 450258 344186 450494
rect 344422 450258 344464 450494
rect 344144 443494 344464 450258
rect 344144 443258 344186 443494
rect 344422 443258 344464 443494
rect 344144 436494 344464 443258
rect 344144 436258 344186 436494
rect 344422 436258 344464 436494
rect 344144 429494 344464 436258
rect 344144 429258 344186 429494
rect 344422 429258 344464 429494
rect 344144 422494 344464 429258
rect 344144 422258 344186 422494
rect 344422 422258 344464 422494
rect 344144 415494 344464 422258
rect 344144 415258 344186 415494
rect 344422 415258 344464 415494
rect 344144 408494 344464 415258
rect 344144 408258 344186 408494
rect 344422 408258 344464 408494
rect 344144 401494 344464 408258
rect 344144 401258 344186 401494
rect 344422 401258 344464 401494
rect 344144 394494 344464 401258
rect 344144 394258 344186 394494
rect 344422 394258 344464 394494
rect 344144 387494 344464 394258
rect 344144 387258 344186 387494
rect 344422 387258 344464 387494
rect 344144 380494 344464 387258
rect 344144 380258 344186 380494
rect 344422 380258 344464 380494
rect 344144 373494 344464 380258
rect 344144 373258 344186 373494
rect 344422 373258 344464 373494
rect 344144 366494 344464 373258
rect 344144 366258 344186 366494
rect 344422 366258 344464 366494
rect 344144 359494 344464 366258
rect 344144 359258 344186 359494
rect 344422 359258 344464 359494
rect 344144 352494 344464 359258
rect 344144 352258 344186 352494
rect 344422 352258 344464 352494
rect 344144 345494 344464 352258
rect 344144 345258 344186 345494
rect 344422 345258 344464 345494
rect 344144 338494 344464 345258
rect 344144 338258 344186 338494
rect 344422 338258 344464 338494
rect 344144 331494 344464 338258
rect 344144 331258 344186 331494
rect 344422 331258 344464 331494
rect 344144 324494 344464 331258
rect 344144 324258 344186 324494
rect 344422 324258 344464 324494
rect 344144 317494 344464 324258
rect 344144 317258 344186 317494
rect 344422 317258 344464 317494
rect 344144 310494 344464 317258
rect 344144 310258 344186 310494
rect 344422 310258 344464 310494
rect 344144 303494 344464 310258
rect 344144 303258 344186 303494
rect 344422 303258 344464 303494
rect 344144 296494 344464 303258
rect 344144 296258 344186 296494
rect 344422 296258 344464 296494
rect 344144 289494 344464 296258
rect 344144 289258 344186 289494
rect 344422 289258 344464 289494
rect 344144 282494 344464 289258
rect 344144 282258 344186 282494
rect 344422 282258 344464 282494
rect 344144 275494 344464 282258
rect 344144 275258 344186 275494
rect 344422 275258 344464 275494
rect 344144 268494 344464 275258
rect 344144 268258 344186 268494
rect 344422 268258 344464 268494
rect 344144 261494 344464 268258
rect 344144 261258 344186 261494
rect 344422 261258 344464 261494
rect 344144 254494 344464 261258
rect 344144 254258 344186 254494
rect 344422 254258 344464 254494
rect 344144 247494 344464 254258
rect 344144 247258 344186 247494
rect 344422 247258 344464 247494
rect 344144 240494 344464 247258
rect 344144 240258 344186 240494
rect 344422 240258 344464 240494
rect 344144 233494 344464 240258
rect 344144 233258 344186 233494
rect 344422 233258 344464 233494
rect 344144 226494 344464 233258
rect 344144 226258 344186 226494
rect 344422 226258 344464 226494
rect 344144 219494 344464 226258
rect 344144 219258 344186 219494
rect 344422 219258 344464 219494
rect 344144 212494 344464 219258
rect 344144 212258 344186 212494
rect 344422 212258 344464 212494
rect 344144 205494 344464 212258
rect 344144 205258 344186 205494
rect 344422 205258 344464 205494
rect 344144 198494 344464 205258
rect 344144 198258 344186 198494
rect 344422 198258 344464 198494
rect 344144 191494 344464 198258
rect 344144 191258 344186 191494
rect 344422 191258 344464 191494
rect 344144 184494 344464 191258
rect 344144 184258 344186 184494
rect 344422 184258 344464 184494
rect 344144 177494 344464 184258
rect 344144 177258 344186 177494
rect 344422 177258 344464 177494
rect 344144 170494 344464 177258
rect 344144 170258 344186 170494
rect 344422 170258 344464 170494
rect 344144 163494 344464 170258
rect 344144 163258 344186 163494
rect 344422 163258 344464 163494
rect 344144 156494 344464 163258
rect 344144 156258 344186 156494
rect 344422 156258 344464 156494
rect 344144 149494 344464 156258
rect 344144 149258 344186 149494
rect 344422 149258 344464 149494
rect 344144 142494 344464 149258
rect 344144 142258 344186 142494
rect 344422 142258 344464 142494
rect 344144 135494 344464 142258
rect 344144 135258 344186 135494
rect 344422 135258 344464 135494
rect 344144 128494 344464 135258
rect 344144 128258 344186 128494
rect 344422 128258 344464 128494
rect 344144 121494 344464 128258
rect 344144 121258 344186 121494
rect 344422 121258 344464 121494
rect 344144 114494 344464 121258
rect 344144 114258 344186 114494
rect 344422 114258 344464 114494
rect 344144 107494 344464 114258
rect 344144 107258 344186 107494
rect 344422 107258 344464 107494
rect 344144 100494 344464 107258
rect 344144 100258 344186 100494
rect 344422 100258 344464 100494
rect 344144 93494 344464 100258
rect 344144 93258 344186 93494
rect 344422 93258 344464 93494
rect 344144 86494 344464 93258
rect 344144 86258 344186 86494
rect 344422 86258 344464 86494
rect 344144 79494 344464 86258
rect 344144 79258 344186 79494
rect 344422 79258 344464 79494
rect 344144 72494 344464 79258
rect 344144 72258 344186 72494
rect 344422 72258 344464 72494
rect 344144 65494 344464 72258
rect 344144 65258 344186 65494
rect 344422 65258 344464 65494
rect 344144 58494 344464 65258
rect 344144 58258 344186 58494
rect 344422 58258 344464 58494
rect 344144 51494 344464 58258
rect 344144 51258 344186 51494
rect 344422 51258 344464 51494
rect 344144 44494 344464 51258
rect 344144 44258 344186 44494
rect 344422 44258 344464 44494
rect 344144 37494 344464 44258
rect 344144 37258 344186 37494
rect 344422 37258 344464 37494
rect 344144 30494 344464 37258
rect 344144 30258 344186 30494
rect 344422 30258 344464 30494
rect 344144 23494 344464 30258
rect 344144 23258 344186 23494
rect 344422 23258 344464 23494
rect 344144 16494 344464 23258
rect 344144 16258 344186 16494
rect 344422 16258 344464 16494
rect 344144 9494 344464 16258
rect 344144 9258 344186 9494
rect 344422 9258 344464 9494
rect 344144 2494 344464 9258
rect 344144 2258 344186 2494
rect 344422 2258 344464 2494
rect 344144 -746 344464 2258
rect 344144 -982 344186 -746
rect 344422 -982 344464 -746
rect 344144 -1066 344464 -982
rect 344144 -1302 344186 -1066
rect 344422 -1302 344464 -1066
rect 344144 -2294 344464 -1302
rect 345876 706198 346196 706230
rect 345876 705962 345918 706198
rect 346154 705962 346196 706198
rect 345876 705878 346196 705962
rect 345876 705642 345918 705878
rect 346154 705642 346196 705878
rect 345876 696561 346196 705642
rect 345876 696325 345918 696561
rect 346154 696325 346196 696561
rect 345876 689561 346196 696325
rect 345876 689325 345918 689561
rect 346154 689325 346196 689561
rect 345876 682561 346196 689325
rect 345876 682325 345918 682561
rect 346154 682325 346196 682561
rect 345876 675561 346196 682325
rect 345876 675325 345918 675561
rect 346154 675325 346196 675561
rect 345876 668561 346196 675325
rect 345876 668325 345918 668561
rect 346154 668325 346196 668561
rect 345876 661561 346196 668325
rect 345876 661325 345918 661561
rect 346154 661325 346196 661561
rect 345876 654561 346196 661325
rect 345876 654325 345918 654561
rect 346154 654325 346196 654561
rect 345876 647561 346196 654325
rect 345876 647325 345918 647561
rect 346154 647325 346196 647561
rect 345876 640561 346196 647325
rect 345876 640325 345918 640561
rect 346154 640325 346196 640561
rect 345876 633561 346196 640325
rect 345876 633325 345918 633561
rect 346154 633325 346196 633561
rect 345876 626561 346196 633325
rect 345876 626325 345918 626561
rect 346154 626325 346196 626561
rect 345876 619561 346196 626325
rect 345876 619325 345918 619561
rect 346154 619325 346196 619561
rect 345876 612561 346196 619325
rect 345876 612325 345918 612561
rect 346154 612325 346196 612561
rect 345876 605561 346196 612325
rect 345876 605325 345918 605561
rect 346154 605325 346196 605561
rect 345876 598561 346196 605325
rect 345876 598325 345918 598561
rect 346154 598325 346196 598561
rect 345876 591561 346196 598325
rect 345876 591325 345918 591561
rect 346154 591325 346196 591561
rect 345876 584561 346196 591325
rect 345876 584325 345918 584561
rect 346154 584325 346196 584561
rect 345876 577561 346196 584325
rect 345876 577325 345918 577561
rect 346154 577325 346196 577561
rect 345876 570561 346196 577325
rect 345876 570325 345918 570561
rect 346154 570325 346196 570561
rect 345876 563561 346196 570325
rect 345876 563325 345918 563561
rect 346154 563325 346196 563561
rect 345876 556561 346196 563325
rect 345876 556325 345918 556561
rect 346154 556325 346196 556561
rect 345876 549561 346196 556325
rect 345876 549325 345918 549561
rect 346154 549325 346196 549561
rect 345876 542561 346196 549325
rect 345876 542325 345918 542561
rect 346154 542325 346196 542561
rect 345876 535561 346196 542325
rect 345876 535325 345918 535561
rect 346154 535325 346196 535561
rect 345876 528561 346196 535325
rect 345876 528325 345918 528561
rect 346154 528325 346196 528561
rect 345876 521561 346196 528325
rect 345876 521325 345918 521561
rect 346154 521325 346196 521561
rect 345876 514561 346196 521325
rect 345876 514325 345918 514561
rect 346154 514325 346196 514561
rect 345876 507561 346196 514325
rect 345876 507325 345918 507561
rect 346154 507325 346196 507561
rect 345876 500561 346196 507325
rect 345876 500325 345918 500561
rect 346154 500325 346196 500561
rect 345876 493561 346196 500325
rect 345876 493325 345918 493561
rect 346154 493325 346196 493561
rect 345876 486561 346196 493325
rect 345876 486325 345918 486561
rect 346154 486325 346196 486561
rect 345876 479561 346196 486325
rect 345876 479325 345918 479561
rect 346154 479325 346196 479561
rect 345876 472561 346196 479325
rect 345876 472325 345918 472561
rect 346154 472325 346196 472561
rect 345876 465561 346196 472325
rect 345876 465325 345918 465561
rect 346154 465325 346196 465561
rect 345876 458561 346196 465325
rect 345876 458325 345918 458561
rect 346154 458325 346196 458561
rect 345876 451561 346196 458325
rect 345876 451325 345918 451561
rect 346154 451325 346196 451561
rect 345876 444561 346196 451325
rect 345876 444325 345918 444561
rect 346154 444325 346196 444561
rect 345876 437561 346196 444325
rect 345876 437325 345918 437561
rect 346154 437325 346196 437561
rect 345876 430561 346196 437325
rect 345876 430325 345918 430561
rect 346154 430325 346196 430561
rect 345876 423561 346196 430325
rect 345876 423325 345918 423561
rect 346154 423325 346196 423561
rect 345876 416561 346196 423325
rect 345876 416325 345918 416561
rect 346154 416325 346196 416561
rect 345876 409561 346196 416325
rect 345876 409325 345918 409561
rect 346154 409325 346196 409561
rect 345876 402561 346196 409325
rect 345876 402325 345918 402561
rect 346154 402325 346196 402561
rect 345876 395561 346196 402325
rect 345876 395325 345918 395561
rect 346154 395325 346196 395561
rect 345876 388561 346196 395325
rect 345876 388325 345918 388561
rect 346154 388325 346196 388561
rect 345876 381561 346196 388325
rect 345876 381325 345918 381561
rect 346154 381325 346196 381561
rect 345876 374561 346196 381325
rect 345876 374325 345918 374561
rect 346154 374325 346196 374561
rect 345876 367561 346196 374325
rect 345876 367325 345918 367561
rect 346154 367325 346196 367561
rect 345876 360561 346196 367325
rect 345876 360325 345918 360561
rect 346154 360325 346196 360561
rect 345876 353561 346196 360325
rect 345876 353325 345918 353561
rect 346154 353325 346196 353561
rect 345876 346561 346196 353325
rect 345876 346325 345918 346561
rect 346154 346325 346196 346561
rect 345876 339561 346196 346325
rect 345876 339325 345918 339561
rect 346154 339325 346196 339561
rect 345876 332561 346196 339325
rect 345876 332325 345918 332561
rect 346154 332325 346196 332561
rect 345876 325561 346196 332325
rect 345876 325325 345918 325561
rect 346154 325325 346196 325561
rect 345876 318561 346196 325325
rect 345876 318325 345918 318561
rect 346154 318325 346196 318561
rect 345876 311561 346196 318325
rect 345876 311325 345918 311561
rect 346154 311325 346196 311561
rect 345876 304561 346196 311325
rect 345876 304325 345918 304561
rect 346154 304325 346196 304561
rect 345876 297561 346196 304325
rect 345876 297325 345918 297561
rect 346154 297325 346196 297561
rect 345876 290561 346196 297325
rect 345876 290325 345918 290561
rect 346154 290325 346196 290561
rect 345876 283561 346196 290325
rect 345876 283325 345918 283561
rect 346154 283325 346196 283561
rect 345876 276561 346196 283325
rect 345876 276325 345918 276561
rect 346154 276325 346196 276561
rect 345876 269561 346196 276325
rect 345876 269325 345918 269561
rect 346154 269325 346196 269561
rect 345876 262561 346196 269325
rect 345876 262325 345918 262561
rect 346154 262325 346196 262561
rect 345876 255561 346196 262325
rect 345876 255325 345918 255561
rect 346154 255325 346196 255561
rect 345876 248561 346196 255325
rect 345876 248325 345918 248561
rect 346154 248325 346196 248561
rect 345876 241561 346196 248325
rect 345876 241325 345918 241561
rect 346154 241325 346196 241561
rect 345876 234561 346196 241325
rect 345876 234325 345918 234561
rect 346154 234325 346196 234561
rect 345876 227561 346196 234325
rect 345876 227325 345918 227561
rect 346154 227325 346196 227561
rect 345876 220561 346196 227325
rect 345876 220325 345918 220561
rect 346154 220325 346196 220561
rect 345876 213561 346196 220325
rect 345876 213325 345918 213561
rect 346154 213325 346196 213561
rect 345876 206561 346196 213325
rect 345876 206325 345918 206561
rect 346154 206325 346196 206561
rect 345876 199561 346196 206325
rect 345876 199325 345918 199561
rect 346154 199325 346196 199561
rect 345876 192561 346196 199325
rect 345876 192325 345918 192561
rect 346154 192325 346196 192561
rect 345876 185561 346196 192325
rect 345876 185325 345918 185561
rect 346154 185325 346196 185561
rect 345876 178561 346196 185325
rect 345876 178325 345918 178561
rect 346154 178325 346196 178561
rect 345876 171561 346196 178325
rect 345876 171325 345918 171561
rect 346154 171325 346196 171561
rect 345876 164561 346196 171325
rect 345876 164325 345918 164561
rect 346154 164325 346196 164561
rect 345876 157561 346196 164325
rect 345876 157325 345918 157561
rect 346154 157325 346196 157561
rect 345876 150561 346196 157325
rect 345876 150325 345918 150561
rect 346154 150325 346196 150561
rect 345876 143561 346196 150325
rect 345876 143325 345918 143561
rect 346154 143325 346196 143561
rect 345876 136561 346196 143325
rect 345876 136325 345918 136561
rect 346154 136325 346196 136561
rect 345876 129561 346196 136325
rect 345876 129325 345918 129561
rect 346154 129325 346196 129561
rect 345876 122561 346196 129325
rect 345876 122325 345918 122561
rect 346154 122325 346196 122561
rect 345876 115561 346196 122325
rect 345876 115325 345918 115561
rect 346154 115325 346196 115561
rect 345876 108561 346196 115325
rect 345876 108325 345918 108561
rect 346154 108325 346196 108561
rect 345876 101561 346196 108325
rect 345876 101325 345918 101561
rect 346154 101325 346196 101561
rect 345876 94561 346196 101325
rect 345876 94325 345918 94561
rect 346154 94325 346196 94561
rect 345876 87561 346196 94325
rect 345876 87325 345918 87561
rect 346154 87325 346196 87561
rect 345876 80561 346196 87325
rect 345876 80325 345918 80561
rect 346154 80325 346196 80561
rect 345876 73561 346196 80325
rect 345876 73325 345918 73561
rect 346154 73325 346196 73561
rect 345876 66561 346196 73325
rect 345876 66325 345918 66561
rect 346154 66325 346196 66561
rect 345876 59561 346196 66325
rect 345876 59325 345918 59561
rect 346154 59325 346196 59561
rect 345876 52561 346196 59325
rect 345876 52325 345918 52561
rect 346154 52325 346196 52561
rect 345876 45561 346196 52325
rect 345876 45325 345918 45561
rect 346154 45325 346196 45561
rect 345876 38561 346196 45325
rect 345876 38325 345918 38561
rect 346154 38325 346196 38561
rect 345876 31561 346196 38325
rect 345876 31325 345918 31561
rect 346154 31325 346196 31561
rect 345876 24561 346196 31325
rect 345876 24325 345918 24561
rect 346154 24325 346196 24561
rect 345876 17561 346196 24325
rect 345876 17325 345918 17561
rect 346154 17325 346196 17561
rect 345876 10561 346196 17325
rect 345876 10325 345918 10561
rect 346154 10325 346196 10561
rect 345876 3561 346196 10325
rect 345876 3325 345918 3561
rect 346154 3325 346196 3561
rect 345876 -1706 346196 3325
rect 345876 -1942 345918 -1706
rect 346154 -1942 346196 -1706
rect 345876 -2026 346196 -1942
rect 345876 -2262 345918 -2026
rect 346154 -2262 346196 -2026
rect 345876 -2294 346196 -2262
rect 351144 705238 351464 706230
rect 351144 705002 351186 705238
rect 351422 705002 351464 705238
rect 351144 704918 351464 705002
rect 351144 704682 351186 704918
rect 351422 704682 351464 704918
rect 351144 695494 351464 704682
rect 351144 695258 351186 695494
rect 351422 695258 351464 695494
rect 351144 688494 351464 695258
rect 351144 688258 351186 688494
rect 351422 688258 351464 688494
rect 351144 681494 351464 688258
rect 351144 681258 351186 681494
rect 351422 681258 351464 681494
rect 351144 674494 351464 681258
rect 351144 674258 351186 674494
rect 351422 674258 351464 674494
rect 351144 667494 351464 674258
rect 351144 667258 351186 667494
rect 351422 667258 351464 667494
rect 351144 660494 351464 667258
rect 351144 660258 351186 660494
rect 351422 660258 351464 660494
rect 351144 653494 351464 660258
rect 351144 653258 351186 653494
rect 351422 653258 351464 653494
rect 351144 646494 351464 653258
rect 351144 646258 351186 646494
rect 351422 646258 351464 646494
rect 351144 639494 351464 646258
rect 351144 639258 351186 639494
rect 351422 639258 351464 639494
rect 351144 632494 351464 639258
rect 351144 632258 351186 632494
rect 351422 632258 351464 632494
rect 351144 625494 351464 632258
rect 351144 625258 351186 625494
rect 351422 625258 351464 625494
rect 351144 618494 351464 625258
rect 351144 618258 351186 618494
rect 351422 618258 351464 618494
rect 351144 611494 351464 618258
rect 351144 611258 351186 611494
rect 351422 611258 351464 611494
rect 351144 604494 351464 611258
rect 351144 604258 351186 604494
rect 351422 604258 351464 604494
rect 351144 597494 351464 604258
rect 351144 597258 351186 597494
rect 351422 597258 351464 597494
rect 351144 590494 351464 597258
rect 351144 590258 351186 590494
rect 351422 590258 351464 590494
rect 351144 583494 351464 590258
rect 351144 583258 351186 583494
rect 351422 583258 351464 583494
rect 351144 576494 351464 583258
rect 351144 576258 351186 576494
rect 351422 576258 351464 576494
rect 351144 569494 351464 576258
rect 351144 569258 351186 569494
rect 351422 569258 351464 569494
rect 351144 562494 351464 569258
rect 351144 562258 351186 562494
rect 351422 562258 351464 562494
rect 351144 555494 351464 562258
rect 351144 555258 351186 555494
rect 351422 555258 351464 555494
rect 351144 548494 351464 555258
rect 351144 548258 351186 548494
rect 351422 548258 351464 548494
rect 351144 541494 351464 548258
rect 351144 541258 351186 541494
rect 351422 541258 351464 541494
rect 351144 534494 351464 541258
rect 351144 534258 351186 534494
rect 351422 534258 351464 534494
rect 351144 527494 351464 534258
rect 351144 527258 351186 527494
rect 351422 527258 351464 527494
rect 351144 520494 351464 527258
rect 351144 520258 351186 520494
rect 351422 520258 351464 520494
rect 351144 513494 351464 520258
rect 351144 513258 351186 513494
rect 351422 513258 351464 513494
rect 351144 506494 351464 513258
rect 351144 506258 351186 506494
rect 351422 506258 351464 506494
rect 351144 499494 351464 506258
rect 351144 499258 351186 499494
rect 351422 499258 351464 499494
rect 351144 492494 351464 499258
rect 351144 492258 351186 492494
rect 351422 492258 351464 492494
rect 351144 485494 351464 492258
rect 351144 485258 351186 485494
rect 351422 485258 351464 485494
rect 351144 478494 351464 485258
rect 351144 478258 351186 478494
rect 351422 478258 351464 478494
rect 351144 471494 351464 478258
rect 351144 471258 351186 471494
rect 351422 471258 351464 471494
rect 351144 464494 351464 471258
rect 351144 464258 351186 464494
rect 351422 464258 351464 464494
rect 351144 457494 351464 464258
rect 351144 457258 351186 457494
rect 351422 457258 351464 457494
rect 351144 450494 351464 457258
rect 351144 450258 351186 450494
rect 351422 450258 351464 450494
rect 351144 443494 351464 450258
rect 351144 443258 351186 443494
rect 351422 443258 351464 443494
rect 351144 436494 351464 443258
rect 351144 436258 351186 436494
rect 351422 436258 351464 436494
rect 351144 429494 351464 436258
rect 351144 429258 351186 429494
rect 351422 429258 351464 429494
rect 351144 422494 351464 429258
rect 351144 422258 351186 422494
rect 351422 422258 351464 422494
rect 351144 415494 351464 422258
rect 351144 415258 351186 415494
rect 351422 415258 351464 415494
rect 351144 408494 351464 415258
rect 351144 408258 351186 408494
rect 351422 408258 351464 408494
rect 351144 401494 351464 408258
rect 351144 401258 351186 401494
rect 351422 401258 351464 401494
rect 351144 394494 351464 401258
rect 351144 394258 351186 394494
rect 351422 394258 351464 394494
rect 351144 387494 351464 394258
rect 351144 387258 351186 387494
rect 351422 387258 351464 387494
rect 351144 380494 351464 387258
rect 351144 380258 351186 380494
rect 351422 380258 351464 380494
rect 351144 373494 351464 380258
rect 351144 373258 351186 373494
rect 351422 373258 351464 373494
rect 351144 366494 351464 373258
rect 351144 366258 351186 366494
rect 351422 366258 351464 366494
rect 351144 359494 351464 366258
rect 351144 359258 351186 359494
rect 351422 359258 351464 359494
rect 351144 352494 351464 359258
rect 351144 352258 351186 352494
rect 351422 352258 351464 352494
rect 351144 345494 351464 352258
rect 351144 345258 351186 345494
rect 351422 345258 351464 345494
rect 351144 338494 351464 345258
rect 351144 338258 351186 338494
rect 351422 338258 351464 338494
rect 351144 331494 351464 338258
rect 351144 331258 351186 331494
rect 351422 331258 351464 331494
rect 351144 324494 351464 331258
rect 351144 324258 351186 324494
rect 351422 324258 351464 324494
rect 351144 317494 351464 324258
rect 351144 317258 351186 317494
rect 351422 317258 351464 317494
rect 351144 310494 351464 317258
rect 351144 310258 351186 310494
rect 351422 310258 351464 310494
rect 351144 303494 351464 310258
rect 351144 303258 351186 303494
rect 351422 303258 351464 303494
rect 351144 296494 351464 303258
rect 351144 296258 351186 296494
rect 351422 296258 351464 296494
rect 351144 289494 351464 296258
rect 351144 289258 351186 289494
rect 351422 289258 351464 289494
rect 351144 282494 351464 289258
rect 351144 282258 351186 282494
rect 351422 282258 351464 282494
rect 351144 275494 351464 282258
rect 351144 275258 351186 275494
rect 351422 275258 351464 275494
rect 351144 268494 351464 275258
rect 351144 268258 351186 268494
rect 351422 268258 351464 268494
rect 351144 261494 351464 268258
rect 351144 261258 351186 261494
rect 351422 261258 351464 261494
rect 351144 254494 351464 261258
rect 351144 254258 351186 254494
rect 351422 254258 351464 254494
rect 351144 247494 351464 254258
rect 351144 247258 351186 247494
rect 351422 247258 351464 247494
rect 351144 240494 351464 247258
rect 351144 240258 351186 240494
rect 351422 240258 351464 240494
rect 351144 233494 351464 240258
rect 351144 233258 351186 233494
rect 351422 233258 351464 233494
rect 351144 226494 351464 233258
rect 351144 226258 351186 226494
rect 351422 226258 351464 226494
rect 351144 219494 351464 226258
rect 351144 219258 351186 219494
rect 351422 219258 351464 219494
rect 351144 212494 351464 219258
rect 351144 212258 351186 212494
rect 351422 212258 351464 212494
rect 351144 205494 351464 212258
rect 351144 205258 351186 205494
rect 351422 205258 351464 205494
rect 351144 198494 351464 205258
rect 351144 198258 351186 198494
rect 351422 198258 351464 198494
rect 351144 191494 351464 198258
rect 351144 191258 351186 191494
rect 351422 191258 351464 191494
rect 351144 184494 351464 191258
rect 351144 184258 351186 184494
rect 351422 184258 351464 184494
rect 351144 177494 351464 184258
rect 351144 177258 351186 177494
rect 351422 177258 351464 177494
rect 351144 170494 351464 177258
rect 351144 170258 351186 170494
rect 351422 170258 351464 170494
rect 351144 163494 351464 170258
rect 351144 163258 351186 163494
rect 351422 163258 351464 163494
rect 351144 156494 351464 163258
rect 351144 156258 351186 156494
rect 351422 156258 351464 156494
rect 351144 149494 351464 156258
rect 351144 149258 351186 149494
rect 351422 149258 351464 149494
rect 351144 142494 351464 149258
rect 351144 142258 351186 142494
rect 351422 142258 351464 142494
rect 351144 135494 351464 142258
rect 351144 135258 351186 135494
rect 351422 135258 351464 135494
rect 351144 128494 351464 135258
rect 351144 128258 351186 128494
rect 351422 128258 351464 128494
rect 351144 121494 351464 128258
rect 351144 121258 351186 121494
rect 351422 121258 351464 121494
rect 351144 114494 351464 121258
rect 351144 114258 351186 114494
rect 351422 114258 351464 114494
rect 351144 107494 351464 114258
rect 351144 107258 351186 107494
rect 351422 107258 351464 107494
rect 351144 100494 351464 107258
rect 351144 100258 351186 100494
rect 351422 100258 351464 100494
rect 351144 93494 351464 100258
rect 351144 93258 351186 93494
rect 351422 93258 351464 93494
rect 351144 86494 351464 93258
rect 351144 86258 351186 86494
rect 351422 86258 351464 86494
rect 351144 79494 351464 86258
rect 351144 79258 351186 79494
rect 351422 79258 351464 79494
rect 351144 72494 351464 79258
rect 351144 72258 351186 72494
rect 351422 72258 351464 72494
rect 351144 65494 351464 72258
rect 351144 65258 351186 65494
rect 351422 65258 351464 65494
rect 351144 58494 351464 65258
rect 351144 58258 351186 58494
rect 351422 58258 351464 58494
rect 351144 51494 351464 58258
rect 351144 51258 351186 51494
rect 351422 51258 351464 51494
rect 351144 44494 351464 51258
rect 351144 44258 351186 44494
rect 351422 44258 351464 44494
rect 351144 37494 351464 44258
rect 351144 37258 351186 37494
rect 351422 37258 351464 37494
rect 351144 30494 351464 37258
rect 351144 30258 351186 30494
rect 351422 30258 351464 30494
rect 351144 23494 351464 30258
rect 351144 23258 351186 23494
rect 351422 23258 351464 23494
rect 351144 16494 351464 23258
rect 351144 16258 351186 16494
rect 351422 16258 351464 16494
rect 351144 9494 351464 16258
rect 351144 9258 351186 9494
rect 351422 9258 351464 9494
rect 351144 2494 351464 9258
rect 351144 2258 351186 2494
rect 351422 2258 351464 2494
rect 351144 -746 351464 2258
rect 351144 -982 351186 -746
rect 351422 -982 351464 -746
rect 351144 -1066 351464 -982
rect 351144 -1302 351186 -1066
rect 351422 -1302 351464 -1066
rect 351144 -2294 351464 -1302
rect 352876 706198 353196 706230
rect 352876 705962 352918 706198
rect 353154 705962 353196 706198
rect 352876 705878 353196 705962
rect 352876 705642 352918 705878
rect 353154 705642 353196 705878
rect 352876 696561 353196 705642
rect 352876 696325 352918 696561
rect 353154 696325 353196 696561
rect 352876 689561 353196 696325
rect 352876 689325 352918 689561
rect 353154 689325 353196 689561
rect 352876 682561 353196 689325
rect 352876 682325 352918 682561
rect 353154 682325 353196 682561
rect 352876 675561 353196 682325
rect 352876 675325 352918 675561
rect 353154 675325 353196 675561
rect 352876 668561 353196 675325
rect 352876 668325 352918 668561
rect 353154 668325 353196 668561
rect 352876 661561 353196 668325
rect 352876 661325 352918 661561
rect 353154 661325 353196 661561
rect 352876 654561 353196 661325
rect 352876 654325 352918 654561
rect 353154 654325 353196 654561
rect 352876 647561 353196 654325
rect 352876 647325 352918 647561
rect 353154 647325 353196 647561
rect 352876 640561 353196 647325
rect 352876 640325 352918 640561
rect 353154 640325 353196 640561
rect 352876 633561 353196 640325
rect 352876 633325 352918 633561
rect 353154 633325 353196 633561
rect 352876 626561 353196 633325
rect 352876 626325 352918 626561
rect 353154 626325 353196 626561
rect 352876 619561 353196 626325
rect 352876 619325 352918 619561
rect 353154 619325 353196 619561
rect 352876 612561 353196 619325
rect 352876 612325 352918 612561
rect 353154 612325 353196 612561
rect 352876 605561 353196 612325
rect 352876 605325 352918 605561
rect 353154 605325 353196 605561
rect 352876 598561 353196 605325
rect 352876 598325 352918 598561
rect 353154 598325 353196 598561
rect 352876 591561 353196 598325
rect 352876 591325 352918 591561
rect 353154 591325 353196 591561
rect 352876 584561 353196 591325
rect 352876 584325 352918 584561
rect 353154 584325 353196 584561
rect 352876 577561 353196 584325
rect 352876 577325 352918 577561
rect 353154 577325 353196 577561
rect 352876 570561 353196 577325
rect 352876 570325 352918 570561
rect 353154 570325 353196 570561
rect 352876 563561 353196 570325
rect 352876 563325 352918 563561
rect 353154 563325 353196 563561
rect 352876 556561 353196 563325
rect 352876 556325 352918 556561
rect 353154 556325 353196 556561
rect 352876 549561 353196 556325
rect 352876 549325 352918 549561
rect 353154 549325 353196 549561
rect 352876 542561 353196 549325
rect 352876 542325 352918 542561
rect 353154 542325 353196 542561
rect 352876 535561 353196 542325
rect 352876 535325 352918 535561
rect 353154 535325 353196 535561
rect 352876 528561 353196 535325
rect 352876 528325 352918 528561
rect 353154 528325 353196 528561
rect 352876 521561 353196 528325
rect 352876 521325 352918 521561
rect 353154 521325 353196 521561
rect 352876 514561 353196 521325
rect 352876 514325 352918 514561
rect 353154 514325 353196 514561
rect 352876 507561 353196 514325
rect 352876 507325 352918 507561
rect 353154 507325 353196 507561
rect 352876 500561 353196 507325
rect 352876 500325 352918 500561
rect 353154 500325 353196 500561
rect 352876 493561 353196 500325
rect 352876 493325 352918 493561
rect 353154 493325 353196 493561
rect 352876 486561 353196 493325
rect 352876 486325 352918 486561
rect 353154 486325 353196 486561
rect 352876 479561 353196 486325
rect 352876 479325 352918 479561
rect 353154 479325 353196 479561
rect 352876 472561 353196 479325
rect 352876 472325 352918 472561
rect 353154 472325 353196 472561
rect 352876 465561 353196 472325
rect 352876 465325 352918 465561
rect 353154 465325 353196 465561
rect 352876 458561 353196 465325
rect 352876 458325 352918 458561
rect 353154 458325 353196 458561
rect 352876 451561 353196 458325
rect 352876 451325 352918 451561
rect 353154 451325 353196 451561
rect 352876 444561 353196 451325
rect 352876 444325 352918 444561
rect 353154 444325 353196 444561
rect 352876 437561 353196 444325
rect 352876 437325 352918 437561
rect 353154 437325 353196 437561
rect 352876 430561 353196 437325
rect 352876 430325 352918 430561
rect 353154 430325 353196 430561
rect 352876 423561 353196 430325
rect 352876 423325 352918 423561
rect 353154 423325 353196 423561
rect 352876 416561 353196 423325
rect 352876 416325 352918 416561
rect 353154 416325 353196 416561
rect 352876 409561 353196 416325
rect 352876 409325 352918 409561
rect 353154 409325 353196 409561
rect 352876 402561 353196 409325
rect 352876 402325 352918 402561
rect 353154 402325 353196 402561
rect 352876 395561 353196 402325
rect 352876 395325 352918 395561
rect 353154 395325 353196 395561
rect 352876 388561 353196 395325
rect 352876 388325 352918 388561
rect 353154 388325 353196 388561
rect 352876 381561 353196 388325
rect 352876 381325 352918 381561
rect 353154 381325 353196 381561
rect 352876 374561 353196 381325
rect 352876 374325 352918 374561
rect 353154 374325 353196 374561
rect 352876 367561 353196 374325
rect 352876 367325 352918 367561
rect 353154 367325 353196 367561
rect 352876 360561 353196 367325
rect 352876 360325 352918 360561
rect 353154 360325 353196 360561
rect 352876 353561 353196 360325
rect 352876 353325 352918 353561
rect 353154 353325 353196 353561
rect 352876 346561 353196 353325
rect 352876 346325 352918 346561
rect 353154 346325 353196 346561
rect 352876 339561 353196 346325
rect 352876 339325 352918 339561
rect 353154 339325 353196 339561
rect 352876 332561 353196 339325
rect 352876 332325 352918 332561
rect 353154 332325 353196 332561
rect 352876 325561 353196 332325
rect 352876 325325 352918 325561
rect 353154 325325 353196 325561
rect 352876 318561 353196 325325
rect 352876 318325 352918 318561
rect 353154 318325 353196 318561
rect 352876 311561 353196 318325
rect 352876 311325 352918 311561
rect 353154 311325 353196 311561
rect 352876 304561 353196 311325
rect 352876 304325 352918 304561
rect 353154 304325 353196 304561
rect 352876 297561 353196 304325
rect 352876 297325 352918 297561
rect 353154 297325 353196 297561
rect 352876 290561 353196 297325
rect 352876 290325 352918 290561
rect 353154 290325 353196 290561
rect 352876 283561 353196 290325
rect 352876 283325 352918 283561
rect 353154 283325 353196 283561
rect 352876 276561 353196 283325
rect 352876 276325 352918 276561
rect 353154 276325 353196 276561
rect 352876 269561 353196 276325
rect 352876 269325 352918 269561
rect 353154 269325 353196 269561
rect 352876 262561 353196 269325
rect 352876 262325 352918 262561
rect 353154 262325 353196 262561
rect 352876 255561 353196 262325
rect 352876 255325 352918 255561
rect 353154 255325 353196 255561
rect 352876 248561 353196 255325
rect 352876 248325 352918 248561
rect 353154 248325 353196 248561
rect 352876 241561 353196 248325
rect 352876 241325 352918 241561
rect 353154 241325 353196 241561
rect 352876 234561 353196 241325
rect 352876 234325 352918 234561
rect 353154 234325 353196 234561
rect 352876 227561 353196 234325
rect 352876 227325 352918 227561
rect 353154 227325 353196 227561
rect 352876 220561 353196 227325
rect 352876 220325 352918 220561
rect 353154 220325 353196 220561
rect 352876 213561 353196 220325
rect 352876 213325 352918 213561
rect 353154 213325 353196 213561
rect 352876 206561 353196 213325
rect 352876 206325 352918 206561
rect 353154 206325 353196 206561
rect 352876 199561 353196 206325
rect 352876 199325 352918 199561
rect 353154 199325 353196 199561
rect 352876 192561 353196 199325
rect 352876 192325 352918 192561
rect 353154 192325 353196 192561
rect 352876 185561 353196 192325
rect 352876 185325 352918 185561
rect 353154 185325 353196 185561
rect 352876 178561 353196 185325
rect 352876 178325 352918 178561
rect 353154 178325 353196 178561
rect 352876 171561 353196 178325
rect 352876 171325 352918 171561
rect 353154 171325 353196 171561
rect 352876 164561 353196 171325
rect 352876 164325 352918 164561
rect 353154 164325 353196 164561
rect 352876 157561 353196 164325
rect 352876 157325 352918 157561
rect 353154 157325 353196 157561
rect 352876 150561 353196 157325
rect 352876 150325 352918 150561
rect 353154 150325 353196 150561
rect 352876 143561 353196 150325
rect 352876 143325 352918 143561
rect 353154 143325 353196 143561
rect 352876 136561 353196 143325
rect 352876 136325 352918 136561
rect 353154 136325 353196 136561
rect 352876 129561 353196 136325
rect 352876 129325 352918 129561
rect 353154 129325 353196 129561
rect 352876 122561 353196 129325
rect 352876 122325 352918 122561
rect 353154 122325 353196 122561
rect 352876 115561 353196 122325
rect 352876 115325 352918 115561
rect 353154 115325 353196 115561
rect 352876 108561 353196 115325
rect 352876 108325 352918 108561
rect 353154 108325 353196 108561
rect 352876 101561 353196 108325
rect 352876 101325 352918 101561
rect 353154 101325 353196 101561
rect 352876 94561 353196 101325
rect 352876 94325 352918 94561
rect 353154 94325 353196 94561
rect 352876 87561 353196 94325
rect 352876 87325 352918 87561
rect 353154 87325 353196 87561
rect 352876 80561 353196 87325
rect 352876 80325 352918 80561
rect 353154 80325 353196 80561
rect 352876 73561 353196 80325
rect 352876 73325 352918 73561
rect 353154 73325 353196 73561
rect 352876 66561 353196 73325
rect 352876 66325 352918 66561
rect 353154 66325 353196 66561
rect 352876 59561 353196 66325
rect 352876 59325 352918 59561
rect 353154 59325 353196 59561
rect 352876 52561 353196 59325
rect 352876 52325 352918 52561
rect 353154 52325 353196 52561
rect 352876 45561 353196 52325
rect 352876 45325 352918 45561
rect 353154 45325 353196 45561
rect 352876 38561 353196 45325
rect 352876 38325 352918 38561
rect 353154 38325 353196 38561
rect 352876 31561 353196 38325
rect 352876 31325 352918 31561
rect 353154 31325 353196 31561
rect 352876 24561 353196 31325
rect 352876 24325 352918 24561
rect 353154 24325 353196 24561
rect 352876 17561 353196 24325
rect 352876 17325 352918 17561
rect 353154 17325 353196 17561
rect 352876 10561 353196 17325
rect 352876 10325 352918 10561
rect 353154 10325 353196 10561
rect 352876 3561 353196 10325
rect 352876 3325 352918 3561
rect 353154 3325 353196 3561
rect 352876 -1706 353196 3325
rect 352876 -1942 352918 -1706
rect 353154 -1942 353196 -1706
rect 352876 -2026 353196 -1942
rect 352876 -2262 352918 -2026
rect 353154 -2262 353196 -2026
rect 352876 -2294 353196 -2262
rect 358144 705238 358464 706230
rect 358144 705002 358186 705238
rect 358422 705002 358464 705238
rect 358144 704918 358464 705002
rect 358144 704682 358186 704918
rect 358422 704682 358464 704918
rect 358144 695494 358464 704682
rect 358144 695258 358186 695494
rect 358422 695258 358464 695494
rect 358144 688494 358464 695258
rect 358144 688258 358186 688494
rect 358422 688258 358464 688494
rect 358144 681494 358464 688258
rect 358144 681258 358186 681494
rect 358422 681258 358464 681494
rect 358144 674494 358464 681258
rect 358144 674258 358186 674494
rect 358422 674258 358464 674494
rect 358144 667494 358464 674258
rect 358144 667258 358186 667494
rect 358422 667258 358464 667494
rect 358144 660494 358464 667258
rect 358144 660258 358186 660494
rect 358422 660258 358464 660494
rect 358144 653494 358464 660258
rect 358144 653258 358186 653494
rect 358422 653258 358464 653494
rect 358144 646494 358464 653258
rect 358144 646258 358186 646494
rect 358422 646258 358464 646494
rect 358144 639494 358464 646258
rect 358144 639258 358186 639494
rect 358422 639258 358464 639494
rect 358144 632494 358464 639258
rect 358144 632258 358186 632494
rect 358422 632258 358464 632494
rect 358144 625494 358464 632258
rect 358144 625258 358186 625494
rect 358422 625258 358464 625494
rect 358144 618494 358464 625258
rect 358144 618258 358186 618494
rect 358422 618258 358464 618494
rect 358144 611494 358464 618258
rect 358144 611258 358186 611494
rect 358422 611258 358464 611494
rect 358144 604494 358464 611258
rect 358144 604258 358186 604494
rect 358422 604258 358464 604494
rect 358144 597494 358464 604258
rect 358144 597258 358186 597494
rect 358422 597258 358464 597494
rect 358144 590494 358464 597258
rect 358144 590258 358186 590494
rect 358422 590258 358464 590494
rect 358144 583494 358464 590258
rect 358144 583258 358186 583494
rect 358422 583258 358464 583494
rect 358144 576494 358464 583258
rect 358144 576258 358186 576494
rect 358422 576258 358464 576494
rect 358144 569494 358464 576258
rect 358144 569258 358186 569494
rect 358422 569258 358464 569494
rect 358144 562494 358464 569258
rect 358144 562258 358186 562494
rect 358422 562258 358464 562494
rect 358144 555494 358464 562258
rect 358144 555258 358186 555494
rect 358422 555258 358464 555494
rect 358144 548494 358464 555258
rect 358144 548258 358186 548494
rect 358422 548258 358464 548494
rect 358144 541494 358464 548258
rect 358144 541258 358186 541494
rect 358422 541258 358464 541494
rect 358144 534494 358464 541258
rect 358144 534258 358186 534494
rect 358422 534258 358464 534494
rect 358144 527494 358464 534258
rect 358144 527258 358186 527494
rect 358422 527258 358464 527494
rect 358144 520494 358464 527258
rect 358144 520258 358186 520494
rect 358422 520258 358464 520494
rect 358144 513494 358464 520258
rect 358144 513258 358186 513494
rect 358422 513258 358464 513494
rect 358144 506494 358464 513258
rect 358144 506258 358186 506494
rect 358422 506258 358464 506494
rect 358144 499494 358464 506258
rect 358144 499258 358186 499494
rect 358422 499258 358464 499494
rect 358144 492494 358464 499258
rect 358144 492258 358186 492494
rect 358422 492258 358464 492494
rect 358144 485494 358464 492258
rect 358144 485258 358186 485494
rect 358422 485258 358464 485494
rect 358144 478494 358464 485258
rect 358144 478258 358186 478494
rect 358422 478258 358464 478494
rect 358144 471494 358464 478258
rect 358144 471258 358186 471494
rect 358422 471258 358464 471494
rect 358144 464494 358464 471258
rect 358144 464258 358186 464494
rect 358422 464258 358464 464494
rect 358144 457494 358464 464258
rect 358144 457258 358186 457494
rect 358422 457258 358464 457494
rect 358144 450494 358464 457258
rect 358144 450258 358186 450494
rect 358422 450258 358464 450494
rect 358144 443494 358464 450258
rect 358144 443258 358186 443494
rect 358422 443258 358464 443494
rect 358144 436494 358464 443258
rect 358144 436258 358186 436494
rect 358422 436258 358464 436494
rect 358144 429494 358464 436258
rect 358144 429258 358186 429494
rect 358422 429258 358464 429494
rect 358144 422494 358464 429258
rect 358144 422258 358186 422494
rect 358422 422258 358464 422494
rect 358144 415494 358464 422258
rect 358144 415258 358186 415494
rect 358422 415258 358464 415494
rect 358144 408494 358464 415258
rect 358144 408258 358186 408494
rect 358422 408258 358464 408494
rect 358144 401494 358464 408258
rect 358144 401258 358186 401494
rect 358422 401258 358464 401494
rect 358144 394494 358464 401258
rect 358144 394258 358186 394494
rect 358422 394258 358464 394494
rect 358144 387494 358464 394258
rect 358144 387258 358186 387494
rect 358422 387258 358464 387494
rect 358144 380494 358464 387258
rect 358144 380258 358186 380494
rect 358422 380258 358464 380494
rect 358144 373494 358464 380258
rect 358144 373258 358186 373494
rect 358422 373258 358464 373494
rect 358144 366494 358464 373258
rect 358144 366258 358186 366494
rect 358422 366258 358464 366494
rect 358144 359494 358464 366258
rect 358144 359258 358186 359494
rect 358422 359258 358464 359494
rect 358144 352494 358464 359258
rect 358144 352258 358186 352494
rect 358422 352258 358464 352494
rect 358144 345494 358464 352258
rect 358144 345258 358186 345494
rect 358422 345258 358464 345494
rect 358144 338494 358464 345258
rect 358144 338258 358186 338494
rect 358422 338258 358464 338494
rect 358144 331494 358464 338258
rect 358144 331258 358186 331494
rect 358422 331258 358464 331494
rect 358144 324494 358464 331258
rect 358144 324258 358186 324494
rect 358422 324258 358464 324494
rect 358144 317494 358464 324258
rect 358144 317258 358186 317494
rect 358422 317258 358464 317494
rect 358144 310494 358464 317258
rect 358144 310258 358186 310494
rect 358422 310258 358464 310494
rect 358144 303494 358464 310258
rect 358144 303258 358186 303494
rect 358422 303258 358464 303494
rect 358144 296494 358464 303258
rect 358144 296258 358186 296494
rect 358422 296258 358464 296494
rect 358144 289494 358464 296258
rect 358144 289258 358186 289494
rect 358422 289258 358464 289494
rect 358144 282494 358464 289258
rect 358144 282258 358186 282494
rect 358422 282258 358464 282494
rect 358144 275494 358464 282258
rect 358144 275258 358186 275494
rect 358422 275258 358464 275494
rect 358144 268494 358464 275258
rect 358144 268258 358186 268494
rect 358422 268258 358464 268494
rect 358144 261494 358464 268258
rect 358144 261258 358186 261494
rect 358422 261258 358464 261494
rect 358144 254494 358464 261258
rect 358144 254258 358186 254494
rect 358422 254258 358464 254494
rect 358144 247494 358464 254258
rect 358144 247258 358186 247494
rect 358422 247258 358464 247494
rect 358144 240494 358464 247258
rect 358144 240258 358186 240494
rect 358422 240258 358464 240494
rect 358144 233494 358464 240258
rect 358144 233258 358186 233494
rect 358422 233258 358464 233494
rect 358144 226494 358464 233258
rect 358144 226258 358186 226494
rect 358422 226258 358464 226494
rect 358144 219494 358464 226258
rect 358144 219258 358186 219494
rect 358422 219258 358464 219494
rect 358144 212494 358464 219258
rect 358144 212258 358186 212494
rect 358422 212258 358464 212494
rect 358144 205494 358464 212258
rect 358144 205258 358186 205494
rect 358422 205258 358464 205494
rect 358144 198494 358464 205258
rect 358144 198258 358186 198494
rect 358422 198258 358464 198494
rect 358144 191494 358464 198258
rect 358144 191258 358186 191494
rect 358422 191258 358464 191494
rect 358144 184494 358464 191258
rect 358144 184258 358186 184494
rect 358422 184258 358464 184494
rect 358144 177494 358464 184258
rect 358144 177258 358186 177494
rect 358422 177258 358464 177494
rect 358144 170494 358464 177258
rect 358144 170258 358186 170494
rect 358422 170258 358464 170494
rect 358144 163494 358464 170258
rect 358144 163258 358186 163494
rect 358422 163258 358464 163494
rect 358144 156494 358464 163258
rect 358144 156258 358186 156494
rect 358422 156258 358464 156494
rect 358144 149494 358464 156258
rect 358144 149258 358186 149494
rect 358422 149258 358464 149494
rect 358144 142494 358464 149258
rect 358144 142258 358186 142494
rect 358422 142258 358464 142494
rect 358144 135494 358464 142258
rect 358144 135258 358186 135494
rect 358422 135258 358464 135494
rect 358144 128494 358464 135258
rect 358144 128258 358186 128494
rect 358422 128258 358464 128494
rect 358144 121494 358464 128258
rect 358144 121258 358186 121494
rect 358422 121258 358464 121494
rect 358144 114494 358464 121258
rect 358144 114258 358186 114494
rect 358422 114258 358464 114494
rect 358144 107494 358464 114258
rect 358144 107258 358186 107494
rect 358422 107258 358464 107494
rect 358144 100494 358464 107258
rect 358144 100258 358186 100494
rect 358422 100258 358464 100494
rect 358144 93494 358464 100258
rect 358144 93258 358186 93494
rect 358422 93258 358464 93494
rect 358144 86494 358464 93258
rect 358144 86258 358186 86494
rect 358422 86258 358464 86494
rect 358144 79494 358464 86258
rect 358144 79258 358186 79494
rect 358422 79258 358464 79494
rect 358144 72494 358464 79258
rect 358144 72258 358186 72494
rect 358422 72258 358464 72494
rect 358144 65494 358464 72258
rect 358144 65258 358186 65494
rect 358422 65258 358464 65494
rect 358144 58494 358464 65258
rect 358144 58258 358186 58494
rect 358422 58258 358464 58494
rect 358144 51494 358464 58258
rect 358144 51258 358186 51494
rect 358422 51258 358464 51494
rect 358144 44494 358464 51258
rect 358144 44258 358186 44494
rect 358422 44258 358464 44494
rect 358144 37494 358464 44258
rect 358144 37258 358186 37494
rect 358422 37258 358464 37494
rect 358144 30494 358464 37258
rect 358144 30258 358186 30494
rect 358422 30258 358464 30494
rect 358144 23494 358464 30258
rect 358144 23258 358186 23494
rect 358422 23258 358464 23494
rect 358144 16494 358464 23258
rect 358144 16258 358186 16494
rect 358422 16258 358464 16494
rect 358144 9494 358464 16258
rect 358144 9258 358186 9494
rect 358422 9258 358464 9494
rect 358144 2494 358464 9258
rect 358144 2258 358186 2494
rect 358422 2258 358464 2494
rect 358144 -746 358464 2258
rect 358144 -982 358186 -746
rect 358422 -982 358464 -746
rect 358144 -1066 358464 -982
rect 358144 -1302 358186 -1066
rect 358422 -1302 358464 -1066
rect 358144 -2294 358464 -1302
rect 359876 706198 360196 706230
rect 359876 705962 359918 706198
rect 360154 705962 360196 706198
rect 359876 705878 360196 705962
rect 359876 705642 359918 705878
rect 360154 705642 360196 705878
rect 359876 696561 360196 705642
rect 359876 696325 359918 696561
rect 360154 696325 360196 696561
rect 359876 689561 360196 696325
rect 359876 689325 359918 689561
rect 360154 689325 360196 689561
rect 359876 682561 360196 689325
rect 359876 682325 359918 682561
rect 360154 682325 360196 682561
rect 359876 675561 360196 682325
rect 359876 675325 359918 675561
rect 360154 675325 360196 675561
rect 359876 668561 360196 675325
rect 359876 668325 359918 668561
rect 360154 668325 360196 668561
rect 359876 661561 360196 668325
rect 359876 661325 359918 661561
rect 360154 661325 360196 661561
rect 359876 654561 360196 661325
rect 359876 654325 359918 654561
rect 360154 654325 360196 654561
rect 359876 647561 360196 654325
rect 359876 647325 359918 647561
rect 360154 647325 360196 647561
rect 359876 640561 360196 647325
rect 359876 640325 359918 640561
rect 360154 640325 360196 640561
rect 359876 633561 360196 640325
rect 359876 633325 359918 633561
rect 360154 633325 360196 633561
rect 359876 626561 360196 633325
rect 359876 626325 359918 626561
rect 360154 626325 360196 626561
rect 359876 619561 360196 626325
rect 359876 619325 359918 619561
rect 360154 619325 360196 619561
rect 359876 612561 360196 619325
rect 359876 612325 359918 612561
rect 360154 612325 360196 612561
rect 359876 605561 360196 612325
rect 359876 605325 359918 605561
rect 360154 605325 360196 605561
rect 359876 598561 360196 605325
rect 359876 598325 359918 598561
rect 360154 598325 360196 598561
rect 359876 591561 360196 598325
rect 359876 591325 359918 591561
rect 360154 591325 360196 591561
rect 359876 584561 360196 591325
rect 359876 584325 359918 584561
rect 360154 584325 360196 584561
rect 359876 577561 360196 584325
rect 359876 577325 359918 577561
rect 360154 577325 360196 577561
rect 359876 570561 360196 577325
rect 359876 570325 359918 570561
rect 360154 570325 360196 570561
rect 359876 563561 360196 570325
rect 359876 563325 359918 563561
rect 360154 563325 360196 563561
rect 359876 556561 360196 563325
rect 359876 556325 359918 556561
rect 360154 556325 360196 556561
rect 359876 549561 360196 556325
rect 359876 549325 359918 549561
rect 360154 549325 360196 549561
rect 359876 542561 360196 549325
rect 359876 542325 359918 542561
rect 360154 542325 360196 542561
rect 359876 535561 360196 542325
rect 359876 535325 359918 535561
rect 360154 535325 360196 535561
rect 359876 528561 360196 535325
rect 359876 528325 359918 528561
rect 360154 528325 360196 528561
rect 359876 521561 360196 528325
rect 359876 521325 359918 521561
rect 360154 521325 360196 521561
rect 359876 514561 360196 521325
rect 359876 514325 359918 514561
rect 360154 514325 360196 514561
rect 359876 507561 360196 514325
rect 359876 507325 359918 507561
rect 360154 507325 360196 507561
rect 359876 500561 360196 507325
rect 359876 500325 359918 500561
rect 360154 500325 360196 500561
rect 359876 493561 360196 500325
rect 359876 493325 359918 493561
rect 360154 493325 360196 493561
rect 359876 486561 360196 493325
rect 359876 486325 359918 486561
rect 360154 486325 360196 486561
rect 359876 479561 360196 486325
rect 359876 479325 359918 479561
rect 360154 479325 360196 479561
rect 359876 472561 360196 479325
rect 359876 472325 359918 472561
rect 360154 472325 360196 472561
rect 359876 465561 360196 472325
rect 359876 465325 359918 465561
rect 360154 465325 360196 465561
rect 359876 458561 360196 465325
rect 359876 458325 359918 458561
rect 360154 458325 360196 458561
rect 359876 451561 360196 458325
rect 359876 451325 359918 451561
rect 360154 451325 360196 451561
rect 359876 444561 360196 451325
rect 359876 444325 359918 444561
rect 360154 444325 360196 444561
rect 359876 437561 360196 444325
rect 359876 437325 359918 437561
rect 360154 437325 360196 437561
rect 359876 430561 360196 437325
rect 359876 430325 359918 430561
rect 360154 430325 360196 430561
rect 359876 423561 360196 430325
rect 359876 423325 359918 423561
rect 360154 423325 360196 423561
rect 359876 416561 360196 423325
rect 359876 416325 359918 416561
rect 360154 416325 360196 416561
rect 359876 409561 360196 416325
rect 359876 409325 359918 409561
rect 360154 409325 360196 409561
rect 359876 402561 360196 409325
rect 359876 402325 359918 402561
rect 360154 402325 360196 402561
rect 359876 395561 360196 402325
rect 359876 395325 359918 395561
rect 360154 395325 360196 395561
rect 359876 388561 360196 395325
rect 359876 388325 359918 388561
rect 360154 388325 360196 388561
rect 359876 381561 360196 388325
rect 359876 381325 359918 381561
rect 360154 381325 360196 381561
rect 359876 374561 360196 381325
rect 359876 374325 359918 374561
rect 360154 374325 360196 374561
rect 359876 367561 360196 374325
rect 359876 367325 359918 367561
rect 360154 367325 360196 367561
rect 359876 360561 360196 367325
rect 359876 360325 359918 360561
rect 360154 360325 360196 360561
rect 359876 353561 360196 360325
rect 359876 353325 359918 353561
rect 360154 353325 360196 353561
rect 359876 346561 360196 353325
rect 359876 346325 359918 346561
rect 360154 346325 360196 346561
rect 359876 339561 360196 346325
rect 359876 339325 359918 339561
rect 360154 339325 360196 339561
rect 359876 332561 360196 339325
rect 359876 332325 359918 332561
rect 360154 332325 360196 332561
rect 359876 325561 360196 332325
rect 359876 325325 359918 325561
rect 360154 325325 360196 325561
rect 359876 318561 360196 325325
rect 359876 318325 359918 318561
rect 360154 318325 360196 318561
rect 359876 311561 360196 318325
rect 359876 311325 359918 311561
rect 360154 311325 360196 311561
rect 359876 304561 360196 311325
rect 359876 304325 359918 304561
rect 360154 304325 360196 304561
rect 359876 297561 360196 304325
rect 359876 297325 359918 297561
rect 360154 297325 360196 297561
rect 359876 290561 360196 297325
rect 359876 290325 359918 290561
rect 360154 290325 360196 290561
rect 359876 283561 360196 290325
rect 359876 283325 359918 283561
rect 360154 283325 360196 283561
rect 359876 276561 360196 283325
rect 359876 276325 359918 276561
rect 360154 276325 360196 276561
rect 359876 269561 360196 276325
rect 359876 269325 359918 269561
rect 360154 269325 360196 269561
rect 359876 262561 360196 269325
rect 359876 262325 359918 262561
rect 360154 262325 360196 262561
rect 359876 255561 360196 262325
rect 359876 255325 359918 255561
rect 360154 255325 360196 255561
rect 359876 248561 360196 255325
rect 359876 248325 359918 248561
rect 360154 248325 360196 248561
rect 359876 241561 360196 248325
rect 359876 241325 359918 241561
rect 360154 241325 360196 241561
rect 359876 234561 360196 241325
rect 359876 234325 359918 234561
rect 360154 234325 360196 234561
rect 359876 227561 360196 234325
rect 359876 227325 359918 227561
rect 360154 227325 360196 227561
rect 359876 220561 360196 227325
rect 359876 220325 359918 220561
rect 360154 220325 360196 220561
rect 359876 213561 360196 220325
rect 359876 213325 359918 213561
rect 360154 213325 360196 213561
rect 359876 206561 360196 213325
rect 359876 206325 359918 206561
rect 360154 206325 360196 206561
rect 359876 199561 360196 206325
rect 359876 199325 359918 199561
rect 360154 199325 360196 199561
rect 359876 192561 360196 199325
rect 359876 192325 359918 192561
rect 360154 192325 360196 192561
rect 359876 185561 360196 192325
rect 359876 185325 359918 185561
rect 360154 185325 360196 185561
rect 359876 178561 360196 185325
rect 359876 178325 359918 178561
rect 360154 178325 360196 178561
rect 359876 171561 360196 178325
rect 359876 171325 359918 171561
rect 360154 171325 360196 171561
rect 359876 164561 360196 171325
rect 359876 164325 359918 164561
rect 360154 164325 360196 164561
rect 359876 157561 360196 164325
rect 359876 157325 359918 157561
rect 360154 157325 360196 157561
rect 359876 150561 360196 157325
rect 359876 150325 359918 150561
rect 360154 150325 360196 150561
rect 359876 143561 360196 150325
rect 359876 143325 359918 143561
rect 360154 143325 360196 143561
rect 359876 136561 360196 143325
rect 359876 136325 359918 136561
rect 360154 136325 360196 136561
rect 359876 129561 360196 136325
rect 359876 129325 359918 129561
rect 360154 129325 360196 129561
rect 359876 122561 360196 129325
rect 359876 122325 359918 122561
rect 360154 122325 360196 122561
rect 359876 115561 360196 122325
rect 359876 115325 359918 115561
rect 360154 115325 360196 115561
rect 359876 108561 360196 115325
rect 359876 108325 359918 108561
rect 360154 108325 360196 108561
rect 359876 101561 360196 108325
rect 359876 101325 359918 101561
rect 360154 101325 360196 101561
rect 359876 94561 360196 101325
rect 359876 94325 359918 94561
rect 360154 94325 360196 94561
rect 359876 87561 360196 94325
rect 359876 87325 359918 87561
rect 360154 87325 360196 87561
rect 359876 80561 360196 87325
rect 359876 80325 359918 80561
rect 360154 80325 360196 80561
rect 359876 73561 360196 80325
rect 359876 73325 359918 73561
rect 360154 73325 360196 73561
rect 359876 66561 360196 73325
rect 359876 66325 359918 66561
rect 360154 66325 360196 66561
rect 359876 59561 360196 66325
rect 359876 59325 359918 59561
rect 360154 59325 360196 59561
rect 359876 52561 360196 59325
rect 359876 52325 359918 52561
rect 360154 52325 360196 52561
rect 359876 45561 360196 52325
rect 359876 45325 359918 45561
rect 360154 45325 360196 45561
rect 359876 38561 360196 45325
rect 359876 38325 359918 38561
rect 360154 38325 360196 38561
rect 359876 31561 360196 38325
rect 359876 31325 359918 31561
rect 360154 31325 360196 31561
rect 359876 24561 360196 31325
rect 359876 24325 359918 24561
rect 360154 24325 360196 24561
rect 359876 17561 360196 24325
rect 359876 17325 359918 17561
rect 360154 17325 360196 17561
rect 359876 10561 360196 17325
rect 359876 10325 359918 10561
rect 360154 10325 360196 10561
rect 359876 3561 360196 10325
rect 359876 3325 359918 3561
rect 360154 3325 360196 3561
rect 359876 -1706 360196 3325
rect 359876 -1942 359918 -1706
rect 360154 -1942 360196 -1706
rect 359876 -2026 360196 -1942
rect 359876 -2262 359918 -2026
rect 360154 -2262 360196 -2026
rect 359876 -2294 360196 -2262
rect 365144 705238 365464 706230
rect 365144 705002 365186 705238
rect 365422 705002 365464 705238
rect 365144 704918 365464 705002
rect 365144 704682 365186 704918
rect 365422 704682 365464 704918
rect 365144 695494 365464 704682
rect 365144 695258 365186 695494
rect 365422 695258 365464 695494
rect 365144 688494 365464 695258
rect 365144 688258 365186 688494
rect 365422 688258 365464 688494
rect 365144 681494 365464 688258
rect 365144 681258 365186 681494
rect 365422 681258 365464 681494
rect 365144 674494 365464 681258
rect 365144 674258 365186 674494
rect 365422 674258 365464 674494
rect 365144 667494 365464 674258
rect 365144 667258 365186 667494
rect 365422 667258 365464 667494
rect 365144 660494 365464 667258
rect 365144 660258 365186 660494
rect 365422 660258 365464 660494
rect 365144 653494 365464 660258
rect 365144 653258 365186 653494
rect 365422 653258 365464 653494
rect 365144 646494 365464 653258
rect 365144 646258 365186 646494
rect 365422 646258 365464 646494
rect 365144 639494 365464 646258
rect 365144 639258 365186 639494
rect 365422 639258 365464 639494
rect 365144 632494 365464 639258
rect 365144 632258 365186 632494
rect 365422 632258 365464 632494
rect 365144 625494 365464 632258
rect 365144 625258 365186 625494
rect 365422 625258 365464 625494
rect 365144 618494 365464 625258
rect 365144 618258 365186 618494
rect 365422 618258 365464 618494
rect 365144 611494 365464 618258
rect 365144 611258 365186 611494
rect 365422 611258 365464 611494
rect 365144 604494 365464 611258
rect 365144 604258 365186 604494
rect 365422 604258 365464 604494
rect 365144 597494 365464 604258
rect 365144 597258 365186 597494
rect 365422 597258 365464 597494
rect 365144 590494 365464 597258
rect 365144 590258 365186 590494
rect 365422 590258 365464 590494
rect 365144 583494 365464 590258
rect 365144 583258 365186 583494
rect 365422 583258 365464 583494
rect 365144 576494 365464 583258
rect 365144 576258 365186 576494
rect 365422 576258 365464 576494
rect 365144 569494 365464 576258
rect 365144 569258 365186 569494
rect 365422 569258 365464 569494
rect 365144 562494 365464 569258
rect 365144 562258 365186 562494
rect 365422 562258 365464 562494
rect 365144 555494 365464 562258
rect 365144 555258 365186 555494
rect 365422 555258 365464 555494
rect 365144 548494 365464 555258
rect 365144 548258 365186 548494
rect 365422 548258 365464 548494
rect 365144 541494 365464 548258
rect 365144 541258 365186 541494
rect 365422 541258 365464 541494
rect 365144 534494 365464 541258
rect 365144 534258 365186 534494
rect 365422 534258 365464 534494
rect 365144 527494 365464 534258
rect 365144 527258 365186 527494
rect 365422 527258 365464 527494
rect 365144 520494 365464 527258
rect 365144 520258 365186 520494
rect 365422 520258 365464 520494
rect 365144 513494 365464 520258
rect 365144 513258 365186 513494
rect 365422 513258 365464 513494
rect 365144 506494 365464 513258
rect 365144 506258 365186 506494
rect 365422 506258 365464 506494
rect 365144 499494 365464 506258
rect 365144 499258 365186 499494
rect 365422 499258 365464 499494
rect 365144 492494 365464 499258
rect 365144 492258 365186 492494
rect 365422 492258 365464 492494
rect 365144 485494 365464 492258
rect 365144 485258 365186 485494
rect 365422 485258 365464 485494
rect 365144 478494 365464 485258
rect 365144 478258 365186 478494
rect 365422 478258 365464 478494
rect 365144 471494 365464 478258
rect 365144 471258 365186 471494
rect 365422 471258 365464 471494
rect 365144 464494 365464 471258
rect 365144 464258 365186 464494
rect 365422 464258 365464 464494
rect 365144 457494 365464 464258
rect 365144 457258 365186 457494
rect 365422 457258 365464 457494
rect 365144 450494 365464 457258
rect 365144 450258 365186 450494
rect 365422 450258 365464 450494
rect 365144 443494 365464 450258
rect 365144 443258 365186 443494
rect 365422 443258 365464 443494
rect 365144 436494 365464 443258
rect 365144 436258 365186 436494
rect 365422 436258 365464 436494
rect 365144 429494 365464 436258
rect 365144 429258 365186 429494
rect 365422 429258 365464 429494
rect 365144 422494 365464 429258
rect 365144 422258 365186 422494
rect 365422 422258 365464 422494
rect 365144 415494 365464 422258
rect 365144 415258 365186 415494
rect 365422 415258 365464 415494
rect 365144 408494 365464 415258
rect 365144 408258 365186 408494
rect 365422 408258 365464 408494
rect 365144 401494 365464 408258
rect 365144 401258 365186 401494
rect 365422 401258 365464 401494
rect 365144 394494 365464 401258
rect 365144 394258 365186 394494
rect 365422 394258 365464 394494
rect 365144 387494 365464 394258
rect 365144 387258 365186 387494
rect 365422 387258 365464 387494
rect 365144 380494 365464 387258
rect 365144 380258 365186 380494
rect 365422 380258 365464 380494
rect 365144 373494 365464 380258
rect 365144 373258 365186 373494
rect 365422 373258 365464 373494
rect 365144 366494 365464 373258
rect 365144 366258 365186 366494
rect 365422 366258 365464 366494
rect 365144 359494 365464 366258
rect 365144 359258 365186 359494
rect 365422 359258 365464 359494
rect 365144 352494 365464 359258
rect 365144 352258 365186 352494
rect 365422 352258 365464 352494
rect 365144 345494 365464 352258
rect 365144 345258 365186 345494
rect 365422 345258 365464 345494
rect 365144 338494 365464 345258
rect 365144 338258 365186 338494
rect 365422 338258 365464 338494
rect 365144 331494 365464 338258
rect 365144 331258 365186 331494
rect 365422 331258 365464 331494
rect 365144 324494 365464 331258
rect 365144 324258 365186 324494
rect 365422 324258 365464 324494
rect 365144 317494 365464 324258
rect 365144 317258 365186 317494
rect 365422 317258 365464 317494
rect 365144 310494 365464 317258
rect 365144 310258 365186 310494
rect 365422 310258 365464 310494
rect 365144 303494 365464 310258
rect 365144 303258 365186 303494
rect 365422 303258 365464 303494
rect 365144 296494 365464 303258
rect 365144 296258 365186 296494
rect 365422 296258 365464 296494
rect 365144 289494 365464 296258
rect 365144 289258 365186 289494
rect 365422 289258 365464 289494
rect 365144 282494 365464 289258
rect 365144 282258 365186 282494
rect 365422 282258 365464 282494
rect 365144 275494 365464 282258
rect 365144 275258 365186 275494
rect 365422 275258 365464 275494
rect 365144 268494 365464 275258
rect 365144 268258 365186 268494
rect 365422 268258 365464 268494
rect 365144 261494 365464 268258
rect 365144 261258 365186 261494
rect 365422 261258 365464 261494
rect 365144 254494 365464 261258
rect 365144 254258 365186 254494
rect 365422 254258 365464 254494
rect 365144 247494 365464 254258
rect 365144 247258 365186 247494
rect 365422 247258 365464 247494
rect 365144 240494 365464 247258
rect 365144 240258 365186 240494
rect 365422 240258 365464 240494
rect 365144 233494 365464 240258
rect 365144 233258 365186 233494
rect 365422 233258 365464 233494
rect 365144 226494 365464 233258
rect 365144 226258 365186 226494
rect 365422 226258 365464 226494
rect 365144 219494 365464 226258
rect 365144 219258 365186 219494
rect 365422 219258 365464 219494
rect 365144 212494 365464 219258
rect 365144 212258 365186 212494
rect 365422 212258 365464 212494
rect 365144 205494 365464 212258
rect 365144 205258 365186 205494
rect 365422 205258 365464 205494
rect 365144 198494 365464 205258
rect 365144 198258 365186 198494
rect 365422 198258 365464 198494
rect 365144 191494 365464 198258
rect 365144 191258 365186 191494
rect 365422 191258 365464 191494
rect 365144 184494 365464 191258
rect 365144 184258 365186 184494
rect 365422 184258 365464 184494
rect 365144 177494 365464 184258
rect 365144 177258 365186 177494
rect 365422 177258 365464 177494
rect 365144 170494 365464 177258
rect 365144 170258 365186 170494
rect 365422 170258 365464 170494
rect 365144 163494 365464 170258
rect 365144 163258 365186 163494
rect 365422 163258 365464 163494
rect 365144 156494 365464 163258
rect 365144 156258 365186 156494
rect 365422 156258 365464 156494
rect 365144 149494 365464 156258
rect 365144 149258 365186 149494
rect 365422 149258 365464 149494
rect 365144 142494 365464 149258
rect 365144 142258 365186 142494
rect 365422 142258 365464 142494
rect 365144 135494 365464 142258
rect 365144 135258 365186 135494
rect 365422 135258 365464 135494
rect 365144 128494 365464 135258
rect 365144 128258 365186 128494
rect 365422 128258 365464 128494
rect 365144 121494 365464 128258
rect 365144 121258 365186 121494
rect 365422 121258 365464 121494
rect 365144 114494 365464 121258
rect 365144 114258 365186 114494
rect 365422 114258 365464 114494
rect 365144 107494 365464 114258
rect 365144 107258 365186 107494
rect 365422 107258 365464 107494
rect 365144 100494 365464 107258
rect 365144 100258 365186 100494
rect 365422 100258 365464 100494
rect 365144 93494 365464 100258
rect 365144 93258 365186 93494
rect 365422 93258 365464 93494
rect 365144 86494 365464 93258
rect 365144 86258 365186 86494
rect 365422 86258 365464 86494
rect 365144 79494 365464 86258
rect 365144 79258 365186 79494
rect 365422 79258 365464 79494
rect 365144 72494 365464 79258
rect 365144 72258 365186 72494
rect 365422 72258 365464 72494
rect 365144 65494 365464 72258
rect 365144 65258 365186 65494
rect 365422 65258 365464 65494
rect 365144 58494 365464 65258
rect 365144 58258 365186 58494
rect 365422 58258 365464 58494
rect 365144 51494 365464 58258
rect 365144 51258 365186 51494
rect 365422 51258 365464 51494
rect 365144 44494 365464 51258
rect 365144 44258 365186 44494
rect 365422 44258 365464 44494
rect 365144 37494 365464 44258
rect 365144 37258 365186 37494
rect 365422 37258 365464 37494
rect 365144 30494 365464 37258
rect 365144 30258 365186 30494
rect 365422 30258 365464 30494
rect 365144 23494 365464 30258
rect 365144 23258 365186 23494
rect 365422 23258 365464 23494
rect 365144 16494 365464 23258
rect 365144 16258 365186 16494
rect 365422 16258 365464 16494
rect 365144 9494 365464 16258
rect 365144 9258 365186 9494
rect 365422 9258 365464 9494
rect 365144 2494 365464 9258
rect 365144 2258 365186 2494
rect 365422 2258 365464 2494
rect 365144 -746 365464 2258
rect 365144 -982 365186 -746
rect 365422 -982 365464 -746
rect 365144 -1066 365464 -982
rect 365144 -1302 365186 -1066
rect 365422 -1302 365464 -1066
rect 365144 -2294 365464 -1302
rect 366876 706198 367196 706230
rect 366876 705962 366918 706198
rect 367154 705962 367196 706198
rect 366876 705878 367196 705962
rect 366876 705642 366918 705878
rect 367154 705642 367196 705878
rect 366876 696561 367196 705642
rect 366876 696325 366918 696561
rect 367154 696325 367196 696561
rect 366876 689561 367196 696325
rect 366876 689325 366918 689561
rect 367154 689325 367196 689561
rect 366876 682561 367196 689325
rect 366876 682325 366918 682561
rect 367154 682325 367196 682561
rect 366876 675561 367196 682325
rect 366876 675325 366918 675561
rect 367154 675325 367196 675561
rect 366876 668561 367196 675325
rect 366876 668325 366918 668561
rect 367154 668325 367196 668561
rect 366876 661561 367196 668325
rect 366876 661325 366918 661561
rect 367154 661325 367196 661561
rect 366876 654561 367196 661325
rect 366876 654325 366918 654561
rect 367154 654325 367196 654561
rect 366876 647561 367196 654325
rect 366876 647325 366918 647561
rect 367154 647325 367196 647561
rect 366876 640561 367196 647325
rect 366876 640325 366918 640561
rect 367154 640325 367196 640561
rect 366876 633561 367196 640325
rect 366876 633325 366918 633561
rect 367154 633325 367196 633561
rect 366876 626561 367196 633325
rect 366876 626325 366918 626561
rect 367154 626325 367196 626561
rect 366876 619561 367196 626325
rect 366876 619325 366918 619561
rect 367154 619325 367196 619561
rect 366876 612561 367196 619325
rect 366876 612325 366918 612561
rect 367154 612325 367196 612561
rect 366876 605561 367196 612325
rect 366876 605325 366918 605561
rect 367154 605325 367196 605561
rect 366876 598561 367196 605325
rect 366876 598325 366918 598561
rect 367154 598325 367196 598561
rect 366876 591561 367196 598325
rect 366876 591325 366918 591561
rect 367154 591325 367196 591561
rect 366876 584561 367196 591325
rect 366876 584325 366918 584561
rect 367154 584325 367196 584561
rect 366876 577561 367196 584325
rect 366876 577325 366918 577561
rect 367154 577325 367196 577561
rect 366876 570561 367196 577325
rect 366876 570325 366918 570561
rect 367154 570325 367196 570561
rect 366876 563561 367196 570325
rect 366876 563325 366918 563561
rect 367154 563325 367196 563561
rect 366876 556561 367196 563325
rect 366876 556325 366918 556561
rect 367154 556325 367196 556561
rect 366876 549561 367196 556325
rect 366876 549325 366918 549561
rect 367154 549325 367196 549561
rect 366876 542561 367196 549325
rect 366876 542325 366918 542561
rect 367154 542325 367196 542561
rect 366876 535561 367196 542325
rect 366876 535325 366918 535561
rect 367154 535325 367196 535561
rect 366876 528561 367196 535325
rect 366876 528325 366918 528561
rect 367154 528325 367196 528561
rect 366876 521561 367196 528325
rect 366876 521325 366918 521561
rect 367154 521325 367196 521561
rect 366876 514561 367196 521325
rect 366876 514325 366918 514561
rect 367154 514325 367196 514561
rect 366876 507561 367196 514325
rect 366876 507325 366918 507561
rect 367154 507325 367196 507561
rect 366876 500561 367196 507325
rect 366876 500325 366918 500561
rect 367154 500325 367196 500561
rect 366876 493561 367196 500325
rect 366876 493325 366918 493561
rect 367154 493325 367196 493561
rect 366876 486561 367196 493325
rect 366876 486325 366918 486561
rect 367154 486325 367196 486561
rect 366876 479561 367196 486325
rect 366876 479325 366918 479561
rect 367154 479325 367196 479561
rect 366876 472561 367196 479325
rect 366876 472325 366918 472561
rect 367154 472325 367196 472561
rect 366876 465561 367196 472325
rect 366876 465325 366918 465561
rect 367154 465325 367196 465561
rect 366876 458561 367196 465325
rect 366876 458325 366918 458561
rect 367154 458325 367196 458561
rect 366876 451561 367196 458325
rect 366876 451325 366918 451561
rect 367154 451325 367196 451561
rect 366876 444561 367196 451325
rect 366876 444325 366918 444561
rect 367154 444325 367196 444561
rect 366876 437561 367196 444325
rect 366876 437325 366918 437561
rect 367154 437325 367196 437561
rect 366876 430561 367196 437325
rect 366876 430325 366918 430561
rect 367154 430325 367196 430561
rect 366876 423561 367196 430325
rect 366876 423325 366918 423561
rect 367154 423325 367196 423561
rect 366876 416561 367196 423325
rect 366876 416325 366918 416561
rect 367154 416325 367196 416561
rect 366876 409561 367196 416325
rect 366876 409325 366918 409561
rect 367154 409325 367196 409561
rect 366876 402561 367196 409325
rect 366876 402325 366918 402561
rect 367154 402325 367196 402561
rect 366876 395561 367196 402325
rect 366876 395325 366918 395561
rect 367154 395325 367196 395561
rect 366876 388561 367196 395325
rect 366876 388325 366918 388561
rect 367154 388325 367196 388561
rect 366876 381561 367196 388325
rect 366876 381325 366918 381561
rect 367154 381325 367196 381561
rect 366876 374561 367196 381325
rect 366876 374325 366918 374561
rect 367154 374325 367196 374561
rect 366876 367561 367196 374325
rect 366876 367325 366918 367561
rect 367154 367325 367196 367561
rect 366876 360561 367196 367325
rect 366876 360325 366918 360561
rect 367154 360325 367196 360561
rect 366876 353561 367196 360325
rect 366876 353325 366918 353561
rect 367154 353325 367196 353561
rect 366876 346561 367196 353325
rect 366876 346325 366918 346561
rect 367154 346325 367196 346561
rect 366876 339561 367196 346325
rect 366876 339325 366918 339561
rect 367154 339325 367196 339561
rect 366876 332561 367196 339325
rect 366876 332325 366918 332561
rect 367154 332325 367196 332561
rect 366876 325561 367196 332325
rect 366876 325325 366918 325561
rect 367154 325325 367196 325561
rect 366876 318561 367196 325325
rect 366876 318325 366918 318561
rect 367154 318325 367196 318561
rect 366876 311561 367196 318325
rect 366876 311325 366918 311561
rect 367154 311325 367196 311561
rect 366876 304561 367196 311325
rect 366876 304325 366918 304561
rect 367154 304325 367196 304561
rect 366876 297561 367196 304325
rect 366876 297325 366918 297561
rect 367154 297325 367196 297561
rect 366876 290561 367196 297325
rect 366876 290325 366918 290561
rect 367154 290325 367196 290561
rect 366876 283561 367196 290325
rect 366876 283325 366918 283561
rect 367154 283325 367196 283561
rect 366876 276561 367196 283325
rect 366876 276325 366918 276561
rect 367154 276325 367196 276561
rect 366876 269561 367196 276325
rect 366876 269325 366918 269561
rect 367154 269325 367196 269561
rect 366876 262561 367196 269325
rect 366876 262325 366918 262561
rect 367154 262325 367196 262561
rect 366876 255561 367196 262325
rect 366876 255325 366918 255561
rect 367154 255325 367196 255561
rect 366876 248561 367196 255325
rect 366876 248325 366918 248561
rect 367154 248325 367196 248561
rect 366876 241561 367196 248325
rect 366876 241325 366918 241561
rect 367154 241325 367196 241561
rect 366876 234561 367196 241325
rect 366876 234325 366918 234561
rect 367154 234325 367196 234561
rect 366876 227561 367196 234325
rect 366876 227325 366918 227561
rect 367154 227325 367196 227561
rect 366876 220561 367196 227325
rect 366876 220325 366918 220561
rect 367154 220325 367196 220561
rect 366876 213561 367196 220325
rect 366876 213325 366918 213561
rect 367154 213325 367196 213561
rect 366876 206561 367196 213325
rect 366876 206325 366918 206561
rect 367154 206325 367196 206561
rect 366876 199561 367196 206325
rect 366876 199325 366918 199561
rect 367154 199325 367196 199561
rect 366876 192561 367196 199325
rect 366876 192325 366918 192561
rect 367154 192325 367196 192561
rect 366876 185561 367196 192325
rect 366876 185325 366918 185561
rect 367154 185325 367196 185561
rect 366876 178561 367196 185325
rect 366876 178325 366918 178561
rect 367154 178325 367196 178561
rect 366876 171561 367196 178325
rect 366876 171325 366918 171561
rect 367154 171325 367196 171561
rect 366876 164561 367196 171325
rect 366876 164325 366918 164561
rect 367154 164325 367196 164561
rect 366876 157561 367196 164325
rect 366876 157325 366918 157561
rect 367154 157325 367196 157561
rect 366876 150561 367196 157325
rect 366876 150325 366918 150561
rect 367154 150325 367196 150561
rect 366876 143561 367196 150325
rect 366876 143325 366918 143561
rect 367154 143325 367196 143561
rect 366876 136561 367196 143325
rect 366876 136325 366918 136561
rect 367154 136325 367196 136561
rect 366876 129561 367196 136325
rect 366876 129325 366918 129561
rect 367154 129325 367196 129561
rect 366876 122561 367196 129325
rect 366876 122325 366918 122561
rect 367154 122325 367196 122561
rect 366876 115561 367196 122325
rect 366876 115325 366918 115561
rect 367154 115325 367196 115561
rect 366876 108561 367196 115325
rect 366876 108325 366918 108561
rect 367154 108325 367196 108561
rect 366876 101561 367196 108325
rect 366876 101325 366918 101561
rect 367154 101325 367196 101561
rect 366876 94561 367196 101325
rect 366876 94325 366918 94561
rect 367154 94325 367196 94561
rect 366876 87561 367196 94325
rect 366876 87325 366918 87561
rect 367154 87325 367196 87561
rect 366876 80561 367196 87325
rect 366876 80325 366918 80561
rect 367154 80325 367196 80561
rect 366876 73561 367196 80325
rect 366876 73325 366918 73561
rect 367154 73325 367196 73561
rect 366876 66561 367196 73325
rect 366876 66325 366918 66561
rect 367154 66325 367196 66561
rect 366876 59561 367196 66325
rect 366876 59325 366918 59561
rect 367154 59325 367196 59561
rect 366876 52561 367196 59325
rect 366876 52325 366918 52561
rect 367154 52325 367196 52561
rect 366876 45561 367196 52325
rect 366876 45325 366918 45561
rect 367154 45325 367196 45561
rect 366876 38561 367196 45325
rect 366876 38325 366918 38561
rect 367154 38325 367196 38561
rect 366876 31561 367196 38325
rect 366876 31325 366918 31561
rect 367154 31325 367196 31561
rect 366876 24561 367196 31325
rect 366876 24325 366918 24561
rect 367154 24325 367196 24561
rect 366876 17561 367196 24325
rect 366876 17325 366918 17561
rect 367154 17325 367196 17561
rect 366876 10561 367196 17325
rect 366876 10325 366918 10561
rect 367154 10325 367196 10561
rect 366876 3561 367196 10325
rect 366876 3325 366918 3561
rect 367154 3325 367196 3561
rect 366876 -1706 367196 3325
rect 366876 -1942 366918 -1706
rect 367154 -1942 367196 -1706
rect 366876 -2026 367196 -1942
rect 366876 -2262 366918 -2026
rect 367154 -2262 367196 -2026
rect 366876 -2294 367196 -2262
rect 372144 705238 372464 706230
rect 372144 705002 372186 705238
rect 372422 705002 372464 705238
rect 372144 704918 372464 705002
rect 372144 704682 372186 704918
rect 372422 704682 372464 704918
rect 372144 695494 372464 704682
rect 372144 695258 372186 695494
rect 372422 695258 372464 695494
rect 372144 688494 372464 695258
rect 372144 688258 372186 688494
rect 372422 688258 372464 688494
rect 372144 681494 372464 688258
rect 372144 681258 372186 681494
rect 372422 681258 372464 681494
rect 372144 674494 372464 681258
rect 372144 674258 372186 674494
rect 372422 674258 372464 674494
rect 372144 667494 372464 674258
rect 372144 667258 372186 667494
rect 372422 667258 372464 667494
rect 372144 660494 372464 667258
rect 372144 660258 372186 660494
rect 372422 660258 372464 660494
rect 372144 653494 372464 660258
rect 372144 653258 372186 653494
rect 372422 653258 372464 653494
rect 372144 646494 372464 653258
rect 372144 646258 372186 646494
rect 372422 646258 372464 646494
rect 372144 639494 372464 646258
rect 372144 639258 372186 639494
rect 372422 639258 372464 639494
rect 372144 632494 372464 639258
rect 372144 632258 372186 632494
rect 372422 632258 372464 632494
rect 372144 625494 372464 632258
rect 372144 625258 372186 625494
rect 372422 625258 372464 625494
rect 372144 618494 372464 625258
rect 372144 618258 372186 618494
rect 372422 618258 372464 618494
rect 372144 611494 372464 618258
rect 372144 611258 372186 611494
rect 372422 611258 372464 611494
rect 372144 604494 372464 611258
rect 372144 604258 372186 604494
rect 372422 604258 372464 604494
rect 372144 597494 372464 604258
rect 372144 597258 372186 597494
rect 372422 597258 372464 597494
rect 372144 590494 372464 597258
rect 372144 590258 372186 590494
rect 372422 590258 372464 590494
rect 372144 583494 372464 590258
rect 372144 583258 372186 583494
rect 372422 583258 372464 583494
rect 372144 576494 372464 583258
rect 372144 576258 372186 576494
rect 372422 576258 372464 576494
rect 372144 569494 372464 576258
rect 372144 569258 372186 569494
rect 372422 569258 372464 569494
rect 372144 562494 372464 569258
rect 372144 562258 372186 562494
rect 372422 562258 372464 562494
rect 372144 555494 372464 562258
rect 372144 555258 372186 555494
rect 372422 555258 372464 555494
rect 372144 548494 372464 555258
rect 372144 548258 372186 548494
rect 372422 548258 372464 548494
rect 372144 541494 372464 548258
rect 372144 541258 372186 541494
rect 372422 541258 372464 541494
rect 372144 534494 372464 541258
rect 372144 534258 372186 534494
rect 372422 534258 372464 534494
rect 372144 527494 372464 534258
rect 372144 527258 372186 527494
rect 372422 527258 372464 527494
rect 372144 520494 372464 527258
rect 372144 520258 372186 520494
rect 372422 520258 372464 520494
rect 372144 513494 372464 520258
rect 372144 513258 372186 513494
rect 372422 513258 372464 513494
rect 372144 506494 372464 513258
rect 372144 506258 372186 506494
rect 372422 506258 372464 506494
rect 372144 499494 372464 506258
rect 372144 499258 372186 499494
rect 372422 499258 372464 499494
rect 372144 492494 372464 499258
rect 372144 492258 372186 492494
rect 372422 492258 372464 492494
rect 372144 485494 372464 492258
rect 372144 485258 372186 485494
rect 372422 485258 372464 485494
rect 372144 478494 372464 485258
rect 372144 478258 372186 478494
rect 372422 478258 372464 478494
rect 372144 471494 372464 478258
rect 372144 471258 372186 471494
rect 372422 471258 372464 471494
rect 372144 464494 372464 471258
rect 372144 464258 372186 464494
rect 372422 464258 372464 464494
rect 372144 457494 372464 464258
rect 372144 457258 372186 457494
rect 372422 457258 372464 457494
rect 372144 450494 372464 457258
rect 372144 450258 372186 450494
rect 372422 450258 372464 450494
rect 372144 443494 372464 450258
rect 372144 443258 372186 443494
rect 372422 443258 372464 443494
rect 372144 436494 372464 443258
rect 372144 436258 372186 436494
rect 372422 436258 372464 436494
rect 372144 429494 372464 436258
rect 372144 429258 372186 429494
rect 372422 429258 372464 429494
rect 372144 422494 372464 429258
rect 372144 422258 372186 422494
rect 372422 422258 372464 422494
rect 372144 415494 372464 422258
rect 372144 415258 372186 415494
rect 372422 415258 372464 415494
rect 372144 408494 372464 415258
rect 372144 408258 372186 408494
rect 372422 408258 372464 408494
rect 372144 401494 372464 408258
rect 372144 401258 372186 401494
rect 372422 401258 372464 401494
rect 372144 394494 372464 401258
rect 372144 394258 372186 394494
rect 372422 394258 372464 394494
rect 372144 387494 372464 394258
rect 372144 387258 372186 387494
rect 372422 387258 372464 387494
rect 372144 380494 372464 387258
rect 372144 380258 372186 380494
rect 372422 380258 372464 380494
rect 372144 373494 372464 380258
rect 372144 373258 372186 373494
rect 372422 373258 372464 373494
rect 372144 366494 372464 373258
rect 372144 366258 372186 366494
rect 372422 366258 372464 366494
rect 372144 359494 372464 366258
rect 372144 359258 372186 359494
rect 372422 359258 372464 359494
rect 372144 352494 372464 359258
rect 372144 352258 372186 352494
rect 372422 352258 372464 352494
rect 372144 345494 372464 352258
rect 372144 345258 372186 345494
rect 372422 345258 372464 345494
rect 372144 338494 372464 345258
rect 372144 338258 372186 338494
rect 372422 338258 372464 338494
rect 372144 331494 372464 338258
rect 372144 331258 372186 331494
rect 372422 331258 372464 331494
rect 372144 324494 372464 331258
rect 372144 324258 372186 324494
rect 372422 324258 372464 324494
rect 372144 317494 372464 324258
rect 372144 317258 372186 317494
rect 372422 317258 372464 317494
rect 372144 310494 372464 317258
rect 372144 310258 372186 310494
rect 372422 310258 372464 310494
rect 372144 303494 372464 310258
rect 372144 303258 372186 303494
rect 372422 303258 372464 303494
rect 372144 296494 372464 303258
rect 372144 296258 372186 296494
rect 372422 296258 372464 296494
rect 372144 289494 372464 296258
rect 372144 289258 372186 289494
rect 372422 289258 372464 289494
rect 372144 282494 372464 289258
rect 372144 282258 372186 282494
rect 372422 282258 372464 282494
rect 372144 275494 372464 282258
rect 372144 275258 372186 275494
rect 372422 275258 372464 275494
rect 372144 268494 372464 275258
rect 372144 268258 372186 268494
rect 372422 268258 372464 268494
rect 372144 261494 372464 268258
rect 372144 261258 372186 261494
rect 372422 261258 372464 261494
rect 372144 254494 372464 261258
rect 372144 254258 372186 254494
rect 372422 254258 372464 254494
rect 372144 247494 372464 254258
rect 372144 247258 372186 247494
rect 372422 247258 372464 247494
rect 372144 240494 372464 247258
rect 372144 240258 372186 240494
rect 372422 240258 372464 240494
rect 372144 233494 372464 240258
rect 372144 233258 372186 233494
rect 372422 233258 372464 233494
rect 372144 226494 372464 233258
rect 372144 226258 372186 226494
rect 372422 226258 372464 226494
rect 372144 219494 372464 226258
rect 372144 219258 372186 219494
rect 372422 219258 372464 219494
rect 372144 212494 372464 219258
rect 372144 212258 372186 212494
rect 372422 212258 372464 212494
rect 372144 205494 372464 212258
rect 372144 205258 372186 205494
rect 372422 205258 372464 205494
rect 372144 198494 372464 205258
rect 372144 198258 372186 198494
rect 372422 198258 372464 198494
rect 372144 191494 372464 198258
rect 372144 191258 372186 191494
rect 372422 191258 372464 191494
rect 372144 184494 372464 191258
rect 372144 184258 372186 184494
rect 372422 184258 372464 184494
rect 372144 177494 372464 184258
rect 372144 177258 372186 177494
rect 372422 177258 372464 177494
rect 372144 170494 372464 177258
rect 372144 170258 372186 170494
rect 372422 170258 372464 170494
rect 372144 163494 372464 170258
rect 372144 163258 372186 163494
rect 372422 163258 372464 163494
rect 372144 156494 372464 163258
rect 372144 156258 372186 156494
rect 372422 156258 372464 156494
rect 372144 149494 372464 156258
rect 372144 149258 372186 149494
rect 372422 149258 372464 149494
rect 372144 142494 372464 149258
rect 372144 142258 372186 142494
rect 372422 142258 372464 142494
rect 372144 135494 372464 142258
rect 372144 135258 372186 135494
rect 372422 135258 372464 135494
rect 372144 128494 372464 135258
rect 372144 128258 372186 128494
rect 372422 128258 372464 128494
rect 372144 121494 372464 128258
rect 372144 121258 372186 121494
rect 372422 121258 372464 121494
rect 372144 114494 372464 121258
rect 372144 114258 372186 114494
rect 372422 114258 372464 114494
rect 372144 107494 372464 114258
rect 372144 107258 372186 107494
rect 372422 107258 372464 107494
rect 372144 100494 372464 107258
rect 372144 100258 372186 100494
rect 372422 100258 372464 100494
rect 372144 93494 372464 100258
rect 372144 93258 372186 93494
rect 372422 93258 372464 93494
rect 372144 86494 372464 93258
rect 372144 86258 372186 86494
rect 372422 86258 372464 86494
rect 372144 79494 372464 86258
rect 372144 79258 372186 79494
rect 372422 79258 372464 79494
rect 372144 72494 372464 79258
rect 372144 72258 372186 72494
rect 372422 72258 372464 72494
rect 372144 65494 372464 72258
rect 372144 65258 372186 65494
rect 372422 65258 372464 65494
rect 372144 58494 372464 65258
rect 372144 58258 372186 58494
rect 372422 58258 372464 58494
rect 372144 51494 372464 58258
rect 372144 51258 372186 51494
rect 372422 51258 372464 51494
rect 372144 44494 372464 51258
rect 372144 44258 372186 44494
rect 372422 44258 372464 44494
rect 372144 37494 372464 44258
rect 372144 37258 372186 37494
rect 372422 37258 372464 37494
rect 372144 30494 372464 37258
rect 372144 30258 372186 30494
rect 372422 30258 372464 30494
rect 372144 23494 372464 30258
rect 372144 23258 372186 23494
rect 372422 23258 372464 23494
rect 372144 16494 372464 23258
rect 372144 16258 372186 16494
rect 372422 16258 372464 16494
rect 372144 9494 372464 16258
rect 372144 9258 372186 9494
rect 372422 9258 372464 9494
rect 372144 2494 372464 9258
rect 372144 2258 372186 2494
rect 372422 2258 372464 2494
rect 372144 -746 372464 2258
rect 372144 -982 372186 -746
rect 372422 -982 372464 -746
rect 372144 -1066 372464 -982
rect 372144 -1302 372186 -1066
rect 372422 -1302 372464 -1066
rect 372144 -2294 372464 -1302
rect 373876 706198 374196 706230
rect 373876 705962 373918 706198
rect 374154 705962 374196 706198
rect 373876 705878 374196 705962
rect 373876 705642 373918 705878
rect 374154 705642 374196 705878
rect 373876 696561 374196 705642
rect 373876 696325 373918 696561
rect 374154 696325 374196 696561
rect 373876 689561 374196 696325
rect 373876 689325 373918 689561
rect 374154 689325 374196 689561
rect 373876 682561 374196 689325
rect 373876 682325 373918 682561
rect 374154 682325 374196 682561
rect 373876 675561 374196 682325
rect 373876 675325 373918 675561
rect 374154 675325 374196 675561
rect 373876 668561 374196 675325
rect 373876 668325 373918 668561
rect 374154 668325 374196 668561
rect 373876 661561 374196 668325
rect 373876 661325 373918 661561
rect 374154 661325 374196 661561
rect 373876 654561 374196 661325
rect 373876 654325 373918 654561
rect 374154 654325 374196 654561
rect 373876 647561 374196 654325
rect 373876 647325 373918 647561
rect 374154 647325 374196 647561
rect 373876 640561 374196 647325
rect 373876 640325 373918 640561
rect 374154 640325 374196 640561
rect 373876 633561 374196 640325
rect 373876 633325 373918 633561
rect 374154 633325 374196 633561
rect 373876 626561 374196 633325
rect 373876 626325 373918 626561
rect 374154 626325 374196 626561
rect 373876 619561 374196 626325
rect 373876 619325 373918 619561
rect 374154 619325 374196 619561
rect 373876 612561 374196 619325
rect 373876 612325 373918 612561
rect 374154 612325 374196 612561
rect 373876 605561 374196 612325
rect 373876 605325 373918 605561
rect 374154 605325 374196 605561
rect 373876 598561 374196 605325
rect 373876 598325 373918 598561
rect 374154 598325 374196 598561
rect 373876 591561 374196 598325
rect 373876 591325 373918 591561
rect 374154 591325 374196 591561
rect 373876 584561 374196 591325
rect 373876 584325 373918 584561
rect 374154 584325 374196 584561
rect 373876 577561 374196 584325
rect 373876 577325 373918 577561
rect 374154 577325 374196 577561
rect 373876 570561 374196 577325
rect 373876 570325 373918 570561
rect 374154 570325 374196 570561
rect 373876 563561 374196 570325
rect 373876 563325 373918 563561
rect 374154 563325 374196 563561
rect 373876 556561 374196 563325
rect 373876 556325 373918 556561
rect 374154 556325 374196 556561
rect 373876 549561 374196 556325
rect 373876 549325 373918 549561
rect 374154 549325 374196 549561
rect 373876 542561 374196 549325
rect 373876 542325 373918 542561
rect 374154 542325 374196 542561
rect 373876 535561 374196 542325
rect 373876 535325 373918 535561
rect 374154 535325 374196 535561
rect 373876 528561 374196 535325
rect 373876 528325 373918 528561
rect 374154 528325 374196 528561
rect 373876 521561 374196 528325
rect 373876 521325 373918 521561
rect 374154 521325 374196 521561
rect 373876 514561 374196 521325
rect 373876 514325 373918 514561
rect 374154 514325 374196 514561
rect 373876 507561 374196 514325
rect 373876 507325 373918 507561
rect 374154 507325 374196 507561
rect 373876 500561 374196 507325
rect 373876 500325 373918 500561
rect 374154 500325 374196 500561
rect 373876 493561 374196 500325
rect 373876 493325 373918 493561
rect 374154 493325 374196 493561
rect 373876 486561 374196 493325
rect 373876 486325 373918 486561
rect 374154 486325 374196 486561
rect 373876 479561 374196 486325
rect 373876 479325 373918 479561
rect 374154 479325 374196 479561
rect 373876 472561 374196 479325
rect 373876 472325 373918 472561
rect 374154 472325 374196 472561
rect 373876 465561 374196 472325
rect 373876 465325 373918 465561
rect 374154 465325 374196 465561
rect 373876 458561 374196 465325
rect 373876 458325 373918 458561
rect 374154 458325 374196 458561
rect 373876 451561 374196 458325
rect 373876 451325 373918 451561
rect 374154 451325 374196 451561
rect 373876 444561 374196 451325
rect 373876 444325 373918 444561
rect 374154 444325 374196 444561
rect 373876 437561 374196 444325
rect 373876 437325 373918 437561
rect 374154 437325 374196 437561
rect 373876 430561 374196 437325
rect 373876 430325 373918 430561
rect 374154 430325 374196 430561
rect 373876 423561 374196 430325
rect 373876 423325 373918 423561
rect 374154 423325 374196 423561
rect 373876 416561 374196 423325
rect 373876 416325 373918 416561
rect 374154 416325 374196 416561
rect 373876 409561 374196 416325
rect 373876 409325 373918 409561
rect 374154 409325 374196 409561
rect 373876 402561 374196 409325
rect 373876 402325 373918 402561
rect 374154 402325 374196 402561
rect 373876 395561 374196 402325
rect 373876 395325 373918 395561
rect 374154 395325 374196 395561
rect 373876 388561 374196 395325
rect 373876 388325 373918 388561
rect 374154 388325 374196 388561
rect 373876 381561 374196 388325
rect 373876 381325 373918 381561
rect 374154 381325 374196 381561
rect 373876 374561 374196 381325
rect 373876 374325 373918 374561
rect 374154 374325 374196 374561
rect 373876 367561 374196 374325
rect 373876 367325 373918 367561
rect 374154 367325 374196 367561
rect 373876 360561 374196 367325
rect 373876 360325 373918 360561
rect 374154 360325 374196 360561
rect 373876 353561 374196 360325
rect 373876 353325 373918 353561
rect 374154 353325 374196 353561
rect 373876 346561 374196 353325
rect 373876 346325 373918 346561
rect 374154 346325 374196 346561
rect 373876 339561 374196 346325
rect 373876 339325 373918 339561
rect 374154 339325 374196 339561
rect 373876 332561 374196 339325
rect 373876 332325 373918 332561
rect 374154 332325 374196 332561
rect 373876 325561 374196 332325
rect 373876 325325 373918 325561
rect 374154 325325 374196 325561
rect 373876 318561 374196 325325
rect 373876 318325 373918 318561
rect 374154 318325 374196 318561
rect 373876 311561 374196 318325
rect 373876 311325 373918 311561
rect 374154 311325 374196 311561
rect 373876 304561 374196 311325
rect 373876 304325 373918 304561
rect 374154 304325 374196 304561
rect 373876 297561 374196 304325
rect 373876 297325 373918 297561
rect 374154 297325 374196 297561
rect 373876 290561 374196 297325
rect 373876 290325 373918 290561
rect 374154 290325 374196 290561
rect 373876 283561 374196 290325
rect 373876 283325 373918 283561
rect 374154 283325 374196 283561
rect 373876 276561 374196 283325
rect 373876 276325 373918 276561
rect 374154 276325 374196 276561
rect 373876 269561 374196 276325
rect 373876 269325 373918 269561
rect 374154 269325 374196 269561
rect 373876 262561 374196 269325
rect 373876 262325 373918 262561
rect 374154 262325 374196 262561
rect 373876 255561 374196 262325
rect 373876 255325 373918 255561
rect 374154 255325 374196 255561
rect 373876 248561 374196 255325
rect 373876 248325 373918 248561
rect 374154 248325 374196 248561
rect 373876 241561 374196 248325
rect 373876 241325 373918 241561
rect 374154 241325 374196 241561
rect 373876 234561 374196 241325
rect 373876 234325 373918 234561
rect 374154 234325 374196 234561
rect 373876 227561 374196 234325
rect 373876 227325 373918 227561
rect 374154 227325 374196 227561
rect 373876 220561 374196 227325
rect 373876 220325 373918 220561
rect 374154 220325 374196 220561
rect 373876 213561 374196 220325
rect 373876 213325 373918 213561
rect 374154 213325 374196 213561
rect 373876 206561 374196 213325
rect 373876 206325 373918 206561
rect 374154 206325 374196 206561
rect 373876 199561 374196 206325
rect 373876 199325 373918 199561
rect 374154 199325 374196 199561
rect 373876 192561 374196 199325
rect 373876 192325 373918 192561
rect 374154 192325 374196 192561
rect 373876 185561 374196 192325
rect 373876 185325 373918 185561
rect 374154 185325 374196 185561
rect 373876 178561 374196 185325
rect 373876 178325 373918 178561
rect 374154 178325 374196 178561
rect 373876 171561 374196 178325
rect 373876 171325 373918 171561
rect 374154 171325 374196 171561
rect 373876 164561 374196 171325
rect 373876 164325 373918 164561
rect 374154 164325 374196 164561
rect 373876 157561 374196 164325
rect 373876 157325 373918 157561
rect 374154 157325 374196 157561
rect 373876 150561 374196 157325
rect 373876 150325 373918 150561
rect 374154 150325 374196 150561
rect 373876 143561 374196 150325
rect 373876 143325 373918 143561
rect 374154 143325 374196 143561
rect 373876 136561 374196 143325
rect 373876 136325 373918 136561
rect 374154 136325 374196 136561
rect 373876 129561 374196 136325
rect 373876 129325 373918 129561
rect 374154 129325 374196 129561
rect 373876 122561 374196 129325
rect 373876 122325 373918 122561
rect 374154 122325 374196 122561
rect 373876 115561 374196 122325
rect 373876 115325 373918 115561
rect 374154 115325 374196 115561
rect 373876 108561 374196 115325
rect 373876 108325 373918 108561
rect 374154 108325 374196 108561
rect 373876 101561 374196 108325
rect 373876 101325 373918 101561
rect 374154 101325 374196 101561
rect 373876 94561 374196 101325
rect 373876 94325 373918 94561
rect 374154 94325 374196 94561
rect 373876 87561 374196 94325
rect 373876 87325 373918 87561
rect 374154 87325 374196 87561
rect 373876 80561 374196 87325
rect 373876 80325 373918 80561
rect 374154 80325 374196 80561
rect 373876 73561 374196 80325
rect 373876 73325 373918 73561
rect 374154 73325 374196 73561
rect 373876 66561 374196 73325
rect 373876 66325 373918 66561
rect 374154 66325 374196 66561
rect 373876 59561 374196 66325
rect 373876 59325 373918 59561
rect 374154 59325 374196 59561
rect 373876 52561 374196 59325
rect 373876 52325 373918 52561
rect 374154 52325 374196 52561
rect 373876 45561 374196 52325
rect 373876 45325 373918 45561
rect 374154 45325 374196 45561
rect 373876 38561 374196 45325
rect 373876 38325 373918 38561
rect 374154 38325 374196 38561
rect 373876 31561 374196 38325
rect 373876 31325 373918 31561
rect 374154 31325 374196 31561
rect 373876 24561 374196 31325
rect 373876 24325 373918 24561
rect 374154 24325 374196 24561
rect 373876 17561 374196 24325
rect 373876 17325 373918 17561
rect 374154 17325 374196 17561
rect 373876 10561 374196 17325
rect 373876 10325 373918 10561
rect 374154 10325 374196 10561
rect 373876 3561 374196 10325
rect 373876 3325 373918 3561
rect 374154 3325 374196 3561
rect 373876 -1706 374196 3325
rect 373876 -1942 373918 -1706
rect 374154 -1942 374196 -1706
rect 373876 -2026 374196 -1942
rect 373876 -2262 373918 -2026
rect 374154 -2262 374196 -2026
rect 373876 -2294 374196 -2262
rect 379144 705238 379464 706230
rect 379144 705002 379186 705238
rect 379422 705002 379464 705238
rect 379144 704918 379464 705002
rect 379144 704682 379186 704918
rect 379422 704682 379464 704918
rect 379144 695494 379464 704682
rect 379144 695258 379186 695494
rect 379422 695258 379464 695494
rect 379144 688494 379464 695258
rect 379144 688258 379186 688494
rect 379422 688258 379464 688494
rect 379144 681494 379464 688258
rect 379144 681258 379186 681494
rect 379422 681258 379464 681494
rect 379144 674494 379464 681258
rect 379144 674258 379186 674494
rect 379422 674258 379464 674494
rect 379144 667494 379464 674258
rect 379144 667258 379186 667494
rect 379422 667258 379464 667494
rect 379144 660494 379464 667258
rect 379144 660258 379186 660494
rect 379422 660258 379464 660494
rect 379144 653494 379464 660258
rect 379144 653258 379186 653494
rect 379422 653258 379464 653494
rect 379144 646494 379464 653258
rect 379144 646258 379186 646494
rect 379422 646258 379464 646494
rect 379144 639494 379464 646258
rect 379144 639258 379186 639494
rect 379422 639258 379464 639494
rect 379144 632494 379464 639258
rect 379144 632258 379186 632494
rect 379422 632258 379464 632494
rect 379144 625494 379464 632258
rect 379144 625258 379186 625494
rect 379422 625258 379464 625494
rect 379144 618494 379464 625258
rect 379144 618258 379186 618494
rect 379422 618258 379464 618494
rect 379144 611494 379464 618258
rect 379144 611258 379186 611494
rect 379422 611258 379464 611494
rect 379144 604494 379464 611258
rect 379144 604258 379186 604494
rect 379422 604258 379464 604494
rect 379144 597494 379464 604258
rect 379144 597258 379186 597494
rect 379422 597258 379464 597494
rect 379144 590494 379464 597258
rect 379144 590258 379186 590494
rect 379422 590258 379464 590494
rect 379144 583494 379464 590258
rect 379144 583258 379186 583494
rect 379422 583258 379464 583494
rect 379144 576494 379464 583258
rect 379144 576258 379186 576494
rect 379422 576258 379464 576494
rect 379144 569494 379464 576258
rect 379144 569258 379186 569494
rect 379422 569258 379464 569494
rect 379144 562494 379464 569258
rect 379144 562258 379186 562494
rect 379422 562258 379464 562494
rect 379144 555494 379464 562258
rect 379144 555258 379186 555494
rect 379422 555258 379464 555494
rect 379144 548494 379464 555258
rect 379144 548258 379186 548494
rect 379422 548258 379464 548494
rect 379144 541494 379464 548258
rect 379144 541258 379186 541494
rect 379422 541258 379464 541494
rect 379144 534494 379464 541258
rect 379144 534258 379186 534494
rect 379422 534258 379464 534494
rect 379144 527494 379464 534258
rect 379144 527258 379186 527494
rect 379422 527258 379464 527494
rect 379144 520494 379464 527258
rect 379144 520258 379186 520494
rect 379422 520258 379464 520494
rect 379144 513494 379464 520258
rect 379144 513258 379186 513494
rect 379422 513258 379464 513494
rect 379144 506494 379464 513258
rect 379144 506258 379186 506494
rect 379422 506258 379464 506494
rect 379144 499494 379464 506258
rect 379144 499258 379186 499494
rect 379422 499258 379464 499494
rect 379144 492494 379464 499258
rect 379144 492258 379186 492494
rect 379422 492258 379464 492494
rect 379144 485494 379464 492258
rect 379144 485258 379186 485494
rect 379422 485258 379464 485494
rect 379144 478494 379464 485258
rect 379144 478258 379186 478494
rect 379422 478258 379464 478494
rect 379144 471494 379464 478258
rect 379144 471258 379186 471494
rect 379422 471258 379464 471494
rect 379144 464494 379464 471258
rect 379144 464258 379186 464494
rect 379422 464258 379464 464494
rect 379144 457494 379464 464258
rect 379144 457258 379186 457494
rect 379422 457258 379464 457494
rect 379144 450494 379464 457258
rect 379144 450258 379186 450494
rect 379422 450258 379464 450494
rect 379144 443494 379464 450258
rect 379144 443258 379186 443494
rect 379422 443258 379464 443494
rect 379144 436494 379464 443258
rect 379144 436258 379186 436494
rect 379422 436258 379464 436494
rect 379144 429494 379464 436258
rect 379144 429258 379186 429494
rect 379422 429258 379464 429494
rect 379144 422494 379464 429258
rect 379144 422258 379186 422494
rect 379422 422258 379464 422494
rect 379144 415494 379464 422258
rect 379144 415258 379186 415494
rect 379422 415258 379464 415494
rect 379144 408494 379464 415258
rect 379144 408258 379186 408494
rect 379422 408258 379464 408494
rect 379144 401494 379464 408258
rect 379144 401258 379186 401494
rect 379422 401258 379464 401494
rect 379144 394494 379464 401258
rect 379144 394258 379186 394494
rect 379422 394258 379464 394494
rect 379144 387494 379464 394258
rect 379144 387258 379186 387494
rect 379422 387258 379464 387494
rect 379144 380494 379464 387258
rect 379144 380258 379186 380494
rect 379422 380258 379464 380494
rect 379144 373494 379464 380258
rect 379144 373258 379186 373494
rect 379422 373258 379464 373494
rect 379144 366494 379464 373258
rect 379144 366258 379186 366494
rect 379422 366258 379464 366494
rect 379144 359494 379464 366258
rect 379144 359258 379186 359494
rect 379422 359258 379464 359494
rect 379144 352494 379464 359258
rect 379144 352258 379186 352494
rect 379422 352258 379464 352494
rect 379144 345494 379464 352258
rect 379144 345258 379186 345494
rect 379422 345258 379464 345494
rect 379144 338494 379464 345258
rect 379144 338258 379186 338494
rect 379422 338258 379464 338494
rect 379144 331494 379464 338258
rect 379144 331258 379186 331494
rect 379422 331258 379464 331494
rect 379144 324494 379464 331258
rect 379144 324258 379186 324494
rect 379422 324258 379464 324494
rect 379144 317494 379464 324258
rect 379144 317258 379186 317494
rect 379422 317258 379464 317494
rect 379144 310494 379464 317258
rect 379144 310258 379186 310494
rect 379422 310258 379464 310494
rect 379144 303494 379464 310258
rect 379144 303258 379186 303494
rect 379422 303258 379464 303494
rect 379144 296494 379464 303258
rect 379144 296258 379186 296494
rect 379422 296258 379464 296494
rect 379144 289494 379464 296258
rect 379144 289258 379186 289494
rect 379422 289258 379464 289494
rect 379144 282494 379464 289258
rect 379144 282258 379186 282494
rect 379422 282258 379464 282494
rect 379144 275494 379464 282258
rect 379144 275258 379186 275494
rect 379422 275258 379464 275494
rect 379144 268494 379464 275258
rect 379144 268258 379186 268494
rect 379422 268258 379464 268494
rect 379144 261494 379464 268258
rect 379144 261258 379186 261494
rect 379422 261258 379464 261494
rect 379144 254494 379464 261258
rect 379144 254258 379186 254494
rect 379422 254258 379464 254494
rect 379144 247494 379464 254258
rect 379144 247258 379186 247494
rect 379422 247258 379464 247494
rect 379144 240494 379464 247258
rect 379144 240258 379186 240494
rect 379422 240258 379464 240494
rect 379144 233494 379464 240258
rect 379144 233258 379186 233494
rect 379422 233258 379464 233494
rect 379144 226494 379464 233258
rect 379144 226258 379186 226494
rect 379422 226258 379464 226494
rect 379144 219494 379464 226258
rect 379144 219258 379186 219494
rect 379422 219258 379464 219494
rect 379144 212494 379464 219258
rect 379144 212258 379186 212494
rect 379422 212258 379464 212494
rect 379144 205494 379464 212258
rect 379144 205258 379186 205494
rect 379422 205258 379464 205494
rect 379144 198494 379464 205258
rect 379144 198258 379186 198494
rect 379422 198258 379464 198494
rect 379144 191494 379464 198258
rect 379144 191258 379186 191494
rect 379422 191258 379464 191494
rect 379144 184494 379464 191258
rect 379144 184258 379186 184494
rect 379422 184258 379464 184494
rect 379144 177494 379464 184258
rect 379144 177258 379186 177494
rect 379422 177258 379464 177494
rect 379144 170494 379464 177258
rect 379144 170258 379186 170494
rect 379422 170258 379464 170494
rect 379144 163494 379464 170258
rect 379144 163258 379186 163494
rect 379422 163258 379464 163494
rect 379144 156494 379464 163258
rect 379144 156258 379186 156494
rect 379422 156258 379464 156494
rect 379144 149494 379464 156258
rect 379144 149258 379186 149494
rect 379422 149258 379464 149494
rect 379144 142494 379464 149258
rect 379144 142258 379186 142494
rect 379422 142258 379464 142494
rect 379144 135494 379464 142258
rect 379144 135258 379186 135494
rect 379422 135258 379464 135494
rect 379144 128494 379464 135258
rect 379144 128258 379186 128494
rect 379422 128258 379464 128494
rect 379144 121494 379464 128258
rect 379144 121258 379186 121494
rect 379422 121258 379464 121494
rect 379144 114494 379464 121258
rect 379144 114258 379186 114494
rect 379422 114258 379464 114494
rect 379144 107494 379464 114258
rect 379144 107258 379186 107494
rect 379422 107258 379464 107494
rect 379144 100494 379464 107258
rect 379144 100258 379186 100494
rect 379422 100258 379464 100494
rect 379144 93494 379464 100258
rect 379144 93258 379186 93494
rect 379422 93258 379464 93494
rect 379144 86494 379464 93258
rect 379144 86258 379186 86494
rect 379422 86258 379464 86494
rect 379144 79494 379464 86258
rect 379144 79258 379186 79494
rect 379422 79258 379464 79494
rect 379144 72494 379464 79258
rect 379144 72258 379186 72494
rect 379422 72258 379464 72494
rect 379144 65494 379464 72258
rect 379144 65258 379186 65494
rect 379422 65258 379464 65494
rect 379144 58494 379464 65258
rect 379144 58258 379186 58494
rect 379422 58258 379464 58494
rect 379144 51494 379464 58258
rect 379144 51258 379186 51494
rect 379422 51258 379464 51494
rect 379144 44494 379464 51258
rect 379144 44258 379186 44494
rect 379422 44258 379464 44494
rect 379144 37494 379464 44258
rect 379144 37258 379186 37494
rect 379422 37258 379464 37494
rect 379144 30494 379464 37258
rect 379144 30258 379186 30494
rect 379422 30258 379464 30494
rect 379144 23494 379464 30258
rect 379144 23258 379186 23494
rect 379422 23258 379464 23494
rect 379144 16494 379464 23258
rect 379144 16258 379186 16494
rect 379422 16258 379464 16494
rect 379144 9494 379464 16258
rect 379144 9258 379186 9494
rect 379422 9258 379464 9494
rect 379144 2494 379464 9258
rect 379144 2258 379186 2494
rect 379422 2258 379464 2494
rect 379144 -746 379464 2258
rect 379144 -982 379186 -746
rect 379422 -982 379464 -746
rect 379144 -1066 379464 -982
rect 379144 -1302 379186 -1066
rect 379422 -1302 379464 -1066
rect 379144 -2294 379464 -1302
rect 380876 706198 381196 706230
rect 380876 705962 380918 706198
rect 381154 705962 381196 706198
rect 380876 705878 381196 705962
rect 380876 705642 380918 705878
rect 381154 705642 381196 705878
rect 380876 696561 381196 705642
rect 380876 696325 380918 696561
rect 381154 696325 381196 696561
rect 380876 689561 381196 696325
rect 380876 689325 380918 689561
rect 381154 689325 381196 689561
rect 380876 682561 381196 689325
rect 380876 682325 380918 682561
rect 381154 682325 381196 682561
rect 380876 675561 381196 682325
rect 380876 675325 380918 675561
rect 381154 675325 381196 675561
rect 380876 668561 381196 675325
rect 380876 668325 380918 668561
rect 381154 668325 381196 668561
rect 380876 661561 381196 668325
rect 380876 661325 380918 661561
rect 381154 661325 381196 661561
rect 380876 654561 381196 661325
rect 380876 654325 380918 654561
rect 381154 654325 381196 654561
rect 380876 647561 381196 654325
rect 380876 647325 380918 647561
rect 381154 647325 381196 647561
rect 380876 640561 381196 647325
rect 380876 640325 380918 640561
rect 381154 640325 381196 640561
rect 380876 633561 381196 640325
rect 380876 633325 380918 633561
rect 381154 633325 381196 633561
rect 380876 626561 381196 633325
rect 380876 626325 380918 626561
rect 381154 626325 381196 626561
rect 380876 619561 381196 626325
rect 380876 619325 380918 619561
rect 381154 619325 381196 619561
rect 380876 612561 381196 619325
rect 380876 612325 380918 612561
rect 381154 612325 381196 612561
rect 380876 605561 381196 612325
rect 380876 605325 380918 605561
rect 381154 605325 381196 605561
rect 380876 598561 381196 605325
rect 380876 598325 380918 598561
rect 381154 598325 381196 598561
rect 380876 591561 381196 598325
rect 380876 591325 380918 591561
rect 381154 591325 381196 591561
rect 380876 584561 381196 591325
rect 380876 584325 380918 584561
rect 381154 584325 381196 584561
rect 380876 577561 381196 584325
rect 380876 577325 380918 577561
rect 381154 577325 381196 577561
rect 380876 570561 381196 577325
rect 380876 570325 380918 570561
rect 381154 570325 381196 570561
rect 380876 563561 381196 570325
rect 380876 563325 380918 563561
rect 381154 563325 381196 563561
rect 380876 556561 381196 563325
rect 380876 556325 380918 556561
rect 381154 556325 381196 556561
rect 380876 549561 381196 556325
rect 380876 549325 380918 549561
rect 381154 549325 381196 549561
rect 380876 542561 381196 549325
rect 380876 542325 380918 542561
rect 381154 542325 381196 542561
rect 380876 535561 381196 542325
rect 380876 535325 380918 535561
rect 381154 535325 381196 535561
rect 380876 528561 381196 535325
rect 380876 528325 380918 528561
rect 381154 528325 381196 528561
rect 380876 521561 381196 528325
rect 380876 521325 380918 521561
rect 381154 521325 381196 521561
rect 380876 514561 381196 521325
rect 380876 514325 380918 514561
rect 381154 514325 381196 514561
rect 380876 507561 381196 514325
rect 380876 507325 380918 507561
rect 381154 507325 381196 507561
rect 380876 500561 381196 507325
rect 380876 500325 380918 500561
rect 381154 500325 381196 500561
rect 380876 493561 381196 500325
rect 380876 493325 380918 493561
rect 381154 493325 381196 493561
rect 380876 486561 381196 493325
rect 380876 486325 380918 486561
rect 381154 486325 381196 486561
rect 380876 479561 381196 486325
rect 380876 479325 380918 479561
rect 381154 479325 381196 479561
rect 380876 472561 381196 479325
rect 380876 472325 380918 472561
rect 381154 472325 381196 472561
rect 380876 465561 381196 472325
rect 380876 465325 380918 465561
rect 381154 465325 381196 465561
rect 380876 458561 381196 465325
rect 380876 458325 380918 458561
rect 381154 458325 381196 458561
rect 380876 451561 381196 458325
rect 380876 451325 380918 451561
rect 381154 451325 381196 451561
rect 380876 444561 381196 451325
rect 380876 444325 380918 444561
rect 381154 444325 381196 444561
rect 380876 437561 381196 444325
rect 380876 437325 380918 437561
rect 381154 437325 381196 437561
rect 380876 430561 381196 437325
rect 380876 430325 380918 430561
rect 381154 430325 381196 430561
rect 380876 423561 381196 430325
rect 380876 423325 380918 423561
rect 381154 423325 381196 423561
rect 380876 416561 381196 423325
rect 380876 416325 380918 416561
rect 381154 416325 381196 416561
rect 380876 409561 381196 416325
rect 380876 409325 380918 409561
rect 381154 409325 381196 409561
rect 380876 402561 381196 409325
rect 380876 402325 380918 402561
rect 381154 402325 381196 402561
rect 380876 395561 381196 402325
rect 380876 395325 380918 395561
rect 381154 395325 381196 395561
rect 380876 388561 381196 395325
rect 380876 388325 380918 388561
rect 381154 388325 381196 388561
rect 380876 381561 381196 388325
rect 380876 381325 380918 381561
rect 381154 381325 381196 381561
rect 380876 374561 381196 381325
rect 380876 374325 380918 374561
rect 381154 374325 381196 374561
rect 380876 367561 381196 374325
rect 380876 367325 380918 367561
rect 381154 367325 381196 367561
rect 380876 360561 381196 367325
rect 380876 360325 380918 360561
rect 381154 360325 381196 360561
rect 380876 353561 381196 360325
rect 380876 353325 380918 353561
rect 381154 353325 381196 353561
rect 380876 346561 381196 353325
rect 380876 346325 380918 346561
rect 381154 346325 381196 346561
rect 380876 339561 381196 346325
rect 380876 339325 380918 339561
rect 381154 339325 381196 339561
rect 380876 332561 381196 339325
rect 380876 332325 380918 332561
rect 381154 332325 381196 332561
rect 380876 325561 381196 332325
rect 380876 325325 380918 325561
rect 381154 325325 381196 325561
rect 380876 318561 381196 325325
rect 380876 318325 380918 318561
rect 381154 318325 381196 318561
rect 380876 311561 381196 318325
rect 380876 311325 380918 311561
rect 381154 311325 381196 311561
rect 380876 304561 381196 311325
rect 380876 304325 380918 304561
rect 381154 304325 381196 304561
rect 380876 297561 381196 304325
rect 380876 297325 380918 297561
rect 381154 297325 381196 297561
rect 380876 290561 381196 297325
rect 380876 290325 380918 290561
rect 381154 290325 381196 290561
rect 380876 283561 381196 290325
rect 380876 283325 380918 283561
rect 381154 283325 381196 283561
rect 380876 276561 381196 283325
rect 380876 276325 380918 276561
rect 381154 276325 381196 276561
rect 380876 269561 381196 276325
rect 380876 269325 380918 269561
rect 381154 269325 381196 269561
rect 380876 262561 381196 269325
rect 380876 262325 380918 262561
rect 381154 262325 381196 262561
rect 380876 255561 381196 262325
rect 380876 255325 380918 255561
rect 381154 255325 381196 255561
rect 380876 248561 381196 255325
rect 380876 248325 380918 248561
rect 381154 248325 381196 248561
rect 380876 241561 381196 248325
rect 380876 241325 380918 241561
rect 381154 241325 381196 241561
rect 380876 234561 381196 241325
rect 380876 234325 380918 234561
rect 381154 234325 381196 234561
rect 380876 227561 381196 234325
rect 380876 227325 380918 227561
rect 381154 227325 381196 227561
rect 380876 220561 381196 227325
rect 380876 220325 380918 220561
rect 381154 220325 381196 220561
rect 380876 213561 381196 220325
rect 380876 213325 380918 213561
rect 381154 213325 381196 213561
rect 380876 206561 381196 213325
rect 380876 206325 380918 206561
rect 381154 206325 381196 206561
rect 380876 199561 381196 206325
rect 380876 199325 380918 199561
rect 381154 199325 381196 199561
rect 380876 192561 381196 199325
rect 380876 192325 380918 192561
rect 381154 192325 381196 192561
rect 380876 185561 381196 192325
rect 380876 185325 380918 185561
rect 381154 185325 381196 185561
rect 380876 178561 381196 185325
rect 380876 178325 380918 178561
rect 381154 178325 381196 178561
rect 380876 171561 381196 178325
rect 380876 171325 380918 171561
rect 381154 171325 381196 171561
rect 380876 164561 381196 171325
rect 380876 164325 380918 164561
rect 381154 164325 381196 164561
rect 380876 157561 381196 164325
rect 380876 157325 380918 157561
rect 381154 157325 381196 157561
rect 380876 150561 381196 157325
rect 380876 150325 380918 150561
rect 381154 150325 381196 150561
rect 380876 143561 381196 150325
rect 380876 143325 380918 143561
rect 381154 143325 381196 143561
rect 380876 136561 381196 143325
rect 380876 136325 380918 136561
rect 381154 136325 381196 136561
rect 380876 129561 381196 136325
rect 380876 129325 380918 129561
rect 381154 129325 381196 129561
rect 380876 122561 381196 129325
rect 380876 122325 380918 122561
rect 381154 122325 381196 122561
rect 380876 115561 381196 122325
rect 380876 115325 380918 115561
rect 381154 115325 381196 115561
rect 380876 108561 381196 115325
rect 380876 108325 380918 108561
rect 381154 108325 381196 108561
rect 380876 101561 381196 108325
rect 380876 101325 380918 101561
rect 381154 101325 381196 101561
rect 380876 94561 381196 101325
rect 380876 94325 380918 94561
rect 381154 94325 381196 94561
rect 380876 87561 381196 94325
rect 380876 87325 380918 87561
rect 381154 87325 381196 87561
rect 380876 80561 381196 87325
rect 380876 80325 380918 80561
rect 381154 80325 381196 80561
rect 380876 73561 381196 80325
rect 380876 73325 380918 73561
rect 381154 73325 381196 73561
rect 380876 66561 381196 73325
rect 380876 66325 380918 66561
rect 381154 66325 381196 66561
rect 380876 59561 381196 66325
rect 380876 59325 380918 59561
rect 381154 59325 381196 59561
rect 380876 52561 381196 59325
rect 380876 52325 380918 52561
rect 381154 52325 381196 52561
rect 380876 45561 381196 52325
rect 380876 45325 380918 45561
rect 381154 45325 381196 45561
rect 380876 38561 381196 45325
rect 380876 38325 380918 38561
rect 381154 38325 381196 38561
rect 380876 31561 381196 38325
rect 380876 31325 380918 31561
rect 381154 31325 381196 31561
rect 380876 24561 381196 31325
rect 380876 24325 380918 24561
rect 381154 24325 381196 24561
rect 380876 17561 381196 24325
rect 380876 17325 380918 17561
rect 381154 17325 381196 17561
rect 380876 10561 381196 17325
rect 380876 10325 380918 10561
rect 381154 10325 381196 10561
rect 380876 3561 381196 10325
rect 380876 3325 380918 3561
rect 381154 3325 381196 3561
rect 380876 -1706 381196 3325
rect 380876 -1942 380918 -1706
rect 381154 -1942 381196 -1706
rect 380876 -2026 381196 -1942
rect 380876 -2262 380918 -2026
rect 381154 -2262 381196 -2026
rect 380876 -2294 381196 -2262
rect 386144 705238 386464 706230
rect 386144 705002 386186 705238
rect 386422 705002 386464 705238
rect 386144 704918 386464 705002
rect 386144 704682 386186 704918
rect 386422 704682 386464 704918
rect 386144 695494 386464 704682
rect 386144 695258 386186 695494
rect 386422 695258 386464 695494
rect 386144 688494 386464 695258
rect 386144 688258 386186 688494
rect 386422 688258 386464 688494
rect 386144 681494 386464 688258
rect 386144 681258 386186 681494
rect 386422 681258 386464 681494
rect 386144 674494 386464 681258
rect 386144 674258 386186 674494
rect 386422 674258 386464 674494
rect 386144 667494 386464 674258
rect 386144 667258 386186 667494
rect 386422 667258 386464 667494
rect 386144 660494 386464 667258
rect 386144 660258 386186 660494
rect 386422 660258 386464 660494
rect 386144 653494 386464 660258
rect 386144 653258 386186 653494
rect 386422 653258 386464 653494
rect 386144 646494 386464 653258
rect 386144 646258 386186 646494
rect 386422 646258 386464 646494
rect 386144 639494 386464 646258
rect 386144 639258 386186 639494
rect 386422 639258 386464 639494
rect 386144 632494 386464 639258
rect 386144 632258 386186 632494
rect 386422 632258 386464 632494
rect 386144 625494 386464 632258
rect 386144 625258 386186 625494
rect 386422 625258 386464 625494
rect 386144 618494 386464 625258
rect 386144 618258 386186 618494
rect 386422 618258 386464 618494
rect 386144 611494 386464 618258
rect 386144 611258 386186 611494
rect 386422 611258 386464 611494
rect 386144 604494 386464 611258
rect 386144 604258 386186 604494
rect 386422 604258 386464 604494
rect 386144 597494 386464 604258
rect 386144 597258 386186 597494
rect 386422 597258 386464 597494
rect 386144 590494 386464 597258
rect 386144 590258 386186 590494
rect 386422 590258 386464 590494
rect 386144 583494 386464 590258
rect 386144 583258 386186 583494
rect 386422 583258 386464 583494
rect 386144 576494 386464 583258
rect 386144 576258 386186 576494
rect 386422 576258 386464 576494
rect 386144 569494 386464 576258
rect 386144 569258 386186 569494
rect 386422 569258 386464 569494
rect 386144 562494 386464 569258
rect 386144 562258 386186 562494
rect 386422 562258 386464 562494
rect 386144 555494 386464 562258
rect 386144 555258 386186 555494
rect 386422 555258 386464 555494
rect 386144 548494 386464 555258
rect 386144 548258 386186 548494
rect 386422 548258 386464 548494
rect 386144 541494 386464 548258
rect 386144 541258 386186 541494
rect 386422 541258 386464 541494
rect 386144 534494 386464 541258
rect 386144 534258 386186 534494
rect 386422 534258 386464 534494
rect 386144 527494 386464 534258
rect 386144 527258 386186 527494
rect 386422 527258 386464 527494
rect 386144 520494 386464 527258
rect 386144 520258 386186 520494
rect 386422 520258 386464 520494
rect 386144 513494 386464 520258
rect 386144 513258 386186 513494
rect 386422 513258 386464 513494
rect 386144 506494 386464 513258
rect 386144 506258 386186 506494
rect 386422 506258 386464 506494
rect 386144 499494 386464 506258
rect 386144 499258 386186 499494
rect 386422 499258 386464 499494
rect 386144 492494 386464 499258
rect 386144 492258 386186 492494
rect 386422 492258 386464 492494
rect 386144 485494 386464 492258
rect 386144 485258 386186 485494
rect 386422 485258 386464 485494
rect 386144 478494 386464 485258
rect 386144 478258 386186 478494
rect 386422 478258 386464 478494
rect 386144 471494 386464 478258
rect 386144 471258 386186 471494
rect 386422 471258 386464 471494
rect 386144 464494 386464 471258
rect 386144 464258 386186 464494
rect 386422 464258 386464 464494
rect 386144 457494 386464 464258
rect 386144 457258 386186 457494
rect 386422 457258 386464 457494
rect 386144 450494 386464 457258
rect 386144 450258 386186 450494
rect 386422 450258 386464 450494
rect 386144 443494 386464 450258
rect 386144 443258 386186 443494
rect 386422 443258 386464 443494
rect 386144 436494 386464 443258
rect 386144 436258 386186 436494
rect 386422 436258 386464 436494
rect 386144 429494 386464 436258
rect 386144 429258 386186 429494
rect 386422 429258 386464 429494
rect 386144 422494 386464 429258
rect 386144 422258 386186 422494
rect 386422 422258 386464 422494
rect 386144 415494 386464 422258
rect 386144 415258 386186 415494
rect 386422 415258 386464 415494
rect 386144 408494 386464 415258
rect 386144 408258 386186 408494
rect 386422 408258 386464 408494
rect 386144 401494 386464 408258
rect 386144 401258 386186 401494
rect 386422 401258 386464 401494
rect 386144 394494 386464 401258
rect 386144 394258 386186 394494
rect 386422 394258 386464 394494
rect 386144 387494 386464 394258
rect 386144 387258 386186 387494
rect 386422 387258 386464 387494
rect 386144 380494 386464 387258
rect 386144 380258 386186 380494
rect 386422 380258 386464 380494
rect 386144 373494 386464 380258
rect 386144 373258 386186 373494
rect 386422 373258 386464 373494
rect 386144 366494 386464 373258
rect 386144 366258 386186 366494
rect 386422 366258 386464 366494
rect 386144 359494 386464 366258
rect 386144 359258 386186 359494
rect 386422 359258 386464 359494
rect 386144 352494 386464 359258
rect 386144 352258 386186 352494
rect 386422 352258 386464 352494
rect 386144 345494 386464 352258
rect 386144 345258 386186 345494
rect 386422 345258 386464 345494
rect 386144 338494 386464 345258
rect 386144 338258 386186 338494
rect 386422 338258 386464 338494
rect 386144 331494 386464 338258
rect 386144 331258 386186 331494
rect 386422 331258 386464 331494
rect 386144 324494 386464 331258
rect 386144 324258 386186 324494
rect 386422 324258 386464 324494
rect 386144 317494 386464 324258
rect 386144 317258 386186 317494
rect 386422 317258 386464 317494
rect 386144 310494 386464 317258
rect 386144 310258 386186 310494
rect 386422 310258 386464 310494
rect 386144 303494 386464 310258
rect 386144 303258 386186 303494
rect 386422 303258 386464 303494
rect 386144 296494 386464 303258
rect 386144 296258 386186 296494
rect 386422 296258 386464 296494
rect 386144 289494 386464 296258
rect 386144 289258 386186 289494
rect 386422 289258 386464 289494
rect 386144 282494 386464 289258
rect 386144 282258 386186 282494
rect 386422 282258 386464 282494
rect 386144 275494 386464 282258
rect 386144 275258 386186 275494
rect 386422 275258 386464 275494
rect 386144 268494 386464 275258
rect 386144 268258 386186 268494
rect 386422 268258 386464 268494
rect 386144 261494 386464 268258
rect 386144 261258 386186 261494
rect 386422 261258 386464 261494
rect 386144 254494 386464 261258
rect 386144 254258 386186 254494
rect 386422 254258 386464 254494
rect 386144 247494 386464 254258
rect 386144 247258 386186 247494
rect 386422 247258 386464 247494
rect 386144 240494 386464 247258
rect 386144 240258 386186 240494
rect 386422 240258 386464 240494
rect 386144 233494 386464 240258
rect 386144 233258 386186 233494
rect 386422 233258 386464 233494
rect 386144 226494 386464 233258
rect 386144 226258 386186 226494
rect 386422 226258 386464 226494
rect 386144 219494 386464 226258
rect 386144 219258 386186 219494
rect 386422 219258 386464 219494
rect 386144 212494 386464 219258
rect 386144 212258 386186 212494
rect 386422 212258 386464 212494
rect 386144 205494 386464 212258
rect 386144 205258 386186 205494
rect 386422 205258 386464 205494
rect 386144 198494 386464 205258
rect 386144 198258 386186 198494
rect 386422 198258 386464 198494
rect 386144 191494 386464 198258
rect 386144 191258 386186 191494
rect 386422 191258 386464 191494
rect 386144 184494 386464 191258
rect 386144 184258 386186 184494
rect 386422 184258 386464 184494
rect 386144 177494 386464 184258
rect 386144 177258 386186 177494
rect 386422 177258 386464 177494
rect 386144 170494 386464 177258
rect 386144 170258 386186 170494
rect 386422 170258 386464 170494
rect 386144 163494 386464 170258
rect 386144 163258 386186 163494
rect 386422 163258 386464 163494
rect 386144 156494 386464 163258
rect 386144 156258 386186 156494
rect 386422 156258 386464 156494
rect 386144 149494 386464 156258
rect 386144 149258 386186 149494
rect 386422 149258 386464 149494
rect 386144 142494 386464 149258
rect 386144 142258 386186 142494
rect 386422 142258 386464 142494
rect 386144 135494 386464 142258
rect 386144 135258 386186 135494
rect 386422 135258 386464 135494
rect 386144 128494 386464 135258
rect 386144 128258 386186 128494
rect 386422 128258 386464 128494
rect 386144 121494 386464 128258
rect 386144 121258 386186 121494
rect 386422 121258 386464 121494
rect 386144 114494 386464 121258
rect 386144 114258 386186 114494
rect 386422 114258 386464 114494
rect 386144 107494 386464 114258
rect 386144 107258 386186 107494
rect 386422 107258 386464 107494
rect 386144 100494 386464 107258
rect 386144 100258 386186 100494
rect 386422 100258 386464 100494
rect 386144 93494 386464 100258
rect 386144 93258 386186 93494
rect 386422 93258 386464 93494
rect 386144 86494 386464 93258
rect 386144 86258 386186 86494
rect 386422 86258 386464 86494
rect 386144 79494 386464 86258
rect 386144 79258 386186 79494
rect 386422 79258 386464 79494
rect 386144 72494 386464 79258
rect 386144 72258 386186 72494
rect 386422 72258 386464 72494
rect 386144 65494 386464 72258
rect 386144 65258 386186 65494
rect 386422 65258 386464 65494
rect 386144 58494 386464 65258
rect 386144 58258 386186 58494
rect 386422 58258 386464 58494
rect 386144 51494 386464 58258
rect 386144 51258 386186 51494
rect 386422 51258 386464 51494
rect 386144 44494 386464 51258
rect 386144 44258 386186 44494
rect 386422 44258 386464 44494
rect 386144 37494 386464 44258
rect 386144 37258 386186 37494
rect 386422 37258 386464 37494
rect 386144 30494 386464 37258
rect 386144 30258 386186 30494
rect 386422 30258 386464 30494
rect 386144 23494 386464 30258
rect 386144 23258 386186 23494
rect 386422 23258 386464 23494
rect 386144 16494 386464 23258
rect 386144 16258 386186 16494
rect 386422 16258 386464 16494
rect 386144 9494 386464 16258
rect 386144 9258 386186 9494
rect 386422 9258 386464 9494
rect 386144 2494 386464 9258
rect 386144 2258 386186 2494
rect 386422 2258 386464 2494
rect 386144 -746 386464 2258
rect 386144 -982 386186 -746
rect 386422 -982 386464 -746
rect 386144 -1066 386464 -982
rect 386144 -1302 386186 -1066
rect 386422 -1302 386464 -1066
rect 386144 -2294 386464 -1302
rect 387876 706198 388196 706230
rect 387876 705962 387918 706198
rect 388154 705962 388196 706198
rect 387876 705878 388196 705962
rect 387876 705642 387918 705878
rect 388154 705642 388196 705878
rect 387876 696561 388196 705642
rect 387876 696325 387918 696561
rect 388154 696325 388196 696561
rect 387876 689561 388196 696325
rect 387876 689325 387918 689561
rect 388154 689325 388196 689561
rect 387876 682561 388196 689325
rect 387876 682325 387918 682561
rect 388154 682325 388196 682561
rect 387876 675561 388196 682325
rect 387876 675325 387918 675561
rect 388154 675325 388196 675561
rect 387876 668561 388196 675325
rect 387876 668325 387918 668561
rect 388154 668325 388196 668561
rect 387876 661561 388196 668325
rect 387876 661325 387918 661561
rect 388154 661325 388196 661561
rect 387876 654561 388196 661325
rect 387876 654325 387918 654561
rect 388154 654325 388196 654561
rect 387876 647561 388196 654325
rect 387876 647325 387918 647561
rect 388154 647325 388196 647561
rect 387876 640561 388196 647325
rect 387876 640325 387918 640561
rect 388154 640325 388196 640561
rect 387876 633561 388196 640325
rect 387876 633325 387918 633561
rect 388154 633325 388196 633561
rect 387876 626561 388196 633325
rect 387876 626325 387918 626561
rect 388154 626325 388196 626561
rect 387876 619561 388196 626325
rect 387876 619325 387918 619561
rect 388154 619325 388196 619561
rect 387876 612561 388196 619325
rect 387876 612325 387918 612561
rect 388154 612325 388196 612561
rect 387876 605561 388196 612325
rect 387876 605325 387918 605561
rect 388154 605325 388196 605561
rect 387876 598561 388196 605325
rect 387876 598325 387918 598561
rect 388154 598325 388196 598561
rect 387876 591561 388196 598325
rect 387876 591325 387918 591561
rect 388154 591325 388196 591561
rect 387876 584561 388196 591325
rect 387876 584325 387918 584561
rect 388154 584325 388196 584561
rect 387876 577561 388196 584325
rect 387876 577325 387918 577561
rect 388154 577325 388196 577561
rect 387876 570561 388196 577325
rect 387876 570325 387918 570561
rect 388154 570325 388196 570561
rect 387876 563561 388196 570325
rect 387876 563325 387918 563561
rect 388154 563325 388196 563561
rect 387876 556561 388196 563325
rect 387876 556325 387918 556561
rect 388154 556325 388196 556561
rect 387876 549561 388196 556325
rect 387876 549325 387918 549561
rect 388154 549325 388196 549561
rect 387876 542561 388196 549325
rect 387876 542325 387918 542561
rect 388154 542325 388196 542561
rect 387876 535561 388196 542325
rect 387876 535325 387918 535561
rect 388154 535325 388196 535561
rect 387876 528561 388196 535325
rect 387876 528325 387918 528561
rect 388154 528325 388196 528561
rect 387876 521561 388196 528325
rect 387876 521325 387918 521561
rect 388154 521325 388196 521561
rect 387876 514561 388196 521325
rect 387876 514325 387918 514561
rect 388154 514325 388196 514561
rect 387876 507561 388196 514325
rect 387876 507325 387918 507561
rect 388154 507325 388196 507561
rect 387876 500561 388196 507325
rect 387876 500325 387918 500561
rect 388154 500325 388196 500561
rect 387876 493561 388196 500325
rect 387876 493325 387918 493561
rect 388154 493325 388196 493561
rect 387876 486561 388196 493325
rect 387876 486325 387918 486561
rect 388154 486325 388196 486561
rect 387876 479561 388196 486325
rect 387876 479325 387918 479561
rect 388154 479325 388196 479561
rect 387876 472561 388196 479325
rect 387876 472325 387918 472561
rect 388154 472325 388196 472561
rect 387876 465561 388196 472325
rect 387876 465325 387918 465561
rect 388154 465325 388196 465561
rect 387876 458561 388196 465325
rect 387876 458325 387918 458561
rect 388154 458325 388196 458561
rect 387876 451561 388196 458325
rect 387876 451325 387918 451561
rect 388154 451325 388196 451561
rect 387876 444561 388196 451325
rect 387876 444325 387918 444561
rect 388154 444325 388196 444561
rect 387876 437561 388196 444325
rect 387876 437325 387918 437561
rect 388154 437325 388196 437561
rect 387876 430561 388196 437325
rect 387876 430325 387918 430561
rect 388154 430325 388196 430561
rect 387876 423561 388196 430325
rect 387876 423325 387918 423561
rect 388154 423325 388196 423561
rect 387876 416561 388196 423325
rect 387876 416325 387918 416561
rect 388154 416325 388196 416561
rect 387876 409561 388196 416325
rect 387876 409325 387918 409561
rect 388154 409325 388196 409561
rect 387876 402561 388196 409325
rect 387876 402325 387918 402561
rect 388154 402325 388196 402561
rect 387876 395561 388196 402325
rect 387876 395325 387918 395561
rect 388154 395325 388196 395561
rect 387876 388561 388196 395325
rect 387876 388325 387918 388561
rect 388154 388325 388196 388561
rect 387876 381561 388196 388325
rect 387876 381325 387918 381561
rect 388154 381325 388196 381561
rect 387876 374561 388196 381325
rect 387876 374325 387918 374561
rect 388154 374325 388196 374561
rect 387876 367561 388196 374325
rect 387876 367325 387918 367561
rect 388154 367325 388196 367561
rect 387876 360561 388196 367325
rect 387876 360325 387918 360561
rect 388154 360325 388196 360561
rect 387876 353561 388196 360325
rect 387876 353325 387918 353561
rect 388154 353325 388196 353561
rect 387876 346561 388196 353325
rect 387876 346325 387918 346561
rect 388154 346325 388196 346561
rect 387876 339561 388196 346325
rect 387876 339325 387918 339561
rect 388154 339325 388196 339561
rect 387876 332561 388196 339325
rect 387876 332325 387918 332561
rect 388154 332325 388196 332561
rect 387876 325561 388196 332325
rect 387876 325325 387918 325561
rect 388154 325325 388196 325561
rect 387876 318561 388196 325325
rect 387876 318325 387918 318561
rect 388154 318325 388196 318561
rect 387876 311561 388196 318325
rect 387876 311325 387918 311561
rect 388154 311325 388196 311561
rect 387876 304561 388196 311325
rect 387876 304325 387918 304561
rect 388154 304325 388196 304561
rect 387876 297561 388196 304325
rect 387876 297325 387918 297561
rect 388154 297325 388196 297561
rect 387876 290561 388196 297325
rect 387876 290325 387918 290561
rect 388154 290325 388196 290561
rect 387876 283561 388196 290325
rect 387876 283325 387918 283561
rect 388154 283325 388196 283561
rect 387876 276561 388196 283325
rect 387876 276325 387918 276561
rect 388154 276325 388196 276561
rect 387876 269561 388196 276325
rect 387876 269325 387918 269561
rect 388154 269325 388196 269561
rect 387876 262561 388196 269325
rect 387876 262325 387918 262561
rect 388154 262325 388196 262561
rect 387876 255561 388196 262325
rect 387876 255325 387918 255561
rect 388154 255325 388196 255561
rect 387876 248561 388196 255325
rect 387876 248325 387918 248561
rect 388154 248325 388196 248561
rect 387876 241561 388196 248325
rect 387876 241325 387918 241561
rect 388154 241325 388196 241561
rect 387876 234561 388196 241325
rect 387876 234325 387918 234561
rect 388154 234325 388196 234561
rect 387876 227561 388196 234325
rect 387876 227325 387918 227561
rect 388154 227325 388196 227561
rect 387876 220561 388196 227325
rect 387876 220325 387918 220561
rect 388154 220325 388196 220561
rect 387876 213561 388196 220325
rect 387876 213325 387918 213561
rect 388154 213325 388196 213561
rect 387876 206561 388196 213325
rect 387876 206325 387918 206561
rect 388154 206325 388196 206561
rect 387876 199561 388196 206325
rect 387876 199325 387918 199561
rect 388154 199325 388196 199561
rect 387876 192561 388196 199325
rect 387876 192325 387918 192561
rect 388154 192325 388196 192561
rect 387876 185561 388196 192325
rect 387876 185325 387918 185561
rect 388154 185325 388196 185561
rect 387876 178561 388196 185325
rect 387876 178325 387918 178561
rect 388154 178325 388196 178561
rect 387876 171561 388196 178325
rect 387876 171325 387918 171561
rect 388154 171325 388196 171561
rect 387876 164561 388196 171325
rect 387876 164325 387918 164561
rect 388154 164325 388196 164561
rect 387876 157561 388196 164325
rect 387876 157325 387918 157561
rect 388154 157325 388196 157561
rect 387876 150561 388196 157325
rect 387876 150325 387918 150561
rect 388154 150325 388196 150561
rect 387876 143561 388196 150325
rect 387876 143325 387918 143561
rect 388154 143325 388196 143561
rect 387876 136561 388196 143325
rect 387876 136325 387918 136561
rect 388154 136325 388196 136561
rect 387876 129561 388196 136325
rect 387876 129325 387918 129561
rect 388154 129325 388196 129561
rect 387876 122561 388196 129325
rect 387876 122325 387918 122561
rect 388154 122325 388196 122561
rect 387876 115561 388196 122325
rect 387876 115325 387918 115561
rect 388154 115325 388196 115561
rect 387876 108561 388196 115325
rect 387876 108325 387918 108561
rect 388154 108325 388196 108561
rect 387876 101561 388196 108325
rect 387876 101325 387918 101561
rect 388154 101325 388196 101561
rect 387876 94561 388196 101325
rect 387876 94325 387918 94561
rect 388154 94325 388196 94561
rect 387876 87561 388196 94325
rect 387876 87325 387918 87561
rect 388154 87325 388196 87561
rect 387876 80561 388196 87325
rect 387876 80325 387918 80561
rect 388154 80325 388196 80561
rect 387876 73561 388196 80325
rect 387876 73325 387918 73561
rect 388154 73325 388196 73561
rect 387876 66561 388196 73325
rect 387876 66325 387918 66561
rect 388154 66325 388196 66561
rect 387876 59561 388196 66325
rect 387876 59325 387918 59561
rect 388154 59325 388196 59561
rect 387876 52561 388196 59325
rect 387876 52325 387918 52561
rect 388154 52325 388196 52561
rect 387876 45561 388196 52325
rect 387876 45325 387918 45561
rect 388154 45325 388196 45561
rect 387876 38561 388196 45325
rect 387876 38325 387918 38561
rect 388154 38325 388196 38561
rect 387876 31561 388196 38325
rect 387876 31325 387918 31561
rect 388154 31325 388196 31561
rect 387876 24561 388196 31325
rect 387876 24325 387918 24561
rect 388154 24325 388196 24561
rect 387876 17561 388196 24325
rect 387876 17325 387918 17561
rect 388154 17325 388196 17561
rect 387876 10561 388196 17325
rect 387876 10325 387918 10561
rect 388154 10325 388196 10561
rect 387876 3561 388196 10325
rect 387876 3325 387918 3561
rect 388154 3325 388196 3561
rect 387876 -1706 388196 3325
rect 387876 -1942 387918 -1706
rect 388154 -1942 388196 -1706
rect 387876 -2026 388196 -1942
rect 387876 -2262 387918 -2026
rect 388154 -2262 388196 -2026
rect 387876 -2294 388196 -2262
rect 393144 705238 393464 706230
rect 393144 705002 393186 705238
rect 393422 705002 393464 705238
rect 393144 704918 393464 705002
rect 393144 704682 393186 704918
rect 393422 704682 393464 704918
rect 393144 695494 393464 704682
rect 393144 695258 393186 695494
rect 393422 695258 393464 695494
rect 393144 688494 393464 695258
rect 393144 688258 393186 688494
rect 393422 688258 393464 688494
rect 393144 681494 393464 688258
rect 393144 681258 393186 681494
rect 393422 681258 393464 681494
rect 393144 674494 393464 681258
rect 393144 674258 393186 674494
rect 393422 674258 393464 674494
rect 393144 667494 393464 674258
rect 393144 667258 393186 667494
rect 393422 667258 393464 667494
rect 393144 660494 393464 667258
rect 393144 660258 393186 660494
rect 393422 660258 393464 660494
rect 393144 653494 393464 660258
rect 393144 653258 393186 653494
rect 393422 653258 393464 653494
rect 393144 646494 393464 653258
rect 393144 646258 393186 646494
rect 393422 646258 393464 646494
rect 393144 639494 393464 646258
rect 393144 639258 393186 639494
rect 393422 639258 393464 639494
rect 393144 632494 393464 639258
rect 393144 632258 393186 632494
rect 393422 632258 393464 632494
rect 393144 625494 393464 632258
rect 393144 625258 393186 625494
rect 393422 625258 393464 625494
rect 393144 618494 393464 625258
rect 393144 618258 393186 618494
rect 393422 618258 393464 618494
rect 393144 611494 393464 618258
rect 393144 611258 393186 611494
rect 393422 611258 393464 611494
rect 393144 604494 393464 611258
rect 393144 604258 393186 604494
rect 393422 604258 393464 604494
rect 393144 597494 393464 604258
rect 393144 597258 393186 597494
rect 393422 597258 393464 597494
rect 393144 590494 393464 597258
rect 393144 590258 393186 590494
rect 393422 590258 393464 590494
rect 393144 583494 393464 590258
rect 393144 583258 393186 583494
rect 393422 583258 393464 583494
rect 393144 576494 393464 583258
rect 393144 576258 393186 576494
rect 393422 576258 393464 576494
rect 393144 569494 393464 576258
rect 393144 569258 393186 569494
rect 393422 569258 393464 569494
rect 393144 562494 393464 569258
rect 393144 562258 393186 562494
rect 393422 562258 393464 562494
rect 393144 555494 393464 562258
rect 393144 555258 393186 555494
rect 393422 555258 393464 555494
rect 393144 548494 393464 555258
rect 393144 548258 393186 548494
rect 393422 548258 393464 548494
rect 393144 541494 393464 548258
rect 393144 541258 393186 541494
rect 393422 541258 393464 541494
rect 393144 534494 393464 541258
rect 393144 534258 393186 534494
rect 393422 534258 393464 534494
rect 393144 527494 393464 534258
rect 393144 527258 393186 527494
rect 393422 527258 393464 527494
rect 393144 520494 393464 527258
rect 393144 520258 393186 520494
rect 393422 520258 393464 520494
rect 393144 513494 393464 520258
rect 393144 513258 393186 513494
rect 393422 513258 393464 513494
rect 393144 506494 393464 513258
rect 393144 506258 393186 506494
rect 393422 506258 393464 506494
rect 393144 499494 393464 506258
rect 393144 499258 393186 499494
rect 393422 499258 393464 499494
rect 393144 492494 393464 499258
rect 393144 492258 393186 492494
rect 393422 492258 393464 492494
rect 393144 485494 393464 492258
rect 393144 485258 393186 485494
rect 393422 485258 393464 485494
rect 393144 478494 393464 485258
rect 393144 478258 393186 478494
rect 393422 478258 393464 478494
rect 393144 471494 393464 478258
rect 393144 471258 393186 471494
rect 393422 471258 393464 471494
rect 393144 464494 393464 471258
rect 393144 464258 393186 464494
rect 393422 464258 393464 464494
rect 393144 457494 393464 464258
rect 393144 457258 393186 457494
rect 393422 457258 393464 457494
rect 393144 450494 393464 457258
rect 393144 450258 393186 450494
rect 393422 450258 393464 450494
rect 393144 443494 393464 450258
rect 393144 443258 393186 443494
rect 393422 443258 393464 443494
rect 393144 436494 393464 443258
rect 393144 436258 393186 436494
rect 393422 436258 393464 436494
rect 393144 429494 393464 436258
rect 393144 429258 393186 429494
rect 393422 429258 393464 429494
rect 393144 422494 393464 429258
rect 393144 422258 393186 422494
rect 393422 422258 393464 422494
rect 393144 415494 393464 422258
rect 393144 415258 393186 415494
rect 393422 415258 393464 415494
rect 393144 408494 393464 415258
rect 393144 408258 393186 408494
rect 393422 408258 393464 408494
rect 393144 401494 393464 408258
rect 393144 401258 393186 401494
rect 393422 401258 393464 401494
rect 393144 394494 393464 401258
rect 393144 394258 393186 394494
rect 393422 394258 393464 394494
rect 393144 387494 393464 394258
rect 393144 387258 393186 387494
rect 393422 387258 393464 387494
rect 393144 380494 393464 387258
rect 393144 380258 393186 380494
rect 393422 380258 393464 380494
rect 393144 373494 393464 380258
rect 393144 373258 393186 373494
rect 393422 373258 393464 373494
rect 393144 366494 393464 373258
rect 393144 366258 393186 366494
rect 393422 366258 393464 366494
rect 393144 359494 393464 366258
rect 393144 359258 393186 359494
rect 393422 359258 393464 359494
rect 393144 352494 393464 359258
rect 393144 352258 393186 352494
rect 393422 352258 393464 352494
rect 393144 345494 393464 352258
rect 393144 345258 393186 345494
rect 393422 345258 393464 345494
rect 393144 338494 393464 345258
rect 393144 338258 393186 338494
rect 393422 338258 393464 338494
rect 393144 331494 393464 338258
rect 393144 331258 393186 331494
rect 393422 331258 393464 331494
rect 393144 324494 393464 331258
rect 393144 324258 393186 324494
rect 393422 324258 393464 324494
rect 393144 317494 393464 324258
rect 393144 317258 393186 317494
rect 393422 317258 393464 317494
rect 393144 310494 393464 317258
rect 393144 310258 393186 310494
rect 393422 310258 393464 310494
rect 393144 303494 393464 310258
rect 393144 303258 393186 303494
rect 393422 303258 393464 303494
rect 393144 296494 393464 303258
rect 393144 296258 393186 296494
rect 393422 296258 393464 296494
rect 393144 289494 393464 296258
rect 393144 289258 393186 289494
rect 393422 289258 393464 289494
rect 393144 282494 393464 289258
rect 393144 282258 393186 282494
rect 393422 282258 393464 282494
rect 393144 275494 393464 282258
rect 393144 275258 393186 275494
rect 393422 275258 393464 275494
rect 393144 268494 393464 275258
rect 393144 268258 393186 268494
rect 393422 268258 393464 268494
rect 393144 261494 393464 268258
rect 393144 261258 393186 261494
rect 393422 261258 393464 261494
rect 393144 254494 393464 261258
rect 393144 254258 393186 254494
rect 393422 254258 393464 254494
rect 393144 247494 393464 254258
rect 393144 247258 393186 247494
rect 393422 247258 393464 247494
rect 393144 240494 393464 247258
rect 393144 240258 393186 240494
rect 393422 240258 393464 240494
rect 393144 233494 393464 240258
rect 393144 233258 393186 233494
rect 393422 233258 393464 233494
rect 393144 226494 393464 233258
rect 393144 226258 393186 226494
rect 393422 226258 393464 226494
rect 393144 219494 393464 226258
rect 393144 219258 393186 219494
rect 393422 219258 393464 219494
rect 393144 212494 393464 219258
rect 393144 212258 393186 212494
rect 393422 212258 393464 212494
rect 393144 205494 393464 212258
rect 393144 205258 393186 205494
rect 393422 205258 393464 205494
rect 393144 198494 393464 205258
rect 393144 198258 393186 198494
rect 393422 198258 393464 198494
rect 393144 191494 393464 198258
rect 393144 191258 393186 191494
rect 393422 191258 393464 191494
rect 393144 184494 393464 191258
rect 393144 184258 393186 184494
rect 393422 184258 393464 184494
rect 393144 177494 393464 184258
rect 393144 177258 393186 177494
rect 393422 177258 393464 177494
rect 393144 170494 393464 177258
rect 393144 170258 393186 170494
rect 393422 170258 393464 170494
rect 393144 163494 393464 170258
rect 393144 163258 393186 163494
rect 393422 163258 393464 163494
rect 393144 156494 393464 163258
rect 393144 156258 393186 156494
rect 393422 156258 393464 156494
rect 393144 149494 393464 156258
rect 393144 149258 393186 149494
rect 393422 149258 393464 149494
rect 393144 142494 393464 149258
rect 393144 142258 393186 142494
rect 393422 142258 393464 142494
rect 393144 135494 393464 142258
rect 393144 135258 393186 135494
rect 393422 135258 393464 135494
rect 393144 128494 393464 135258
rect 393144 128258 393186 128494
rect 393422 128258 393464 128494
rect 393144 121494 393464 128258
rect 393144 121258 393186 121494
rect 393422 121258 393464 121494
rect 393144 114494 393464 121258
rect 393144 114258 393186 114494
rect 393422 114258 393464 114494
rect 393144 107494 393464 114258
rect 393144 107258 393186 107494
rect 393422 107258 393464 107494
rect 393144 100494 393464 107258
rect 393144 100258 393186 100494
rect 393422 100258 393464 100494
rect 393144 93494 393464 100258
rect 393144 93258 393186 93494
rect 393422 93258 393464 93494
rect 393144 86494 393464 93258
rect 393144 86258 393186 86494
rect 393422 86258 393464 86494
rect 393144 79494 393464 86258
rect 393144 79258 393186 79494
rect 393422 79258 393464 79494
rect 393144 72494 393464 79258
rect 393144 72258 393186 72494
rect 393422 72258 393464 72494
rect 393144 65494 393464 72258
rect 393144 65258 393186 65494
rect 393422 65258 393464 65494
rect 393144 58494 393464 65258
rect 393144 58258 393186 58494
rect 393422 58258 393464 58494
rect 393144 51494 393464 58258
rect 393144 51258 393186 51494
rect 393422 51258 393464 51494
rect 393144 44494 393464 51258
rect 393144 44258 393186 44494
rect 393422 44258 393464 44494
rect 393144 37494 393464 44258
rect 393144 37258 393186 37494
rect 393422 37258 393464 37494
rect 393144 30494 393464 37258
rect 393144 30258 393186 30494
rect 393422 30258 393464 30494
rect 393144 23494 393464 30258
rect 393144 23258 393186 23494
rect 393422 23258 393464 23494
rect 393144 16494 393464 23258
rect 393144 16258 393186 16494
rect 393422 16258 393464 16494
rect 393144 9494 393464 16258
rect 393144 9258 393186 9494
rect 393422 9258 393464 9494
rect 393144 2494 393464 9258
rect 393144 2258 393186 2494
rect 393422 2258 393464 2494
rect 393144 -746 393464 2258
rect 393144 -982 393186 -746
rect 393422 -982 393464 -746
rect 393144 -1066 393464 -982
rect 393144 -1302 393186 -1066
rect 393422 -1302 393464 -1066
rect 393144 -2294 393464 -1302
rect 394876 706198 395196 706230
rect 394876 705962 394918 706198
rect 395154 705962 395196 706198
rect 394876 705878 395196 705962
rect 394876 705642 394918 705878
rect 395154 705642 395196 705878
rect 394876 696561 395196 705642
rect 394876 696325 394918 696561
rect 395154 696325 395196 696561
rect 394876 689561 395196 696325
rect 394876 689325 394918 689561
rect 395154 689325 395196 689561
rect 394876 682561 395196 689325
rect 394876 682325 394918 682561
rect 395154 682325 395196 682561
rect 394876 675561 395196 682325
rect 394876 675325 394918 675561
rect 395154 675325 395196 675561
rect 394876 668561 395196 675325
rect 394876 668325 394918 668561
rect 395154 668325 395196 668561
rect 394876 661561 395196 668325
rect 394876 661325 394918 661561
rect 395154 661325 395196 661561
rect 394876 654561 395196 661325
rect 394876 654325 394918 654561
rect 395154 654325 395196 654561
rect 394876 647561 395196 654325
rect 394876 647325 394918 647561
rect 395154 647325 395196 647561
rect 394876 640561 395196 647325
rect 394876 640325 394918 640561
rect 395154 640325 395196 640561
rect 394876 633561 395196 640325
rect 394876 633325 394918 633561
rect 395154 633325 395196 633561
rect 394876 626561 395196 633325
rect 394876 626325 394918 626561
rect 395154 626325 395196 626561
rect 394876 619561 395196 626325
rect 394876 619325 394918 619561
rect 395154 619325 395196 619561
rect 394876 612561 395196 619325
rect 394876 612325 394918 612561
rect 395154 612325 395196 612561
rect 394876 605561 395196 612325
rect 394876 605325 394918 605561
rect 395154 605325 395196 605561
rect 394876 598561 395196 605325
rect 394876 598325 394918 598561
rect 395154 598325 395196 598561
rect 394876 591561 395196 598325
rect 394876 591325 394918 591561
rect 395154 591325 395196 591561
rect 394876 584561 395196 591325
rect 394876 584325 394918 584561
rect 395154 584325 395196 584561
rect 394876 577561 395196 584325
rect 394876 577325 394918 577561
rect 395154 577325 395196 577561
rect 394876 570561 395196 577325
rect 394876 570325 394918 570561
rect 395154 570325 395196 570561
rect 394876 563561 395196 570325
rect 394876 563325 394918 563561
rect 395154 563325 395196 563561
rect 394876 556561 395196 563325
rect 394876 556325 394918 556561
rect 395154 556325 395196 556561
rect 394876 549561 395196 556325
rect 394876 549325 394918 549561
rect 395154 549325 395196 549561
rect 394876 542561 395196 549325
rect 394876 542325 394918 542561
rect 395154 542325 395196 542561
rect 394876 535561 395196 542325
rect 394876 535325 394918 535561
rect 395154 535325 395196 535561
rect 394876 528561 395196 535325
rect 394876 528325 394918 528561
rect 395154 528325 395196 528561
rect 394876 521561 395196 528325
rect 394876 521325 394918 521561
rect 395154 521325 395196 521561
rect 394876 514561 395196 521325
rect 394876 514325 394918 514561
rect 395154 514325 395196 514561
rect 394876 507561 395196 514325
rect 394876 507325 394918 507561
rect 395154 507325 395196 507561
rect 394876 500561 395196 507325
rect 394876 500325 394918 500561
rect 395154 500325 395196 500561
rect 394876 493561 395196 500325
rect 394876 493325 394918 493561
rect 395154 493325 395196 493561
rect 394876 486561 395196 493325
rect 394876 486325 394918 486561
rect 395154 486325 395196 486561
rect 394876 479561 395196 486325
rect 394876 479325 394918 479561
rect 395154 479325 395196 479561
rect 394876 472561 395196 479325
rect 394876 472325 394918 472561
rect 395154 472325 395196 472561
rect 394876 465561 395196 472325
rect 394876 465325 394918 465561
rect 395154 465325 395196 465561
rect 394876 458561 395196 465325
rect 394876 458325 394918 458561
rect 395154 458325 395196 458561
rect 394876 451561 395196 458325
rect 394876 451325 394918 451561
rect 395154 451325 395196 451561
rect 394876 444561 395196 451325
rect 394876 444325 394918 444561
rect 395154 444325 395196 444561
rect 394876 437561 395196 444325
rect 394876 437325 394918 437561
rect 395154 437325 395196 437561
rect 394876 430561 395196 437325
rect 394876 430325 394918 430561
rect 395154 430325 395196 430561
rect 394876 423561 395196 430325
rect 394876 423325 394918 423561
rect 395154 423325 395196 423561
rect 394876 416561 395196 423325
rect 394876 416325 394918 416561
rect 395154 416325 395196 416561
rect 394876 409561 395196 416325
rect 394876 409325 394918 409561
rect 395154 409325 395196 409561
rect 394876 402561 395196 409325
rect 394876 402325 394918 402561
rect 395154 402325 395196 402561
rect 394876 395561 395196 402325
rect 394876 395325 394918 395561
rect 395154 395325 395196 395561
rect 394876 388561 395196 395325
rect 394876 388325 394918 388561
rect 395154 388325 395196 388561
rect 394876 381561 395196 388325
rect 394876 381325 394918 381561
rect 395154 381325 395196 381561
rect 394876 374561 395196 381325
rect 394876 374325 394918 374561
rect 395154 374325 395196 374561
rect 394876 367561 395196 374325
rect 394876 367325 394918 367561
rect 395154 367325 395196 367561
rect 394876 360561 395196 367325
rect 394876 360325 394918 360561
rect 395154 360325 395196 360561
rect 394876 353561 395196 360325
rect 394876 353325 394918 353561
rect 395154 353325 395196 353561
rect 394876 346561 395196 353325
rect 394876 346325 394918 346561
rect 395154 346325 395196 346561
rect 394876 339561 395196 346325
rect 394876 339325 394918 339561
rect 395154 339325 395196 339561
rect 394876 332561 395196 339325
rect 394876 332325 394918 332561
rect 395154 332325 395196 332561
rect 394876 325561 395196 332325
rect 394876 325325 394918 325561
rect 395154 325325 395196 325561
rect 394876 318561 395196 325325
rect 394876 318325 394918 318561
rect 395154 318325 395196 318561
rect 394876 311561 395196 318325
rect 394876 311325 394918 311561
rect 395154 311325 395196 311561
rect 394876 304561 395196 311325
rect 394876 304325 394918 304561
rect 395154 304325 395196 304561
rect 394876 297561 395196 304325
rect 394876 297325 394918 297561
rect 395154 297325 395196 297561
rect 394876 290561 395196 297325
rect 394876 290325 394918 290561
rect 395154 290325 395196 290561
rect 394876 283561 395196 290325
rect 394876 283325 394918 283561
rect 395154 283325 395196 283561
rect 394876 276561 395196 283325
rect 394876 276325 394918 276561
rect 395154 276325 395196 276561
rect 394876 269561 395196 276325
rect 394876 269325 394918 269561
rect 395154 269325 395196 269561
rect 394876 262561 395196 269325
rect 394876 262325 394918 262561
rect 395154 262325 395196 262561
rect 394876 255561 395196 262325
rect 394876 255325 394918 255561
rect 395154 255325 395196 255561
rect 394876 248561 395196 255325
rect 394876 248325 394918 248561
rect 395154 248325 395196 248561
rect 394876 241561 395196 248325
rect 394876 241325 394918 241561
rect 395154 241325 395196 241561
rect 394876 234561 395196 241325
rect 394876 234325 394918 234561
rect 395154 234325 395196 234561
rect 394876 227561 395196 234325
rect 394876 227325 394918 227561
rect 395154 227325 395196 227561
rect 394876 220561 395196 227325
rect 394876 220325 394918 220561
rect 395154 220325 395196 220561
rect 394876 213561 395196 220325
rect 394876 213325 394918 213561
rect 395154 213325 395196 213561
rect 394876 206561 395196 213325
rect 394876 206325 394918 206561
rect 395154 206325 395196 206561
rect 394876 199561 395196 206325
rect 394876 199325 394918 199561
rect 395154 199325 395196 199561
rect 394876 192561 395196 199325
rect 394876 192325 394918 192561
rect 395154 192325 395196 192561
rect 394876 185561 395196 192325
rect 394876 185325 394918 185561
rect 395154 185325 395196 185561
rect 394876 178561 395196 185325
rect 394876 178325 394918 178561
rect 395154 178325 395196 178561
rect 394876 171561 395196 178325
rect 394876 171325 394918 171561
rect 395154 171325 395196 171561
rect 394876 164561 395196 171325
rect 394876 164325 394918 164561
rect 395154 164325 395196 164561
rect 394876 157561 395196 164325
rect 394876 157325 394918 157561
rect 395154 157325 395196 157561
rect 394876 150561 395196 157325
rect 394876 150325 394918 150561
rect 395154 150325 395196 150561
rect 394876 143561 395196 150325
rect 394876 143325 394918 143561
rect 395154 143325 395196 143561
rect 394876 136561 395196 143325
rect 394876 136325 394918 136561
rect 395154 136325 395196 136561
rect 394876 129561 395196 136325
rect 394876 129325 394918 129561
rect 395154 129325 395196 129561
rect 394876 122561 395196 129325
rect 394876 122325 394918 122561
rect 395154 122325 395196 122561
rect 394876 115561 395196 122325
rect 394876 115325 394918 115561
rect 395154 115325 395196 115561
rect 394876 108561 395196 115325
rect 394876 108325 394918 108561
rect 395154 108325 395196 108561
rect 394876 101561 395196 108325
rect 394876 101325 394918 101561
rect 395154 101325 395196 101561
rect 394876 94561 395196 101325
rect 394876 94325 394918 94561
rect 395154 94325 395196 94561
rect 394876 87561 395196 94325
rect 394876 87325 394918 87561
rect 395154 87325 395196 87561
rect 394876 80561 395196 87325
rect 394876 80325 394918 80561
rect 395154 80325 395196 80561
rect 394876 73561 395196 80325
rect 394876 73325 394918 73561
rect 395154 73325 395196 73561
rect 394876 66561 395196 73325
rect 394876 66325 394918 66561
rect 395154 66325 395196 66561
rect 394876 59561 395196 66325
rect 394876 59325 394918 59561
rect 395154 59325 395196 59561
rect 394876 52561 395196 59325
rect 394876 52325 394918 52561
rect 395154 52325 395196 52561
rect 394876 45561 395196 52325
rect 394876 45325 394918 45561
rect 395154 45325 395196 45561
rect 394876 38561 395196 45325
rect 394876 38325 394918 38561
rect 395154 38325 395196 38561
rect 394876 31561 395196 38325
rect 394876 31325 394918 31561
rect 395154 31325 395196 31561
rect 394876 24561 395196 31325
rect 394876 24325 394918 24561
rect 395154 24325 395196 24561
rect 394876 17561 395196 24325
rect 394876 17325 394918 17561
rect 395154 17325 395196 17561
rect 394876 10561 395196 17325
rect 394876 10325 394918 10561
rect 395154 10325 395196 10561
rect 394876 3561 395196 10325
rect 394876 3325 394918 3561
rect 395154 3325 395196 3561
rect 394876 -1706 395196 3325
rect 394876 -1942 394918 -1706
rect 395154 -1942 395196 -1706
rect 394876 -2026 395196 -1942
rect 394876 -2262 394918 -2026
rect 395154 -2262 395196 -2026
rect 394876 -2294 395196 -2262
rect 400144 705238 400464 706230
rect 400144 705002 400186 705238
rect 400422 705002 400464 705238
rect 400144 704918 400464 705002
rect 400144 704682 400186 704918
rect 400422 704682 400464 704918
rect 400144 695494 400464 704682
rect 400144 695258 400186 695494
rect 400422 695258 400464 695494
rect 400144 688494 400464 695258
rect 400144 688258 400186 688494
rect 400422 688258 400464 688494
rect 400144 681494 400464 688258
rect 400144 681258 400186 681494
rect 400422 681258 400464 681494
rect 400144 674494 400464 681258
rect 400144 674258 400186 674494
rect 400422 674258 400464 674494
rect 400144 667494 400464 674258
rect 400144 667258 400186 667494
rect 400422 667258 400464 667494
rect 400144 660494 400464 667258
rect 400144 660258 400186 660494
rect 400422 660258 400464 660494
rect 400144 653494 400464 660258
rect 400144 653258 400186 653494
rect 400422 653258 400464 653494
rect 400144 646494 400464 653258
rect 400144 646258 400186 646494
rect 400422 646258 400464 646494
rect 400144 639494 400464 646258
rect 400144 639258 400186 639494
rect 400422 639258 400464 639494
rect 400144 632494 400464 639258
rect 400144 632258 400186 632494
rect 400422 632258 400464 632494
rect 400144 625494 400464 632258
rect 400144 625258 400186 625494
rect 400422 625258 400464 625494
rect 400144 618494 400464 625258
rect 400144 618258 400186 618494
rect 400422 618258 400464 618494
rect 400144 611494 400464 618258
rect 400144 611258 400186 611494
rect 400422 611258 400464 611494
rect 400144 604494 400464 611258
rect 400144 604258 400186 604494
rect 400422 604258 400464 604494
rect 400144 597494 400464 604258
rect 400144 597258 400186 597494
rect 400422 597258 400464 597494
rect 400144 590494 400464 597258
rect 400144 590258 400186 590494
rect 400422 590258 400464 590494
rect 400144 583494 400464 590258
rect 400144 583258 400186 583494
rect 400422 583258 400464 583494
rect 400144 576494 400464 583258
rect 400144 576258 400186 576494
rect 400422 576258 400464 576494
rect 400144 569494 400464 576258
rect 400144 569258 400186 569494
rect 400422 569258 400464 569494
rect 400144 562494 400464 569258
rect 400144 562258 400186 562494
rect 400422 562258 400464 562494
rect 400144 555494 400464 562258
rect 400144 555258 400186 555494
rect 400422 555258 400464 555494
rect 400144 548494 400464 555258
rect 400144 548258 400186 548494
rect 400422 548258 400464 548494
rect 400144 541494 400464 548258
rect 400144 541258 400186 541494
rect 400422 541258 400464 541494
rect 400144 534494 400464 541258
rect 400144 534258 400186 534494
rect 400422 534258 400464 534494
rect 400144 527494 400464 534258
rect 400144 527258 400186 527494
rect 400422 527258 400464 527494
rect 400144 520494 400464 527258
rect 400144 520258 400186 520494
rect 400422 520258 400464 520494
rect 400144 513494 400464 520258
rect 400144 513258 400186 513494
rect 400422 513258 400464 513494
rect 400144 506494 400464 513258
rect 400144 506258 400186 506494
rect 400422 506258 400464 506494
rect 400144 499494 400464 506258
rect 400144 499258 400186 499494
rect 400422 499258 400464 499494
rect 400144 492494 400464 499258
rect 400144 492258 400186 492494
rect 400422 492258 400464 492494
rect 400144 485494 400464 492258
rect 400144 485258 400186 485494
rect 400422 485258 400464 485494
rect 400144 478494 400464 485258
rect 400144 478258 400186 478494
rect 400422 478258 400464 478494
rect 400144 471494 400464 478258
rect 400144 471258 400186 471494
rect 400422 471258 400464 471494
rect 400144 464494 400464 471258
rect 400144 464258 400186 464494
rect 400422 464258 400464 464494
rect 400144 457494 400464 464258
rect 400144 457258 400186 457494
rect 400422 457258 400464 457494
rect 400144 450494 400464 457258
rect 400144 450258 400186 450494
rect 400422 450258 400464 450494
rect 400144 443494 400464 450258
rect 400144 443258 400186 443494
rect 400422 443258 400464 443494
rect 400144 436494 400464 443258
rect 400144 436258 400186 436494
rect 400422 436258 400464 436494
rect 400144 429494 400464 436258
rect 400144 429258 400186 429494
rect 400422 429258 400464 429494
rect 400144 422494 400464 429258
rect 400144 422258 400186 422494
rect 400422 422258 400464 422494
rect 400144 415494 400464 422258
rect 400144 415258 400186 415494
rect 400422 415258 400464 415494
rect 400144 408494 400464 415258
rect 400144 408258 400186 408494
rect 400422 408258 400464 408494
rect 400144 401494 400464 408258
rect 400144 401258 400186 401494
rect 400422 401258 400464 401494
rect 400144 394494 400464 401258
rect 400144 394258 400186 394494
rect 400422 394258 400464 394494
rect 400144 387494 400464 394258
rect 400144 387258 400186 387494
rect 400422 387258 400464 387494
rect 400144 380494 400464 387258
rect 400144 380258 400186 380494
rect 400422 380258 400464 380494
rect 400144 373494 400464 380258
rect 400144 373258 400186 373494
rect 400422 373258 400464 373494
rect 400144 366494 400464 373258
rect 400144 366258 400186 366494
rect 400422 366258 400464 366494
rect 400144 359494 400464 366258
rect 400144 359258 400186 359494
rect 400422 359258 400464 359494
rect 400144 352494 400464 359258
rect 400144 352258 400186 352494
rect 400422 352258 400464 352494
rect 400144 345494 400464 352258
rect 400144 345258 400186 345494
rect 400422 345258 400464 345494
rect 400144 338494 400464 345258
rect 400144 338258 400186 338494
rect 400422 338258 400464 338494
rect 400144 331494 400464 338258
rect 400144 331258 400186 331494
rect 400422 331258 400464 331494
rect 400144 324494 400464 331258
rect 400144 324258 400186 324494
rect 400422 324258 400464 324494
rect 400144 317494 400464 324258
rect 400144 317258 400186 317494
rect 400422 317258 400464 317494
rect 400144 310494 400464 317258
rect 400144 310258 400186 310494
rect 400422 310258 400464 310494
rect 400144 303494 400464 310258
rect 400144 303258 400186 303494
rect 400422 303258 400464 303494
rect 400144 296494 400464 303258
rect 400144 296258 400186 296494
rect 400422 296258 400464 296494
rect 400144 289494 400464 296258
rect 400144 289258 400186 289494
rect 400422 289258 400464 289494
rect 400144 282494 400464 289258
rect 400144 282258 400186 282494
rect 400422 282258 400464 282494
rect 400144 275494 400464 282258
rect 400144 275258 400186 275494
rect 400422 275258 400464 275494
rect 400144 268494 400464 275258
rect 400144 268258 400186 268494
rect 400422 268258 400464 268494
rect 400144 261494 400464 268258
rect 400144 261258 400186 261494
rect 400422 261258 400464 261494
rect 400144 254494 400464 261258
rect 400144 254258 400186 254494
rect 400422 254258 400464 254494
rect 400144 247494 400464 254258
rect 400144 247258 400186 247494
rect 400422 247258 400464 247494
rect 400144 240494 400464 247258
rect 400144 240258 400186 240494
rect 400422 240258 400464 240494
rect 400144 233494 400464 240258
rect 400144 233258 400186 233494
rect 400422 233258 400464 233494
rect 400144 226494 400464 233258
rect 400144 226258 400186 226494
rect 400422 226258 400464 226494
rect 400144 219494 400464 226258
rect 400144 219258 400186 219494
rect 400422 219258 400464 219494
rect 400144 212494 400464 219258
rect 400144 212258 400186 212494
rect 400422 212258 400464 212494
rect 400144 205494 400464 212258
rect 400144 205258 400186 205494
rect 400422 205258 400464 205494
rect 400144 198494 400464 205258
rect 400144 198258 400186 198494
rect 400422 198258 400464 198494
rect 400144 191494 400464 198258
rect 400144 191258 400186 191494
rect 400422 191258 400464 191494
rect 400144 184494 400464 191258
rect 400144 184258 400186 184494
rect 400422 184258 400464 184494
rect 400144 177494 400464 184258
rect 400144 177258 400186 177494
rect 400422 177258 400464 177494
rect 400144 170494 400464 177258
rect 400144 170258 400186 170494
rect 400422 170258 400464 170494
rect 400144 163494 400464 170258
rect 400144 163258 400186 163494
rect 400422 163258 400464 163494
rect 400144 156494 400464 163258
rect 400144 156258 400186 156494
rect 400422 156258 400464 156494
rect 400144 149494 400464 156258
rect 400144 149258 400186 149494
rect 400422 149258 400464 149494
rect 400144 142494 400464 149258
rect 400144 142258 400186 142494
rect 400422 142258 400464 142494
rect 400144 135494 400464 142258
rect 400144 135258 400186 135494
rect 400422 135258 400464 135494
rect 400144 128494 400464 135258
rect 400144 128258 400186 128494
rect 400422 128258 400464 128494
rect 400144 121494 400464 128258
rect 400144 121258 400186 121494
rect 400422 121258 400464 121494
rect 400144 114494 400464 121258
rect 400144 114258 400186 114494
rect 400422 114258 400464 114494
rect 400144 107494 400464 114258
rect 400144 107258 400186 107494
rect 400422 107258 400464 107494
rect 400144 100494 400464 107258
rect 400144 100258 400186 100494
rect 400422 100258 400464 100494
rect 400144 93494 400464 100258
rect 400144 93258 400186 93494
rect 400422 93258 400464 93494
rect 400144 86494 400464 93258
rect 400144 86258 400186 86494
rect 400422 86258 400464 86494
rect 400144 79494 400464 86258
rect 400144 79258 400186 79494
rect 400422 79258 400464 79494
rect 400144 72494 400464 79258
rect 400144 72258 400186 72494
rect 400422 72258 400464 72494
rect 400144 65494 400464 72258
rect 400144 65258 400186 65494
rect 400422 65258 400464 65494
rect 400144 58494 400464 65258
rect 400144 58258 400186 58494
rect 400422 58258 400464 58494
rect 400144 51494 400464 58258
rect 400144 51258 400186 51494
rect 400422 51258 400464 51494
rect 400144 44494 400464 51258
rect 400144 44258 400186 44494
rect 400422 44258 400464 44494
rect 400144 37494 400464 44258
rect 400144 37258 400186 37494
rect 400422 37258 400464 37494
rect 400144 30494 400464 37258
rect 400144 30258 400186 30494
rect 400422 30258 400464 30494
rect 400144 23494 400464 30258
rect 400144 23258 400186 23494
rect 400422 23258 400464 23494
rect 400144 16494 400464 23258
rect 400144 16258 400186 16494
rect 400422 16258 400464 16494
rect 400144 9494 400464 16258
rect 400144 9258 400186 9494
rect 400422 9258 400464 9494
rect 400144 2494 400464 9258
rect 400144 2258 400186 2494
rect 400422 2258 400464 2494
rect 400144 -746 400464 2258
rect 400144 -982 400186 -746
rect 400422 -982 400464 -746
rect 400144 -1066 400464 -982
rect 400144 -1302 400186 -1066
rect 400422 -1302 400464 -1066
rect 400144 -2294 400464 -1302
rect 401876 706198 402196 706230
rect 401876 705962 401918 706198
rect 402154 705962 402196 706198
rect 401876 705878 402196 705962
rect 401876 705642 401918 705878
rect 402154 705642 402196 705878
rect 401876 696561 402196 705642
rect 401876 696325 401918 696561
rect 402154 696325 402196 696561
rect 401876 689561 402196 696325
rect 401876 689325 401918 689561
rect 402154 689325 402196 689561
rect 401876 682561 402196 689325
rect 401876 682325 401918 682561
rect 402154 682325 402196 682561
rect 401876 675561 402196 682325
rect 401876 675325 401918 675561
rect 402154 675325 402196 675561
rect 401876 668561 402196 675325
rect 401876 668325 401918 668561
rect 402154 668325 402196 668561
rect 401876 661561 402196 668325
rect 401876 661325 401918 661561
rect 402154 661325 402196 661561
rect 401876 654561 402196 661325
rect 401876 654325 401918 654561
rect 402154 654325 402196 654561
rect 401876 647561 402196 654325
rect 401876 647325 401918 647561
rect 402154 647325 402196 647561
rect 401876 640561 402196 647325
rect 401876 640325 401918 640561
rect 402154 640325 402196 640561
rect 401876 633561 402196 640325
rect 401876 633325 401918 633561
rect 402154 633325 402196 633561
rect 401876 626561 402196 633325
rect 401876 626325 401918 626561
rect 402154 626325 402196 626561
rect 401876 619561 402196 626325
rect 401876 619325 401918 619561
rect 402154 619325 402196 619561
rect 401876 612561 402196 619325
rect 401876 612325 401918 612561
rect 402154 612325 402196 612561
rect 401876 605561 402196 612325
rect 401876 605325 401918 605561
rect 402154 605325 402196 605561
rect 401876 598561 402196 605325
rect 401876 598325 401918 598561
rect 402154 598325 402196 598561
rect 401876 591561 402196 598325
rect 401876 591325 401918 591561
rect 402154 591325 402196 591561
rect 401876 584561 402196 591325
rect 401876 584325 401918 584561
rect 402154 584325 402196 584561
rect 401876 577561 402196 584325
rect 401876 577325 401918 577561
rect 402154 577325 402196 577561
rect 401876 570561 402196 577325
rect 401876 570325 401918 570561
rect 402154 570325 402196 570561
rect 401876 563561 402196 570325
rect 401876 563325 401918 563561
rect 402154 563325 402196 563561
rect 401876 556561 402196 563325
rect 401876 556325 401918 556561
rect 402154 556325 402196 556561
rect 401876 549561 402196 556325
rect 401876 549325 401918 549561
rect 402154 549325 402196 549561
rect 401876 542561 402196 549325
rect 401876 542325 401918 542561
rect 402154 542325 402196 542561
rect 401876 535561 402196 542325
rect 401876 535325 401918 535561
rect 402154 535325 402196 535561
rect 401876 528561 402196 535325
rect 401876 528325 401918 528561
rect 402154 528325 402196 528561
rect 401876 521561 402196 528325
rect 401876 521325 401918 521561
rect 402154 521325 402196 521561
rect 401876 514561 402196 521325
rect 401876 514325 401918 514561
rect 402154 514325 402196 514561
rect 401876 507561 402196 514325
rect 401876 507325 401918 507561
rect 402154 507325 402196 507561
rect 401876 500561 402196 507325
rect 401876 500325 401918 500561
rect 402154 500325 402196 500561
rect 401876 493561 402196 500325
rect 401876 493325 401918 493561
rect 402154 493325 402196 493561
rect 401876 486561 402196 493325
rect 401876 486325 401918 486561
rect 402154 486325 402196 486561
rect 401876 479561 402196 486325
rect 401876 479325 401918 479561
rect 402154 479325 402196 479561
rect 401876 472561 402196 479325
rect 401876 472325 401918 472561
rect 402154 472325 402196 472561
rect 401876 465561 402196 472325
rect 401876 465325 401918 465561
rect 402154 465325 402196 465561
rect 401876 458561 402196 465325
rect 401876 458325 401918 458561
rect 402154 458325 402196 458561
rect 401876 451561 402196 458325
rect 401876 451325 401918 451561
rect 402154 451325 402196 451561
rect 401876 444561 402196 451325
rect 401876 444325 401918 444561
rect 402154 444325 402196 444561
rect 401876 437561 402196 444325
rect 401876 437325 401918 437561
rect 402154 437325 402196 437561
rect 401876 430561 402196 437325
rect 401876 430325 401918 430561
rect 402154 430325 402196 430561
rect 401876 423561 402196 430325
rect 401876 423325 401918 423561
rect 402154 423325 402196 423561
rect 401876 416561 402196 423325
rect 401876 416325 401918 416561
rect 402154 416325 402196 416561
rect 401876 409561 402196 416325
rect 401876 409325 401918 409561
rect 402154 409325 402196 409561
rect 401876 402561 402196 409325
rect 401876 402325 401918 402561
rect 402154 402325 402196 402561
rect 401876 395561 402196 402325
rect 401876 395325 401918 395561
rect 402154 395325 402196 395561
rect 401876 388561 402196 395325
rect 401876 388325 401918 388561
rect 402154 388325 402196 388561
rect 401876 381561 402196 388325
rect 401876 381325 401918 381561
rect 402154 381325 402196 381561
rect 401876 374561 402196 381325
rect 401876 374325 401918 374561
rect 402154 374325 402196 374561
rect 401876 367561 402196 374325
rect 401876 367325 401918 367561
rect 402154 367325 402196 367561
rect 401876 360561 402196 367325
rect 401876 360325 401918 360561
rect 402154 360325 402196 360561
rect 401876 353561 402196 360325
rect 401876 353325 401918 353561
rect 402154 353325 402196 353561
rect 401876 346561 402196 353325
rect 401876 346325 401918 346561
rect 402154 346325 402196 346561
rect 401876 339561 402196 346325
rect 401876 339325 401918 339561
rect 402154 339325 402196 339561
rect 401876 332561 402196 339325
rect 401876 332325 401918 332561
rect 402154 332325 402196 332561
rect 401876 325561 402196 332325
rect 401876 325325 401918 325561
rect 402154 325325 402196 325561
rect 401876 318561 402196 325325
rect 401876 318325 401918 318561
rect 402154 318325 402196 318561
rect 401876 311561 402196 318325
rect 401876 311325 401918 311561
rect 402154 311325 402196 311561
rect 401876 304561 402196 311325
rect 401876 304325 401918 304561
rect 402154 304325 402196 304561
rect 401876 297561 402196 304325
rect 401876 297325 401918 297561
rect 402154 297325 402196 297561
rect 401876 290561 402196 297325
rect 401876 290325 401918 290561
rect 402154 290325 402196 290561
rect 401876 283561 402196 290325
rect 401876 283325 401918 283561
rect 402154 283325 402196 283561
rect 401876 276561 402196 283325
rect 401876 276325 401918 276561
rect 402154 276325 402196 276561
rect 401876 269561 402196 276325
rect 401876 269325 401918 269561
rect 402154 269325 402196 269561
rect 401876 262561 402196 269325
rect 401876 262325 401918 262561
rect 402154 262325 402196 262561
rect 401876 255561 402196 262325
rect 401876 255325 401918 255561
rect 402154 255325 402196 255561
rect 401876 248561 402196 255325
rect 401876 248325 401918 248561
rect 402154 248325 402196 248561
rect 401876 241561 402196 248325
rect 401876 241325 401918 241561
rect 402154 241325 402196 241561
rect 401876 234561 402196 241325
rect 401876 234325 401918 234561
rect 402154 234325 402196 234561
rect 401876 227561 402196 234325
rect 401876 227325 401918 227561
rect 402154 227325 402196 227561
rect 401876 220561 402196 227325
rect 401876 220325 401918 220561
rect 402154 220325 402196 220561
rect 401876 213561 402196 220325
rect 401876 213325 401918 213561
rect 402154 213325 402196 213561
rect 401876 206561 402196 213325
rect 401876 206325 401918 206561
rect 402154 206325 402196 206561
rect 401876 199561 402196 206325
rect 401876 199325 401918 199561
rect 402154 199325 402196 199561
rect 401876 192561 402196 199325
rect 401876 192325 401918 192561
rect 402154 192325 402196 192561
rect 401876 185561 402196 192325
rect 401876 185325 401918 185561
rect 402154 185325 402196 185561
rect 401876 178561 402196 185325
rect 401876 178325 401918 178561
rect 402154 178325 402196 178561
rect 401876 171561 402196 178325
rect 401876 171325 401918 171561
rect 402154 171325 402196 171561
rect 401876 164561 402196 171325
rect 401876 164325 401918 164561
rect 402154 164325 402196 164561
rect 401876 157561 402196 164325
rect 401876 157325 401918 157561
rect 402154 157325 402196 157561
rect 401876 150561 402196 157325
rect 401876 150325 401918 150561
rect 402154 150325 402196 150561
rect 401876 143561 402196 150325
rect 401876 143325 401918 143561
rect 402154 143325 402196 143561
rect 401876 136561 402196 143325
rect 401876 136325 401918 136561
rect 402154 136325 402196 136561
rect 401876 129561 402196 136325
rect 401876 129325 401918 129561
rect 402154 129325 402196 129561
rect 401876 122561 402196 129325
rect 401876 122325 401918 122561
rect 402154 122325 402196 122561
rect 401876 115561 402196 122325
rect 401876 115325 401918 115561
rect 402154 115325 402196 115561
rect 401876 108561 402196 115325
rect 401876 108325 401918 108561
rect 402154 108325 402196 108561
rect 401876 101561 402196 108325
rect 401876 101325 401918 101561
rect 402154 101325 402196 101561
rect 401876 94561 402196 101325
rect 401876 94325 401918 94561
rect 402154 94325 402196 94561
rect 401876 87561 402196 94325
rect 401876 87325 401918 87561
rect 402154 87325 402196 87561
rect 401876 80561 402196 87325
rect 401876 80325 401918 80561
rect 402154 80325 402196 80561
rect 401876 73561 402196 80325
rect 401876 73325 401918 73561
rect 402154 73325 402196 73561
rect 401876 66561 402196 73325
rect 401876 66325 401918 66561
rect 402154 66325 402196 66561
rect 401876 59561 402196 66325
rect 401876 59325 401918 59561
rect 402154 59325 402196 59561
rect 401876 52561 402196 59325
rect 401876 52325 401918 52561
rect 402154 52325 402196 52561
rect 401876 45561 402196 52325
rect 401876 45325 401918 45561
rect 402154 45325 402196 45561
rect 401876 38561 402196 45325
rect 401876 38325 401918 38561
rect 402154 38325 402196 38561
rect 401876 31561 402196 38325
rect 401876 31325 401918 31561
rect 402154 31325 402196 31561
rect 401876 24561 402196 31325
rect 401876 24325 401918 24561
rect 402154 24325 402196 24561
rect 401876 17561 402196 24325
rect 401876 17325 401918 17561
rect 402154 17325 402196 17561
rect 401876 10561 402196 17325
rect 401876 10325 401918 10561
rect 402154 10325 402196 10561
rect 401876 3561 402196 10325
rect 401876 3325 401918 3561
rect 402154 3325 402196 3561
rect 401876 -1706 402196 3325
rect 401876 -1942 401918 -1706
rect 402154 -1942 402196 -1706
rect 401876 -2026 402196 -1942
rect 401876 -2262 401918 -2026
rect 402154 -2262 402196 -2026
rect 401876 -2294 402196 -2262
rect 407144 705238 407464 706230
rect 407144 705002 407186 705238
rect 407422 705002 407464 705238
rect 407144 704918 407464 705002
rect 407144 704682 407186 704918
rect 407422 704682 407464 704918
rect 407144 695494 407464 704682
rect 407144 695258 407186 695494
rect 407422 695258 407464 695494
rect 407144 688494 407464 695258
rect 407144 688258 407186 688494
rect 407422 688258 407464 688494
rect 407144 681494 407464 688258
rect 407144 681258 407186 681494
rect 407422 681258 407464 681494
rect 407144 674494 407464 681258
rect 407144 674258 407186 674494
rect 407422 674258 407464 674494
rect 407144 667494 407464 674258
rect 407144 667258 407186 667494
rect 407422 667258 407464 667494
rect 407144 660494 407464 667258
rect 407144 660258 407186 660494
rect 407422 660258 407464 660494
rect 407144 653494 407464 660258
rect 407144 653258 407186 653494
rect 407422 653258 407464 653494
rect 407144 646494 407464 653258
rect 407144 646258 407186 646494
rect 407422 646258 407464 646494
rect 407144 639494 407464 646258
rect 407144 639258 407186 639494
rect 407422 639258 407464 639494
rect 407144 632494 407464 639258
rect 407144 632258 407186 632494
rect 407422 632258 407464 632494
rect 407144 625494 407464 632258
rect 407144 625258 407186 625494
rect 407422 625258 407464 625494
rect 407144 618494 407464 625258
rect 407144 618258 407186 618494
rect 407422 618258 407464 618494
rect 407144 611494 407464 618258
rect 407144 611258 407186 611494
rect 407422 611258 407464 611494
rect 407144 604494 407464 611258
rect 407144 604258 407186 604494
rect 407422 604258 407464 604494
rect 407144 597494 407464 604258
rect 407144 597258 407186 597494
rect 407422 597258 407464 597494
rect 407144 590494 407464 597258
rect 407144 590258 407186 590494
rect 407422 590258 407464 590494
rect 407144 583494 407464 590258
rect 407144 583258 407186 583494
rect 407422 583258 407464 583494
rect 407144 576494 407464 583258
rect 407144 576258 407186 576494
rect 407422 576258 407464 576494
rect 407144 569494 407464 576258
rect 407144 569258 407186 569494
rect 407422 569258 407464 569494
rect 407144 562494 407464 569258
rect 407144 562258 407186 562494
rect 407422 562258 407464 562494
rect 407144 555494 407464 562258
rect 407144 555258 407186 555494
rect 407422 555258 407464 555494
rect 407144 548494 407464 555258
rect 407144 548258 407186 548494
rect 407422 548258 407464 548494
rect 407144 541494 407464 548258
rect 407144 541258 407186 541494
rect 407422 541258 407464 541494
rect 407144 534494 407464 541258
rect 407144 534258 407186 534494
rect 407422 534258 407464 534494
rect 407144 527494 407464 534258
rect 407144 527258 407186 527494
rect 407422 527258 407464 527494
rect 407144 520494 407464 527258
rect 407144 520258 407186 520494
rect 407422 520258 407464 520494
rect 407144 513494 407464 520258
rect 407144 513258 407186 513494
rect 407422 513258 407464 513494
rect 407144 506494 407464 513258
rect 407144 506258 407186 506494
rect 407422 506258 407464 506494
rect 407144 499494 407464 506258
rect 407144 499258 407186 499494
rect 407422 499258 407464 499494
rect 407144 492494 407464 499258
rect 407144 492258 407186 492494
rect 407422 492258 407464 492494
rect 407144 485494 407464 492258
rect 407144 485258 407186 485494
rect 407422 485258 407464 485494
rect 407144 478494 407464 485258
rect 407144 478258 407186 478494
rect 407422 478258 407464 478494
rect 407144 471494 407464 478258
rect 407144 471258 407186 471494
rect 407422 471258 407464 471494
rect 407144 464494 407464 471258
rect 407144 464258 407186 464494
rect 407422 464258 407464 464494
rect 407144 457494 407464 464258
rect 407144 457258 407186 457494
rect 407422 457258 407464 457494
rect 407144 450494 407464 457258
rect 407144 450258 407186 450494
rect 407422 450258 407464 450494
rect 407144 443494 407464 450258
rect 407144 443258 407186 443494
rect 407422 443258 407464 443494
rect 407144 436494 407464 443258
rect 407144 436258 407186 436494
rect 407422 436258 407464 436494
rect 407144 429494 407464 436258
rect 407144 429258 407186 429494
rect 407422 429258 407464 429494
rect 407144 422494 407464 429258
rect 407144 422258 407186 422494
rect 407422 422258 407464 422494
rect 407144 415494 407464 422258
rect 407144 415258 407186 415494
rect 407422 415258 407464 415494
rect 407144 408494 407464 415258
rect 407144 408258 407186 408494
rect 407422 408258 407464 408494
rect 407144 401494 407464 408258
rect 407144 401258 407186 401494
rect 407422 401258 407464 401494
rect 407144 394494 407464 401258
rect 407144 394258 407186 394494
rect 407422 394258 407464 394494
rect 407144 387494 407464 394258
rect 407144 387258 407186 387494
rect 407422 387258 407464 387494
rect 407144 380494 407464 387258
rect 407144 380258 407186 380494
rect 407422 380258 407464 380494
rect 407144 373494 407464 380258
rect 407144 373258 407186 373494
rect 407422 373258 407464 373494
rect 407144 366494 407464 373258
rect 407144 366258 407186 366494
rect 407422 366258 407464 366494
rect 407144 359494 407464 366258
rect 407144 359258 407186 359494
rect 407422 359258 407464 359494
rect 407144 352494 407464 359258
rect 407144 352258 407186 352494
rect 407422 352258 407464 352494
rect 407144 345494 407464 352258
rect 407144 345258 407186 345494
rect 407422 345258 407464 345494
rect 407144 338494 407464 345258
rect 407144 338258 407186 338494
rect 407422 338258 407464 338494
rect 407144 331494 407464 338258
rect 407144 331258 407186 331494
rect 407422 331258 407464 331494
rect 407144 324494 407464 331258
rect 407144 324258 407186 324494
rect 407422 324258 407464 324494
rect 407144 317494 407464 324258
rect 407144 317258 407186 317494
rect 407422 317258 407464 317494
rect 407144 310494 407464 317258
rect 407144 310258 407186 310494
rect 407422 310258 407464 310494
rect 407144 303494 407464 310258
rect 407144 303258 407186 303494
rect 407422 303258 407464 303494
rect 407144 296494 407464 303258
rect 407144 296258 407186 296494
rect 407422 296258 407464 296494
rect 407144 289494 407464 296258
rect 407144 289258 407186 289494
rect 407422 289258 407464 289494
rect 407144 282494 407464 289258
rect 407144 282258 407186 282494
rect 407422 282258 407464 282494
rect 407144 275494 407464 282258
rect 407144 275258 407186 275494
rect 407422 275258 407464 275494
rect 407144 268494 407464 275258
rect 407144 268258 407186 268494
rect 407422 268258 407464 268494
rect 407144 261494 407464 268258
rect 407144 261258 407186 261494
rect 407422 261258 407464 261494
rect 407144 254494 407464 261258
rect 407144 254258 407186 254494
rect 407422 254258 407464 254494
rect 407144 247494 407464 254258
rect 407144 247258 407186 247494
rect 407422 247258 407464 247494
rect 407144 240494 407464 247258
rect 407144 240258 407186 240494
rect 407422 240258 407464 240494
rect 407144 233494 407464 240258
rect 407144 233258 407186 233494
rect 407422 233258 407464 233494
rect 407144 226494 407464 233258
rect 407144 226258 407186 226494
rect 407422 226258 407464 226494
rect 407144 219494 407464 226258
rect 407144 219258 407186 219494
rect 407422 219258 407464 219494
rect 407144 212494 407464 219258
rect 407144 212258 407186 212494
rect 407422 212258 407464 212494
rect 407144 205494 407464 212258
rect 407144 205258 407186 205494
rect 407422 205258 407464 205494
rect 407144 198494 407464 205258
rect 407144 198258 407186 198494
rect 407422 198258 407464 198494
rect 407144 191494 407464 198258
rect 407144 191258 407186 191494
rect 407422 191258 407464 191494
rect 407144 184494 407464 191258
rect 407144 184258 407186 184494
rect 407422 184258 407464 184494
rect 407144 177494 407464 184258
rect 407144 177258 407186 177494
rect 407422 177258 407464 177494
rect 407144 170494 407464 177258
rect 407144 170258 407186 170494
rect 407422 170258 407464 170494
rect 407144 163494 407464 170258
rect 407144 163258 407186 163494
rect 407422 163258 407464 163494
rect 407144 156494 407464 163258
rect 407144 156258 407186 156494
rect 407422 156258 407464 156494
rect 407144 149494 407464 156258
rect 407144 149258 407186 149494
rect 407422 149258 407464 149494
rect 407144 142494 407464 149258
rect 407144 142258 407186 142494
rect 407422 142258 407464 142494
rect 407144 135494 407464 142258
rect 407144 135258 407186 135494
rect 407422 135258 407464 135494
rect 407144 128494 407464 135258
rect 407144 128258 407186 128494
rect 407422 128258 407464 128494
rect 407144 121494 407464 128258
rect 407144 121258 407186 121494
rect 407422 121258 407464 121494
rect 407144 114494 407464 121258
rect 407144 114258 407186 114494
rect 407422 114258 407464 114494
rect 407144 107494 407464 114258
rect 407144 107258 407186 107494
rect 407422 107258 407464 107494
rect 407144 100494 407464 107258
rect 407144 100258 407186 100494
rect 407422 100258 407464 100494
rect 407144 93494 407464 100258
rect 407144 93258 407186 93494
rect 407422 93258 407464 93494
rect 407144 86494 407464 93258
rect 407144 86258 407186 86494
rect 407422 86258 407464 86494
rect 407144 79494 407464 86258
rect 407144 79258 407186 79494
rect 407422 79258 407464 79494
rect 407144 72494 407464 79258
rect 407144 72258 407186 72494
rect 407422 72258 407464 72494
rect 407144 65494 407464 72258
rect 407144 65258 407186 65494
rect 407422 65258 407464 65494
rect 407144 58494 407464 65258
rect 407144 58258 407186 58494
rect 407422 58258 407464 58494
rect 407144 51494 407464 58258
rect 407144 51258 407186 51494
rect 407422 51258 407464 51494
rect 407144 44494 407464 51258
rect 407144 44258 407186 44494
rect 407422 44258 407464 44494
rect 407144 37494 407464 44258
rect 407144 37258 407186 37494
rect 407422 37258 407464 37494
rect 407144 30494 407464 37258
rect 407144 30258 407186 30494
rect 407422 30258 407464 30494
rect 407144 23494 407464 30258
rect 407144 23258 407186 23494
rect 407422 23258 407464 23494
rect 407144 16494 407464 23258
rect 407144 16258 407186 16494
rect 407422 16258 407464 16494
rect 407144 9494 407464 16258
rect 407144 9258 407186 9494
rect 407422 9258 407464 9494
rect 407144 2494 407464 9258
rect 407144 2258 407186 2494
rect 407422 2258 407464 2494
rect 407144 -746 407464 2258
rect 407144 -982 407186 -746
rect 407422 -982 407464 -746
rect 407144 -1066 407464 -982
rect 407144 -1302 407186 -1066
rect 407422 -1302 407464 -1066
rect 407144 -2294 407464 -1302
rect 408876 706198 409196 706230
rect 408876 705962 408918 706198
rect 409154 705962 409196 706198
rect 408876 705878 409196 705962
rect 408876 705642 408918 705878
rect 409154 705642 409196 705878
rect 408876 696561 409196 705642
rect 408876 696325 408918 696561
rect 409154 696325 409196 696561
rect 408876 689561 409196 696325
rect 408876 689325 408918 689561
rect 409154 689325 409196 689561
rect 408876 682561 409196 689325
rect 408876 682325 408918 682561
rect 409154 682325 409196 682561
rect 408876 675561 409196 682325
rect 408876 675325 408918 675561
rect 409154 675325 409196 675561
rect 408876 668561 409196 675325
rect 408876 668325 408918 668561
rect 409154 668325 409196 668561
rect 408876 661561 409196 668325
rect 408876 661325 408918 661561
rect 409154 661325 409196 661561
rect 408876 654561 409196 661325
rect 408876 654325 408918 654561
rect 409154 654325 409196 654561
rect 408876 647561 409196 654325
rect 408876 647325 408918 647561
rect 409154 647325 409196 647561
rect 408876 640561 409196 647325
rect 408876 640325 408918 640561
rect 409154 640325 409196 640561
rect 408876 633561 409196 640325
rect 408876 633325 408918 633561
rect 409154 633325 409196 633561
rect 408876 626561 409196 633325
rect 408876 626325 408918 626561
rect 409154 626325 409196 626561
rect 408876 619561 409196 626325
rect 408876 619325 408918 619561
rect 409154 619325 409196 619561
rect 408876 612561 409196 619325
rect 408876 612325 408918 612561
rect 409154 612325 409196 612561
rect 408876 605561 409196 612325
rect 408876 605325 408918 605561
rect 409154 605325 409196 605561
rect 408876 598561 409196 605325
rect 408876 598325 408918 598561
rect 409154 598325 409196 598561
rect 408876 591561 409196 598325
rect 408876 591325 408918 591561
rect 409154 591325 409196 591561
rect 408876 584561 409196 591325
rect 408876 584325 408918 584561
rect 409154 584325 409196 584561
rect 408876 577561 409196 584325
rect 408876 577325 408918 577561
rect 409154 577325 409196 577561
rect 408876 570561 409196 577325
rect 408876 570325 408918 570561
rect 409154 570325 409196 570561
rect 408876 563561 409196 570325
rect 408876 563325 408918 563561
rect 409154 563325 409196 563561
rect 408876 556561 409196 563325
rect 408876 556325 408918 556561
rect 409154 556325 409196 556561
rect 408876 549561 409196 556325
rect 408876 549325 408918 549561
rect 409154 549325 409196 549561
rect 408876 542561 409196 549325
rect 408876 542325 408918 542561
rect 409154 542325 409196 542561
rect 408876 535561 409196 542325
rect 408876 535325 408918 535561
rect 409154 535325 409196 535561
rect 408876 528561 409196 535325
rect 408876 528325 408918 528561
rect 409154 528325 409196 528561
rect 408876 521561 409196 528325
rect 408876 521325 408918 521561
rect 409154 521325 409196 521561
rect 408876 514561 409196 521325
rect 408876 514325 408918 514561
rect 409154 514325 409196 514561
rect 408876 507561 409196 514325
rect 408876 507325 408918 507561
rect 409154 507325 409196 507561
rect 408876 500561 409196 507325
rect 408876 500325 408918 500561
rect 409154 500325 409196 500561
rect 408876 493561 409196 500325
rect 408876 493325 408918 493561
rect 409154 493325 409196 493561
rect 408876 486561 409196 493325
rect 408876 486325 408918 486561
rect 409154 486325 409196 486561
rect 408876 479561 409196 486325
rect 408876 479325 408918 479561
rect 409154 479325 409196 479561
rect 408876 472561 409196 479325
rect 408876 472325 408918 472561
rect 409154 472325 409196 472561
rect 408876 465561 409196 472325
rect 408876 465325 408918 465561
rect 409154 465325 409196 465561
rect 408876 458561 409196 465325
rect 408876 458325 408918 458561
rect 409154 458325 409196 458561
rect 408876 451561 409196 458325
rect 408876 451325 408918 451561
rect 409154 451325 409196 451561
rect 408876 444561 409196 451325
rect 408876 444325 408918 444561
rect 409154 444325 409196 444561
rect 408876 437561 409196 444325
rect 408876 437325 408918 437561
rect 409154 437325 409196 437561
rect 408876 430561 409196 437325
rect 408876 430325 408918 430561
rect 409154 430325 409196 430561
rect 408876 423561 409196 430325
rect 408876 423325 408918 423561
rect 409154 423325 409196 423561
rect 408876 416561 409196 423325
rect 408876 416325 408918 416561
rect 409154 416325 409196 416561
rect 408876 409561 409196 416325
rect 408876 409325 408918 409561
rect 409154 409325 409196 409561
rect 408876 402561 409196 409325
rect 408876 402325 408918 402561
rect 409154 402325 409196 402561
rect 408876 395561 409196 402325
rect 408876 395325 408918 395561
rect 409154 395325 409196 395561
rect 408876 388561 409196 395325
rect 408876 388325 408918 388561
rect 409154 388325 409196 388561
rect 408876 381561 409196 388325
rect 408876 381325 408918 381561
rect 409154 381325 409196 381561
rect 408876 374561 409196 381325
rect 408876 374325 408918 374561
rect 409154 374325 409196 374561
rect 408876 367561 409196 374325
rect 408876 367325 408918 367561
rect 409154 367325 409196 367561
rect 408876 360561 409196 367325
rect 408876 360325 408918 360561
rect 409154 360325 409196 360561
rect 408876 353561 409196 360325
rect 408876 353325 408918 353561
rect 409154 353325 409196 353561
rect 408876 346561 409196 353325
rect 408876 346325 408918 346561
rect 409154 346325 409196 346561
rect 408876 339561 409196 346325
rect 408876 339325 408918 339561
rect 409154 339325 409196 339561
rect 408876 332561 409196 339325
rect 408876 332325 408918 332561
rect 409154 332325 409196 332561
rect 408876 325561 409196 332325
rect 408876 325325 408918 325561
rect 409154 325325 409196 325561
rect 408876 318561 409196 325325
rect 408876 318325 408918 318561
rect 409154 318325 409196 318561
rect 408876 311561 409196 318325
rect 408876 311325 408918 311561
rect 409154 311325 409196 311561
rect 408876 304561 409196 311325
rect 408876 304325 408918 304561
rect 409154 304325 409196 304561
rect 408876 297561 409196 304325
rect 408876 297325 408918 297561
rect 409154 297325 409196 297561
rect 408876 290561 409196 297325
rect 408876 290325 408918 290561
rect 409154 290325 409196 290561
rect 408876 283561 409196 290325
rect 408876 283325 408918 283561
rect 409154 283325 409196 283561
rect 408876 276561 409196 283325
rect 408876 276325 408918 276561
rect 409154 276325 409196 276561
rect 408876 269561 409196 276325
rect 408876 269325 408918 269561
rect 409154 269325 409196 269561
rect 408876 262561 409196 269325
rect 408876 262325 408918 262561
rect 409154 262325 409196 262561
rect 408876 255561 409196 262325
rect 408876 255325 408918 255561
rect 409154 255325 409196 255561
rect 408876 248561 409196 255325
rect 408876 248325 408918 248561
rect 409154 248325 409196 248561
rect 408876 241561 409196 248325
rect 408876 241325 408918 241561
rect 409154 241325 409196 241561
rect 408876 234561 409196 241325
rect 408876 234325 408918 234561
rect 409154 234325 409196 234561
rect 408876 227561 409196 234325
rect 408876 227325 408918 227561
rect 409154 227325 409196 227561
rect 408876 220561 409196 227325
rect 408876 220325 408918 220561
rect 409154 220325 409196 220561
rect 408876 213561 409196 220325
rect 408876 213325 408918 213561
rect 409154 213325 409196 213561
rect 408876 206561 409196 213325
rect 408876 206325 408918 206561
rect 409154 206325 409196 206561
rect 408876 199561 409196 206325
rect 408876 199325 408918 199561
rect 409154 199325 409196 199561
rect 408876 192561 409196 199325
rect 408876 192325 408918 192561
rect 409154 192325 409196 192561
rect 408876 185561 409196 192325
rect 408876 185325 408918 185561
rect 409154 185325 409196 185561
rect 408876 178561 409196 185325
rect 408876 178325 408918 178561
rect 409154 178325 409196 178561
rect 408876 171561 409196 178325
rect 408876 171325 408918 171561
rect 409154 171325 409196 171561
rect 408876 164561 409196 171325
rect 408876 164325 408918 164561
rect 409154 164325 409196 164561
rect 408876 157561 409196 164325
rect 408876 157325 408918 157561
rect 409154 157325 409196 157561
rect 408876 150561 409196 157325
rect 408876 150325 408918 150561
rect 409154 150325 409196 150561
rect 408876 143561 409196 150325
rect 408876 143325 408918 143561
rect 409154 143325 409196 143561
rect 408876 136561 409196 143325
rect 408876 136325 408918 136561
rect 409154 136325 409196 136561
rect 408876 129561 409196 136325
rect 408876 129325 408918 129561
rect 409154 129325 409196 129561
rect 408876 122561 409196 129325
rect 408876 122325 408918 122561
rect 409154 122325 409196 122561
rect 408876 115561 409196 122325
rect 408876 115325 408918 115561
rect 409154 115325 409196 115561
rect 408876 108561 409196 115325
rect 408876 108325 408918 108561
rect 409154 108325 409196 108561
rect 408876 101561 409196 108325
rect 408876 101325 408918 101561
rect 409154 101325 409196 101561
rect 408876 94561 409196 101325
rect 408876 94325 408918 94561
rect 409154 94325 409196 94561
rect 408876 87561 409196 94325
rect 408876 87325 408918 87561
rect 409154 87325 409196 87561
rect 408876 80561 409196 87325
rect 408876 80325 408918 80561
rect 409154 80325 409196 80561
rect 408876 73561 409196 80325
rect 408876 73325 408918 73561
rect 409154 73325 409196 73561
rect 408876 66561 409196 73325
rect 408876 66325 408918 66561
rect 409154 66325 409196 66561
rect 408876 59561 409196 66325
rect 408876 59325 408918 59561
rect 409154 59325 409196 59561
rect 408876 52561 409196 59325
rect 408876 52325 408918 52561
rect 409154 52325 409196 52561
rect 408876 45561 409196 52325
rect 408876 45325 408918 45561
rect 409154 45325 409196 45561
rect 408876 38561 409196 45325
rect 408876 38325 408918 38561
rect 409154 38325 409196 38561
rect 408876 31561 409196 38325
rect 408876 31325 408918 31561
rect 409154 31325 409196 31561
rect 408876 24561 409196 31325
rect 408876 24325 408918 24561
rect 409154 24325 409196 24561
rect 408876 17561 409196 24325
rect 408876 17325 408918 17561
rect 409154 17325 409196 17561
rect 408876 10561 409196 17325
rect 408876 10325 408918 10561
rect 409154 10325 409196 10561
rect 408876 3561 409196 10325
rect 408876 3325 408918 3561
rect 409154 3325 409196 3561
rect 408876 -1706 409196 3325
rect 408876 -1942 408918 -1706
rect 409154 -1942 409196 -1706
rect 408876 -2026 409196 -1942
rect 408876 -2262 408918 -2026
rect 409154 -2262 409196 -2026
rect 408876 -2294 409196 -2262
rect 414144 705238 414464 706230
rect 414144 705002 414186 705238
rect 414422 705002 414464 705238
rect 414144 704918 414464 705002
rect 414144 704682 414186 704918
rect 414422 704682 414464 704918
rect 414144 695494 414464 704682
rect 414144 695258 414186 695494
rect 414422 695258 414464 695494
rect 414144 688494 414464 695258
rect 414144 688258 414186 688494
rect 414422 688258 414464 688494
rect 414144 681494 414464 688258
rect 414144 681258 414186 681494
rect 414422 681258 414464 681494
rect 414144 674494 414464 681258
rect 414144 674258 414186 674494
rect 414422 674258 414464 674494
rect 414144 667494 414464 674258
rect 414144 667258 414186 667494
rect 414422 667258 414464 667494
rect 414144 660494 414464 667258
rect 414144 660258 414186 660494
rect 414422 660258 414464 660494
rect 414144 653494 414464 660258
rect 414144 653258 414186 653494
rect 414422 653258 414464 653494
rect 414144 646494 414464 653258
rect 414144 646258 414186 646494
rect 414422 646258 414464 646494
rect 414144 639494 414464 646258
rect 414144 639258 414186 639494
rect 414422 639258 414464 639494
rect 414144 632494 414464 639258
rect 414144 632258 414186 632494
rect 414422 632258 414464 632494
rect 414144 625494 414464 632258
rect 414144 625258 414186 625494
rect 414422 625258 414464 625494
rect 414144 618494 414464 625258
rect 414144 618258 414186 618494
rect 414422 618258 414464 618494
rect 414144 611494 414464 618258
rect 414144 611258 414186 611494
rect 414422 611258 414464 611494
rect 414144 604494 414464 611258
rect 414144 604258 414186 604494
rect 414422 604258 414464 604494
rect 414144 597494 414464 604258
rect 414144 597258 414186 597494
rect 414422 597258 414464 597494
rect 414144 590494 414464 597258
rect 414144 590258 414186 590494
rect 414422 590258 414464 590494
rect 414144 583494 414464 590258
rect 414144 583258 414186 583494
rect 414422 583258 414464 583494
rect 414144 576494 414464 583258
rect 414144 576258 414186 576494
rect 414422 576258 414464 576494
rect 414144 569494 414464 576258
rect 414144 569258 414186 569494
rect 414422 569258 414464 569494
rect 414144 562494 414464 569258
rect 414144 562258 414186 562494
rect 414422 562258 414464 562494
rect 414144 555494 414464 562258
rect 414144 555258 414186 555494
rect 414422 555258 414464 555494
rect 414144 548494 414464 555258
rect 414144 548258 414186 548494
rect 414422 548258 414464 548494
rect 414144 541494 414464 548258
rect 414144 541258 414186 541494
rect 414422 541258 414464 541494
rect 414144 534494 414464 541258
rect 414144 534258 414186 534494
rect 414422 534258 414464 534494
rect 414144 527494 414464 534258
rect 414144 527258 414186 527494
rect 414422 527258 414464 527494
rect 414144 520494 414464 527258
rect 414144 520258 414186 520494
rect 414422 520258 414464 520494
rect 414144 513494 414464 520258
rect 414144 513258 414186 513494
rect 414422 513258 414464 513494
rect 414144 506494 414464 513258
rect 414144 506258 414186 506494
rect 414422 506258 414464 506494
rect 414144 499494 414464 506258
rect 414144 499258 414186 499494
rect 414422 499258 414464 499494
rect 414144 492494 414464 499258
rect 414144 492258 414186 492494
rect 414422 492258 414464 492494
rect 414144 485494 414464 492258
rect 414144 485258 414186 485494
rect 414422 485258 414464 485494
rect 414144 478494 414464 485258
rect 414144 478258 414186 478494
rect 414422 478258 414464 478494
rect 414144 471494 414464 478258
rect 414144 471258 414186 471494
rect 414422 471258 414464 471494
rect 414144 464494 414464 471258
rect 414144 464258 414186 464494
rect 414422 464258 414464 464494
rect 414144 457494 414464 464258
rect 414144 457258 414186 457494
rect 414422 457258 414464 457494
rect 414144 450494 414464 457258
rect 414144 450258 414186 450494
rect 414422 450258 414464 450494
rect 414144 443494 414464 450258
rect 414144 443258 414186 443494
rect 414422 443258 414464 443494
rect 414144 436494 414464 443258
rect 414144 436258 414186 436494
rect 414422 436258 414464 436494
rect 414144 429494 414464 436258
rect 414144 429258 414186 429494
rect 414422 429258 414464 429494
rect 414144 422494 414464 429258
rect 414144 422258 414186 422494
rect 414422 422258 414464 422494
rect 414144 415494 414464 422258
rect 414144 415258 414186 415494
rect 414422 415258 414464 415494
rect 414144 408494 414464 415258
rect 414144 408258 414186 408494
rect 414422 408258 414464 408494
rect 414144 401494 414464 408258
rect 414144 401258 414186 401494
rect 414422 401258 414464 401494
rect 414144 394494 414464 401258
rect 414144 394258 414186 394494
rect 414422 394258 414464 394494
rect 414144 387494 414464 394258
rect 414144 387258 414186 387494
rect 414422 387258 414464 387494
rect 414144 380494 414464 387258
rect 414144 380258 414186 380494
rect 414422 380258 414464 380494
rect 414144 373494 414464 380258
rect 414144 373258 414186 373494
rect 414422 373258 414464 373494
rect 414144 366494 414464 373258
rect 414144 366258 414186 366494
rect 414422 366258 414464 366494
rect 414144 359494 414464 366258
rect 414144 359258 414186 359494
rect 414422 359258 414464 359494
rect 414144 352494 414464 359258
rect 414144 352258 414186 352494
rect 414422 352258 414464 352494
rect 414144 345494 414464 352258
rect 414144 345258 414186 345494
rect 414422 345258 414464 345494
rect 414144 338494 414464 345258
rect 414144 338258 414186 338494
rect 414422 338258 414464 338494
rect 414144 331494 414464 338258
rect 414144 331258 414186 331494
rect 414422 331258 414464 331494
rect 414144 324494 414464 331258
rect 414144 324258 414186 324494
rect 414422 324258 414464 324494
rect 414144 317494 414464 324258
rect 414144 317258 414186 317494
rect 414422 317258 414464 317494
rect 414144 310494 414464 317258
rect 414144 310258 414186 310494
rect 414422 310258 414464 310494
rect 414144 303494 414464 310258
rect 414144 303258 414186 303494
rect 414422 303258 414464 303494
rect 414144 296494 414464 303258
rect 414144 296258 414186 296494
rect 414422 296258 414464 296494
rect 414144 289494 414464 296258
rect 414144 289258 414186 289494
rect 414422 289258 414464 289494
rect 414144 282494 414464 289258
rect 414144 282258 414186 282494
rect 414422 282258 414464 282494
rect 414144 275494 414464 282258
rect 414144 275258 414186 275494
rect 414422 275258 414464 275494
rect 414144 268494 414464 275258
rect 414144 268258 414186 268494
rect 414422 268258 414464 268494
rect 414144 261494 414464 268258
rect 414144 261258 414186 261494
rect 414422 261258 414464 261494
rect 414144 254494 414464 261258
rect 414144 254258 414186 254494
rect 414422 254258 414464 254494
rect 414144 247494 414464 254258
rect 414144 247258 414186 247494
rect 414422 247258 414464 247494
rect 414144 240494 414464 247258
rect 414144 240258 414186 240494
rect 414422 240258 414464 240494
rect 414144 233494 414464 240258
rect 414144 233258 414186 233494
rect 414422 233258 414464 233494
rect 414144 226494 414464 233258
rect 414144 226258 414186 226494
rect 414422 226258 414464 226494
rect 414144 219494 414464 226258
rect 414144 219258 414186 219494
rect 414422 219258 414464 219494
rect 414144 212494 414464 219258
rect 414144 212258 414186 212494
rect 414422 212258 414464 212494
rect 414144 205494 414464 212258
rect 414144 205258 414186 205494
rect 414422 205258 414464 205494
rect 414144 198494 414464 205258
rect 414144 198258 414186 198494
rect 414422 198258 414464 198494
rect 414144 191494 414464 198258
rect 414144 191258 414186 191494
rect 414422 191258 414464 191494
rect 414144 184494 414464 191258
rect 414144 184258 414186 184494
rect 414422 184258 414464 184494
rect 414144 177494 414464 184258
rect 414144 177258 414186 177494
rect 414422 177258 414464 177494
rect 414144 170494 414464 177258
rect 414144 170258 414186 170494
rect 414422 170258 414464 170494
rect 414144 163494 414464 170258
rect 414144 163258 414186 163494
rect 414422 163258 414464 163494
rect 414144 156494 414464 163258
rect 414144 156258 414186 156494
rect 414422 156258 414464 156494
rect 414144 149494 414464 156258
rect 414144 149258 414186 149494
rect 414422 149258 414464 149494
rect 414144 142494 414464 149258
rect 414144 142258 414186 142494
rect 414422 142258 414464 142494
rect 414144 135494 414464 142258
rect 414144 135258 414186 135494
rect 414422 135258 414464 135494
rect 414144 128494 414464 135258
rect 414144 128258 414186 128494
rect 414422 128258 414464 128494
rect 414144 121494 414464 128258
rect 414144 121258 414186 121494
rect 414422 121258 414464 121494
rect 414144 114494 414464 121258
rect 414144 114258 414186 114494
rect 414422 114258 414464 114494
rect 414144 107494 414464 114258
rect 414144 107258 414186 107494
rect 414422 107258 414464 107494
rect 414144 100494 414464 107258
rect 414144 100258 414186 100494
rect 414422 100258 414464 100494
rect 414144 93494 414464 100258
rect 414144 93258 414186 93494
rect 414422 93258 414464 93494
rect 414144 86494 414464 93258
rect 414144 86258 414186 86494
rect 414422 86258 414464 86494
rect 414144 79494 414464 86258
rect 414144 79258 414186 79494
rect 414422 79258 414464 79494
rect 414144 72494 414464 79258
rect 414144 72258 414186 72494
rect 414422 72258 414464 72494
rect 414144 65494 414464 72258
rect 414144 65258 414186 65494
rect 414422 65258 414464 65494
rect 414144 58494 414464 65258
rect 414144 58258 414186 58494
rect 414422 58258 414464 58494
rect 414144 51494 414464 58258
rect 414144 51258 414186 51494
rect 414422 51258 414464 51494
rect 414144 44494 414464 51258
rect 414144 44258 414186 44494
rect 414422 44258 414464 44494
rect 414144 37494 414464 44258
rect 414144 37258 414186 37494
rect 414422 37258 414464 37494
rect 414144 30494 414464 37258
rect 414144 30258 414186 30494
rect 414422 30258 414464 30494
rect 414144 23494 414464 30258
rect 414144 23258 414186 23494
rect 414422 23258 414464 23494
rect 414144 16494 414464 23258
rect 414144 16258 414186 16494
rect 414422 16258 414464 16494
rect 414144 9494 414464 16258
rect 414144 9258 414186 9494
rect 414422 9258 414464 9494
rect 414144 2494 414464 9258
rect 414144 2258 414186 2494
rect 414422 2258 414464 2494
rect 414144 -746 414464 2258
rect 414144 -982 414186 -746
rect 414422 -982 414464 -746
rect 414144 -1066 414464 -982
rect 414144 -1302 414186 -1066
rect 414422 -1302 414464 -1066
rect 414144 -2294 414464 -1302
rect 415876 706198 416196 706230
rect 415876 705962 415918 706198
rect 416154 705962 416196 706198
rect 415876 705878 416196 705962
rect 415876 705642 415918 705878
rect 416154 705642 416196 705878
rect 415876 696561 416196 705642
rect 415876 696325 415918 696561
rect 416154 696325 416196 696561
rect 415876 689561 416196 696325
rect 415876 689325 415918 689561
rect 416154 689325 416196 689561
rect 415876 682561 416196 689325
rect 415876 682325 415918 682561
rect 416154 682325 416196 682561
rect 415876 675561 416196 682325
rect 415876 675325 415918 675561
rect 416154 675325 416196 675561
rect 415876 668561 416196 675325
rect 415876 668325 415918 668561
rect 416154 668325 416196 668561
rect 415876 661561 416196 668325
rect 415876 661325 415918 661561
rect 416154 661325 416196 661561
rect 415876 654561 416196 661325
rect 415876 654325 415918 654561
rect 416154 654325 416196 654561
rect 415876 647561 416196 654325
rect 415876 647325 415918 647561
rect 416154 647325 416196 647561
rect 415876 640561 416196 647325
rect 415876 640325 415918 640561
rect 416154 640325 416196 640561
rect 415876 633561 416196 640325
rect 415876 633325 415918 633561
rect 416154 633325 416196 633561
rect 415876 626561 416196 633325
rect 415876 626325 415918 626561
rect 416154 626325 416196 626561
rect 415876 619561 416196 626325
rect 415876 619325 415918 619561
rect 416154 619325 416196 619561
rect 415876 612561 416196 619325
rect 415876 612325 415918 612561
rect 416154 612325 416196 612561
rect 415876 605561 416196 612325
rect 415876 605325 415918 605561
rect 416154 605325 416196 605561
rect 415876 598561 416196 605325
rect 415876 598325 415918 598561
rect 416154 598325 416196 598561
rect 415876 591561 416196 598325
rect 415876 591325 415918 591561
rect 416154 591325 416196 591561
rect 415876 584561 416196 591325
rect 415876 584325 415918 584561
rect 416154 584325 416196 584561
rect 415876 577561 416196 584325
rect 415876 577325 415918 577561
rect 416154 577325 416196 577561
rect 415876 570561 416196 577325
rect 415876 570325 415918 570561
rect 416154 570325 416196 570561
rect 415876 563561 416196 570325
rect 415876 563325 415918 563561
rect 416154 563325 416196 563561
rect 415876 556561 416196 563325
rect 415876 556325 415918 556561
rect 416154 556325 416196 556561
rect 415876 549561 416196 556325
rect 415876 549325 415918 549561
rect 416154 549325 416196 549561
rect 415876 542561 416196 549325
rect 415876 542325 415918 542561
rect 416154 542325 416196 542561
rect 415876 535561 416196 542325
rect 415876 535325 415918 535561
rect 416154 535325 416196 535561
rect 415876 528561 416196 535325
rect 415876 528325 415918 528561
rect 416154 528325 416196 528561
rect 415876 521561 416196 528325
rect 415876 521325 415918 521561
rect 416154 521325 416196 521561
rect 415876 514561 416196 521325
rect 415876 514325 415918 514561
rect 416154 514325 416196 514561
rect 415876 507561 416196 514325
rect 415876 507325 415918 507561
rect 416154 507325 416196 507561
rect 415876 500561 416196 507325
rect 415876 500325 415918 500561
rect 416154 500325 416196 500561
rect 415876 493561 416196 500325
rect 415876 493325 415918 493561
rect 416154 493325 416196 493561
rect 415876 486561 416196 493325
rect 415876 486325 415918 486561
rect 416154 486325 416196 486561
rect 415876 479561 416196 486325
rect 415876 479325 415918 479561
rect 416154 479325 416196 479561
rect 415876 472561 416196 479325
rect 415876 472325 415918 472561
rect 416154 472325 416196 472561
rect 415876 465561 416196 472325
rect 415876 465325 415918 465561
rect 416154 465325 416196 465561
rect 415876 458561 416196 465325
rect 415876 458325 415918 458561
rect 416154 458325 416196 458561
rect 415876 451561 416196 458325
rect 415876 451325 415918 451561
rect 416154 451325 416196 451561
rect 415876 444561 416196 451325
rect 415876 444325 415918 444561
rect 416154 444325 416196 444561
rect 415876 437561 416196 444325
rect 415876 437325 415918 437561
rect 416154 437325 416196 437561
rect 415876 430561 416196 437325
rect 415876 430325 415918 430561
rect 416154 430325 416196 430561
rect 415876 423561 416196 430325
rect 415876 423325 415918 423561
rect 416154 423325 416196 423561
rect 415876 416561 416196 423325
rect 415876 416325 415918 416561
rect 416154 416325 416196 416561
rect 415876 409561 416196 416325
rect 415876 409325 415918 409561
rect 416154 409325 416196 409561
rect 415876 402561 416196 409325
rect 415876 402325 415918 402561
rect 416154 402325 416196 402561
rect 415876 395561 416196 402325
rect 415876 395325 415918 395561
rect 416154 395325 416196 395561
rect 415876 388561 416196 395325
rect 415876 388325 415918 388561
rect 416154 388325 416196 388561
rect 415876 381561 416196 388325
rect 415876 381325 415918 381561
rect 416154 381325 416196 381561
rect 415876 374561 416196 381325
rect 415876 374325 415918 374561
rect 416154 374325 416196 374561
rect 415876 367561 416196 374325
rect 415876 367325 415918 367561
rect 416154 367325 416196 367561
rect 415876 360561 416196 367325
rect 415876 360325 415918 360561
rect 416154 360325 416196 360561
rect 415876 353561 416196 360325
rect 415876 353325 415918 353561
rect 416154 353325 416196 353561
rect 415876 346561 416196 353325
rect 415876 346325 415918 346561
rect 416154 346325 416196 346561
rect 415876 339561 416196 346325
rect 415876 339325 415918 339561
rect 416154 339325 416196 339561
rect 415876 332561 416196 339325
rect 415876 332325 415918 332561
rect 416154 332325 416196 332561
rect 415876 325561 416196 332325
rect 415876 325325 415918 325561
rect 416154 325325 416196 325561
rect 415876 318561 416196 325325
rect 415876 318325 415918 318561
rect 416154 318325 416196 318561
rect 415876 311561 416196 318325
rect 415876 311325 415918 311561
rect 416154 311325 416196 311561
rect 415876 304561 416196 311325
rect 415876 304325 415918 304561
rect 416154 304325 416196 304561
rect 415876 297561 416196 304325
rect 415876 297325 415918 297561
rect 416154 297325 416196 297561
rect 415876 290561 416196 297325
rect 415876 290325 415918 290561
rect 416154 290325 416196 290561
rect 415876 283561 416196 290325
rect 415876 283325 415918 283561
rect 416154 283325 416196 283561
rect 415876 276561 416196 283325
rect 415876 276325 415918 276561
rect 416154 276325 416196 276561
rect 415876 269561 416196 276325
rect 415876 269325 415918 269561
rect 416154 269325 416196 269561
rect 415876 262561 416196 269325
rect 415876 262325 415918 262561
rect 416154 262325 416196 262561
rect 415876 255561 416196 262325
rect 415876 255325 415918 255561
rect 416154 255325 416196 255561
rect 415876 248561 416196 255325
rect 415876 248325 415918 248561
rect 416154 248325 416196 248561
rect 415876 241561 416196 248325
rect 415876 241325 415918 241561
rect 416154 241325 416196 241561
rect 415876 234561 416196 241325
rect 415876 234325 415918 234561
rect 416154 234325 416196 234561
rect 415876 227561 416196 234325
rect 415876 227325 415918 227561
rect 416154 227325 416196 227561
rect 415876 220561 416196 227325
rect 415876 220325 415918 220561
rect 416154 220325 416196 220561
rect 415876 213561 416196 220325
rect 415876 213325 415918 213561
rect 416154 213325 416196 213561
rect 415876 206561 416196 213325
rect 415876 206325 415918 206561
rect 416154 206325 416196 206561
rect 415876 199561 416196 206325
rect 415876 199325 415918 199561
rect 416154 199325 416196 199561
rect 415876 192561 416196 199325
rect 415876 192325 415918 192561
rect 416154 192325 416196 192561
rect 415876 185561 416196 192325
rect 415876 185325 415918 185561
rect 416154 185325 416196 185561
rect 415876 178561 416196 185325
rect 415876 178325 415918 178561
rect 416154 178325 416196 178561
rect 415876 171561 416196 178325
rect 415876 171325 415918 171561
rect 416154 171325 416196 171561
rect 415876 164561 416196 171325
rect 415876 164325 415918 164561
rect 416154 164325 416196 164561
rect 415876 157561 416196 164325
rect 415876 157325 415918 157561
rect 416154 157325 416196 157561
rect 415876 150561 416196 157325
rect 415876 150325 415918 150561
rect 416154 150325 416196 150561
rect 415876 143561 416196 150325
rect 415876 143325 415918 143561
rect 416154 143325 416196 143561
rect 415876 136561 416196 143325
rect 415876 136325 415918 136561
rect 416154 136325 416196 136561
rect 415876 129561 416196 136325
rect 415876 129325 415918 129561
rect 416154 129325 416196 129561
rect 415876 122561 416196 129325
rect 415876 122325 415918 122561
rect 416154 122325 416196 122561
rect 415876 115561 416196 122325
rect 415876 115325 415918 115561
rect 416154 115325 416196 115561
rect 415876 108561 416196 115325
rect 415876 108325 415918 108561
rect 416154 108325 416196 108561
rect 415876 101561 416196 108325
rect 415876 101325 415918 101561
rect 416154 101325 416196 101561
rect 415876 94561 416196 101325
rect 415876 94325 415918 94561
rect 416154 94325 416196 94561
rect 415876 87561 416196 94325
rect 415876 87325 415918 87561
rect 416154 87325 416196 87561
rect 415876 80561 416196 87325
rect 415876 80325 415918 80561
rect 416154 80325 416196 80561
rect 415876 73561 416196 80325
rect 415876 73325 415918 73561
rect 416154 73325 416196 73561
rect 415876 66561 416196 73325
rect 415876 66325 415918 66561
rect 416154 66325 416196 66561
rect 415876 59561 416196 66325
rect 415876 59325 415918 59561
rect 416154 59325 416196 59561
rect 415876 52561 416196 59325
rect 415876 52325 415918 52561
rect 416154 52325 416196 52561
rect 415876 45561 416196 52325
rect 415876 45325 415918 45561
rect 416154 45325 416196 45561
rect 415876 38561 416196 45325
rect 415876 38325 415918 38561
rect 416154 38325 416196 38561
rect 415876 31561 416196 38325
rect 415876 31325 415918 31561
rect 416154 31325 416196 31561
rect 415876 24561 416196 31325
rect 415876 24325 415918 24561
rect 416154 24325 416196 24561
rect 415876 17561 416196 24325
rect 415876 17325 415918 17561
rect 416154 17325 416196 17561
rect 415876 10561 416196 17325
rect 415876 10325 415918 10561
rect 416154 10325 416196 10561
rect 415876 3561 416196 10325
rect 415876 3325 415918 3561
rect 416154 3325 416196 3561
rect 415876 -1706 416196 3325
rect 415876 -1942 415918 -1706
rect 416154 -1942 416196 -1706
rect 415876 -2026 416196 -1942
rect 415876 -2262 415918 -2026
rect 416154 -2262 416196 -2026
rect 415876 -2294 416196 -2262
rect 421144 705238 421464 706230
rect 421144 705002 421186 705238
rect 421422 705002 421464 705238
rect 421144 704918 421464 705002
rect 421144 704682 421186 704918
rect 421422 704682 421464 704918
rect 421144 695494 421464 704682
rect 421144 695258 421186 695494
rect 421422 695258 421464 695494
rect 421144 688494 421464 695258
rect 421144 688258 421186 688494
rect 421422 688258 421464 688494
rect 421144 681494 421464 688258
rect 421144 681258 421186 681494
rect 421422 681258 421464 681494
rect 421144 674494 421464 681258
rect 421144 674258 421186 674494
rect 421422 674258 421464 674494
rect 421144 667494 421464 674258
rect 421144 667258 421186 667494
rect 421422 667258 421464 667494
rect 421144 660494 421464 667258
rect 421144 660258 421186 660494
rect 421422 660258 421464 660494
rect 421144 653494 421464 660258
rect 421144 653258 421186 653494
rect 421422 653258 421464 653494
rect 421144 646494 421464 653258
rect 421144 646258 421186 646494
rect 421422 646258 421464 646494
rect 421144 639494 421464 646258
rect 421144 639258 421186 639494
rect 421422 639258 421464 639494
rect 421144 632494 421464 639258
rect 421144 632258 421186 632494
rect 421422 632258 421464 632494
rect 421144 625494 421464 632258
rect 421144 625258 421186 625494
rect 421422 625258 421464 625494
rect 421144 618494 421464 625258
rect 421144 618258 421186 618494
rect 421422 618258 421464 618494
rect 421144 611494 421464 618258
rect 421144 611258 421186 611494
rect 421422 611258 421464 611494
rect 421144 604494 421464 611258
rect 421144 604258 421186 604494
rect 421422 604258 421464 604494
rect 421144 597494 421464 604258
rect 421144 597258 421186 597494
rect 421422 597258 421464 597494
rect 421144 590494 421464 597258
rect 421144 590258 421186 590494
rect 421422 590258 421464 590494
rect 421144 583494 421464 590258
rect 421144 583258 421186 583494
rect 421422 583258 421464 583494
rect 421144 576494 421464 583258
rect 421144 576258 421186 576494
rect 421422 576258 421464 576494
rect 421144 569494 421464 576258
rect 421144 569258 421186 569494
rect 421422 569258 421464 569494
rect 421144 562494 421464 569258
rect 421144 562258 421186 562494
rect 421422 562258 421464 562494
rect 421144 555494 421464 562258
rect 421144 555258 421186 555494
rect 421422 555258 421464 555494
rect 421144 548494 421464 555258
rect 421144 548258 421186 548494
rect 421422 548258 421464 548494
rect 421144 541494 421464 548258
rect 421144 541258 421186 541494
rect 421422 541258 421464 541494
rect 421144 534494 421464 541258
rect 421144 534258 421186 534494
rect 421422 534258 421464 534494
rect 421144 527494 421464 534258
rect 421144 527258 421186 527494
rect 421422 527258 421464 527494
rect 421144 520494 421464 527258
rect 421144 520258 421186 520494
rect 421422 520258 421464 520494
rect 421144 513494 421464 520258
rect 421144 513258 421186 513494
rect 421422 513258 421464 513494
rect 421144 506494 421464 513258
rect 421144 506258 421186 506494
rect 421422 506258 421464 506494
rect 421144 499494 421464 506258
rect 421144 499258 421186 499494
rect 421422 499258 421464 499494
rect 421144 492494 421464 499258
rect 421144 492258 421186 492494
rect 421422 492258 421464 492494
rect 421144 485494 421464 492258
rect 421144 485258 421186 485494
rect 421422 485258 421464 485494
rect 421144 478494 421464 485258
rect 421144 478258 421186 478494
rect 421422 478258 421464 478494
rect 421144 471494 421464 478258
rect 421144 471258 421186 471494
rect 421422 471258 421464 471494
rect 421144 464494 421464 471258
rect 421144 464258 421186 464494
rect 421422 464258 421464 464494
rect 421144 457494 421464 464258
rect 421144 457258 421186 457494
rect 421422 457258 421464 457494
rect 421144 450494 421464 457258
rect 421144 450258 421186 450494
rect 421422 450258 421464 450494
rect 421144 443494 421464 450258
rect 421144 443258 421186 443494
rect 421422 443258 421464 443494
rect 421144 436494 421464 443258
rect 421144 436258 421186 436494
rect 421422 436258 421464 436494
rect 421144 429494 421464 436258
rect 421144 429258 421186 429494
rect 421422 429258 421464 429494
rect 421144 422494 421464 429258
rect 421144 422258 421186 422494
rect 421422 422258 421464 422494
rect 421144 415494 421464 422258
rect 421144 415258 421186 415494
rect 421422 415258 421464 415494
rect 421144 408494 421464 415258
rect 421144 408258 421186 408494
rect 421422 408258 421464 408494
rect 421144 401494 421464 408258
rect 421144 401258 421186 401494
rect 421422 401258 421464 401494
rect 421144 394494 421464 401258
rect 421144 394258 421186 394494
rect 421422 394258 421464 394494
rect 421144 387494 421464 394258
rect 421144 387258 421186 387494
rect 421422 387258 421464 387494
rect 421144 380494 421464 387258
rect 421144 380258 421186 380494
rect 421422 380258 421464 380494
rect 421144 373494 421464 380258
rect 421144 373258 421186 373494
rect 421422 373258 421464 373494
rect 421144 366494 421464 373258
rect 421144 366258 421186 366494
rect 421422 366258 421464 366494
rect 421144 359494 421464 366258
rect 421144 359258 421186 359494
rect 421422 359258 421464 359494
rect 421144 352494 421464 359258
rect 421144 352258 421186 352494
rect 421422 352258 421464 352494
rect 421144 345494 421464 352258
rect 421144 345258 421186 345494
rect 421422 345258 421464 345494
rect 421144 338494 421464 345258
rect 421144 338258 421186 338494
rect 421422 338258 421464 338494
rect 421144 331494 421464 338258
rect 421144 331258 421186 331494
rect 421422 331258 421464 331494
rect 421144 324494 421464 331258
rect 421144 324258 421186 324494
rect 421422 324258 421464 324494
rect 421144 317494 421464 324258
rect 421144 317258 421186 317494
rect 421422 317258 421464 317494
rect 421144 310494 421464 317258
rect 421144 310258 421186 310494
rect 421422 310258 421464 310494
rect 421144 303494 421464 310258
rect 421144 303258 421186 303494
rect 421422 303258 421464 303494
rect 421144 296494 421464 303258
rect 421144 296258 421186 296494
rect 421422 296258 421464 296494
rect 421144 289494 421464 296258
rect 421144 289258 421186 289494
rect 421422 289258 421464 289494
rect 421144 282494 421464 289258
rect 421144 282258 421186 282494
rect 421422 282258 421464 282494
rect 421144 275494 421464 282258
rect 421144 275258 421186 275494
rect 421422 275258 421464 275494
rect 421144 268494 421464 275258
rect 421144 268258 421186 268494
rect 421422 268258 421464 268494
rect 421144 261494 421464 268258
rect 421144 261258 421186 261494
rect 421422 261258 421464 261494
rect 421144 254494 421464 261258
rect 421144 254258 421186 254494
rect 421422 254258 421464 254494
rect 421144 247494 421464 254258
rect 421144 247258 421186 247494
rect 421422 247258 421464 247494
rect 421144 240494 421464 247258
rect 421144 240258 421186 240494
rect 421422 240258 421464 240494
rect 421144 233494 421464 240258
rect 421144 233258 421186 233494
rect 421422 233258 421464 233494
rect 421144 226494 421464 233258
rect 421144 226258 421186 226494
rect 421422 226258 421464 226494
rect 421144 219494 421464 226258
rect 421144 219258 421186 219494
rect 421422 219258 421464 219494
rect 421144 212494 421464 219258
rect 421144 212258 421186 212494
rect 421422 212258 421464 212494
rect 421144 205494 421464 212258
rect 421144 205258 421186 205494
rect 421422 205258 421464 205494
rect 421144 198494 421464 205258
rect 421144 198258 421186 198494
rect 421422 198258 421464 198494
rect 421144 191494 421464 198258
rect 421144 191258 421186 191494
rect 421422 191258 421464 191494
rect 421144 184494 421464 191258
rect 421144 184258 421186 184494
rect 421422 184258 421464 184494
rect 421144 177494 421464 184258
rect 421144 177258 421186 177494
rect 421422 177258 421464 177494
rect 421144 170494 421464 177258
rect 421144 170258 421186 170494
rect 421422 170258 421464 170494
rect 421144 163494 421464 170258
rect 421144 163258 421186 163494
rect 421422 163258 421464 163494
rect 421144 156494 421464 163258
rect 421144 156258 421186 156494
rect 421422 156258 421464 156494
rect 421144 149494 421464 156258
rect 421144 149258 421186 149494
rect 421422 149258 421464 149494
rect 421144 142494 421464 149258
rect 421144 142258 421186 142494
rect 421422 142258 421464 142494
rect 421144 135494 421464 142258
rect 421144 135258 421186 135494
rect 421422 135258 421464 135494
rect 421144 128494 421464 135258
rect 421144 128258 421186 128494
rect 421422 128258 421464 128494
rect 421144 121494 421464 128258
rect 421144 121258 421186 121494
rect 421422 121258 421464 121494
rect 421144 114494 421464 121258
rect 421144 114258 421186 114494
rect 421422 114258 421464 114494
rect 421144 107494 421464 114258
rect 421144 107258 421186 107494
rect 421422 107258 421464 107494
rect 421144 100494 421464 107258
rect 421144 100258 421186 100494
rect 421422 100258 421464 100494
rect 421144 93494 421464 100258
rect 421144 93258 421186 93494
rect 421422 93258 421464 93494
rect 421144 86494 421464 93258
rect 421144 86258 421186 86494
rect 421422 86258 421464 86494
rect 421144 79494 421464 86258
rect 421144 79258 421186 79494
rect 421422 79258 421464 79494
rect 421144 72494 421464 79258
rect 421144 72258 421186 72494
rect 421422 72258 421464 72494
rect 421144 65494 421464 72258
rect 421144 65258 421186 65494
rect 421422 65258 421464 65494
rect 421144 58494 421464 65258
rect 421144 58258 421186 58494
rect 421422 58258 421464 58494
rect 421144 51494 421464 58258
rect 421144 51258 421186 51494
rect 421422 51258 421464 51494
rect 421144 44494 421464 51258
rect 421144 44258 421186 44494
rect 421422 44258 421464 44494
rect 421144 37494 421464 44258
rect 421144 37258 421186 37494
rect 421422 37258 421464 37494
rect 421144 30494 421464 37258
rect 421144 30258 421186 30494
rect 421422 30258 421464 30494
rect 421144 23494 421464 30258
rect 421144 23258 421186 23494
rect 421422 23258 421464 23494
rect 421144 16494 421464 23258
rect 421144 16258 421186 16494
rect 421422 16258 421464 16494
rect 421144 9494 421464 16258
rect 421144 9258 421186 9494
rect 421422 9258 421464 9494
rect 421144 2494 421464 9258
rect 421144 2258 421186 2494
rect 421422 2258 421464 2494
rect 421144 -746 421464 2258
rect 421144 -982 421186 -746
rect 421422 -982 421464 -746
rect 421144 -1066 421464 -982
rect 421144 -1302 421186 -1066
rect 421422 -1302 421464 -1066
rect 421144 -2294 421464 -1302
rect 422876 706198 423196 706230
rect 422876 705962 422918 706198
rect 423154 705962 423196 706198
rect 422876 705878 423196 705962
rect 422876 705642 422918 705878
rect 423154 705642 423196 705878
rect 422876 696561 423196 705642
rect 422876 696325 422918 696561
rect 423154 696325 423196 696561
rect 422876 689561 423196 696325
rect 422876 689325 422918 689561
rect 423154 689325 423196 689561
rect 422876 682561 423196 689325
rect 422876 682325 422918 682561
rect 423154 682325 423196 682561
rect 422876 675561 423196 682325
rect 422876 675325 422918 675561
rect 423154 675325 423196 675561
rect 422876 668561 423196 675325
rect 422876 668325 422918 668561
rect 423154 668325 423196 668561
rect 422876 661561 423196 668325
rect 422876 661325 422918 661561
rect 423154 661325 423196 661561
rect 422876 654561 423196 661325
rect 422876 654325 422918 654561
rect 423154 654325 423196 654561
rect 422876 647561 423196 654325
rect 422876 647325 422918 647561
rect 423154 647325 423196 647561
rect 422876 640561 423196 647325
rect 422876 640325 422918 640561
rect 423154 640325 423196 640561
rect 422876 633561 423196 640325
rect 422876 633325 422918 633561
rect 423154 633325 423196 633561
rect 422876 626561 423196 633325
rect 422876 626325 422918 626561
rect 423154 626325 423196 626561
rect 422876 619561 423196 626325
rect 422876 619325 422918 619561
rect 423154 619325 423196 619561
rect 422876 612561 423196 619325
rect 422876 612325 422918 612561
rect 423154 612325 423196 612561
rect 422876 605561 423196 612325
rect 422876 605325 422918 605561
rect 423154 605325 423196 605561
rect 422876 598561 423196 605325
rect 422876 598325 422918 598561
rect 423154 598325 423196 598561
rect 422876 591561 423196 598325
rect 422876 591325 422918 591561
rect 423154 591325 423196 591561
rect 422876 584561 423196 591325
rect 422876 584325 422918 584561
rect 423154 584325 423196 584561
rect 422876 577561 423196 584325
rect 422876 577325 422918 577561
rect 423154 577325 423196 577561
rect 422876 570561 423196 577325
rect 422876 570325 422918 570561
rect 423154 570325 423196 570561
rect 422876 563561 423196 570325
rect 422876 563325 422918 563561
rect 423154 563325 423196 563561
rect 422876 556561 423196 563325
rect 422876 556325 422918 556561
rect 423154 556325 423196 556561
rect 422876 549561 423196 556325
rect 422876 549325 422918 549561
rect 423154 549325 423196 549561
rect 422876 542561 423196 549325
rect 422876 542325 422918 542561
rect 423154 542325 423196 542561
rect 422876 535561 423196 542325
rect 422876 535325 422918 535561
rect 423154 535325 423196 535561
rect 422876 528561 423196 535325
rect 422876 528325 422918 528561
rect 423154 528325 423196 528561
rect 422876 521561 423196 528325
rect 422876 521325 422918 521561
rect 423154 521325 423196 521561
rect 422876 514561 423196 521325
rect 422876 514325 422918 514561
rect 423154 514325 423196 514561
rect 422876 507561 423196 514325
rect 422876 507325 422918 507561
rect 423154 507325 423196 507561
rect 422876 500561 423196 507325
rect 422876 500325 422918 500561
rect 423154 500325 423196 500561
rect 422876 493561 423196 500325
rect 422876 493325 422918 493561
rect 423154 493325 423196 493561
rect 422876 486561 423196 493325
rect 422876 486325 422918 486561
rect 423154 486325 423196 486561
rect 422876 479561 423196 486325
rect 422876 479325 422918 479561
rect 423154 479325 423196 479561
rect 422876 472561 423196 479325
rect 422876 472325 422918 472561
rect 423154 472325 423196 472561
rect 422876 465561 423196 472325
rect 422876 465325 422918 465561
rect 423154 465325 423196 465561
rect 422876 458561 423196 465325
rect 422876 458325 422918 458561
rect 423154 458325 423196 458561
rect 422876 451561 423196 458325
rect 422876 451325 422918 451561
rect 423154 451325 423196 451561
rect 422876 444561 423196 451325
rect 422876 444325 422918 444561
rect 423154 444325 423196 444561
rect 422876 437561 423196 444325
rect 422876 437325 422918 437561
rect 423154 437325 423196 437561
rect 422876 430561 423196 437325
rect 422876 430325 422918 430561
rect 423154 430325 423196 430561
rect 422876 423561 423196 430325
rect 422876 423325 422918 423561
rect 423154 423325 423196 423561
rect 422876 416561 423196 423325
rect 422876 416325 422918 416561
rect 423154 416325 423196 416561
rect 422876 409561 423196 416325
rect 422876 409325 422918 409561
rect 423154 409325 423196 409561
rect 422876 402561 423196 409325
rect 422876 402325 422918 402561
rect 423154 402325 423196 402561
rect 422876 395561 423196 402325
rect 422876 395325 422918 395561
rect 423154 395325 423196 395561
rect 422876 388561 423196 395325
rect 422876 388325 422918 388561
rect 423154 388325 423196 388561
rect 422876 381561 423196 388325
rect 422876 381325 422918 381561
rect 423154 381325 423196 381561
rect 422876 374561 423196 381325
rect 422876 374325 422918 374561
rect 423154 374325 423196 374561
rect 422876 367561 423196 374325
rect 422876 367325 422918 367561
rect 423154 367325 423196 367561
rect 422876 360561 423196 367325
rect 422876 360325 422918 360561
rect 423154 360325 423196 360561
rect 422876 353561 423196 360325
rect 422876 353325 422918 353561
rect 423154 353325 423196 353561
rect 422876 346561 423196 353325
rect 422876 346325 422918 346561
rect 423154 346325 423196 346561
rect 422876 339561 423196 346325
rect 422876 339325 422918 339561
rect 423154 339325 423196 339561
rect 422876 332561 423196 339325
rect 422876 332325 422918 332561
rect 423154 332325 423196 332561
rect 422876 325561 423196 332325
rect 422876 325325 422918 325561
rect 423154 325325 423196 325561
rect 422876 318561 423196 325325
rect 422876 318325 422918 318561
rect 423154 318325 423196 318561
rect 422876 311561 423196 318325
rect 422876 311325 422918 311561
rect 423154 311325 423196 311561
rect 422876 304561 423196 311325
rect 422876 304325 422918 304561
rect 423154 304325 423196 304561
rect 422876 297561 423196 304325
rect 422876 297325 422918 297561
rect 423154 297325 423196 297561
rect 422876 290561 423196 297325
rect 422876 290325 422918 290561
rect 423154 290325 423196 290561
rect 422876 283561 423196 290325
rect 422876 283325 422918 283561
rect 423154 283325 423196 283561
rect 422876 276561 423196 283325
rect 422876 276325 422918 276561
rect 423154 276325 423196 276561
rect 422876 269561 423196 276325
rect 422876 269325 422918 269561
rect 423154 269325 423196 269561
rect 422876 262561 423196 269325
rect 422876 262325 422918 262561
rect 423154 262325 423196 262561
rect 422876 255561 423196 262325
rect 422876 255325 422918 255561
rect 423154 255325 423196 255561
rect 422876 248561 423196 255325
rect 422876 248325 422918 248561
rect 423154 248325 423196 248561
rect 422876 241561 423196 248325
rect 422876 241325 422918 241561
rect 423154 241325 423196 241561
rect 422876 234561 423196 241325
rect 422876 234325 422918 234561
rect 423154 234325 423196 234561
rect 422876 227561 423196 234325
rect 422876 227325 422918 227561
rect 423154 227325 423196 227561
rect 422876 220561 423196 227325
rect 422876 220325 422918 220561
rect 423154 220325 423196 220561
rect 422876 213561 423196 220325
rect 422876 213325 422918 213561
rect 423154 213325 423196 213561
rect 422876 206561 423196 213325
rect 422876 206325 422918 206561
rect 423154 206325 423196 206561
rect 422876 199561 423196 206325
rect 422876 199325 422918 199561
rect 423154 199325 423196 199561
rect 422876 192561 423196 199325
rect 422876 192325 422918 192561
rect 423154 192325 423196 192561
rect 422876 185561 423196 192325
rect 422876 185325 422918 185561
rect 423154 185325 423196 185561
rect 422876 178561 423196 185325
rect 422876 178325 422918 178561
rect 423154 178325 423196 178561
rect 422876 171561 423196 178325
rect 422876 171325 422918 171561
rect 423154 171325 423196 171561
rect 422876 164561 423196 171325
rect 422876 164325 422918 164561
rect 423154 164325 423196 164561
rect 422876 157561 423196 164325
rect 422876 157325 422918 157561
rect 423154 157325 423196 157561
rect 422876 150561 423196 157325
rect 422876 150325 422918 150561
rect 423154 150325 423196 150561
rect 422876 143561 423196 150325
rect 422876 143325 422918 143561
rect 423154 143325 423196 143561
rect 422876 136561 423196 143325
rect 422876 136325 422918 136561
rect 423154 136325 423196 136561
rect 422876 129561 423196 136325
rect 422876 129325 422918 129561
rect 423154 129325 423196 129561
rect 422876 122561 423196 129325
rect 422876 122325 422918 122561
rect 423154 122325 423196 122561
rect 422876 115561 423196 122325
rect 422876 115325 422918 115561
rect 423154 115325 423196 115561
rect 422876 108561 423196 115325
rect 422876 108325 422918 108561
rect 423154 108325 423196 108561
rect 422876 101561 423196 108325
rect 422876 101325 422918 101561
rect 423154 101325 423196 101561
rect 422876 94561 423196 101325
rect 422876 94325 422918 94561
rect 423154 94325 423196 94561
rect 422876 87561 423196 94325
rect 422876 87325 422918 87561
rect 423154 87325 423196 87561
rect 422876 80561 423196 87325
rect 422876 80325 422918 80561
rect 423154 80325 423196 80561
rect 422876 73561 423196 80325
rect 422876 73325 422918 73561
rect 423154 73325 423196 73561
rect 422876 66561 423196 73325
rect 422876 66325 422918 66561
rect 423154 66325 423196 66561
rect 422876 59561 423196 66325
rect 422876 59325 422918 59561
rect 423154 59325 423196 59561
rect 422876 52561 423196 59325
rect 422876 52325 422918 52561
rect 423154 52325 423196 52561
rect 422876 45561 423196 52325
rect 422876 45325 422918 45561
rect 423154 45325 423196 45561
rect 422876 38561 423196 45325
rect 422876 38325 422918 38561
rect 423154 38325 423196 38561
rect 422876 31561 423196 38325
rect 422876 31325 422918 31561
rect 423154 31325 423196 31561
rect 422876 24561 423196 31325
rect 422876 24325 422918 24561
rect 423154 24325 423196 24561
rect 422876 17561 423196 24325
rect 422876 17325 422918 17561
rect 423154 17325 423196 17561
rect 422876 10561 423196 17325
rect 422876 10325 422918 10561
rect 423154 10325 423196 10561
rect 422876 3561 423196 10325
rect 422876 3325 422918 3561
rect 423154 3325 423196 3561
rect 422876 -1706 423196 3325
rect 422876 -1942 422918 -1706
rect 423154 -1942 423196 -1706
rect 422876 -2026 423196 -1942
rect 422876 -2262 422918 -2026
rect 423154 -2262 423196 -2026
rect 422876 -2294 423196 -2262
rect 428144 705238 428464 706230
rect 428144 705002 428186 705238
rect 428422 705002 428464 705238
rect 428144 704918 428464 705002
rect 428144 704682 428186 704918
rect 428422 704682 428464 704918
rect 428144 695494 428464 704682
rect 428144 695258 428186 695494
rect 428422 695258 428464 695494
rect 428144 688494 428464 695258
rect 428144 688258 428186 688494
rect 428422 688258 428464 688494
rect 428144 681494 428464 688258
rect 428144 681258 428186 681494
rect 428422 681258 428464 681494
rect 428144 674494 428464 681258
rect 428144 674258 428186 674494
rect 428422 674258 428464 674494
rect 428144 667494 428464 674258
rect 428144 667258 428186 667494
rect 428422 667258 428464 667494
rect 428144 660494 428464 667258
rect 428144 660258 428186 660494
rect 428422 660258 428464 660494
rect 428144 653494 428464 660258
rect 428144 653258 428186 653494
rect 428422 653258 428464 653494
rect 428144 646494 428464 653258
rect 428144 646258 428186 646494
rect 428422 646258 428464 646494
rect 428144 639494 428464 646258
rect 428144 639258 428186 639494
rect 428422 639258 428464 639494
rect 428144 632494 428464 639258
rect 428144 632258 428186 632494
rect 428422 632258 428464 632494
rect 428144 625494 428464 632258
rect 428144 625258 428186 625494
rect 428422 625258 428464 625494
rect 428144 618494 428464 625258
rect 428144 618258 428186 618494
rect 428422 618258 428464 618494
rect 428144 611494 428464 618258
rect 428144 611258 428186 611494
rect 428422 611258 428464 611494
rect 428144 604494 428464 611258
rect 428144 604258 428186 604494
rect 428422 604258 428464 604494
rect 428144 597494 428464 604258
rect 428144 597258 428186 597494
rect 428422 597258 428464 597494
rect 428144 590494 428464 597258
rect 428144 590258 428186 590494
rect 428422 590258 428464 590494
rect 428144 583494 428464 590258
rect 428144 583258 428186 583494
rect 428422 583258 428464 583494
rect 428144 576494 428464 583258
rect 428144 576258 428186 576494
rect 428422 576258 428464 576494
rect 428144 569494 428464 576258
rect 428144 569258 428186 569494
rect 428422 569258 428464 569494
rect 428144 562494 428464 569258
rect 428144 562258 428186 562494
rect 428422 562258 428464 562494
rect 428144 555494 428464 562258
rect 428144 555258 428186 555494
rect 428422 555258 428464 555494
rect 428144 548494 428464 555258
rect 428144 548258 428186 548494
rect 428422 548258 428464 548494
rect 428144 541494 428464 548258
rect 428144 541258 428186 541494
rect 428422 541258 428464 541494
rect 428144 534494 428464 541258
rect 428144 534258 428186 534494
rect 428422 534258 428464 534494
rect 428144 527494 428464 534258
rect 428144 527258 428186 527494
rect 428422 527258 428464 527494
rect 428144 520494 428464 527258
rect 428144 520258 428186 520494
rect 428422 520258 428464 520494
rect 428144 513494 428464 520258
rect 428144 513258 428186 513494
rect 428422 513258 428464 513494
rect 428144 506494 428464 513258
rect 428144 506258 428186 506494
rect 428422 506258 428464 506494
rect 428144 499494 428464 506258
rect 428144 499258 428186 499494
rect 428422 499258 428464 499494
rect 428144 492494 428464 499258
rect 428144 492258 428186 492494
rect 428422 492258 428464 492494
rect 428144 485494 428464 492258
rect 428144 485258 428186 485494
rect 428422 485258 428464 485494
rect 428144 478494 428464 485258
rect 428144 478258 428186 478494
rect 428422 478258 428464 478494
rect 428144 471494 428464 478258
rect 428144 471258 428186 471494
rect 428422 471258 428464 471494
rect 428144 464494 428464 471258
rect 428144 464258 428186 464494
rect 428422 464258 428464 464494
rect 428144 457494 428464 464258
rect 428144 457258 428186 457494
rect 428422 457258 428464 457494
rect 428144 450494 428464 457258
rect 428144 450258 428186 450494
rect 428422 450258 428464 450494
rect 428144 443494 428464 450258
rect 428144 443258 428186 443494
rect 428422 443258 428464 443494
rect 428144 436494 428464 443258
rect 428144 436258 428186 436494
rect 428422 436258 428464 436494
rect 428144 429494 428464 436258
rect 428144 429258 428186 429494
rect 428422 429258 428464 429494
rect 428144 422494 428464 429258
rect 428144 422258 428186 422494
rect 428422 422258 428464 422494
rect 428144 415494 428464 422258
rect 428144 415258 428186 415494
rect 428422 415258 428464 415494
rect 428144 408494 428464 415258
rect 428144 408258 428186 408494
rect 428422 408258 428464 408494
rect 428144 401494 428464 408258
rect 428144 401258 428186 401494
rect 428422 401258 428464 401494
rect 428144 394494 428464 401258
rect 428144 394258 428186 394494
rect 428422 394258 428464 394494
rect 428144 387494 428464 394258
rect 428144 387258 428186 387494
rect 428422 387258 428464 387494
rect 428144 380494 428464 387258
rect 428144 380258 428186 380494
rect 428422 380258 428464 380494
rect 428144 373494 428464 380258
rect 428144 373258 428186 373494
rect 428422 373258 428464 373494
rect 428144 366494 428464 373258
rect 428144 366258 428186 366494
rect 428422 366258 428464 366494
rect 428144 359494 428464 366258
rect 428144 359258 428186 359494
rect 428422 359258 428464 359494
rect 428144 352494 428464 359258
rect 428144 352258 428186 352494
rect 428422 352258 428464 352494
rect 428144 345494 428464 352258
rect 428144 345258 428186 345494
rect 428422 345258 428464 345494
rect 428144 338494 428464 345258
rect 428144 338258 428186 338494
rect 428422 338258 428464 338494
rect 428144 331494 428464 338258
rect 428144 331258 428186 331494
rect 428422 331258 428464 331494
rect 428144 324494 428464 331258
rect 428144 324258 428186 324494
rect 428422 324258 428464 324494
rect 428144 317494 428464 324258
rect 428144 317258 428186 317494
rect 428422 317258 428464 317494
rect 428144 310494 428464 317258
rect 428144 310258 428186 310494
rect 428422 310258 428464 310494
rect 428144 303494 428464 310258
rect 428144 303258 428186 303494
rect 428422 303258 428464 303494
rect 428144 296494 428464 303258
rect 428144 296258 428186 296494
rect 428422 296258 428464 296494
rect 428144 289494 428464 296258
rect 428144 289258 428186 289494
rect 428422 289258 428464 289494
rect 428144 282494 428464 289258
rect 428144 282258 428186 282494
rect 428422 282258 428464 282494
rect 428144 275494 428464 282258
rect 428144 275258 428186 275494
rect 428422 275258 428464 275494
rect 428144 268494 428464 275258
rect 428144 268258 428186 268494
rect 428422 268258 428464 268494
rect 428144 261494 428464 268258
rect 428144 261258 428186 261494
rect 428422 261258 428464 261494
rect 428144 254494 428464 261258
rect 428144 254258 428186 254494
rect 428422 254258 428464 254494
rect 428144 247494 428464 254258
rect 428144 247258 428186 247494
rect 428422 247258 428464 247494
rect 428144 240494 428464 247258
rect 428144 240258 428186 240494
rect 428422 240258 428464 240494
rect 428144 233494 428464 240258
rect 428144 233258 428186 233494
rect 428422 233258 428464 233494
rect 428144 226494 428464 233258
rect 428144 226258 428186 226494
rect 428422 226258 428464 226494
rect 428144 219494 428464 226258
rect 428144 219258 428186 219494
rect 428422 219258 428464 219494
rect 428144 212494 428464 219258
rect 428144 212258 428186 212494
rect 428422 212258 428464 212494
rect 428144 205494 428464 212258
rect 428144 205258 428186 205494
rect 428422 205258 428464 205494
rect 428144 198494 428464 205258
rect 428144 198258 428186 198494
rect 428422 198258 428464 198494
rect 428144 191494 428464 198258
rect 428144 191258 428186 191494
rect 428422 191258 428464 191494
rect 428144 184494 428464 191258
rect 428144 184258 428186 184494
rect 428422 184258 428464 184494
rect 428144 177494 428464 184258
rect 428144 177258 428186 177494
rect 428422 177258 428464 177494
rect 428144 170494 428464 177258
rect 428144 170258 428186 170494
rect 428422 170258 428464 170494
rect 428144 163494 428464 170258
rect 428144 163258 428186 163494
rect 428422 163258 428464 163494
rect 428144 156494 428464 163258
rect 428144 156258 428186 156494
rect 428422 156258 428464 156494
rect 428144 149494 428464 156258
rect 428144 149258 428186 149494
rect 428422 149258 428464 149494
rect 428144 142494 428464 149258
rect 428144 142258 428186 142494
rect 428422 142258 428464 142494
rect 428144 135494 428464 142258
rect 428144 135258 428186 135494
rect 428422 135258 428464 135494
rect 428144 128494 428464 135258
rect 428144 128258 428186 128494
rect 428422 128258 428464 128494
rect 428144 121494 428464 128258
rect 428144 121258 428186 121494
rect 428422 121258 428464 121494
rect 428144 114494 428464 121258
rect 428144 114258 428186 114494
rect 428422 114258 428464 114494
rect 428144 107494 428464 114258
rect 428144 107258 428186 107494
rect 428422 107258 428464 107494
rect 428144 100494 428464 107258
rect 428144 100258 428186 100494
rect 428422 100258 428464 100494
rect 428144 93494 428464 100258
rect 428144 93258 428186 93494
rect 428422 93258 428464 93494
rect 428144 86494 428464 93258
rect 428144 86258 428186 86494
rect 428422 86258 428464 86494
rect 428144 79494 428464 86258
rect 428144 79258 428186 79494
rect 428422 79258 428464 79494
rect 428144 72494 428464 79258
rect 428144 72258 428186 72494
rect 428422 72258 428464 72494
rect 428144 65494 428464 72258
rect 428144 65258 428186 65494
rect 428422 65258 428464 65494
rect 428144 58494 428464 65258
rect 428144 58258 428186 58494
rect 428422 58258 428464 58494
rect 428144 51494 428464 58258
rect 428144 51258 428186 51494
rect 428422 51258 428464 51494
rect 428144 44494 428464 51258
rect 428144 44258 428186 44494
rect 428422 44258 428464 44494
rect 428144 37494 428464 44258
rect 428144 37258 428186 37494
rect 428422 37258 428464 37494
rect 428144 30494 428464 37258
rect 428144 30258 428186 30494
rect 428422 30258 428464 30494
rect 428144 23494 428464 30258
rect 428144 23258 428186 23494
rect 428422 23258 428464 23494
rect 428144 16494 428464 23258
rect 428144 16258 428186 16494
rect 428422 16258 428464 16494
rect 428144 9494 428464 16258
rect 428144 9258 428186 9494
rect 428422 9258 428464 9494
rect 428144 2494 428464 9258
rect 428144 2258 428186 2494
rect 428422 2258 428464 2494
rect 428144 -746 428464 2258
rect 428144 -982 428186 -746
rect 428422 -982 428464 -746
rect 428144 -1066 428464 -982
rect 428144 -1302 428186 -1066
rect 428422 -1302 428464 -1066
rect 428144 -2294 428464 -1302
rect 429876 706198 430196 706230
rect 429876 705962 429918 706198
rect 430154 705962 430196 706198
rect 429876 705878 430196 705962
rect 429876 705642 429918 705878
rect 430154 705642 430196 705878
rect 429876 696561 430196 705642
rect 429876 696325 429918 696561
rect 430154 696325 430196 696561
rect 429876 689561 430196 696325
rect 429876 689325 429918 689561
rect 430154 689325 430196 689561
rect 429876 682561 430196 689325
rect 429876 682325 429918 682561
rect 430154 682325 430196 682561
rect 429876 675561 430196 682325
rect 429876 675325 429918 675561
rect 430154 675325 430196 675561
rect 429876 668561 430196 675325
rect 429876 668325 429918 668561
rect 430154 668325 430196 668561
rect 429876 661561 430196 668325
rect 429876 661325 429918 661561
rect 430154 661325 430196 661561
rect 429876 654561 430196 661325
rect 429876 654325 429918 654561
rect 430154 654325 430196 654561
rect 429876 647561 430196 654325
rect 429876 647325 429918 647561
rect 430154 647325 430196 647561
rect 429876 640561 430196 647325
rect 429876 640325 429918 640561
rect 430154 640325 430196 640561
rect 429876 633561 430196 640325
rect 429876 633325 429918 633561
rect 430154 633325 430196 633561
rect 429876 626561 430196 633325
rect 429876 626325 429918 626561
rect 430154 626325 430196 626561
rect 429876 619561 430196 626325
rect 429876 619325 429918 619561
rect 430154 619325 430196 619561
rect 429876 612561 430196 619325
rect 429876 612325 429918 612561
rect 430154 612325 430196 612561
rect 429876 605561 430196 612325
rect 429876 605325 429918 605561
rect 430154 605325 430196 605561
rect 429876 598561 430196 605325
rect 429876 598325 429918 598561
rect 430154 598325 430196 598561
rect 429876 591561 430196 598325
rect 429876 591325 429918 591561
rect 430154 591325 430196 591561
rect 429876 584561 430196 591325
rect 429876 584325 429918 584561
rect 430154 584325 430196 584561
rect 429876 577561 430196 584325
rect 429876 577325 429918 577561
rect 430154 577325 430196 577561
rect 429876 570561 430196 577325
rect 429876 570325 429918 570561
rect 430154 570325 430196 570561
rect 429876 563561 430196 570325
rect 429876 563325 429918 563561
rect 430154 563325 430196 563561
rect 429876 556561 430196 563325
rect 429876 556325 429918 556561
rect 430154 556325 430196 556561
rect 429876 549561 430196 556325
rect 429876 549325 429918 549561
rect 430154 549325 430196 549561
rect 429876 542561 430196 549325
rect 429876 542325 429918 542561
rect 430154 542325 430196 542561
rect 429876 535561 430196 542325
rect 429876 535325 429918 535561
rect 430154 535325 430196 535561
rect 429876 528561 430196 535325
rect 429876 528325 429918 528561
rect 430154 528325 430196 528561
rect 429876 521561 430196 528325
rect 429876 521325 429918 521561
rect 430154 521325 430196 521561
rect 429876 514561 430196 521325
rect 429876 514325 429918 514561
rect 430154 514325 430196 514561
rect 429876 507561 430196 514325
rect 429876 507325 429918 507561
rect 430154 507325 430196 507561
rect 429876 500561 430196 507325
rect 429876 500325 429918 500561
rect 430154 500325 430196 500561
rect 429876 493561 430196 500325
rect 429876 493325 429918 493561
rect 430154 493325 430196 493561
rect 429876 486561 430196 493325
rect 429876 486325 429918 486561
rect 430154 486325 430196 486561
rect 429876 479561 430196 486325
rect 429876 479325 429918 479561
rect 430154 479325 430196 479561
rect 429876 472561 430196 479325
rect 429876 472325 429918 472561
rect 430154 472325 430196 472561
rect 429876 465561 430196 472325
rect 429876 465325 429918 465561
rect 430154 465325 430196 465561
rect 429876 458561 430196 465325
rect 429876 458325 429918 458561
rect 430154 458325 430196 458561
rect 429876 451561 430196 458325
rect 429876 451325 429918 451561
rect 430154 451325 430196 451561
rect 429876 444561 430196 451325
rect 429876 444325 429918 444561
rect 430154 444325 430196 444561
rect 429876 437561 430196 444325
rect 429876 437325 429918 437561
rect 430154 437325 430196 437561
rect 429876 430561 430196 437325
rect 429876 430325 429918 430561
rect 430154 430325 430196 430561
rect 429876 423561 430196 430325
rect 429876 423325 429918 423561
rect 430154 423325 430196 423561
rect 429876 416561 430196 423325
rect 429876 416325 429918 416561
rect 430154 416325 430196 416561
rect 429876 409561 430196 416325
rect 429876 409325 429918 409561
rect 430154 409325 430196 409561
rect 429876 402561 430196 409325
rect 429876 402325 429918 402561
rect 430154 402325 430196 402561
rect 429876 395561 430196 402325
rect 429876 395325 429918 395561
rect 430154 395325 430196 395561
rect 429876 388561 430196 395325
rect 429876 388325 429918 388561
rect 430154 388325 430196 388561
rect 429876 381561 430196 388325
rect 429876 381325 429918 381561
rect 430154 381325 430196 381561
rect 429876 374561 430196 381325
rect 429876 374325 429918 374561
rect 430154 374325 430196 374561
rect 429876 367561 430196 374325
rect 429876 367325 429918 367561
rect 430154 367325 430196 367561
rect 429876 360561 430196 367325
rect 429876 360325 429918 360561
rect 430154 360325 430196 360561
rect 429876 353561 430196 360325
rect 429876 353325 429918 353561
rect 430154 353325 430196 353561
rect 429876 346561 430196 353325
rect 429876 346325 429918 346561
rect 430154 346325 430196 346561
rect 429876 339561 430196 346325
rect 429876 339325 429918 339561
rect 430154 339325 430196 339561
rect 429876 332561 430196 339325
rect 429876 332325 429918 332561
rect 430154 332325 430196 332561
rect 429876 325561 430196 332325
rect 429876 325325 429918 325561
rect 430154 325325 430196 325561
rect 429876 318561 430196 325325
rect 429876 318325 429918 318561
rect 430154 318325 430196 318561
rect 429876 311561 430196 318325
rect 429876 311325 429918 311561
rect 430154 311325 430196 311561
rect 429876 304561 430196 311325
rect 429876 304325 429918 304561
rect 430154 304325 430196 304561
rect 429876 297561 430196 304325
rect 429876 297325 429918 297561
rect 430154 297325 430196 297561
rect 429876 290561 430196 297325
rect 429876 290325 429918 290561
rect 430154 290325 430196 290561
rect 429876 283561 430196 290325
rect 429876 283325 429918 283561
rect 430154 283325 430196 283561
rect 429876 276561 430196 283325
rect 429876 276325 429918 276561
rect 430154 276325 430196 276561
rect 429876 269561 430196 276325
rect 429876 269325 429918 269561
rect 430154 269325 430196 269561
rect 429876 262561 430196 269325
rect 429876 262325 429918 262561
rect 430154 262325 430196 262561
rect 429876 255561 430196 262325
rect 429876 255325 429918 255561
rect 430154 255325 430196 255561
rect 429876 248561 430196 255325
rect 429876 248325 429918 248561
rect 430154 248325 430196 248561
rect 429876 241561 430196 248325
rect 429876 241325 429918 241561
rect 430154 241325 430196 241561
rect 429876 234561 430196 241325
rect 429876 234325 429918 234561
rect 430154 234325 430196 234561
rect 429876 227561 430196 234325
rect 429876 227325 429918 227561
rect 430154 227325 430196 227561
rect 429876 220561 430196 227325
rect 429876 220325 429918 220561
rect 430154 220325 430196 220561
rect 429876 213561 430196 220325
rect 429876 213325 429918 213561
rect 430154 213325 430196 213561
rect 429876 206561 430196 213325
rect 429876 206325 429918 206561
rect 430154 206325 430196 206561
rect 429876 199561 430196 206325
rect 429876 199325 429918 199561
rect 430154 199325 430196 199561
rect 429876 192561 430196 199325
rect 429876 192325 429918 192561
rect 430154 192325 430196 192561
rect 429876 185561 430196 192325
rect 429876 185325 429918 185561
rect 430154 185325 430196 185561
rect 429876 178561 430196 185325
rect 429876 178325 429918 178561
rect 430154 178325 430196 178561
rect 429876 171561 430196 178325
rect 429876 171325 429918 171561
rect 430154 171325 430196 171561
rect 429876 164561 430196 171325
rect 429876 164325 429918 164561
rect 430154 164325 430196 164561
rect 429876 157561 430196 164325
rect 429876 157325 429918 157561
rect 430154 157325 430196 157561
rect 429876 150561 430196 157325
rect 429876 150325 429918 150561
rect 430154 150325 430196 150561
rect 429876 143561 430196 150325
rect 429876 143325 429918 143561
rect 430154 143325 430196 143561
rect 429876 136561 430196 143325
rect 429876 136325 429918 136561
rect 430154 136325 430196 136561
rect 429876 129561 430196 136325
rect 429876 129325 429918 129561
rect 430154 129325 430196 129561
rect 429876 122561 430196 129325
rect 429876 122325 429918 122561
rect 430154 122325 430196 122561
rect 429876 115561 430196 122325
rect 429876 115325 429918 115561
rect 430154 115325 430196 115561
rect 429876 108561 430196 115325
rect 429876 108325 429918 108561
rect 430154 108325 430196 108561
rect 429876 101561 430196 108325
rect 429876 101325 429918 101561
rect 430154 101325 430196 101561
rect 429876 94561 430196 101325
rect 429876 94325 429918 94561
rect 430154 94325 430196 94561
rect 429876 87561 430196 94325
rect 429876 87325 429918 87561
rect 430154 87325 430196 87561
rect 429876 80561 430196 87325
rect 429876 80325 429918 80561
rect 430154 80325 430196 80561
rect 429876 73561 430196 80325
rect 429876 73325 429918 73561
rect 430154 73325 430196 73561
rect 429876 66561 430196 73325
rect 429876 66325 429918 66561
rect 430154 66325 430196 66561
rect 429876 59561 430196 66325
rect 429876 59325 429918 59561
rect 430154 59325 430196 59561
rect 429876 52561 430196 59325
rect 429876 52325 429918 52561
rect 430154 52325 430196 52561
rect 429876 45561 430196 52325
rect 429876 45325 429918 45561
rect 430154 45325 430196 45561
rect 429876 38561 430196 45325
rect 429876 38325 429918 38561
rect 430154 38325 430196 38561
rect 429876 31561 430196 38325
rect 429876 31325 429918 31561
rect 430154 31325 430196 31561
rect 429876 24561 430196 31325
rect 429876 24325 429918 24561
rect 430154 24325 430196 24561
rect 429876 17561 430196 24325
rect 429876 17325 429918 17561
rect 430154 17325 430196 17561
rect 429876 10561 430196 17325
rect 429876 10325 429918 10561
rect 430154 10325 430196 10561
rect 429876 3561 430196 10325
rect 429876 3325 429918 3561
rect 430154 3325 430196 3561
rect 429876 -1706 430196 3325
rect 429876 -1942 429918 -1706
rect 430154 -1942 430196 -1706
rect 429876 -2026 430196 -1942
rect 429876 -2262 429918 -2026
rect 430154 -2262 430196 -2026
rect 429876 -2294 430196 -2262
rect 435144 705238 435464 706230
rect 435144 705002 435186 705238
rect 435422 705002 435464 705238
rect 435144 704918 435464 705002
rect 435144 704682 435186 704918
rect 435422 704682 435464 704918
rect 435144 695494 435464 704682
rect 435144 695258 435186 695494
rect 435422 695258 435464 695494
rect 435144 688494 435464 695258
rect 435144 688258 435186 688494
rect 435422 688258 435464 688494
rect 435144 681494 435464 688258
rect 435144 681258 435186 681494
rect 435422 681258 435464 681494
rect 435144 674494 435464 681258
rect 435144 674258 435186 674494
rect 435422 674258 435464 674494
rect 435144 667494 435464 674258
rect 435144 667258 435186 667494
rect 435422 667258 435464 667494
rect 435144 660494 435464 667258
rect 435144 660258 435186 660494
rect 435422 660258 435464 660494
rect 435144 653494 435464 660258
rect 435144 653258 435186 653494
rect 435422 653258 435464 653494
rect 435144 646494 435464 653258
rect 435144 646258 435186 646494
rect 435422 646258 435464 646494
rect 435144 639494 435464 646258
rect 435144 639258 435186 639494
rect 435422 639258 435464 639494
rect 435144 632494 435464 639258
rect 435144 632258 435186 632494
rect 435422 632258 435464 632494
rect 435144 625494 435464 632258
rect 435144 625258 435186 625494
rect 435422 625258 435464 625494
rect 435144 618494 435464 625258
rect 435144 618258 435186 618494
rect 435422 618258 435464 618494
rect 435144 611494 435464 618258
rect 435144 611258 435186 611494
rect 435422 611258 435464 611494
rect 435144 604494 435464 611258
rect 435144 604258 435186 604494
rect 435422 604258 435464 604494
rect 435144 597494 435464 604258
rect 435144 597258 435186 597494
rect 435422 597258 435464 597494
rect 435144 590494 435464 597258
rect 435144 590258 435186 590494
rect 435422 590258 435464 590494
rect 435144 583494 435464 590258
rect 435144 583258 435186 583494
rect 435422 583258 435464 583494
rect 435144 576494 435464 583258
rect 435144 576258 435186 576494
rect 435422 576258 435464 576494
rect 435144 569494 435464 576258
rect 435144 569258 435186 569494
rect 435422 569258 435464 569494
rect 435144 562494 435464 569258
rect 435144 562258 435186 562494
rect 435422 562258 435464 562494
rect 435144 555494 435464 562258
rect 435144 555258 435186 555494
rect 435422 555258 435464 555494
rect 435144 548494 435464 555258
rect 435144 548258 435186 548494
rect 435422 548258 435464 548494
rect 435144 541494 435464 548258
rect 435144 541258 435186 541494
rect 435422 541258 435464 541494
rect 435144 534494 435464 541258
rect 435144 534258 435186 534494
rect 435422 534258 435464 534494
rect 435144 527494 435464 534258
rect 435144 527258 435186 527494
rect 435422 527258 435464 527494
rect 435144 520494 435464 527258
rect 435144 520258 435186 520494
rect 435422 520258 435464 520494
rect 435144 513494 435464 520258
rect 435144 513258 435186 513494
rect 435422 513258 435464 513494
rect 435144 506494 435464 513258
rect 435144 506258 435186 506494
rect 435422 506258 435464 506494
rect 435144 499494 435464 506258
rect 435144 499258 435186 499494
rect 435422 499258 435464 499494
rect 435144 492494 435464 499258
rect 435144 492258 435186 492494
rect 435422 492258 435464 492494
rect 435144 485494 435464 492258
rect 435144 485258 435186 485494
rect 435422 485258 435464 485494
rect 435144 478494 435464 485258
rect 435144 478258 435186 478494
rect 435422 478258 435464 478494
rect 435144 471494 435464 478258
rect 435144 471258 435186 471494
rect 435422 471258 435464 471494
rect 435144 464494 435464 471258
rect 435144 464258 435186 464494
rect 435422 464258 435464 464494
rect 435144 457494 435464 464258
rect 435144 457258 435186 457494
rect 435422 457258 435464 457494
rect 435144 450494 435464 457258
rect 435144 450258 435186 450494
rect 435422 450258 435464 450494
rect 435144 443494 435464 450258
rect 435144 443258 435186 443494
rect 435422 443258 435464 443494
rect 435144 436494 435464 443258
rect 435144 436258 435186 436494
rect 435422 436258 435464 436494
rect 435144 429494 435464 436258
rect 435144 429258 435186 429494
rect 435422 429258 435464 429494
rect 435144 422494 435464 429258
rect 435144 422258 435186 422494
rect 435422 422258 435464 422494
rect 435144 415494 435464 422258
rect 435144 415258 435186 415494
rect 435422 415258 435464 415494
rect 435144 408494 435464 415258
rect 435144 408258 435186 408494
rect 435422 408258 435464 408494
rect 435144 401494 435464 408258
rect 435144 401258 435186 401494
rect 435422 401258 435464 401494
rect 435144 394494 435464 401258
rect 435144 394258 435186 394494
rect 435422 394258 435464 394494
rect 435144 387494 435464 394258
rect 435144 387258 435186 387494
rect 435422 387258 435464 387494
rect 435144 380494 435464 387258
rect 435144 380258 435186 380494
rect 435422 380258 435464 380494
rect 435144 373494 435464 380258
rect 435144 373258 435186 373494
rect 435422 373258 435464 373494
rect 435144 366494 435464 373258
rect 435144 366258 435186 366494
rect 435422 366258 435464 366494
rect 435144 359494 435464 366258
rect 435144 359258 435186 359494
rect 435422 359258 435464 359494
rect 435144 352494 435464 359258
rect 435144 352258 435186 352494
rect 435422 352258 435464 352494
rect 435144 345494 435464 352258
rect 435144 345258 435186 345494
rect 435422 345258 435464 345494
rect 435144 338494 435464 345258
rect 435144 338258 435186 338494
rect 435422 338258 435464 338494
rect 435144 331494 435464 338258
rect 435144 331258 435186 331494
rect 435422 331258 435464 331494
rect 435144 324494 435464 331258
rect 435144 324258 435186 324494
rect 435422 324258 435464 324494
rect 435144 317494 435464 324258
rect 435144 317258 435186 317494
rect 435422 317258 435464 317494
rect 435144 310494 435464 317258
rect 435144 310258 435186 310494
rect 435422 310258 435464 310494
rect 435144 303494 435464 310258
rect 435144 303258 435186 303494
rect 435422 303258 435464 303494
rect 435144 296494 435464 303258
rect 435144 296258 435186 296494
rect 435422 296258 435464 296494
rect 435144 289494 435464 296258
rect 435144 289258 435186 289494
rect 435422 289258 435464 289494
rect 435144 282494 435464 289258
rect 435144 282258 435186 282494
rect 435422 282258 435464 282494
rect 435144 275494 435464 282258
rect 435144 275258 435186 275494
rect 435422 275258 435464 275494
rect 435144 268494 435464 275258
rect 435144 268258 435186 268494
rect 435422 268258 435464 268494
rect 435144 261494 435464 268258
rect 435144 261258 435186 261494
rect 435422 261258 435464 261494
rect 435144 254494 435464 261258
rect 435144 254258 435186 254494
rect 435422 254258 435464 254494
rect 435144 247494 435464 254258
rect 435144 247258 435186 247494
rect 435422 247258 435464 247494
rect 435144 240494 435464 247258
rect 435144 240258 435186 240494
rect 435422 240258 435464 240494
rect 435144 233494 435464 240258
rect 435144 233258 435186 233494
rect 435422 233258 435464 233494
rect 435144 226494 435464 233258
rect 435144 226258 435186 226494
rect 435422 226258 435464 226494
rect 435144 219494 435464 226258
rect 435144 219258 435186 219494
rect 435422 219258 435464 219494
rect 435144 212494 435464 219258
rect 435144 212258 435186 212494
rect 435422 212258 435464 212494
rect 435144 205494 435464 212258
rect 435144 205258 435186 205494
rect 435422 205258 435464 205494
rect 435144 198494 435464 205258
rect 435144 198258 435186 198494
rect 435422 198258 435464 198494
rect 435144 191494 435464 198258
rect 435144 191258 435186 191494
rect 435422 191258 435464 191494
rect 435144 184494 435464 191258
rect 435144 184258 435186 184494
rect 435422 184258 435464 184494
rect 435144 177494 435464 184258
rect 435144 177258 435186 177494
rect 435422 177258 435464 177494
rect 435144 170494 435464 177258
rect 435144 170258 435186 170494
rect 435422 170258 435464 170494
rect 435144 163494 435464 170258
rect 435144 163258 435186 163494
rect 435422 163258 435464 163494
rect 435144 156494 435464 163258
rect 435144 156258 435186 156494
rect 435422 156258 435464 156494
rect 435144 149494 435464 156258
rect 435144 149258 435186 149494
rect 435422 149258 435464 149494
rect 435144 142494 435464 149258
rect 435144 142258 435186 142494
rect 435422 142258 435464 142494
rect 435144 135494 435464 142258
rect 435144 135258 435186 135494
rect 435422 135258 435464 135494
rect 435144 128494 435464 135258
rect 435144 128258 435186 128494
rect 435422 128258 435464 128494
rect 435144 121494 435464 128258
rect 435144 121258 435186 121494
rect 435422 121258 435464 121494
rect 435144 114494 435464 121258
rect 435144 114258 435186 114494
rect 435422 114258 435464 114494
rect 435144 107494 435464 114258
rect 435144 107258 435186 107494
rect 435422 107258 435464 107494
rect 435144 100494 435464 107258
rect 435144 100258 435186 100494
rect 435422 100258 435464 100494
rect 435144 93494 435464 100258
rect 435144 93258 435186 93494
rect 435422 93258 435464 93494
rect 435144 86494 435464 93258
rect 435144 86258 435186 86494
rect 435422 86258 435464 86494
rect 435144 79494 435464 86258
rect 435144 79258 435186 79494
rect 435422 79258 435464 79494
rect 435144 72494 435464 79258
rect 435144 72258 435186 72494
rect 435422 72258 435464 72494
rect 435144 65494 435464 72258
rect 435144 65258 435186 65494
rect 435422 65258 435464 65494
rect 435144 58494 435464 65258
rect 435144 58258 435186 58494
rect 435422 58258 435464 58494
rect 435144 51494 435464 58258
rect 435144 51258 435186 51494
rect 435422 51258 435464 51494
rect 435144 44494 435464 51258
rect 435144 44258 435186 44494
rect 435422 44258 435464 44494
rect 435144 37494 435464 44258
rect 435144 37258 435186 37494
rect 435422 37258 435464 37494
rect 435144 30494 435464 37258
rect 435144 30258 435186 30494
rect 435422 30258 435464 30494
rect 435144 23494 435464 30258
rect 435144 23258 435186 23494
rect 435422 23258 435464 23494
rect 435144 16494 435464 23258
rect 435144 16258 435186 16494
rect 435422 16258 435464 16494
rect 435144 9494 435464 16258
rect 435144 9258 435186 9494
rect 435422 9258 435464 9494
rect 435144 2494 435464 9258
rect 435144 2258 435186 2494
rect 435422 2258 435464 2494
rect 435144 -746 435464 2258
rect 435144 -982 435186 -746
rect 435422 -982 435464 -746
rect 435144 -1066 435464 -982
rect 435144 -1302 435186 -1066
rect 435422 -1302 435464 -1066
rect 435144 -2294 435464 -1302
rect 436876 706198 437196 706230
rect 436876 705962 436918 706198
rect 437154 705962 437196 706198
rect 436876 705878 437196 705962
rect 436876 705642 436918 705878
rect 437154 705642 437196 705878
rect 436876 696561 437196 705642
rect 436876 696325 436918 696561
rect 437154 696325 437196 696561
rect 436876 689561 437196 696325
rect 436876 689325 436918 689561
rect 437154 689325 437196 689561
rect 436876 682561 437196 689325
rect 436876 682325 436918 682561
rect 437154 682325 437196 682561
rect 436876 675561 437196 682325
rect 436876 675325 436918 675561
rect 437154 675325 437196 675561
rect 436876 668561 437196 675325
rect 436876 668325 436918 668561
rect 437154 668325 437196 668561
rect 436876 661561 437196 668325
rect 436876 661325 436918 661561
rect 437154 661325 437196 661561
rect 436876 654561 437196 661325
rect 436876 654325 436918 654561
rect 437154 654325 437196 654561
rect 436876 647561 437196 654325
rect 436876 647325 436918 647561
rect 437154 647325 437196 647561
rect 436876 640561 437196 647325
rect 436876 640325 436918 640561
rect 437154 640325 437196 640561
rect 436876 633561 437196 640325
rect 436876 633325 436918 633561
rect 437154 633325 437196 633561
rect 436876 626561 437196 633325
rect 436876 626325 436918 626561
rect 437154 626325 437196 626561
rect 436876 619561 437196 626325
rect 436876 619325 436918 619561
rect 437154 619325 437196 619561
rect 436876 612561 437196 619325
rect 436876 612325 436918 612561
rect 437154 612325 437196 612561
rect 436876 605561 437196 612325
rect 436876 605325 436918 605561
rect 437154 605325 437196 605561
rect 436876 598561 437196 605325
rect 436876 598325 436918 598561
rect 437154 598325 437196 598561
rect 436876 591561 437196 598325
rect 436876 591325 436918 591561
rect 437154 591325 437196 591561
rect 436876 584561 437196 591325
rect 436876 584325 436918 584561
rect 437154 584325 437196 584561
rect 436876 577561 437196 584325
rect 436876 577325 436918 577561
rect 437154 577325 437196 577561
rect 436876 570561 437196 577325
rect 436876 570325 436918 570561
rect 437154 570325 437196 570561
rect 436876 563561 437196 570325
rect 436876 563325 436918 563561
rect 437154 563325 437196 563561
rect 436876 556561 437196 563325
rect 436876 556325 436918 556561
rect 437154 556325 437196 556561
rect 436876 549561 437196 556325
rect 436876 549325 436918 549561
rect 437154 549325 437196 549561
rect 436876 542561 437196 549325
rect 436876 542325 436918 542561
rect 437154 542325 437196 542561
rect 436876 535561 437196 542325
rect 436876 535325 436918 535561
rect 437154 535325 437196 535561
rect 436876 528561 437196 535325
rect 436876 528325 436918 528561
rect 437154 528325 437196 528561
rect 436876 521561 437196 528325
rect 436876 521325 436918 521561
rect 437154 521325 437196 521561
rect 436876 514561 437196 521325
rect 436876 514325 436918 514561
rect 437154 514325 437196 514561
rect 436876 507561 437196 514325
rect 436876 507325 436918 507561
rect 437154 507325 437196 507561
rect 436876 500561 437196 507325
rect 436876 500325 436918 500561
rect 437154 500325 437196 500561
rect 436876 493561 437196 500325
rect 436876 493325 436918 493561
rect 437154 493325 437196 493561
rect 436876 486561 437196 493325
rect 436876 486325 436918 486561
rect 437154 486325 437196 486561
rect 436876 479561 437196 486325
rect 436876 479325 436918 479561
rect 437154 479325 437196 479561
rect 436876 472561 437196 479325
rect 436876 472325 436918 472561
rect 437154 472325 437196 472561
rect 436876 465561 437196 472325
rect 436876 465325 436918 465561
rect 437154 465325 437196 465561
rect 436876 458561 437196 465325
rect 436876 458325 436918 458561
rect 437154 458325 437196 458561
rect 436876 451561 437196 458325
rect 436876 451325 436918 451561
rect 437154 451325 437196 451561
rect 436876 444561 437196 451325
rect 436876 444325 436918 444561
rect 437154 444325 437196 444561
rect 436876 437561 437196 444325
rect 436876 437325 436918 437561
rect 437154 437325 437196 437561
rect 436876 430561 437196 437325
rect 436876 430325 436918 430561
rect 437154 430325 437196 430561
rect 436876 423561 437196 430325
rect 436876 423325 436918 423561
rect 437154 423325 437196 423561
rect 436876 416561 437196 423325
rect 436876 416325 436918 416561
rect 437154 416325 437196 416561
rect 436876 409561 437196 416325
rect 436876 409325 436918 409561
rect 437154 409325 437196 409561
rect 436876 402561 437196 409325
rect 436876 402325 436918 402561
rect 437154 402325 437196 402561
rect 436876 395561 437196 402325
rect 436876 395325 436918 395561
rect 437154 395325 437196 395561
rect 436876 388561 437196 395325
rect 436876 388325 436918 388561
rect 437154 388325 437196 388561
rect 436876 381561 437196 388325
rect 436876 381325 436918 381561
rect 437154 381325 437196 381561
rect 436876 374561 437196 381325
rect 436876 374325 436918 374561
rect 437154 374325 437196 374561
rect 436876 367561 437196 374325
rect 436876 367325 436918 367561
rect 437154 367325 437196 367561
rect 436876 360561 437196 367325
rect 436876 360325 436918 360561
rect 437154 360325 437196 360561
rect 436876 353561 437196 360325
rect 436876 353325 436918 353561
rect 437154 353325 437196 353561
rect 436876 346561 437196 353325
rect 436876 346325 436918 346561
rect 437154 346325 437196 346561
rect 436876 339561 437196 346325
rect 436876 339325 436918 339561
rect 437154 339325 437196 339561
rect 436876 332561 437196 339325
rect 436876 332325 436918 332561
rect 437154 332325 437196 332561
rect 436876 325561 437196 332325
rect 436876 325325 436918 325561
rect 437154 325325 437196 325561
rect 436876 318561 437196 325325
rect 436876 318325 436918 318561
rect 437154 318325 437196 318561
rect 436876 311561 437196 318325
rect 436876 311325 436918 311561
rect 437154 311325 437196 311561
rect 436876 304561 437196 311325
rect 436876 304325 436918 304561
rect 437154 304325 437196 304561
rect 436876 297561 437196 304325
rect 436876 297325 436918 297561
rect 437154 297325 437196 297561
rect 436876 290561 437196 297325
rect 436876 290325 436918 290561
rect 437154 290325 437196 290561
rect 436876 283561 437196 290325
rect 436876 283325 436918 283561
rect 437154 283325 437196 283561
rect 436876 276561 437196 283325
rect 436876 276325 436918 276561
rect 437154 276325 437196 276561
rect 436876 269561 437196 276325
rect 436876 269325 436918 269561
rect 437154 269325 437196 269561
rect 436876 262561 437196 269325
rect 436876 262325 436918 262561
rect 437154 262325 437196 262561
rect 436876 255561 437196 262325
rect 436876 255325 436918 255561
rect 437154 255325 437196 255561
rect 436876 248561 437196 255325
rect 436876 248325 436918 248561
rect 437154 248325 437196 248561
rect 436876 241561 437196 248325
rect 436876 241325 436918 241561
rect 437154 241325 437196 241561
rect 436876 234561 437196 241325
rect 436876 234325 436918 234561
rect 437154 234325 437196 234561
rect 436876 227561 437196 234325
rect 436876 227325 436918 227561
rect 437154 227325 437196 227561
rect 436876 220561 437196 227325
rect 436876 220325 436918 220561
rect 437154 220325 437196 220561
rect 436876 213561 437196 220325
rect 436876 213325 436918 213561
rect 437154 213325 437196 213561
rect 436876 206561 437196 213325
rect 436876 206325 436918 206561
rect 437154 206325 437196 206561
rect 436876 199561 437196 206325
rect 436876 199325 436918 199561
rect 437154 199325 437196 199561
rect 436876 192561 437196 199325
rect 436876 192325 436918 192561
rect 437154 192325 437196 192561
rect 436876 185561 437196 192325
rect 436876 185325 436918 185561
rect 437154 185325 437196 185561
rect 436876 178561 437196 185325
rect 436876 178325 436918 178561
rect 437154 178325 437196 178561
rect 436876 171561 437196 178325
rect 436876 171325 436918 171561
rect 437154 171325 437196 171561
rect 436876 164561 437196 171325
rect 436876 164325 436918 164561
rect 437154 164325 437196 164561
rect 436876 157561 437196 164325
rect 436876 157325 436918 157561
rect 437154 157325 437196 157561
rect 436876 150561 437196 157325
rect 436876 150325 436918 150561
rect 437154 150325 437196 150561
rect 436876 143561 437196 150325
rect 436876 143325 436918 143561
rect 437154 143325 437196 143561
rect 436876 136561 437196 143325
rect 436876 136325 436918 136561
rect 437154 136325 437196 136561
rect 436876 129561 437196 136325
rect 436876 129325 436918 129561
rect 437154 129325 437196 129561
rect 436876 122561 437196 129325
rect 436876 122325 436918 122561
rect 437154 122325 437196 122561
rect 436876 115561 437196 122325
rect 436876 115325 436918 115561
rect 437154 115325 437196 115561
rect 436876 108561 437196 115325
rect 436876 108325 436918 108561
rect 437154 108325 437196 108561
rect 436876 101561 437196 108325
rect 436876 101325 436918 101561
rect 437154 101325 437196 101561
rect 436876 94561 437196 101325
rect 436876 94325 436918 94561
rect 437154 94325 437196 94561
rect 436876 87561 437196 94325
rect 436876 87325 436918 87561
rect 437154 87325 437196 87561
rect 436876 80561 437196 87325
rect 436876 80325 436918 80561
rect 437154 80325 437196 80561
rect 436876 73561 437196 80325
rect 436876 73325 436918 73561
rect 437154 73325 437196 73561
rect 436876 66561 437196 73325
rect 436876 66325 436918 66561
rect 437154 66325 437196 66561
rect 436876 59561 437196 66325
rect 436876 59325 436918 59561
rect 437154 59325 437196 59561
rect 436876 52561 437196 59325
rect 436876 52325 436918 52561
rect 437154 52325 437196 52561
rect 436876 45561 437196 52325
rect 436876 45325 436918 45561
rect 437154 45325 437196 45561
rect 436876 38561 437196 45325
rect 436876 38325 436918 38561
rect 437154 38325 437196 38561
rect 436876 31561 437196 38325
rect 436876 31325 436918 31561
rect 437154 31325 437196 31561
rect 436876 24561 437196 31325
rect 436876 24325 436918 24561
rect 437154 24325 437196 24561
rect 436876 17561 437196 24325
rect 436876 17325 436918 17561
rect 437154 17325 437196 17561
rect 436876 10561 437196 17325
rect 436876 10325 436918 10561
rect 437154 10325 437196 10561
rect 436876 3561 437196 10325
rect 436876 3325 436918 3561
rect 437154 3325 437196 3561
rect 436876 -1706 437196 3325
rect 436876 -1942 436918 -1706
rect 437154 -1942 437196 -1706
rect 436876 -2026 437196 -1942
rect 436876 -2262 436918 -2026
rect 437154 -2262 437196 -2026
rect 436876 -2294 437196 -2262
rect 442144 705238 442464 706230
rect 442144 705002 442186 705238
rect 442422 705002 442464 705238
rect 442144 704918 442464 705002
rect 442144 704682 442186 704918
rect 442422 704682 442464 704918
rect 442144 695494 442464 704682
rect 442144 695258 442186 695494
rect 442422 695258 442464 695494
rect 442144 688494 442464 695258
rect 442144 688258 442186 688494
rect 442422 688258 442464 688494
rect 442144 681494 442464 688258
rect 442144 681258 442186 681494
rect 442422 681258 442464 681494
rect 442144 674494 442464 681258
rect 442144 674258 442186 674494
rect 442422 674258 442464 674494
rect 442144 667494 442464 674258
rect 442144 667258 442186 667494
rect 442422 667258 442464 667494
rect 442144 660494 442464 667258
rect 442144 660258 442186 660494
rect 442422 660258 442464 660494
rect 442144 653494 442464 660258
rect 442144 653258 442186 653494
rect 442422 653258 442464 653494
rect 442144 646494 442464 653258
rect 442144 646258 442186 646494
rect 442422 646258 442464 646494
rect 442144 639494 442464 646258
rect 442144 639258 442186 639494
rect 442422 639258 442464 639494
rect 442144 632494 442464 639258
rect 442144 632258 442186 632494
rect 442422 632258 442464 632494
rect 442144 625494 442464 632258
rect 442144 625258 442186 625494
rect 442422 625258 442464 625494
rect 442144 618494 442464 625258
rect 442144 618258 442186 618494
rect 442422 618258 442464 618494
rect 442144 611494 442464 618258
rect 442144 611258 442186 611494
rect 442422 611258 442464 611494
rect 442144 604494 442464 611258
rect 442144 604258 442186 604494
rect 442422 604258 442464 604494
rect 442144 597494 442464 604258
rect 442144 597258 442186 597494
rect 442422 597258 442464 597494
rect 442144 590494 442464 597258
rect 442144 590258 442186 590494
rect 442422 590258 442464 590494
rect 442144 583494 442464 590258
rect 442144 583258 442186 583494
rect 442422 583258 442464 583494
rect 442144 576494 442464 583258
rect 442144 576258 442186 576494
rect 442422 576258 442464 576494
rect 442144 569494 442464 576258
rect 442144 569258 442186 569494
rect 442422 569258 442464 569494
rect 442144 562494 442464 569258
rect 442144 562258 442186 562494
rect 442422 562258 442464 562494
rect 442144 555494 442464 562258
rect 442144 555258 442186 555494
rect 442422 555258 442464 555494
rect 442144 548494 442464 555258
rect 442144 548258 442186 548494
rect 442422 548258 442464 548494
rect 442144 541494 442464 548258
rect 442144 541258 442186 541494
rect 442422 541258 442464 541494
rect 442144 534494 442464 541258
rect 442144 534258 442186 534494
rect 442422 534258 442464 534494
rect 442144 527494 442464 534258
rect 442144 527258 442186 527494
rect 442422 527258 442464 527494
rect 442144 520494 442464 527258
rect 442144 520258 442186 520494
rect 442422 520258 442464 520494
rect 442144 513494 442464 520258
rect 442144 513258 442186 513494
rect 442422 513258 442464 513494
rect 442144 506494 442464 513258
rect 442144 506258 442186 506494
rect 442422 506258 442464 506494
rect 442144 499494 442464 506258
rect 442144 499258 442186 499494
rect 442422 499258 442464 499494
rect 442144 492494 442464 499258
rect 442144 492258 442186 492494
rect 442422 492258 442464 492494
rect 442144 485494 442464 492258
rect 442144 485258 442186 485494
rect 442422 485258 442464 485494
rect 442144 478494 442464 485258
rect 442144 478258 442186 478494
rect 442422 478258 442464 478494
rect 442144 471494 442464 478258
rect 442144 471258 442186 471494
rect 442422 471258 442464 471494
rect 442144 464494 442464 471258
rect 442144 464258 442186 464494
rect 442422 464258 442464 464494
rect 442144 457494 442464 464258
rect 442144 457258 442186 457494
rect 442422 457258 442464 457494
rect 442144 450494 442464 457258
rect 442144 450258 442186 450494
rect 442422 450258 442464 450494
rect 442144 443494 442464 450258
rect 442144 443258 442186 443494
rect 442422 443258 442464 443494
rect 442144 436494 442464 443258
rect 442144 436258 442186 436494
rect 442422 436258 442464 436494
rect 442144 429494 442464 436258
rect 442144 429258 442186 429494
rect 442422 429258 442464 429494
rect 442144 422494 442464 429258
rect 442144 422258 442186 422494
rect 442422 422258 442464 422494
rect 442144 415494 442464 422258
rect 442144 415258 442186 415494
rect 442422 415258 442464 415494
rect 442144 408494 442464 415258
rect 442144 408258 442186 408494
rect 442422 408258 442464 408494
rect 442144 401494 442464 408258
rect 442144 401258 442186 401494
rect 442422 401258 442464 401494
rect 442144 394494 442464 401258
rect 442144 394258 442186 394494
rect 442422 394258 442464 394494
rect 442144 387494 442464 394258
rect 442144 387258 442186 387494
rect 442422 387258 442464 387494
rect 442144 380494 442464 387258
rect 442144 380258 442186 380494
rect 442422 380258 442464 380494
rect 442144 373494 442464 380258
rect 442144 373258 442186 373494
rect 442422 373258 442464 373494
rect 442144 366494 442464 373258
rect 442144 366258 442186 366494
rect 442422 366258 442464 366494
rect 442144 359494 442464 366258
rect 442144 359258 442186 359494
rect 442422 359258 442464 359494
rect 442144 352494 442464 359258
rect 442144 352258 442186 352494
rect 442422 352258 442464 352494
rect 442144 345494 442464 352258
rect 442144 345258 442186 345494
rect 442422 345258 442464 345494
rect 442144 338494 442464 345258
rect 442144 338258 442186 338494
rect 442422 338258 442464 338494
rect 442144 331494 442464 338258
rect 442144 331258 442186 331494
rect 442422 331258 442464 331494
rect 442144 324494 442464 331258
rect 442144 324258 442186 324494
rect 442422 324258 442464 324494
rect 442144 317494 442464 324258
rect 442144 317258 442186 317494
rect 442422 317258 442464 317494
rect 442144 310494 442464 317258
rect 442144 310258 442186 310494
rect 442422 310258 442464 310494
rect 442144 303494 442464 310258
rect 442144 303258 442186 303494
rect 442422 303258 442464 303494
rect 442144 296494 442464 303258
rect 442144 296258 442186 296494
rect 442422 296258 442464 296494
rect 442144 289494 442464 296258
rect 442144 289258 442186 289494
rect 442422 289258 442464 289494
rect 442144 282494 442464 289258
rect 442144 282258 442186 282494
rect 442422 282258 442464 282494
rect 442144 275494 442464 282258
rect 442144 275258 442186 275494
rect 442422 275258 442464 275494
rect 442144 268494 442464 275258
rect 442144 268258 442186 268494
rect 442422 268258 442464 268494
rect 442144 261494 442464 268258
rect 442144 261258 442186 261494
rect 442422 261258 442464 261494
rect 442144 254494 442464 261258
rect 442144 254258 442186 254494
rect 442422 254258 442464 254494
rect 442144 247494 442464 254258
rect 442144 247258 442186 247494
rect 442422 247258 442464 247494
rect 442144 240494 442464 247258
rect 442144 240258 442186 240494
rect 442422 240258 442464 240494
rect 442144 233494 442464 240258
rect 442144 233258 442186 233494
rect 442422 233258 442464 233494
rect 442144 226494 442464 233258
rect 442144 226258 442186 226494
rect 442422 226258 442464 226494
rect 442144 219494 442464 226258
rect 442144 219258 442186 219494
rect 442422 219258 442464 219494
rect 442144 212494 442464 219258
rect 442144 212258 442186 212494
rect 442422 212258 442464 212494
rect 442144 205494 442464 212258
rect 442144 205258 442186 205494
rect 442422 205258 442464 205494
rect 442144 198494 442464 205258
rect 442144 198258 442186 198494
rect 442422 198258 442464 198494
rect 442144 191494 442464 198258
rect 442144 191258 442186 191494
rect 442422 191258 442464 191494
rect 442144 184494 442464 191258
rect 442144 184258 442186 184494
rect 442422 184258 442464 184494
rect 442144 177494 442464 184258
rect 442144 177258 442186 177494
rect 442422 177258 442464 177494
rect 442144 170494 442464 177258
rect 442144 170258 442186 170494
rect 442422 170258 442464 170494
rect 442144 163494 442464 170258
rect 442144 163258 442186 163494
rect 442422 163258 442464 163494
rect 442144 156494 442464 163258
rect 442144 156258 442186 156494
rect 442422 156258 442464 156494
rect 442144 149494 442464 156258
rect 442144 149258 442186 149494
rect 442422 149258 442464 149494
rect 442144 142494 442464 149258
rect 442144 142258 442186 142494
rect 442422 142258 442464 142494
rect 442144 135494 442464 142258
rect 442144 135258 442186 135494
rect 442422 135258 442464 135494
rect 442144 128494 442464 135258
rect 442144 128258 442186 128494
rect 442422 128258 442464 128494
rect 442144 121494 442464 128258
rect 442144 121258 442186 121494
rect 442422 121258 442464 121494
rect 442144 114494 442464 121258
rect 442144 114258 442186 114494
rect 442422 114258 442464 114494
rect 442144 107494 442464 114258
rect 442144 107258 442186 107494
rect 442422 107258 442464 107494
rect 442144 100494 442464 107258
rect 442144 100258 442186 100494
rect 442422 100258 442464 100494
rect 442144 93494 442464 100258
rect 442144 93258 442186 93494
rect 442422 93258 442464 93494
rect 442144 86494 442464 93258
rect 442144 86258 442186 86494
rect 442422 86258 442464 86494
rect 442144 79494 442464 86258
rect 442144 79258 442186 79494
rect 442422 79258 442464 79494
rect 442144 72494 442464 79258
rect 442144 72258 442186 72494
rect 442422 72258 442464 72494
rect 442144 65494 442464 72258
rect 442144 65258 442186 65494
rect 442422 65258 442464 65494
rect 442144 58494 442464 65258
rect 442144 58258 442186 58494
rect 442422 58258 442464 58494
rect 442144 51494 442464 58258
rect 442144 51258 442186 51494
rect 442422 51258 442464 51494
rect 442144 44494 442464 51258
rect 442144 44258 442186 44494
rect 442422 44258 442464 44494
rect 442144 37494 442464 44258
rect 442144 37258 442186 37494
rect 442422 37258 442464 37494
rect 442144 30494 442464 37258
rect 442144 30258 442186 30494
rect 442422 30258 442464 30494
rect 442144 23494 442464 30258
rect 442144 23258 442186 23494
rect 442422 23258 442464 23494
rect 442144 16494 442464 23258
rect 442144 16258 442186 16494
rect 442422 16258 442464 16494
rect 442144 9494 442464 16258
rect 442144 9258 442186 9494
rect 442422 9258 442464 9494
rect 442144 2494 442464 9258
rect 442144 2258 442186 2494
rect 442422 2258 442464 2494
rect 442144 -746 442464 2258
rect 442144 -982 442186 -746
rect 442422 -982 442464 -746
rect 442144 -1066 442464 -982
rect 442144 -1302 442186 -1066
rect 442422 -1302 442464 -1066
rect 442144 -2294 442464 -1302
rect 443876 706198 444196 706230
rect 443876 705962 443918 706198
rect 444154 705962 444196 706198
rect 443876 705878 444196 705962
rect 443876 705642 443918 705878
rect 444154 705642 444196 705878
rect 443876 696561 444196 705642
rect 443876 696325 443918 696561
rect 444154 696325 444196 696561
rect 443876 689561 444196 696325
rect 443876 689325 443918 689561
rect 444154 689325 444196 689561
rect 443876 682561 444196 689325
rect 443876 682325 443918 682561
rect 444154 682325 444196 682561
rect 443876 675561 444196 682325
rect 443876 675325 443918 675561
rect 444154 675325 444196 675561
rect 443876 668561 444196 675325
rect 443876 668325 443918 668561
rect 444154 668325 444196 668561
rect 443876 661561 444196 668325
rect 443876 661325 443918 661561
rect 444154 661325 444196 661561
rect 443876 654561 444196 661325
rect 443876 654325 443918 654561
rect 444154 654325 444196 654561
rect 443876 647561 444196 654325
rect 443876 647325 443918 647561
rect 444154 647325 444196 647561
rect 443876 640561 444196 647325
rect 443876 640325 443918 640561
rect 444154 640325 444196 640561
rect 443876 633561 444196 640325
rect 443876 633325 443918 633561
rect 444154 633325 444196 633561
rect 443876 626561 444196 633325
rect 443876 626325 443918 626561
rect 444154 626325 444196 626561
rect 443876 619561 444196 626325
rect 443876 619325 443918 619561
rect 444154 619325 444196 619561
rect 443876 612561 444196 619325
rect 443876 612325 443918 612561
rect 444154 612325 444196 612561
rect 443876 605561 444196 612325
rect 443876 605325 443918 605561
rect 444154 605325 444196 605561
rect 443876 598561 444196 605325
rect 443876 598325 443918 598561
rect 444154 598325 444196 598561
rect 443876 591561 444196 598325
rect 443876 591325 443918 591561
rect 444154 591325 444196 591561
rect 443876 584561 444196 591325
rect 443876 584325 443918 584561
rect 444154 584325 444196 584561
rect 443876 577561 444196 584325
rect 443876 577325 443918 577561
rect 444154 577325 444196 577561
rect 443876 570561 444196 577325
rect 443876 570325 443918 570561
rect 444154 570325 444196 570561
rect 443876 563561 444196 570325
rect 443876 563325 443918 563561
rect 444154 563325 444196 563561
rect 443876 556561 444196 563325
rect 443876 556325 443918 556561
rect 444154 556325 444196 556561
rect 443876 549561 444196 556325
rect 443876 549325 443918 549561
rect 444154 549325 444196 549561
rect 443876 542561 444196 549325
rect 443876 542325 443918 542561
rect 444154 542325 444196 542561
rect 443876 535561 444196 542325
rect 443876 535325 443918 535561
rect 444154 535325 444196 535561
rect 443876 528561 444196 535325
rect 443876 528325 443918 528561
rect 444154 528325 444196 528561
rect 443876 521561 444196 528325
rect 443876 521325 443918 521561
rect 444154 521325 444196 521561
rect 443876 514561 444196 521325
rect 443876 514325 443918 514561
rect 444154 514325 444196 514561
rect 443876 507561 444196 514325
rect 443876 507325 443918 507561
rect 444154 507325 444196 507561
rect 443876 500561 444196 507325
rect 443876 500325 443918 500561
rect 444154 500325 444196 500561
rect 443876 493561 444196 500325
rect 443876 493325 443918 493561
rect 444154 493325 444196 493561
rect 443876 486561 444196 493325
rect 443876 486325 443918 486561
rect 444154 486325 444196 486561
rect 443876 479561 444196 486325
rect 443876 479325 443918 479561
rect 444154 479325 444196 479561
rect 443876 472561 444196 479325
rect 443876 472325 443918 472561
rect 444154 472325 444196 472561
rect 443876 465561 444196 472325
rect 443876 465325 443918 465561
rect 444154 465325 444196 465561
rect 443876 458561 444196 465325
rect 443876 458325 443918 458561
rect 444154 458325 444196 458561
rect 443876 451561 444196 458325
rect 443876 451325 443918 451561
rect 444154 451325 444196 451561
rect 443876 444561 444196 451325
rect 443876 444325 443918 444561
rect 444154 444325 444196 444561
rect 443876 437561 444196 444325
rect 443876 437325 443918 437561
rect 444154 437325 444196 437561
rect 443876 430561 444196 437325
rect 443876 430325 443918 430561
rect 444154 430325 444196 430561
rect 443876 423561 444196 430325
rect 443876 423325 443918 423561
rect 444154 423325 444196 423561
rect 443876 416561 444196 423325
rect 443876 416325 443918 416561
rect 444154 416325 444196 416561
rect 443876 409561 444196 416325
rect 443876 409325 443918 409561
rect 444154 409325 444196 409561
rect 443876 402561 444196 409325
rect 443876 402325 443918 402561
rect 444154 402325 444196 402561
rect 443876 395561 444196 402325
rect 443876 395325 443918 395561
rect 444154 395325 444196 395561
rect 443876 388561 444196 395325
rect 443876 388325 443918 388561
rect 444154 388325 444196 388561
rect 443876 381561 444196 388325
rect 443876 381325 443918 381561
rect 444154 381325 444196 381561
rect 443876 374561 444196 381325
rect 443876 374325 443918 374561
rect 444154 374325 444196 374561
rect 443876 367561 444196 374325
rect 443876 367325 443918 367561
rect 444154 367325 444196 367561
rect 443876 360561 444196 367325
rect 443876 360325 443918 360561
rect 444154 360325 444196 360561
rect 443876 353561 444196 360325
rect 443876 353325 443918 353561
rect 444154 353325 444196 353561
rect 443876 346561 444196 353325
rect 443876 346325 443918 346561
rect 444154 346325 444196 346561
rect 443876 339561 444196 346325
rect 443876 339325 443918 339561
rect 444154 339325 444196 339561
rect 443876 332561 444196 339325
rect 443876 332325 443918 332561
rect 444154 332325 444196 332561
rect 443876 325561 444196 332325
rect 443876 325325 443918 325561
rect 444154 325325 444196 325561
rect 443876 318561 444196 325325
rect 443876 318325 443918 318561
rect 444154 318325 444196 318561
rect 443876 311561 444196 318325
rect 443876 311325 443918 311561
rect 444154 311325 444196 311561
rect 443876 304561 444196 311325
rect 443876 304325 443918 304561
rect 444154 304325 444196 304561
rect 443876 297561 444196 304325
rect 443876 297325 443918 297561
rect 444154 297325 444196 297561
rect 443876 290561 444196 297325
rect 443876 290325 443918 290561
rect 444154 290325 444196 290561
rect 443876 283561 444196 290325
rect 443876 283325 443918 283561
rect 444154 283325 444196 283561
rect 443876 276561 444196 283325
rect 443876 276325 443918 276561
rect 444154 276325 444196 276561
rect 443876 269561 444196 276325
rect 443876 269325 443918 269561
rect 444154 269325 444196 269561
rect 443876 262561 444196 269325
rect 443876 262325 443918 262561
rect 444154 262325 444196 262561
rect 443876 255561 444196 262325
rect 443876 255325 443918 255561
rect 444154 255325 444196 255561
rect 443876 248561 444196 255325
rect 443876 248325 443918 248561
rect 444154 248325 444196 248561
rect 443876 241561 444196 248325
rect 443876 241325 443918 241561
rect 444154 241325 444196 241561
rect 443876 234561 444196 241325
rect 443876 234325 443918 234561
rect 444154 234325 444196 234561
rect 443876 227561 444196 234325
rect 443876 227325 443918 227561
rect 444154 227325 444196 227561
rect 443876 220561 444196 227325
rect 443876 220325 443918 220561
rect 444154 220325 444196 220561
rect 443876 213561 444196 220325
rect 443876 213325 443918 213561
rect 444154 213325 444196 213561
rect 443876 206561 444196 213325
rect 443876 206325 443918 206561
rect 444154 206325 444196 206561
rect 443876 199561 444196 206325
rect 443876 199325 443918 199561
rect 444154 199325 444196 199561
rect 443876 192561 444196 199325
rect 443876 192325 443918 192561
rect 444154 192325 444196 192561
rect 443876 185561 444196 192325
rect 443876 185325 443918 185561
rect 444154 185325 444196 185561
rect 443876 178561 444196 185325
rect 443876 178325 443918 178561
rect 444154 178325 444196 178561
rect 443876 171561 444196 178325
rect 443876 171325 443918 171561
rect 444154 171325 444196 171561
rect 443876 164561 444196 171325
rect 443876 164325 443918 164561
rect 444154 164325 444196 164561
rect 443876 157561 444196 164325
rect 443876 157325 443918 157561
rect 444154 157325 444196 157561
rect 443876 150561 444196 157325
rect 443876 150325 443918 150561
rect 444154 150325 444196 150561
rect 443876 143561 444196 150325
rect 443876 143325 443918 143561
rect 444154 143325 444196 143561
rect 443876 136561 444196 143325
rect 443876 136325 443918 136561
rect 444154 136325 444196 136561
rect 443876 129561 444196 136325
rect 443876 129325 443918 129561
rect 444154 129325 444196 129561
rect 443876 122561 444196 129325
rect 443876 122325 443918 122561
rect 444154 122325 444196 122561
rect 443876 115561 444196 122325
rect 443876 115325 443918 115561
rect 444154 115325 444196 115561
rect 443876 108561 444196 115325
rect 443876 108325 443918 108561
rect 444154 108325 444196 108561
rect 443876 101561 444196 108325
rect 443876 101325 443918 101561
rect 444154 101325 444196 101561
rect 443876 94561 444196 101325
rect 443876 94325 443918 94561
rect 444154 94325 444196 94561
rect 443876 87561 444196 94325
rect 443876 87325 443918 87561
rect 444154 87325 444196 87561
rect 443876 80561 444196 87325
rect 443876 80325 443918 80561
rect 444154 80325 444196 80561
rect 443876 73561 444196 80325
rect 443876 73325 443918 73561
rect 444154 73325 444196 73561
rect 443876 66561 444196 73325
rect 443876 66325 443918 66561
rect 444154 66325 444196 66561
rect 443876 59561 444196 66325
rect 443876 59325 443918 59561
rect 444154 59325 444196 59561
rect 443876 52561 444196 59325
rect 443876 52325 443918 52561
rect 444154 52325 444196 52561
rect 443876 45561 444196 52325
rect 443876 45325 443918 45561
rect 444154 45325 444196 45561
rect 443876 38561 444196 45325
rect 443876 38325 443918 38561
rect 444154 38325 444196 38561
rect 443876 31561 444196 38325
rect 443876 31325 443918 31561
rect 444154 31325 444196 31561
rect 443876 24561 444196 31325
rect 443876 24325 443918 24561
rect 444154 24325 444196 24561
rect 443876 17561 444196 24325
rect 443876 17325 443918 17561
rect 444154 17325 444196 17561
rect 443876 10561 444196 17325
rect 443876 10325 443918 10561
rect 444154 10325 444196 10561
rect 443876 3561 444196 10325
rect 443876 3325 443918 3561
rect 444154 3325 444196 3561
rect 443876 -1706 444196 3325
rect 443876 -1942 443918 -1706
rect 444154 -1942 444196 -1706
rect 443876 -2026 444196 -1942
rect 443876 -2262 443918 -2026
rect 444154 -2262 444196 -2026
rect 443876 -2294 444196 -2262
rect 449144 705238 449464 706230
rect 449144 705002 449186 705238
rect 449422 705002 449464 705238
rect 449144 704918 449464 705002
rect 449144 704682 449186 704918
rect 449422 704682 449464 704918
rect 449144 695494 449464 704682
rect 449144 695258 449186 695494
rect 449422 695258 449464 695494
rect 449144 688494 449464 695258
rect 449144 688258 449186 688494
rect 449422 688258 449464 688494
rect 449144 681494 449464 688258
rect 449144 681258 449186 681494
rect 449422 681258 449464 681494
rect 449144 674494 449464 681258
rect 449144 674258 449186 674494
rect 449422 674258 449464 674494
rect 449144 667494 449464 674258
rect 449144 667258 449186 667494
rect 449422 667258 449464 667494
rect 449144 660494 449464 667258
rect 449144 660258 449186 660494
rect 449422 660258 449464 660494
rect 449144 653494 449464 660258
rect 449144 653258 449186 653494
rect 449422 653258 449464 653494
rect 449144 646494 449464 653258
rect 449144 646258 449186 646494
rect 449422 646258 449464 646494
rect 449144 639494 449464 646258
rect 449144 639258 449186 639494
rect 449422 639258 449464 639494
rect 449144 632494 449464 639258
rect 449144 632258 449186 632494
rect 449422 632258 449464 632494
rect 449144 625494 449464 632258
rect 449144 625258 449186 625494
rect 449422 625258 449464 625494
rect 449144 618494 449464 625258
rect 449144 618258 449186 618494
rect 449422 618258 449464 618494
rect 449144 611494 449464 618258
rect 449144 611258 449186 611494
rect 449422 611258 449464 611494
rect 449144 604494 449464 611258
rect 449144 604258 449186 604494
rect 449422 604258 449464 604494
rect 449144 597494 449464 604258
rect 449144 597258 449186 597494
rect 449422 597258 449464 597494
rect 449144 590494 449464 597258
rect 449144 590258 449186 590494
rect 449422 590258 449464 590494
rect 449144 583494 449464 590258
rect 449144 583258 449186 583494
rect 449422 583258 449464 583494
rect 449144 576494 449464 583258
rect 449144 576258 449186 576494
rect 449422 576258 449464 576494
rect 449144 569494 449464 576258
rect 449144 569258 449186 569494
rect 449422 569258 449464 569494
rect 449144 562494 449464 569258
rect 449144 562258 449186 562494
rect 449422 562258 449464 562494
rect 449144 555494 449464 562258
rect 449144 555258 449186 555494
rect 449422 555258 449464 555494
rect 449144 548494 449464 555258
rect 449144 548258 449186 548494
rect 449422 548258 449464 548494
rect 449144 541494 449464 548258
rect 449144 541258 449186 541494
rect 449422 541258 449464 541494
rect 449144 534494 449464 541258
rect 449144 534258 449186 534494
rect 449422 534258 449464 534494
rect 449144 527494 449464 534258
rect 449144 527258 449186 527494
rect 449422 527258 449464 527494
rect 449144 520494 449464 527258
rect 449144 520258 449186 520494
rect 449422 520258 449464 520494
rect 449144 513494 449464 520258
rect 449144 513258 449186 513494
rect 449422 513258 449464 513494
rect 449144 506494 449464 513258
rect 449144 506258 449186 506494
rect 449422 506258 449464 506494
rect 449144 499494 449464 506258
rect 449144 499258 449186 499494
rect 449422 499258 449464 499494
rect 449144 492494 449464 499258
rect 449144 492258 449186 492494
rect 449422 492258 449464 492494
rect 449144 485494 449464 492258
rect 449144 485258 449186 485494
rect 449422 485258 449464 485494
rect 449144 478494 449464 485258
rect 449144 478258 449186 478494
rect 449422 478258 449464 478494
rect 449144 471494 449464 478258
rect 449144 471258 449186 471494
rect 449422 471258 449464 471494
rect 449144 464494 449464 471258
rect 449144 464258 449186 464494
rect 449422 464258 449464 464494
rect 449144 457494 449464 464258
rect 449144 457258 449186 457494
rect 449422 457258 449464 457494
rect 449144 450494 449464 457258
rect 449144 450258 449186 450494
rect 449422 450258 449464 450494
rect 449144 443494 449464 450258
rect 449144 443258 449186 443494
rect 449422 443258 449464 443494
rect 449144 436494 449464 443258
rect 449144 436258 449186 436494
rect 449422 436258 449464 436494
rect 449144 429494 449464 436258
rect 449144 429258 449186 429494
rect 449422 429258 449464 429494
rect 449144 422494 449464 429258
rect 449144 422258 449186 422494
rect 449422 422258 449464 422494
rect 449144 415494 449464 422258
rect 449144 415258 449186 415494
rect 449422 415258 449464 415494
rect 449144 408494 449464 415258
rect 449144 408258 449186 408494
rect 449422 408258 449464 408494
rect 449144 401494 449464 408258
rect 449144 401258 449186 401494
rect 449422 401258 449464 401494
rect 449144 394494 449464 401258
rect 449144 394258 449186 394494
rect 449422 394258 449464 394494
rect 449144 387494 449464 394258
rect 449144 387258 449186 387494
rect 449422 387258 449464 387494
rect 449144 380494 449464 387258
rect 449144 380258 449186 380494
rect 449422 380258 449464 380494
rect 449144 373494 449464 380258
rect 449144 373258 449186 373494
rect 449422 373258 449464 373494
rect 449144 366494 449464 373258
rect 449144 366258 449186 366494
rect 449422 366258 449464 366494
rect 449144 359494 449464 366258
rect 449144 359258 449186 359494
rect 449422 359258 449464 359494
rect 449144 352494 449464 359258
rect 449144 352258 449186 352494
rect 449422 352258 449464 352494
rect 449144 345494 449464 352258
rect 449144 345258 449186 345494
rect 449422 345258 449464 345494
rect 449144 338494 449464 345258
rect 449144 338258 449186 338494
rect 449422 338258 449464 338494
rect 449144 331494 449464 338258
rect 449144 331258 449186 331494
rect 449422 331258 449464 331494
rect 449144 324494 449464 331258
rect 449144 324258 449186 324494
rect 449422 324258 449464 324494
rect 449144 317494 449464 324258
rect 449144 317258 449186 317494
rect 449422 317258 449464 317494
rect 449144 310494 449464 317258
rect 449144 310258 449186 310494
rect 449422 310258 449464 310494
rect 449144 303494 449464 310258
rect 449144 303258 449186 303494
rect 449422 303258 449464 303494
rect 449144 296494 449464 303258
rect 449144 296258 449186 296494
rect 449422 296258 449464 296494
rect 449144 289494 449464 296258
rect 449144 289258 449186 289494
rect 449422 289258 449464 289494
rect 449144 282494 449464 289258
rect 449144 282258 449186 282494
rect 449422 282258 449464 282494
rect 449144 275494 449464 282258
rect 449144 275258 449186 275494
rect 449422 275258 449464 275494
rect 449144 268494 449464 275258
rect 449144 268258 449186 268494
rect 449422 268258 449464 268494
rect 449144 261494 449464 268258
rect 449144 261258 449186 261494
rect 449422 261258 449464 261494
rect 449144 254494 449464 261258
rect 449144 254258 449186 254494
rect 449422 254258 449464 254494
rect 449144 247494 449464 254258
rect 449144 247258 449186 247494
rect 449422 247258 449464 247494
rect 449144 240494 449464 247258
rect 449144 240258 449186 240494
rect 449422 240258 449464 240494
rect 449144 233494 449464 240258
rect 449144 233258 449186 233494
rect 449422 233258 449464 233494
rect 449144 226494 449464 233258
rect 449144 226258 449186 226494
rect 449422 226258 449464 226494
rect 449144 219494 449464 226258
rect 449144 219258 449186 219494
rect 449422 219258 449464 219494
rect 449144 212494 449464 219258
rect 449144 212258 449186 212494
rect 449422 212258 449464 212494
rect 449144 205494 449464 212258
rect 449144 205258 449186 205494
rect 449422 205258 449464 205494
rect 449144 198494 449464 205258
rect 449144 198258 449186 198494
rect 449422 198258 449464 198494
rect 449144 191494 449464 198258
rect 449144 191258 449186 191494
rect 449422 191258 449464 191494
rect 449144 184494 449464 191258
rect 449144 184258 449186 184494
rect 449422 184258 449464 184494
rect 449144 177494 449464 184258
rect 449144 177258 449186 177494
rect 449422 177258 449464 177494
rect 449144 170494 449464 177258
rect 449144 170258 449186 170494
rect 449422 170258 449464 170494
rect 449144 163494 449464 170258
rect 449144 163258 449186 163494
rect 449422 163258 449464 163494
rect 449144 156494 449464 163258
rect 449144 156258 449186 156494
rect 449422 156258 449464 156494
rect 449144 149494 449464 156258
rect 449144 149258 449186 149494
rect 449422 149258 449464 149494
rect 449144 142494 449464 149258
rect 449144 142258 449186 142494
rect 449422 142258 449464 142494
rect 449144 135494 449464 142258
rect 449144 135258 449186 135494
rect 449422 135258 449464 135494
rect 449144 128494 449464 135258
rect 449144 128258 449186 128494
rect 449422 128258 449464 128494
rect 449144 121494 449464 128258
rect 449144 121258 449186 121494
rect 449422 121258 449464 121494
rect 449144 114494 449464 121258
rect 449144 114258 449186 114494
rect 449422 114258 449464 114494
rect 449144 107494 449464 114258
rect 449144 107258 449186 107494
rect 449422 107258 449464 107494
rect 449144 100494 449464 107258
rect 449144 100258 449186 100494
rect 449422 100258 449464 100494
rect 449144 93494 449464 100258
rect 449144 93258 449186 93494
rect 449422 93258 449464 93494
rect 449144 86494 449464 93258
rect 449144 86258 449186 86494
rect 449422 86258 449464 86494
rect 449144 79494 449464 86258
rect 449144 79258 449186 79494
rect 449422 79258 449464 79494
rect 449144 72494 449464 79258
rect 449144 72258 449186 72494
rect 449422 72258 449464 72494
rect 449144 65494 449464 72258
rect 449144 65258 449186 65494
rect 449422 65258 449464 65494
rect 449144 58494 449464 65258
rect 449144 58258 449186 58494
rect 449422 58258 449464 58494
rect 449144 51494 449464 58258
rect 449144 51258 449186 51494
rect 449422 51258 449464 51494
rect 449144 44494 449464 51258
rect 449144 44258 449186 44494
rect 449422 44258 449464 44494
rect 449144 37494 449464 44258
rect 449144 37258 449186 37494
rect 449422 37258 449464 37494
rect 449144 30494 449464 37258
rect 449144 30258 449186 30494
rect 449422 30258 449464 30494
rect 449144 23494 449464 30258
rect 449144 23258 449186 23494
rect 449422 23258 449464 23494
rect 449144 16494 449464 23258
rect 449144 16258 449186 16494
rect 449422 16258 449464 16494
rect 449144 9494 449464 16258
rect 449144 9258 449186 9494
rect 449422 9258 449464 9494
rect 449144 2494 449464 9258
rect 449144 2258 449186 2494
rect 449422 2258 449464 2494
rect 449144 -746 449464 2258
rect 449144 -982 449186 -746
rect 449422 -982 449464 -746
rect 449144 -1066 449464 -982
rect 449144 -1302 449186 -1066
rect 449422 -1302 449464 -1066
rect 449144 -2294 449464 -1302
rect 450876 706198 451196 706230
rect 450876 705962 450918 706198
rect 451154 705962 451196 706198
rect 450876 705878 451196 705962
rect 450876 705642 450918 705878
rect 451154 705642 451196 705878
rect 450876 696561 451196 705642
rect 450876 696325 450918 696561
rect 451154 696325 451196 696561
rect 450876 689561 451196 696325
rect 450876 689325 450918 689561
rect 451154 689325 451196 689561
rect 450876 682561 451196 689325
rect 450876 682325 450918 682561
rect 451154 682325 451196 682561
rect 450876 675561 451196 682325
rect 450876 675325 450918 675561
rect 451154 675325 451196 675561
rect 450876 668561 451196 675325
rect 450876 668325 450918 668561
rect 451154 668325 451196 668561
rect 450876 661561 451196 668325
rect 450876 661325 450918 661561
rect 451154 661325 451196 661561
rect 450876 654561 451196 661325
rect 450876 654325 450918 654561
rect 451154 654325 451196 654561
rect 450876 647561 451196 654325
rect 450876 647325 450918 647561
rect 451154 647325 451196 647561
rect 450876 640561 451196 647325
rect 450876 640325 450918 640561
rect 451154 640325 451196 640561
rect 450876 633561 451196 640325
rect 450876 633325 450918 633561
rect 451154 633325 451196 633561
rect 450876 626561 451196 633325
rect 450876 626325 450918 626561
rect 451154 626325 451196 626561
rect 450876 619561 451196 626325
rect 450876 619325 450918 619561
rect 451154 619325 451196 619561
rect 450876 612561 451196 619325
rect 450876 612325 450918 612561
rect 451154 612325 451196 612561
rect 450876 605561 451196 612325
rect 450876 605325 450918 605561
rect 451154 605325 451196 605561
rect 450876 598561 451196 605325
rect 450876 598325 450918 598561
rect 451154 598325 451196 598561
rect 450876 591561 451196 598325
rect 450876 591325 450918 591561
rect 451154 591325 451196 591561
rect 450876 584561 451196 591325
rect 450876 584325 450918 584561
rect 451154 584325 451196 584561
rect 450876 577561 451196 584325
rect 450876 577325 450918 577561
rect 451154 577325 451196 577561
rect 450876 570561 451196 577325
rect 450876 570325 450918 570561
rect 451154 570325 451196 570561
rect 450876 563561 451196 570325
rect 450876 563325 450918 563561
rect 451154 563325 451196 563561
rect 450876 556561 451196 563325
rect 450876 556325 450918 556561
rect 451154 556325 451196 556561
rect 450876 549561 451196 556325
rect 450876 549325 450918 549561
rect 451154 549325 451196 549561
rect 450876 542561 451196 549325
rect 450876 542325 450918 542561
rect 451154 542325 451196 542561
rect 450876 535561 451196 542325
rect 450876 535325 450918 535561
rect 451154 535325 451196 535561
rect 450876 528561 451196 535325
rect 450876 528325 450918 528561
rect 451154 528325 451196 528561
rect 450876 521561 451196 528325
rect 450876 521325 450918 521561
rect 451154 521325 451196 521561
rect 450876 514561 451196 521325
rect 450876 514325 450918 514561
rect 451154 514325 451196 514561
rect 450876 507561 451196 514325
rect 450876 507325 450918 507561
rect 451154 507325 451196 507561
rect 450876 500561 451196 507325
rect 450876 500325 450918 500561
rect 451154 500325 451196 500561
rect 450876 493561 451196 500325
rect 450876 493325 450918 493561
rect 451154 493325 451196 493561
rect 450876 486561 451196 493325
rect 450876 486325 450918 486561
rect 451154 486325 451196 486561
rect 450876 479561 451196 486325
rect 450876 479325 450918 479561
rect 451154 479325 451196 479561
rect 450876 472561 451196 479325
rect 450876 472325 450918 472561
rect 451154 472325 451196 472561
rect 450876 465561 451196 472325
rect 450876 465325 450918 465561
rect 451154 465325 451196 465561
rect 450876 458561 451196 465325
rect 450876 458325 450918 458561
rect 451154 458325 451196 458561
rect 450876 451561 451196 458325
rect 450876 451325 450918 451561
rect 451154 451325 451196 451561
rect 450876 444561 451196 451325
rect 450876 444325 450918 444561
rect 451154 444325 451196 444561
rect 450876 437561 451196 444325
rect 450876 437325 450918 437561
rect 451154 437325 451196 437561
rect 450876 430561 451196 437325
rect 450876 430325 450918 430561
rect 451154 430325 451196 430561
rect 450876 423561 451196 430325
rect 450876 423325 450918 423561
rect 451154 423325 451196 423561
rect 450876 416561 451196 423325
rect 450876 416325 450918 416561
rect 451154 416325 451196 416561
rect 450876 409561 451196 416325
rect 450876 409325 450918 409561
rect 451154 409325 451196 409561
rect 450876 402561 451196 409325
rect 450876 402325 450918 402561
rect 451154 402325 451196 402561
rect 450876 395561 451196 402325
rect 450876 395325 450918 395561
rect 451154 395325 451196 395561
rect 450876 388561 451196 395325
rect 450876 388325 450918 388561
rect 451154 388325 451196 388561
rect 450876 381561 451196 388325
rect 450876 381325 450918 381561
rect 451154 381325 451196 381561
rect 450876 374561 451196 381325
rect 450876 374325 450918 374561
rect 451154 374325 451196 374561
rect 450876 367561 451196 374325
rect 450876 367325 450918 367561
rect 451154 367325 451196 367561
rect 450876 360561 451196 367325
rect 450876 360325 450918 360561
rect 451154 360325 451196 360561
rect 450876 353561 451196 360325
rect 450876 353325 450918 353561
rect 451154 353325 451196 353561
rect 450876 346561 451196 353325
rect 450876 346325 450918 346561
rect 451154 346325 451196 346561
rect 450876 339561 451196 346325
rect 450876 339325 450918 339561
rect 451154 339325 451196 339561
rect 450876 332561 451196 339325
rect 450876 332325 450918 332561
rect 451154 332325 451196 332561
rect 450876 325561 451196 332325
rect 450876 325325 450918 325561
rect 451154 325325 451196 325561
rect 450876 318561 451196 325325
rect 450876 318325 450918 318561
rect 451154 318325 451196 318561
rect 450876 311561 451196 318325
rect 450876 311325 450918 311561
rect 451154 311325 451196 311561
rect 450876 304561 451196 311325
rect 450876 304325 450918 304561
rect 451154 304325 451196 304561
rect 450876 297561 451196 304325
rect 450876 297325 450918 297561
rect 451154 297325 451196 297561
rect 450876 290561 451196 297325
rect 450876 290325 450918 290561
rect 451154 290325 451196 290561
rect 450876 283561 451196 290325
rect 450876 283325 450918 283561
rect 451154 283325 451196 283561
rect 450876 276561 451196 283325
rect 450876 276325 450918 276561
rect 451154 276325 451196 276561
rect 450876 269561 451196 276325
rect 450876 269325 450918 269561
rect 451154 269325 451196 269561
rect 450876 262561 451196 269325
rect 450876 262325 450918 262561
rect 451154 262325 451196 262561
rect 450876 255561 451196 262325
rect 450876 255325 450918 255561
rect 451154 255325 451196 255561
rect 450876 248561 451196 255325
rect 450876 248325 450918 248561
rect 451154 248325 451196 248561
rect 450876 241561 451196 248325
rect 450876 241325 450918 241561
rect 451154 241325 451196 241561
rect 450876 234561 451196 241325
rect 450876 234325 450918 234561
rect 451154 234325 451196 234561
rect 450876 227561 451196 234325
rect 450876 227325 450918 227561
rect 451154 227325 451196 227561
rect 450876 220561 451196 227325
rect 450876 220325 450918 220561
rect 451154 220325 451196 220561
rect 450876 213561 451196 220325
rect 450876 213325 450918 213561
rect 451154 213325 451196 213561
rect 450876 206561 451196 213325
rect 450876 206325 450918 206561
rect 451154 206325 451196 206561
rect 450876 199561 451196 206325
rect 450876 199325 450918 199561
rect 451154 199325 451196 199561
rect 450876 192561 451196 199325
rect 450876 192325 450918 192561
rect 451154 192325 451196 192561
rect 450876 185561 451196 192325
rect 450876 185325 450918 185561
rect 451154 185325 451196 185561
rect 450876 178561 451196 185325
rect 450876 178325 450918 178561
rect 451154 178325 451196 178561
rect 450876 171561 451196 178325
rect 450876 171325 450918 171561
rect 451154 171325 451196 171561
rect 450876 164561 451196 171325
rect 450876 164325 450918 164561
rect 451154 164325 451196 164561
rect 450876 157561 451196 164325
rect 450876 157325 450918 157561
rect 451154 157325 451196 157561
rect 450876 150561 451196 157325
rect 450876 150325 450918 150561
rect 451154 150325 451196 150561
rect 450876 143561 451196 150325
rect 450876 143325 450918 143561
rect 451154 143325 451196 143561
rect 450876 136561 451196 143325
rect 450876 136325 450918 136561
rect 451154 136325 451196 136561
rect 450876 129561 451196 136325
rect 450876 129325 450918 129561
rect 451154 129325 451196 129561
rect 450876 122561 451196 129325
rect 450876 122325 450918 122561
rect 451154 122325 451196 122561
rect 450876 115561 451196 122325
rect 450876 115325 450918 115561
rect 451154 115325 451196 115561
rect 450876 108561 451196 115325
rect 450876 108325 450918 108561
rect 451154 108325 451196 108561
rect 450876 101561 451196 108325
rect 450876 101325 450918 101561
rect 451154 101325 451196 101561
rect 450876 94561 451196 101325
rect 450876 94325 450918 94561
rect 451154 94325 451196 94561
rect 450876 87561 451196 94325
rect 450876 87325 450918 87561
rect 451154 87325 451196 87561
rect 450876 80561 451196 87325
rect 450876 80325 450918 80561
rect 451154 80325 451196 80561
rect 450876 73561 451196 80325
rect 450876 73325 450918 73561
rect 451154 73325 451196 73561
rect 450876 66561 451196 73325
rect 450876 66325 450918 66561
rect 451154 66325 451196 66561
rect 450876 59561 451196 66325
rect 450876 59325 450918 59561
rect 451154 59325 451196 59561
rect 450876 52561 451196 59325
rect 450876 52325 450918 52561
rect 451154 52325 451196 52561
rect 450876 45561 451196 52325
rect 450876 45325 450918 45561
rect 451154 45325 451196 45561
rect 450876 38561 451196 45325
rect 450876 38325 450918 38561
rect 451154 38325 451196 38561
rect 450876 31561 451196 38325
rect 450876 31325 450918 31561
rect 451154 31325 451196 31561
rect 450876 24561 451196 31325
rect 450876 24325 450918 24561
rect 451154 24325 451196 24561
rect 450876 17561 451196 24325
rect 450876 17325 450918 17561
rect 451154 17325 451196 17561
rect 450876 10561 451196 17325
rect 450876 10325 450918 10561
rect 451154 10325 451196 10561
rect 450876 3561 451196 10325
rect 450876 3325 450918 3561
rect 451154 3325 451196 3561
rect 450876 -1706 451196 3325
rect 450876 -1942 450918 -1706
rect 451154 -1942 451196 -1706
rect 450876 -2026 451196 -1942
rect 450876 -2262 450918 -2026
rect 451154 -2262 451196 -2026
rect 450876 -2294 451196 -2262
rect 456144 705238 456464 706230
rect 456144 705002 456186 705238
rect 456422 705002 456464 705238
rect 456144 704918 456464 705002
rect 456144 704682 456186 704918
rect 456422 704682 456464 704918
rect 456144 695494 456464 704682
rect 456144 695258 456186 695494
rect 456422 695258 456464 695494
rect 456144 688494 456464 695258
rect 456144 688258 456186 688494
rect 456422 688258 456464 688494
rect 456144 681494 456464 688258
rect 456144 681258 456186 681494
rect 456422 681258 456464 681494
rect 456144 674494 456464 681258
rect 456144 674258 456186 674494
rect 456422 674258 456464 674494
rect 456144 667494 456464 674258
rect 456144 667258 456186 667494
rect 456422 667258 456464 667494
rect 456144 660494 456464 667258
rect 456144 660258 456186 660494
rect 456422 660258 456464 660494
rect 456144 653494 456464 660258
rect 456144 653258 456186 653494
rect 456422 653258 456464 653494
rect 456144 646494 456464 653258
rect 456144 646258 456186 646494
rect 456422 646258 456464 646494
rect 456144 639494 456464 646258
rect 456144 639258 456186 639494
rect 456422 639258 456464 639494
rect 456144 632494 456464 639258
rect 456144 632258 456186 632494
rect 456422 632258 456464 632494
rect 456144 625494 456464 632258
rect 456144 625258 456186 625494
rect 456422 625258 456464 625494
rect 456144 618494 456464 625258
rect 456144 618258 456186 618494
rect 456422 618258 456464 618494
rect 456144 611494 456464 618258
rect 456144 611258 456186 611494
rect 456422 611258 456464 611494
rect 456144 604494 456464 611258
rect 456144 604258 456186 604494
rect 456422 604258 456464 604494
rect 456144 597494 456464 604258
rect 456144 597258 456186 597494
rect 456422 597258 456464 597494
rect 456144 590494 456464 597258
rect 456144 590258 456186 590494
rect 456422 590258 456464 590494
rect 456144 583494 456464 590258
rect 456144 583258 456186 583494
rect 456422 583258 456464 583494
rect 456144 576494 456464 583258
rect 456144 576258 456186 576494
rect 456422 576258 456464 576494
rect 456144 569494 456464 576258
rect 456144 569258 456186 569494
rect 456422 569258 456464 569494
rect 456144 562494 456464 569258
rect 456144 562258 456186 562494
rect 456422 562258 456464 562494
rect 456144 555494 456464 562258
rect 456144 555258 456186 555494
rect 456422 555258 456464 555494
rect 456144 548494 456464 555258
rect 456144 548258 456186 548494
rect 456422 548258 456464 548494
rect 456144 541494 456464 548258
rect 456144 541258 456186 541494
rect 456422 541258 456464 541494
rect 456144 534494 456464 541258
rect 456144 534258 456186 534494
rect 456422 534258 456464 534494
rect 456144 527494 456464 534258
rect 456144 527258 456186 527494
rect 456422 527258 456464 527494
rect 456144 520494 456464 527258
rect 456144 520258 456186 520494
rect 456422 520258 456464 520494
rect 456144 513494 456464 520258
rect 456144 513258 456186 513494
rect 456422 513258 456464 513494
rect 456144 506494 456464 513258
rect 456144 506258 456186 506494
rect 456422 506258 456464 506494
rect 456144 499494 456464 506258
rect 456144 499258 456186 499494
rect 456422 499258 456464 499494
rect 456144 492494 456464 499258
rect 456144 492258 456186 492494
rect 456422 492258 456464 492494
rect 456144 485494 456464 492258
rect 456144 485258 456186 485494
rect 456422 485258 456464 485494
rect 456144 478494 456464 485258
rect 456144 478258 456186 478494
rect 456422 478258 456464 478494
rect 456144 471494 456464 478258
rect 456144 471258 456186 471494
rect 456422 471258 456464 471494
rect 456144 464494 456464 471258
rect 456144 464258 456186 464494
rect 456422 464258 456464 464494
rect 456144 457494 456464 464258
rect 456144 457258 456186 457494
rect 456422 457258 456464 457494
rect 456144 450494 456464 457258
rect 456144 450258 456186 450494
rect 456422 450258 456464 450494
rect 456144 443494 456464 450258
rect 456144 443258 456186 443494
rect 456422 443258 456464 443494
rect 456144 436494 456464 443258
rect 456144 436258 456186 436494
rect 456422 436258 456464 436494
rect 456144 429494 456464 436258
rect 456144 429258 456186 429494
rect 456422 429258 456464 429494
rect 456144 422494 456464 429258
rect 456144 422258 456186 422494
rect 456422 422258 456464 422494
rect 456144 415494 456464 422258
rect 456144 415258 456186 415494
rect 456422 415258 456464 415494
rect 456144 408494 456464 415258
rect 456144 408258 456186 408494
rect 456422 408258 456464 408494
rect 456144 401494 456464 408258
rect 456144 401258 456186 401494
rect 456422 401258 456464 401494
rect 456144 394494 456464 401258
rect 456144 394258 456186 394494
rect 456422 394258 456464 394494
rect 456144 387494 456464 394258
rect 456144 387258 456186 387494
rect 456422 387258 456464 387494
rect 456144 380494 456464 387258
rect 456144 380258 456186 380494
rect 456422 380258 456464 380494
rect 456144 373494 456464 380258
rect 456144 373258 456186 373494
rect 456422 373258 456464 373494
rect 456144 366494 456464 373258
rect 456144 366258 456186 366494
rect 456422 366258 456464 366494
rect 456144 359494 456464 366258
rect 456144 359258 456186 359494
rect 456422 359258 456464 359494
rect 456144 352494 456464 359258
rect 456144 352258 456186 352494
rect 456422 352258 456464 352494
rect 456144 345494 456464 352258
rect 456144 345258 456186 345494
rect 456422 345258 456464 345494
rect 456144 338494 456464 345258
rect 456144 338258 456186 338494
rect 456422 338258 456464 338494
rect 456144 331494 456464 338258
rect 456144 331258 456186 331494
rect 456422 331258 456464 331494
rect 456144 324494 456464 331258
rect 456144 324258 456186 324494
rect 456422 324258 456464 324494
rect 456144 317494 456464 324258
rect 456144 317258 456186 317494
rect 456422 317258 456464 317494
rect 456144 310494 456464 317258
rect 456144 310258 456186 310494
rect 456422 310258 456464 310494
rect 456144 303494 456464 310258
rect 456144 303258 456186 303494
rect 456422 303258 456464 303494
rect 456144 296494 456464 303258
rect 456144 296258 456186 296494
rect 456422 296258 456464 296494
rect 456144 289494 456464 296258
rect 456144 289258 456186 289494
rect 456422 289258 456464 289494
rect 456144 282494 456464 289258
rect 456144 282258 456186 282494
rect 456422 282258 456464 282494
rect 456144 275494 456464 282258
rect 456144 275258 456186 275494
rect 456422 275258 456464 275494
rect 456144 268494 456464 275258
rect 456144 268258 456186 268494
rect 456422 268258 456464 268494
rect 456144 261494 456464 268258
rect 456144 261258 456186 261494
rect 456422 261258 456464 261494
rect 456144 254494 456464 261258
rect 456144 254258 456186 254494
rect 456422 254258 456464 254494
rect 456144 247494 456464 254258
rect 456144 247258 456186 247494
rect 456422 247258 456464 247494
rect 456144 240494 456464 247258
rect 456144 240258 456186 240494
rect 456422 240258 456464 240494
rect 456144 233494 456464 240258
rect 456144 233258 456186 233494
rect 456422 233258 456464 233494
rect 456144 226494 456464 233258
rect 456144 226258 456186 226494
rect 456422 226258 456464 226494
rect 456144 219494 456464 226258
rect 456144 219258 456186 219494
rect 456422 219258 456464 219494
rect 456144 212494 456464 219258
rect 456144 212258 456186 212494
rect 456422 212258 456464 212494
rect 456144 205494 456464 212258
rect 456144 205258 456186 205494
rect 456422 205258 456464 205494
rect 456144 198494 456464 205258
rect 456144 198258 456186 198494
rect 456422 198258 456464 198494
rect 456144 191494 456464 198258
rect 456144 191258 456186 191494
rect 456422 191258 456464 191494
rect 456144 184494 456464 191258
rect 456144 184258 456186 184494
rect 456422 184258 456464 184494
rect 456144 177494 456464 184258
rect 456144 177258 456186 177494
rect 456422 177258 456464 177494
rect 456144 170494 456464 177258
rect 456144 170258 456186 170494
rect 456422 170258 456464 170494
rect 456144 163494 456464 170258
rect 456144 163258 456186 163494
rect 456422 163258 456464 163494
rect 456144 156494 456464 163258
rect 456144 156258 456186 156494
rect 456422 156258 456464 156494
rect 456144 149494 456464 156258
rect 456144 149258 456186 149494
rect 456422 149258 456464 149494
rect 456144 142494 456464 149258
rect 456144 142258 456186 142494
rect 456422 142258 456464 142494
rect 456144 135494 456464 142258
rect 456144 135258 456186 135494
rect 456422 135258 456464 135494
rect 456144 128494 456464 135258
rect 456144 128258 456186 128494
rect 456422 128258 456464 128494
rect 456144 121494 456464 128258
rect 456144 121258 456186 121494
rect 456422 121258 456464 121494
rect 456144 114494 456464 121258
rect 456144 114258 456186 114494
rect 456422 114258 456464 114494
rect 456144 107494 456464 114258
rect 456144 107258 456186 107494
rect 456422 107258 456464 107494
rect 456144 100494 456464 107258
rect 456144 100258 456186 100494
rect 456422 100258 456464 100494
rect 456144 93494 456464 100258
rect 456144 93258 456186 93494
rect 456422 93258 456464 93494
rect 456144 86494 456464 93258
rect 456144 86258 456186 86494
rect 456422 86258 456464 86494
rect 456144 79494 456464 86258
rect 456144 79258 456186 79494
rect 456422 79258 456464 79494
rect 456144 72494 456464 79258
rect 456144 72258 456186 72494
rect 456422 72258 456464 72494
rect 456144 65494 456464 72258
rect 456144 65258 456186 65494
rect 456422 65258 456464 65494
rect 456144 58494 456464 65258
rect 456144 58258 456186 58494
rect 456422 58258 456464 58494
rect 456144 51494 456464 58258
rect 456144 51258 456186 51494
rect 456422 51258 456464 51494
rect 456144 44494 456464 51258
rect 456144 44258 456186 44494
rect 456422 44258 456464 44494
rect 456144 37494 456464 44258
rect 456144 37258 456186 37494
rect 456422 37258 456464 37494
rect 456144 30494 456464 37258
rect 456144 30258 456186 30494
rect 456422 30258 456464 30494
rect 456144 23494 456464 30258
rect 456144 23258 456186 23494
rect 456422 23258 456464 23494
rect 456144 16494 456464 23258
rect 456144 16258 456186 16494
rect 456422 16258 456464 16494
rect 456144 9494 456464 16258
rect 456144 9258 456186 9494
rect 456422 9258 456464 9494
rect 456144 2494 456464 9258
rect 456144 2258 456186 2494
rect 456422 2258 456464 2494
rect 456144 -746 456464 2258
rect 456144 -982 456186 -746
rect 456422 -982 456464 -746
rect 456144 -1066 456464 -982
rect 456144 -1302 456186 -1066
rect 456422 -1302 456464 -1066
rect 456144 -2294 456464 -1302
rect 457876 706198 458196 706230
rect 457876 705962 457918 706198
rect 458154 705962 458196 706198
rect 457876 705878 458196 705962
rect 457876 705642 457918 705878
rect 458154 705642 458196 705878
rect 457876 696561 458196 705642
rect 457876 696325 457918 696561
rect 458154 696325 458196 696561
rect 457876 689561 458196 696325
rect 457876 689325 457918 689561
rect 458154 689325 458196 689561
rect 457876 682561 458196 689325
rect 457876 682325 457918 682561
rect 458154 682325 458196 682561
rect 457876 675561 458196 682325
rect 457876 675325 457918 675561
rect 458154 675325 458196 675561
rect 457876 668561 458196 675325
rect 457876 668325 457918 668561
rect 458154 668325 458196 668561
rect 457876 661561 458196 668325
rect 457876 661325 457918 661561
rect 458154 661325 458196 661561
rect 457876 654561 458196 661325
rect 457876 654325 457918 654561
rect 458154 654325 458196 654561
rect 457876 647561 458196 654325
rect 457876 647325 457918 647561
rect 458154 647325 458196 647561
rect 457876 640561 458196 647325
rect 457876 640325 457918 640561
rect 458154 640325 458196 640561
rect 457876 633561 458196 640325
rect 457876 633325 457918 633561
rect 458154 633325 458196 633561
rect 457876 626561 458196 633325
rect 457876 626325 457918 626561
rect 458154 626325 458196 626561
rect 457876 619561 458196 626325
rect 457876 619325 457918 619561
rect 458154 619325 458196 619561
rect 457876 612561 458196 619325
rect 457876 612325 457918 612561
rect 458154 612325 458196 612561
rect 457876 605561 458196 612325
rect 457876 605325 457918 605561
rect 458154 605325 458196 605561
rect 457876 598561 458196 605325
rect 457876 598325 457918 598561
rect 458154 598325 458196 598561
rect 457876 591561 458196 598325
rect 457876 591325 457918 591561
rect 458154 591325 458196 591561
rect 457876 584561 458196 591325
rect 457876 584325 457918 584561
rect 458154 584325 458196 584561
rect 457876 577561 458196 584325
rect 457876 577325 457918 577561
rect 458154 577325 458196 577561
rect 457876 570561 458196 577325
rect 457876 570325 457918 570561
rect 458154 570325 458196 570561
rect 457876 563561 458196 570325
rect 457876 563325 457918 563561
rect 458154 563325 458196 563561
rect 457876 556561 458196 563325
rect 457876 556325 457918 556561
rect 458154 556325 458196 556561
rect 457876 549561 458196 556325
rect 457876 549325 457918 549561
rect 458154 549325 458196 549561
rect 457876 542561 458196 549325
rect 457876 542325 457918 542561
rect 458154 542325 458196 542561
rect 457876 535561 458196 542325
rect 457876 535325 457918 535561
rect 458154 535325 458196 535561
rect 457876 528561 458196 535325
rect 457876 528325 457918 528561
rect 458154 528325 458196 528561
rect 457876 521561 458196 528325
rect 457876 521325 457918 521561
rect 458154 521325 458196 521561
rect 457876 514561 458196 521325
rect 457876 514325 457918 514561
rect 458154 514325 458196 514561
rect 457876 507561 458196 514325
rect 457876 507325 457918 507561
rect 458154 507325 458196 507561
rect 457876 500561 458196 507325
rect 457876 500325 457918 500561
rect 458154 500325 458196 500561
rect 457876 493561 458196 500325
rect 457876 493325 457918 493561
rect 458154 493325 458196 493561
rect 457876 486561 458196 493325
rect 457876 486325 457918 486561
rect 458154 486325 458196 486561
rect 457876 479561 458196 486325
rect 457876 479325 457918 479561
rect 458154 479325 458196 479561
rect 457876 472561 458196 479325
rect 457876 472325 457918 472561
rect 458154 472325 458196 472561
rect 457876 465561 458196 472325
rect 457876 465325 457918 465561
rect 458154 465325 458196 465561
rect 457876 458561 458196 465325
rect 457876 458325 457918 458561
rect 458154 458325 458196 458561
rect 457876 451561 458196 458325
rect 457876 451325 457918 451561
rect 458154 451325 458196 451561
rect 457876 444561 458196 451325
rect 457876 444325 457918 444561
rect 458154 444325 458196 444561
rect 457876 437561 458196 444325
rect 457876 437325 457918 437561
rect 458154 437325 458196 437561
rect 457876 430561 458196 437325
rect 457876 430325 457918 430561
rect 458154 430325 458196 430561
rect 457876 423561 458196 430325
rect 457876 423325 457918 423561
rect 458154 423325 458196 423561
rect 457876 416561 458196 423325
rect 457876 416325 457918 416561
rect 458154 416325 458196 416561
rect 457876 409561 458196 416325
rect 457876 409325 457918 409561
rect 458154 409325 458196 409561
rect 457876 402561 458196 409325
rect 457876 402325 457918 402561
rect 458154 402325 458196 402561
rect 457876 395561 458196 402325
rect 457876 395325 457918 395561
rect 458154 395325 458196 395561
rect 457876 388561 458196 395325
rect 457876 388325 457918 388561
rect 458154 388325 458196 388561
rect 457876 381561 458196 388325
rect 457876 381325 457918 381561
rect 458154 381325 458196 381561
rect 457876 374561 458196 381325
rect 457876 374325 457918 374561
rect 458154 374325 458196 374561
rect 457876 367561 458196 374325
rect 457876 367325 457918 367561
rect 458154 367325 458196 367561
rect 457876 360561 458196 367325
rect 457876 360325 457918 360561
rect 458154 360325 458196 360561
rect 457876 353561 458196 360325
rect 457876 353325 457918 353561
rect 458154 353325 458196 353561
rect 457876 346561 458196 353325
rect 457876 346325 457918 346561
rect 458154 346325 458196 346561
rect 457876 339561 458196 346325
rect 457876 339325 457918 339561
rect 458154 339325 458196 339561
rect 457876 332561 458196 339325
rect 457876 332325 457918 332561
rect 458154 332325 458196 332561
rect 457876 325561 458196 332325
rect 457876 325325 457918 325561
rect 458154 325325 458196 325561
rect 457876 318561 458196 325325
rect 457876 318325 457918 318561
rect 458154 318325 458196 318561
rect 457876 311561 458196 318325
rect 457876 311325 457918 311561
rect 458154 311325 458196 311561
rect 457876 304561 458196 311325
rect 457876 304325 457918 304561
rect 458154 304325 458196 304561
rect 457876 297561 458196 304325
rect 457876 297325 457918 297561
rect 458154 297325 458196 297561
rect 457876 290561 458196 297325
rect 457876 290325 457918 290561
rect 458154 290325 458196 290561
rect 457876 283561 458196 290325
rect 457876 283325 457918 283561
rect 458154 283325 458196 283561
rect 457876 276561 458196 283325
rect 457876 276325 457918 276561
rect 458154 276325 458196 276561
rect 457876 269561 458196 276325
rect 457876 269325 457918 269561
rect 458154 269325 458196 269561
rect 457876 262561 458196 269325
rect 457876 262325 457918 262561
rect 458154 262325 458196 262561
rect 457876 255561 458196 262325
rect 457876 255325 457918 255561
rect 458154 255325 458196 255561
rect 457876 248561 458196 255325
rect 457876 248325 457918 248561
rect 458154 248325 458196 248561
rect 457876 241561 458196 248325
rect 457876 241325 457918 241561
rect 458154 241325 458196 241561
rect 457876 234561 458196 241325
rect 457876 234325 457918 234561
rect 458154 234325 458196 234561
rect 457876 227561 458196 234325
rect 457876 227325 457918 227561
rect 458154 227325 458196 227561
rect 457876 220561 458196 227325
rect 457876 220325 457918 220561
rect 458154 220325 458196 220561
rect 457876 213561 458196 220325
rect 457876 213325 457918 213561
rect 458154 213325 458196 213561
rect 457876 206561 458196 213325
rect 457876 206325 457918 206561
rect 458154 206325 458196 206561
rect 457876 199561 458196 206325
rect 457876 199325 457918 199561
rect 458154 199325 458196 199561
rect 457876 192561 458196 199325
rect 457876 192325 457918 192561
rect 458154 192325 458196 192561
rect 457876 185561 458196 192325
rect 457876 185325 457918 185561
rect 458154 185325 458196 185561
rect 457876 178561 458196 185325
rect 457876 178325 457918 178561
rect 458154 178325 458196 178561
rect 457876 171561 458196 178325
rect 457876 171325 457918 171561
rect 458154 171325 458196 171561
rect 457876 164561 458196 171325
rect 457876 164325 457918 164561
rect 458154 164325 458196 164561
rect 457876 157561 458196 164325
rect 457876 157325 457918 157561
rect 458154 157325 458196 157561
rect 457876 150561 458196 157325
rect 457876 150325 457918 150561
rect 458154 150325 458196 150561
rect 457876 143561 458196 150325
rect 457876 143325 457918 143561
rect 458154 143325 458196 143561
rect 457876 136561 458196 143325
rect 457876 136325 457918 136561
rect 458154 136325 458196 136561
rect 457876 129561 458196 136325
rect 457876 129325 457918 129561
rect 458154 129325 458196 129561
rect 457876 122561 458196 129325
rect 457876 122325 457918 122561
rect 458154 122325 458196 122561
rect 457876 115561 458196 122325
rect 457876 115325 457918 115561
rect 458154 115325 458196 115561
rect 457876 108561 458196 115325
rect 457876 108325 457918 108561
rect 458154 108325 458196 108561
rect 457876 101561 458196 108325
rect 457876 101325 457918 101561
rect 458154 101325 458196 101561
rect 457876 94561 458196 101325
rect 457876 94325 457918 94561
rect 458154 94325 458196 94561
rect 457876 87561 458196 94325
rect 457876 87325 457918 87561
rect 458154 87325 458196 87561
rect 457876 80561 458196 87325
rect 457876 80325 457918 80561
rect 458154 80325 458196 80561
rect 457876 73561 458196 80325
rect 457876 73325 457918 73561
rect 458154 73325 458196 73561
rect 457876 66561 458196 73325
rect 457876 66325 457918 66561
rect 458154 66325 458196 66561
rect 457876 59561 458196 66325
rect 457876 59325 457918 59561
rect 458154 59325 458196 59561
rect 457876 52561 458196 59325
rect 457876 52325 457918 52561
rect 458154 52325 458196 52561
rect 457876 45561 458196 52325
rect 457876 45325 457918 45561
rect 458154 45325 458196 45561
rect 457876 38561 458196 45325
rect 457876 38325 457918 38561
rect 458154 38325 458196 38561
rect 457876 31561 458196 38325
rect 457876 31325 457918 31561
rect 458154 31325 458196 31561
rect 457876 24561 458196 31325
rect 457876 24325 457918 24561
rect 458154 24325 458196 24561
rect 457876 17561 458196 24325
rect 457876 17325 457918 17561
rect 458154 17325 458196 17561
rect 457876 10561 458196 17325
rect 457876 10325 457918 10561
rect 458154 10325 458196 10561
rect 457876 3561 458196 10325
rect 457876 3325 457918 3561
rect 458154 3325 458196 3561
rect 457876 -1706 458196 3325
rect 457876 -1942 457918 -1706
rect 458154 -1942 458196 -1706
rect 457876 -2026 458196 -1942
rect 457876 -2262 457918 -2026
rect 458154 -2262 458196 -2026
rect 457876 -2294 458196 -2262
rect 463144 705238 463464 706230
rect 463144 705002 463186 705238
rect 463422 705002 463464 705238
rect 463144 704918 463464 705002
rect 463144 704682 463186 704918
rect 463422 704682 463464 704918
rect 463144 695494 463464 704682
rect 463144 695258 463186 695494
rect 463422 695258 463464 695494
rect 463144 688494 463464 695258
rect 463144 688258 463186 688494
rect 463422 688258 463464 688494
rect 463144 681494 463464 688258
rect 463144 681258 463186 681494
rect 463422 681258 463464 681494
rect 463144 674494 463464 681258
rect 463144 674258 463186 674494
rect 463422 674258 463464 674494
rect 463144 667494 463464 674258
rect 463144 667258 463186 667494
rect 463422 667258 463464 667494
rect 463144 660494 463464 667258
rect 463144 660258 463186 660494
rect 463422 660258 463464 660494
rect 463144 653494 463464 660258
rect 463144 653258 463186 653494
rect 463422 653258 463464 653494
rect 463144 646494 463464 653258
rect 463144 646258 463186 646494
rect 463422 646258 463464 646494
rect 463144 639494 463464 646258
rect 463144 639258 463186 639494
rect 463422 639258 463464 639494
rect 463144 632494 463464 639258
rect 463144 632258 463186 632494
rect 463422 632258 463464 632494
rect 463144 625494 463464 632258
rect 463144 625258 463186 625494
rect 463422 625258 463464 625494
rect 463144 618494 463464 625258
rect 463144 618258 463186 618494
rect 463422 618258 463464 618494
rect 463144 611494 463464 618258
rect 463144 611258 463186 611494
rect 463422 611258 463464 611494
rect 463144 604494 463464 611258
rect 463144 604258 463186 604494
rect 463422 604258 463464 604494
rect 463144 597494 463464 604258
rect 463144 597258 463186 597494
rect 463422 597258 463464 597494
rect 463144 590494 463464 597258
rect 463144 590258 463186 590494
rect 463422 590258 463464 590494
rect 463144 583494 463464 590258
rect 463144 583258 463186 583494
rect 463422 583258 463464 583494
rect 463144 576494 463464 583258
rect 463144 576258 463186 576494
rect 463422 576258 463464 576494
rect 463144 569494 463464 576258
rect 463144 569258 463186 569494
rect 463422 569258 463464 569494
rect 463144 562494 463464 569258
rect 463144 562258 463186 562494
rect 463422 562258 463464 562494
rect 463144 555494 463464 562258
rect 463144 555258 463186 555494
rect 463422 555258 463464 555494
rect 463144 548494 463464 555258
rect 463144 548258 463186 548494
rect 463422 548258 463464 548494
rect 463144 541494 463464 548258
rect 463144 541258 463186 541494
rect 463422 541258 463464 541494
rect 463144 534494 463464 541258
rect 463144 534258 463186 534494
rect 463422 534258 463464 534494
rect 463144 527494 463464 534258
rect 463144 527258 463186 527494
rect 463422 527258 463464 527494
rect 463144 520494 463464 527258
rect 463144 520258 463186 520494
rect 463422 520258 463464 520494
rect 463144 513494 463464 520258
rect 463144 513258 463186 513494
rect 463422 513258 463464 513494
rect 463144 506494 463464 513258
rect 463144 506258 463186 506494
rect 463422 506258 463464 506494
rect 463144 499494 463464 506258
rect 463144 499258 463186 499494
rect 463422 499258 463464 499494
rect 463144 492494 463464 499258
rect 463144 492258 463186 492494
rect 463422 492258 463464 492494
rect 463144 485494 463464 492258
rect 463144 485258 463186 485494
rect 463422 485258 463464 485494
rect 463144 478494 463464 485258
rect 463144 478258 463186 478494
rect 463422 478258 463464 478494
rect 463144 471494 463464 478258
rect 463144 471258 463186 471494
rect 463422 471258 463464 471494
rect 463144 464494 463464 471258
rect 463144 464258 463186 464494
rect 463422 464258 463464 464494
rect 463144 457494 463464 464258
rect 463144 457258 463186 457494
rect 463422 457258 463464 457494
rect 463144 450494 463464 457258
rect 463144 450258 463186 450494
rect 463422 450258 463464 450494
rect 463144 443494 463464 450258
rect 463144 443258 463186 443494
rect 463422 443258 463464 443494
rect 463144 436494 463464 443258
rect 463144 436258 463186 436494
rect 463422 436258 463464 436494
rect 463144 429494 463464 436258
rect 463144 429258 463186 429494
rect 463422 429258 463464 429494
rect 463144 422494 463464 429258
rect 463144 422258 463186 422494
rect 463422 422258 463464 422494
rect 463144 415494 463464 422258
rect 463144 415258 463186 415494
rect 463422 415258 463464 415494
rect 463144 408494 463464 415258
rect 463144 408258 463186 408494
rect 463422 408258 463464 408494
rect 463144 401494 463464 408258
rect 463144 401258 463186 401494
rect 463422 401258 463464 401494
rect 463144 394494 463464 401258
rect 463144 394258 463186 394494
rect 463422 394258 463464 394494
rect 463144 387494 463464 394258
rect 463144 387258 463186 387494
rect 463422 387258 463464 387494
rect 463144 380494 463464 387258
rect 463144 380258 463186 380494
rect 463422 380258 463464 380494
rect 463144 373494 463464 380258
rect 463144 373258 463186 373494
rect 463422 373258 463464 373494
rect 463144 366494 463464 373258
rect 463144 366258 463186 366494
rect 463422 366258 463464 366494
rect 463144 359494 463464 366258
rect 463144 359258 463186 359494
rect 463422 359258 463464 359494
rect 463144 352494 463464 359258
rect 463144 352258 463186 352494
rect 463422 352258 463464 352494
rect 463144 345494 463464 352258
rect 463144 345258 463186 345494
rect 463422 345258 463464 345494
rect 463144 338494 463464 345258
rect 463144 338258 463186 338494
rect 463422 338258 463464 338494
rect 463144 331494 463464 338258
rect 463144 331258 463186 331494
rect 463422 331258 463464 331494
rect 463144 324494 463464 331258
rect 463144 324258 463186 324494
rect 463422 324258 463464 324494
rect 463144 317494 463464 324258
rect 463144 317258 463186 317494
rect 463422 317258 463464 317494
rect 463144 310494 463464 317258
rect 463144 310258 463186 310494
rect 463422 310258 463464 310494
rect 463144 303494 463464 310258
rect 463144 303258 463186 303494
rect 463422 303258 463464 303494
rect 463144 296494 463464 303258
rect 463144 296258 463186 296494
rect 463422 296258 463464 296494
rect 463144 289494 463464 296258
rect 463144 289258 463186 289494
rect 463422 289258 463464 289494
rect 463144 282494 463464 289258
rect 463144 282258 463186 282494
rect 463422 282258 463464 282494
rect 463144 275494 463464 282258
rect 463144 275258 463186 275494
rect 463422 275258 463464 275494
rect 463144 268494 463464 275258
rect 463144 268258 463186 268494
rect 463422 268258 463464 268494
rect 463144 261494 463464 268258
rect 463144 261258 463186 261494
rect 463422 261258 463464 261494
rect 463144 254494 463464 261258
rect 463144 254258 463186 254494
rect 463422 254258 463464 254494
rect 463144 247494 463464 254258
rect 463144 247258 463186 247494
rect 463422 247258 463464 247494
rect 463144 240494 463464 247258
rect 463144 240258 463186 240494
rect 463422 240258 463464 240494
rect 463144 233494 463464 240258
rect 463144 233258 463186 233494
rect 463422 233258 463464 233494
rect 463144 226494 463464 233258
rect 463144 226258 463186 226494
rect 463422 226258 463464 226494
rect 463144 219494 463464 226258
rect 463144 219258 463186 219494
rect 463422 219258 463464 219494
rect 463144 212494 463464 219258
rect 463144 212258 463186 212494
rect 463422 212258 463464 212494
rect 463144 205494 463464 212258
rect 463144 205258 463186 205494
rect 463422 205258 463464 205494
rect 463144 198494 463464 205258
rect 463144 198258 463186 198494
rect 463422 198258 463464 198494
rect 463144 191494 463464 198258
rect 463144 191258 463186 191494
rect 463422 191258 463464 191494
rect 463144 184494 463464 191258
rect 463144 184258 463186 184494
rect 463422 184258 463464 184494
rect 463144 177494 463464 184258
rect 463144 177258 463186 177494
rect 463422 177258 463464 177494
rect 463144 170494 463464 177258
rect 463144 170258 463186 170494
rect 463422 170258 463464 170494
rect 463144 163494 463464 170258
rect 463144 163258 463186 163494
rect 463422 163258 463464 163494
rect 463144 156494 463464 163258
rect 463144 156258 463186 156494
rect 463422 156258 463464 156494
rect 463144 149494 463464 156258
rect 463144 149258 463186 149494
rect 463422 149258 463464 149494
rect 463144 142494 463464 149258
rect 463144 142258 463186 142494
rect 463422 142258 463464 142494
rect 463144 135494 463464 142258
rect 463144 135258 463186 135494
rect 463422 135258 463464 135494
rect 463144 128494 463464 135258
rect 463144 128258 463186 128494
rect 463422 128258 463464 128494
rect 463144 121494 463464 128258
rect 463144 121258 463186 121494
rect 463422 121258 463464 121494
rect 463144 114494 463464 121258
rect 463144 114258 463186 114494
rect 463422 114258 463464 114494
rect 463144 107494 463464 114258
rect 463144 107258 463186 107494
rect 463422 107258 463464 107494
rect 463144 100494 463464 107258
rect 463144 100258 463186 100494
rect 463422 100258 463464 100494
rect 463144 93494 463464 100258
rect 463144 93258 463186 93494
rect 463422 93258 463464 93494
rect 463144 86494 463464 93258
rect 463144 86258 463186 86494
rect 463422 86258 463464 86494
rect 463144 79494 463464 86258
rect 463144 79258 463186 79494
rect 463422 79258 463464 79494
rect 463144 72494 463464 79258
rect 463144 72258 463186 72494
rect 463422 72258 463464 72494
rect 463144 65494 463464 72258
rect 463144 65258 463186 65494
rect 463422 65258 463464 65494
rect 463144 58494 463464 65258
rect 463144 58258 463186 58494
rect 463422 58258 463464 58494
rect 463144 51494 463464 58258
rect 463144 51258 463186 51494
rect 463422 51258 463464 51494
rect 463144 44494 463464 51258
rect 463144 44258 463186 44494
rect 463422 44258 463464 44494
rect 463144 37494 463464 44258
rect 463144 37258 463186 37494
rect 463422 37258 463464 37494
rect 463144 30494 463464 37258
rect 463144 30258 463186 30494
rect 463422 30258 463464 30494
rect 463144 23494 463464 30258
rect 463144 23258 463186 23494
rect 463422 23258 463464 23494
rect 463144 16494 463464 23258
rect 463144 16258 463186 16494
rect 463422 16258 463464 16494
rect 463144 9494 463464 16258
rect 463144 9258 463186 9494
rect 463422 9258 463464 9494
rect 463144 2494 463464 9258
rect 463144 2258 463186 2494
rect 463422 2258 463464 2494
rect 463144 -746 463464 2258
rect 463144 -982 463186 -746
rect 463422 -982 463464 -746
rect 463144 -1066 463464 -982
rect 463144 -1302 463186 -1066
rect 463422 -1302 463464 -1066
rect 463144 -2294 463464 -1302
rect 464876 706198 465196 706230
rect 464876 705962 464918 706198
rect 465154 705962 465196 706198
rect 464876 705878 465196 705962
rect 464876 705642 464918 705878
rect 465154 705642 465196 705878
rect 464876 696561 465196 705642
rect 464876 696325 464918 696561
rect 465154 696325 465196 696561
rect 464876 689561 465196 696325
rect 464876 689325 464918 689561
rect 465154 689325 465196 689561
rect 464876 682561 465196 689325
rect 464876 682325 464918 682561
rect 465154 682325 465196 682561
rect 464876 675561 465196 682325
rect 464876 675325 464918 675561
rect 465154 675325 465196 675561
rect 464876 668561 465196 675325
rect 464876 668325 464918 668561
rect 465154 668325 465196 668561
rect 464876 661561 465196 668325
rect 464876 661325 464918 661561
rect 465154 661325 465196 661561
rect 464876 654561 465196 661325
rect 464876 654325 464918 654561
rect 465154 654325 465196 654561
rect 464876 647561 465196 654325
rect 464876 647325 464918 647561
rect 465154 647325 465196 647561
rect 464876 640561 465196 647325
rect 464876 640325 464918 640561
rect 465154 640325 465196 640561
rect 464876 633561 465196 640325
rect 464876 633325 464918 633561
rect 465154 633325 465196 633561
rect 464876 626561 465196 633325
rect 464876 626325 464918 626561
rect 465154 626325 465196 626561
rect 464876 619561 465196 626325
rect 464876 619325 464918 619561
rect 465154 619325 465196 619561
rect 464876 612561 465196 619325
rect 464876 612325 464918 612561
rect 465154 612325 465196 612561
rect 464876 605561 465196 612325
rect 464876 605325 464918 605561
rect 465154 605325 465196 605561
rect 464876 598561 465196 605325
rect 464876 598325 464918 598561
rect 465154 598325 465196 598561
rect 464876 591561 465196 598325
rect 464876 591325 464918 591561
rect 465154 591325 465196 591561
rect 464876 584561 465196 591325
rect 464876 584325 464918 584561
rect 465154 584325 465196 584561
rect 464876 577561 465196 584325
rect 464876 577325 464918 577561
rect 465154 577325 465196 577561
rect 464876 570561 465196 577325
rect 464876 570325 464918 570561
rect 465154 570325 465196 570561
rect 464876 563561 465196 570325
rect 464876 563325 464918 563561
rect 465154 563325 465196 563561
rect 464876 556561 465196 563325
rect 464876 556325 464918 556561
rect 465154 556325 465196 556561
rect 464876 549561 465196 556325
rect 464876 549325 464918 549561
rect 465154 549325 465196 549561
rect 464876 542561 465196 549325
rect 464876 542325 464918 542561
rect 465154 542325 465196 542561
rect 464876 535561 465196 542325
rect 464876 535325 464918 535561
rect 465154 535325 465196 535561
rect 464876 528561 465196 535325
rect 464876 528325 464918 528561
rect 465154 528325 465196 528561
rect 464876 521561 465196 528325
rect 464876 521325 464918 521561
rect 465154 521325 465196 521561
rect 464876 514561 465196 521325
rect 464876 514325 464918 514561
rect 465154 514325 465196 514561
rect 464876 507561 465196 514325
rect 464876 507325 464918 507561
rect 465154 507325 465196 507561
rect 464876 500561 465196 507325
rect 464876 500325 464918 500561
rect 465154 500325 465196 500561
rect 464876 493561 465196 500325
rect 464876 493325 464918 493561
rect 465154 493325 465196 493561
rect 464876 486561 465196 493325
rect 464876 486325 464918 486561
rect 465154 486325 465196 486561
rect 464876 479561 465196 486325
rect 464876 479325 464918 479561
rect 465154 479325 465196 479561
rect 464876 472561 465196 479325
rect 464876 472325 464918 472561
rect 465154 472325 465196 472561
rect 464876 465561 465196 472325
rect 464876 465325 464918 465561
rect 465154 465325 465196 465561
rect 464876 458561 465196 465325
rect 464876 458325 464918 458561
rect 465154 458325 465196 458561
rect 464876 451561 465196 458325
rect 464876 451325 464918 451561
rect 465154 451325 465196 451561
rect 464876 444561 465196 451325
rect 464876 444325 464918 444561
rect 465154 444325 465196 444561
rect 464876 437561 465196 444325
rect 464876 437325 464918 437561
rect 465154 437325 465196 437561
rect 464876 430561 465196 437325
rect 464876 430325 464918 430561
rect 465154 430325 465196 430561
rect 464876 423561 465196 430325
rect 464876 423325 464918 423561
rect 465154 423325 465196 423561
rect 464876 416561 465196 423325
rect 464876 416325 464918 416561
rect 465154 416325 465196 416561
rect 464876 409561 465196 416325
rect 464876 409325 464918 409561
rect 465154 409325 465196 409561
rect 464876 402561 465196 409325
rect 464876 402325 464918 402561
rect 465154 402325 465196 402561
rect 464876 395561 465196 402325
rect 464876 395325 464918 395561
rect 465154 395325 465196 395561
rect 464876 388561 465196 395325
rect 464876 388325 464918 388561
rect 465154 388325 465196 388561
rect 464876 381561 465196 388325
rect 464876 381325 464918 381561
rect 465154 381325 465196 381561
rect 464876 374561 465196 381325
rect 464876 374325 464918 374561
rect 465154 374325 465196 374561
rect 464876 367561 465196 374325
rect 464876 367325 464918 367561
rect 465154 367325 465196 367561
rect 464876 360561 465196 367325
rect 464876 360325 464918 360561
rect 465154 360325 465196 360561
rect 464876 353561 465196 360325
rect 464876 353325 464918 353561
rect 465154 353325 465196 353561
rect 464876 346561 465196 353325
rect 464876 346325 464918 346561
rect 465154 346325 465196 346561
rect 464876 339561 465196 346325
rect 464876 339325 464918 339561
rect 465154 339325 465196 339561
rect 464876 332561 465196 339325
rect 464876 332325 464918 332561
rect 465154 332325 465196 332561
rect 464876 325561 465196 332325
rect 464876 325325 464918 325561
rect 465154 325325 465196 325561
rect 464876 318561 465196 325325
rect 464876 318325 464918 318561
rect 465154 318325 465196 318561
rect 464876 311561 465196 318325
rect 464876 311325 464918 311561
rect 465154 311325 465196 311561
rect 464876 304561 465196 311325
rect 464876 304325 464918 304561
rect 465154 304325 465196 304561
rect 464876 297561 465196 304325
rect 464876 297325 464918 297561
rect 465154 297325 465196 297561
rect 464876 290561 465196 297325
rect 464876 290325 464918 290561
rect 465154 290325 465196 290561
rect 464876 283561 465196 290325
rect 464876 283325 464918 283561
rect 465154 283325 465196 283561
rect 464876 276561 465196 283325
rect 464876 276325 464918 276561
rect 465154 276325 465196 276561
rect 464876 269561 465196 276325
rect 464876 269325 464918 269561
rect 465154 269325 465196 269561
rect 464876 262561 465196 269325
rect 464876 262325 464918 262561
rect 465154 262325 465196 262561
rect 464876 255561 465196 262325
rect 464876 255325 464918 255561
rect 465154 255325 465196 255561
rect 464876 248561 465196 255325
rect 464876 248325 464918 248561
rect 465154 248325 465196 248561
rect 464876 241561 465196 248325
rect 464876 241325 464918 241561
rect 465154 241325 465196 241561
rect 464876 234561 465196 241325
rect 464876 234325 464918 234561
rect 465154 234325 465196 234561
rect 464876 227561 465196 234325
rect 464876 227325 464918 227561
rect 465154 227325 465196 227561
rect 464876 220561 465196 227325
rect 464876 220325 464918 220561
rect 465154 220325 465196 220561
rect 464876 213561 465196 220325
rect 464876 213325 464918 213561
rect 465154 213325 465196 213561
rect 464876 206561 465196 213325
rect 464876 206325 464918 206561
rect 465154 206325 465196 206561
rect 464876 199561 465196 206325
rect 464876 199325 464918 199561
rect 465154 199325 465196 199561
rect 464876 192561 465196 199325
rect 464876 192325 464918 192561
rect 465154 192325 465196 192561
rect 464876 185561 465196 192325
rect 464876 185325 464918 185561
rect 465154 185325 465196 185561
rect 464876 178561 465196 185325
rect 464876 178325 464918 178561
rect 465154 178325 465196 178561
rect 464876 171561 465196 178325
rect 464876 171325 464918 171561
rect 465154 171325 465196 171561
rect 464876 164561 465196 171325
rect 464876 164325 464918 164561
rect 465154 164325 465196 164561
rect 464876 157561 465196 164325
rect 464876 157325 464918 157561
rect 465154 157325 465196 157561
rect 464876 150561 465196 157325
rect 464876 150325 464918 150561
rect 465154 150325 465196 150561
rect 464876 143561 465196 150325
rect 464876 143325 464918 143561
rect 465154 143325 465196 143561
rect 464876 136561 465196 143325
rect 464876 136325 464918 136561
rect 465154 136325 465196 136561
rect 464876 129561 465196 136325
rect 464876 129325 464918 129561
rect 465154 129325 465196 129561
rect 464876 122561 465196 129325
rect 464876 122325 464918 122561
rect 465154 122325 465196 122561
rect 464876 115561 465196 122325
rect 464876 115325 464918 115561
rect 465154 115325 465196 115561
rect 464876 108561 465196 115325
rect 464876 108325 464918 108561
rect 465154 108325 465196 108561
rect 464876 101561 465196 108325
rect 464876 101325 464918 101561
rect 465154 101325 465196 101561
rect 464876 94561 465196 101325
rect 464876 94325 464918 94561
rect 465154 94325 465196 94561
rect 464876 87561 465196 94325
rect 464876 87325 464918 87561
rect 465154 87325 465196 87561
rect 464876 80561 465196 87325
rect 464876 80325 464918 80561
rect 465154 80325 465196 80561
rect 464876 73561 465196 80325
rect 464876 73325 464918 73561
rect 465154 73325 465196 73561
rect 464876 66561 465196 73325
rect 464876 66325 464918 66561
rect 465154 66325 465196 66561
rect 464876 59561 465196 66325
rect 464876 59325 464918 59561
rect 465154 59325 465196 59561
rect 464876 52561 465196 59325
rect 464876 52325 464918 52561
rect 465154 52325 465196 52561
rect 464876 45561 465196 52325
rect 464876 45325 464918 45561
rect 465154 45325 465196 45561
rect 464876 38561 465196 45325
rect 464876 38325 464918 38561
rect 465154 38325 465196 38561
rect 464876 31561 465196 38325
rect 464876 31325 464918 31561
rect 465154 31325 465196 31561
rect 464876 24561 465196 31325
rect 464876 24325 464918 24561
rect 465154 24325 465196 24561
rect 464876 17561 465196 24325
rect 464876 17325 464918 17561
rect 465154 17325 465196 17561
rect 464876 10561 465196 17325
rect 464876 10325 464918 10561
rect 465154 10325 465196 10561
rect 464876 3561 465196 10325
rect 464876 3325 464918 3561
rect 465154 3325 465196 3561
rect 464876 -1706 465196 3325
rect 464876 -1942 464918 -1706
rect 465154 -1942 465196 -1706
rect 464876 -2026 465196 -1942
rect 464876 -2262 464918 -2026
rect 465154 -2262 465196 -2026
rect 464876 -2294 465196 -2262
rect 470144 705238 470464 706230
rect 470144 705002 470186 705238
rect 470422 705002 470464 705238
rect 470144 704918 470464 705002
rect 470144 704682 470186 704918
rect 470422 704682 470464 704918
rect 470144 695494 470464 704682
rect 470144 695258 470186 695494
rect 470422 695258 470464 695494
rect 470144 688494 470464 695258
rect 470144 688258 470186 688494
rect 470422 688258 470464 688494
rect 470144 681494 470464 688258
rect 470144 681258 470186 681494
rect 470422 681258 470464 681494
rect 470144 674494 470464 681258
rect 470144 674258 470186 674494
rect 470422 674258 470464 674494
rect 470144 667494 470464 674258
rect 470144 667258 470186 667494
rect 470422 667258 470464 667494
rect 470144 660494 470464 667258
rect 470144 660258 470186 660494
rect 470422 660258 470464 660494
rect 470144 653494 470464 660258
rect 470144 653258 470186 653494
rect 470422 653258 470464 653494
rect 470144 646494 470464 653258
rect 470144 646258 470186 646494
rect 470422 646258 470464 646494
rect 470144 639494 470464 646258
rect 470144 639258 470186 639494
rect 470422 639258 470464 639494
rect 470144 632494 470464 639258
rect 470144 632258 470186 632494
rect 470422 632258 470464 632494
rect 470144 625494 470464 632258
rect 470144 625258 470186 625494
rect 470422 625258 470464 625494
rect 470144 618494 470464 625258
rect 470144 618258 470186 618494
rect 470422 618258 470464 618494
rect 470144 611494 470464 618258
rect 470144 611258 470186 611494
rect 470422 611258 470464 611494
rect 470144 604494 470464 611258
rect 470144 604258 470186 604494
rect 470422 604258 470464 604494
rect 470144 597494 470464 604258
rect 470144 597258 470186 597494
rect 470422 597258 470464 597494
rect 470144 590494 470464 597258
rect 470144 590258 470186 590494
rect 470422 590258 470464 590494
rect 470144 583494 470464 590258
rect 470144 583258 470186 583494
rect 470422 583258 470464 583494
rect 470144 576494 470464 583258
rect 470144 576258 470186 576494
rect 470422 576258 470464 576494
rect 470144 569494 470464 576258
rect 470144 569258 470186 569494
rect 470422 569258 470464 569494
rect 470144 562494 470464 569258
rect 470144 562258 470186 562494
rect 470422 562258 470464 562494
rect 470144 555494 470464 562258
rect 470144 555258 470186 555494
rect 470422 555258 470464 555494
rect 470144 548494 470464 555258
rect 470144 548258 470186 548494
rect 470422 548258 470464 548494
rect 470144 541494 470464 548258
rect 470144 541258 470186 541494
rect 470422 541258 470464 541494
rect 470144 534494 470464 541258
rect 470144 534258 470186 534494
rect 470422 534258 470464 534494
rect 470144 527494 470464 534258
rect 470144 527258 470186 527494
rect 470422 527258 470464 527494
rect 470144 520494 470464 527258
rect 470144 520258 470186 520494
rect 470422 520258 470464 520494
rect 470144 513494 470464 520258
rect 470144 513258 470186 513494
rect 470422 513258 470464 513494
rect 470144 506494 470464 513258
rect 470144 506258 470186 506494
rect 470422 506258 470464 506494
rect 470144 499494 470464 506258
rect 470144 499258 470186 499494
rect 470422 499258 470464 499494
rect 470144 492494 470464 499258
rect 470144 492258 470186 492494
rect 470422 492258 470464 492494
rect 470144 485494 470464 492258
rect 470144 485258 470186 485494
rect 470422 485258 470464 485494
rect 470144 478494 470464 485258
rect 470144 478258 470186 478494
rect 470422 478258 470464 478494
rect 470144 471494 470464 478258
rect 470144 471258 470186 471494
rect 470422 471258 470464 471494
rect 470144 464494 470464 471258
rect 470144 464258 470186 464494
rect 470422 464258 470464 464494
rect 470144 457494 470464 464258
rect 470144 457258 470186 457494
rect 470422 457258 470464 457494
rect 470144 450494 470464 457258
rect 470144 450258 470186 450494
rect 470422 450258 470464 450494
rect 470144 443494 470464 450258
rect 470144 443258 470186 443494
rect 470422 443258 470464 443494
rect 470144 436494 470464 443258
rect 470144 436258 470186 436494
rect 470422 436258 470464 436494
rect 470144 429494 470464 436258
rect 470144 429258 470186 429494
rect 470422 429258 470464 429494
rect 470144 422494 470464 429258
rect 470144 422258 470186 422494
rect 470422 422258 470464 422494
rect 470144 415494 470464 422258
rect 470144 415258 470186 415494
rect 470422 415258 470464 415494
rect 470144 408494 470464 415258
rect 470144 408258 470186 408494
rect 470422 408258 470464 408494
rect 470144 401494 470464 408258
rect 470144 401258 470186 401494
rect 470422 401258 470464 401494
rect 470144 394494 470464 401258
rect 470144 394258 470186 394494
rect 470422 394258 470464 394494
rect 470144 387494 470464 394258
rect 470144 387258 470186 387494
rect 470422 387258 470464 387494
rect 470144 380494 470464 387258
rect 470144 380258 470186 380494
rect 470422 380258 470464 380494
rect 470144 373494 470464 380258
rect 470144 373258 470186 373494
rect 470422 373258 470464 373494
rect 470144 366494 470464 373258
rect 470144 366258 470186 366494
rect 470422 366258 470464 366494
rect 470144 359494 470464 366258
rect 470144 359258 470186 359494
rect 470422 359258 470464 359494
rect 470144 352494 470464 359258
rect 470144 352258 470186 352494
rect 470422 352258 470464 352494
rect 470144 345494 470464 352258
rect 470144 345258 470186 345494
rect 470422 345258 470464 345494
rect 470144 338494 470464 345258
rect 470144 338258 470186 338494
rect 470422 338258 470464 338494
rect 470144 331494 470464 338258
rect 470144 331258 470186 331494
rect 470422 331258 470464 331494
rect 470144 324494 470464 331258
rect 470144 324258 470186 324494
rect 470422 324258 470464 324494
rect 470144 317494 470464 324258
rect 470144 317258 470186 317494
rect 470422 317258 470464 317494
rect 470144 310494 470464 317258
rect 470144 310258 470186 310494
rect 470422 310258 470464 310494
rect 470144 303494 470464 310258
rect 470144 303258 470186 303494
rect 470422 303258 470464 303494
rect 470144 296494 470464 303258
rect 470144 296258 470186 296494
rect 470422 296258 470464 296494
rect 470144 289494 470464 296258
rect 470144 289258 470186 289494
rect 470422 289258 470464 289494
rect 470144 282494 470464 289258
rect 470144 282258 470186 282494
rect 470422 282258 470464 282494
rect 470144 275494 470464 282258
rect 470144 275258 470186 275494
rect 470422 275258 470464 275494
rect 470144 268494 470464 275258
rect 470144 268258 470186 268494
rect 470422 268258 470464 268494
rect 470144 261494 470464 268258
rect 470144 261258 470186 261494
rect 470422 261258 470464 261494
rect 470144 254494 470464 261258
rect 470144 254258 470186 254494
rect 470422 254258 470464 254494
rect 470144 247494 470464 254258
rect 470144 247258 470186 247494
rect 470422 247258 470464 247494
rect 470144 240494 470464 247258
rect 470144 240258 470186 240494
rect 470422 240258 470464 240494
rect 470144 233494 470464 240258
rect 470144 233258 470186 233494
rect 470422 233258 470464 233494
rect 470144 226494 470464 233258
rect 470144 226258 470186 226494
rect 470422 226258 470464 226494
rect 470144 219494 470464 226258
rect 470144 219258 470186 219494
rect 470422 219258 470464 219494
rect 470144 212494 470464 219258
rect 470144 212258 470186 212494
rect 470422 212258 470464 212494
rect 470144 205494 470464 212258
rect 470144 205258 470186 205494
rect 470422 205258 470464 205494
rect 470144 198494 470464 205258
rect 470144 198258 470186 198494
rect 470422 198258 470464 198494
rect 470144 191494 470464 198258
rect 470144 191258 470186 191494
rect 470422 191258 470464 191494
rect 470144 184494 470464 191258
rect 470144 184258 470186 184494
rect 470422 184258 470464 184494
rect 470144 177494 470464 184258
rect 470144 177258 470186 177494
rect 470422 177258 470464 177494
rect 470144 170494 470464 177258
rect 470144 170258 470186 170494
rect 470422 170258 470464 170494
rect 470144 163494 470464 170258
rect 470144 163258 470186 163494
rect 470422 163258 470464 163494
rect 470144 156494 470464 163258
rect 470144 156258 470186 156494
rect 470422 156258 470464 156494
rect 470144 149494 470464 156258
rect 470144 149258 470186 149494
rect 470422 149258 470464 149494
rect 470144 142494 470464 149258
rect 470144 142258 470186 142494
rect 470422 142258 470464 142494
rect 470144 135494 470464 142258
rect 470144 135258 470186 135494
rect 470422 135258 470464 135494
rect 470144 128494 470464 135258
rect 470144 128258 470186 128494
rect 470422 128258 470464 128494
rect 470144 121494 470464 128258
rect 470144 121258 470186 121494
rect 470422 121258 470464 121494
rect 470144 114494 470464 121258
rect 470144 114258 470186 114494
rect 470422 114258 470464 114494
rect 470144 107494 470464 114258
rect 470144 107258 470186 107494
rect 470422 107258 470464 107494
rect 470144 100494 470464 107258
rect 470144 100258 470186 100494
rect 470422 100258 470464 100494
rect 470144 93494 470464 100258
rect 470144 93258 470186 93494
rect 470422 93258 470464 93494
rect 470144 86494 470464 93258
rect 470144 86258 470186 86494
rect 470422 86258 470464 86494
rect 470144 79494 470464 86258
rect 470144 79258 470186 79494
rect 470422 79258 470464 79494
rect 470144 72494 470464 79258
rect 470144 72258 470186 72494
rect 470422 72258 470464 72494
rect 470144 65494 470464 72258
rect 470144 65258 470186 65494
rect 470422 65258 470464 65494
rect 470144 58494 470464 65258
rect 470144 58258 470186 58494
rect 470422 58258 470464 58494
rect 470144 51494 470464 58258
rect 470144 51258 470186 51494
rect 470422 51258 470464 51494
rect 470144 44494 470464 51258
rect 470144 44258 470186 44494
rect 470422 44258 470464 44494
rect 470144 37494 470464 44258
rect 470144 37258 470186 37494
rect 470422 37258 470464 37494
rect 470144 30494 470464 37258
rect 470144 30258 470186 30494
rect 470422 30258 470464 30494
rect 470144 23494 470464 30258
rect 470144 23258 470186 23494
rect 470422 23258 470464 23494
rect 470144 16494 470464 23258
rect 470144 16258 470186 16494
rect 470422 16258 470464 16494
rect 470144 9494 470464 16258
rect 470144 9258 470186 9494
rect 470422 9258 470464 9494
rect 470144 2494 470464 9258
rect 470144 2258 470186 2494
rect 470422 2258 470464 2494
rect 470144 -746 470464 2258
rect 470144 -982 470186 -746
rect 470422 -982 470464 -746
rect 470144 -1066 470464 -982
rect 470144 -1302 470186 -1066
rect 470422 -1302 470464 -1066
rect 470144 -2294 470464 -1302
rect 471876 706198 472196 706230
rect 471876 705962 471918 706198
rect 472154 705962 472196 706198
rect 471876 705878 472196 705962
rect 471876 705642 471918 705878
rect 472154 705642 472196 705878
rect 471876 696561 472196 705642
rect 471876 696325 471918 696561
rect 472154 696325 472196 696561
rect 471876 689561 472196 696325
rect 471876 689325 471918 689561
rect 472154 689325 472196 689561
rect 471876 682561 472196 689325
rect 471876 682325 471918 682561
rect 472154 682325 472196 682561
rect 471876 675561 472196 682325
rect 471876 675325 471918 675561
rect 472154 675325 472196 675561
rect 471876 668561 472196 675325
rect 471876 668325 471918 668561
rect 472154 668325 472196 668561
rect 471876 661561 472196 668325
rect 471876 661325 471918 661561
rect 472154 661325 472196 661561
rect 471876 654561 472196 661325
rect 471876 654325 471918 654561
rect 472154 654325 472196 654561
rect 471876 647561 472196 654325
rect 471876 647325 471918 647561
rect 472154 647325 472196 647561
rect 471876 640561 472196 647325
rect 471876 640325 471918 640561
rect 472154 640325 472196 640561
rect 471876 633561 472196 640325
rect 471876 633325 471918 633561
rect 472154 633325 472196 633561
rect 471876 626561 472196 633325
rect 471876 626325 471918 626561
rect 472154 626325 472196 626561
rect 471876 619561 472196 626325
rect 471876 619325 471918 619561
rect 472154 619325 472196 619561
rect 471876 612561 472196 619325
rect 471876 612325 471918 612561
rect 472154 612325 472196 612561
rect 471876 605561 472196 612325
rect 471876 605325 471918 605561
rect 472154 605325 472196 605561
rect 471876 598561 472196 605325
rect 471876 598325 471918 598561
rect 472154 598325 472196 598561
rect 471876 591561 472196 598325
rect 471876 591325 471918 591561
rect 472154 591325 472196 591561
rect 471876 584561 472196 591325
rect 471876 584325 471918 584561
rect 472154 584325 472196 584561
rect 471876 577561 472196 584325
rect 471876 577325 471918 577561
rect 472154 577325 472196 577561
rect 471876 570561 472196 577325
rect 471876 570325 471918 570561
rect 472154 570325 472196 570561
rect 471876 563561 472196 570325
rect 471876 563325 471918 563561
rect 472154 563325 472196 563561
rect 471876 556561 472196 563325
rect 471876 556325 471918 556561
rect 472154 556325 472196 556561
rect 471876 549561 472196 556325
rect 471876 549325 471918 549561
rect 472154 549325 472196 549561
rect 471876 542561 472196 549325
rect 471876 542325 471918 542561
rect 472154 542325 472196 542561
rect 471876 535561 472196 542325
rect 471876 535325 471918 535561
rect 472154 535325 472196 535561
rect 471876 528561 472196 535325
rect 471876 528325 471918 528561
rect 472154 528325 472196 528561
rect 471876 521561 472196 528325
rect 471876 521325 471918 521561
rect 472154 521325 472196 521561
rect 471876 514561 472196 521325
rect 471876 514325 471918 514561
rect 472154 514325 472196 514561
rect 471876 507561 472196 514325
rect 471876 507325 471918 507561
rect 472154 507325 472196 507561
rect 471876 500561 472196 507325
rect 471876 500325 471918 500561
rect 472154 500325 472196 500561
rect 471876 493561 472196 500325
rect 471876 493325 471918 493561
rect 472154 493325 472196 493561
rect 471876 486561 472196 493325
rect 471876 486325 471918 486561
rect 472154 486325 472196 486561
rect 471876 479561 472196 486325
rect 471876 479325 471918 479561
rect 472154 479325 472196 479561
rect 471876 472561 472196 479325
rect 471876 472325 471918 472561
rect 472154 472325 472196 472561
rect 471876 465561 472196 472325
rect 471876 465325 471918 465561
rect 472154 465325 472196 465561
rect 471876 458561 472196 465325
rect 471876 458325 471918 458561
rect 472154 458325 472196 458561
rect 471876 451561 472196 458325
rect 471876 451325 471918 451561
rect 472154 451325 472196 451561
rect 471876 444561 472196 451325
rect 471876 444325 471918 444561
rect 472154 444325 472196 444561
rect 471876 437561 472196 444325
rect 471876 437325 471918 437561
rect 472154 437325 472196 437561
rect 471876 430561 472196 437325
rect 471876 430325 471918 430561
rect 472154 430325 472196 430561
rect 471876 423561 472196 430325
rect 471876 423325 471918 423561
rect 472154 423325 472196 423561
rect 471876 416561 472196 423325
rect 471876 416325 471918 416561
rect 472154 416325 472196 416561
rect 471876 409561 472196 416325
rect 471876 409325 471918 409561
rect 472154 409325 472196 409561
rect 471876 402561 472196 409325
rect 471876 402325 471918 402561
rect 472154 402325 472196 402561
rect 471876 395561 472196 402325
rect 471876 395325 471918 395561
rect 472154 395325 472196 395561
rect 471876 388561 472196 395325
rect 471876 388325 471918 388561
rect 472154 388325 472196 388561
rect 471876 381561 472196 388325
rect 471876 381325 471918 381561
rect 472154 381325 472196 381561
rect 471876 374561 472196 381325
rect 471876 374325 471918 374561
rect 472154 374325 472196 374561
rect 471876 367561 472196 374325
rect 471876 367325 471918 367561
rect 472154 367325 472196 367561
rect 471876 360561 472196 367325
rect 471876 360325 471918 360561
rect 472154 360325 472196 360561
rect 471876 353561 472196 360325
rect 471876 353325 471918 353561
rect 472154 353325 472196 353561
rect 471876 346561 472196 353325
rect 471876 346325 471918 346561
rect 472154 346325 472196 346561
rect 471876 339561 472196 346325
rect 471876 339325 471918 339561
rect 472154 339325 472196 339561
rect 471876 332561 472196 339325
rect 471876 332325 471918 332561
rect 472154 332325 472196 332561
rect 471876 325561 472196 332325
rect 471876 325325 471918 325561
rect 472154 325325 472196 325561
rect 471876 318561 472196 325325
rect 471876 318325 471918 318561
rect 472154 318325 472196 318561
rect 471876 311561 472196 318325
rect 471876 311325 471918 311561
rect 472154 311325 472196 311561
rect 471876 304561 472196 311325
rect 471876 304325 471918 304561
rect 472154 304325 472196 304561
rect 471876 297561 472196 304325
rect 471876 297325 471918 297561
rect 472154 297325 472196 297561
rect 471876 290561 472196 297325
rect 471876 290325 471918 290561
rect 472154 290325 472196 290561
rect 471876 283561 472196 290325
rect 471876 283325 471918 283561
rect 472154 283325 472196 283561
rect 471876 276561 472196 283325
rect 471876 276325 471918 276561
rect 472154 276325 472196 276561
rect 471876 269561 472196 276325
rect 471876 269325 471918 269561
rect 472154 269325 472196 269561
rect 471876 262561 472196 269325
rect 471876 262325 471918 262561
rect 472154 262325 472196 262561
rect 471876 255561 472196 262325
rect 471876 255325 471918 255561
rect 472154 255325 472196 255561
rect 471876 248561 472196 255325
rect 471876 248325 471918 248561
rect 472154 248325 472196 248561
rect 471876 241561 472196 248325
rect 471876 241325 471918 241561
rect 472154 241325 472196 241561
rect 471876 234561 472196 241325
rect 471876 234325 471918 234561
rect 472154 234325 472196 234561
rect 471876 227561 472196 234325
rect 471876 227325 471918 227561
rect 472154 227325 472196 227561
rect 471876 220561 472196 227325
rect 471876 220325 471918 220561
rect 472154 220325 472196 220561
rect 471876 213561 472196 220325
rect 471876 213325 471918 213561
rect 472154 213325 472196 213561
rect 471876 206561 472196 213325
rect 471876 206325 471918 206561
rect 472154 206325 472196 206561
rect 471876 199561 472196 206325
rect 471876 199325 471918 199561
rect 472154 199325 472196 199561
rect 471876 192561 472196 199325
rect 471876 192325 471918 192561
rect 472154 192325 472196 192561
rect 471876 185561 472196 192325
rect 471876 185325 471918 185561
rect 472154 185325 472196 185561
rect 471876 178561 472196 185325
rect 471876 178325 471918 178561
rect 472154 178325 472196 178561
rect 471876 171561 472196 178325
rect 471876 171325 471918 171561
rect 472154 171325 472196 171561
rect 471876 164561 472196 171325
rect 471876 164325 471918 164561
rect 472154 164325 472196 164561
rect 471876 157561 472196 164325
rect 471876 157325 471918 157561
rect 472154 157325 472196 157561
rect 471876 150561 472196 157325
rect 471876 150325 471918 150561
rect 472154 150325 472196 150561
rect 471876 143561 472196 150325
rect 471876 143325 471918 143561
rect 472154 143325 472196 143561
rect 471876 136561 472196 143325
rect 471876 136325 471918 136561
rect 472154 136325 472196 136561
rect 471876 129561 472196 136325
rect 471876 129325 471918 129561
rect 472154 129325 472196 129561
rect 471876 122561 472196 129325
rect 471876 122325 471918 122561
rect 472154 122325 472196 122561
rect 471876 115561 472196 122325
rect 471876 115325 471918 115561
rect 472154 115325 472196 115561
rect 471876 108561 472196 115325
rect 471876 108325 471918 108561
rect 472154 108325 472196 108561
rect 471876 101561 472196 108325
rect 471876 101325 471918 101561
rect 472154 101325 472196 101561
rect 471876 94561 472196 101325
rect 471876 94325 471918 94561
rect 472154 94325 472196 94561
rect 471876 87561 472196 94325
rect 471876 87325 471918 87561
rect 472154 87325 472196 87561
rect 471876 80561 472196 87325
rect 471876 80325 471918 80561
rect 472154 80325 472196 80561
rect 471876 73561 472196 80325
rect 471876 73325 471918 73561
rect 472154 73325 472196 73561
rect 471876 66561 472196 73325
rect 471876 66325 471918 66561
rect 472154 66325 472196 66561
rect 471876 59561 472196 66325
rect 471876 59325 471918 59561
rect 472154 59325 472196 59561
rect 471876 52561 472196 59325
rect 471876 52325 471918 52561
rect 472154 52325 472196 52561
rect 471876 45561 472196 52325
rect 471876 45325 471918 45561
rect 472154 45325 472196 45561
rect 471876 38561 472196 45325
rect 471876 38325 471918 38561
rect 472154 38325 472196 38561
rect 471876 31561 472196 38325
rect 471876 31325 471918 31561
rect 472154 31325 472196 31561
rect 471876 24561 472196 31325
rect 471876 24325 471918 24561
rect 472154 24325 472196 24561
rect 471876 17561 472196 24325
rect 471876 17325 471918 17561
rect 472154 17325 472196 17561
rect 471876 10561 472196 17325
rect 471876 10325 471918 10561
rect 472154 10325 472196 10561
rect 471876 3561 472196 10325
rect 471876 3325 471918 3561
rect 472154 3325 472196 3561
rect 471876 -1706 472196 3325
rect 471876 -1942 471918 -1706
rect 472154 -1942 472196 -1706
rect 471876 -2026 472196 -1942
rect 471876 -2262 471918 -2026
rect 472154 -2262 472196 -2026
rect 471876 -2294 472196 -2262
rect 477144 705238 477464 706230
rect 477144 705002 477186 705238
rect 477422 705002 477464 705238
rect 477144 704918 477464 705002
rect 477144 704682 477186 704918
rect 477422 704682 477464 704918
rect 477144 695494 477464 704682
rect 477144 695258 477186 695494
rect 477422 695258 477464 695494
rect 477144 688494 477464 695258
rect 477144 688258 477186 688494
rect 477422 688258 477464 688494
rect 477144 681494 477464 688258
rect 477144 681258 477186 681494
rect 477422 681258 477464 681494
rect 477144 674494 477464 681258
rect 477144 674258 477186 674494
rect 477422 674258 477464 674494
rect 477144 667494 477464 674258
rect 477144 667258 477186 667494
rect 477422 667258 477464 667494
rect 477144 660494 477464 667258
rect 477144 660258 477186 660494
rect 477422 660258 477464 660494
rect 477144 653494 477464 660258
rect 477144 653258 477186 653494
rect 477422 653258 477464 653494
rect 477144 646494 477464 653258
rect 477144 646258 477186 646494
rect 477422 646258 477464 646494
rect 477144 639494 477464 646258
rect 477144 639258 477186 639494
rect 477422 639258 477464 639494
rect 477144 632494 477464 639258
rect 477144 632258 477186 632494
rect 477422 632258 477464 632494
rect 477144 625494 477464 632258
rect 477144 625258 477186 625494
rect 477422 625258 477464 625494
rect 477144 618494 477464 625258
rect 477144 618258 477186 618494
rect 477422 618258 477464 618494
rect 477144 611494 477464 618258
rect 477144 611258 477186 611494
rect 477422 611258 477464 611494
rect 477144 604494 477464 611258
rect 477144 604258 477186 604494
rect 477422 604258 477464 604494
rect 477144 597494 477464 604258
rect 477144 597258 477186 597494
rect 477422 597258 477464 597494
rect 477144 590494 477464 597258
rect 477144 590258 477186 590494
rect 477422 590258 477464 590494
rect 477144 583494 477464 590258
rect 477144 583258 477186 583494
rect 477422 583258 477464 583494
rect 477144 576494 477464 583258
rect 477144 576258 477186 576494
rect 477422 576258 477464 576494
rect 477144 569494 477464 576258
rect 477144 569258 477186 569494
rect 477422 569258 477464 569494
rect 477144 562494 477464 569258
rect 477144 562258 477186 562494
rect 477422 562258 477464 562494
rect 477144 555494 477464 562258
rect 477144 555258 477186 555494
rect 477422 555258 477464 555494
rect 477144 548494 477464 555258
rect 477144 548258 477186 548494
rect 477422 548258 477464 548494
rect 477144 541494 477464 548258
rect 477144 541258 477186 541494
rect 477422 541258 477464 541494
rect 477144 534494 477464 541258
rect 477144 534258 477186 534494
rect 477422 534258 477464 534494
rect 477144 527494 477464 534258
rect 477144 527258 477186 527494
rect 477422 527258 477464 527494
rect 477144 520494 477464 527258
rect 477144 520258 477186 520494
rect 477422 520258 477464 520494
rect 477144 513494 477464 520258
rect 477144 513258 477186 513494
rect 477422 513258 477464 513494
rect 477144 506494 477464 513258
rect 477144 506258 477186 506494
rect 477422 506258 477464 506494
rect 477144 499494 477464 506258
rect 477144 499258 477186 499494
rect 477422 499258 477464 499494
rect 477144 492494 477464 499258
rect 477144 492258 477186 492494
rect 477422 492258 477464 492494
rect 477144 485494 477464 492258
rect 477144 485258 477186 485494
rect 477422 485258 477464 485494
rect 477144 478494 477464 485258
rect 477144 478258 477186 478494
rect 477422 478258 477464 478494
rect 477144 471494 477464 478258
rect 477144 471258 477186 471494
rect 477422 471258 477464 471494
rect 477144 464494 477464 471258
rect 477144 464258 477186 464494
rect 477422 464258 477464 464494
rect 477144 457494 477464 464258
rect 477144 457258 477186 457494
rect 477422 457258 477464 457494
rect 477144 450494 477464 457258
rect 477144 450258 477186 450494
rect 477422 450258 477464 450494
rect 477144 443494 477464 450258
rect 477144 443258 477186 443494
rect 477422 443258 477464 443494
rect 477144 436494 477464 443258
rect 477144 436258 477186 436494
rect 477422 436258 477464 436494
rect 477144 429494 477464 436258
rect 477144 429258 477186 429494
rect 477422 429258 477464 429494
rect 477144 422494 477464 429258
rect 477144 422258 477186 422494
rect 477422 422258 477464 422494
rect 477144 415494 477464 422258
rect 477144 415258 477186 415494
rect 477422 415258 477464 415494
rect 477144 408494 477464 415258
rect 477144 408258 477186 408494
rect 477422 408258 477464 408494
rect 477144 401494 477464 408258
rect 477144 401258 477186 401494
rect 477422 401258 477464 401494
rect 477144 394494 477464 401258
rect 477144 394258 477186 394494
rect 477422 394258 477464 394494
rect 477144 387494 477464 394258
rect 477144 387258 477186 387494
rect 477422 387258 477464 387494
rect 477144 380494 477464 387258
rect 477144 380258 477186 380494
rect 477422 380258 477464 380494
rect 477144 373494 477464 380258
rect 477144 373258 477186 373494
rect 477422 373258 477464 373494
rect 477144 366494 477464 373258
rect 477144 366258 477186 366494
rect 477422 366258 477464 366494
rect 477144 359494 477464 366258
rect 477144 359258 477186 359494
rect 477422 359258 477464 359494
rect 477144 352494 477464 359258
rect 477144 352258 477186 352494
rect 477422 352258 477464 352494
rect 477144 345494 477464 352258
rect 477144 345258 477186 345494
rect 477422 345258 477464 345494
rect 477144 338494 477464 345258
rect 477144 338258 477186 338494
rect 477422 338258 477464 338494
rect 477144 331494 477464 338258
rect 477144 331258 477186 331494
rect 477422 331258 477464 331494
rect 477144 324494 477464 331258
rect 477144 324258 477186 324494
rect 477422 324258 477464 324494
rect 477144 317494 477464 324258
rect 477144 317258 477186 317494
rect 477422 317258 477464 317494
rect 477144 310494 477464 317258
rect 477144 310258 477186 310494
rect 477422 310258 477464 310494
rect 477144 303494 477464 310258
rect 477144 303258 477186 303494
rect 477422 303258 477464 303494
rect 477144 296494 477464 303258
rect 477144 296258 477186 296494
rect 477422 296258 477464 296494
rect 477144 289494 477464 296258
rect 477144 289258 477186 289494
rect 477422 289258 477464 289494
rect 477144 282494 477464 289258
rect 477144 282258 477186 282494
rect 477422 282258 477464 282494
rect 477144 275494 477464 282258
rect 477144 275258 477186 275494
rect 477422 275258 477464 275494
rect 477144 268494 477464 275258
rect 477144 268258 477186 268494
rect 477422 268258 477464 268494
rect 477144 261494 477464 268258
rect 477144 261258 477186 261494
rect 477422 261258 477464 261494
rect 477144 254494 477464 261258
rect 477144 254258 477186 254494
rect 477422 254258 477464 254494
rect 477144 247494 477464 254258
rect 477144 247258 477186 247494
rect 477422 247258 477464 247494
rect 477144 240494 477464 247258
rect 477144 240258 477186 240494
rect 477422 240258 477464 240494
rect 477144 233494 477464 240258
rect 477144 233258 477186 233494
rect 477422 233258 477464 233494
rect 477144 226494 477464 233258
rect 477144 226258 477186 226494
rect 477422 226258 477464 226494
rect 477144 219494 477464 226258
rect 477144 219258 477186 219494
rect 477422 219258 477464 219494
rect 477144 212494 477464 219258
rect 477144 212258 477186 212494
rect 477422 212258 477464 212494
rect 477144 205494 477464 212258
rect 477144 205258 477186 205494
rect 477422 205258 477464 205494
rect 477144 198494 477464 205258
rect 477144 198258 477186 198494
rect 477422 198258 477464 198494
rect 477144 191494 477464 198258
rect 477144 191258 477186 191494
rect 477422 191258 477464 191494
rect 477144 184494 477464 191258
rect 477144 184258 477186 184494
rect 477422 184258 477464 184494
rect 477144 177494 477464 184258
rect 477144 177258 477186 177494
rect 477422 177258 477464 177494
rect 477144 170494 477464 177258
rect 477144 170258 477186 170494
rect 477422 170258 477464 170494
rect 477144 163494 477464 170258
rect 477144 163258 477186 163494
rect 477422 163258 477464 163494
rect 477144 156494 477464 163258
rect 477144 156258 477186 156494
rect 477422 156258 477464 156494
rect 477144 149494 477464 156258
rect 477144 149258 477186 149494
rect 477422 149258 477464 149494
rect 477144 142494 477464 149258
rect 477144 142258 477186 142494
rect 477422 142258 477464 142494
rect 477144 135494 477464 142258
rect 477144 135258 477186 135494
rect 477422 135258 477464 135494
rect 477144 128494 477464 135258
rect 477144 128258 477186 128494
rect 477422 128258 477464 128494
rect 477144 121494 477464 128258
rect 477144 121258 477186 121494
rect 477422 121258 477464 121494
rect 477144 114494 477464 121258
rect 477144 114258 477186 114494
rect 477422 114258 477464 114494
rect 477144 107494 477464 114258
rect 477144 107258 477186 107494
rect 477422 107258 477464 107494
rect 477144 100494 477464 107258
rect 477144 100258 477186 100494
rect 477422 100258 477464 100494
rect 477144 93494 477464 100258
rect 477144 93258 477186 93494
rect 477422 93258 477464 93494
rect 477144 86494 477464 93258
rect 477144 86258 477186 86494
rect 477422 86258 477464 86494
rect 477144 79494 477464 86258
rect 477144 79258 477186 79494
rect 477422 79258 477464 79494
rect 477144 72494 477464 79258
rect 477144 72258 477186 72494
rect 477422 72258 477464 72494
rect 477144 65494 477464 72258
rect 477144 65258 477186 65494
rect 477422 65258 477464 65494
rect 477144 58494 477464 65258
rect 477144 58258 477186 58494
rect 477422 58258 477464 58494
rect 477144 51494 477464 58258
rect 477144 51258 477186 51494
rect 477422 51258 477464 51494
rect 477144 44494 477464 51258
rect 477144 44258 477186 44494
rect 477422 44258 477464 44494
rect 477144 37494 477464 44258
rect 477144 37258 477186 37494
rect 477422 37258 477464 37494
rect 477144 30494 477464 37258
rect 477144 30258 477186 30494
rect 477422 30258 477464 30494
rect 477144 23494 477464 30258
rect 477144 23258 477186 23494
rect 477422 23258 477464 23494
rect 477144 16494 477464 23258
rect 477144 16258 477186 16494
rect 477422 16258 477464 16494
rect 477144 9494 477464 16258
rect 477144 9258 477186 9494
rect 477422 9258 477464 9494
rect 477144 2494 477464 9258
rect 477144 2258 477186 2494
rect 477422 2258 477464 2494
rect 477144 -746 477464 2258
rect 477144 -982 477186 -746
rect 477422 -982 477464 -746
rect 477144 -1066 477464 -982
rect 477144 -1302 477186 -1066
rect 477422 -1302 477464 -1066
rect 477144 -2294 477464 -1302
rect 478876 706198 479196 706230
rect 478876 705962 478918 706198
rect 479154 705962 479196 706198
rect 478876 705878 479196 705962
rect 478876 705642 478918 705878
rect 479154 705642 479196 705878
rect 478876 696561 479196 705642
rect 478876 696325 478918 696561
rect 479154 696325 479196 696561
rect 478876 689561 479196 696325
rect 478876 689325 478918 689561
rect 479154 689325 479196 689561
rect 478876 682561 479196 689325
rect 478876 682325 478918 682561
rect 479154 682325 479196 682561
rect 478876 675561 479196 682325
rect 478876 675325 478918 675561
rect 479154 675325 479196 675561
rect 478876 668561 479196 675325
rect 478876 668325 478918 668561
rect 479154 668325 479196 668561
rect 478876 661561 479196 668325
rect 478876 661325 478918 661561
rect 479154 661325 479196 661561
rect 478876 654561 479196 661325
rect 478876 654325 478918 654561
rect 479154 654325 479196 654561
rect 478876 647561 479196 654325
rect 478876 647325 478918 647561
rect 479154 647325 479196 647561
rect 478876 640561 479196 647325
rect 478876 640325 478918 640561
rect 479154 640325 479196 640561
rect 478876 633561 479196 640325
rect 478876 633325 478918 633561
rect 479154 633325 479196 633561
rect 478876 626561 479196 633325
rect 478876 626325 478918 626561
rect 479154 626325 479196 626561
rect 478876 619561 479196 626325
rect 478876 619325 478918 619561
rect 479154 619325 479196 619561
rect 478876 612561 479196 619325
rect 478876 612325 478918 612561
rect 479154 612325 479196 612561
rect 478876 605561 479196 612325
rect 478876 605325 478918 605561
rect 479154 605325 479196 605561
rect 478876 598561 479196 605325
rect 478876 598325 478918 598561
rect 479154 598325 479196 598561
rect 478876 591561 479196 598325
rect 478876 591325 478918 591561
rect 479154 591325 479196 591561
rect 478876 584561 479196 591325
rect 478876 584325 478918 584561
rect 479154 584325 479196 584561
rect 478876 577561 479196 584325
rect 478876 577325 478918 577561
rect 479154 577325 479196 577561
rect 478876 570561 479196 577325
rect 478876 570325 478918 570561
rect 479154 570325 479196 570561
rect 478876 563561 479196 570325
rect 478876 563325 478918 563561
rect 479154 563325 479196 563561
rect 478876 556561 479196 563325
rect 478876 556325 478918 556561
rect 479154 556325 479196 556561
rect 478876 549561 479196 556325
rect 478876 549325 478918 549561
rect 479154 549325 479196 549561
rect 478876 542561 479196 549325
rect 478876 542325 478918 542561
rect 479154 542325 479196 542561
rect 478876 535561 479196 542325
rect 478876 535325 478918 535561
rect 479154 535325 479196 535561
rect 478876 528561 479196 535325
rect 478876 528325 478918 528561
rect 479154 528325 479196 528561
rect 478876 521561 479196 528325
rect 478876 521325 478918 521561
rect 479154 521325 479196 521561
rect 478876 514561 479196 521325
rect 478876 514325 478918 514561
rect 479154 514325 479196 514561
rect 478876 507561 479196 514325
rect 478876 507325 478918 507561
rect 479154 507325 479196 507561
rect 478876 500561 479196 507325
rect 478876 500325 478918 500561
rect 479154 500325 479196 500561
rect 478876 493561 479196 500325
rect 478876 493325 478918 493561
rect 479154 493325 479196 493561
rect 478876 486561 479196 493325
rect 478876 486325 478918 486561
rect 479154 486325 479196 486561
rect 478876 479561 479196 486325
rect 478876 479325 478918 479561
rect 479154 479325 479196 479561
rect 478876 472561 479196 479325
rect 478876 472325 478918 472561
rect 479154 472325 479196 472561
rect 478876 465561 479196 472325
rect 478876 465325 478918 465561
rect 479154 465325 479196 465561
rect 478876 458561 479196 465325
rect 478876 458325 478918 458561
rect 479154 458325 479196 458561
rect 478876 451561 479196 458325
rect 478876 451325 478918 451561
rect 479154 451325 479196 451561
rect 478876 444561 479196 451325
rect 478876 444325 478918 444561
rect 479154 444325 479196 444561
rect 478876 437561 479196 444325
rect 478876 437325 478918 437561
rect 479154 437325 479196 437561
rect 478876 430561 479196 437325
rect 478876 430325 478918 430561
rect 479154 430325 479196 430561
rect 478876 423561 479196 430325
rect 478876 423325 478918 423561
rect 479154 423325 479196 423561
rect 478876 416561 479196 423325
rect 478876 416325 478918 416561
rect 479154 416325 479196 416561
rect 478876 409561 479196 416325
rect 478876 409325 478918 409561
rect 479154 409325 479196 409561
rect 478876 402561 479196 409325
rect 478876 402325 478918 402561
rect 479154 402325 479196 402561
rect 478876 395561 479196 402325
rect 478876 395325 478918 395561
rect 479154 395325 479196 395561
rect 478876 388561 479196 395325
rect 478876 388325 478918 388561
rect 479154 388325 479196 388561
rect 478876 381561 479196 388325
rect 478876 381325 478918 381561
rect 479154 381325 479196 381561
rect 478876 374561 479196 381325
rect 478876 374325 478918 374561
rect 479154 374325 479196 374561
rect 478876 367561 479196 374325
rect 478876 367325 478918 367561
rect 479154 367325 479196 367561
rect 478876 360561 479196 367325
rect 478876 360325 478918 360561
rect 479154 360325 479196 360561
rect 478876 353561 479196 360325
rect 478876 353325 478918 353561
rect 479154 353325 479196 353561
rect 478876 346561 479196 353325
rect 478876 346325 478918 346561
rect 479154 346325 479196 346561
rect 478876 339561 479196 346325
rect 478876 339325 478918 339561
rect 479154 339325 479196 339561
rect 478876 332561 479196 339325
rect 478876 332325 478918 332561
rect 479154 332325 479196 332561
rect 478876 325561 479196 332325
rect 478876 325325 478918 325561
rect 479154 325325 479196 325561
rect 478876 318561 479196 325325
rect 478876 318325 478918 318561
rect 479154 318325 479196 318561
rect 478876 311561 479196 318325
rect 478876 311325 478918 311561
rect 479154 311325 479196 311561
rect 478876 304561 479196 311325
rect 478876 304325 478918 304561
rect 479154 304325 479196 304561
rect 478876 297561 479196 304325
rect 478876 297325 478918 297561
rect 479154 297325 479196 297561
rect 478876 290561 479196 297325
rect 478876 290325 478918 290561
rect 479154 290325 479196 290561
rect 478876 283561 479196 290325
rect 478876 283325 478918 283561
rect 479154 283325 479196 283561
rect 478876 276561 479196 283325
rect 478876 276325 478918 276561
rect 479154 276325 479196 276561
rect 478876 269561 479196 276325
rect 478876 269325 478918 269561
rect 479154 269325 479196 269561
rect 478876 262561 479196 269325
rect 478876 262325 478918 262561
rect 479154 262325 479196 262561
rect 478876 255561 479196 262325
rect 478876 255325 478918 255561
rect 479154 255325 479196 255561
rect 478876 248561 479196 255325
rect 478876 248325 478918 248561
rect 479154 248325 479196 248561
rect 478876 241561 479196 248325
rect 478876 241325 478918 241561
rect 479154 241325 479196 241561
rect 478876 234561 479196 241325
rect 478876 234325 478918 234561
rect 479154 234325 479196 234561
rect 478876 227561 479196 234325
rect 478876 227325 478918 227561
rect 479154 227325 479196 227561
rect 478876 220561 479196 227325
rect 478876 220325 478918 220561
rect 479154 220325 479196 220561
rect 478876 213561 479196 220325
rect 478876 213325 478918 213561
rect 479154 213325 479196 213561
rect 478876 206561 479196 213325
rect 478876 206325 478918 206561
rect 479154 206325 479196 206561
rect 478876 199561 479196 206325
rect 478876 199325 478918 199561
rect 479154 199325 479196 199561
rect 478876 192561 479196 199325
rect 478876 192325 478918 192561
rect 479154 192325 479196 192561
rect 478876 185561 479196 192325
rect 478876 185325 478918 185561
rect 479154 185325 479196 185561
rect 478876 178561 479196 185325
rect 478876 178325 478918 178561
rect 479154 178325 479196 178561
rect 478876 171561 479196 178325
rect 478876 171325 478918 171561
rect 479154 171325 479196 171561
rect 478876 164561 479196 171325
rect 478876 164325 478918 164561
rect 479154 164325 479196 164561
rect 478876 157561 479196 164325
rect 478876 157325 478918 157561
rect 479154 157325 479196 157561
rect 478876 150561 479196 157325
rect 478876 150325 478918 150561
rect 479154 150325 479196 150561
rect 478876 143561 479196 150325
rect 478876 143325 478918 143561
rect 479154 143325 479196 143561
rect 478876 136561 479196 143325
rect 478876 136325 478918 136561
rect 479154 136325 479196 136561
rect 478876 129561 479196 136325
rect 478876 129325 478918 129561
rect 479154 129325 479196 129561
rect 478876 122561 479196 129325
rect 478876 122325 478918 122561
rect 479154 122325 479196 122561
rect 478876 115561 479196 122325
rect 478876 115325 478918 115561
rect 479154 115325 479196 115561
rect 478876 108561 479196 115325
rect 478876 108325 478918 108561
rect 479154 108325 479196 108561
rect 478876 101561 479196 108325
rect 478876 101325 478918 101561
rect 479154 101325 479196 101561
rect 478876 94561 479196 101325
rect 478876 94325 478918 94561
rect 479154 94325 479196 94561
rect 478876 87561 479196 94325
rect 478876 87325 478918 87561
rect 479154 87325 479196 87561
rect 478876 80561 479196 87325
rect 478876 80325 478918 80561
rect 479154 80325 479196 80561
rect 478876 73561 479196 80325
rect 478876 73325 478918 73561
rect 479154 73325 479196 73561
rect 478876 66561 479196 73325
rect 478876 66325 478918 66561
rect 479154 66325 479196 66561
rect 478876 59561 479196 66325
rect 478876 59325 478918 59561
rect 479154 59325 479196 59561
rect 478876 52561 479196 59325
rect 478876 52325 478918 52561
rect 479154 52325 479196 52561
rect 478876 45561 479196 52325
rect 478876 45325 478918 45561
rect 479154 45325 479196 45561
rect 478876 38561 479196 45325
rect 478876 38325 478918 38561
rect 479154 38325 479196 38561
rect 478876 31561 479196 38325
rect 478876 31325 478918 31561
rect 479154 31325 479196 31561
rect 478876 24561 479196 31325
rect 478876 24325 478918 24561
rect 479154 24325 479196 24561
rect 478876 17561 479196 24325
rect 478876 17325 478918 17561
rect 479154 17325 479196 17561
rect 478876 10561 479196 17325
rect 478876 10325 478918 10561
rect 479154 10325 479196 10561
rect 478876 3561 479196 10325
rect 478876 3325 478918 3561
rect 479154 3325 479196 3561
rect 478876 -1706 479196 3325
rect 478876 -1942 478918 -1706
rect 479154 -1942 479196 -1706
rect 478876 -2026 479196 -1942
rect 478876 -2262 478918 -2026
rect 479154 -2262 479196 -2026
rect 478876 -2294 479196 -2262
rect 484144 705238 484464 706230
rect 484144 705002 484186 705238
rect 484422 705002 484464 705238
rect 484144 704918 484464 705002
rect 484144 704682 484186 704918
rect 484422 704682 484464 704918
rect 484144 695494 484464 704682
rect 484144 695258 484186 695494
rect 484422 695258 484464 695494
rect 484144 688494 484464 695258
rect 484144 688258 484186 688494
rect 484422 688258 484464 688494
rect 484144 681494 484464 688258
rect 484144 681258 484186 681494
rect 484422 681258 484464 681494
rect 484144 674494 484464 681258
rect 484144 674258 484186 674494
rect 484422 674258 484464 674494
rect 484144 667494 484464 674258
rect 484144 667258 484186 667494
rect 484422 667258 484464 667494
rect 484144 660494 484464 667258
rect 484144 660258 484186 660494
rect 484422 660258 484464 660494
rect 484144 653494 484464 660258
rect 484144 653258 484186 653494
rect 484422 653258 484464 653494
rect 484144 646494 484464 653258
rect 484144 646258 484186 646494
rect 484422 646258 484464 646494
rect 484144 639494 484464 646258
rect 484144 639258 484186 639494
rect 484422 639258 484464 639494
rect 484144 632494 484464 639258
rect 484144 632258 484186 632494
rect 484422 632258 484464 632494
rect 484144 625494 484464 632258
rect 484144 625258 484186 625494
rect 484422 625258 484464 625494
rect 484144 618494 484464 625258
rect 484144 618258 484186 618494
rect 484422 618258 484464 618494
rect 484144 611494 484464 618258
rect 484144 611258 484186 611494
rect 484422 611258 484464 611494
rect 484144 604494 484464 611258
rect 484144 604258 484186 604494
rect 484422 604258 484464 604494
rect 484144 597494 484464 604258
rect 484144 597258 484186 597494
rect 484422 597258 484464 597494
rect 484144 590494 484464 597258
rect 484144 590258 484186 590494
rect 484422 590258 484464 590494
rect 484144 583494 484464 590258
rect 484144 583258 484186 583494
rect 484422 583258 484464 583494
rect 484144 576494 484464 583258
rect 484144 576258 484186 576494
rect 484422 576258 484464 576494
rect 484144 569494 484464 576258
rect 484144 569258 484186 569494
rect 484422 569258 484464 569494
rect 484144 562494 484464 569258
rect 484144 562258 484186 562494
rect 484422 562258 484464 562494
rect 484144 555494 484464 562258
rect 484144 555258 484186 555494
rect 484422 555258 484464 555494
rect 484144 548494 484464 555258
rect 484144 548258 484186 548494
rect 484422 548258 484464 548494
rect 484144 541494 484464 548258
rect 484144 541258 484186 541494
rect 484422 541258 484464 541494
rect 484144 534494 484464 541258
rect 484144 534258 484186 534494
rect 484422 534258 484464 534494
rect 484144 527494 484464 534258
rect 484144 527258 484186 527494
rect 484422 527258 484464 527494
rect 484144 520494 484464 527258
rect 484144 520258 484186 520494
rect 484422 520258 484464 520494
rect 484144 513494 484464 520258
rect 484144 513258 484186 513494
rect 484422 513258 484464 513494
rect 484144 506494 484464 513258
rect 484144 506258 484186 506494
rect 484422 506258 484464 506494
rect 484144 499494 484464 506258
rect 484144 499258 484186 499494
rect 484422 499258 484464 499494
rect 484144 492494 484464 499258
rect 484144 492258 484186 492494
rect 484422 492258 484464 492494
rect 484144 485494 484464 492258
rect 484144 485258 484186 485494
rect 484422 485258 484464 485494
rect 484144 478494 484464 485258
rect 484144 478258 484186 478494
rect 484422 478258 484464 478494
rect 484144 471494 484464 478258
rect 484144 471258 484186 471494
rect 484422 471258 484464 471494
rect 484144 464494 484464 471258
rect 484144 464258 484186 464494
rect 484422 464258 484464 464494
rect 484144 457494 484464 464258
rect 484144 457258 484186 457494
rect 484422 457258 484464 457494
rect 484144 450494 484464 457258
rect 484144 450258 484186 450494
rect 484422 450258 484464 450494
rect 484144 443494 484464 450258
rect 484144 443258 484186 443494
rect 484422 443258 484464 443494
rect 484144 436494 484464 443258
rect 484144 436258 484186 436494
rect 484422 436258 484464 436494
rect 484144 429494 484464 436258
rect 484144 429258 484186 429494
rect 484422 429258 484464 429494
rect 484144 422494 484464 429258
rect 484144 422258 484186 422494
rect 484422 422258 484464 422494
rect 484144 415494 484464 422258
rect 484144 415258 484186 415494
rect 484422 415258 484464 415494
rect 484144 408494 484464 415258
rect 484144 408258 484186 408494
rect 484422 408258 484464 408494
rect 484144 401494 484464 408258
rect 484144 401258 484186 401494
rect 484422 401258 484464 401494
rect 484144 394494 484464 401258
rect 484144 394258 484186 394494
rect 484422 394258 484464 394494
rect 484144 387494 484464 394258
rect 484144 387258 484186 387494
rect 484422 387258 484464 387494
rect 484144 380494 484464 387258
rect 484144 380258 484186 380494
rect 484422 380258 484464 380494
rect 484144 373494 484464 380258
rect 484144 373258 484186 373494
rect 484422 373258 484464 373494
rect 484144 366494 484464 373258
rect 484144 366258 484186 366494
rect 484422 366258 484464 366494
rect 484144 359494 484464 366258
rect 484144 359258 484186 359494
rect 484422 359258 484464 359494
rect 484144 352494 484464 359258
rect 484144 352258 484186 352494
rect 484422 352258 484464 352494
rect 484144 345494 484464 352258
rect 484144 345258 484186 345494
rect 484422 345258 484464 345494
rect 484144 338494 484464 345258
rect 484144 338258 484186 338494
rect 484422 338258 484464 338494
rect 484144 331494 484464 338258
rect 484144 331258 484186 331494
rect 484422 331258 484464 331494
rect 484144 324494 484464 331258
rect 484144 324258 484186 324494
rect 484422 324258 484464 324494
rect 484144 317494 484464 324258
rect 484144 317258 484186 317494
rect 484422 317258 484464 317494
rect 484144 310494 484464 317258
rect 484144 310258 484186 310494
rect 484422 310258 484464 310494
rect 484144 303494 484464 310258
rect 484144 303258 484186 303494
rect 484422 303258 484464 303494
rect 484144 296494 484464 303258
rect 484144 296258 484186 296494
rect 484422 296258 484464 296494
rect 484144 289494 484464 296258
rect 484144 289258 484186 289494
rect 484422 289258 484464 289494
rect 484144 282494 484464 289258
rect 484144 282258 484186 282494
rect 484422 282258 484464 282494
rect 484144 275494 484464 282258
rect 484144 275258 484186 275494
rect 484422 275258 484464 275494
rect 484144 268494 484464 275258
rect 484144 268258 484186 268494
rect 484422 268258 484464 268494
rect 484144 261494 484464 268258
rect 484144 261258 484186 261494
rect 484422 261258 484464 261494
rect 484144 254494 484464 261258
rect 484144 254258 484186 254494
rect 484422 254258 484464 254494
rect 484144 247494 484464 254258
rect 484144 247258 484186 247494
rect 484422 247258 484464 247494
rect 484144 240494 484464 247258
rect 484144 240258 484186 240494
rect 484422 240258 484464 240494
rect 484144 233494 484464 240258
rect 484144 233258 484186 233494
rect 484422 233258 484464 233494
rect 484144 226494 484464 233258
rect 484144 226258 484186 226494
rect 484422 226258 484464 226494
rect 484144 219494 484464 226258
rect 484144 219258 484186 219494
rect 484422 219258 484464 219494
rect 484144 212494 484464 219258
rect 484144 212258 484186 212494
rect 484422 212258 484464 212494
rect 484144 205494 484464 212258
rect 484144 205258 484186 205494
rect 484422 205258 484464 205494
rect 484144 198494 484464 205258
rect 484144 198258 484186 198494
rect 484422 198258 484464 198494
rect 484144 191494 484464 198258
rect 484144 191258 484186 191494
rect 484422 191258 484464 191494
rect 484144 184494 484464 191258
rect 484144 184258 484186 184494
rect 484422 184258 484464 184494
rect 484144 177494 484464 184258
rect 484144 177258 484186 177494
rect 484422 177258 484464 177494
rect 484144 170494 484464 177258
rect 484144 170258 484186 170494
rect 484422 170258 484464 170494
rect 484144 163494 484464 170258
rect 484144 163258 484186 163494
rect 484422 163258 484464 163494
rect 484144 156494 484464 163258
rect 484144 156258 484186 156494
rect 484422 156258 484464 156494
rect 484144 149494 484464 156258
rect 484144 149258 484186 149494
rect 484422 149258 484464 149494
rect 484144 142494 484464 149258
rect 484144 142258 484186 142494
rect 484422 142258 484464 142494
rect 484144 135494 484464 142258
rect 484144 135258 484186 135494
rect 484422 135258 484464 135494
rect 484144 128494 484464 135258
rect 484144 128258 484186 128494
rect 484422 128258 484464 128494
rect 484144 121494 484464 128258
rect 484144 121258 484186 121494
rect 484422 121258 484464 121494
rect 484144 114494 484464 121258
rect 484144 114258 484186 114494
rect 484422 114258 484464 114494
rect 484144 107494 484464 114258
rect 484144 107258 484186 107494
rect 484422 107258 484464 107494
rect 484144 100494 484464 107258
rect 484144 100258 484186 100494
rect 484422 100258 484464 100494
rect 484144 93494 484464 100258
rect 484144 93258 484186 93494
rect 484422 93258 484464 93494
rect 484144 86494 484464 93258
rect 484144 86258 484186 86494
rect 484422 86258 484464 86494
rect 484144 79494 484464 86258
rect 484144 79258 484186 79494
rect 484422 79258 484464 79494
rect 484144 72494 484464 79258
rect 484144 72258 484186 72494
rect 484422 72258 484464 72494
rect 484144 65494 484464 72258
rect 484144 65258 484186 65494
rect 484422 65258 484464 65494
rect 484144 58494 484464 65258
rect 484144 58258 484186 58494
rect 484422 58258 484464 58494
rect 484144 51494 484464 58258
rect 484144 51258 484186 51494
rect 484422 51258 484464 51494
rect 484144 44494 484464 51258
rect 484144 44258 484186 44494
rect 484422 44258 484464 44494
rect 484144 37494 484464 44258
rect 484144 37258 484186 37494
rect 484422 37258 484464 37494
rect 484144 30494 484464 37258
rect 484144 30258 484186 30494
rect 484422 30258 484464 30494
rect 484144 23494 484464 30258
rect 484144 23258 484186 23494
rect 484422 23258 484464 23494
rect 484144 16494 484464 23258
rect 484144 16258 484186 16494
rect 484422 16258 484464 16494
rect 484144 9494 484464 16258
rect 484144 9258 484186 9494
rect 484422 9258 484464 9494
rect 484144 2494 484464 9258
rect 484144 2258 484186 2494
rect 484422 2258 484464 2494
rect 484144 -746 484464 2258
rect 484144 -982 484186 -746
rect 484422 -982 484464 -746
rect 484144 -1066 484464 -982
rect 484144 -1302 484186 -1066
rect 484422 -1302 484464 -1066
rect 484144 -2294 484464 -1302
rect 485876 706198 486196 706230
rect 485876 705962 485918 706198
rect 486154 705962 486196 706198
rect 485876 705878 486196 705962
rect 485876 705642 485918 705878
rect 486154 705642 486196 705878
rect 485876 696561 486196 705642
rect 485876 696325 485918 696561
rect 486154 696325 486196 696561
rect 485876 689561 486196 696325
rect 485876 689325 485918 689561
rect 486154 689325 486196 689561
rect 485876 682561 486196 689325
rect 485876 682325 485918 682561
rect 486154 682325 486196 682561
rect 485876 675561 486196 682325
rect 485876 675325 485918 675561
rect 486154 675325 486196 675561
rect 485876 668561 486196 675325
rect 485876 668325 485918 668561
rect 486154 668325 486196 668561
rect 485876 661561 486196 668325
rect 485876 661325 485918 661561
rect 486154 661325 486196 661561
rect 485876 654561 486196 661325
rect 485876 654325 485918 654561
rect 486154 654325 486196 654561
rect 485876 647561 486196 654325
rect 485876 647325 485918 647561
rect 486154 647325 486196 647561
rect 485876 640561 486196 647325
rect 485876 640325 485918 640561
rect 486154 640325 486196 640561
rect 485876 633561 486196 640325
rect 485876 633325 485918 633561
rect 486154 633325 486196 633561
rect 485876 626561 486196 633325
rect 485876 626325 485918 626561
rect 486154 626325 486196 626561
rect 485876 619561 486196 626325
rect 485876 619325 485918 619561
rect 486154 619325 486196 619561
rect 485876 612561 486196 619325
rect 485876 612325 485918 612561
rect 486154 612325 486196 612561
rect 485876 605561 486196 612325
rect 485876 605325 485918 605561
rect 486154 605325 486196 605561
rect 485876 598561 486196 605325
rect 485876 598325 485918 598561
rect 486154 598325 486196 598561
rect 485876 591561 486196 598325
rect 485876 591325 485918 591561
rect 486154 591325 486196 591561
rect 485876 584561 486196 591325
rect 485876 584325 485918 584561
rect 486154 584325 486196 584561
rect 485876 577561 486196 584325
rect 485876 577325 485918 577561
rect 486154 577325 486196 577561
rect 485876 570561 486196 577325
rect 485876 570325 485918 570561
rect 486154 570325 486196 570561
rect 485876 563561 486196 570325
rect 485876 563325 485918 563561
rect 486154 563325 486196 563561
rect 485876 556561 486196 563325
rect 485876 556325 485918 556561
rect 486154 556325 486196 556561
rect 485876 549561 486196 556325
rect 485876 549325 485918 549561
rect 486154 549325 486196 549561
rect 485876 542561 486196 549325
rect 485876 542325 485918 542561
rect 486154 542325 486196 542561
rect 485876 535561 486196 542325
rect 485876 535325 485918 535561
rect 486154 535325 486196 535561
rect 485876 528561 486196 535325
rect 485876 528325 485918 528561
rect 486154 528325 486196 528561
rect 485876 521561 486196 528325
rect 485876 521325 485918 521561
rect 486154 521325 486196 521561
rect 485876 514561 486196 521325
rect 485876 514325 485918 514561
rect 486154 514325 486196 514561
rect 485876 507561 486196 514325
rect 485876 507325 485918 507561
rect 486154 507325 486196 507561
rect 485876 500561 486196 507325
rect 485876 500325 485918 500561
rect 486154 500325 486196 500561
rect 485876 493561 486196 500325
rect 485876 493325 485918 493561
rect 486154 493325 486196 493561
rect 485876 486561 486196 493325
rect 485876 486325 485918 486561
rect 486154 486325 486196 486561
rect 485876 479561 486196 486325
rect 485876 479325 485918 479561
rect 486154 479325 486196 479561
rect 485876 472561 486196 479325
rect 485876 472325 485918 472561
rect 486154 472325 486196 472561
rect 485876 465561 486196 472325
rect 485876 465325 485918 465561
rect 486154 465325 486196 465561
rect 485876 458561 486196 465325
rect 485876 458325 485918 458561
rect 486154 458325 486196 458561
rect 485876 451561 486196 458325
rect 485876 451325 485918 451561
rect 486154 451325 486196 451561
rect 485876 444561 486196 451325
rect 485876 444325 485918 444561
rect 486154 444325 486196 444561
rect 485876 437561 486196 444325
rect 485876 437325 485918 437561
rect 486154 437325 486196 437561
rect 485876 430561 486196 437325
rect 485876 430325 485918 430561
rect 486154 430325 486196 430561
rect 485876 423561 486196 430325
rect 485876 423325 485918 423561
rect 486154 423325 486196 423561
rect 485876 416561 486196 423325
rect 485876 416325 485918 416561
rect 486154 416325 486196 416561
rect 485876 409561 486196 416325
rect 485876 409325 485918 409561
rect 486154 409325 486196 409561
rect 485876 402561 486196 409325
rect 485876 402325 485918 402561
rect 486154 402325 486196 402561
rect 485876 395561 486196 402325
rect 485876 395325 485918 395561
rect 486154 395325 486196 395561
rect 485876 388561 486196 395325
rect 485876 388325 485918 388561
rect 486154 388325 486196 388561
rect 485876 381561 486196 388325
rect 485876 381325 485918 381561
rect 486154 381325 486196 381561
rect 485876 374561 486196 381325
rect 485876 374325 485918 374561
rect 486154 374325 486196 374561
rect 485876 367561 486196 374325
rect 485876 367325 485918 367561
rect 486154 367325 486196 367561
rect 485876 360561 486196 367325
rect 485876 360325 485918 360561
rect 486154 360325 486196 360561
rect 485876 353561 486196 360325
rect 485876 353325 485918 353561
rect 486154 353325 486196 353561
rect 485876 346561 486196 353325
rect 485876 346325 485918 346561
rect 486154 346325 486196 346561
rect 485876 339561 486196 346325
rect 485876 339325 485918 339561
rect 486154 339325 486196 339561
rect 485876 332561 486196 339325
rect 485876 332325 485918 332561
rect 486154 332325 486196 332561
rect 485876 325561 486196 332325
rect 485876 325325 485918 325561
rect 486154 325325 486196 325561
rect 485876 318561 486196 325325
rect 485876 318325 485918 318561
rect 486154 318325 486196 318561
rect 485876 311561 486196 318325
rect 485876 311325 485918 311561
rect 486154 311325 486196 311561
rect 485876 304561 486196 311325
rect 485876 304325 485918 304561
rect 486154 304325 486196 304561
rect 485876 297561 486196 304325
rect 485876 297325 485918 297561
rect 486154 297325 486196 297561
rect 485876 290561 486196 297325
rect 485876 290325 485918 290561
rect 486154 290325 486196 290561
rect 485876 283561 486196 290325
rect 485876 283325 485918 283561
rect 486154 283325 486196 283561
rect 485876 276561 486196 283325
rect 485876 276325 485918 276561
rect 486154 276325 486196 276561
rect 485876 269561 486196 276325
rect 485876 269325 485918 269561
rect 486154 269325 486196 269561
rect 485876 262561 486196 269325
rect 485876 262325 485918 262561
rect 486154 262325 486196 262561
rect 485876 255561 486196 262325
rect 485876 255325 485918 255561
rect 486154 255325 486196 255561
rect 485876 248561 486196 255325
rect 485876 248325 485918 248561
rect 486154 248325 486196 248561
rect 485876 241561 486196 248325
rect 485876 241325 485918 241561
rect 486154 241325 486196 241561
rect 485876 234561 486196 241325
rect 485876 234325 485918 234561
rect 486154 234325 486196 234561
rect 485876 227561 486196 234325
rect 485876 227325 485918 227561
rect 486154 227325 486196 227561
rect 485876 220561 486196 227325
rect 485876 220325 485918 220561
rect 486154 220325 486196 220561
rect 485876 213561 486196 220325
rect 485876 213325 485918 213561
rect 486154 213325 486196 213561
rect 485876 206561 486196 213325
rect 485876 206325 485918 206561
rect 486154 206325 486196 206561
rect 485876 199561 486196 206325
rect 485876 199325 485918 199561
rect 486154 199325 486196 199561
rect 485876 192561 486196 199325
rect 485876 192325 485918 192561
rect 486154 192325 486196 192561
rect 485876 185561 486196 192325
rect 485876 185325 485918 185561
rect 486154 185325 486196 185561
rect 485876 178561 486196 185325
rect 485876 178325 485918 178561
rect 486154 178325 486196 178561
rect 485876 171561 486196 178325
rect 485876 171325 485918 171561
rect 486154 171325 486196 171561
rect 485876 164561 486196 171325
rect 485876 164325 485918 164561
rect 486154 164325 486196 164561
rect 485876 157561 486196 164325
rect 485876 157325 485918 157561
rect 486154 157325 486196 157561
rect 485876 150561 486196 157325
rect 485876 150325 485918 150561
rect 486154 150325 486196 150561
rect 485876 143561 486196 150325
rect 485876 143325 485918 143561
rect 486154 143325 486196 143561
rect 485876 136561 486196 143325
rect 485876 136325 485918 136561
rect 486154 136325 486196 136561
rect 485876 129561 486196 136325
rect 485876 129325 485918 129561
rect 486154 129325 486196 129561
rect 485876 122561 486196 129325
rect 485876 122325 485918 122561
rect 486154 122325 486196 122561
rect 485876 115561 486196 122325
rect 485876 115325 485918 115561
rect 486154 115325 486196 115561
rect 485876 108561 486196 115325
rect 485876 108325 485918 108561
rect 486154 108325 486196 108561
rect 485876 101561 486196 108325
rect 485876 101325 485918 101561
rect 486154 101325 486196 101561
rect 485876 94561 486196 101325
rect 485876 94325 485918 94561
rect 486154 94325 486196 94561
rect 485876 87561 486196 94325
rect 485876 87325 485918 87561
rect 486154 87325 486196 87561
rect 485876 80561 486196 87325
rect 485876 80325 485918 80561
rect 486154 80325 486196 80561
rect 485876 73561 486196 80325
rect 485876 73325 485918 73561
rect 486154 73325 486196 73561
rect 485876 66561 486196 73325
rect 485876 66325 485918 66561
rect 486154 66325 486196 66561
rect 485876 59561 486196 66325
rect 485876 59325 485918 59561
rect 486154 59325 486196 59561
rect 485876 52561 486196 59325
rect 485876 52325 485918 52561
rect 486154 52325 486196 52561
rect 485876 45561 486196 52325
rect 485876 45325 485918 45561
rect 486154 45325 486196 45561
rect 485876 38561 486196 45325
rect 485876 38325 485918 38561
rect 486154 38325 486196 38561
rect 485876 31561 486196 38325
rect 485876 31325 485918 31561
rect 486154 31325 486196 31561
rect 485876 24561 486196 31325
rect 485876 24325 485918 24561
rect 486154 24325 486196 24561
rect 485876 17561 486196 24325
rect 485876 17325 485918 17561
rect 486154 17325 486196 17561
rect 485876 10561 486196 17325
rect 485876 10325 485918 10561
rect 486154 10325 486196 10561
rect 485876 3561 486196 10325
rect 485876 3325 485918 3561
rect 486154 3325 486196 3561
rect 485876 -1706 486196 3325
rect 485876 -1942 485918 -1706
rect 486154 -1942 486196 -1706
rect 485876 -2026 486196 -1942
rect 485876 -2262 485918 -2026
rect 486154 -2262 486196 -2026
rect 485876 -2294 486196 -2262
rect 491144 705238 491464 706230
rect 491144 705002 491186 705238
rect 491422 705002 491464 705238
rect 491144 704918 491464 705002
rect 491144 704682 491186 704918
rect 491422 704682 491464 704918
rect 491144 695494 491464 704682
rect 491144 695258 491186 695494
rect 491422 695258 491464 695494
rect 491144 688494 491464 695258
rect 491144 688258 491186 688494
rect 491422 688258 491464 688494
rect 491144 681494 491464 688258
rect 491144 681258 491186 681494
rect 491422 681258 491464 681494
rect 491144 674494 491464 681258
rect 491144 674258 491186 674494
rect 491422 674258 491464 674494
rect 491144 667494 491464 674258
rect 491144 667258 491186 667494
rect 491422 667258 491464 667494
rect 491144 660494 491464 667258
rect 491144 660258 491186 660494
rect 491422 660258 491464 660494
rect 491144 653494 491464 660258
rect 491144 653258 491186 653494
rect 491422 653258 491464 653494
rect 491144 646494 491464 653258
rect 491144 646258 491186 646494
rect 491422 646258 491464 646494
rect 491144 639494 491464 646258
rect 491144 639258 491186 639494
rect 491422 639258 491464 639494
rect 491144 632494 491464 639258
rect 491144 632258 491186 632494
rect 491422 632258 491464 632494
rect 491144 625494 491464 632258
rect 491144 625258 491186 625494
rect 491422 625258 491464 625494
rect 491144 618494 491464 625258
rect 491144 618258 491186 618494
rect 491422 618258 491464 618494
rect 491144 611494 491464 618258
rect 491144 611258 491186 611494
rect 491422 611258 491464 611494
rect 491144 604494 491464 611258
rect 491144 604258 491186 604494
rect 491422 604258 491464 604494
rect 491144 597494 491464 604258
rect 491144 597258 491186 597494
rect 491422 597258 491464 597494
rect 491144 590494 491464 597258
rect 491144 590258 491186 590494
rect 491422 590258 491464 590494
rect 491144 583494 491464 590258
rect 491144 583258 491186 583494
rect 491422 583258 491464 583494
rect 491144 576494 491464 583258
rect 491144 576258 491186 576494
rect 491422 576258 491464 576494
rect 491144 569494 491464 576258
rect 491144 569258 491186 569494
rect 491422 569258 491464 569494
rect 491144 562494 491464 569258
rect 491144 562258 491186 562494
rect 491422 562258 491464 562494
rect 491144 555494 491464 562258
rect 491144 555258 491186 555494
rect 491422 555258 491464 555494
rect 491144 548494 491464 555258
rect 491144 548258 491186 548494
rect 491422 548258 491464 548494
rect 491144 541494 491464 548258
rect 491144 541258 491186 541494
rect 491422 541258 491464 541494
rect 491144 534494 491464 541258
rect 491144 534258 491186 534494
rect 491422 534258 491464 534494
rect 491144 527494 491464 534258
rect 491144 527258 491186 527494
rect 491422 527258 491464 527494
rect 491144 520494 491464 527258
rect 491144 520258 491186 520494
rect 491422 520258 491464 520494
rect 491144 513494 491464 520258
rect 491144 513258 491186 513494
rect 491422 513258 491464 513494
rect 491144 506494 491464 513258
rect 491144 506258 491186 506494
rect 491422 506258 491464 506494
rect 491144 499494 491464 506258
rect 491144 499258 491186 499494
rect 491422 499258 491464 499494
rect 491144 492494 491464 499258
rect 491144 492258 491186 492494
rect 491422 492258 491464 492494
rect 491144 485494 491464 492258
rect 491144 485258 491186 485494
rect 491422 485258 491464 485494
rect 491144 478494 491464 485258
rect 491144 478258 491186 478494
rect 491422 478258 491464 478494
rect 491144 471494 491464 478258
rect 491144 471258 491186 471494
rect 491422 471258 491464 471494
rect 491144 464494 491464 471258
rect 491144 464258 491186 464494
rect 491422 464258 491464 464494
rect 491144 457494 491464 464258
rect 491144 457258 491186 457494
rect 491422 457258 491464 457494
rect 491144 450494 491464 457258
rect 491144 450258 491186 450494
rect 491422 450258 491464 450494
rect 491144 443494 491464 450258
rect 491144 443258 491186 443494
rect 491422 443258 491464 443494
rect 491144 436494 491464 443258
rect 491144 436258 491186 436494
rect 491422 436258 491464 436494
rect 491144 429494 491464 436258
rect 491144 429258 491186 429494
rect 491422 429258 491464 429494
rect 491144 422494 491464 429258
rect 491144 422258 491186 422494
rect 491422 422258 491464 422494
rect 491144 415494 491464 422258
rect 491144 415258 491186 415494
rect 491422 415258 491464 415494
rect 491144 408494 491464 415258
rect 491144 408258 491186 408494
rect 491422 408258 491464 408494
rect 491144 401494 491464 408258
rect 491144 401258 491186 401494
rect 491422 401258 491464 401494
rect 491144 394494 491464 401258
rect 491144 394258 491186 394494
rect 491422 394258 491464 394494
rect 491144 387494 491464 394258
rect 491144 387258 491186 387494
rect 491422 387258 491464 387494
rect 491144 380494 491464 387258
rect 491144 380258 491186 380494
rect 491422 380258 491464 380494
rect 491144 373494 491464 380258
rect 491144 373258 491186 373494
rect 491422 373258 491464 373494
rect 491144 366494 491464 373258
rect 491144 366258 491186 366494
rect 491422 366258 491464 366494
rect 491144 359494 491464 366258
rect 491144 359258 491186 359494
rect 491422 359258 491464 359494
rect 491144 352494 491464 359258
rect 491144 352258 491186 352494
rect 491422 352258 491464 352494
rect 491144 345494 491464 352258
rect 491144 345258 491186 345494
rect 491422 345258 491464 345494
rect 491144 338494 491464 345258
rect 491144 338258 491186 338494
rect 491422 338258 491464 338494
rect 491144 331494 491464 338258
rect 491144 331258 491186 331494
rect 491422 331258 491464 331494
rect 491144 324494 491464 331258
rect 491144 324258 491186 324494
rect 491422 324258 491464 324494
rect 491144 317494 491464 324258
rect 491144 317258 491186 317494
rect 491422 317258 491464 317494
rect 491144 310494 491464 317258
rect 491144 310258 491186 310494
rect 491422 310258 491464 310494
rect 491144 303494 491464 310258
rect 491144 303258 491186 303494
rect 491422 303258 491464 303494
rect 491144 296494 491464 303258
rect 491144 296258 491186 296494
rect 491422 296258 491464 296494
rect 491144 289494 491464 296258
rect 491144 289258 491186 289494
rect 491422 289258 491464 289494
rect 491144 282494 491464 289258
rect 491144 282258 491186 282494
rect 491422 282258 491464 282494
rect 491144 275494 491464 282258
rect 491144 275258 491186 275494
rect 491422 275258 491464 275494
rect 491144 268494 491464 275258
rect 491144 268258 491186 268494
rect 491422 268258 491464 268494
rect 491144 261494 491464 268258
rect 491144 261258 491186 261494
rect 491422 261258 491464 261494
rect 491144 254494 491464 261258
rect 491144 254258 491186 254494
rect 491422 254258 491464 254494
rect 491144 247494 491464 254258
rect 491144 247258 491186 247494
rect 491422 247258 491464 247494
rect 491144 240494 491464 247258
rect 491144 240258 491186 240494
rect 491422 240258 491464 240494
rect 491144 233494 491464 240258
rect 491144 233258 491186 233494
rect 491422 233258 491464 233494
rect 491144 226494 491464 233258
rect 491144 226258 491186 226494
rect 491422 226258 491464 226494
rect 491144 219494 491464 226258
rect 491144 219258 491186 219494
rect 491422 219258 491464 219494
rect 491144 212494 491464 219258
rect 491144 212258 491186 212494
rect 491422 212258 491464 212494
rect 491144 205494 491464 212258
rect 491144 205258 491186 205494
rect 491422 205258 491464 205494
rect 491144 198494 491464 205258
rect 491144 198258 491186 198494
rect 491422 198258 491464 198494
rect 491144 191494 491464 198258
rect 491144 191258 491186 191494
rect 491422 191258 491464 191494
rect 491144 184494 491464 191258
rect 491144 184258 491186 184494
rect 491422 184258 491464 184494
rect 491144 177494 491464 184258
rect 491144 177258 491186 177494
rect 491422 177258 491464 177494
rect 491144 170494 491464 177258
rect 491144 170258 491186 170494
rect 491422 170258 491464 170494
rect 491144 163494 491464 170258
rect 491144 163258 491186 163494
rect 491422 163258 491464 163494
rect 491144 156494 491464 163258
rect 491144 156258 491186 156494
rect 491422 156258 491464 156494
rect 491144 149494 491464 156258
rect 491144 149258 491186 149494
rect 491422 149258 491464 149494
rect 491144 142494 491464 149258
rect 491144 142258 491186 142494
rect 491422 142258 491464 142494
rect 491144 135494 491464 142258
rect 491144 135258 491186 135494
rect 491422 135258 491464 135494
rect 491144 128494 491464 135258
rect 491144 128258 491186 128494
rect 491422 128258 491464 128494
rect 491144 121494 491464 128258
rect 491144 121258 491186 121494
rect 491422 121258 491464 121494
rect 491144 114494 491464 121258
rect 491144 114258 491186 114494
rect 491422 114258 491464 114494
rect 491144 107494 491464 114258
rect 491144 107258 491186 107494
rect 491422 107258 491464 107494
rect 491144 100494 491464 107258
rect 491144 100258 491186 100494
rect 491422 100258 491464 100494
rect 491144 93494 491464 100258
rect 491144 93258 491186 93494
rect 491422 93258 491464 93494
rect 491144 86494 491464 93258
rect 491144 86258 491186 86494
rect 491422 86258 491464 86494
rect 491144 79494 491464 86258
rect 491144 79258 491186 79494
rect 491422 79258 491464 79494
rect 491144 72494 491464 79258
rect 491144 72258 491186 72494
rect 491422 72258 491464 72494
rect 491144 65494 491464 72258
rect 491144 65258 491186 65494
rect 491422 65258 491464 65494
rect 491144 58494 491464 65258
rect 491144 58258 491186 58494
rect 491422 58258 491464 58494
rect 491144 51494 491464 58258
rect 491144 51258 491186 51494
rect 491422 51258 491464 51494
rect 491144 44494 491464 51258
rect 491144 44258 491186 44494
rect 491422 44258 491464 44494
rect 491144 37494 491464 44258
rect 491144 37258 491186 37494
rect 491422 37258 491464 37494
rect 491144 30494 491464 37258
rect 491144 30258 491186 30494
rect 491422 30258 491464 30494
rect 491144 23494 491464 30258
rect 491144 23258 491186 23494
rect 491422 23258 491464 23494
rect 491144 16494 491464 23258
rect 491144 16258 491186 16494
rect 491422 16258 491464 16494
rect 491144 9494 491464 16258
rect 491144 9258 491186 9494
rect 491422 9258 491464 9494
rect 491144 2494 491464 9258
rect 491144 2258 491186 2494
rect 491422 2258 491464 2494
rect 491144 -746 491464 2258
rect 491144 -982 491186 -746
rect 491422 -982 491464 -746
rect 491144 -1066 491464 -982
rect 491144 -1302 491186 -1066
rect 491422 -1302 491464 -1066
rect 491144 -2294 491464 -1302
rect 492876 706198 493196 706230
rect 492876 705962 492918 706198
rect 493154 705962 493196 706198
rect 492876 705878 493196 705962
rect 492876 705642 492918 705878
rect 493154 705642 493196 705878
rect 492876 696561 493196 705642
rect 492876 696325 492918 696561
rect 493154 696325 493196 696561
rect 492876 689561 493196 696325
rect 492876 689325 492918 689561
rect 493154 689325 493196 689561
rect 492876 682561 493196 689325
rect 492876 682325 492918 682561
rect 493154 682325 493196 682561
rect 492876 675561 493196 682325
rect 492876 675325 492918 675561
rect 493154 675325 493196 675561
rect 492876 668561 493196 675325
rect 492876 668325 492918 668561
rect 493154 668325 493196 668561
rect 492876 661561 493196 668325
rect 492876 661325 492918 661561
rect 493154 661325 493196 661561
rect 492876 654561 493196 661325
rect 492876 654325 492918 654561
rect 493154 654325 493196 654561
rect 492876 647561 493196 654325
rect 492876 647325 492918 647561
rect 493154 647325 493196 647561
rect 492876 640561 493196 647325
rect 492876 640325 492918 640561
rect 493154 640325 493196 640561
rect 492876 633561 493196 640325
rect 492876 633325 492918 633561
rect 493154 633325 493196 633561
rect 492876 626561 493196 633325
rect 492876 626325 492918 626561
rect 493154 626325 493196 626561
rect 492876 619561 493196 626325
rect 492876 619325 492918 619561
rect 493154 619325 493196 619561
rect 492876 612561 493196 619325
rect 492876 612325 492918 612561
rect 493154 612325 493196 612561
rect 492876 605561 493196 612325
rect 492876 605325 492918 605561
rect 493154 605325 493196 605561
rect 492876 598561 493196 605325
rect 492876 598325 492918 598561
rect 493154 598325 493196 598561
rect 492876 591561 493196 598325
rect 492876 591325 492918 591561
rect 493154 591325 493196 591561
rect 492876 584561 493196 591325
rect 492876 584325 492918 584561
rect 493154 584325 493196 584561
rect 492876 577561 493196 584325
rect 492876 577325 492918 577561
rect 493154 577325 493196 577561
rect 492876 570561 493196 577325
rect 492876 570325 492918 570561
rect 493154 570325 493196 570561
rect 492876 563561 493196 570325
rect 492876 563325 492918 563561
rect 493154 563325 493196 563561
rect 492876 556561 493196 563325
rect 492876 556325 492918 556561
rect 493154 556325 493196 556561
rect 492876 549561 493196 556325
rect 492876 549325 492918 549561
rect 493154 549325 493196 549561
rect 492876 542561 493196 549325
rect 492876 542325 492918 542561
rect 493154 542325 493196 542561
rect 492876 535561 493196 542325
rect 492876 535325 492918 535561
rect 493154 535325 493196 535561
rect 492876 528561 493196 535325
rect 492876 528325 492918 528561
rect 493154 528325 493196 528561
rect 492876 521561 493196 528325
rect 492876 521325 492918 521561
rect 493154 521325 493196 521561
rect 492876 514561 493196 521325
rect 492876 514325 492918 514561
rect 493154 514325 493196 514561
rect 492876 507561 493196 514325
rect 492876 507325 492918 507561
rect 493154 507325 493196 507561
rect 492876 500561 493196 507325
rect 492876 500325 492918 500561
rect 493154 500325 493196 500561
rect 492876 493561 493196 500325
rect 492876 493325 492918 493561
rect 493154 493325 493196 493561
rect 492876 486561 493196 493325
rect 492876 486325 492918 486561
rect 493154 486325 493196 486561
rect 492876 479561 493196 486325
rect 492876 479325 492918 479561
rect 493154 479325 493196 479561
rect 492876 472561 493196 479325
rect 492876 472325 492918 472561
rect 493154 472325 493196 472561
rect 492876 465561 493196 472325
rect 492876 465325 492918 465561
rect 493154 465325 493196 465561
rect 492876 458561 493196 465325
rect 492876 458325 492918 458561
rect 493154 458325 493196 458561
rect 492876 451561 493196 458325
rect 492876 451325 492918 451561
rect 493154 451325 493196 451561
rect 492876 444561 493196 451325
rect 492876 444325 492918 444561
rect 493154 444325 493196 444561
rect 492876 437561 493196 444325
rect 492876 437325 492918 437561
rect 493154 437325 493196 437561
rect 492876 430561 493196 437325
rect 492876 430325 492918 430561
rect 493154 430325 493196 430561
rect 492876 423561 493196 430325
rect 492876 423325 492918 423561
rect 493154 423325 493196 423561
rect 492876 416561 493196 423325
rect 492876 416325 492918 416561
rect 493154 416325 493196 416561
rect 492876 409561 493196 416325
rect 492876 409325 492918 409561
rect 493154 409325 493196 409561
rect 492876 402561 493196 409325
rect 492876 402325 492918 402561
rect 493154 402325 493196 402561
rect 492876 395561 493196 402325
rect 492876 395325 492918 395561
rect 493154 395325 493196 395561
rect 492876 388561 493196 395325
rect 492876 388325 492918 388561
rect 493154 388325 493196 388561
rect 492876 381561 493196 388325
rect 492876 381325 492918 381561
rect 493154 381325 493196 381561
rect 492876 374561 493196 381325
rect 492876 374325 492918 374561
rect 493154 374325 493196 374561
rect 492876 367561 493196 374325
rect 492876 367325 492918 367561
rect 493154 367325 493196 367561
rect 492876 360561 493196 367325
rect 492876 360325 492918 360561
rect 493154 360325 493196 360561
rect 492876 353561 493196 360325
rect 492876 353325 492918 353561
rect 493154 353325 493196 353561
rect 492876 346561 493196 353325
rect 492876 346325 492918 346561
rect 493154 346325 493196 346561
rect 492876 339561 493196 346325
rect 492876 339325 492918 339561
rect 493154 339325 493196 339561
rect 492876 332561 493196 339325
rect 492876 332325 492918 332561
rect 493154 332325 493196 332561
rect 492876 325561 493196 332325
rect 492876 325325 492918 325561
rect 493154 325325 493196 325561
rect 492876 318561 493196 325325
rect 492876 318325 492918 318561
rect 493154 318325 493196 318561
rect 492876 311561 493196 318325
rect 492876 311325 492918 311561
rect 493154 311325 493196 311561
rect 492876 304561 493196 311325
rect 492876 304325 492918 304561
rect 493154 304325 493196 304561
rect 492876 297561 493196 304325
rect 492876 297325 492918 297561
rect 493154 297325 493196 297561
rect 492876 290561 493196 297325
rect 492876 290325 492918 290561
rect 493154 290325 493196 290561
rect 492876 283561 493196 290325
rect 492876 283325 492918 283561
rect 493154 283325 493196 283561
rect 492876 276561 493196 283325
rect 492876 276325 492918 276561
rect 493154 276325 493196 276561
rect 492876 269561 493196 276325
rect 492876 269325 492918 269561
rect 493154 269325 493196 269561
rect 492876 262561 493196 269325
rect 492876 262325 492918 262561
rect 493154 262325 493196 262561
rect 492876 255561 493196 262325
rect 492876 255325 492918 255561
rect 493154 255325 493196 255561
rect 492876 248561 493196 255325
rect 492876 248325 492918 248561
rect 493154 248325 493196 248561
rect 492876 241561 493196 248325
rect 492876 241325 492918 241561
rect 493154 241325 493196 241561
rect 492876 234561 493196 241325
rect 492876 234325 492918 234561
rect 493154 234325 493196 234561
rect 492876 227561 493196 234325
rect 492876 227325 492918 227561
rect 493154 227325 493196 227561
rect 492876 220561 493196 227325
rect 492876 220325 492918 220561
rect 493154 220325 493196 220561
rect 492876 213561 493196 220325
rect 492876 213325 492918 213561
rect 493154 213325 493196 213561
rect 492876 206561 493196 213325
rect 492876 206325 492918 206561
rect 493154 206325 493196 206561
rect 492876 199561 493196 206325
rect 492876 199325 492918 199561
rect 493154 199325 493196 199561
rect 492876 192561 493196 199325
rect 492876 192325 492918 192561
rect 493154 192325 493196 192561
rect 492876 185561 493196 192325
rect 492876 185325 492918 185561
rect 493154 185325 493196 185561
rect 492876 178561 493196 185325
rect 492876 178325 492918 178561
rect 493154 178325 493196 178561
rect 492876 171561 493196 178325
rect 492876 171325 492918 171561
rect 493154 171325 493196 171561
rect 492876 164561 493196 171325
rect 492876 164325 492918 164561
rect 493154 164325 493196 164561
rect 492876 157561 493196 164325
rect 492876 157325 492918 157561
rect 493154 157325 493196 157561
rect 492876 150561 493196 157325
rect 492876 150325 492918 150561
rect 493154 150325 493196 150561
rect 492876 143561 493196 150325
rect 492876 143325 492918 143561
rect 493154 143325 493196 143561
rect 492876 136561 493196 143325
rect 492876 136325 492918 136561
rect 493154 136325 493196 136561
rect 492876 129561 493196 136325
rect 492876 129325 492918 129561
rect 493154 129325 493196 129561
rect 492876 122561 493196 129325
rect 492876 122325 492918 122561
rect 493154 122325 493196 122561
rect 492876 115561 493196 122325
rect 492876 115325 492918 115561
rect 493154 115325 493196 115561
rect 492876 108561 493196 115325
rect 492876 108325 492918 108561
rect 493154 108325 493196 108561
rect 492876 101561 493196 108325
rect 492876 101325 492918 101561
rect 493154 101325 493196 101561
rect 492876 94561 493196 101325
rect 492876 94325 492918 94561
rect 493154 94325 493196 94561
rect 492876 87561 493196 94325
rect 492876 87325 492918 87561
rect 493154 87325 493196 87561
rect 492876 80561 493196 87325
rect 492876 80325 492918 80561
rect 493154 80325 493196 80561
rect 492876 73561 493196 80325
rect 492876 73325 492918 73561
rect 493154 73325 493196 73561
rect 492876 66561 493196 73325
rect 492876 66325 492918 66561
rect 493154 66325 493196 66561
rect 492876 59561 493196 66325
rect 492876 59325 492918 59561
rect 493154 59325 493196 59561
rect 492876 52561 493196 59325
rect 492876 52325 492918 52561
rect 493154 52325 493196 52561
rect 492876 45561 493196 52325
rect 492876 45325 492918 45561
rect 493154 45325 493196 45561
rect 492876 38561 493196 45325
rect 492876 38325 492918 38561
rect 493154 38325 493196 38561
rect 492876 31561 493196 38325
rect 492876 31325 492918 31561
rect 493154 31325 493196 31561
rect 492876 24561 493196 31325
rect 492876 24325 492918 24561
rect 493154 24325 493196 24561
rect 492876 17561 493196 24325
rect 492876 17325 492918 17561
rect 493154 17325 493196 17561
rect 492876 10561 493196 17325
rect 492876 10325 492918 10561
rect 493154 10325 493196 10561
rect 492876 3561 493196 10325
rect 492876 3325 492918 3561
rect 493154 3325 493196 3561
rect 492876 -1706 493196 3325
rect 492876 -1942 492918 -1706
rect 493154 -1942 493196 -1706
rect 492876 -2026 493196 -1942
rect 492876 -2262 492918 -2026
rect 493154 -2262 493196 -2026
rect 492876 -2294 493196 -2262
rect 498144 705238 498464 706230
rect 498144 705002 498186 705238
rect 498422 705002 498464 705238
rect 498144 704918 498464 705002
rect 498144 704682 498186 704918
rect 498422 704682 498464 704918
rect 498144 695494 498464 704682
rect 498144 695258 498186 695494
rect 498422 695258 498464 695494
rect 498144 688494 498464 695258
rect 498144 688258 498186 688494
rect 498422 688258 498464 688494
rect 498144 681494 498464 688258
rect 498144 681258 498186 681494
rect 498422 681258 498464 681494
rect 498144 674494 498464 681258
rect 498144 674258 498186 674494
rect 498422 674258 498464 674494
rect 498144 667494 498464 674258
rect 498144 667258 498186 667494
rect 498422 667258 498464 667494
rect 498144 660494 498464 667258
rect 498144 660258 498186 660494
rect 498422 660258 498464 660494
rect 498144 653494 498464 660258
rect 498144 653258 498186 653494
rect 498422 653258 498464 653494
rect 498144 646494 498464 653258
rect 498144 646258 498186 646494
rect 498422 646258 498464 646494
rect 498144 639494 498464 646258
rect 498144 639258 498186 639494
rect 498422 639258 498464 639494
rect 498144 632494 498464 639258
rect 498144 632258 498186 632494
rect 498422 632258 498464 632494
rect 498144 625494 498464 632258
rect 498144 625258 498186 625494
rect 498422 625258 498464 625494
rect 498144 618494 498464 625258
rect 498144 618258 498186 618494
rect 498422 618258 498464 618494
rect 498144 611494 498464 618258
rect 498144 611258 498186 611494
rect 498422 611258 498464 611494
rect 498144 604494 498464 611258
rect 498144 604258 498186 604494
rect 498422 604258 498464 604494
rect 498144 597494 498464 604258
rect 498144 597258 498186 597494
rect 498422 597258 498464 597494
rect 498144 590494 498464 597258
rect 498144 590258 498186 590494
rect 498422 590258 498464 590494
rect 498144 583494 498464 590258
rect 498144 583258 498186 583494
rect 498422 583258 498464 583494
rect 498144 576494 498464 583258
rect 498144 576258 498186 576494
rect 498422 576258 498464 576494
rect 498144 569494 498464 576258
rect 498144 569258 498186 569494
rect 498422 569258 498464 569494
rect 498144 562494 498464 569258
rect 498144 562258 498186 562494
rect 498422 562258 498464 562494
rect 498144 555494 498464 562258
rect 498144 555258 498186 555494
rect 498422 555258 498464 555494
rect 498144 548494 498464 555258
rect 498144 548258 498186 548494
rect 498422 548258 498464 548494
rect 498144 541494 498464 548258
rect 498144 541258 498186 541494
rect 498422 541258 498464 541494
rect 498144 534494 498464 541258
rect 498144 534258 498186 534494
rect 498422 534258 498464 534494
rect 498144 527494 498464 534258
rect 498144 527258 498186 527494
rect 498422 527258 498464 527494
rect 498144 520494 498464 527258
rect 498144 520258 498186 520494
rect 498422 520258 498464 520494
rect 498144 513494 498464 520258
rect 498144 513258 498186 513494
rect 498422 513258 498464 513494
rect 498144 506494 498464 513258
rect 498144 506258 498186 506494
rect 498422 506258 498464 506494
rect 498144 499494 498464 506258
rect 498144 499258 498186 499494
rect 498422 499258 498464 499494
rect 498144 492494 498464 499258
rect 498144 492258 498186 492494
rect 498422 492258 498464 492494
rect 498144 485494 498464 492258
rect 498144 485258 498186 485494
rect 498422 485258 498464 485494
rect 498144 478494 498464 485258
rect 498144 478258 498186 478494
rect 498422 478258 498464 478494
rect 498144 471494 498464 478258
rect 498144 471258 498186 471494
rect 498422 471258 498464 471494
rect 498144 464494 498464 471258
rect 498144 464258 498186 464494
rect 498422 464258 498464 464494
rect 498144 457494 498464 464258
rect 498144 457258 498186 457494
rect 498422 457258 498464 457494
rect 498144 450494 498464 457258
rect 498144 450258 498186 450494
rect 498422 450258 498464 450494
rect 498144 443494 498464 450258
rect 498144 443258 498186 443494
rect 498422 443258 498464 443494
rect 498144 436494 498464 443258
rect 498144 436258 498186 436494
rect 498422 436258 498464 436494
rect 498144 429494 498464 436258
rect 498144 429258 498186 429494
rect 498422 429258 498464 429494
rect 498144 422494 498464 429258
rect 498144 422258 498186 422494
rect 498422 422258 498464 422494
rect 498144 415494 498464 422258
rect 498144 415258 498186 415494
rect 498422 415258 498464 415494
rect 498144 408494 498464 415258
rect 498144 408258 498186 408494
rect 498422 408258 498464 408494
rect 498144 401494 498464 408258
rect 498144 401258 498186 401494
rect 498422 401258 498464 401494
rect 498144 394494 498464 401258
rect 498144 394258 498186 394494
rect 498422 394258 498464 394494
rect 498144 387494 498464 394258
rect 498144 387258 498186 387494
rect 498422 387258 498464 387494
rect 498144 380494 498464 387258
rect 498144 380258 498186 380494
rect 498422 380258 498464 380494
rect 498144 373494 498464 380258
rect 498144 373258 498186 373494
rect 498422 373258 498464 373494
rect 498144 366494 498464 373258
rect 498144 366258 498186 366494
rect 498422 366258 498464 366494
rect 498144 359494 498464 366258
rect 498144 359258 498186 359494
rect 498422 359258 498464 359494
rect 498144 352494 498464 359258
rect 498144 352258 498186 352494
rect 498422 352258 498464 352494
rect 498144 345494 498464 352258
rect 498144 345258 498186 345494
rect 498422 345258 498464 345494
rect 498144 338494 498464 345258
rect 498144 338258 498186 338494
rect 498422 338258 498464 338494
rect 498144 331494 498464 338258
rect 498144 331258 498186 331494
rect 498422 331258 498464 331494
rect 498144 324494 498464 331258
rect 498144 324258 498186 324494
rect 498422 324258 498464 324494
rect 498144 317494 498464 324258
rect 498144 317258 498186 317494
rect 498422 317258 498464 317494
rect 498144 310494 498464 317258
rect 498144 310258 498186 310494
rect 498422 310258 498464 310494
rect 498144 303494 498464 310258
rect 498144 303258 498186 303494
rect 498422 303258 498464 303494
rect 498144 296494 498464 303258
rect 498144 296258 498186 296494
rect 498422 296258 498464 296494
rect 498144 289494 498464 296258
rect 498144 289258 498186 289494
rect 498422 289258 498464 289494
rect 498144 282494 498464 289258
rect 498144 282258 498186 282494
rect 498422 282258 498464 282494
rect 498144 275494 498464 282258
rect 498144 275258 498186 275494
rect 498422 275258 498464 275494
rect 498144 268494 498464 275258
rect 498144 268258 498186 268494
rect 498422 268258 498464 268494
rect 498144 261494 498464 268258
rect 498144 261258 498186 261494
rect 498422 261258 498464 261494
rect 498144 254494 498464 261258
rect 498144 254258 498186 254494
rect 498422 254258 498464 254494
rect 498144 247494 498464 254258
rect 498144 247258 498186 247494
rect 498422 247258 498464 247494
rect 498144 240494 498464 247258
rect 498144 240258 498186 240494
rect 498422 240258 498464 240494
rect 498144 233494 498464 240258
rect 498144 233258 498186 233494
rect 498422 233258 498464 233494
rect 498144 226494 498464 233258
rect 498144 226258 498186 226494
rect 498422 226258 498464 226494
rect 498144 219494 498464 226258
rect 498144 219258 498186 219494
rect 498422 219258 498464 219494
rect 498144 212494 498464 219258
rect 498144 212258 498186 212494
rect 498422 212258 498464 212494
rect 498144 205494 498464 212258
rect 498144 205258 498186 205494
rect 498422 205258 498464 205494
rect 498144 198494 498464 205258
rect 498144 198258 498186 198494
rect 498422 198258 498464 198494
rect 498144 191494 498464 198258
rect 498144 191258 498186 191494
rect 498422 191258 498464 191494
rect 498144 184494 498464 191258
rect 498144 184258 498186 184494
rect 498422 184258 498464 184494
rect 498144 177494 498464 184258
rect 498144 177258 498186 177494
rect 498422 177258 498464 177494
rect 498144 170494 498464 177258
rect 498144 170258 498186 170494
rect 498422 170258 498464 170494
rect 498144 163494 498464 170258
rect 498144 163258 498186 163494
rect 498422 163258 498464 163494
rect 498144 156494 498464 163258
rect 498144 156258 498186 156494
rect 498422 156258 498464 156494
rect 498144 149494 498464 156258
rect 498144 149258 498186 149494
rect 498422 149258 498464 149494
rect 498144 142494 498464 149258
rect 498144 142258 498186 142494
rect 498422 142258 498464 142494
rect 498144 135494 498464 142258
rect 498144 135258 498186 135494
rect 498422 135258 498464 135494
rect 498144 128494 498464 135258
rect 498144 128258 498186 128494
rect 498422 128258 498464 128494
rect 498144 121494 498464 128258
rect 498144 121258 498186 121494
rect 498422 121258 498464 121494
rect 498144 114494 498464 121258
rect 498144 114258 498186 114494
rect 498422 114258 498464 114494
rect 498144 107494 498464 114258
rect 498144 107258 498186 107494
rect 498422 107258 498464 107494
rect 498144 100494 498464 107258
rect 498144 100258 498186 100494
rect 498422 100258 498464 100494
rect 498144 93494 498464 100258
rect 498144 93258 498186 93494
rect 498422 93258 498464 93494
rect 498144 86494 498464 93258
rect 498144 86258 498186 86494
rect 498422 86258 498464 86494
rect 498144 79494 498464 86258
rect 498144 79258 498186 79494
rect 498422 79258 498464 79494
rect 498144 72494 498464 79258
rect 498144 72258 498186 72494
rect 498422 72258 498464 72494
rect 498144 65494 498464 72258
rect 498144 65258 498186 65494
rect 498422 65258 498464 65494
rect 498144 58494 498464 65258
rect 498144 58258 498186 58494
rect 498422 58258 498464 58494
rect 498144 51494 498464 58258
rect 498144 51258 498186 51494
rect 498422 51258 498464 51494
rect 498144 44494 498464 51258
rect 498144 44258 498186 44494
rect 498422 44258 498464 44494
rect 498144 37494 498464 44258
rect 498144 37258 498186 37494
rect 498422 37258 498464 37494
rect 498144 30494 498464 37258
rect 498144 30258 498186 30494
rect 498422 30258 498464 30494
rect 498144 23494 498464 30258
rect 498144 23258 498186 23494
rect 498422 23258 498464 23494
rect 498144 16494 498464 23258
rect 498144 16258 498186 16494
rect 498422 16258 498464 16494
rect 498144 9494 498464 16258
rect 498144 9258 498186 9494
rect 498422 9258 498464 9494
rect 498144 2494 498464 9258
rect 498144 2258 498186 2494
rect 498422 2258 498464 2494
rect 498144 -746 498464 2258
rect 498144 -982 498186 -746
rect 498422 -982 498464 -746
rect 498144 -1066 498464 -982
rect 498144 -1302 498186 -1066
rect 498422 -1302 498464 -1066
rect 498144 -2294 498464 -1302
rect 499876 706198 500196 706230
rect 499876 705962 499918 706198
rect 500154 705962 500196 706198
rect 499876 705878 500196 705962
rect 499876 705642 499918 705878
rect 500154 705642 500196 705878
rect 499876 696561 500196 705642
rect 499876 696325 499918 696561
rect 500154 696325 500196 696561
rect 499876 689561 500196 696325
rect 499876 689325 499918 689561
rect 500154 689325 500196 689561
rect 499876 682561 500196 689325
rect 499876 682325 499918 682561
rect 500154 682325 500196 682561
rect 499876 675561 500196 682325
rect 499876 675325 499918 675561
rect 500154 675325 500196 675561
rect 499876 668561 500196 675325
rect 499876 668325 499918 668561
rect 500154 668325 500196 668561
rect 499876 661561 500196 668325
rect 499876 661325 499918 661561
rect 500154 661325 500196 661561
rect 499876 654561 500196 661325
rect 499876 654325 499918 654561
rect 500154 654325 500196 654561
rect 499876 647561 500196 654325
rect 499876 647325 499918 647561
rect 500154 647325 500196 647561
rect 499876 640561 500196 647325
rect 499876 640325 499918 640561
rect 500154 640325 500196 640561
rect 499876 633561 500196 640325
rect 499876 633325 499918 633561
rect 500154 633325 500196 633561
rect 499876 626561 500196 633325
rect 499876 626325 499918 626561
rect 500154 626325 500196 626561
rect 499876 619561 500196 626325
rect 499876 619325 499918 619561
rect 500154 619325 500196 619561
rect 499876 612561 500196 619325
rect 499876 612325 499918 612561
rect 500154 612325 500196 612561
rect 499876 605561 500196 612325
rect 499876 605325 499918 605561
rect 500154 605325 500196 605561
rect 499876 598561 500196 605325
rect 499876 598325 499918 598561
rect 500154 598325 500196 598561
rect 499876 591561 500196 598325
rect 499876 591325 499918 591561
rect 500154 591325 500196 591561
rect 499876 584561 500196 591325
rect 499876 584325 499918 584561
rect 500154 584325 500196 584561
rect 499876 577561 500196 584325
rect 499876 577325 499918 577561
rect 500154 577325 500196 577561
rect 499876 570561 500196 577325
rect 499876 570325 499918 570561
rect 500154 570325 500196 570561
rect 499876 563561 500196 570325
rect 499876 563325 499918 563561
rect 500154 563325 500196 563561
rect 499876 556561 500196 563325
rect 499876 556325 499918 556561
rect 500154 556325 500196 556561
rect 499876 549561 500196 556325
rect 499876 549325 499918 549561
rect 500154 549325 500196 549561
rect 499876 542561 500196 549325
rect 499876 542325 499918 542561
rect 500154 542325 500196 542561
rect 499876 535561 500196 542325
rect 499876 535325 499918 535561
rect 500154 535325 500196 535561
rect 499876 528561 500196 535325
rect 499876 528325 499918 528561
rect 500154 528325 500196 528561
rect 499876 521561 500196 528325
rect 499876 521325 499918 521561
rect 500154 521325 500196 521561
rect 499876 514561 500196 521325
rect 499876 514325 499918 514561
rect 500154 514325 500196 514561
rect 499876 507561 500196 514325
rect 499876 507325 499918 507561
rect 500154 507325 500196 507561
rect 499876 500561 500196 507325
rect 499876 500325 499918 500561
rect 500154 500325 500196 500561
rect 499876 493561 500196 500325
rect 499876 493325 499918 493561
rect 500154 493325 500196 493561
rect 499876 486561 500196 493325
rect 499876 486325 499918 486561
rect 500154 486325 500196 486561
rect 499876 479561 500196 486325
rect 499876 479325 499918 479561
rect 500154 479325 500196 479561
rect 499876 472561 500196 479325
rect 499876 472325 499918 472561
rect 500154 472325 500196 472561
rect 499876 465561 500196 472325
rect 499876 465325 499918 465561
rect 500154 465325 500196 465561
rect 499876 458561 500196 465325
rect 499876 458325 499918 458561
rect 500154 458325 500196 458561
rect 499876 451561 500196 458325
rect 499876 451325 499918 451561
rect 500154 451325 500196 451561
rect 499876 444561 500196 451325
rect 499876 444325 499918 444561
rect 500154 444325 500196 444561
rect 499876 437561 500196 444325
rect 499876 437325 499918 437561
rect 500154 437325 500196 437561
rect 499876 430561 500196 437325
rect 499876 430325 499918 430561
rect 500154 430325 500196 430561
rect 499876 423561 500196 430325
rect 499876 423325 499918 423561
rect 500154 423325 500196 423561
rect 499876 416561 500196 423325
rect 499876 416325 499918 416561
rect 500154 416325 500196 416561
rect 499876 409561 500196 416325
rect 499876 409325 499918 409561
rect 500154 409325 500196 409561
rect 499876 402561 500196 409325
rect 499876 402325 499918 402561
rect 500154 402325 500196 402561
rect 499876 395561 500196 402325
rect 499876 395325 499918 395561
rect 500154 395325 500196 395561
rect 499876 388561 500196 395325
rect 499876 388325 499918 388561
rect 500154 388325 500196 388561
rect 499876 381561 500196 388325
rect 499876 381325 499918 381561
rect 500154 381325 500196 381561
rect 499876 374561 500196 381325
rect 499876 374325 499918 374561
rect 500154 374325 500196 374561
rect 499876 367561 500196 374325
rect 499876 367325 499918 367561
rect 500154 367325 500196 367561
rect 499876 360561 500196 367325
rect 499876 360325 499918 360561
rect 500154 360325 500196 360561
rect 499876 353561 500196 360325
rect 499876 353325 499918 353561
rect 500154 353325 500196 353561
rect 499876 346561 500196 353325
rect 499876 346325 499918 346561
rect 500154 346325 500196 346561
rect 499876 339561 500196 346325
rect 499876 339325 499918 339561
rect 500154 339325 500196 339561
rect 499876 332561 500196 339325
rect 499876 332325 499918 332561
rect 500154 332325 500196 332561
rect 499876 325561 500196 332325
rect 499876 325325 499918 325561
rect 500154 325325 500196 325561
rect 499876 318561 500196 325325
rect 499876 318325 499918 318561
rect 500154 318325 500196 318561
rect 499876 311561 500196 318325
rect 499876 311325 499918 311561
rect 500154 311325 500196 311561
rect 499876 304561 500196 311325
rect 499876 304325 499918 304561
rect 500154 304325 500196 304561
rect 499876 297561 500196 304325
rect 499876 297325 499918 297561
rect 500154 297325 500196 297561
rect 499876 290561 500196 297325
rect 499876 290325 499918 290561
rect 500154 290325 500196 290561
rect 499876 283561 500196 290325
rect 499876 283325 499918 283561
rect 500154 283325 500196 283561
rect 499876 276561 500196 283325
rect 499876 276325 499918 276561
rect 500154 276325 500196 276561
rect 499876 269561 500196 276325
rect 499876 269325 499918 269561
rect 500154 269325 500196 269561
rect 499876 262561 500196 269325
rect 499876 262325 499918 262561
rect 500154 262325 500196 262561
rect 499876 255561 500196 262325
rect 499876 255325 499918 255561
rect 500154 255325 500196 255561
rect 499876 248561 500196 255325
rect 499876 248325 499918 248561
rect 500154 248325 500196 248561
rect 499876 241561 500196 248325
rect 499876 241325 499918 241561
rect 500154 241325 500196 241561
rect 499876 234561 500196 241325
rect 499876 234325 499918 234561
rect 500154 234325 500196 234561
rect 499876 227561 500196 234325
rect 499876 227325 499918 227561
rect 500154 227325 500196 227561
rect 499876 220561 500196 227325
rect 499876 220325 499918 220561
rect 500154 220325 500196 220561
rect 499876 213561 500196 220325
rect 499876 213325 499918 213561
rect 500154 213325 500196 213561
rect 499876 206561 500196 213325
rect 499876 206325 499918 206561
rect 500154 206325 500196 206561
rect 499876 199561 500196 206325
rect 499876 199325 499918 199561
rect 500154 199325 500196 199561
rect 499876 192561 500196 199325
rect 499876 192325 499918 192561
rect 500154 192325 500196 192561
rect 499876 185561 500196 192325
rect 499876 185325 499918 185561
rect 500154 185325 500196 185561
rect 499876 178561 500196 185325
rect 499876 178325 499918 178561
rect 500154 178325 500196 178561
rect 499876 171561 500196 178325
rect 499876 171325 499918 171561
rect 500154 171325 500196 171561
rect 499876 164561 500196 171325
rect 499876 164325 499918 164561
rect 500154 164325 500196 164561
rect 499876 157561 500196 164325
rect 499876 157325 499918 157561
rect 500154 157325 500196 157561
rect 499876 150561 500196 157325
rect 499876 150325 499918 150561
rect 500154 150325 500196 150561
rect 499876 143561 500196 150325
rect 499876 143325 499918 143561
rect 500154 143325 500196 143561
rect 499876 136561 500196 143325
rect 499876 136325 499918 136561
rect 500154 136325 500196 136561
rect 499876 129561 500196 136325
rect 499876 129325 499918 129561
rect 500154 129325 500196 129561
rect 499876 122561 500196 129325
rect 499876 122325 499918 122561
rect 500154 122325 500196 122561
rect 499876 115561 500196 122325
rect 499876 115325 499918 115561
rect 500154 115325 500196 115561
rect 499876 108561 500196 115325
rect 499876 108325 499918 108561
rect 500154 108325 500196 108561
rect 499876 101561 500196 108325
rect 499876 101325 499918 101561
rect 500154 101325 500196 101561
rect 499876 94561 500196 101325
rect 499876 94325 499918 94561
rect 500154 94325 500196 94561
rect 499876 87561 500196 94325
rect 499876 87325 499918 87561
rect 500154 87325 500196 87561
rect 499876 80561 500196 87325
rect 499876 80325 499918 80561
rect 500154 80325 500196 80561
rect 499876 73561 500196 80325
rect 499876 73325 499918 73561
rect 500154 73325 500196 73561
rect 499876 66561 500196 73325
rect 499876 66325 499918 66561
rect 500154 66325 500196 66561
rect 499876 59561 500196 66325
rect 499876 59325 499918 59561
rect 500154 59325 500196 59561
rect 499876 52561 500196 59325
rect 499876 52325 499918 52561
rect 500154 52325 500196 52561
rect 499876 45561 500196 52325
rect 499876 45325 499918 45561
rect 500154 45325 500196 45561
rect 499876 38561 500196 45325
rect 499876 38325 499918 38561
rect 500154 38325 500196 38561
rect 499876 31561 500196 38325
rect 499876 31325 499918 31561
rect 500154 31325 500196 31561
rect 499876 24561 500196 31325
rect 499876 24325 499918 24561
rect 500154 24325 500196 24561
rect 499876 17561 500196 24325
rect 499876 17325 499918 17561
rect 500154 17325 500196 17561
rect 499876 10561 500196 17325
rect 499876 10325 499918 10561
rect 500154 10325 500196 10561
rect 499876 3561 500196 10325
rect 499876 3325 499918 3561
rect 500154 3325 500196 3561
rect 499876 -1706 500196 3325
rect 499876 -1942 499918 -1706
rect 500154 -1942 500196 -1706
rect 499876 -2026 500196 -1942
rect 499876 -2262 499918 -2026
rect 500154 -2262 500196 -2026
rect 499876 -2294 500196 -2262
rect 505144 705238 505464 706230
rect 505144 705002 505186 705238
rect 505422 705002 505464 705238
rect 505144 704918 505464 705002
rect 505144 704682 505186 704918
rect 505422 704682 505464 704918
rect 505144 695494 505464 704682
rect 505144 695258 505186 695494
rect 505422 695258 505464 695494
rect 505144 688494 505464 695258
rect 505144 688258 505186 688494
rect 505422 688258 505464 688494
rect 505144 681494 505464 688258
rect 505144 681258 505186 681494
rect 505422 681258 505464 681494
rect 505144 674494 505464 681258
rect 505144 674258 505186 674494
rect 505422 674258 505464 674494
rect 505144 667494 505464 674258
rect 505144 667258 505186 667494
rect 505422 667258 505464 667494
rect 505144 660494 505464 667258
rect 505144 660258 505186 660494
rect 505422 660258 505464 660494
rect 505144 653494 505464 660258
rect 505144 653258 505186 653494
rect 505422 653258 505464 653494
rect 505144 646494 505464 653258
rect 505144 646258 505186 646494
rect 505422 646258 505464 646494
rect 505144 639494 505464 646258
rect 505144 639258 505186 639494
rect 505422 639258 505464 639494
rect 505144 632494 505464 639258
rect 505144 632258 505186 632494
rect 505422 632258 505464 632494
rect 505144 625494 505464 632258
rect 505144 625258 505186 625494
rect 505422 625258 505464 625494
rect 505144 618494 505464 625258
rect 505144 618258 505186 618494
rect 505422 618258 505464 618494
rect 505144 611494 505464 618258
rect 505144 611258 505186 611494
rect 505422 611258 505464 611494
rect 505144 604494 505464 611258
rect 505144 604258 505186 604494
rect 505422 604258 505464 604494
rect 505144 597494 505464 604258
rect 505144 597258 505186 597494
rect 505422 597258 505464 597494
rect 505144 590494 505464 597258
rect 505144 590258 505186 590494
rect 505422 590258 505464 590494
rect 505144 583494 505464 590258
rect 505144 583258 505186 583494
rect 505422 583258 505464 583494
rect 505144 576494 505464 583258
rect 505144 576258 505186 576494
rect 505422 576258 505464 576494
rect 505144 569494 505464 576258
rect 505144 569258 505186 569494
rect 505422 569258 505464 569494
rect 505144 562494 505464 569258
rect 505144 562258 505186 562494
rect 505422 562258 505464 562494
rect 505144 555494 505464 562258
rect 505144 555258 505186 555494
rect 505422 555258 505464 555494
rect 505144 548494 505464 555258
rect 505144 548258 505186 548494
rect 505422 548258 505464 548494
rect 505144 541494 505464 548258
rect 505144 541258 505186 541494
rect 505422 541258 505464 541494
rect 505144 534494 505464 541258
rect 505144 534258 505186 534494
rect 505422 534258 505464 534494
rect 505144 527494 505464 534258
rect 505144 527258 505186 527494
rect 505422 527258 505464 527494
rect 505144 520494 505464 527258
rect 505144 520258 505186 520494
rect 505422 520258 505464 520494
rect 505144 513494 505464 520258
rect 505144 513258 505186 513494
rect 505422 513258 505464 513494
rect 505144 506494 505464 513258
rect 505144 506258 505186 506494
rect 505422 506258 505464 506494
rect 505144 499494 505464 506258
rect 505144 499258 505186 499494
rect 505422 499258 505464 499494
rect 505144 492494 505464 499258
rect 505144 492258 505186 492494
rect 505422 492258 505464 492494
rect 505144 485494 505464 492258
rect 505144 485258 505186 485494
rect 505422 485258 505464 485494
rect 505144 478494 505464 485258
rect 505144 478258 505186 478494
rect 505422 478258 505464 478494
rect 505144 471494 505464 478258
rect 505144 471258 505186 471494
rect 505422 471258 505464 471494
rect 505144 464494 505464 471258
rect 505144 464258 505186 464494
rect 505422 464258 505464 464494
rect 505144 457494 505464 464258
rect 505144 457258 505186 457494
rect 505422 457258 505464 457494
rect 505144 450494 505464 457258
rect 505144 450258 505186 450494
rect 505422 450258 505464 450494
rect 505144 443494 505464 450258
rect 505144 443258 505186 443494
rect 505422 443258 505464 443494
rect 505144 436494 505464 443258
rect 505144 436258 505186 436494
rect 505422 436258 505464 436494
rect 505144 429494 505464 436258
rect 505144 429258 505186 429494
rect 505422 429258 505464 429494
rect 505144 422494 505464 429258
rect 505144 422258 505186 422494
rect 505422 422258 505464 422494
rect 505144 415494 505464 422258
rect 505144 415258 505186 415494
rect 505422 415258 505464 415494
rect 505144 408494 505464 415258
rect 505144 408258 505186 408494
rect 505422 408258 505464 408494
rect 505144 401494 505464 408258
rect 505144 401258 505186 401494
rect 505422 401258 505464 401494
rect 505144 394494 505464 401258
rect 505144 394258 505186 394494
rect 505422 394258 505464 394494
rect 505144 387494 505464 394258
rect 505144 387258 505186 387494
rect 505422 387258 505464 387494
rect 505144 380494 505464 387258
rect 505144 380258 505186 380494
rect 505422 380258 505464 380494
rect 505144 373494 505464 380258
rect 505144 373258 505186 373494
rect 505422 373258 505464 373494
rect 505144 366494 505464 373258
rect 505144 366258 505186 366494
rect 505422 366258 505464 366494
rect 505144 359494 505464 366258
rect 505144 359258 505186 359494
rect 505422 359258 505464 359494
rect 505144 352494 505464 359258
rect 505144 352258 505186 352494
rect 505422 352258 505464 352494
rect 505144 345494 505464 352258
rect 505144 345258 505186 345494
rect 505422 345258 505464 345494
rect 505144 338494 505464 345258
rect 505144 338258 505186 338494
rect 505422 338258 505464 338494
rect 505144 331494 505464 338258
rect 505144 331258 505186 331494
rect 505422 331258 505464 331494
rect 505144 324494 505464 331258
rect 505144 324258 505186 324494
rect 505422 324258 505464 324494
rect 505144 317494 505464 324258
rect 505144 317258 505186 317494
rect 505422 317258 505464 317494
rect 505144 310494 505464 317258
rect 505144 310258 505186 310494
rect 505422 310258 505464 310494
rect 505144 303494 505464 310258
rect 505144 303258 505186 303494
rect 505422 303258 505464 303494
rect 505144 296494 505464 303258
rect 505144 296258 505186 296494
rect 505422 296258 505464 296494
rect 505144 289494 505464 296258
rect 505144 289258 505186 289494
rect 505422 289258 505464 289494
rect 505144 282494 505464 289258
rect 505144 282258 505186 282494
rect 505422 282258 505464 282494
rect 505144 275494 505464 282258
rect 505144 275258 505186 275494
rect 505422 275258 505464 275494
rect 505144 268494 505464 275258
rect 505144 268258 505186 268494
rect 505422 268258 505464 268494
rect 505144 261494 505464 268258
rect 505144 261258 505186 261494
rect 505422 261258 505464 261494
rect 505144 254494 505464 261258
rect 505144 254258 505186 254494
rect 505422 254258 505464 254494
rect 505144 247494 505464 254258
rect 505144 247258 505186 247494
rect 505422 247258 505464 247494
rect 505144 240494 505464 247258
rect 505144 240258 505186 240494
rect 505422 240258 505464 240494
rect 505144 233494 505464 240258
rect 505144 233258 505186 233494
rect 505422 233258 505464 233494
rect 505144 226494 505464 233258
rect 505144 226258 505186 226494
rect 505422 226258 505464 226494
rect 505144 219494 505464 226258
rect 505144 219258 505186 219494
rect 505422 219258 505464 219494
rect 505144 212494 505464 219258
rect 505144 212258 505186 212494
rect 505422 212258 505464 212494
rect 505144 205494 505464 212258
rect 505144 205258 505186 205494
rect 505422 205258 505464 205494
rect 505144 198494 505464 205258
rect 505144 198258 505186 198494
rect 505422 198258 505464 198494
rect 505144 191494 505464 198258
rect 505144 191258 505186 191494
rect 505422 191258 505464 191494
rect 505144 184494 505464 191258
rect 505144 184258 505186 184494
rect 505422 184258 505464 184494
rect 505144 177494 505464 184258
rect 505144 177258 505186 177494
rect 505422 177258 505464 177494
rect 505144 170494 505464 177258
rect 505144 170258 505186 170494
rect 505422 170258 505464 170494
rect 505144 163494 505464 170258
rect 505144 163258 505186 163494
rect 505422 163258 505464 163494
rect 505144 156494 505464 163258
rect 505144 156258 505186 156494
rect 505422 156258 505464 156494
rect 505144 149494 505464 156258
rect 505144 149258 505186 149494
rect 505422 149258 505464 149494
rect 505144 142494 505464 149258
rect 505144 142258 505186 142494
rect 505422 142258 505464 142494
rect 505144 135494 505464 142258
rect 505144 135258 505186 135494
rect 505422 135258 505464 135494
rect 505144 128494 505464 135258
rect 505144 128258 505186 128494
rect 505422 128258 505464 128494
rect 505144 121494 505464 128258
rect 505144 121258 505186 121494
rect 505422 121258 505464 121494
rect 505144 114494 505464 121258
rect 505144 114258 505186 114494
rect 505422 114258 505464 114494
rect 505144 107494 505464 114258
rect 505144 107258 505186 107494
rect 505422 107258 505464 107494
rect 505144 100494 505464 107258
rect 505144 100258 505186 100494
rect 505422 100258 505464 100494
rect 505144 93494 505464 100258
rect 505144 93258 505186 93494
rect 505422 93258 505464 93494
rect 505144 86494 505464 93258
rect 505144 86258 505186 86494
rect 505422 86258 505464 86494
rect 505144 79494 505464 86258
rect 505144 79258 505186 79494
rect 505422 79258 505464 79494
rect 505144 72494 505464 79258
rect 505144 72258 505186 72494
rect 505422 72258 505464 72494
rect 505144 65494 505464 72258
rect 505144 65258 505186 65494
rect 505422 65258 505464 65494
rect 505144 58494 505464 65258
rect 505144 58258 505186 58494
rect 505422 58258 505464 58494
rect 505144 51494 505464 58258
rect 505144 51258 505186 51494
rect 505422 51258 505464 51494
rect 505144 44494 505464 51258
rect 505144 44258 505186 44494
rect 505422 44258 505464 44494
rect 505144 37494 505464 44258
rect 505144 37258 505186 37494
rect 505422 37258 505464 37494
rect 505144 30494 505464 37258
rect 505144 30258 505186 30494
rect 505422 30258 505464 30494
rect 505144 23494 505464 30258
rect 505144 23258 505186 23494
rect 505422 23258 505464 23494
rect 505144 16494 505464 23258
rect 505144 16258 505186 16494
rect 505422 16258 505464 16494
rect 505144 9494 505464 16258
rect 505144 9258 505186 9494
rect 505422 9258 505464 9494
rect 505144 2494 505464 9258
rect 505144 2258 505186 2494
rect 505422 2258 505464 2494
rect 505144 -746 505464 2258
rect 505144 -982 505186 -746
rect 505422 -982 505464 -746
rect 505144 -1066 505464 -982
rect 505144 -1302 505186 -1066
rect 505422 -1302 505464 -1066
rect 505144 -2294 505464 -1302
rect 506876 706198 507196 706230
rect 506876 705962 506918 706198
rect 507154 705962 507196 706198
rect 506876 705878 507196 705962
rect 506876 705642 506918 705878
rect 507154 705642 507196 705878
rect 506876 696561 507196 705642
rect 506876 696325 506918 696561
rect 507154 696325 507196 696561
rect 506876 689561 507196 696325
rect 506876 689325 506918 689561
rect 507154 689325 507196 689561
rect 506876 682561 507196 689325
rect 506876 682325 506918 682561
rect 507154 682325 507196 682561
rect 506876 675561 507196 682325
rect 506876 675325 506918 675561
rect 507154 675325 507196 675561
rect 506876 668561 507196 675325
rect 506876 668325 506918 668561
rect 507154 668325 507196 668561
rect 506876 661561 507196 668325
rect 506876 661325 506918 661561
rect 507154 661325 507196 661561
rect 506876 654561 507196 661325
rect 506876 654325 506918 654561
rect 507154 654325 507196 654561
rect 506876 647561 507196 654325
rect 506876 647325 506918 647561
rect 507154 647325 507196 647561
rect 506876 640561 507196 647325
rect 506876 640325 506918 640561
rect 507154 640325 507196 640561
rect 506876 633561 507196 640325
rect 506876 633325 506918 633561
rect 507154 633325 507196 633561
rect 506876 626561 507196 633325
rect 506876 626325 506918 626561
rect 507154 626325 507196 626561
rect 506876 619561 507196 626325
rect 506876 619325 506918 619561
rect 507154 619325 507196 619561
rect 506876 612561 507196 619325
rect 506876 612325 506918 612561
rect 507154 612325 507196 612561
rect 506876 605561 507196 612325
rect 506876 605325 506918 605561
rect 507154 605325 507196 605561
rect 506876 598561 507196 605325
rect 506876 598325 506918 598561
rect 507154 598325 507196 598561
rect 506876 591561 507196 598325
rect 506876 591325 506918 591561
rect 507154 591325 507196 591561
rect 506876 584561 507196 591325
rect 506876 584325 506918 584561
rect 507154 584325 507196 584561
rect 506876 577561 507196 584325
rect 506876 577325 506918 577561
rect 507154 577325 507196 577561
rect 506876 570561 507196 577325
rect 506876 570325 506918 570561
rect 507154 570325 507196 570561
rect 506876 563561 507196 570325
rect 506876 563325 506918 563561
rect 507154 563325 507196 563561
rect 506876 556561 507196 563325
rect 506876 556325 506918 556561
rect 507154 556325 507196 556561
rect 506876 549561 507196 556325
rect 506876 549325 506918 549561
rect 507154 549325 507196 549561
rect 506876 542561 507196 549325
rect 506876 542325 506918 542561
rect 507154 542325 507196 542561
rect 506876 535561 507196 542325
rect 506876 535325 506918 535561
rect 507154 535325 507196 535561
rect 506876 528561 507196 535325
rect 506876 528325 506918 528561
rect 507154 528325 507196 528561
rect 506876 521561 507196 528325
rect 506876 521325 506918 521561
rect 507154 521325 507196 521561
rect 506876 514561 507196 521325
rect 506876 514325 506918 514561
rect 507154 514325 507196 514561
rect 506876 507561 507196 514325
rect 506876 507325 506918 507561
rect 507154 507325 507196 507561
rect 506876 500561 507196 507325
rect 506876 500325 506918 500561
rect 507154 500325 507196 500561
rect 506876 493561 507196 500325
rect 506876 493325 506918 493561
rect 507154 493325 507196 493561
rect 506876 486561 507196 493325
rect 506876 486325 506918 486561
rect 507154 486325 507196 486561
rect 506876 479561 507196 486325
rect 506876 479325 506918 479561
rect 507154 479325 507196 479561
rect 506876 472561 507196 479325
rect 506876 472325 506918 472561
rect 507154 472325 507196 472561
rect 506876 465561 507196 472325
rect 506876 465325 506918 465561
rect 507154 465325 507196 465561
rect 506876 458561 507196 465325
rect 506876 458325 506918 458561
rect 507154 458325 507196 458561
rect 506876 451561 507196 458325
rect 506876 451325 506918 451561
rect 507154 451325 507196 451561
rect 506876 444561 507196 451325
rect 506876 444325 506918 444561
rect 507154 444325 507196 444561
rect 506876 437561 507196 444325
rect 506876 437325 506918 437561
rect 507154 437325 507196 437561
rect 506876 430561 507196 437325
rect 506876 430325 506918 430561
rect 507154 430325 507196 430561
rect 506876 423561 507196 430325
rect 506876 423325 506918 423561
rect 507154 423325 507196 423561
rect 506876 416561 507196 423325
rect 506876 416325 506918 416561
rect 507154 416325 507196 416561
rect 506876 409561 507196 416325
rect 506876 409325 506918 409561
rect 507154 409325 507196 409561
rect 506876 402561 507196 409325
rect 506876 402325 506918 402561
rect 507154 402325 507196 402561
rect 506876 395561 507196 402325
rect 506876 395325 506918 395561
rect 507154 395325 507196 395561
rect 506876 388561 507196 395325
rect 506876 388325 506918 388561
rect 507154 388325 507196 388561
rect 506876 381561 507196 388325
rect 506876 381325 506918 381561
rect 507154 381325 507196 381561
rect 506876 374561 507196 381325
rect 506876 374325 506918 374561
rect 507154 374325 507196 374561
rect 506876 367561 507196 374325
rect 506876 367325 506918 367561
rect 507154 367325 507196 367561
rect 506876 360561 507196 367325
rect 506876 360325 506918 360561
rect 507154 360325 507196 360561
rect 506876 353561 507196 360325
rect 506876 353325 506918 353561
rect 507154 353325 507196 353561
rect 506876 346561 507196 353325
rect 506876 346325 506918 346561
rect 507154 346325 507196 346561
rect 506876 339561 507196 346325
rect 506876 339325 506918 339561
rect 507154 339325 507196 339561
rect 506876 332561 507196 339325
rect 506876 332325 506918 332561
rect 507154 332325 507196 332561
rect 506876 325561 507196 332325
rect 506876 325325 506918 325561
rect 507154 325325 507196 325561
rect 506876 318561 507196 325325
rect 506876 318325 506918 318561
rect 507154 318325 507196 318561
rect 506876 311561 507196 318325
rect 506876 311325 506918 311561
rect 507154 311325 507196 311561
rect 506876 304561 507196 311325
rect 506876 304325 506918 304561
rect 507154 304325 507196 304561
rect 506876 297561 507196 304325
rect 506876 297325 506918 297561
rect 507154 297325 507196 297561
rect 506876 290561 507196 297325
rect 506876 290325 506918 290561
rect 507154 290325 507196 290561
rect 506876 283561 507196 290325
rect 506876 283325 506918 283561
rect 507154 283325 507196 283561
rect 506876 276561 507196 283325
rect 506876 276325 506918 276561
rect 507154 276325 507196 276561
rect 506876 269561 507196 276325
rect 506876 269325 506918 269561
rect 507154 269325 507196 269561
rect 506876 262561 507196 269325
rect 506876 262325 506918 262561
rect 507154 262325 507196 262561
rect 506876 255561 507196 262325
rect 506876 255325 506918 255561
rect 507154 255325 507196 255561
rect 506876 248561 507196 255325
rect 506876 248325 506918 248561
rect 507154 248325 507196 248561
rect 506876 241561 507196 248325
rect 506876 241325 506918 241561
rect 507154 241325 507196 241561
rect 506876 234561 507196 241325
rect 506876 234325 506918 234561
rect 507154 234325 507196 234561
rect 506876 227561 507196 234325
rect 506876 227325 506918 227561
rect 507154 227325 507196 227561
rect 506876 220561 507196 227325
rect 506876 220325 506918 220561
rect 507154 220325 507196 220561
rect 506876 213561 507196 220325
rect 506876 213325 506918 213561
rect 507154 213325 507196 213561
rect 506876 206561 507196 213325
rect 506876 206325 506918 206561
rect 507154 206325 507196 206561
rect 506876 199561 507196 206325
rect 506876 199325 506918 199561
rect 507154 199325 507196 199561
rect 506876 192561 507196 199325
rect 506876 192325 506918 192561
rect 507154 192325 507196 192561
rect 506876 185561 507196 192325
rect 506876 185325 506918 185561
rect 507154 185325 507196 185561
rect 506876 178561 507196 185325
rect 506876 178325 506918 178561
rect 507154 178325 507196 178561
rect 506876 171561 507196 178325
rect 506876 171325 506918 171561
rect 507154 171325 507196 171561
rect 506876 164561 507196 171325
rect 506876 164325 506918 164561
rect 507154 164325 507196 164561
rect 506876 157561 507196 164325
rect 506876 157325 506918 157561
rect 507154 157325 507196 157561
rect 506876 150561 507196 157325
rect 506876 150325 506918 150561
rect 507154 150325 507196 150561
rect 506876 143561 507196 150325
rect 506876 143325 506918 143561
rect 507154 143325 507196 143561
rect 506876 136561 507196 143325
rect 506876 136325 506918 136561
rect 507154 136325 507196 136561
rect 506876 129561 507196 136325
rect 506876 129325 506918 129561
rect 507154 129325 507196 129561
rect 506876 122561 507196 129325
rect 506876 122325 506918 122561
rect 507154 122325 507196 122561
rect 506876 115561 507196 122325
rect 506876 115325 506918 115561
rect 507154 115325 507196 115561
rect 506876 108561 507196 115325
rect 506876 108325 506918 108561
rect 507154 108325 507196 108561
rect 506876 101561 507196 108325
rect 506876 101325 506918 101561
rect 507154 101325 507196 101561
rect 506876 94561 507196 101325
rect 506876 94325 506918 94561
rect 507154 94325 507196 94561
rect 506876 87561 507196 94325
rect 506876 87325 506918 87561
rect 507154 87325 507196 87561
rect 506876 80561 507196 87325
rect 506876 80325 506918 80561
rect 507154 80325 507196 80561
rect 506876 73561 507196 80325
rect 506876 73325 506918 73561
rect 507154 73325 507196 73561
rect 506876 66561 507196 73325
rect 506876 66325 506918 66561
rect 507154 66325 507196 66561
rect 506876 59561 507196 66325
rect 506876 59325 506918 59561
rect 507154 59325 507196 59561
rect 506876 52561 507196 59325
rect 506876 52325 506918 52561
rect 507154 52325 507196 52561
rect 506876 45561 507196 52325
rect 506876 45325 506918 45561
rect 507154 45325 507196 45561
rect 506876 38561 507196 45325
rect 506876 38325 506918 38561
rect 507154 38325 507196 38561
rect 506876 31561 507196 38325
rect 506876 31325 506918 31561
rect 507154 31325 507196 31561
rect 506876 24561 507196 31325
rect 506876 24325 506918 24561
rect 507154 24325 507196 24561
rect 506876 17561 507196 24325
rect 506876 17325 506918 17561
rect 507154 17325 507196 17561
rect 506876 10561 507196 17325
rect 506876 10325 506918 10561
rect 507154 10325 507196 10561
rect 506876 3561 507196 10325
rect 506876 3325 506918 3561
rect 507154 3325 507196 3561
rect 506876 -1706 507196 3325
rect 506876 -1942 506918 -1706
rect 507154 -1942 507196 -1706
rect 506876 -2026 507196 -1942
rect 506876 -2262 506918 -2026
rect 507154 -2262 507196 -2026
rect 506876 -2294 507196 -2262
rect 512144 705238 512464 706230
rect 512144 705002 512186 705238
rect 512422 705002 512464 705238
rect 512144 704918 512464 705002
rect 512144 704682 512186 704918
rect 512422 704682 512464 704918
rect 512144 695494 512464 704682
rect 512144 695258 512186 695494
rect 512422 695258 512464 695494
rect 512144 688494 512464 695258
rect 512144 688258 512186 688494
rect 512422 688258 512464 688494
rect 512144 681494 512464 688258
rect 512144 681258 512186 681494
rect 512422 681258 512464 681494
rect 512144 674494 512464 681258
rect 512144 674258 512186 674494
rect 512422 674258 512464 674494
rect 512144 667494 512464 674258
rect 512144 667258 512186 667494
rect 512422 667258 512464 667494
rect 512144 660494 512464 667258
rect 512144 660258 512186 660494
rect 512422 660258 512464 660494
rect 512144 653494 512464 660258
rect 512144 653258 512186 653494
rect 512422 653258 512464 653494
rect 512144 646494 512464 653258
rect 512144 646258 512186 646494
rect 512422 646258 512464 646494
rect 512144 639494 512464 646258
rect 512144 639258 512186 639494
rect 512422 639258 512464 639494
rect 512144 632494 512464 639258
rect 512144 632258 512186 632494
rect 512422 632258 512464 632494
rect 512144 625494 512464 632258
rect 512144 625258 512186 625494
rect 512422 625258 512464 625494
rect 512144 618494 512464 625258
rect 512144 618258 512186 618494
rect 512422 618258 512464 618494
rect 512144 611494 512464 618258
rect 512144 611258 512186 611494
rect 512422 611258 512464 611494
rect 512144 604494 512464 611258
rect 512144 604258 512186 604494
rect 512422 604258 512464 604494
rect 512144 597494 512464 604258
rect 512144 597258 512186 597494
rect 512422 597258 512464 597494
rect 512144 590494 512464 597258
rect 512144 590258 512186 590494
rect 512422 590258 512464 590494
rect 512144 583494 512464 590258
rect 512144 583258 512186 583494
rect 512422 583258 512464 583494
rect 512144 576494 512464 583258
rect 512144 576258 512186 576494
rect 512422 576258 512464 576494
rect 512144 569494 512464 576258
rect 512144 569258 512186 569494
rect 512422 569258 512464 569494
rect 512144 562494 512464 569258
rect 512144 562258 512186 562494
rect 512422 562258 512464 562494
rect 512144 555494 512464 562258
rect 512144 555258 512186 555494
rect 512422 555258 512464 555494
rect 512144 548494 512464 555258
rect 512144 548258 512186 548494
rect 512422 548258 512464 548494
rect 512144 541494 512464 548258
rect 512144 541258 512186 541494
rect 512422 541258 512464 541494
rect 512144 534494 512464 541258
rect 512144 534258 512186 534494
rect 512422 534258 512464 534494
rect 512144 527494 512464 534258
rect 512144 527258 512186 527494
rect 512422 527258 512464 527494
rect 512144 520494 512464 527258
rect 512144 520258 512186 520494
rect 512422 520258 512464 520494
rect 512144 513494 512464 520258
rect 512144 513258 512186 513494
rect 512422 513258 512464 513494
rect 512144 506494 512464 513258
rect 512144 506258 512186 506494
rect 512422 506258 512464 506494
rect 512144 499494 512464 506258
rect 512144 499258 512186 499494
rect 512422 499258 512464 499494
rect 512144 492494 512464 499258
rect 512144 492258 512186 492494
rect 512422 492258 512464 492494
rect 512144 485494 512464 492258
rect 512144 485258 512186 485494
rect 512422 485258 512464 485494
rect 512144 478494 512464 485258
rect 512144 478258 512186 478494
rect 512422 478258 512464 478494
rect 512144 471494 512464 478258
rect 512144 471258 512186 471494
rect 512422 471258 512464 471494
rect 512144 464494 512464 471258
rect 512144 464258 512186 464494
rect 512422 464258 512464 464494
rect 512144 457494 512464 464258
rect 512144 457258 512186 457494
rect 512422 457258 512464 457494
rect 512144 450494 512464 457258
rect 512144 450258 512186 450494
rect 512422 450258 512464 450494
rect 512144 443494 512464 450258
rect 512144 443258 512186 443494
rect 512422 443258 512464 443494
rect 512144 436494 512464 443258
rect 512144 436258 512186 436494
rect 512422 436258 512464 436494
rect 512144 429494 512464 436258
rect 512144 429258 512186 429494
rect 512422 429258 512464 429494
rect 512144 422494 512464 429258
rect 512144 422258 512186 422494
rect 512422 422258 512464 422494
rect 512144 415494 512464 422258
rect 512144 415258 512186 415494
rect 512422 415258 512464 415494
rect 512144 408494 512464 415258
rect 512144 408258 512186 408494
rect 512422 408258 512464 408494
rect 512144 401494 512464 408258
rect 512144 401258 512186 401494
rect 512422 401258 512464 401494
rect 512144 394494 512464 401258
rect 512144 394258 512186 394494
rect 512422 394258 512464 394494
rect 512144 387494 512464 394258
rect 512144 387258 512186 387494
rect 512422 387258 512464 387494
rect 512144 380494 512464 387258
rect 512144 380258 512186 380494
rect 512422 380258 512464 380494
rect 512144 373494 512464 380258
rect 512144 373258 512186 373494
rect 512422 373258 512464 373494
rect 512144 366494 512464 373258
rect 512144 366258 512186 366494
rect 512422 366258 512464 366494
rect 512144 359494 512464 366258
rect 512144 359258 512186 359494
rect 512422 359258 512464 359494
rect 512144 352494 512464 359258
rect 512144 352258 512186 352494
rect 512422 352258 512464 352494
rect 512144 345494 512464 352258
rect 512144 345258 512186 345494
rect 512422 345258 512464 345494
rect 512144 338494 512464 345258
rect 512144 338258 512186 338494
rect 512422 338258 512464 338494
rect 512144 331494 512464 338258
rect 512144 331258 512186 331494
rect 512422 331258 512464 331494
rect 512144 324494 512464 331258
rect 512144 324258 512186 324494
rect 512422 324258 512464 324494
rect 512144 317494 512464 324258
rect 512144 317258 512186 317494
rect 512422 317258 512464 317494
rect 512144 310494 512464 317258
rect 512144 310258 512186 310494
rect 512422 310258 512464 310494
rect 512144 303494 512464 310258
rect 512144 303258 512186 303494
rect 512422 303258 512464 303494
rect 512144 296494 512464 303258
rect 512144 296258 512186 296494
rect 512422 296258 512464 296494
rect 512144 289494 512464 296258
rect 512144 289258 512186 289494
rect 512422 289258 512464 289494
rect 512144 282494 512464 289258
rect 512144 282258 512186 282494
rect 512422 282258 512464 282494
rect 512144 275494 512464 282258
rect 512144 275258 512186 275494
rect 512422 275258 512464 275494
rect 512144 268494 512464 275258
rect 512144 268258 512186 268494
rect 512422 268258 512464 268494
rect 512144 261494 512464 268258
rect 512144 261258 512186 261494
rect 512422 261258 512464 261494
rect 512144 254494 512464 261258
rect 512144 254258 512186 254494
rect 512422 254258 512464 254494
rect 512144 247494 512464 254258
rect 512144 247258 512186 247494
rect 512422 247258 512464 247494
rect 512144 240494 512464 247258
rect 512144 240258 512186 240494
rect 512422 240258 512464 240494
rect 512144 233494 512464 240258
rect 512144 233258 512186 233494
rect 512422 233258 512464 233494
rect 512144 226494 512464 233258
rect 512144 226258 512186 226494
rect 512422 226258 512464 226494
rect 512144 219494 512464 226258
rect 512144 219258 512186 219494
rect 512422 219258 512464 219494
rect 512144 212494 512464 219258
rect 512144 212258 512186 212494
rect 512422 212258 512464 212494
rect 512144 205494 512464 212258
rect 512144 205258 512186 205494
rect 512422 205258 512464 205494
rect 512144 198494 512464 205258
rect 512144 198258 512186 198494
rect 512422 198258 512464 198494
rect 512144 191494 512464 198258
rect 512144 191258 512186 191494
rect 512422 191258 512464 191494
rect 512144 184494 512464 191258
rect 512144 184258 512186 184494
rect 512422 184258 512464 184494
rect 512144 177494 512464 184258
rect 512144 177258 512186 177494
rect 512422 177258 512464 177494
rect 512144 170494 512464 177258
rect 512144 170258 512186 170494
rect 512422 170258 512464 170494
rect 512144 163494 512464 170258
rect 512144 163258 512186 163494
rect 512422 163258 512464 163494
rect 512144 156494 512464 163258
rect 512144 156258 512186 156494
rect 512422 156258 512464 156494
rect 512144 149494 512464 156258
rect 512144 149258 512186 149494
rect 512422 149258 512464 149494
rect 512144 142494 512464 149258
rect 512144 142258 512186 142494
rect 512422 142258 512464 142494
rect 512144 135494 512464 142258
rect 512144 135258 512186 135494
rect 512422 135258 512464 135494
rect 512144 128494 512464 135258
rect 512144 128258 512186 128494
rect 512422 128258 512464 128494
rect 512144 121494 512464 128258
rect 512144 121258 512186 121494
rect 512422 121258 512464 121494
rect 512144 114494 512464 121258
rect 512144 114258 512186 114494
rect 512422 114258 512464 114494
rect 512144 107494 512464 114258
rect 512144 107258 512186 107494
rect 512422 107258 512464 107494
rect 512144 100494 512464 107258
rect 512144 100258 512186 100494
rect 512422 100258 512464 100494
rect 512144 93494 512464 100258
rect 512144 93258 512186 93494
rect 512422 93258 512464 93494
rect 512144 86494 512464 93258
rect 512144 86258 512186 86494
rect 512422 86258 512464 86494
rect 512144 79494 512464 86258
rect 512144 79258 512186 79494
rect 512422 79258 512464 79494
rect 512144 72494 512464 79258
rect 512144 72258 512186 72494
rect 512422 72258 512464 72494
rect 512144 65494 512464 72258
rect 512144 65258 512186 65494
rect 512422 65258 512464 65494
rect 512144 58494 512464 65258
rect 512144 58258 512186 58494
rect 512422 58258 512464 58494
rect 512144 51494 512464 58258
rect 512144 51258 512186 51494
rect 512422 51258 512464 51494
rect 512144 44494 512464 51258
rect 512144 44258 512186 44494
rect 512422 44258 512464 44494
rect 512144 37494 512464 44258
rect 512144 37258 512186 37494
rect 512422 37258 512464 37494
rect 512144 30494 512464 37258
rect 512144 30258 512186 30494
rect 512422 30258 512464 30494
rect 512144 23494 512464 30258
rect 512144 23258 512186 23494
rect 512422 23258 512464 23494
rect 512144 16494 512464 23258
rect 512144 16258 512186 16494
rect 512422 16258 512464 16494
rect 512144 9494 512464 16258
rect 512144 9258 512186 9494
rect 512422 9258 512464 9494
rect 512144 2494 512464 9258
rect 512144 2258 512186 2494
rect 512422 2258 512464 2494
rect 512144 -746 512464 2258
rect 512144 -982 512186 -746
rect 512422 -982 512464 -746
rect 512144 -1066 512464 -982
rect 512144 -1302 512186 -1066
rect 512422 -1302 512464 -1066
rect 512144 -2294 512464 -1302
rect 513876 706198 514196 706230
rect 513876 705962 513918 706198
rect 514154 705962 514196 706198
rect 513876 705878 514196 705962
rect 513876 705642 513918 705878
rect 514154 705642 514196 705878
rect 513876 696561 514196 705642
rect 513876 696325 513918 696561
rect 514154 696325 514196 696561
rect 513876 689561 514196 696325
rect 513876 689325 513918 689561
rect 514154 689325 514196 689561
rect 513876 682561 514196 689325
rect 513876 682325 513918 682561
rect 514154 682325 514196 682561
rect 513876 675561 514196 682325
rect 513876 675325 513918 675561
rect 514154 675325 514196 675561
rect 513876 668561 514196 675325
rect 513876 668325 513918 668561
rect 514154 668325 514196 668561
rect 513876 661561 514196 668325
rect 513876 661325 513918 661561
rect 514154 661325 514196 661561
rect 513876 654561 514196 661325
rect 513876 654325 513918 654561
rect 514154 654325 514196 654561
rect 513876 647561 514196 654325
rect 513876 647325 513918 647561
rect 514154 647325 514196 647561
rect 513876 640561 514196 647325
rect 513876 640325 513918 640561
rect 514154 640325 514196 640561
rect 513876 633561 514196 640325
rect 513876 633325 513918 633561
rect 514154 633325 514196 633561
rect 513876 626561 514196 633325
rect 513876 626325 513918 626561
rect 514154 626325 514196 626561
rect 513876 619561 514196 626325
rect 513876 619325 513918 619561
rect 514154 619325 514196 619561
rect 513876 612561 514196 619325
rect 513876 612325 513918 612561
rect 514154 612325 514196 612561
rect 513876 605561 514196 612325
rect 513876 605325 513918 605561
rect 514154 605325 514196 605561
rect 513876 598561 514196 605325
rect 513876 598325 513918 598561
rect 514154 598325 514196 598561
rect 513876 591561 514196 598325
rect 513876 591325 513918 591561
rect 514154 591325 514196 591561
rect 513876 584561 514196 591325
rect 513876 584325 513918 584561
rect 514154 584325 514196 584561
rect 513876 577561 514196 584325
rect 513876 577325 513918 577561
rect 514154 577325 514196 577561
rect 513876 570561 514196 577325
rect 513876 570325 513918 570561
rect 514154 570325 514196 570561
rect 513876 563561 514196 570325
rect 513876 563325 513918 563561
rect 514154 563325 514196 563561
rect 513876 556561 514196 563325
rect 513876 556325 513918 556561
rect 514154 556325 514196 556561
rect 513876 549561 514196 556325
rect 513876 549325 513918 549561
rect 514154 549325 514196 549561
rect 513876 542561 514196 549325
rect 513876 542325 513918 542561
rect 514154 542325 514196 542561
rect 513876 535561 514196 542325
rect 513876 535325 513918 535561
rect 514154 535325 514196 535561
rect 513876 528561 514196 535325
rect 513876 528325 513918 528561
rect 514154 528325 514196 528561
rect 513876 521561 514196 528325
rect 513876 521325 513918 521561
rect 514154 521325 514196 521561
rect 513876 514561 514196 521325
rect 513876 514325 513918 514561
rect 514154 514325 514196 514561
rect 513876 507561 514196 514325
rect 513876 507325 513918 507561
rect 514154 507325 514196 507561
rect 513876 500561 514196 507325
rect 513876 500325 513918 500561
rect 514154 500325 514196 500561
rect 513876 493561 514196 500325
rect 513876 493325 513918 493561
rect 514154 493325 514196 493561
rect 513876 486561 514196 493325
rect 513876 486325 513918 486561
rect 514154 486325 514196 486561
rect 513876 479561 514196 486325
rect 513876 479325 513918 479561
rect 514154 479325 514196 479561
rect 513876 472561 514196 479325
rect 513876 472325 513918 472561
rect 514154 472325 514196 472561
rect 513876 465561 514196 472325
rect 513876 465325 513918 465561
rect 514154 465325 514196 465561
rect 513876 458561 514196 465325
rect 513876 458325 513918 458561
rect 514154 458325 514196 458561
rect 513876 451561 514196 458325
rect 513876 451325 513918 451561
rect 514154 451325 514196 451561
rect 513876 444561 514196 451325
rect 513876 444325 513918 444561
rect 514154 444325 514196 444561
rect 513876 437561 514196 444325
rect 513876 437325 513918 437561
rect 514154 437325 514196 437561
rect 513876 430561 514196 437325
rect 513876 430325 513918 430561
rect 514154 430325 514196 430561
rect 513876 423561 514196 430325
rect 513876 423325 513918 423561
rect 514154 423325 514196 423561
rect 513876 416561 514196 423325
rect 513876 416325 513918 416561
rect 514154 416325 514196 416561
rect 513876 409561 514196 416325
rect 513876 409325 513918 409561
rect 514154 409325 514196 409561
rect 513876 402561 514196 409325
rect 513876 402325 513918 402561
rect 514154 402325 514196 402561
rect 513876 395561 514196 402325
rect 513876 395325 513918 395561
rect 514154 395325 514196 395561
rect 513876 388561 514196 395325
rect 513876 388325 513918 388561
rect 514154 388325 514196 388561
rect 513876 381561 514196 388325
rect 513876 381325 513918 381561
rect 514154 381325 514196 381561
rect 513876 374561 514196 381325
rect 513876 374325 513918 374561
rect 514154 374325 514196 374561
rect 513876 367561 514196 374325
rect 513876 367325 513918 367561
rect 514154 367325 514196 367561
rect 513876 360561 514196 367325
rect 513876 360325 513918 360561
rect 514154 360325 514196 360561
rect 513876 353561 514196 360325
rect 513876 353325 513918 353561
rect 514154 353325 514196 353561
rect 513876 346561 514196 353325
rect 513876 346325 513918 346561
rect 514154 346325 514196 346561
rect 513876 339561 514196 346325
rect 513876 339325 513918 339561
rect 514154 339325 514196 339561
rect 513876 332561 514196 339325
rect 513876 332325 513918 332561
rect 514154 332325 514196 332561
rect 513876 325561 514196 332325
rect 513876 325325 513918 325561
rect 514154 325325 514196 325561
rect 513876 318561 514196 325325
rect 513876 318325 513918 318561
rect 514154 318325 514196 318561
rect 513876 311561 514196 318325
rect 513876 311325 513918 311561
rect 514154 311325 514196 311561
rect 513876 304561 514196 311325
rect 513876 304325 513918 304561
rect 514154 304325 514196 304561
rect 513876 297561 514196 304325
rect 513876 297325 513918 297561
rect 514154 297325 514196 297561
rect 513876 290561 514196 297325
rect 513876 290325 513918 290561
rect 514154 290325 514196 290561
rect 513876 283561 514196 290325
rect 513876 283325 513918 283561
rect 514154 283325 514196 283561
rect 513876 276561 514196 283325
rect 513876 276325 513918 276561
rect 514154 276325 514196 276561
rect 513876 269561 514196 276325
rect 513876 269325 513918 269561
rect 514154 269325 514196 269561
rect 513876 262561 514196 269325
rect 513876 262325 513918 262561
rect 514154 262325 514196 262561
rect 513876 255561 514196 262325
rect 513876 255325 513918 255561
rect 514154 255325 514196 255561
rect 513876 248561 514196 255325
rect 513876 248325 513918 248561
rect 514154 248325 514196 248561
rect 513876 241561 514196 248325
rect 513876 241325 513918 241561
rect 514154 241325 514196 241561
rect 513876 234561 514196 241325
rect 513876 234325 513918 234561
rect 514154 234325 514196 234561
rect 513876 227561 514196 234325
rect 513876 227325 513918 227561
rect 514154 227325 514196 227561
rect 513876 220561 514196 227325
rect 513876 220325 513918 220561
rect 514154 220325 514196 220561
rect 513876 213561 514196 220325
rect 513876 213325 513918 213561
rect 514154 213325 514196 213561
rect 513876 206561 514196 213325
rect 513876 206325 513918 206561
rect 514154 206325 514196 206561
rect 513876 199561 514196 206325
rect 513876 199325 513918 199561
rect 514154 199325 514196 199561
rect 513876 192561 514196 199325
rect 513876 192325 513918 192561
rect 514154 192325 514196 192561
rect 513876 185561 514196 192325
rect 513876 185325 513918 185561
rect 514154 185325 514196 185561
rect 513876 178561 514196 185325
rect 513876 178325 513918 178561
rect 514154 178325 514196 178561
rect 513876 171561 514196 178325
rect 513876 171325 513918 171561
rect 514154 171325 514196 171561
rect 513876 164561 514196 171325
rect 513876 164325 513918 164561
rect 514154 164325 514196 164561
rect 513876 157561 514196 164325
rect 513876 157325 513918 157561
rect 514154 157325 514196 157561
rect 513876 150561 514196 157325
rect 513876 150325 513918 150561
rect 514154 150325 514196 150561
rect 513876 143561 514196 150325
rect 513876 143325 513918 143561
rect 514154 143325 514196 143561
rect 513876 136561 514196 143325
rect 513876 136325 513918 136561
rect 514154 136325 514196 136561
rect 513876 129561 514196 136325
rect 513876 129325 513918 129561
rect 514154 129325 514196 129561
rect 513876 122561 514196 129325
rect 513876 122325 513918 122561
rect 514154 122325 514196 122561
rect 513876 115561 514196 122325
rect 513876 115325 513918 115561
rect 514154 115325 514196 115561
rect 513876 108561 514196 115325
rect 513876 108325 513918 108561
rect 514154 108325 514196 108561
rect 513876 101561 514196 108325
rect 513876 101325 513918 101561
rect 514154 101325 514196 101561
rect 513876 94561 514196 101325
rect 513876 94325 513918 94561
rect 514154 94325 514196 94561
rect 513876 87561 514196 94325
rect 513876 87325 513918 87561
rect 514154 87325 514196 87561
rect 513876 80561 514196 87325
rect 513876 80325 513918 80561
rect 514154 80325 514196 80561
rect 513876 73561 514196 80325
rect 513876 73325 513918 73561
rect 514154 73325 514196 73561
rect 513876 66561 514196 73325
rect 513876 66325 513918 66561
rect 514154 66325 514196 66561
rect 513876 59561 514196 66325
rect 513876 59325 513918 59561
rect 514154 59325 514196 59561
rect 513876 52561 514196 59325
rect 513876 52325 513918 52561
rect 514154 52325 514196 52561
rect 513876 45561 514196 52325
rect 513876 45325 513918 45561
rect 514154 45325 514196 45561
rect 513876 38561 514196 45325
rect 513876 38325 513918 38561
rect 514154 38325 514196 38561
rect 513876 31561 514196 38325
rect 513876 31325 513918 31561
rect 514154 31325 514196 31561
rect 513876 24561 514196 31325
rect 513876 24325 513918 24561
rect 514154 24325 514196 24561
rect 513876 17561 514196 24325
rect 513876 17325 513918 17561
rect 514154 17325 514196 17561
rect 513876 10561 514196 17325
rect 513876 10325 513918 10561
rect 514154 10325 514196 10561
rect 513876 3561 514196 10325
rect 513876 3325 513918 3561
rect 514154 3325 514196 3561
rect 513876 -1706 514196 3325
rect 513876 -1942 513918 -1706
rect 514154 -1942 514196 -1706
rect 513876 -2026 514196 -1942
rect 513876 -2262 513918 -2026
rect 514154 -2262 514196 -2026
rect 513876 -2294 514196 -2262
rect 519144 705238 519464 706230
rect 519144 705002 519186 705238
rect 519422 705002 519464 705238
rect 519144 704918 519464 705002
rect 519144 704682 519186 704918
rect 519422 704682 519464 704918
rect 519144 695494 519464 704682
rect 519144 695258 519186 695494
rect 519422 695258 519464 695494
rect 519144 688494 519464 695258
rect 519144 688258 519186 688494
rect 519422 688258 519464 688494
rect 519144 681494 519464 688258
rect 519144 681258 519186 681494
rect 519422 681258 519464 681494
rect 519144 674494 519464 681258
rect 519144 674258 519186 674494
rect 519422 674258 519464 674494
rect 519144 667494 519464 674258
rect 519144 667258 519186 667494
rect 519422 667258 519464 667494
rect 519144 660494 519464 667258
rect 519144 660258 519186 660494
rect 519422 660258 519464 660494
rect 519144 653494 519464 660258
rect 519144 653258 519186 653494
rect 519422 653258 519464 653494
rect 519144 646494 519464 653258
rect 519144 646258 519186 646494
rect 519422 646258 519464 646494
rect 519144 639494 519464 646258
rect 519144 639258 519186 639494
rect 519422 639258 519464 639494
rect 519144 632494 519464 639258
rect 519144 632258 519186 632494
rect 519422 632258 519464 632494
rect 519144 625494 519464 632258
rect 519144 625258 519186 625494
rect 519422 625258 519464 625494
rect 519144 618494 519464 625258
rect 519144 618258 519186 618494
rect 519422 618258 519464 618494
rect 519144 611494 519464 618258
rect 519144 611258 519186 611494
rect 519422 611258 519464 611494
rect 519144 604494 519464 611258
rect 519144 604258 519186 604494
rect 519422 604258 519464 604494
rect 519144 597494 519464 604258
rect 519144 597258 519186 597494
rect 519422 597258 519464 597494
rect 519144 590494 519464 597258
rect 519144 590258 519186 590494
rect 519422 590258 519464 590494
rect 519144 583494 519464 590258
rect 519144 583258 519186 583494
rect 519422 583258 519464 583494
rect 519144 576494 519464 583258
rect 519144 576258 519186 576494
rect 519422 576258 519464 576494
rect 519144 569494 519464 576258
rect 519144 569258 519186 569494
rect 519422 569258 519464 569494
rect 519144 562494 519464 569258
rect 519144 562258 519186 562494
rect 519422 562258 519464 562494
rect 519144 555494 519464 562258
rect 519144 555258 519186 555494
rect 519422 555258 519464 555494
rect 519144 548494 519464 555258
rect 519144 548258 519186 548494
rect 519422 548258 519464 548494
rect 519144 541494 519464 548258
rect 519144 541258 519186 541494
rect 519422 541258 519464 541494
rect 519144 534494 519464 541258
rect 519144 534258 519186 534494
rect 519422 534258 519464 534494
rect 519144 527494 519464 534258
rect 519144 527258 519186 527494
rect 519422 527258 519464 527494
rect 519144 520494 519464 527258
rect 519144 520258 519186 520494
rect 519422 520258 519464 520494
rect 519144 513494 519464 520258
rect 519144 513258 519186 513494
rect 519422 513258 519464 513494
rect 519144 506494 519464 513258
rect 519144 506258 519186 506494
rect 519422 506258 519464 506494
rect 519144 499494 519464 506258
rect 519144 499258 519186 499494
rect 519422 499258 519464 499494
rect 519144 492494 519464 499258
rect 519144 492258 519186 492494
rect 519422 492258 519464 492494
rect 519144 485494 519464 492258
rect 519144 485258 519186 485494
rect 519422 485258 519464 485494
rect 519144 478494 519464 485258
rect 519144 478258 519186 478494
rect 519422 478258 519464 478494
rect 519144 471494 519464 478258
rect 519144 471258 519186 471494
rect 519422 471258 519464 471494
rect 519144 464494 519464 471258
rect 519144 464258 519186 464494
rect 519422 464258 519464 464494
rect 519144 457494 519464 464258
rect 519144 457258 519186 457494
rect 519422 457258 519464 457494
rect 519144 450494 519464 457258
rect 519144 450258 519186 450494
rect 519422 450258 519464 450494
rect 519144 443494 519464 450258
rect 519144 443258 519186 443494
rect 519422 443258 519464 443494
rect 519144 436494 519464 443258
rect 519144 436258 519186 436494
rect 519422 436258 519464 436494
rect 519144 429494 519464 436258
rect 519144 429258 519186 429494
rect 519422 429258 519464 429494
rect 519144 422494 519464 429258
rect 519144 422258 519186 422494
rect 519422 422258 519464 422494
rect 519144 415494 519464 422258
rect 520876 706198 521196 706230
rect 520876 705962 520918 706198
rect 521154 705962 521196 706198
rect 520876 705878 521196 705962
rect 520876 705642 520918 705878
rect 521154 705642 521196 705878
rect 520876 696561 521196 705642
rect 520876 696325 520918 696561
rect 521154 696325 521196 696561
rect 520876 689561 521196 696325
rect 520876 689325 520918 689561
rect 521154 689325 521196 689561
rect 520876 682561 521196 689325
rect 520876 682325 520918 682561
rect 521154 682325 521196 682561
rect 520876 675561 521196 682325
rect 520876 675325 520918 675561
rect 521154 675325 521196 675561
rect 520876 668561 521196 675325
rect 520876 668325 520918 668561
rect 521154 668325 521196 668561
rect 520876 661561 521196 668325
rect 520876 661325 520918 661561
rect 521154 661325 521196 661561
rect 520876 654561 521196 661325
rect 520876 654325 520918 654561
rect 521154 654325 521196 654561
rect 520876 647561 521196 654325
rect 520876 647325 520918 647561
rect 521154 647325 521196 647561
rect 520876 640561 521196 647325
rect 520876 640325 520918 640561
rect 521154 640325 521196 640561
rect 520876 633561 521196 640325
rect 520876 633325 520918 633561
rect 521154 633325 521196 633561
rect 520876 626561 521196 633325
rect 520876 626325 520918 626561
rect 521154 626325 521196 626561
rect 520876 619561 521196 626325
rect 520876 619325 520918 619561
rect 521154 619325 521196 619561
rect 520876 612561 521196 619325
rect 520876 612325 520918 612561
rect 521154 612325 521196 612561
rect 520876 605561 521196 612325
rect 520876 605325 520918 605561
rect 521154 605325 521196 605561
rect 520876 598561 521196 605325
rect 520876 598325 520918 598561
rect 521154 598325 521196 598561
rect 520876 591561 521196 598325
rect 520876 591325 520918 591561
rect 521154 591325 521196 591561
rect 520876 584561 521196 591325
rect 520876 584325 520918 584561
rect 521154 584325 521196 584561
rect 520876 577561 521196 584325
rect 520876 577325 520918 577561
rect 521154 577325 521196 577561
rect 520876 570561 521196 577325
rect 520876 570325 520918 570561
rect 521154 570325 521196 570561
rect 520876 563561 521196 570325
rect 520876 563325 520918 563561
rect 521154 563325 521196 563561
rect 520876 556561 521196 563325
rect 520876 556325 520918 556561
rect 521154 556325 521196 556561
rect 520876 549561 521196 556325
rect 520876 549325 520918 549561
rect 521154 549325 521196 549561
rect 520876 542561 521196 549325
rect 520876 542325 520918 542561
rect 521154 542325 521196 542561
rect 520876 535561 521196 542325
rect 520876 535325 520918 535561
rect 521154 535325 521196 535561
rect 520876 528561 521196 535325
rect 520876 528325 520918 528561
rect 521154 528325 521196 528561
rect 520876 521561 521196 528325
rect 520876 521325 520918 521561
rect 521154 521325 521196 521561
rect 520876 514561 521196 521325
rect 520876 514325 520918 514561
rect 521154 514325 521196 514561
rect 520876 507561 521196 514325
rect 520876 507325 520918 507561
rect 521154 507325 521196 507561
rect 520876 500561 521196 507325
rect 520876 500325 520918 500561
rect 521154 500325 521196 500561
rect 520876 493561 521196 500325
rect 520876 493325 520918 493561
rect 521154 493325 521196 493561
rect 520876 486561 521196 493325
rect 520876 486325 520918 486561
rect 521154 486325 521196 486561
rect 520876 479561 521196 486325
rect 520876 479325 520918 479561
rect 521154 479325 521196 479561
rect 520876 472561 521196 479325
rect 520876 472325 520918 472561
rect 521154 472325 521196 472561
rect 520876 465561 521196 472325
rect 520876 465325 520918 465561
rect 521154 465325 521196 465561
rect 520876 458561 521196 465325
rect 520876 458325 520918 458561
rect 521154 458325 521196 458561
rect 520876 451561 521196 458325
rect 520876 451325 520918 451561
rect 521154 451325 521196 451561
rect 520876 444561 521196 451325
rect 520876 444325 520918 444561
rect 521154 444325 521196 444561
rect 520876 437561 521196 444325
rect 520876 437325 520918 437561
rect 521154 437325 521196 437561
rect 520876 430561 521196 437325
rect 520876 430325 520918 430561
rect 521154 430325 521196 430561
rect 520876 423561 521196 430325
rect 520876 423325 520918 423561
rect 521154 423325 521196 423561
rect 520876 421752 521196 423325
rect 526144 705238 526464 706230
rect 526144 705002 526186 705238
rect 526422 705002 526464 705238
rect 526144 704918 526464 705002
rect 526144 704682 526186 704918
rect 526422 704682 526464 704918
rect 526144 695494 526464 704682
rect 526144 695258 526186 695494
rect 526422 695258 526464 695494
rect 526144 688494 526464 695258
rect 526144 688258 526186 688494
rect 526422 688258 526464 688494
rect 526144 681494 526464 688258
rect 526144 681258 526186 681494
rect 526422 681258 526464 681494
rect 526144 674494 526464 681258
rect 526144 674258 526186 674494
rect 526422 674258 526464 674494
rect 526144 667494 526464 674258
rect 526144 667258 526186 667494
rect 526422 667258 526464 667494
rect 526144 660494 526464 667258
rect 526144 660258 526186 660494
rect 526422 660258 526464 660494
rect 526144 653494 526464 660258
rect 526144 653258 526186 653494
rect 526422 653258 526464 653494
rect 526144 646494 526464 653258
rect 526144 646258 526186 646494
rect 526422 646258 526464 646494
rect 526144 639494 526464 646258
rect 526144 639258 526186 639494
rect 526422 639258 526464 639494
rect 526144 632494 526464 639258
rect 526144 632258 526186 632494
rect 526422 632258 526464 632494
rect 526144 625494 526464 632258
rect 526144 625258 526186 625494
rect 526422 625258 526464 625494
rect 526144 618494 526464 625258
rect 526144 618258 526186 618494
rect 526422 618258 526464 618494
rect 526144 611494 526464 618258
rect 526144 611258 526186 611494
rect 526422 611258 526464 611494
rect 526144 604494 526464 611258
rect 526144 604258 526186 604494
rect 526422 604258 526464 604494
rect 526144 597494 526464 604258
rect 526144 597258 526186 597494
rect 526422 597258 526464 597494
rect 526144 590494 526464 597258
rect 526144 590258 526186 590494
rect 526422 590258 526464 590494
rect 526144 583494 526464 590258
rect 526144 583258 526186 583494
rect 526422 583258 526464 583494
rect 526144 576494 526464 583258
rect 526144 576258 526186 576494
rect 526422 576258 526464 576494
rect 526144 569494 526464 576258
rect 526144 569258 526186 569494
rect 526422 569258 526464 569494
rect 526144 562494 526464 569258
rect 526144 562258 526186 562494
rect 526422 562258 526464 562494
rect 526144 555494 526464 562258
rect 526144 555258 526186 555494
rect 526422 555258 526464 555494
rect 526144 548494 526464 555258
rect 526144 548258 526186 548494
rect 526422 548258 526464 548494
rect 526144 541494 526464 548258
rect 526144 541258 526186 541494
rect 526422 541258 526464 541494
rect 526144 534494 526464 541258
rect 526144 534258 526186 534494
rect 526422 534258 526464 534494
rect 526144 527494 526464 534258
rect 526144 527258 526186 527494
rect 526422 527258 526464 527494
rect 526144 520494 526464 527258
rect 526144 520258 526186 520494
rect 526422 520258 526464 520494
rect 526144 513494 526464 520258
rect 526144 513258 526186 513494
rect 526422 513258 526464 513494
rect 526144 506494 526464 513258
rect 526144 506258 526186 506494
rect 526422 506258 526464 506494
rect 526144 499494 526464 506258
rect 526144 499258 526186 499494
rect 526422 499258 526464 499494
rect 526144 492494 526464 499258
rect 526144 492258 526186 492494
rect 526422 492258 526464 492494
rect 526144 485494 526464 492258
rect 526144 485258 526186 485494
rect 526422 485258 526464 485494
rect 526144 478494 526464 485258
rect 526144 478258 526186 478494
rect 526422 478258 526464 478494
rect 526144 471494 526464 478258
rect 526144 471258 526186 471494
rect 526422 471258 526464 471494
rect 526144 464494 526464 471258
rect 526144 464258 526186 464494
rect 526422 464258 526464 464494
rect 526144 457494 526464 464258
rect 526144 457258 526186 457494
rect 526422 457258 526464 457494
rect 526144 450494 526464 457258
rect 526144 450258 526186 450494
rect 526422 450258 526464 450494
rect 526144 443494 526464 450258
rect 526144 443258 526186 443494
rect 526422 443258 526464 443494
rect 526144 436494 526464 443258
rect 526144 436258 526186 436494
rect 526422 436258 526464 436494
rect 526144 429494 526464 436258
rect 526144 429258 526186 429494
rect 526422 429258 526464 429494
rect 526144 422494 526464 429258
rect 526144 422258 526186 422494
rect 526422 422258 526464 422494
rect 526144 421752 526464 422258
rect 527876 706198 528196 706230
rect 527876 705962 527918 706198
rect 528154 705962 528196 706198
rect 527876 705878 528196 705962
rect 527876 705642 527918 705878
rect 528154 705642 528196 705878
rect 527876 696561 528196 705642
rect 527876 696325 527918 696561
rect 528154 696325 528196 696561
rect 527876 689561 528196 696325
rect 527876 689325 527918 689561
rect 528154 689325 528196 689561
rect 527876 682561 528196 689325
rect 527876 682325 527918 682561
rect 528154 682325 528196 682561
rect 527876 675561 528196 682325
rect 527876 675325 527918 675561
rect 528154 675325 528196 675561
rect 527876 668561 528196 675325
rect 527876 668325 527918 668561
rect 528154 668325 528196 668561
rect 527876 661561 528196 668325
rect 527876 661325 527918 661561
rect 528154 661325 528196 661561
rect 527876 654561 528196 661325
rect 527876 654325 527918 654561
rect 528154 654325 528196 654561
rect 527876 647561 528196 654325
rect 527876 647325 527918 647561
rect 528154 647325 528196 647561
rect 527876 640561 528196 647325
rect 527876 640325 527918 640561
rect 528154 640325 528196 640561
rect 527876 633561 528196 640325
rect 527876 633325 527918 633561
rect 528154 633325 528196 633561
rect 527876 626561 528196 633325
rect 527876 626325 527918 626561
rect 528154 626325 528196 626561
rect 527876 619561 528196 626325
rect 527876 619325 527918 619561
rect 528154 619325 528196 619561
rect 527876 612561 528196 619325
rect 527876 612325 527918 612561
rect 528154 612325 528196 612561
rect 527876 605561 528196 612325
rect 527876 605325 527918 605561
rect 528154 605325 528196 605561
rect 527876 598561 528196 605325
rect 527876 598325 527918 598561
rect 528154 598325 528196 598561
rect 527876 591561 528196 598325
rect 527876 591325 527918 591561
rect 528154 591325 528196 591561
rect 527876 584561 528196 591325
rect 527876 584325 527918 584561
rect 528154 584325 528196 584561
rect 527876 577561 528196 584325
rect 527876 577325 527918 577561
rect 528154 577325 528196 577561
rect 527876 570561 528196 577325
rect 527876 570325 527918 570561
rect 528154 570325 528196 570561
rect 527876 563561 528196 570325
rect 527876 563325 527918 563561
rect 528154 563325 528196 563561
rect 527876 556561 528196 563325
rect 527876 556325 527918 556561
rect 528154 556325 528196 556561
rect 527876 549561 528196 556325
rect 527876 549325 527918 549561
rect 528154 549325 528196 549561
rect 527876 542561 528196 549325
rect 527876 542325 527918 542561
rect 528154 542325 528196 542561
rect 527876 535561 528196 542325
rect 527876 535325 527918 535561
rect 528154 535325 528196 535561
rect 527876 528561 528196 535325
rect 527876 528325 527918 528561
rect 528154 528325 528196 528561
rect 527876 521561 528196 528325
rect 527876 521325 527918 521561
rect 528154 521325 528196 521561
rect 527876 514561 528196 521325
rect 527876 514325 527918 514561
rect 528154 514325 528196 514561
rect 527876 507561 528196 514325
rect 527876 507325 527918 507561
rect 528154 507325 528196 507561
rect 527876 500561 528196 507325
rect 527876 500325 527918 500561
rect 528154 500325 528196 500561
rect 527876 493561 528196 500325
rect 527876 493325 527918 493561
rect 528154 493325 528196 493561
rect 527876 486561 528196 493325
rect 527876 486325 527918 486561
rect 528154 486325 528196 486561
rect 527876 479561 528196 486325
rect 527876 479325 527918 479561
rect 528154 479325 528196 479561
rect 527876 472561 528196 479325
rect 527876 472325 527918 472561
rect 528154 472325 528196 472561
rect 527876 465561 528196 472325
rect 527876 465325 527918 465561
rect 528154 465325 528196 465561
rect 527876 458561 528196 465325
rect 527876 458325 527918 458561
rect 528154 458325 528196 458561
rect 527876 451561 528196 458325
rect 527876 451325 527918 451561
rect 528154 451325 528196 451561
rect 527876 444561 528196 451325
rect 527876 444325 527918 444561
rect 528154 444325 528196 444561
rect 527876 437561 528196 444325
rect 527876 437325 527918 437561
rect 528154 437325 528196 437561
rect 527876 430561 528196 437325
rect 527876 430325 527918 430561
rect 528154 430325 528196 430561
rect 527876 423561 528196 430325
rect 527876 423325 527918 423561
rect 528154 423325 528196 423561
rect 527876 416561 528196 423325
rect 520876 416325 520918 416561
rect 521154 416325 521196 416561
rect 522808 416325 522850 416561
rect 523086 416325 523128 416561
rect 524740 416325 524782 416561
rect 525018 416325 525060 416561
rect 526672 416325 526714 416561
rect 526950 416325 526992 416561
rect 527876 416325 527918 416561
rect 528154 416325 528196 416561
rect 519144 415258 519186 415494
rect 519422 415258 519464 415494
rect 519910 415258 519952 415494
rect 520188 415258 520230 415494
rect 521842 415258 521884 415494
rect 522120 415258 522162 415494
rect 523774 415258 523816 415494
rect 524052 415258 524094 415494
rect 525706 415258 525748 415494
rect 525984 415258 526026 415494
rect 519144 408494 519464 415258
rect 527876 409561 528196 416325
rect 520876 409325 520918 409561
rect 521154 409325 521196 409561
rect 522808 409325 522850 409561
rect 523086 409325 523128 409561
rect 524740 409325 524782 409561
rect 525018 409325 525060 409561
rect 526672 409325 526714 409561
rect 526950 409325 526992 409561
rect 527876 409325 527918 409561
rect 528154 409325 528196 409561
rect 519144 408258 519186 408494
rect 519422 408258 519464 408494
rect 519910 408258 519952 408494
rect 520188 408258 520230 408494
rect 521842 408258 521884 408494
rect 522120 408258 522162 408494
rect 523774 408258 523816 408494
rect 524052 408258 524094 408494
rect 525706 408258 525748 408494
rect 525984 408258 526026 408494
rect 519144 401494 519464 408258
rect 527876 402561 528196 409325
rect 520876 402325 520918 402561
rect 521154 402325 521196 402561
rect 522808 402325 522850 402561
rect 523086 402325 523128 402561
rect 524740 402325 524782 402561
rect 525018 402325 525060 402561
rect 526672 402325 526714 402561
rect 526950 402325 526992 402561
rect 527876 402325 527918 402561
rect 528154 402325 528196 402561
rect 519144 401258 519186 401494
rect 519422 401258 519464 401494
rect 519144 394494 519464 401258
rect 519144 394258 519186 394494
rect 519422 394258 519464 394494
rect 519144 387494 519464 394258
rect 519144 387258 519186 387494
rect 519422 387258 519464 387494
rect 519144 380494 519464 387258
rect 520876 395561 521196 400008
rect 520876 395325 520918 395561
rect 521154 395325 521196 395561
rect 520876 388561 521196 395325
rect 520876 388325 520918 388561
rect 521154 388325 521196 388561
rect 520876 381752 521196 388325
rect 526144 394494 526464 400008
rect 526144 394258 526186 394494
rect 526422 394258 526464 394494
rect 526144 387494 526464 394258
rect 526144 387258 526186 387494
rect 526422 387258 526464 387494
rect 526144 381752 526464 387258
rect 527876 395561 528196 402325
rect 527876 395325 527918 395561
rect 528154 395325 528196 395561
rect 527876 388561 528196 395325
rect 527876 388325 527918 388561
rect 528154 388325 528196 388561
rect 519144 380258 519186 380494
rect 519422 380258 519464 380494
rect 519144 373494 519464 380258
rect 527876 381561 528196 388325
rect 527876 381325 527918 381561
rect 528154 381325 528196 381561
rect 527876 374561 528196 381325
rect 520876 374325 520918 374561
rect 521154 374325 521196 374561
rect 522808 374325 522850 374561
rect 523086 374325 523128 374561
rect 524740 374325 524782 374561
rect 525018 374325 525060 374561
rect 526672 374325 526714 374561
rect 526950 374325 526992 374561
rect 527876 374325 527918 374561
rect 528154 374325 528196 374561
rect 519144 373258 519186 373494
rect 519422 373258 519464 373494
rect 519910 373258 519952 373494
rect 520188 373258 520230 373494
rect 521842 373258 521884 373494
rect 522120 373258 522162 373494
rect 523774 373258 523816 373494
rect 524052 373258 524094 373494
rect 525706 373258 525748 373494
rect 525984 373258 526026 373494
rect 519144 366494 519464 373258
rect 527876 367561 528196 374325
rect 520876 367325 520918 367561
rect 521154 367325 521196 367561
rect 522808 367325 522850 367561
rect 523086 367325 523128 367561
rect 524740 367325 524782 367561
rect 525018 367325 525060 367561
rect 526672 367325 526714 367561
rect 526950 367325 526992 367561
rect 527876 367325 527918 367561
rect 528154 367325 528196 367561
rect 519144 366258 519186 366494
rect 519422 366258 519464 366494
rect 519910 366258 519952 366494
rect 520188 366258 520230 366494
rect 521842 366258 521884 366494
rect 522120 366258 522162 366494
rect 523774 366258 523816 366494
rect 524052 366258 524094 366494
rect 525706 366258 525748 366494
rect 525984 366258 526026 366494
rect 519144 359494 519464 366258
rect 527876 360561 528196 367325
rect 527876 360325 527918 360561
rect 528154 360325 528196 360561
rect 519144 359258 519186 359494
rect 519422 359258 519464 359494
rect 519144 352494 519464 359258
rect 519144 352258 519186 352494
rect 519422 352258 519464 352494
rect 519144 345494 519464 352258
rect 519144 345258 519186 345494
rect 519422 345258 519464 345494
rect 519144 338494 519464 345258
rect 520876 353561 521196 360008
rect 520876 353325 520918 353561
rect 521154 353325 521196 353561
rect 520876 346561 521196 353325
rect 520876 346325 520918 346561
rect 521154 346325 521196 346561
rect 520876 341752 521196 346325
rect 526144 359494 526464 360008
rect 526144 359258 526186 359494
rect 526422 359258 526464 359494
rect 526144 352494 526464 359258
rect 526144 352258 526186 352494
rect 526422 352258 526464 352494
rect 526144 345494 526464 352258
rect 526144 345258 526186 345494
rect 526422 345258 526464 345494
rect 526144 341752 526464 345258
rect 527876 353561 528196 360325
rect 527876 353325 527918 353561
rect 528154 353325 528196 353561
rect 527876 346561 528196 353325
rect 527876 346325 527918 346561
rect 528154 346325 528196 346561
rect 527876 339561 528196 346325
rect 520876 339325 520918 339561
rect 521154 339325 521196 339561
rect 522808 339325 522850 339561
rect 523086 339325 523128 339561
rect 524740 339325 524782 339561
rect 525018 339325 525060 339561
rect 526672 339325 526714 339561
rect 526950 339325 526992 339561
rect 527876 339325 527918 339561
rect 528154 339325 528196 339561
rect 519144 338258 519186 338494
rect 519422 338258 519464 338494
rect 519910 338258 519952 338494
rect 520188 338258 520230 338494
rect 521842 338258 521884 338494
rect 522120 338258 522162 338494
rect 523774 338258 523816 338494
rect 524052 338258 524094 338494
rect 525706 338258 525748 338494
rect 525984 338258 526026 338494
rect 519144 331494 519464 338258
rect 527876 332561 528196 339325
rect 520876 332325 520918 332561
rect 521154 332325 521196 332561
rect 522808 332325 522850 332561
rect 523086 332325 523128 332561
rect 524740 332325 524782 332561
rect 525018 332325 525060 332561
rect 526672 332325 526714 332561
rect 526950 332325 526992 332561
rect 527876 332325 527918 332561
rect 528154 332325 528196 332561
rect 519144 331258 519186 331494
rect 519422 331258 519464 331494
rect 519910 331258 519952 331494
rect 520188 331258 520230 331494
rect 521842 331258 521884 331494
rect 522120 331258 522162 331494
rect 523774 331258 523816 331494
rect 524052 331258 524094 331494
rect 525706 331258 525748 331494
rect 525984 331258 526026 331494
rect 519144 324494 519464 331258
rect 527876 325561 528196 332325
rect 520876 325325 520918 325561
rect 521154 325325 521196 325561
rect 522808 325325 522850 325561
rect 523086 325325 523128 325561
rect 524740 325325 524782 325561
rect 525018 325325 525060 325561
rect 526672 325325 526714 325561
rect 526950 325325 526992 325561
rect 527876 325325 527918 325561
rect 528154 325325 528196 325561
rect 519144 324258 519186 324494
rect 519422 324258 519464 324494
rect 519910 324258 519952 324494
rect 520188 324258 520230 324494
rect 521842 324258 521884 324494
rect 522120 324258 522162 324494
rect 523774 324258 523816 324494
rect 524052 324258 524094 324494
rect 525706 324258 525748 324494
rect 525984 324258 526026 324494
rect 519144 317494 519464 324258
rect 519144 317258 519186 317494
rect 519422 317258 519464 317494
rect 519144 310494 519464 317258
rect 519144 310258 519186 310494
rect 519422 310258 519464 310494
rect 519144 303494 519464 310258
rect 519144 303258 519186 303494
rect 519422 303258 519464 303494
rect 519144 296494 519464 303258
rect 520876 318561 521196 320008
rect 520876 318325 520918 318561
rect 521154 318325 521196 318561
rect 520876 311561 521196 318325
rect 520876 311325 520918 311561
rect 521154 311325 521196 311561
rect 520876 304561 521196 311325
rect 520876 304325 520918 304561
rect 521154 304325 521196 304561
rect 520876 301752 521196 304325
rect 526144 317494 526464 320008
rect 526144 317258 526186 317494
rect 526422 317258 526464 317494
rect 526144 310494 526464 317258
rect 526144 310258 526186 310494
rect 526422 310258 526464 310494
rect 526144 303494 526464 310258
rect 526144 303258 526186 303494
rect 526422 303258 526464 303494
rect 526144 301752 526464 303258
rect 527876 318561 528196 325325
rect 527876 318325 527918 318561
rect 528154 318325 528196 318561
rect 527876 311561 528196 318325
rect 527876 311325 527918 311561
rect 528154 311325 528196 311561
rect 527876 304561 528196 311325
rect 527876 304325 527918 304561
rect 528154 304325 528196 304561
rect 527876 297561 528196 304325
rect 520876 297325 520918 297561
rect 521154 297325 521196 297561
rect 522808 297325 522850 297561
rect 523086 297325 523128 297561
rect 524740 297325 524782 297561
rect 525018 297325 525060 297561
rect 526672 297325 526714 297561
rect 526950 297325 526992 297561
rect 527876 297325 527918 297561
rect 528154 297325 528196 297561
rect 519144 296258 519186 296494
rect 519422 296258 519464 296494
rect 519910 296258 519952 296494
rect 520188 296258 520230 296494
rect 521842 296258 521884 296494
rect 522120 296258 522162 296494
rect 523774 296258 523816 296494
rect 524052 296258 524094 296494
rect 525706 296258 525748 296494
rect 525984 296258 526026 296494
rect 519144 289494 519464 296258
rect 527876 290561 528196 297325
rect 520876 290325 520918 290561
rect 521154 290325 521196 290561
rect 522808 290325 522850 290561
rect 523086 290325 523128 290561
rect 524740 290325 524782 290561
rect 525018 290325 525060 290561
rect 526672 290325 526714 290561
rect 526950 290325 526992 290561
rect 527876 290325 527918 290561
rect 528154 290325 528196 290561
rect 519144 289258 519186 289494
rect 519422 289258 519464 289494
rect 519910 289258 519952 289494
rect 520188 289258 520230 289494
rect 521842 289258 521884 289494
rect 522120 289258 522162 289494
rect 523774 289258 523816 289494
rect 524052 289258 524094 289494
rect 525706 289258 525748 289494
rect 525984 289258 526026 289494
rect 519144 282494 519464 289258
rect 527876 283561 528196 290325
rect 520876 283325 520918 283561
rect 521154 283325 521196 283561
rect 522808 283325 522850 283561
rect 523086 283325 523128 283561
rect 524740 283325 524782 283561
rect 525018 283325 525060 283561
rect 526672 283325 526714 283561
rect 526950 283325 526992 283561
rect 527876 283325 527918 283561
rect 528154 283325 528196 283561
rect 519144 282258 519186 282494
rect 519422 282258 519464 282494
rect 519910 282258 519952 282494
rect 520188 282258 520230 282494
rect 521842 282258 521884 282494
rect 522120 282258 522162 282494
rect 523774 282258 523816 282494
rect 524052 282258 524094 282494
rect 525706 282258 525748 282494
rect 525984 282258 526026 282494
rect 519144 275494 519464 282258
rect 519144 275258 519186 275494
rect 519422 275258 519464 275494
rect 519144 268494 519464 275258
rect 519144 268258 519186 268494
rect 519422 268258 519464 268494
rect 519144 261494 519464 268258
rect 520876 276561 521196 280008
rect 520876 276325 520918 276561
rect 521154 276325 521196 276561
rect 520876 269561 521196 276325
rect 520876 269325 520918 269561
rect 521154 269325 521196 269561
rect 520876 262561 521196 269325
rect 520876 262325 520918 262561
rect 521154 262325 521196 262561
rect 520876 261752 521196 262325
rect 526144 275494 526464 280008
rect 526144 275258 526186 275494
rect 526422 275258 526464 275494
rect 526144 268494 526464 275258
rect 526144 268258 526186 268494
rect 526422 268258 526464 268494
rect 526144 261752 526464 268258
rect 527876 276561 528196 283325
rect 527876 276325 527918 276561
rect 528154 276325 528196 276561
rect 527876 269561 528196 276325
rect 527876 269325 527918 269561
rect 528154 269325 528196 269561
rect 527876 262561 528196 269325
rect 527876 262325 527918 262561
rect 528154 262325 528196 262561
rect 519144 261258 519186 261494
rect 519422 261258 519464 261494
rect 519144 254494 519464 261258
rect 527876 255561 528196 262325
rect 520876 255325 520918 255561
rect 521154 255325 521196 255561
rect 522808 255325 522850 255561
rect 523086 255325 523128 255561
rect 524740 255325 524782 255561
rect 525018 255325 525060 255561
rect 526672 255325 526714 255561
rect 526950 255325 526992 255561
rect 527876 255325 527918 255561
rect 528154 255325 528196 255561
rect 519144 254258 519186 254494
rect 519422 254258 519464 254494
rect 519910 254258 519952 254494
rect 520188 254258 520230 254494
rect 521842 254258 521884 254494
rect 522120 254258 522162 254494
rect 523774 254258 523816 254494
rect 524052 254258 524094 254494
rect 525706 254258 525748 254494
rect 525984 254258 526026 254494
rect 519144 247494 519464 254258
rect 527876 248561 528196 255325
rect 520876 248325 520918 248561
rect 521154 248325 521196 248561
rect 522808 248325 522850 248561
rect 523086 248325 523128 248561
rect 524740 248325 524782 248561
rect 525018 248325 525060 248561
rect 526672 248325 526714 248561
rect 526950 248325 526992 248561
rect 527876 248325 527918 248561
rect 528154 248325 528196 248561
rect 519144 247258 519186 247494
rect 519422 247258 519464 247494
rect 519910 247258 519952 247494
rect 520188 247258 520230 247494
rect 521842 247258 521884 247494
rect 522120 247258 522162 247494
rect 523774 247258 523816 247494
rect 524052 247258 524094 247494
rect 525706 247258 525748 247494
rect 525984 247258 526026 247494
rect 519144 240494 519464 247258
rect 519144 240258 519186 240494
rect 519422 240258 519464 240494
rect 519144 233494 519464 240258
rect 527876 241561 528196 248325
rect 527876 241325 527918 241561
rect 528154 241325 528196 241561
rect 519144 233258 519186 233494
rect 519422 233258 519464 233494
rect 519144 226494 519464 233258
rect 519144 226258 519186 226494
rect 519422 226258 519464 226494
rect 519144 219494 519464 226258
rect 519144 219258 519186 219494
rect 519422 219258 519464 219494
rect 519144 212494 519464 219258
rect 519144 212258 519186 212494
rect 519422 212258 519464 212494
rect 519144 205494 519464 212258
rect 519144 205258 519186 205494
rect 519422 205258 519464 205494
rect 519144 198494 519464 205258
rect 519144 198258 519186 198494
rect 519422 198258 519464 198494
rect 519144 191494 519464 198258
rect 519144 191258 519186 191494
rect 519422 191258 519464 191494
rect 519144 184494 519464 191258
rect 519144 184258 519186 184494
rect 519422 184258 519464 184494
rect 519144 177494 519464 184258
rect 519144 177258 519186 177494
rect 519422 177258 519464 177494
rect 519144 170494 519464 177258
rect 519144 170258 519186 170494
rect 519422 170258 519464 170494
rect 519144 163494 519464 170258
rect 519144 163258 519186 163494
rect 519422 163258 519464 163494
rect 519144 156494 519464 163258
rect 519144 156258 519186 156494
rect 519422 156258 519464 156494
rect 519144 149494 519464 156258
rect 519144 149258 519186 149494
rect 519422 149258 519464 149494
rect 519144 142494 519464 149258
rect 519144 142258 519186 142494
rect 519422 142258 519464 142494
rect 519144 135494 519464 142258
rect 519144 135258 519186 135494
rect 519422 135258 519464 135494
rect 519144 128494 519464 135258
rect 519144 128258 519186 128494
rect 519422 128258 519464 128494
rect 519144 121494 519464 128258
rect 519144 121258 519186 121494
rect 519422 121258 519464 121494
rect 519144 114494 519464 121258
rect 519144 114258 519186 114494
rect 519422 114258 519464 114494
rect 519144 107494 519464 114258
rect 519144 107258 519186 107494
rect 519422 107258 519464 107494
rect 519144 100494 519464 107258
rect 519144 100258 519186 100494
rect 519422 100258 519464 100494
rect 519144 93494 519464 100258
rect 519144 93258 519186 93494
rect 519422 93258 519464 93494
rect 519144 86494 519464 93258
rect 519144 86258 519186 86494
rect 519422 86258 519464 86494
rect 519144 79494 519464 86258
rect 519144 79258 519186 79494
rect 519422 79258 519464 79494
rect 519144 72494 519464 79258
rect 519144 72258 519186 72494
rect 519422 72258 519464 72494
rect 519144 65494 519464 72258
rect 519144 65258 519186 65494
rect 519422 65258 519464 65494
rect 519144 58494 519464 65258
rect 519144 58258 519186 58494
rect 519422 58258 519464 58494
rect 519144 51494 519464 58258
rect 519144 51258 519186 51494
rect 519422 51258 519464 51494
rect 519144 44494 519464 51258
rect 519144 44258 519186 44494
rect 519422 44258 519464 44494
rect 519144 37494 519464 44258
rect 519144 37258 519186 37494
rect 519422 37258 519464 37494
rect 519144 30494 519464 37258
rect 519144 30258 519186 30494
rect 519422 30258 519464 30494
rect 519144 23494 519464 30258
rect 519144 23258 519186 23494
rect 519422 23258 519464 23494
rect 519144 16494 519464 23258
rect 519144 16258 519186 16494
rect 519422 16258 519464 16494
rect 519144 9494 519464 16258
rect 519144 9258 519186 9494
rect 519422 9258 519464 9494
rect 519144 2494 519464 9258
rect 519144 2258 519186 2494
rect 519422 2258 519464 2494
rect 519144 -746 519464 2258
rect 519144 -982 519186 -746
rect 519422 -982 519464 -746
rect 519144 -1066 519464 -982
rect 519144 -1302 519186 -1066
rect 519422 -1302 519464 -1066
rect 519144 -2294 519464 -1302
rect 520876 234561 521196 240008
rect 520876 234325 520918 234561
rect 521154 234325 521196 234561
rect 520876 227561 521196 234325
rect 520876 227325 520918 227561
rect 521154 227325 521196 227561
rect 520876 220561 521196 227325
rect 520876 220325 520918 220561
rect 521154 220325 521196 220561
rect 520876 213561 521196 220325
rect 520876 213325 520918 213561
rect 521154 213325 521196 213561
rect 520876 206561 521196 213325
rect 520876 206325 520918 206561
rect 521154 206325 521196 206561
rect 520876 199561 521196 206325
rect 520876 199325 520918 199561
rect 521154 199325 521196 199561
rect 520876 192561 521196 199325
rect 520876 192325 520918 192561
rect 521154 192325 521196 192561
rect 520876 185561 521196 192325
rect 520876 185325 520918 185561
rect 521154 185325 521196 185561
rect 520876 178561 521196 185325
rect 520876 178325 520918 178561
rect 521154 178325 521196 178561
rect 520876 171561 521196 178325
rect 520876 171325 520918 171561
rect 521154 171325 521196 171561
rect 520876 164561 521196 171325
rect 520876 164325 520918 164561
rect 521154 164325 521196 164561
rect 520876 157561 521196 164325
rect 520876 157325 520918 157561
rect 521154 157325 521196 157561
rect 520876 150561 521196 157325
rect 520876 150325 520918 150561
rect 521154 150325 521196 150561
rect 520876 143561 521196 150325
rect 520876 143325 520918 143561
rect 521154 143325 521196 143561
rect 520876 136561 521196 143325
rect 520876 136325 520918 136561
rect 521154 136325 521196 136561
rect 520876 129561 521196 136325
rect 520876 129325 520918 129561
rect 521154 129325 521196 129561
rect 520876 122561 521196 129325
rect 520876 122325 520918 122561
rect 521154 122325 521196 122561
rect 520876 115561 521196 122325
rect 520876 115325 520918 115561
rect 521154 115325 521196 115561
rect 520876 108561 521196 115325
rect 520876 108325 520918 108561
rect 521154 108325 521196 108561
rect 520876 101561 521196 108325
rect 520876 101325 520918 101561
rect 521154 101325 521196 101561
rect 520876 94561 521196 101325
rect 520876 94325 520918 94561
rect 521154 94325 521196 94561
rect 520876 87561 521196 94325
rect 520876 87325 520918 87561
rect 521154 87325 521196 87561
rect 520876 80561 521196 87325
rect 520876 80325 520918 80561
rect 521154 80325 521196 80561
rect 520876 73561 521196 80325
rect 520876 73325 520918 73561
rect 521154 73325 521196 73561
rect 520876 66561 521196 73325
rect 520876 66325 520918 66561
rect 521154 66325 521196 66561
rect 520876 59561 521196 66325
rect 520876 59325 520918 59561
rect 521154 59325 521196 59561
rect 520876 52561 521196 59325
rect 520876 52325 520918 52561
rect 521154 52325 521196 52561
rect 520876 45561 521196 52325
rect 520876 45325 520918 45561
rect 521154 45325 521196 45561
rect 520876 38561 521196 45325
rect 520876 38325 520918 38561
rect 521154 38325 521196 38561
rect 520876 31561 521196 38325
rect 520876 31325 520918 31561
rect 521154 31325 521196 31561
rect 520876 24561 521196 31325
rect 520876 24325 520918 24561
rect 521154 24325 521196 24561
rect 520876 17561 521196 24325
rect 520876 17325 520918 17561
rect 521154 17325 521196 17561
rect 520876 10561 521196 17325
rect 520876 10325 520918 10561
rect 521154 10325 521196 10561
rect 520876 3561 521196 10325
rect 520876 3325 520918 3561
rect 521154 3325 521196 3561
rect 520876 -1706 521196 3325
rect 520876 -1942 520918 -1706
rect 521154 -1942 521196 -1706
rect 520876 -2026 521196 -1942
rect 520876 -2262 520918 -2026
rect 521154 -2262 521196 -2026
rect 520876 -2294 521196 -2262
rect 526144 233494 526464 240008
rect 526144 233258 526186 233494
rect 526422 233258 526464 233494
rect 526144 226494 526464 233258
rect 526144 226258 526186 226494
rect 526422 226258 526464 226494
rect 526144 219494 526464 226258
rect 526144 219258 526186 219494
rect 526422 219258 526464 219494
rect 526144 212494 526464 219258
rect 526144 212258 526186 212494
rect 526422 212258 526464 212494
rect 526144 205494 526464 212258
rect 526144 205258 526186 205494
rect 526422 205258 526464 205494
rect 526144 198494 526464 205258
rect 526144 198258 526186 198494
rect 526422 198258 526464 198494
rect 526144 191494 526464 198258
rect 526144 191258 526186 191494
rect 526422 191258 526464 191494
rect 526144 184494 526464 191258
rect 526144 184258 526186 184494
rect 526422 184258 526464 184494
rect 526144 177494 526464 184258
rect 526144 177258 526186 177494
rect 526422 177258 526464 177494
rect 526144 170494 526464 177258
rect 526144 170258 526186 170494
rect 526422 170258 526464 170494
rect 526144 163494 526464 170258
rect 526144 163258 526186 163494
rect 526422 163258 526464 163494
rect 526144 156494 526464 163258
rect 526144 156258 526186 156494
rect 526422 156258 526464 156494
rect 526144 149494 526464 156258
rect 526144 149258 526186 149494
rect 526422 149258 526464 149494
rect 526144 142494 526464 149258
rect 526144 142258 526186 142494
rect 526422 142258 526464 142494
rect 526144 135494 526464 142258
rect 526144 135258 526186 135494
rect 526422 135258 526464 135494
rect 526144 128494 526464 135258
rect 526144 128258 526186 128494
rect 526422 128258 526464 128494
rect 526144 121494 526464 128258
rect 526144 121258 526186 121494
rect 526422 121258 526464 121494
rect 526144 114494 526464 121258
rect 526144 114258 526186 114494
rect 526422 114258 526464 114494
rect 526144 107494 526464 114258
rect 526144 107258 526186 107494
rect 526422 107258 526464 107494
rect 526144 100494 526464 107258
rect 526144 100258 526186 100494
rect 526422 100258 526464 100494
rect 526144 93494 526464 100258
rect 526144 93258 526186 93494
rect 526422 93258 526464 93494
rect 526144 86494 526464 93258
rect 526144 86258 526186 86494
rect 526422 86258 526464 86494
rect 526144 79494 526464 86258
rect 526144 79258 526186 79494
rect 526422 79258 526464 79494
rect 526144 72494 526464 79258
rect 526144 72258 526186 72494
rect 526422 72258 526464 72494
rect 526144 65494 526464 72258
rect 526144 65258 526186 65494
rect 526422 65258 526464 65494
rect 526144 58494 526464 65258
rect 526144 58258 526186 58494
rect 526422 58258 526464 58494
rect 526144 51494 526464 58258
rect 526144 51258 526186 51494
rect 526422 51258 526464 51494
rect 526144 44494 526464 51258
rect 526144 44258 526186 44494
rect 526422 44258 526464 44494
rect 526144 37494 526464 44258
rect 526144 37258 526186 37494
rect 526422 37258 526464 37494
rect 526144 30494 526464 37258
rect 526144 30258 526186 30494
rect 526422 30258 526464 30494
rect 526144 23494 526464 30258
rect 526144 23258 526186 23494
rect 526422 23258 526464 23494
rect 526144 16494 526464 23258
rect 526144 16258 526186 16494
rect 526422 16258 526464 16494
rect 526144 9494 526464 16258
rect 526144 9258 526186 9494
rect 526422 9258 526464 9494
rect 526144 2494 526464 9258
rect 526144 2258 526186 2494
rect 526422 2258 526464 2494
rect 526144 -746 526464 2258
rect 526144 -982 526186 -746
rect 526422 -982 526464 -746
rect 526144 -1066 526464 -982
rect 526144 -1302 526186 -1066
rect 526422 -1302 526464 -1066
rect 526144 -2294 526464 -1302
rect 527876 234561 528196 241325
rect 527876 234325 527918 234561
rect 528154 234325 528196 234561
rect 527876 227561 528196 234325
rect 527876 227325 527918 227561
rect 528154 227325 528196 227561
rect 527876 220561 528196 227325
rect 527876 220325 527918 220561
rect 528154 220325 528196 220561
rect 527876 213561 528196 220325
rect 527876 213325 527918 213561
rect 528154 213325 528196 213561
rect 527876 206561 528196 213325
rect 527876 206325 527918 206561
rect 528154 206325 528196 206561
rect 527876 199561 528196 206325
rect 527876 199325 527918 199561
rect 528154 199325 528196 199561
rect 527876 192561 528196 199325
rect 527876 192325 527918 192561
rect 528154 192325 528196 192561
rect 527876 185561 528196 192325
rect 527876 185325 527918 185561
rect 528154 185325 528196 185561
rect 527876 178561 528196 185325
rect 527876 178325 527918 178561
rect 528154 178325 528196 178561
rect 527876 171561 528196 178325
rect 527876 171325 527918 171561
rect 528154 171325 528196 171561
rect 527876 164561 528196 171325
rect 527876 164325 527918 164561
rect 528154 164325 528196 164561
rect 527876 157561 528196 164325
rect 527876 157325 527918 157561
rect 528154 157325 528196 157561
rect 527876 150561 528196 157325
rect 527876 150325 527918 150561
rect 528154 150325 528196 150561
rect 527876 143561 528196 150325
rect 527876 143325 527918 143561
rect 528154 143325 528196 143561
rect 527876 136561 528196 143325
rect 527876 136325 527918 136561
rect 528154 136325 528196 136561
rect 527876 129561 528196 136325
rect 527876 129325 527918 129561
rect 528154 129325 528196 129561
rect 527876 122561 528196 129325
rect 527876 122325 527918 122561
rect 528154 122325 528196 122561
rect 527876 115561 528196 122325
rect 527876 115325 527918 115561
rect 528154 115325 528196 115561
rect 527876 108561 528196 115325
rect 527876 108325 527918 108561
rect 528154 108325 528196 108561
rect 527876 101561 528196 108325
rect 527876 101325 527918 101561
rect 528154 101325 528196 101561
rect 527876 94561 528196 101325
rect 527876 94325 527918 94561
rect 528154 94325 528196 94561
rect 527876 87561 528196 94325
rect 527876 87325 527918 87561
rect 528154 87325 528196 87561
rect 527876 80561 528196 87325
rect 527876 80325 527918 80561
rect 528154 80325 528196 80561
rect 527876 73561 528196 80325
rect 527876 73325 527918 73561
rect 528154 73325 528196 73561
rect 527876 66561 528196 73325
rect 527876 66325 527918 66561
rect 528154 66325 528196 66561
rect 527876 59561 528196 66325
rect 527876 59325 527918 59561
rect 528154 59325 528196 59561
rect 527876 52561 528196 59325
rect 527876 52325 527918 52561
rect 528154 52325 528196 52561
rect 527876 45561 528196 52325
rect 527876 45325 527918 45561
rect 528154 45325 528196 45561
rect 527876 38561 528196 45325
rect 527876 38325 527918 38561
rect 528154 38325 528196 38561
rect 527876 31561 528196 38325
rect 527876 31325 527918 31561
rect 528154 31325 528196 31561
rect 527876 24561 528196 31325
rect 527876 24325 527918 24561
rect 528154 24325 528196 24561
rect 527876 17561 528196 24325
rect 527876 17325 527918 17561
rect 528154 17325 528196 17561
rect 527876 10561 528196 17325
rect 527876 10325 527918 10561
rect 528154 10325 528196 10561
rect 527876 3561 528196 10325
rect 527876 3325 527918 3561
rect 528154 3325 528196 3561
rect 527876 -1706 528196 3325
rect 527876 -1942 527918 -1706
rect 528154 -1942 528196 -1706
rect 527876 -2026 528196 -1942
rect 527876 -2262 527918 -2026
rect 528154 -2262 528196 -2026
rect 527876 -2294 528196 -2262
rect 533144 705238 533464 706230
rect 533144 705002 533186 705238
rect 533422 705002 533464 705238
rect 533144 704918 533464 705002
rect 533144 704682 533186 704918
rect 533422 704682 533464 704918
rect 533144 695494 533464 704682
rect 533144 695258 533186 695494
rect 533422 695258 533464 695494
rect 533144 688494 533464 695258
rect 533144 688258 533186 688494
rect 533422 688258 533464 688494
rect 533144 681494 533464 688258
rect 533144 681258 533186 681494
rect 533422 681258 533464 681494
rect 533144 674494 533464 681258
rect 533144 674258 533186 674494
rect 533422 674258 533464 674494
rect 533144 667494 533464 674258
rect 533144 667258 533186 667494
rect 533422 667258 533464 667494
rect 533144 660494 533464 667258
rect 533144 660258 533186 660494
rect 533422 660258 533464 660494
rect 533144 653494 533464 660258
rect 533144 653258 533186 653494
rect 533422 653258 533464 653494
rect 533144 646494 533464 653258
rect 533144 646258 533186 646494
rect 533422 646258 533464 646494
rect 533144 639494 533464 646258
rect 533144 639258 533186 639494
rect 533422 639258 533464 639494
rect 533144 632494 533464 639258
rect 533144 632258 533186 632494
rect 533422 632258 533464 632494
rect 533144 625494 533464 632258
rect 533144 625258 533186 625494
rect 533422 625258 533464 625494
rect 533144 618494 533464 625258
rect 533144 618258 533186 618494
rect 533422 618258 533464 618494
rect 533144 611494 533464 618258
rect 533144 611258 533186 611494
rect 533422 611258 533464 611494
rect 533144 604494 533464 611258
rect 533144 604258 533186 604494
rect 533422 604258 533464 604494
rect 533144 597494 533464 604258
rect 533144 597258 533186 597494
rect 533422 597258 533464 597494
rect 533144 590494 533464 597258
rect 533144 590258 533186 590494
rect 533422 590258 533464 590494
rect 533144 583494 533464 590258
rect 533144 583258 533186 583494
rect 533422 583258 533464 583494
rect 533144 576494 533464 583258
rect 533144 576258 533186 576494
rect 533422 576258 533464 576494
rect 533144 569494 533464 576258
rect 533144 569258 533186 569494
rect 533422 569258 533464 569494
rect 533144 562494 533464 569258
rect 533144 562258 533186 562494
rect 533422 562258 533464 562494
rect 533144 555494 533464 562258
rect 533144 555258 533186 555494
rect 533422 555258 533464 555494
rect 533144 548494 533464 555258
rect 533144 548258 533186 548494
rect 533422 548258 533464 548494
rect 533144 541494 533464 548258
rect 533144 541258 533186 541494
rect 533422 541258 533464 541494
rect 533144 534494 533464 541258
rect 533144 534258 533186 534494
rect 533422 534258 533464 534494
rect 533144 527494 533464 534258
rect 533144 527258 533186 527494
rect 533422 527258 533464 527494
rect 533144 520494 533464 527258
rect 533144 520258 533186 520494
rect 533422 520258 533464 520494
rect 533144 513494 533464 520258
rect 533144 513258 533186 513494
rect 533422 513258 533464 513494
rect 533144 506494 533464 513258
rect 533144 506258 533186 506494
rect 533422 506258 533464 506494
rect 533144 499494 533464 506258
rect 533144 499258 533186 499494
rect 533422 499258 533464 499494
rect 533144 492494 533464 499258
rect 533144 492258 533186 492494
rect 533422 492258 533464 492494
rect 533144 485494 533464 492258
rect 533144 485258 533186 485494
rect 533422 485258 533464 485494
rect 533144 478494 533464 485258
rect 533144 478258 533186 478494
rect 533422 478258 533464 478494
rect 533144 471494 533464 478258
rect 533144 471258 533186 471494
rect 533422 471258 533464 471494
rect 533144 464494 533464 471258
rect 533144 464258 533186 464494
rect 533422 464258 533464 464494
rect 533144 457494 533464 464258
rect 533144 457258 533186 457494
rect 533422 457258 533464 457494
rect 533144 450494 533464 457258
rect 533144 450258 533186 450494
rect 533422 450258 533464 450494
rect 533144 443494 533464 450258
rect 533144 443258 533186 443494
rect 533422 443258 533464 443494
rect 533144 436494 533464 443258
rect 533144 436258 533186 436494
rect 533422 436258 533464 436494
rect 533144 429494 533464 436258
rect 533144 429258 533186 429494
rect 533422 429258 533464 429494
rect 533144 422494 533464 429258
rect 533144 422258 533186 422494
rect 533422 422258 533464 422494
rect 533144 415494 533464 422258
rect 533144 415258 533186 415494
rect 533422 415258 533464 415494
rect 533144 408494 533464 415258
rect 533144 408258 533186 408494
rect 533422 408258 533464 408494
rect 533144 401494 533464 408258
rect 533144 401258 533186 401494
rect 533422 401258 533464 401494
rect 533144 394494 533464 401258
rect 533144 394258 533186 394494
rect 533422 394258 533464 394494
rect 533144 387494 533464 394258
rect 533144 387258 533186 387494
rect 533422 387258 533464 387494
rect 533144 380494 533464 387258
rect 533144 380258 533186 380494
rect 533422 380258 533464 380494
rect 533144 373494 533464 380258
rect 533144 373258 533186 373494
rect 533422 373258 533464 373494
rect 533144 366494 533464 373258
rect 533144 366258 533186 366494
rect 533422 366258 533464 366494
rect 533144 359494 533464 366258
rect 533144 359258 533186 359494
rect 533422 359258 533464 359494
rect 533144 352494 533464 359258
rect 533144 352258 533186 352494
rect 533422 352258 533464 352494
rect 533144 345494 533464 352258
rect 533144 345258 533186 345494
rect 533422 345258 533464 345494
rect 533144 338494 533464 345258
rect 533144 338258 533186 338494
rect 533422 338258 533464 338494
rect 533144 331494 533464 338258
rect 533144 331258 533186 331494
rect 533422 331258 533464 331494
rect 533144 324494 533464 331258
rect 533144 324258 533186 324494
rect 533422 324258 533464 324494
rect 533144 317494 533464 324258
rect 533144 317258 533186 317494
rect 533422 317258 533464 317494
rect 533144 310494 533464 317258
rect 533144 310258 533186 310494
rect 533422 310258 533464 310494
rect 533144 303494 533464 310258
rect 533144 303258 533186 303494
rect 533422 303258 533464 303494
rect 533144 296494 533464 303258
rect 533144 296258 533186 296494
rect 533422 296258 533464 296494
rect 533144 289494 533464 296258
rect 533144 289258 533186 289494
rect 533422 289258 533464 289494
rect 533144 282494 533464 289258
rect 533144 282258 533186 282494
rect 533422 282258 533464 282494
rect 533144 275494 533464 282258
rect 533144 275258 533186 275494
rect 533422 275258 533464 275494
rect 533144 268494 533464 275258
rect 533144 268258 533186 268494
rect 533422 268258 533464 268494
rect 533144 261494 533464 268258
rect 533144 261258 533186 261494
rect 533422 261258 533464 261494
rect 533144 254494 533464 261258
rect 533144 254258 533186 254494
rect 533422 254258 533464 254494
rect 533144 247494 533464 254258
rect 533144 247258 533186 247494
rect 533422 247258 533464 247494
rect 533144 240494 533464 247258
rect 533144 240258 533186 240494
rect 533422 240258 533464 240494
rect 533144 233494 533464 240258
rect 533144 233258 533186 233494
rect 533422 233258 533464 233494
rect 533144 226494 533464 233258
rect 533144 226258 533186 226494
rect 533422 226258 533464 226494
rect 533144 219494 533464 226258
rect 533144 219258 533186 219494
rect 533422 219258 533464 219494
rect 533144 212494 533464 219258
rect 533144 212258 533186 212494
rect 533422 212258 533464 212494
rect 533144 205494 533464 212258
rect 533144 205258 533186 205494
rect 533422 205258 533464 205494
rect 533144 198494 533464 205258
rect 533144 198258 533186 198494
rect 533422 198258 533464 198494
rect 533144 191494 533464 198258
rect 533144 191258 533186 191494
rect 533422 191258 533464 191494
rect 533144 184494 533464 191258
rect 533144 184258 533186 184494
rect 533422 184258 533464 184494
rect 533144 177494 533464 184258
rect 533144 177258 533186 177494
rect 533422 177258 533464 177494
rect 533144 170494 533464 177258
rect 533144 170258 533186 170494
rect 533422 170258 533464 170494
rect 533144 163494 533464 170258
rect 533144 163258 533186 163494
rect 533422 163258 533464 163494
rect 533144 156494 533464 163258
rect 533144 156258 533186 156494
rect 533422 156258 533464 156494
rect 533144 149494 533464 156258
rect 533144 149258 533186 149494
rect 533422 149258 533464 149494
rect 533144 142494 533464 149258
rect 533144 142258 533186 142494
rect 533422 142258 533464 142494
rect 533144 135494 533464 142258
rect 533144 135258 533186 135494
rect 533422 135258 533464 135494
rect 533144 128494 533464 135258
rect 533144 128258 533186 128494
rect 533422 128258 533464 128494
rect 533144 121494 533464 128258
rect 533144 121258 533186 121494
rect 533422 121258 533464 121494
rect 533144 114494 533464 121258
rect 533144 114258 533186 114494
rect 533422 114258 533464 114494
rect 533144 107494 533464 114258
rect 533144 107258 533186 107494
rect 533422 107258 533464 107494
rect 533144 100494 533464 107258
rect 533144 100258 533186 100494
rect 533422 100258 533464 100494
rect 533144 93494 533464 100258
rect 533144 93258 533186 93494
rect 533422 93258 533464 93494
rect 533144 86494 533464 93258
rect 533144 86258 533186 86494
rect 533422 86258 533464 86494
rect 533144 79494 533464 86258
rect 533144 79258 533186 79494
rect 533422 79258 533464 79494
rect 533144 72494 533464 79258
rect 533144 72258 533186 72494
rect 533422 72258 533464 72494
rect 533144 65494 533464 72258
rect 533144 65258 533186 65494
rect 533422 65258 533464 65494
rect 533144 58494 533464 65258
rect 533144 58258 533186 58494
rect 533422 58258 533464 58494
rect 533144 51494 533464 58258
rect 533144 51258 533186 51494
rect 533422 51258 533464 51494
rect 533144 44494 533464 51258
rect 533144 44258 533186 44494
rect 533422 44258 533464 44494
rect 533144 37494 533464 44258
rect 533144 37258 533186 37494
rect 533422 37258 533464 37494
rect 533144 30494 533464 37258
rect 533144 30258 533186 30494
rect 533422 30258 533464 30494
rect 533144 23494 533464 30258
rect 533144 23258 533186 23494
rect 533422 23258 533464 23494
rect 533144 16494 533464 23258
rect 533144 16258 533186 16494
rect 533422 16258 533464 16494
rect 533144 9494 533464 16258
rect 533144 9258 533186 9494
rect 533422 9258 533464 9494
rect 533144 2494 533464 9258
rect 533144 2258 533186 2494
rect 533422 2258 533464 2494
rect 533144 -746 533464 2258
rect 533144 -982 533186 -746
rect 533422 -982 533464 -746
rect 533144 -1066 533464 -982
rect 533144 -1302 533186 -1066
rect 533422 -1302 533464 -1066
rect 533144 -2294 533464 -1302
rect 534876 706198 535196 706230
rect 534876 705962 534918 706198
rect 535154 705962 535196 706198
rect 534876 705878 535196 705962
rect 534876 705642 534918 705878
rect 535154 705642 535196 705878
rect 534876 696561 535196 705642
rect 534876 696325 534918 696561
rect 535154 696325 535196 696561
rect 534876 689561 535196 696325
rect 534876 689325 534918 689561
rect 535154 689325 535196 689561
rect 534876 682561 535196 689325
rect 534876 682325 534918 682561
rect 535154 682325 535196 682561
rect 534876 675561 535196 682325
rect 534876 675325 534918 675561
rect 535154 675325 535196 675561
rect 534876 668561 535196 675325
rect 534876 668325 534918 668561
rect 535154 668325 535196 668561
rect 534876 661561 535196 668325
rect 534876 661325 534918 661561
rect 535154 661325 535196 661561
rect 534876 654561 535196 661325
rect 534876 654325 534918 654561
rect 535154 654325 535196 654561
rect 534876 647561 535196 654325
rect 534876 647325 534918 647561
rect 535154 647325 535196 647561
rect 534876 640561 535196 647325
rect 534876 640325 534918 640561
rect 535154 640325 535196 640561
rect 534876 633561 535196 640325
rect 534876 633325 534918 633561
rect 535154 633325 535196 633561
rect 534876 626561 535196 633325
rect 534876 626325 534918 626561
rect 535154 626325 535196 626561
rect 534876 619561 535196 626325
rect 534876 619325 534918 619561
rect 535154 619325 535196 619561
rect 534876 612561 535196 619325
rect 534876 612325 534918 612561
rect 535154 612325 535196 612561
rect 534876 605561 535196 612325
rect 534876 605325 534918 605561
rect 535154 605325 535196 605561
rect 534876 598561 535196 605325
rect 534876 598325 534918 598561
rect 535154 598325 535196 598561
rect 534876 591561 535196 598325
rect 534876 591325 534918 591561
rect 535154 591325 535196 591561
rect 534876 584561 535196 591325
rect 534876 584325 534918 584561
rect 535154 584325 535196 584561
rect 534876 577561 535196 584325
rect 534876 577325 534918 577561
rect 535154 577325 535196 577561
rect 534876 570561 535196 577325
rect 534876 570325 534918 570561
rect 535154 570325 535196 570561
rect 534876 563561 535196 570325
rect 534876 563325 534918 563561
rect 535154 563325 535196 563561
rect 534876 556561 535196 563325
rect 534876 556325 534918 556561
rect 535154 556325 535196 556561
rect 534876 549561 535196 556325
rect 534876 549325 534918 549561
rect 535154 549325 535196 549561
rect 534876 542561 535196 549325
rect 534876 542325 534918 542561
rect 535154 542325 535196 542561
rect 534876 535561 535196 542325
rect 534876 535325 534918 535561
rect 535154 535325 535196 535561
rect 534876 528561 535196 535325
rect 534876 528325 534918 528561
rect 535154 528325 535196 528561
rect 534876 521561 535196 528325
rect 534876 521325 534918 521561
rect 535154 521325 535196 521561
rect 534876 514561 535196 521325
rect 534876 514325 534918 514561
rect 535154 514325 535196 514561
rect 534876 507561 535196 514325
rect 534876 507325 534918 507561
rect 535154 507325 535196 507561
rect 534876 500561 535196 507325
rect 534876 500325 534918 500561
rect 535154 500325 535196 500561
rect 534876 493561 535196 500325
rect 534876 493325 534918 493561
rect 535154 493325 535196 493561
rect 534876 486561 535196 493325
rect 534876 486325 534918 486561
rect 535154 486325 535196 486561
rect 534876 479561 535196 486325
rect 534876 479325 534918 479561
rect 535154 479325 535196 479561
rect 534876 472561 535196 479325
rect 534876 472325 534918 472561
rect 535154 472325 535196 472561
rect 534876 465561 535196 472325
rect 534876 465325 534918 465561
rect 535154 465325 535196 465561
rect 534876 458561 535196 465325
rect 534876 458325 534918 458561
rect 535154 458325 535196 458561
rect 534876 451561 535196 458325
rect 534876 451325 534918 451561
rect 535154 451325 535196 451561
rect 534876 444561 535196 451325
rect 534876 444325 534918 444561
rect 535154 444325 535196 444561
rect 534876 437561 535196 444325
rect 534876 437325 534918 437561
rect 535154 437325 535196 437561
rect 534876 430561 535196 437325
rect 534876 430325 534918 430561
rect 535154 430325 535196 430561
rect 534876 423561 535196 430325
rect 534876 423325 534918 423561
rect 535154 423325 535196 423561
rect 534876 416561 535196 423325
rect 534876 416325 534918 416561
rect 535154 416325 535196 416561
rect 534876 409561 535196 416325
rect 534876 409325 534918 409561
rect 535154 409325 535196 409561
rect 534876 402561 535196 409325
rect 534876 402325 534918 402561
rect 535154 402325 535196 402561
rect 534876 395561 535196 402325
rect 534876 395325 534918 395561
rect 535154 395325 535196 395561
rect 534876 388561 535196 395325
rect 534876 388325 534918 388561
rect 535154 388325 535196 388561
rect 534876 381561 535196 388325
rect 534876 381325 534918 381561
rect 535154 381325 535196 381561
rect 534876 374561 535196 381325
rect 534876 374325 534918 374561
rect 535154 374325 535196 374561
rect 534876 367561 535196 374325
rect 534876 367325 534918 367561
rect 535154 367325 535196 367561
rect 534876 360561 535196 367325
rect 534876 360325 534918 360561
rect 535154 360325 535196 360561
rect 534876 353561 535196 360325
rect 534876 353325 534918 353561
rect 535154 353325 535196 353561
rect 534876 346561 535196 353325
rect 534876 346325 534918 346561
rect 535154 346325 535196 346561
rect 534876 339561 535196 346325
rect 534876 339325 534918 339561
rect 535154 339325 535196 339561
rect 534876 332561 535196 339325
rect 534876 332325 534918 332561
rect 535154 332325 535196 332561
rect 534876 325561 535196 332325
rect 534876 325325 534918 325561
rect 535154 325325 535196 325561
rect 534876 318561 535196 325325
rect 534876 318325 534918 318561
rect 535154 318325 535196 318561
rect 534876 311561 535196 318325
rect 534876 311325 534918 311561
rect 535154 311325 535196 311561
rect 534876 304561 535196 311325
rect 534876 304325 534918 304561
rect 535154 304325 535196 304561
rect 534876 297561 535196 304325
rect 534876 297325 534918 297561
rect 535154 297325 535196 297561
rect 534876 290561 535196 297325
rect 534876 290325 534918 290561
rect 535154 290325 535196 290561
rect 534876 283561 535196 290325
rect 534876 283325 534918 283561
rect 535154 283325 535196 283561
rect 534876 276561 535196 283325
rect 534876 276325 534918 276561
rect 535154 276325 535196 276561
rect 534876 269561 535196 276325
rect 534876 269325 534918 269561
rect 535154 269325 535196 269561
rect 534876 262561 535196 269325
rect 534876 262325 534918 262561
rect 535154 262325 535196 262561
rect 534876 255561 535196 262325
rect 534876 255325 534918 255561
rect 535154 255325 535196 255561
rect 534876 248561 535196 255325
rect 534876 248325 534918 248561
rect 535154 248325 535196 248561
rect 534876 241561 535196 248325
rect 534876 241325 534918 241561
rect 535154 241325 535196 241561
rect 534876 234561 535196 241325
rect 534876 234325 534918 234561
rect 535154 234325 535196 234561
rect 534876 227561 535196 234325
rect 534876 227325 534918 227561
rect 535154 227325 535196 227561
rect 534876 220561 535196 227325
rect 534876 220325 534918 220561
rect 535154 220325 535196 220561
rect 534876 213561 535196 220325
rect 534876 213325 534918 213561
rect 535154 213325 535196 213561
rect 534876 206561 535196 213325
rect 534876 206325 534918 206561
rect 535154 206325 535196 206561
rect 534876 199561 535196 206325
rect 534876 199325 534918 199561
rect 535154 199325 535196 199561
rect 534876 192561 535196 199325
rect 534876 192325 534918 192561
rect 535154 192325 535196 192561
rect 534876 185561 535196 192325
rect 534876 185325 534918 185561
rect 535154 185325 535196 185561
rect 534876 178561 535196 185325
rect 534876 178325 534918 178561
rect 535154 178325 535196 178561
rect 534876 171561 535196 178325
rect 534876 171325 534918 171561
rect 535154 171325 535196 171561
rect 534876 164561 535196 171325
rect 534876 164325 534918 164561
rect 535154 164325 535196 164561
rect 534876 157561 535196 164325
rect 534876 157325 534918 157561
rect 535154 157325 535196 157561
rect 534876 150561 535196 157325
rect 534876 150325 534918 150561
rect 535154 150325 535196 150561
rect 534876 143561 535196 150325
rect 534876 143325 534918 143561
rect 535154 143325 535196 143561
rect 534876 136561 535196 143325
rect 534876 136325 534918 136561
rect 535154 136325 535196 136561
rect 534876 129561 535196 136325
rect 534876 129325 534918 129561
rect 535154 129325 535196 129561
rect 534876 122561 535196 129325
rect 534876 122325 534918 122561
rect 535154 122325 535196 122561
rect 534876 115561 535196 122325
rect 534876 115325 534918 115561
rect 535154 115325 535196 115561
rect 534876 108561 535196 115325
rect 534876 108325 534918 108561
rect 535154 108325 535196 108561
rect 534876 101561 535196 108325
rect 534876 101325 534918 101561
rect 535154 101325 535196 101561
rect 534876 94561 535196 101325
rect 534876 94325 534918 94561
rect 535154 94325 535196 94561
rect 534876 87561 535196 94325
rect 534876 87325 534918 87561
rect 535154 87325 535196 87561
rect 534876 80561 535196 87325
rect 534876 80325 534918 80561
rect 535154 80325 535196 80561
rect 534876 73561 535196 80325
rect 534876 73325 534918 73561
rect 535154 73325 535196 73561
rect 534876 66561 535196 73325
rect 534876 66325 534918 66561
rect 535154 66325 535196 66561
rect 534876 59561 535196 66325
rect 534876 59325 534918 59561
rect 535154 59325 535196 59561
rect 534876 52561 535196 59325
rect 534876 52325 534918 52561
rect 535154 52325 535196 52561
rect 534876 45561 535196 52325
rect 534876 45325 534918 45561
rect 535154 45325 535196 45561
rect 534876 38561 535196 45325
rect 534876 38325 534918 38561
rect 535154 38325 535196 38561
rect 534876 31561 535196 38325
rect 534876 31325 534918 31561
rect 535154 31325 535196 31561
rect 534876 24561 535196 31325
rect 534876 24325 534918 24561
rect 535154 24325 535196 24561
rect 534876 17561 535196 24325
rect 534876 17325 534918 17561
rect 535154 17325 535196 17561
rect 534876 10561 535196 17325
rect 534876 10325 534918 10561
rect 535154 10325 535196 10561
rect 534876 3561 535196 10325
rect 534876 3325 534918 3561
rect 535154 3325 535196 3561
rect 534876 -1706 535196 3325
rect 534876 -1942 534918 -1706
rect 535154 -1942 535196 -1706
rect 534876 -2026 535196 -1942
rect 534876 -2262 534918 -2026
rect 535154 -2262 535196 -2026
rect 534876 -2294 535196 -2262
rect 540144 705238 540464 706230
rect 540144 705002 540186 705238
rect 540422 705002 540464 705238
rect 540144 704918 540464 705002
rect 540144 704682 540186 704918
rect 540422 704682 540464 704918
rect 540144 695494 540464 704682
rect 540144 695258 540186 695494
rect 540422 695258 540464 695494
rect 540144 688494 540464 695258
rect 540144 688258 540186 688494
rect 540422 688258 540464 688494
rect 540144 681494 540464 688258
rect 540144 681258 540186 681494
rect 540422 681258 540464 681494
rect 540144 674494 540464 681258
rect 540144 674258 540186 674494
rect 540422 674258 540464 674494
rect 540144 667494 540464 674258
rect 540144 667258 540186 667494
rect 540422 667258 540464 667494
rect 540144 660494 540464 667258
rect 540144 660258 540186 660494
rect 540422 660258 540464 660494
rect 540144 653494 540464 660258
rect 540144 653258 540186 653494
rect 540422 653258 540464 653494
rect 540144 646494 540464 653258
rect 540144 646258 540186 646494
rect 540422 646258 540464 646494
rect 540144 639494 540464 646258
rect 540144 639258 540186 639494
rect 540422 639258 540464 639494
rect 540144 632494 540464 639258
rect 540144 632258 540186 632494
rect 540422 632258 540464 632494
rect 540144 625494 540464 632258
rect 540144 625258 540186 625494
rect 540422 625258 540464 625494
rect 540144 618494 540464 625258
rect 540144 618258 540186 618494
rect 540422 618258 540464 618494
rect 540144 611494 540464 618258
rect 540144 611258 540186 611494
rect 540422 611258 540464 611494
rect 540144 604494 540464 611258
rect 540144 604258 540186 604494
rect 540422 604258 540464 604494
rect 540144 597494 540464 604258
rect 540144 597258 540186 597494
rect 540422 597258 540464 597494
rect 540144 590494 540464 597258
rect 540144 590258 540186 590494
rect 540422 590258 540464 590494
rect 540144 583494 540464 590258
rect 540144 583258 540186 583494
rect 540422 583258 540464 583494
rect 540144 576494 540464 583258
rect 540144 576258 540186 576494
rect 540422 576258 540464 576494
rect 540144 569494 540464 576258
rect 540144 569258 540186 569494
rect 540422 569258 540464 569494
rect 540144 562494 540464 569258
rect 540144 562258 540186 562494
rect 540422 562258 540464 562494
rect 540144 555494 540464 562258
rect 540144 555258 540186 555494
rect 540422 555258 540464 555494
rect 540144 548494 540464 555258
rect 540144 548258 540186 548494
rect 540422 548258 540464 548494
rect 540144 541494 540464 548258
rect 540144 541258 540186 541494
rect 540422 541258 540464 541494
rect 540144 534494 540464 541258
rect 540144 534258 540186 534494
rect 540422 534258 540464 534494
rect 540144 527494 540464 534258
rect 540144 527258 540186 527494
rect 540422 527258 540464 527494
rect 540144 520494 540464 527258
rect 540144 520258 540186 520494
rect 540422 520258 540464 520494
rect 540144 513494 540464 520258
rect 540144 513258 540186 513494
rect 540422 513258 540464 513494
rect 540144 506494 540464 513258
rect 540144 506258 540186 506494
rect 540422 506258 540464 506494
rect 540144 499494 540464 506258
rect 540144 499258 540186 499494
rect 540422 499258 540464 499494
rect 540144 492494 540464 499258
rect 540144 492258 540186 492494
rect 540422 492258 540464 492494
rect 540144 485494 540464 492258
rect 540144 485258 540186 485494
rect 540422 485258 540464 485494
rect 540144 478494 540464 485258
rect 540144 478258 540186 478494
rect 540422 478258 540464 478494
rect 540144 471494 540464 478258
rect 540144 471258 540186 471494
rect 540422 471258 540464 471494
rect 540144 464494 540464 471258
rect 540144 464258 540186 464494
rect 540422 464258 540464 464494
rect 540144 457494 540464 464258
rect 540144 457258 540186 457494
rect 540422 457258 540464 457494
rect 540144 450494 540464 457258
rect 540144 450258 540186 450494
rect 540422 450258 540464 450494
rect 540144 443494 540464 450258
rect 540144 443258 540186 443494
rect 540422 443258 540464 443494
rect 540144 436494 540464 443258
rect 540144 436258 540186 436494
rect 540422 436258 540464 436494
rect 540144 429494 540464 436258
rect 540144 429258 540186 429494
rect 540422 429258 540464 429494
rect 540144 422494 540464 429258
rect 540144 422258 540186 422494
rect 540422 422258 540464 422494
rect 540144 415494 540464 422258
rect 540144 415258 540186 415494
rect 540422 415258 540464 415494
rect 540144 408494 540464 415258
rect 540144 408258 540186 408494
rect 540422 408258 540464 408494
rect 540144 401494 540464 408258
rect 540144 401258 540186 401494
rect 540422 401258 540464 401494
rect 540144 394494 540464 401258
rect 540144 394258 540186 394494
rect 540422 394258 540464 394494
rect 540144 387494 540464 394258
rect 540144 387258 540186 387494
rect 540422 387258 540464 387494
rect 540144 380494 540464 387258
rect 540144 380258 540186 380494
rect 540422 380258 540464 380494
rect 540144 373494 540464 380258
rect 540144 373258 540186 373494
rect 540422 373258 540464 373494
rect 540144 366494 540464 373258
rect 540144 366258 540186 366494
rect 540422 366258 540464 366494
rect 540144 359494 540464 366258
rect 540144 359258 540186 359494
rect 540422 359258 540464 359494
rect 540144 352494 540464 359258
rect 540144 352258 540186 352494
rect 540422 352258 540464 352494
rect 540144 345494 540464 352258
rect 540144 345258 540186 345494
rect 540422 345258 540464 345494
rect 540144 338494 540464 345258
rect 540144 338258 540186 338494
rect 540422 338258 540464 338494
rect 540144 331494 540464 338258
rect 540144 331258 540186 331494
rect 540422 331258 540464 331494
rect 540144 324494 540464 331258
rect 540144 324258 540186 324494
rect 540422 324258 540464 324494
rect 540144 317494 540464 324258
rect 540144 317258 540186 317494
rect 540422 317258 540464 317494
rect 540144 310494 540464 317258
rect 540144 310258 540186 310494
rect 540422 310258 540464 310494
rect 540144 303494 540464 310258
rect 540144 303258 540186 303494
rect 540422 303258 540464 303494
rect 540144 296494 540464 303258
rect 540144 296258 540186 296494
rect 540422 296258 540464 296494
rect 540144 289494 540464 296258
rect 540144 289258 540186 289494
rect 540422 289258 540464 289494
rect 540144 282494 540464 289258
rect 540144 282258 540186 282494
rect 540422 282258 540464 282494
rect 540144 275494 540464 282258
rect 540144 275258 540186 275494
rect 540422 275258 540464 275494
rect 540144 268494 540464 275258
rect 540144 268258 540186 268494
rect 540422 268258 540464 268494
rect 540144 261494 540464 268258
rect 540144 261258 540186 261494
rect 540422 261258 540464 261494
rect 540144 254494 540464 261258
rect 540144 254258 540186 254494
rect 540422 254258 540464 254494
rect 540144 247494 540464 254258
rect 540144 247258 540186 247494
rect 540422 247258 540464 247494
rect 540144 240494 540464 247258
rect 540144 240258 540186 240494
rect 540422 240258 540464 240494
rect 540144 233494 540464 240258
rect 540144 233258 540186 233494
rect 540422 233258 540464 233494
rect 540144 226494 540464 233258
rect 540144 226258 540186 226494
rect 540422 226258 540464 226494
rect 540144 219494 540464 226258
rect 540144 219258 540186 219494
rect 540422 219258 540464 219494
rect 540144 212494 540464 219258
rect 540144 212258 540186 212494
rect 540422 212258 540464 212494
rect 540144 205494 540464 212258
rect 540144 205258 540186 205494
rect 540422 205258 540464 205494
rect 540144 198494 540464 205258
rect 540144 198258 540186 198494
rect 540422 198258 540464 198494
rect 540144 191494 540464 198258
rect 540144 191258 540186 191494
rect 540422 191258 540464 191494
rect 540144 184494 540464 191258
rect 540144 184258 540186 184494
rect 540422 184258 540464 184494
rect 540144 177494 540464 184258
rect 540144 177258 540186 177494
rect 540422 177258 540464 177494
rect 540144 170494 540464 177258
rect 540144 170258 540186 170494
rect 540422 170258 540464 170494
rect 540144 163494 540464 170258
rect 540144 163258 540186 163494
rect 540422 163258 540464 163494
rect 540144 156494 540464 163258
rect 540144 156258 540186 156494
rect 540422 156258 540464 156494
rect 540144 149494 540464 156258
rect 540144 149258 540186 149494
rect 540422 149258 540464 149494
rect 540144 142494 540464 149258
rect 540144 142258 540186 142494
rect 540422 142258 540464 142494
rect 540144 135494 540464 142258
rect 540144 135258 540186 135494
rect 540422 135258 540464 135494
rect 540144 128494 540464 135258
rect 540144 128258 540186 128494
rect 540422 128258 540464 128494
rect 540144 121494 540464 128258
rect 540144 121258 540186 121494
rect 540422 121258 540464 121494
rect 540144 114494 540464 121258
rect 540144 114258 540186 114494
rect 540422 114258 540464 114494
rect 540144 107494 540464 114258
rect 540144 107258 540186 107494
rect 540422 107258 540464 107494
rect 540144 100494 540464 107258
rect 540144 100258 540186 100494
rect 540422 100258 540464 100494
rect 540144 93494 540464 100258
rect 540144 93258 540186 93494
rect 540422 93258 540464 93494
rect 540144 86494 540464 93258
rect 540144 86258 540186 86494
rect 540422 86258 540464 86494
rect 540144 79494 540464 86258
rect 540144 79258 540186 79494
rect 540422 79258 540464 79494
rect 540144 72494 540464 79258
rect 540144 72258 540186 72494
rect 540422 72258 540464 72494
rect 540144 65494 540464 72258
rect 540144 65258 540186 65494
rect 540422 65258 540464 65494
rect 540144 58494 540464 65258
rect 540144 58258 540186 58494
rect 540422 58258 540464 58494
rect 540144 51494 540464 58258
rect 540144 51258 540186 51494
rect 540422 51258 540464 51494
rect 540144 44494 540464 51258
rect 540144 44258 540186 44494
rect 540422 44258 540464 44494
rect 540144 37494 540464 44258
rect 540144 37258 540186 37494
rect 540422 37258 540464 37494
rect 540144 30494 540464 37258
rect 540144 30258 540186 30494
rect 540422 30258 540464 30494
rect 540144 23494 540464 30258
rect 540144 23258 540186 23494
rect 540422 23258 540464 23494
rect 540144 16494 540464 23258
rect 540144 16258 540186 16494
rect 540422 16258 540464 16494
rect 540144 9494 540464 16258
rect 540144 9258 540186 9494
rect 540422 9258 540464 9494
rect 540144 2494 540464 9258
rect 540144 2258 540186 2494
rect 540422 2258 540464 2494
rect 540144 -746 540464 2258
rect 540144 -982 540186 -746
rect 540422 -982 540464 -746
rect 540144 -1066 540464 -982
rect 540144 -1302 540186 -1066
rect 540422 -1302 540464 -1066
rect 540144 -2294 540464 -1302
rect 541876 706198 542196 706230
rect 541876 705962 541918 706198
rect 542154 705962 542196 706198
rect 541876 705878 542196 705962
rect 541876 705642 541918 705878
rect 542154 705642 542196 705878
rect 541876 696561 542196 705642
rect 541876 696325 541918 696561
rect 542154 696325 542196 696561
rect 541876 689561 542196 696325
rect 541876 689325 541918 689561
rect 542154 689325 542196 689561
rect 541876 682561 542196 689325
rect 541876 682325 541918 682561
rect 542154 682325 542196 682561
rect 541876 675561 542196 682325
rect 541876 675325 541918 675561
rect 542154 675325 542196 675561
rect 541876 668561 542196 675325
rect 541876 668325 541918 668561
rect 542154 668325 542196 668561
rect 541876 661561 542196 668325
rect 541876 661325 541918 661561
rect 542154 661325 542196 661561
rect 541876 654561 542196 661325
rect 541876 654325 541918 654561
rect 542154 654325 542196 654561
rect 541876 647561 542196 654325
rect 541876 647325 541918 647561
rect 542154 647325 542196 647561
rect 541876 640561 542196 647325
rect 541876 640325 541918 640561
rect 542154 640325 542196 640561
rect 541876 633561 542196 640325
rect 541876 633325 541918 633561
rect 542154 633325 542196 633561
rect 541876 626561 542196 633325
rect 541876 626325 541918 626561
rect 542154 626325 542196 626561
rect 541876 619561 542196 626325
rect 541876 619325 541918 619561
rect 542154 619325 542196 619561
rect 541876 612561 542196 619325
rect 541876 612325 541918 612561
rect 542154 612325 542196 612561
rect 541876 605561 542196 612325
rect 541876 605325 541918 605561
rect 542154 605325 542196 605561
rect 541876 598561 542196 605325
rect 541876 598325 541918 598561
rect 542154 598325 542196 598561
rect 541876 591561 542196 598325
rect 541876 591325 541918 591561
rect 542154 591325 542196 591561
rect 541876 584561 542196 591325
rect 541876 584325 541918 584561
rect 542154 584325 542196 584561
rect 541876 577561 542196 584325
rect 541876 577325 541918 577561
rect 542154 577325 542196 577561
rect 541876 570561 542196 577325
rect 541876 570325 541918 570561
rect 542154 570325 542196 570561
rect 541876 563561 542196 570325
rect 541876 563325 541918 563561
rect 542154 563325 542196 563561
rect 541876 556561 542196 563325
rect 541876 556325 541918 556561
rect 542154 556325 542196 556561
rect 541876 549561 542196 556325
rect 541876 549325 541918 549561
rect 542154 549325 542196 549561
rect 541876 542561 542196 549325
rect 541876 542325 541918 542561
rect 542154 542325 542196 542561
rect 541876 535561 542196 542325
rect 541876 535325 541918 535561
rect 542154 535325 542196 535561
rect 541876 528561 542196 535325
rect 541876 528325 541918 528561
rect 542154 528325 542196 528561
rect 541876 521561 542196 528325
rect 541876 521325 541918 521561
rect 542154 521325 542196 521561
rect 541876 514561 542196 521325
rect 541876 514325 541918 514561
rect 542154 514325 542196 514561
rect 541876 507561 542196 514325
rect 541876 507325 541918 507561
rect 542154 507325 542196 507561
rect 541876 500561 542196 507325
rect 541876 500325 541918 500561
rect 542154 500325 542196 500561
rect 541876 493561 542196 500325
rect 541876 493325 541918 493561
rect 542154 493325 542196 493561
rect 541876 486561 542196 493325
rect 541876 486325 541918 486561
rect 542154 486325 542196 486561
rect 541876 479561 542196 486325
rect 541876 479325 541918 479561
rect 542154 479325 542196 479561
rect 541876 472561 542196 479325
rect 541876 472325 541918 472561
rect 542154 472325 542196 472561
rect 541876 465561 542196 472325
rect 541876 465325 541918 465561
rect 542154 465325 542196 465561
rect 541876 458561 542196 465325
rect 541876 458325 541918 458561
rect 542154 458325 542196 458561
rect 541876 451561 542196 458325
rect 541876 451325 541918 451561
rect 542154 451325 542196 451561
rect 541876 444561 542196 451325
rect 541876 444325 541918 444561
rect 542154 444325 542196 444561
rect 541876 437561 542196 444325
rect 541876 437325 541918 437561
rect 542154 437325 542196 437561
rect 541876 430561 542196 437325
rect 541876 430325 541918 430561
rect 542154 430325 542196 430561
rect 541876 423561 542196 430325
rect 541876 423325 541918 423561
rect 542154 423325 542196 423561
rect 541876 416561 542196 423325
rect 541876 416325 541918 416561
rect 542154 416325 542196 416561
rect 541876 409561 542196 416325
rect 541876 409325 541918 409561
rect 542154 409325 542196 409561
rect 541876 402561 542196 409325
rect 541876 402325 541918 402561
rect 542154 402325 542196 402561
rect 541876 395561 542196 402325
rect 541876 395325 541918 395561
rect 542154 395325 542196 395561
rect 541876 388561 542196 395325
rect 541876 388325 541918 388561
rect 542154 388325 542196 388561
rect 541876 381561 542196 388325
rect 541876 381325 541918 381561
rect 542154 381325 542196 381561
rect 541876 374561 542196 381325
rect 541876 374325 541918 374561
rect 542154 374325 542196 374561
rect 541876 367561 542196 374325
rect 541876 367325 541918 367561
rect 542154 367325 542196 367561
rect 541876 360561 542196 367325
rect 541876 360325 541918 360561
rect 542154 360325 542196 360561
rect 541876 353561 542196 360325
rect 541876 353325 541918 353561
rect 542154 353325 542196 353561
rect 541876 346561 542196 353325
rect 541876 346325 541918 346561
rect 542154 346325 542196 346561
rect 541876 339561 542196 346325
rect 541876 339325 541918 339561
rect 542154 339325 542196 339561
rect 541876 332561 542196 339325
rect 541876 332325 541918 332561
rect 542154 332325 542196 332561
rect 541876 325561 542196 332325
rect 541876 325325 541918 325561
rect 542154 325325 542196 325561
rect 541876 318561 542196 325325
rect 541876 318325 541918 318561
rect 542154 318325 542196 318561
rect 541876 311561 542196 318325
rect 541876 311325 541918 311561
rect 542154 311325 542196 311561
rect 541876 304561 542196 311325
rect 541876 304325 541918 304561
rect 542154 304325 542196 304561
rect 541876 297561 542196 304325
rect 541876 297325 541918 297561
rect 542154 297325 542196 297561
rect 541876 290561 542196 297325
rect 541876 290325 541918 290561
rect 542154 290325 542196 290561
rect 541876 283561 542196 290325
rect 541876 283325 541918 283561
rect 542154 283325 542196 283561
rect 541876 276561 542196 283325
rect 541876 276325 541918 276561
rect 542154 276325 542196 276561
rect 541876 269561 542196 276325
rect 541876 269325 541918 269561
rect 542154 269325 542196 269561
rect 541876 262561 542196 269325
rect 541876 262325 541918 262561
rect 542154 262325 542196 262561
rect 541876 255561 542196 262325
rect 541876 255325 541918 255561
rect 542154 255325 542196 255561
rect 541876 248561 542196 255325
rect 541876 248325 541918 248561
rect 542154 248325 542196 248561
rect 541876 241561 542196 248325
rect 541876 241325 541918 241561
rect 542154 241325 542196 241561
rect 541876 234561 542196 241325
rect 541876 234325 541918 234561
rect 542154 234325 542196 234561
rect 541876 227561 542196 234325
rect 541876 227325 541918 227561
rect 542154 227325 542196 227561
rect 541876 220561 542196 227325
rect 541876 220325 541918 220561
rect 542154 220325 542196 220561
rect 541876 213561 542196 220325
rect 541876 213325 541918 213561
rect 542154 213325 542196 213561
rect 541876 206561 542196 213325
rect 541876 206325 541918 206561
rect 542154 206325 542196 206561
rect 541876 199561 542196 206325
rect 541876 199325 541918 199561
rect 542154 199325 542196 199561
rect 541876 192561 542196 199325
rect 541876 192325 541918 192561
rect 542154 192325 542196 192561
rect 541876 185561 542196 192325
rect 541876 185325 541918 185561
rect 542154 185325 542196 185561
rect 541876 178561 542196 185325
rect 541876 178325 541918 178561
rect 542154 178325 542196 178561
rect 541876 171561 542196 178325
rect 541876 171325 541918 171561
rect 542154 171325 542196 171561
rect 541876 164561 542196 171325
rect 541876 164325 541918 164561
rect 542154 164325 542196 164561
rect 541876 157561 542196 164325
rect 541876 157325 541918 157561
rect 542154 157325 542196 157561
rect 541876 150561 542196 157325
rect 541876 150325 541918 150561
rect 542154 150325 542196 150561
rect 541876 143561 542196 150325
rect 541876 143325 541918 143561
rect 542154 143325 542196 143561
rect 541876 136561 542196 143325
rect 541876 136325 541918 136561
rect 542154 136325 542196 136561
rect 541876 129561 542196 136325
rect 541876 129325 541918 129561
rect 542154 129325 542196 129561
rect 541876 122561 542196 129325
rect 541876 122325 541918 122561
rect 542154 122325 542196 122561
rect 541876 115561 542196 122325
rect 541876 115325 541918 115561
rect 542154 115325 542196 115561
rect 541876 108561 542196 115325
rect 541876 108325 541918 108561
rect 542154 108325 542196 108561
rect 541876 101561 542196 108325
rect 541876 101325 541918 101561
rect 542154 101325 542196 101561
rect 541876 94561 542196 101325
rect 541876 94325 541918 94561
rect 542154 94325 542196 94561
rect 541876 87561 542196 94325
rect 541876 87325 541918 87561
rect 542154 87325 542196 87561
rect 541876 80561 542196 87325
rect 541876 80325 541918 80561
rect 542154 80325 542196 80561
rect 541876 73561 542196 80325
rect 541876 73325 541918 73561
rect 542154 73325 542196 73561
rect 541876 66561 542196 73325
rect 541876 66325 541918 66561
rect 542154 66325 542196 66561
rect 541876 59561 542196 66325
rect 541876 59325 541918 59561
rect 542154 59325 542196 59561
rect 541876 52561 542196 59325
rect 541876 52325 541918 52561
rect 542154 52325 542196 52561
rect 541876 45561 542196 52325
rect 541876 45325 541918 45561
rect 542154 45325 542196 45561
rect 541876 38561 542196 45325
rect 541876 38325 541918 38561
rect 542154 38325 542196 38561
rect 541876 31561 542196 38325
rect 541876 31325 541918 31561
rect 542154 31325 542196 31561
rect 541876 24561 542196 31325
rect 541876 24325 541918 24561
rect 542154 24325 542196 24561
rect 541876 17561 542196 24325
rect 541876 17325 541918 17561
rect 542154 17325 542196 17561
rect 541876 10561 542196 17325
rect 541876 10325 541918 10561
rect 542154 10325 542196 10561
rect 541876 3561 542196 10325
rect 541876 3325 541918 3561
rect 542154 3325 542196 3561
rect 541876 -1706 542196 3325
rect 541876 -1942 541918 -1706
rect 542154 -1942 542196 -1706
rect 541876 -2026 542196 -1942
rect 541876 -2262 541918 -2026
rect 542154 -2262 542196 -2026
rect 541876 -2294 542196 -2262
rect 547144 705238 547464 706230
rect 547144 705002 547186 705238
rect 547422 705002 547464 705238
rect 547144 704918 547464 705002
rect 547144 704682 547186 704918
rect 547422 704682 547464 704918
rect 547144 695494 547464 704682
rect 547144 695258 547186 695494
rect 547422 695258 547464 695494
rect 547144 688494 547464 695258
rect 547144 688258 547186 688494
rect 547422 688258 547464 688494
rect 547144 681494 547464 688258
rect 547144 681258 547186 681494
rect 547422 681258 547464 681494
rect 547144 674494 547464 681258
rect 547144 674258 547186 674494
rect 547422 674258 547464 674494
rect 547144 667494 547464 674258
rect 547144 667258 547186 667494
rect 547422 667258 547464 667494
rect 547144 660494 547464 667258
rect 547144 660258 547186 660494
rect 547422 660258 547464 660494
rect 547144 653494 547464 660258
rect 547144 653258 547186 653494
rect 547422 653258 547464 653494
rect 547144 646494 547464 653258
rect 547144 646258 547186 646494
rect 547422 646258 547464 646494
rect 547144 639494 547464 646258
rect 547144 639258 547186 639494
rect 547422 639258 547464 639494
rect 547144 632494 547464 639258
rect 547144 632258 547186 632494
rect 547422 632258 547464 632494
rect 547144 625494 547464 632258
rect 547144 625258 547186 625494
rect 547422 625258 547464 625494
rect 547144 618494 547464 625258
rect 547144 618258 547186 618494
rect 547422 618258 547464 618494
rect 547144 611494 547464 618258
rect 547144 611258 547186 611494
rect 547422 611258 547464 611494
rect 547144 604494 547464 611258
rect 547144 604258 547186 604494
rect 547422 604258 547464 604494
rect 547144 597494 547464 604258
rect 547144 597258 547186 597494
rect 547422 597258 547464 597494
rect 547144 590494 547464 597258
rect 547144 590258 547186 590494
rect 547422 590258 547464 590494
rect 547144 583494 547464 590258
rect 547144 583258 547186 583494
rect 547422 583258 547464 583494
rect 547144 576494 547464 583258
rect 547144 576258 547186 576494
rect 547422 576258 547464 576494
rect 547144 569494 547464 576258
rect 547144 569258 547186 569494
rect 547422 569258 547464 569494
rect 547144 562494 547464 569258
rect 547144 562258 547186 562494
rect 547422 562258 547464 562494
rect 547144 555494 547464 562258
rect 547144 555258 547186 555494
rect 547422 555258 547464 555494
rect 547144 548494 547464 555258
rect 547144 548258 547186 548494
rect 547422 548258 547464 548494
rect 547144 541494 547464 548258
rect 547144 541258 547186 541494
rect 547422 541258 547464 541494
rect 547144 534494 547464 541258
rect 547144 534258 547186 534494
rect 547422 534258 547464 534494
rect 547144 527494 547464 534258
rect 547144 527258 547186 527494
rect 547422 527258 547464 527494
rect 547144 520494 547464 527258
rect 547144 520258 547186 520494
rect 547422 520258 547464 520494
rect 547144 513494 547464 520258
rect 547144 513258 547186 513494
rect 547422 513258 547464 513494
rect 547144 506494 547464 513258
rect 547144 506258 547186 506494
rect 547422 506258 547464 506494
rect 547144 499494 547464 506258
rect 547144 499258 547186 499494
rect 547422 499258 547464 499494
rect 547144 492494 547464 499258
rect 547144 492258 547186 492494
rect 547422 492258 547464 492494
rect 547144 485494 547464 492258
rect 547144 485258 547186 485494
rect 547422 485258 547464 485494
rect 547144 478494 547464 485258
rect 547144 478258 547186 478494
rect 547422 478258 547464 478494
rect 547144 471494 547464 478258
rect 547144 471258 547186 471494
rect 547422 471258 547464 471494
rect 547144 464494 547464 471258
rect 547144 464258 547186 464494
rect 547422 464258 547464 464494
rect 547144 457494 547464 464258
rect 547144 457258 547186 457494
rect 547422 457258 547464 457494
rect 547144 450494 547464 457258
rect 547144 450258 547186 450494
rect 547422 450258 547464 450494
rect 547144 443494 547464 450258
rect 547144 443258 547186 443494
rect 547422 443258 547464 443494
rect 547144 436494 547464 443258
rect 547144 436258 547186 436494
rect 547422 436258 547464 436494
rect 547144 429494 547464 436258
rect 547144 429258 547186 429494
rect 547422 429258 547464 429494
rect 547144 422494 547464 429258
rect 547144 422258 547186 422494
rect 547422 422258 547464 422494
rect 547144 415494 547464 422258
rect 547144 415258 547186 415494
rect 547422 415258 547464 415494
rect 547144 408494 547464 415258
rect 547144 408258 547186 408494
rect 547422 408258 547464 408494
rect 547144 401494 547464 408258
rect 547144 401258 547186 401494
rect 547422 401258 547464 401494
rect 547144 394494 547464 401258
rect 547144 394258 547186 394494
rect 547422 394258 547464 394494
rect 547144 387494 547464 394258
rect 547144 387258 547186 387494
rect 547422 387258 547464 387494
rect 547144 380494 547464 387258
rect 547144 380258 547186 380494
rect 547422 380258 547464 380494
rect 547144 373494 547464 380258
rect 547144 373258 547186 373494
rect 547422 373258 547464 373494
rect 547144 366494 547464 373258
rect 547144 366258 547186 366494
rect 547422 366258 547464 366494
rect 547144 359494 547464 366258
rect 547144 359258 547186 359494
rect 547422 359258 547464 359494
rect 547144 352494 547464 359258
rect 547144 352258 547186 352494
rect 547422 352258 547464 352494
rect 547144 345494 547464 352258
rect 547144 345258 547186 345494
rect 547422 345258 547464 345494
rect 547144 338494 547464 345258
rect 547144 338258 547186 338494
rect 547422 338258 547464 338494
rect 547144 331494 547464 338258
rect 547144 331258 547186 331494
rect 547422 331258 547464 331494
rect 547144 324494 547464 331258
rect 547144 324258 547186 324494
rect 547422 324258 547464 324494
rect 547144 317494 547464 324258
rect 547144 317258 547186 317494
rect 547422 317258 547464 317494
rect 547144 310494 547464 317258
rect 547144 310258 547186 310494
rect 547422 310258 547464 310494
rect 547144 303494 547464 310258
rect 547144 303258 547186 303494
rect 547422 303258 547464 303494
rect 547144 296494 547464 303258
rect 547144 296258 547186 296494
rect 547422 296258 547464 296494
rect 547144 289494 547464 296258
rect 547144 289258 547186 289494
rect 547422 289258 547464 289494
rect 547144 282494 547464 289258
rect 547144 282258 547186 282494
rect 547422 282258 547464 282494
rect 547144 275494 547464 282258
rect 547144 275258 547186 275494
rect 547422 275258 547464 275494
rect 547144 268494 547464 275258
rect 547144 268258 547186 268494
rect 547422 268258 547464 268494
rect 547144 261494 547464 268258
rect 547144 261258 547186 261494
rect 547422 261258 547464 261494
rect 547144 254494 547464 261258
rect 547144 254258 547186 254494
rect 547422 254258 547464 254494
rect 547144 247494 547464 254258
rect 547144 247258 547186 247494
rect 547422 247258 547464 247494
rect 547144 240494 547464 247258
rect 547144 240258 547186 240494
rect 547422 240258 547464 240494
rect 547144 233494 547464 240258
rect 547144 233258 547186 233494
rect 547422 233258 547464 233494
rect 547144 226494 547464 233258
rect 547144 226258 547186 226494
rect 547422 226258 547464 226494
rect 547144 219494 547464 226258
rect 547144 219258 547186 219494
rect 547422 219258 547464 219494
rect 547144 212494 547464 219258
rect 547144 212258 547186 212494
rect 547422 212258 547464 212494
rect 547144 205494 547464 212258
rect 547144 205258 547186 205494
rect 547422 205258 547464 205494
rect 547144 198494 547464 205258
rect 547144 198258 547186 198494
rect 547422 198258 547464 198494
rect 547144 191494 547464 198258
rect 547144 191258 547186 191494
rect 547422 191258 547464 191494
rect 547144 184494 547464 191258
rect 547144 184258 547186 184494
rect 547422 184258 547464 184494
rect 547144 177494 547464 184258
rect 547144 177258 547186 177494
rect 547422 177258 547464 177494
rect 547144 170494 547464 177258
rect 547144 170258 547186 170494
rect 547422 170258 547464 170494
rect 547144 163494 547464 170258
rect 547144 163258 547186 163494
rect 547422 163258 547464 163494
rect 547144 156494 547464 163258
rect 547144 156258 547186 156494
rect 547422 156258 547464 156494
rect 547144 149494 547464 156258
rect 547144 149258 547186 149494
rect 547422 149258 547464 149494
rect 547144 142494 547464 149258
rect 547144 142258 547186 142494
rect 547422 142258 547464 142494
rect 547144 135494 547464 142258
rect 547144 135258 547186 135494
rect 547422 135258 547464 135494
rect 547144 128494 547464 135258
rect 547144 128258 547186 128494
rect 547422 128258 547464 128494
rect 547144 121494 547464 128258
rect 547144 121258 547186 121494
rect 547422 121258 547464 121494
rect 547144 114494 547464 121258
rect 547144 114258 547186 114494
rect 547422 114258 547464 114494
rect 547144 107494 547464 114258
rect 547144 107258 547186 107494
rect 547422 107258 547464 107494
rect 547144 100494 547464 107258
rect 547144 100258 547186 100494
rect 547422 100258 547464 100494
rect 547144 93494 547464 100258
rect 547144 93258 547186 93494
rect 547422 93258 547464 93494
rect 547144 86494 547464 93258
rect 547144 86258 547186 86494
rect 547422 86258 547464 86494
rect 547144 79494 547464 86258
rect 547144 79258 547186 79494
rect 547422 79258 547464 79494
rect 547144 72494 547464 79258
rect 547144 72258 547186 72494
rect 547422 72258 547464 72494
rect 547144 65494 547464 72258
rect 547144 65258 547186 65494
rect 547422 65258 547464 65494
rect 547144 58494 547464 65258
rect 547144 58258 547186 58494
rect 547422 58258 547464 58494
rect 547144 51494 547464 58258
rect 547144 51258 547186 51494
rect 547422 51258 547464 51494
rect 547144 44494 547464 51258
rect 547144 44258 547186 44494
rect 547422 44258 547464 44494
rect 547144 37494 547464 44258
rect 547144 37258 547186 37494
rect 547422 37258 547464 37494
rect 547144 30494 547464 37258
rect 547144 30258 547186 30494
rect 547422 30258 547464 30494
rect 547144 23494 547464 30258
rect 547144 23258 547186 23494
rect 547422 23258 547464 23494
rect 547144 16494 547464 23258
rect 547144 16258 547186 16494
rect 547422 16258 547464 16494
rect 547144 9494 547464 16258
rect 547144 9258 547186 9494
rect 547422 9258 547464 9494
rect 547144 2494 547464 9258
rect 547144 2258 547186 2494
rect 547422 2258 547464 2494
rect 547144 -746 547464 2258
rect 547144 -982 547186 -746
rect 547422 -982 547464 -746
rect 547144 -1066 547464 -982
rect 547144 -1302 547186 -1066
rect 547422 -1302 547464 -1066
rect 547144 -2294 547464 -1302
rect 548876 706198 549196 706230
rect 548876 705962 548918 706198
rect 549154 705962 549196 706198
rect 548876 705878 549196 705962
rect 548876 705642 548918 705878
rect 549154 705642 549196 705878
rect 548876 696561 549196 705642
rect 548876 696325 548918 696561
rect 549154 696325 549196 696561
rect 548876 689561 549196 696325
rect 548876 689325 548918 689561
rect 549154 689325 549196 689561
rect 548876 682561 549196 689325
rect 548876 682325 548918 682561
rect 549154 682325 549196 682561
rect 548876 675561 549196 682325
rect 548876 675325 548918 675561
rect 549154 675325 549196 675561
rect 548876 668561 549196 675325
rect 548876 668325 548918 668561
rect 549154 668325 549196 668561
rect 548876 661561 549196 668325
rect 548876 661325 548918 661561
rect 549154 661325 549196 661561
rect 548876 654561 549196 661325
rect 548876 654325 548918 654561
rect 549154 654325 549196 654561
rect 548876 647561 549196 654325
rect 548876 647325 548918 647561
rect 549154 647325 549196 647561
rect 548876 640561 549196 647325
rect 548876 640325 548918 640561
rect 549154 640325 549196 640561
rect 548876 633561 549196 640325
rect 548876 633325 548918 633561
rect 549154 633325 549196 633561
rect 548876 626561 549196 633325
rect 548876 626325 548918 626561
rect 549154 626325 549196 626561
rect 548876 619561 549196 626325
rect 548876 619325 548918 619561
rect 549154 619325 549196 619561
rect 548876 612561 549196 619325
rect 548876 612325 548918 612561
rect 549154 612325 549196 612561
rect 548876 605561 549196 612325
rect 548876 605325 548918 605561
rect 549154 605325 549196 605561
rect 548876 598561 549196 605325
rect 548876 598325 548918 598561
rect 549154 598325 549196 598561
rect 548876 591561 549196 598325
rect 548876 591325 548918 591561
rect 549154 591325 549196 591561
rect 548876 584561 549196 591325
rect 548876 584325 548918 584561
rect 549154 584325 549196 584561
rect 548876 577561 549196 584325
rect 548876 577325 548918 577561
rect 549154 577325 549196 577561
rect 548876 570561 549196 577325
rect 548876 570325 548918 570561
rect 549154 570325 549196 570561
rect 548876 563561 549196 570325
rect 548876 563325 548918 563561
rect 549154 563325 549196 563561
rect 548876 556561 549196 563325
rect 548876 556325 548918 556561
rect 549154 556325 549196 556561
rect 548876 549561 549196 556325
rect 548876 549325 548918 549561
rect 549154 549325 549196 549561
rect 548876 542561 549196 549325
rect 548876 542325 548918 542561
rect 549154 542325 549196 542561
rect 548876 535561 549196 542325
rect 548876 535325 548918 535561
rect 549154 535325 549196 535561
rect 548876 528561 549196 535325
rect 548876 528325 548918 528561
rect 549154 528325 549196 528561
rect 548876 521561 549196 528325
rect 548876 521325 548918 521561
rect 549154 521325 549196 521561
rect 548876 514561 549196 521325
rect 548876 514325 548918 514561
rect 549154 514325 549196 514561
rect 548876 507561 549196 514325
rect 548876 507325 548918 507561
rect 549154 507325 549196 507561
rect 548876 500561 549196 507325
rect 548876 500325 548918 500561
rect 549154 500325 549196 500561
rect 548876 493561 549196 500325
rect 548876 493325 548918 493561
rect 549154 493325 549196 493561
rect 548876 486561 549196 493325
rect 548876 486325 548918 486561
rect 549154 486325 549196 486561
rect 548876 479561 549196 486325
rect 548876 479325 548918 479561
rect 549154 479325 549196 479561
rect 548876 472561 549196 479325
rect 548876 472325 548918 472561
rect 549154 472325 549196 472561
rect 548876 465561 549196 472325
rect 548876 465325 548918 465561
rect 549154 465325 549196 465561
rect 548876 458561 549196 465325
rect 548876 458325 548918 458561
rect 549154 458325 549196 458561
rect 548876 451561 549196 458325
rect 548876 451325 548918 451561
rect 549154 451325 549196 451561
rect 548876 444561 549196 451325
rect 548876 444325 548918 444561
rect 549154 444325 549196 444561
rect 548876 437561 549196 444325
rect 548876 437325 548918 437561
rect 549154 437325 549196 437561
rect 548876 430561 549196 437325
rect 548876 430325 548918 430561
rect 549154 430325 549196 430561
rect 548876 423561 549196 430325
rect 548876 423325 548918 423561
rect 549154 423325 549196 423561
rect 548876 416561 549196 423325
rect 548876 416325 548918 416561
rect 549154 416325 549196 416561
rect 548876 409561 549196 416325
rect 548876 409325 548918 409561
rect 549154 409325 549196 409561
rect 548876 402561 549196 409325
rect 548876 402325 548918 402561
rect 549154 402325 549196 402561
rect 548876 395561 549196 402325
rect 548876 395325 548918 395561
rect 549154 395325 549196 395561
rect 548876 388561 549196 395325
rect 548876 388325 548918 388561
rect 549154 388325 549196 388561
rect 548876 381561 549196 388325
rect 548876 381325 548918 381561
rect 549154 381325 549196 381561
rect 548876 374561 549196 381325
rect 548876 374325 548918 374561
rect 549154 374325 549196 374561
rect 548876 367561 549196 374325
rect 548876 367325 548918 367561
rect 549154 367325 549196 367561
rect 548876 360561 549196 367325
rect 548876 360325 548918 360561
rect 549154 360325 549196 360561
rect 548876 353561 549196 360325
rect 548876 353325 548918 353561
rect 549154 353325 549196 353561
rect 548876 346561 549196 353325
rect 548876 346325 548918 346561
rect 549154 346325 549196 346561
rect 548876 339561 549196 346325
rect 548876 339325 548918 339561
rect 549154 339325 549196 339561
rect 548876 332561 549196 339325
rect 548876 332325 548918 332561
rect 549154 332325 549196 332561
rect 548876 325561 549196 332325
rect 548876 325325 548918 325561
rect 549154 325325 549196 325561
rect 548876 318561 549196 325325
rect 548876 318325 548918 318561
rect 549154 318325 549196 318561
rect 548876 311561 549196 318325
rect 548876 311325 548918 311561
rect 549154 311325 549196 311561
rect 548876 304561 549196 311325
rect 548876 304325 548918 304561
rect 549154 304325 549196 304561
rect 548876 297561 549196 304325
rect 548876 297325 548918 297561
rect 549154 297325 549196 297561
rect 548876 290561 549196 297325
rect 548876 290325 548918 290561
rect 549154 290325 549196 290561
rect 548876 283561 549196 290325
rect 548876 283325 548918 283561
rect 549154 283325 549196 283561
rect 548876 276561 549196 283325
rect 548876 276325 548918 276561
rect 549154 276325 549196 276561
rect 548876 269561 549196 276325
rect 548876 269325 548918 269561
rect 549154 269325 549196 269561
rect 548876 262561 549196 269325
rect 548876 262325 548918 262561
rect 549154 262325 549196 262561
rect 548876 255561 549196 262325
rect 548876 255325 548918 255561
rect 549154 255325 549196 255561
rect 548876 248561 549196 255325
rect 548876 248325 548918 248561
rect 549154 248325 549196 248561
rect 548876 241561 549196 248325
rect 548876 241325 548918 241561
rect 549154 241325 549196 241561
rect 548876 234561 549196 241325
rect 548876 234325 548918 234561
rect 549154 234325 549196 234561
rect 548876 227561 549196 234325
rect 548876 227325 548918 227561
rect 549154 227325 549196 227561
rect 548876 220561 549196 227325
rect 548876 220325 548918 220561
rect 549154 220325 549196 220561
rect 548876 213561 549196 220325
rect 548876 213325 548918 213561
rect 549154 213325 549196 213561
rect 548876 206561 549196 213325
rect 548876 206325 548918 206561
rect 549154 206325 549196 206561
rect 548876 199561 549196 206325
rect 548876 199325 548918 199561
rect 549154 199325 549196 199561
rect 548876 192561 549196 199325
rect 548876 192325 548918 192561
rect 549154 192325 549196 192561
rect 548876 185561 549196 192325
rect 548876 185325 548918 185561
rect 549154 185325 549196 185561
rect 548876 178561 549196 185325
rect 548876 178325 548918 178561
rect 549154 178325 549196 178561
rect 548876 171561 549196 178325
rect 548876 171325 548918 171561
rect 549154 171325 549196 171561
rect 548876 164561 549196 171325
rect 548876 164325 548918 164561
rect 549154 164325 549196 164561
rect 548876 157561 549196 164325
rect 548876 157325 548918 157561
rect 549154 157325 549196 157561
rect 548876 150561 549196 157325
rect 548876 150325 548918 150561
rect 549154 150325 549196 150561
rect 548876 143561 549196 150325
rect 548876 143325 548918 143561
rect 549154 143325 549196 143561
rect 548876 136561 549196 143325
rect 548876 136325 548918 136561
rect 549154 136325 549196 136561
rect 548876 129561 549196 136325
rect 548876 129325 548918 129561
rect 549154 129325 549196 129561
rect 548876 122561 549196 129325
rect 548876 122325 548918 122561
rect 549154 122325 549196 122561
rect 548876 115561 549196 122325
rect 548876 115325 548918 115561
rect 549154 115325 549196 115561
rect 548876 108561 549196 115325
rect 548876 108325 548918 108561
rect 549154 108325 549196 108561
rect 548876 101561 549196 108325
rect 548876 101325 548918 101561
rect 549154 101325 549196 101561
rect 548876 94561 549196 101325
rect 548876 94325 548918 94561
rect 549154 94325 549196 94561
rect 548876 87561 549196 94325
rect 548876 87325 548918 87561
rect 549154 87325 549196 87561
rect 548876 80561 549196 87325
rect 548876 80325 548918 80561
rect 549154 80325 549196 80561
rect 548876 73561 549196 80325
rect 548876 73325 548918 73561
rect 549154 73325 549196 73561
rect 548876 66561 549196 73325
rect 548876 66325 548918 66561
rect 549154 66325 549196 66561
rect 548876 59561 549196 66325
rect 548876 59325 548918 59561
rect 549154 59325 549196 59561
rect 548876 52561 549196 59325
rect 548876 52325 548918 52561
rect 549154 52325 549196 52561
rect 548876 45561 549196 52325
rect 548876 45325 548918 45561
rect 549154 45325 549196 45561
rect 548876 38561 549196 45325
rect 548876 38325 548918 38561
rect 549154 38325 549196 38561
rect 548876 31561 549196 38325
rect 548876 31325 548918 31561
rect 549154 31325 549196 31561
rect 548876 24561 549196 31325
rect 548876 24325 548918 24561
rect 549154 24325 549196 24561
rect 548876 17561 549196 24325
rect 548876 17325 548918 17561
rect 549154 17325 549196 17561
rect 548876 10561 549196 17325
rect 548876 10325 548918 10561
rect 549154 10325 549196 10561
rect 548876 3561 549196 10325
rect 548876 3325 548918 3561
rect 549154 3325 549196 3561
rect 548876 -1706 549196 3325
rect 548876 -1942 548918 -1706
rect 549154 -1942 549196 -1706
rect 548876 -2026 549196 -1942
rect 548876 -2262 548918 -2026
rect 549154 -2262 549196 -2026
rect 548876 -2294 549196 -2262
rect 554144 705238 554464 706230
rect 554144 705002 554186 705238
rect 554422 705002 554464 705238
rect 554144 704918 554464 705002
rect 554144 704682 554186 704918
rect 554422 704682 554464 704918
rect 554144 695494 554464 704682
rect 554144 695258 554186 695494
rect 554422 695258 554464 695494
rect 554144 688494 554464 695258
rect 554144 688258 554186 688494
rect 554422 688258 554464 688494
rect 554144 681494 554464 688258
rect 554144 681258 554186 681494
rect 554422 681258 554464 681494
rect 554144 674494 554464 681258
rect 554144 674258 554186 674494
rect 554422 674258 554464 674494
rect 554144 667494 554464 674258
rect 554144 667258 554186 667494
rect 554422 667258 554464 667494
rect 554144 660494 554464 667258
rect 554144 660258 554186 660494
rect 554422 660258 554464 660494
rect 554144 653494 554464 660258
rect 554144 653258 554186 653494
rect 554422 653258 554464 653494
rect 554144 646494 554464 653258
rect 554144 646258 554186 646494
rect 554422 646258 554464 646494
rect 554144 639494 554464 646258
rect 554144 639258 554186 639494
rect 554422 639258 554464 639494
rect 554144 632494 554464 639258
rect 554144 632258 554186 632494
rect 554422 632258 554464 632494
rect 554144 625494 554464 632258
rect 554144 625258 554186 625494
rect 554422 625258 554464 625494
rect 554144 618494 554464 625258
rect 554144 618258 554186 618494
rect 554422 618258 554464 618494
rect 554144 611494 554464 618258
rect 554144 611258 554186 611494
rect 554422 611258 554464 611494
rect 554144 604494 554464 611258
rect 554144 604258 554186 604494
rect 554422 604258 554464 604494
rect 554144 597494 554464 604258
rect 554144 597258 554186 597494
rect 554422 597258 554464 597494
rect 554144 590494 554464 597258
rect 554144 590258 554186 590494
rect 554422 590258 554464 590494
rect 554144 583494 554464 590258
rect 554144 583258 554186 583494
rect 554422 583258 554464 583494
rect 554144 576494 554464 583258
rect 554144 576258 554186 576494
rect 554422 576258 554464 576494
rect 554144 569494 554464 576258
rect 554144 569258 554186 569494
rect 554422 569258 554464 569494
rect 554144 562494 554464 569258
rect 554144 562258 554186 562494
rect 554422 562258 554464 562494
rect 554144 555494 554464 562258
rect 554144 555258 554186 555494
rect 554422 555258 554464 555494
rect 554144 548494 554464 555258
rect 554144 548258 554186 548494
rect 554422 548258 554464 548494
rect 554144 541494 554464 548258
rect 554144 541258 554186 541494
rect 554422 541258 554464 541494
rect 554144 534494 554464 541258
rect 554144 534258 554186 534494
rect 554422 534258 554464 534494
rect 554144 527494 554464 534258
rect 554144 527258 554186 527494
rect 554422 527258 554464 527494
rect 554144 520494 554464 527258
rect 554144 520258 554186 520494
rect 554422 520258 554464 520494
rect 554144 513494 554464 520258
rect 554144 513258 554186 513494
rect 554422 513258 554464 513494
rect 554144 506494 554464 513258
rect 554144 506258 554186 506494
rect 554422 506258 554464 506494
rect 554144 499494 554464 506258
rect 554144 499258 554186 499494
rect 554422 499258 554464 499494
rect 554144 492494 554464 499258
rect 554144 492258 554186 492494
rect 554422 492258 554464 492494
rect 554144 485494 554464 492258
rect 554144 485258 554186 485494
rect 554422 485258 554464 485494
rect 554144 478494 554464 485258
rect 554144 478258 554186 478494
rect 554422 478258 554464 478494
rect 554144 471494 554464 478258
rect 554144 471258 554186 471494
rect 554422 471258 554464 471494
rect 554144 464494 554464 471258
rect 554144 464258 554186 464494
rect 554422 464258 554464 464494
rect 554144 457494 554464 464258
rect 554144 457258 554186 457494
rect 554422 457258 554464 457494
rect 554144 450494 554464 457258
rect 554144 450258 554186 450494
rect 554422 450258 554464 450494
rect 554144 443494 554464 450258
rect 554144 443258 554186 443494
rect 554422 443258 554464 443494
rect 554144 436494 554464 443258
rect 554144 436258 554186 436494
rect 554422 436258 554464 436494
rect 554144 429494 554464 436258
rect 554144 429258 554186 429494
rect 554422 429258 554464 429494
rect 554144 422494 554464 429258
rect 554144 422258 554186 422494
rect 554422 422258 554464 422494
rect 554144 415494 554464 422258
rect 554144 415258 554186 415494
rect 554422 415258 554464 415494
rect 554144 408494 554464 415258
rect 554144 408258 554186 408494
rect 554422 408258 554464 408494
rect 554144 401494 554464 408258
rect 554144 401258 554186 401494
rect 554422 401258 554464 401494
rect 554144 394494 554464 401258
rect 554144 394258 554186 394494
rect 554422 394258 554464 394494
rect 554144 387494 554464 394258
rect 554144 387258 554186 387494
rect 554422 387258 554464 387494
rect 554144 380494 554464 387258
rect 554144 380258 554186 380494
rect 554422 380258 554464 380494
rect 554144 373494 554464 380258
rect 554144 373258 554186 373494
rect 554422 373258 554464 373494
rect 554144 366494 554464 373258
rect 554144 366258 554186 366494
rect 554422 366258 554464 366494
rect 554144 359494 554464 366258
rect 554144 359258 554186 359494
rect 554422 359258 554464 359494
rect 554144 352494 554464 359258
rect 554144 352258 554186 352494
rect 554422 352258 554464 352494
rect 554144 345494 554464 352258
rect 554144 345258 554186 345494
rect 554422 345258 554464 345494
rect 554144 338494 554464 345258
rect 554144 338258 554186 338494
rect 554422 338258 554464 338494
rect 554144 331494 554464 338258
rect 554144 331258 554186 331494
rect 554422 331258 554464 331494
rect 554144 324494 554464 331258
rect 554144 324258 554186 324494
rect 554422 324258 554464 324494
rect 554144 317494 554464 324258
rect 554144 317258 554186 317494
rect 554422 317258 554464 317494
rect 554144 310494 554464 317258
rect 554144 310258 554186 310494
rect 554422 310258 554464 310494
rect 554144 303494 554464 310258
rect 554144 303258 554186 303494
rect 554422 303258 554464 303494
rect 554144 296494 554464 303258
rect 554144 296258 554186 296494
rect 554422 296258 554464 296494
rect 554144 289494 554464 296258
rect 554144 289258 554186 289494
rect 554422 289258 554464 289494
rect 554144 282494 554464 289258
rect 554144 282258 554186 282494
rect 554422 282258 554464 282494
rect 554144 275494 554464 282258
rect 554144 275258 554186 275494
rect 554422 275258 554464 275494
rect 554144 268494 554464 275258
rect 554144 268258 554186 268494
rect 554422 268258 554464 268494
rect 554144 261494 554464 268258
rect 554144 261258 554186 261494
rect 554422 261258 554464 261494
rect 554144 254494 554464 261258
rect 554144 254258 554186 254494
rect 554422 254258 554464 254494
rect 554144 247494 554464 254258
rect 554144 247258 554186 247494
rect 554422 247258 554464 247494
rect 554144 240494 554464 247258
rect 554144 240258 554186 240494
rect 554422 240258 554464 240494
rect 554144 233494 554464 240258
rect 554144 233258 554186 233494
rect 554422 233258 554464 233494
rect 554144 226494 554464 233258
rect 554144 226258 554186 226494
rect 554422 226258 554464 226494
rect 554144 219494 554464 226258
rect 554144 219258 554186 219494
rect 554422 219258 554464 219494
rect 554144 212494 554464 219258
rect 554144 212258 554186 212494
rect 554422 212258 554464 212494
rect 554144 205494 554464 212258
rect 554144 205258 554186 205494
rect 554422 205258 554464 205494
rect 554144 198494 554464 205258
rect 554144 198258 554186 198494
rect 554422 198258 554464 198494
rect 554144 191494 554464 198258
rect 554144 191258 554186 191494
rect 554422 191258 554464 191494
rect 554144 184494 554464 191258
rect 554144 184258 554186 184494
rect 554422 184258 554464 184494
rect 554144 177494 554464 184258
rect 554144 177258 554186 177494
rect 554422 177258 554464 177494
rect 554144 170494 554464 177258
rect 554144 170258 554186 170494
rect 554422 170258 554464 170494
rect 554144 163494 554464 170258
rect 554144 163258 554186 163494
rect 554422 163258 554464 163494
rect 554144 156494 554464 163258
rect 554144 156258 554186 156494
rect 554422 156258 554464 156494
rect 554144 149494 554464 156258
rect 554144 149258 554186 149494
rect 554422 149258 554464 149494
rect 554144 142494 554464 149258
rect 554144 142258 554186 142494
rect 554422 142258 554464 142494
rect 554144 135494 554464 142258
rect 554144 135258 554186 135494
rect 554422 135258 554464 135494
rect 554144 128494 554464 135258
rect 554144 128258 554186 128494
rect 554422 128258 554464 128494
rect 554144 121494 554464 128258
rect 554144 121258 554186 121494
rect 554422 121258 554464 121494
rect 554144 114494 554464 121258
rect 554144 114258 554186 114494
rect 554422 114258 554464 114494
rect 554144 107494 554464 114258
rect 554144 107258 554186 107494
rect 554422 107258 554464 107494
rect 554144 100494 554464 107258
rect 554144 100258 554186 100494
rect 554422 100258 554464 100494
rect 554144 93494 554464 100258
rect 554144 93258 554186 93494
rect 554422 93258 554464 93494
rect 554144 86494 554464 93258
rect 554144 86258 554186 86494
rect 554422 86258 554464 86494
rect 554144 79494 554464 86258
rect 554144 79258 554186 79494
rect 554422 79258 554464 79494
rect 554144 72494 554464 79258
rect 554144 72258 554186 72494
rect 554422 72258 554464 72494
rect 554144 65494 554464 72258
rect 554144 65258 554186 65494
rect 554422 65258 554464 65494
rect 554144 58494 554464 65258
rect 554144 58258 554186 58494
rect 554422 58258 554464 58494
rect 554144 51494 554464 58258
rect 554144 51258 554186 51494
rect 554422 51258 554464 51494
rect 554144 44494 554464 51258
rect 554144 44258 554186 44494
rect 554422 44258 554464 44494
rect 554144 37494 554464 44258
rect 554144 37258 554186 37494
rect 554422 37258 554464 37494
rect 554144 30494 554464 37258
rect 554144 30258 554186 30494
rect 554422 30258 554464 30494
rect 554144 23494 554464 30258
rect 554144 23258 554186 23494
rect 554422 23258 554464 23494
rect 554144 16494 554464 23258
rect 554144 16258 554186 16494
rect 554422 16258 554464 16494
rect 554144 9494 554464 16258
rect 554144 9258 554186 9494
rect 554422 9258 554464 9494
rect 554144 2494 554464 9258
rect 554144 2258 554186 2494
rect 554422 2258 554464 2494
rect 554144 -746 554464 2258
rect 554144 -982 554186 -746
rect 554422 -982 554464 -746
rect 554144 -1066 554464 -982
rect 554144 -1302 554186 -1066
rect 554422 -1302 554464 -1066
rect 554144 -2294 554464 -1302
rect 555876 706198 556196 706230
rect 555876 705962 555918 706198
rect 556154 705962 556196 706198
rect 555876 705878 556196 705962
rect 555876 705642 555918 705878
rect 556154 705642 556196 705878
rect 555876 696561 556196 705642
rect 555876 696325 555918 696561
rect 556154 696325 556196 696561
rect 555876 689561 556196 696325
rect 555876 689325 555918 689561
rect 556154 689325 556196 689561
rect 555876 682561 556196 689325
rect 555876 682325 555918 682561
rect 556154 682325 556196 682561
rect 555876 675561 556196 682325
rect 555876 675325 555918 675561
rect 556154 675325 556196 675561
rect 555876 668561 556196 675325
rect 555876 668325 555918 668561
rect 556154 668325 556196 668561
rect 555876 661561 556196 668325
rect 555876 661325 555918 661561
rect 556154 661325 556196 661561
rect 555876 654561 556196 661325
rect 555876 654325 555918 654561
rect 556154 654325 556196 654561
rect 555876 647561 556196 654325
rect 555876 647325 555918 647561
rect 556154 647325 556196 647561
rect 555876 640561 556196 647325
rect 555876 640325 555918 640561
rect 556154 640325 556196 640561
rect 555876 633561 556196 640325
rect 555876 633325 555918 633561
rect 556154 633325 556196 633561
rect 555876 626561 556196 633325
rect 555876 626325 555918 626561
rect 556154 626325 556196 626561
rect 555876 619561 556196 626325
rect 555876 619325 555918 619561
rect 556154 619325 556196 619561
rect 555876 612561 556196 619325
rect 555876 612325 555918 612561
rect 556154 612325 556196 612561
rect 555876 605561 556196 612325
rect 555876 605325 555918 605561
rect 556154 605325 556196 605561
rect 555876 598561 556196 605325
rect 555876 598325 555918 598561
rect 556154 598325 556196 598561
rect 555876 591561 556196 598325
rect 555876 591325 555918 591561
rect 556154 591325 556196 591561
rect 555876 584561 556196 591325
rect 555876 584325 555918 584561
rect 556154 584325 556196 584561
rect 555876 577561 556196 584325
rect 555876 577325 555918 577561
rect 556154 577325 556196 577561
rect 555876 570561 556196 577325
rect 555876 570325 555918 570561
rect 556154 570325 556196 570561
rect 555876 563561 556196 570325
rect 555876 563325 555918 563561
rect 556154 563325 556196 563561
rect 555876 556561 556196 563325
rect 555876 556325 555918 556561
rect 556154 556325 556196 556561
rect 555876 549561 556196 556325
rect 555876 549325 555918 549561
rect 556154 549325 556196 549561
rect 555876 542561 556196 549325
rect 555876 542325 555918 542561
rect 556154 542325 556196 542561
rect 555876 535561 556196 542325
rect 555876 535325 555918 535561
rect 556154 535325 556196 535561
rect 555876 528561 556196 535325
rect 555876 528325 555918 528561
rect 556154 528325 556196 528561
rect 555876 521561 556196 528325
rect 555876 521325 555918 521561
rect 556154 521325 556196 521561
rect 555876 514561 556196 521325
rect 555876 514325 555918 514561
rect 556154 514325 556196 514561
rect 555876 507561 556196 514325
rect 555876 507325 555918 507561
rect 556154 507325 556196 507561
rect 555876 500561 556196 507325
rect 555876 500325 555918 500561
rect 556154 500325 556196 500561
rect 555876 493561 556196 500325
rect 555876 493325 555918 493561
rect 556154 493325 556196 493561
rect 555876 486561 556196 493325
rect 555876 486325 555918 486561
rect 556154 486325 556196 486561
rect 555876 479561 556196 486325
rect 555876 479325 555918 479561
rect 556154 479325 556196 479561
rect 555876 472561 556196 479325
rect 555876 472325 555918 472561
rect 556154 472325 556196 472561
rect 555876 465561 556196 472325
rect 555876 465325 555918 465561
rect 556154 465325 556196 465561
rect 555876 458561 556196 465325
rect 555876 458325 555918 458561
rect 556154 458325 556196 458561
rect 555876 451561 556196 458325
rect 555876 451325 555918 451561
rect 556154 451325 556196 451561
rect 555876 444561 556196 451325
rect 555876 444325 555918 444561
rect 556154 444325 556196 444561
rect 555876 437561 556196 444325
rect 555876 437325 555918 437561
rect 556154 437325 556196 437561
rect 555876 430561 556196 437325
rect 555876 430325 555918 430561
rect 556154 430325 556196 430561
rect 555876 423561 556196 430325
rect 555876 423325 555918 423561
rect 556154 423325 556196 423561
rect 555876 416561 556196 423325
rect 555876 416325 555918 416561
rect 556154 416325 556196 416561
rect 555876 409561 556196 416325
rect 555876 409325 555918 409561
rect 556154 409325 556196 409561
rect 555876 402561 556196 409325
rect 555876 402325 555918 402561
rect 556154 402325 556196 402561
rect 555876 395561 556196 402325
rect 555876 395325 555918 395561
rect 556154 395325 556196 395561
rect 555876 388561 556196 395325
rect 555876 388325 555918 388561
rect 556154 388325 556196 388561
rect 555876 381561 556196 388325
rect 555876 381325 555918 381561
rect 556154 381325 556196 381561
rect 555876 374561 556196 381325
rect 555876 374325 555918 374561
rect 556154 374325 556196 374561
rect 555876 367561 556196 374325
rect 555876 367325 555918 367561
rect 556154 367325 556196 367561
rect 555876 360561 556196 367325
rect 555876 360325 555918 360561
rect 556154 360325 556196 360561
rect 555876 353561 556196 360325
rect 555876 353325 555918 353561
rect 556154 353325 556196 353561
rect 555876 346561 556196 353325
rect 555876 346325 555918 346561
rect 556154 346325 556196 346561
rect 555876 339561 556196 346325
rect 555876 339325 555918 339561
rect 556154 339325 556196 339561
rect 555876 332561 556196 339325
rect 555876 332325 555918 332561
rect 556154 332325 556196 332561
rect 555876 325561 556196 332325
rect 555876 325325 555918 325561
rect 556154 325325 556196 325561
rect 555876 318561 556196 325325
rect 555876 318325 555918 318561
rect 556154 318325 556196 318561
rect 555876 311561 556196 318325
rect 555876 311325 555918 311561
rect 556154 311325 556196 311561
rect 555876 304561 556196 311325
rect 555876 304325 555918 304561
rect 556154 304325 556196 304561
rect 555876 297561 556196 304325
rect 555876 297325 555918 297561
rect 556154 297325 556196 297561
rect 555876 290561 556196 297325
rect 555876 290325 555918 290561
rect 556154 290325 556196 290561
rect 555876 283561 556196 290325
rect 555876 283325 555918 283561
rect 556154 283325 556196 283561
rect 555876 276561 556196 283325
rect 555876 276325 555918 276561
rect 556154 276325 556196 276561
rect 555876 269561 556196 276325
rect 555876 269325 555918 269561
rect 556154 269325 556196 269561
rect 555876 262561 556196 269325
rect 555876 262325 555918 262561
rect 556154 262325 556196 262561
rect 555876 255561 556196 262325
rect 555876 255325 555918 255561
rect 556154 255325 556196 255561
rect 555876 248561 556196 255325
rect 555876 248325 555918 248561
rect 556154 248325 556196 248561
rect 555876 241561 556196 248325
rect 555876 241325 555918 241561
rect 556154 241325 556196 241561
rect 555876 234561 556196 241325
rect 555876 234325 555918 234561
rect 556154 234325 556196 234561
rect 555876 227561 556196 234325
rect 555876 227325 555918 227561
rect 556154 227325 556196 227561
rect 555876 220561 556196 227325
rect 555876 220325 555918 220561
rect 556154 220325 556196 220561
rect 555876 213561 556196 220325
rect 555876 213325 555918 213561
rect 556154 213325 556196 213561
rect 555876 206561 556196 213325
rect 555876 206325 555918 206561
rect 556154 206325 556196 206561
rect 555876 199561 556196 206325
rect 555876 199325 555918 199561
rect 556154 199325 556196 199561
rect 555876 192561 556196 199325
rect 555876 192325 555918 192561
rect 556154 192325 556196 192561
rect 555876 185561 556196 192325
rect 555876 185325 555918 185561
rect 556154 185325 556196 185561
rect 555876 178561 556196 185325
rect 555876 178325 555918 178561
rect 556154 178325 556196 178561
rect 555876 171561 556196 178325
rect 555876 171325 555918 171561
rect 556154 171325 556196 171561
rect 555876 164561 556196 171325
rect 555876 164325 555918 164561
rect 556154 164325 556196 164561
rect 555876 157561 556196 164325
rect 555876 157325 555918 157561
rect 556154 157325 556196 157561
rect 555876 150561 556196 157325
rect 555876 150325 555918 150561
rect 556154 150325 556196 150561
rect 555876 143561 556196 150325
rect 555876 143325 555918 143561
rect 556154 143325 556196 143561
rect 555876 136561 556196 143325
rect 555876 136325 555918 136561
rect 556154 136325 556196 136561
rect 555876 129561 556196 136325
rect 555876 129325 555918 129561
rect 556154 129325 556196 129561
rect 555876 122561 556196 129325
rect 555876 122325 555918 122561
rect 556154 122325 556196 122561
rect 555876 115561 556196 122325
rect 555876 115325 555918 115561
rect 556154 115325 556196 115561
rect 555876 108561 556196 115325
rect 555876 108325 555918 108561
rect 556154 108325 556196 108561
rect 555876 101561 556196 108325
rect 555876 101325 555918 101561
rect 556154 101325 556196 101561
rect 555876 94561 556196 101325
rect 555876 94325 555918 94561
rect 556154 94325 556196 94561
rect 555876 87561 556196 94325
rect 555876 87325 555918 87561
rect 556154 87325 556196 87561
rect 555876 80561 556196 87325
rect 555876 80325 555918 80561
rect 556154 80325 556196 80561
rect 555876 73561 556196 80325
rect 555876 73325 555918 73561
rect 556154 73325 556196 73561
rect 555876 66561 556196 73325
rect 555876 66325 555918 66561
rect 556154 66325 556196 66561
rect 555876 59561 556196 66325
rect 555876 59325 555918 59561
rect 556154 59325 556196 59561
rect 555876 52561 556196 59325
rect 555876 52325 555918 52561
rect 556154 52325 556196 52561
rect 555876 45561 556196 52325
rect 555876 45325 555918 45561
rect 556154 45325 556196 45561
rect 555876 38561 556196 45325
rect 555876 38325 555918 38561
rect 556154 38325 556196 38561
rect 555876 31561 556196 38325
rect 555876 31325 555918 31561
rect 556154 31325 556196 31561
rect 555876 24561 556196 31325
rect 555876 24325 555918 24561
rect 556154 24325 556196 24561
rect 555876 17561 556196 24325
rect 555876 17325 555918 17561
rect 556154 17325 556196 17561
rect 555876 10561 556196 17325
rect 555876 10325 555918 10561
rect 556154 10325 556196 10561
rect 555876 3561 556196 10325
rect 555876 3325 555918 3561
rect 556154 3325 556196 3561
rect 555876 -1706 556196 3325
rect 555876 -1942 555918 -1706
rect 556154 -1942 556196 -1706
rect 555876 -2026 556196 -1942
rect 555876 -2262 555918 -2026
rect 556154 -2262 556196 -2026
rect 555876 -2294 556196 -2262
rect 561144 705238 561464 706230
rect 561144 705002 561186 705238
rect 561422 705002 561464 705238
rect 561144 704918 561464 705002
rect 561144 704682 561186 704918
rect 561422 704682 561464 704918
rect 561144 695494 561464 704682
rect 561144 695258 561186 695494
rect 561422 695258 561464 695494
rect 561144 688494 561464 695258
rect 561144 688258 561186 688494
rect 561422 688258 561464 688494
rect 561144 681494 561464 688258
rect 561144 681258 561186 681494
rect 561422 681258 561464 681494
rect 561144 674494 561464 681258
rect 561144 674258 561186 674494
rect 561422 674258 561464 674494
rect 561144 667494 561464 674258
rect 561144 667258 561186 667494
rect 561422 667258 561464 667494
rect 561144 660494 561464 667258
rect 561144 660258 561186 660494
rect 561422 660258 561464 660494
rect 561144 653494 561464 660258
rect 561144 653258 561186 653494
rect 561422 653258 561464 653494
rect 561144 646494 561464 653258
rect 561144 646258 561186 646494
rect 561422 646258 561464 646494
rect 561144 639494 561464 646258
rect 561144 639258 561186 639494
rect 561422 639258 561464 639494
rect 561144 632494 561464 639258
rect 561144 632258 561186 632494
rect 561422 632258 561464 632494
rect 561144 625494 561464 632258
rect 561144 625258 561186 625494
rect 561422 625258 561464 625494
rect 561144 618494 561464 625258
rect 561144 618258 561186 618494
rect 561422 618258 561464 618494
rect 561144 611494 561464 618258
rect 561144 611258 561186 611494
rect 561422 611258 561464 611494
rect 561144 604494 561464 611258
rect 561144 604258 561186 604494
rect 561422 604258 561464 604494
rect 561144 597494 561464 604258
rect 561144 597258 561186 597494
rect 561422 597258 561464 597494
rect 561144 590494 561464 597258
rect 561144 590258 561186 590494
rect 561422 590258 561464 590494
rect 561144 583494 561464 590258
rect 561144 583258 561186 583494
rect 561422 583258 561464 583494
rect 561144 576494 561464 583258
rect 561144 576258 561186 576494
rect 561422 576258 561464 576494
rect 561144 569494 561464 576258
rect 561144 569258 561186 569494
rect 561422 569258 561464 569494
rect 561144 562494 561464 569258
rect 561144 562258 561186 562494
rect 561422 562258 561464 562494
rect 561144 555494 561464 562258
rect 561144 555258 561186 555494
rect 561422 555258 561464 555494
rect 561144 548494 561464 555258
rect 561144 548258 561186 548494
rect 561422 548258 561464 548494
rect 561144 541494 561464 548258
rect 561144 541258 561186 541494
rect 561422 541258 561464 541494
rect 561144 534494 561464 541258
rect 561144 534258 561186 534494
rect 561422 534258 561464 534494
rect 561144 527494 561464 534258
rect 561144 527258 561186 527494
rect 561422 527258 561464 527494
rect 561144 520494 561464 527258
rect 561144 520258 561186 520494
rect 561422 520258 561464 520494
rect 561144 513494 561464 520258
rect 561144 513258 561186 513494
rect 561422 513258 561464 513494
rect 561144 506494 561464 513258
rect 561144 506258 561186 506494
rect 561422 506258 561464 506494
rect 561144 499494 561464 506258
rect 561144 499258 561186 499494
rect 561422 499258 561464 499494
rect 561144 492494 561464 499258
rect 561144 492258 561186 492494
rect 561422 492258 561464 492494
rect 561144 485494 561464 492258
rect 561144 485258 561186 485494
rect 561422 485258 561464 485494
rect 561144 478494 561464 485258
rect 561144 478258 561186 478494
rect 561422 478258 561464 478494
rect 561144 471494 561464 478258
rect 561144 471258 561186 471494
rect 561422 471258 561464 471494
rect 561144 464494 561464 471258
rect 561144 464258 561186 464494
rect 561422 464258 561464 464494
rect 561144 457494 561464 464258
rect 561144 457258 561186 457494
rect 561422 457258 561464 457494
rect 561144 450494 561464 457258
rect 561144 450258 561186 450494
rect 561422 450258 561464 450494
rect 561144 443494 561464 450258
rect 561144 443258 561186 443494
rect 561422 443258 561464 443494
rect 561144 436494 561464 443258
rect 561144 436258 561186 436494
rect 561422 436258 561464 436494
rect 561144 429494 561464 436258
rect 561144 429258 561186 429494
rect 561422 429258 561464 429494
rect 561144 422494 561464 429258
rect 561144 422258 561186 422494
rect 561422 422258 561464 422494
rect 561144 415494 561464 422258
rect 561144 415258 561186 415494
rect 561422 415258 561464 415494
rect 561144 408494 561464 415258
rect 561144 408258 561186 408494
rect 561422 408258 561464 408494
rect 561144 401494 561464 408258
rect 561144 401258 561186 401494
rect 561422 401258 561464 401494
rect 561144 394494 561464 401258
rect 561144 394258 561186 394494
rect 561422 394258 561464 394494
rect 561144 387494 561464 394258
rect 561144 387258 561186 387494
rect 561422 387258 561464 387494
rect 561144 380494 561464 387258
rect 561144 380258 561186 380494
rect 561422 380258 561464 380494
rect 561144 373494 561464 380258
rect 561144 373258 561186 373494
rect 561422 373258 561464 373494
rect 561144 366494 561464 373258
rect 561144 366258 561186 366494
rect 561422 366258 561464 366494
rect 561144 359494 561464 366258
rect 561144 359258 561186 359494
rect 561422 359258 561464 359494
rect 561144 352494 561464 359258
rect 561144 352258 561186 352494
rect 561422 352258 561464 352494
rect 561144 345494 561464 352258
rect 561144 345258 561186 345494
rect 561422 345258 561464 345494
rect 561144 338494 561464 345258
rect 561144 338258 561186 338494
rect 561422 338258 561464 338494
rect 561144 331494 561464 338258
rect 561144 331258 561186 331494
rect 561422 331258 561464 331494
rect 561144 324494 561464 331258
rect 561144 324258 561186 324494
rect 561422 324258 561464 324494
rect 561144 317494 561464 324258
rect 561144 317258 561186 317494
rect 561422 317258 561464 317494
rect 561144 310494 561464 317258
rect 561144 310258 561186 310494
rect 561422 310258 561464 310494
rect 561144 303494 561464 310258
rect 561144 303258 561186 303494
rect 561422 303258 561464 303494
rect 561144 296494 561464 303258
rect 561144 296258 561186 296494
rect 561422 296258 561464 296494
rect 561144 289494 561464 296258
rect 561144 289258 561186 289494
rect 561422 289258 561464 289494
rect 561144 282494 561464 289258
rect 561144 282258 561186 282494
rect 561422 282258 561464 282494
rect 561144 275494 561464 282258
rect 561144 275258 561186 275494
rect 561422 275258 561464 275494
rect 561144 268494 561464 275258
rect 561144 268258 561186 268494
rect 561422 268258 561464 268494
rect 561144 261494 561464 268258
rect 561144 261258 561186 261494
rect 561422 261258 561464 261494
rect 561144 254494 561464 261258
rect 561144 254258 561186 254494
rect 561422 254258 561464 254494
rect 561144 247494 561464 254258
rect 561144 247258 561186 247494
rect 561422 247258 561464 247494
rect 561144 240494 561464 247258
rect 561144 240258 561186 240494
rect 561422 240258 561464 240494
rect 561144 233494 561464 240258
rect 561144 233258 561186 233494
rect 561422 233258 561464 233494
rect 561144 226494 561464 233258
rect 561144 226258 561186 226494
rect 561422 226258 561464 226494
rect 561144 219494 561464 226258
rect 561144 219258 561186 219494
rect 561422 219258 561464 219494
rect 561144 212494 561464 219258
rect 561144 212258 561186 212494
rect 561422 212258 561464 212494
rect 561144 205494 561464 212258
rect 561144 205258 561186 205494
rect 561422 205258 561464 205494
rect 561144 198494 561464 205258
rect 561144 198258 561186 198494
rect 561422 198258 561464 198494
rect 561144 191494 561464 198258
rect 561144 191258 561186 191494
rect 561422 191258 561464 191494
rect 561144 184494 561464 191258
rect 561144 184258 561186 184494
rect 561422 184258 561464 184494
rect 561144 177494 561464 184258
rect 561144 177258 561186 177494
rect 561422 177258 561464 177494
rect 561144 170494 561464 177258
rect 561144 170258 561186 170494
rect 561422 170258 561464 170494
rect 561144 163494 561464 170258
rect 561144 163258 561186 163494
rect 561422 163258 561464 163494
rect 561144 156494 561464 163258
rect 561144 156258 561186 156494
rect 561422 156258 561464 156494
rect 561144 149494 561464 156258
rect 561144 149258 561186 149494
rect 561422 149258 561464 149494
rect 561144 142494 561464 149258
rect 561144 142258 561186 142494
rect 561422 142258 561464 142494
rect 561144 135494 561464 142258
rect 561144 135258 561186 135494
rect 561422 135258 561464 135494
rect 561144 128494 561464 135258
rect 561144 128258 561186 128494
rect 561422 128258 561464 128494
rect 561144 121494 561464 128258
rect 561144 121258 561186 121494
rect 561422 121258 561464 121494
rect 561144 114494 561464 121258
rect 561144 114258 561186 114494
rect 561422 114258 561464 114494
rect 561144 107494 561464 114258
rect 561144 107258 561186 107494
rect 561422 107258 561464 107494
rect 561144 100494 561464 107258
rect 561144 100258 561186 100494
rect 561422 100258 561464 100494
rect 561144 93494 561464 100258
rect 561144 93258 561186 93494
rect 561422 93258 561464 93494
rect 561144 86494 561464 93258
rect 561144 86258 561186 86494
rect 561422 86258 561464 86494
rect 561144 79494 561464 86258
rect 561144 79258 561186 79494
rect 561422 79258 561464 79494
rect 561144 72494 561464 79258
rect 561144 72258 561186 72494
rect 561422 72258 561464 72494
rect 561144 65494 561464 72258
rect 561144 65258 561186 65494
rect 561422 65258 561464 65494
rect 561144 58494 561464 65258
rect 561144 58258 561186 58494
rect 561422 58258 561464 58494
rect 561144 51494 561464 58258
rect 561144 51258 561186 51494
rect 561422 51258 561464 51494
rect 561144 44494 561464 51258
rect 561144 44258 561186 44494
rect 561422 44258 561464 44494
rect 561144 37494 561464 44258
rect 561144 37258 561186 37494
rect 561422 37258 561464 37494
rect 561144 30494 561464 37258
rect 561144 30258 561186 30494
rect 561422 30258 561464 30494
rect 561144 23494 561464 30258
rect 561144 23258 561186 23494
rect 561422 23258 561464 23494
rect 561144 16494 561464 23258
rect 561144 16258 561186 16494
rect 561422 16258 561464 16494
rect 561144 9494 561464 16258
rect 561144 9258 561186 9494
rect 561422 9258 561464 9494
rect 561144 2494 561464 9258
rect 561144 2258 561186 2494
rect 561422 2258 561464 2494
rect 561144 -746 561464 2258
rect 561144 -982 561186 -746
rect 561422 -982 561464 -746
rect 561144 -1066 561464 -982
rect 561144 -1302 561186 -1066
rect 561422 -1302 561464 -1066
rect 561144 -2294 561464 -1302
rect 562876 706198 563196 706230
rect 562876 705962 562918 706198
rect 563154 705962 563196 706198
rect 562876 705878 563196 705962
rect 562876 705642 562918 705878
rect 563154 705642 563196 705878
rect 562876 696561 563196 705642
rect 562876 696325 562918 696561
rect 563154 696325 563196 696561
rect 562876 689561 563196 696325
rect 562876 689325 562918 689561
rect 563154 689325 563196 689561
rect 562876 682561 563196 689325
rect 562876 682325 562918 682561
rect 563154 682325 563196 682561
rect 562876 675561 563196 682325
rect 562876 675325 562918 675561
rect 563154 675325 563196 675561
rect 562876 668561 563196 675325
rect 562876 668325 562918 668561
rect 563154 668325 563196 668561
rect 562876 661561 563196 668325
rect 562876 661325 562918 661561
rect 563154 661325 563196 661561
rect 562876 654561 563196 661325
rect 562876 654325 562918 654561
rect 563154 654325 563196 654561
rect 562876 647561 563196 654325
rect 562876 647325 562918 647561
rect 563154 647325 563196 647561
rect 562876 640561 563196 647325
rect 562876 640325 562918 640561
rect 563154 640325 563196 640561
rect 562876 633561 563196 640325
rect 562876 633325 562918 633561
rect 563154 633325 563196 633561
rect 562876 626561 563196 633325
rect 562876 626325 562918 626561
rect 563154 626325 563196 626561
rect 562876 619561 563196 626325
rect 562876 619325 562918 619561
rect 563154 619325 563196 619561
rect 562876 612561 563196 619325
rect 562876 612325 562918 612561
rect 563154 612325 563196 612561
rect 562876 605561 563196 612325
rect 562876 605325 562918 605561
rect 563154 605325 563196 605561
rect 562876 598561 563196 605325
rect 562876 598325 562918 598561
rect 563154 598325 563196 598561
rect 562876 591561 563196 598325
rect 562876 591325 562918 591561
rect 563154 591325 563196 591561
rect 562876 584561 563196 591325
rect 562876 584325 562918 584561
rect 563154 584325 563196 584561
rect 562876 577561 563196 584325
rect 562876 577325 562918 577561
rect 563154 577325 563196 577561
rect 562876 570561 563196 577325
rect 562876 570325 562918 570561
rect 563154 570325 563196 570561
rect 562876 563561 563196 570325
rect 562876 563325 562918 563561
rect 563154 563325 563196 563561
rect 562876 556561 563196 563325
rect 562876 556325 562918 556561
rect 563154 556325 563196 556561
rect 562876 549561 563196 556325
rect 562876 549325 562918 549561
rect 563154 549325 563196 549561
rect 562876 542561 563196 549325
rect 562876 542325 562918 542561
rect 563154 542325 563196 542561
rect 562876 535561 563196 542325
rect 562876 535325 562918 535561
rect 563154 535325 563196 535561
rect 562876 528561 563196 535325
rect 562876 528325 562918 528561
rect 563154 528325 563196 528561
rect 562876 521561 563196 528325
rect 562876 521325 562918 521561
rect 563154 521325 563196 521561
rect 562876 514561 563196 521325
rect 562876 514325 562918 514561
rect 563154 514325 563196 514561
rect 562876 507561 563196 514325
rect 562876 507325 562918 507561
rect 563154 507325 563196 507561
rect 562876 500561 563196 507325
rect 562876 500325 562918 500561
rect 563154 500325 563196 500561
rect 562876 493561 563196 500325
rect 562876 493325 562918 493561
rect 563154 493325 563196 493561
rect 562876 486561 563196 493325
rect 562876 486325 562918 486561
rect 563154 486325 563196 486561
rect 562876 479561 563196 486325
rect 562876 479325 562918 479561
rect 563154 479325 563196 479561
rect 562876 472561 563196 479325
rect 562876 472325 562918 472561
rect 563154 472325 563196 472561
rect 562876 465561 563196 472325
rect 562876 465325 562918 465561
rect 563154 465325 563196 465561
rect 562876 458561 563196 465325
rect 562876 458325 562918 458561
rect 563154 458325 563196 458561
rect 562876 451561 563196 458325
rect 562876 451325 562918 451561
rect 563154 451325 563196 451561
rect 562876 444561 563196 451325
rect 562876 444325 562918 444561
rect 563154 444325 563196 444561
rect 562876 437561 563196 444325
rect 562876 437325 562918 437561
rect 563154 437325 563196 437561
rect 562876 430561 563196 437325
rect 562876 430325 562918 430561
rect 563154 430325 563196 430561
rect 562876 423561 563196 430325
rect 562876 423325 562918 423561
rect 563154 423325 563196 423561
rect 562876 416561 563196 423325
rect 562876 416325 562918 416561
rect 563154 416325 563196 416561
rect 562876 409561 563196 416325
rect 562876 409325 562918 409561
rect 563154 409325 563196 409561
rect 562876 402561 563196 409325
rect 562876 402325 562918 402561
rect 563154 402325 563196 402561
rect 562876 395561 563196 402325
rect 562876 395325 562918 395561
rect 563154 395325 563196 395561
rect 562876 388561 563196 395325
rect 562876 388325 562918 388561
rect 563154 388325 563196 388561
rect 562876 381561 563196 388325
rect 562876 381325 562918 381561
rect 563154 381325 563196 381561
rect 562876 374561 563196 381325
rect 562876 374325 562918 374561
rect 563154 374325 563196 374561
rect 562876 367561 563196 374325
rect 562876 367325 562918 367561
rect 563154 367325 563196 367561
rect 562876 360561 563196 367325
rect 562876 360325 562918 360561
rect 563154 360325 563196 360561
rect 562876 353561 563196 360325
rect 562876 353325 562918 353561
rect 563154 353325 563196 353561
rect 562876 346561 563196 353325
rect 562876 346325 562918 346561
rect 563154 346325 563196 346561
rect 562876 339561 563196 346325
rect 562876 339325 562918 339561
rect 563154 339325 563196 339561
rect 562876 332561 563196 339325
rect 562876 332325 562918 332561
rect 563154 332325 563196 332561
rect 562876 325561 563196 332325
rect 562876 325325 562918 325561
rect 563154 325325 563196 325561
rect 562876 318561 563196 325325
rect 562876 318325 562918 318561
rect 563154 318325 563196 318561
rect 562876 311561 563196 318325
rect 562876 311325 562918 311561
rect 563154 311325 563196 311561
rect 562876 304561 563196 311325
rect 562876 304325 562918 304561
rect 563154 304325 563196 304561
rect 562876 297561 563196 304325
rect 562876 297325 562918 297561
rect 563154 297325 563196 297561
rect 562876 290561 563196 297325
rect 562876 290325 562918 290561
rect 563154 290325 563196 290561
rect 562876 283561 563196 290325
rect 562876 283325 562918 283561
rect 563154 283325 563196 283561
rect 562876 276561 563196 283325
rect 562876 276325 562918 276561
rect 563154 276325 563196 276561
rect 562876 269561 563196 276325
rect 562876 269325 562918 269561
rect 563154 269325 563196 269561
rect 562876 262561 563196 269325
rect 562876 262325 562918 262561
rect 563154 262325 563196 262561
rect 562876 255561 563196 262325
rect 562876 255325 562918 255561
rect 563154 255325 563196 255561
rect 562876 248561 563196 255325
rect 562876 248325 562918 248561
rect 563154 248325 563196 248561
rect 562876 241561 563196 248325
rect 562876 241325 562918 241561
rect 563154 241325 563196 241561
rect 562876 234561 563196 241325
rect 562876 234325 562918 234561
rect 563154 234325 563196 234561
rect 562876 227561 563196 234325
rect 562876 227325 562918 227561
rect 563154 227325 563196 227561
rect 562876 220561 563196 227325
rect 562876 220325 562918 220561
rect 563154 220325 563196 220561
rect 562876 213561 563196 220325
rect 562876 213325 562918 213561
rect 563154 213325 563196 213561
rect 562876 206561 563196 213325
rect 562876 206325 562918 206561
rect 563154 206325 563196 206561
rect 562876 199561 563196 206325
rect 562876 199325 562918 199561
rect 563154 199325 563196 199561
rect 562876 192561 563196 199325
rect 562876 192325 562918 192561
rect 563154 192325 563196 192561
rect 562876 185561 563196 192325
rect 562876 185325 562918 185561
rect 563154 185325 563196 185561
rect 562876 178561 563196 185325
rect 562876 178325 562918 178561
rect 563154 178325 563196 178561
rect 562876 171561 563196 178325
rect 562876 171325 562918 171561
rect 563154 171325 563196 171561
rect 562876 164561 563196 171325
rect 562876 164325 562918 164561
rect 563154 164325 563196 164561
rect 562876 157561 563196 164325
rect 562876 157325 562918 157561
rect 563154 157325 563196 157561
rect 562876 150561 563196 157325
rect 562876 150325 562918 150561
rect 563154 150325 563196 150561
rect 562876 143561 563196 150325
rect 562876 143325 562918 143561
rect 563154 143325 563196 143561
rect 562876 136561 563196 143325
rect 562876 136325 562918 136561
rect 563154 136325 563196 136561
rect 562876 129561 563196 136325
rect 562876 129325 562918 129561
rect 563154 129325 563196 129561
rect 562876 122561 563196 129325
rect 562876 122325 562918 122561
rect 563154 122325 563196 122561
rect 562876 115561 563196 122325
rect 562876 115325 562918 115561
rect 563154 115325 563196 115561
rect 562876 108561 563196 115325
rect 562876 108325 562918 108561
rect 563154 108325 563196 108561
rect 562876 101561 563196 108325
rect 562876 101325 562918 101561
rect 563154 101325 563196 101561
rect 562876 94561 563196 101325
rect 562876 94325 562918 94561
rect 563154 94325 563196 94561
rect 562876 87561 563196 94325
rect 562876 87325 562918 87561
rect 563154 87325 563196 87561
rect 562876 80561 563196 87325
rect 562876 80325 562918 80561
rect 563154 80325 563196 80561
rect 562876 73561 563196 80325
rect 562876 73325 562918 73561
rect 563154 73325 563196 73561
rect 562876 66561 563196 73325
rect 562876 66325 562918 66561
rect 563154 66325 563196 66561
rect 562876 59561 563196 66325
rect 562876 59325 562918 59561
rect 563154 59325 563196 59561
rect 562876 52561 563196 59325
rect 562876 52325 562918 52561
rect 563154 52325 563196 52561
rect 562876 45561 563196 52325
rect 562876 45325 562918 45561
rect 563154 45325 563196 45561
rect 562876 38561 563196 45325
rect 562876 38325 562918 38561
rect 563154 38325 563196 38561
rect 562876 31561 563196 38325
rect 562876 31325 562918 31561
rect 563154 31325 563196 31561
rect 562876 24561 563196 31325
rect 562876 24325 562918 24561
rect 563154 24325 563196 24561
rect 562876 17561 563196 24325
rect 562876 17325 562918 17561
rect 563154 17325 563196 17561
rect 562876 10561 563196 17325
rect 562876 10325 562918 10561
rect 563154 10325 563196 10561
rect 562876 3561 563196 10325
rect 562876 3325 562918 3561
rect 563154 3325 563196 3561
rect 562876 -1706 563196 3325
rect 562876 -1942 562918 -1706
rect 563154 -1942 563196 -1706
rect 562876 -2026 563196 -1942
rect 562876 -2262 562918 -2026
rect 563154 -2262 563196 -2026
rect 562876 -2294 563196 -2262
rect 568144 705238 568464 706230
rect 568144 705002 568186 705238
rect 568422 705002 568464 705238
rect 568144 704918 568464 705002
rect 568144 704682 568186 704918
rect 568422 704682 568464 704918
rect 568144 695494 568464 704682
rect 568144 695258 568186 695494
rect 568422 695258 568464 695494
rect 568144 688494 568464 695258
rect 568144 688258 568186 688494
rect 568422 688258 568464 688494
rect 568144 681494 568464 688258
rect 568144 681258 568186 681494
rect 568422 681258 568464 681494
rect 568144 674494 568464 681258
rect 568144 674258 568186 674494
rect 568422 674258 568464 674494
rect 568144 667494 568464 674258
rect 568144 667258 568186 667494
rect 568422 667258 568464 667494
rect 568144 660494 568464 667258
rect 568144 660258 568186 660494
rect 568422 660258 568464 660494
rect 568144 653494 568464 660258
rect 568144 653258 568186 653494
rect 568422 653258 568464 653494
rect 568144 646494 568464 653258
rect 568144 646258 568186 646494
rect 568422 646258 568464 646494
rect 568144 639494 568464 646258
rect 568144 639258 568186 639494
rect 568422 639258 568464 639494
rect 568144 632494 568464 639258
rect 568144 632258 568186 632494
rect 568422 632258 568464 632494
rect 568144 625494 568464 632258
rect 568144 625258 568186 625494
rect 568422 625258 568464 625494
rect 568144 618494 568464 625258
rect 568144 618258 568186 618494
rect 568422 618258 568464 618494
rect 568144 611494 568464 618258
rect 568144 611258 568186 611494
rect 568422 611258 568464 611494
rect 568144 604494 568464 611258
rect 568144 604258 568186 604494
rect 568422 604258 568464 604494
rect 568144 597494 568464 604258
rect 568144 597258 568186 597494
rect 568422 597258 568464 597494
rect 568144 590494 568464 597258
rect 568144 590258 568186 590494
rect 568422 590258 568464 590494
rect 568144 583494 568464 590258
rect 568144 583258 568186 583494
rect 568422 583258 568464 583494
rect 568144 576494 568464 583258
rect 568144 576258 568186 576494
rect 568422 576258 568464 576494
rect 568144 569494 568464 576258
rect 568144 569258 568186 569494
rect 568422 569258 568464 569494
rect 568144 562494 568464 569258
rect 568144 562258 568186 562494
rect 568422 562258 568464 562494
rect 568144 555494 568464 562258
rect 568144 555258 568186 555494
rect 568422 555258 568464 555494
rect 568144 548494 568464 555258
rect 568144 548258 568186 548494
rect 568422 548258 568464 548494
rect 568144 541494 568464 548258
rect 568144 541258 568186 541494
rect 568422 541258 568464 541494
rect 568144 534494 568464 541258
rect 568144 534258 568186 534494
rect 568422 534258 568464 534494
rect 568144 527494 568464 534258
rect 568144 527258 568186 527494
rect 568422 527258 568464 527494
rect 568144 520494 568464 527258
rect 568144 520258 568186 520494
rect 568422 520258 568464 520494
rect 568144 513494 568464 520258
rect 568144 513258 568186 513494
rect 568422 513258 568464 513494
rect 568144 506494 568464 513258
rect 568144 506258 568186 506494
rect 568422 506258 568464 506494
rect 568144 499494 568464 506258
rect 568144 499258 568186 499494
rect 568422 499258 568464 499494
rect 568144 492494 568464 499258
rect 568144 492258 568186 492494
rect 568422 492258 568464 492494
rect 568144 485494 568464 492258
rect 568144 485258 568186 485494
rect 568422 485258 568464 485494
rect 568144 478494 568464 485258
rect 568144 478258 568186 478494
rect 568422 478258 568464 478494
rect 568144 471494 568464 478258
rect 568144 471258 568186 471494
rect 568422 471258 568464 471494
rect 568144 464494 568464 471258
rect 568144 464258 568186 464494
rect 568422 464258 568464 464494
rect 568144 457494 568464 464258
rect 568144 457258 568186 457494
rect 568422 457258 568464 457494
rect 568144 450494 568464 457258
rect 568144 450258 568186 450494
rect 568422 450258 568464 450494
rect 568144 443494 568464 450258
rect 568144 443258 568186 443494
rect 568422 443258 568464 443494
rect 568144 436494 568464 443258
rect 568144 436258 568186 436494
rect 568422 436258 568464 436494
rect 568144 429494 568464 436258
rect 568144 429258 568186 429494
rect 568422 429258 568464 429494
rect 568144 422494 568464 429258
rect 568144 422258 568186 422494
rect 568422 422258 568464 422494
rect 568144 415494 568464 422258
rect 568144 415258 568186 415494
rect 568422 415258 568464 415494
rect 568144 408494 568464 415258
rect 568144 408258 568186 408494
rect 568422 408258 568464 408494
rect 568144 401494 568464 408258
rect 568144 401258 568186 401494
rect 568422 401258 568464 401494
rect 568144 394494 568464 401258
rect 568144 394258 568186 394494
rect 568422 394258 568464 394494
rect 568144 387494 568464 394258
rect 568144 387258 568186 387494
rect 568422 387258 568464 387494
rect 568144 380494 568464 387258
rect 568144 380258 568186 380494
rect 568422 380258 568464 380494
rect 568144 373494 568464 380258
rect 568144 373258 568186 373494
rect 568422 373258 568464 373494
rect 568144 366494 568464 373258
rect 568144 366258 568186 366494
rect 568422 366258 568464 366494
rect 568144 359494 568464 366258
rect 568144 359258 568186 359494
rect 568422 359258 568464 359494
rect 568144 352494 568464 359258
rect 568144 352258 568186 352494
rect 568422 352258 568464 352494
rect 568144 345494 568464 352258
rect 568144 345258 568186 345494
rect 568422 345258 568464 345494
rect 568144 338494 568464 345258
rect 568144 338258 568186 338494
rect 568422 338258 568464 338494
rect 568144 331494 568464 338258
rect 568144 331258 568186 331494
rect 568422 331258 568464 331494
rect 568144 324494 568464 331258
rect 568144 324258 568186 324494
rect 568422 324258 568464 324494
rect 568144 317494 568464 324258
rect 568144 317258 568186 317494
rect 568422 317258 568464 317494
rect 568144 310494 568464 317258
rect 568144 310258 568186 310494
rect 568422 310258 568464 310494
rect 568144 303494 568464 310258
rect 568144 303258 568186 303494
rect 568422 303258 568464 303494
rect 568144 296494 568464 303258
rect 568144 296258 568186 296494
rect 568422 296258 568464 296494
rect 568144 289494 568464 296258
rect 568144 289258 568186 289494
rect 568422 289258 568464 289494
rect 568144 282494 568464 289258
rect 568144 282258 568186 282494
rect 568422 282258 568464 282494
rect 568144 275494 568464 282258
rect 568144 275258 568186 275494
rect 568422 275258 568464 275494
rect 568144 268494 568464 275258
rect 568144 268258 568186 268494
rect 568422 268258 568464 268494
rect 568144 261494 568464 268258
rect 568144 261258 568186 261494
rect 568422 261258 568464 261494
rect 568144 254494 568464 261258
rect 568144 254258 568186 254494
rect 568422 254258 568464 254494
rect 568144 247494 568464 254258
rect 568144 247258 568186 247494
rect 568422 247258 568464 247494
rect 568144 240494 568464 247258
rect 568144 240258 568186 240494
rect 568422 240258 568464 240494
rect 568144 233494 568464 240258
rect 568144 233258 568186 233494
rect 568422 233258 568464 233494
rect 568144 226494 568464 233258
rect 568144 226258 568186 226494
rect 568422 226258 568464 226494
rect 568144 219494 568464 226258
rect 568144 219258 568186 219494
rect 568422 219258 568464 219494
rect 568144 212494 568464 219258
rect 568144 212258 568186 212494
rect 568422 212258 568464 212494
rect 568144 205494 568464 212258
rect 568144 205258 568186 205494
rect 568422 205258 568464 205494
rect 568144 198494 568464 205258
rect 568144 198258 568186 198494
rect 568422 198258 568464 198494
rect 568144 191494 568464 198258
rect 568144 191258 568186 191494
rect 568422 191258 568464 191494
rect 568144 184494 568464 191258
rect 568144 184258 568186 184494
rect 568422 184258 568464 184494
rect 568144 177494 568464 184258
rect 568144 177258 568186 177494
rect 568422 177258 568464 177494
rect 568144 170494 568464 177258
rect 568144 170258 568186 170494
rect 568422 170258 568464 170494
rect 568144 163494 568464 170258
rect 568144 163258 568186 163494
rect 568422 163258 568464 163494
rect 568144 156494 568464 163258
rect 568144 156258 568186 156494
rect 568422 156258 568464 156494
rect 568144 149494 568464 156258
rect 568144 149258 568186 149494
rect 568422 149258 568464 149494
rect 568144 142494 568464 149258
rect 568144 142258 568186 142494
rect 568422 142258 568464 142494
rect 568144 135494 568464 142258
rect 568144 135258 568186 135494
rect 568422 135258 568464 135494
rect 568144 128494 568464 135258
rect 568144 128258 568186 128494
rect 568422 128258 568464 128494
rect 568144 121494 568464 128258
rect 568144 121258 568186 121494
rect 568422 121258 568464 121494
rect 568144 114494 568464 121258
rect 568144 114258 568186 114494
rect 568422 114258 568464 114494
rect 568144 107494 568464 114258
rect 568144 107258 568186 107494
rect 568422 107258 568464 107494
rect 568144 100494 568464 107258
rect 568144 100258 568186 100494
rect 568422 100258 568464 100494
rect 568144 93494 568464 100258
rect 568144 93258 568186 93494
rect 568422 93258 568464 93494
rect 568144 86494 568464 93258
rect 568144 86258 568186 86494
rect 568422 86258 568464 86494
rect 568144 79494 568464 86258
rect 568144 79258 568186 79494
rect 568422 79258 568464 79494
rect 568144 72494 568464 79258
rect 568144 72258 568186 72494
rect 568422 72258 568464 72494
rect 568144 65494 568464 72258
rect 568144 65258 568186 65494
rect 568422 65258 568464 65494
rect 568144 58494 568464 65258
rect 568144 58258 568186 58494
rect 568422 58258 568464 58494
rect 568144 51494 568464 58258
rect 568144 51258 568186 51494
rect 568422 51258 568464 51494
rect 568144 44494 568464 51258
rect 568144 44258 568186 44494
rect 568422 44258 568464 44494
rect 568144 37494 568464 44258
rect 568144 37258 568186 37494
rect 568422 37258 568464 37494
rect 568144 30494 568464 37258
rect 568144 30258 568186 30494
rect 568422 30258 568464 30494
rect 568144 23494 568464 30258
rect 568144 23258 568186 23494
rect 568422 23258 568464 23494
rect 568144 16494 568464 23258
rect 568144 16258 568186 16494
rect 568422 16258 568464 16494
rect 568144 9494 568464 16258
rect 568144 9258 568186 9494
rect 568422 9258 568464 9494
rect 568144 2494 568464 9258
rect 568144 2258 568186 2494
rect 568422 2258 568464 2494
rect 568144 -746 568464 2258
rect 568144 -982 568186 -746
rect 568422 -982 568464 -746
rect 568144 -1066 568464 -982
rect 568144 -1302 568186 -1066
rect 568422 -1302 568464 -1066
rect 568144 -2294 568464 -1302
rect 569876 706198 570196 706230
rect 569876 705962 569918 706198
rect 570154 705962 570196 706198
rect 569876 705878 570196 705962
rect 569876 705642 569918 705878
rect 570154 705642 570196 705878
rect 569876 696561 570196 705642
rect 569876 696325 569918 696561
rect 570154 696325 570196 696561
rect 569876 689561 570196 696325
rect 569876 689325 569918 689561
rect 570154 689325 570196 689561
rect 569876 682561 570196 689325
rect 569876 682325 569918 682561
rect 570154 682325 570196 682561
rect 569876 675561 570196 682325
rect 569876 675325 569918 675561
rect 570154 675325 570196 675561
rect 569876 668561 570196 675325
rect 569876 668325 569918 668561
rect 570154 668325 570196 668561
rect 569876 661561 570196 668325
rect 569876 661325 569918 661561
rect 570154 661325 570196 661561
rect 569876 654561 570196 661325
rect 569876 654325 569918 654561
rect 570154 654325 570196 654561
rect 569876 647561 570196 654325
rect 569876 647325 569918 647561
rect 570154 647325 570196 647561
rect 569876 640561 570196 647325
rect 569876 640325 569918 640561
rect 570154 640325 570196 640561
rect 569876 633561 570196 640325
rect 569876 633325 569918 633561
rect 570154 633325 570196 633561
rect 569876 626561 570196 633325
rect 569876 626325 569918 626561
rect 570154 626325 570196 626561
rect 569876 619561 570196 626325
rect 569876 619325 569918 619561
rect 570154 619325 570196 619561
rect 569876 612561 570196 619325
rect 569876 612325 569918 612561
rect 570154 612325 570196 612561
rect 569876 605561 570196 612325
rect 569876 605325 569918 605561
rect 570154 605325 570196 605561
rect 569876 598561 570196 605325
rect 569876 598325 569918 598561
rect 570154 598325 570196 598561
rect 569876 591561 570196 598325
rect 569876 591325 569918 591561
rect 570154 591325 570196 591561
rect 569876 584561 570196 591325
rect 569876 584325 569918 584561
rect 570154 584325 570196 584561
rect 569876 577561 570196 584325
rect 569876 577325 569918 577561
rect 570154 577325 570196 577561
rect 569876 570561 570196 577325
rect 569876 570325 569918 570561
rect 570154 570325 570196 570561
rect 569876 563561 570196 570325
rect 569876 563325 569918 563561
rect 570154 563325 570196 563561
rect 569876 556561 570196 563325
rect 569876 556325 569918 556561
rect 570154 556325 570196 556561
rect 569876 549561 570196 556325
rect 569876 549325 569918 549561
rect 570154 549325 570196 549561
rect 569876 542561 570196 549325
rect 569876 542325 569918 542561
rect 570154 542325 570196 542561
rect 569876 535561 570196 542325
rect 569876 535325 569918 535561
rect 570154 535325 570196 535561
rect 569876 528561 570196 535325
rect 569876 528325 569918 528561
rect 570154 528325 570196 528561
rect 569876 521561 570196 528325
rect 569876 521325 569918 521561
rect 570154 521325 570196 521561
rect 569876 514561 570196 521325
rect 569876 514325 569918 514561
rect 570154 514325 570196 514561
rect 569876 507561 570196 514325
rect 569876 507325 569918 507561
rect 570154 507325 570196 507561
rect 569876 500561 570196 507325
rect 569876 500325 569918 500561
rect 570154 500325 570196 500561
rect 569876 493561 570196 500325
rect 569876 493325 569918 493561
rect 570154 493325 570196 493561
rect 569876 486561 570196 493325
rect 569876 486325 569918 486561
rect 570154 486325 570196 486561
rect 569876 479561 570196 486325
rect 569876 479325 569918 479561
rect 570154 479325 570196 479561
rect 569876 472561 570196 479325
rect 569876 472325 569918 472561
rect 570154 472325 570196 472561
rect 569876 465561 570196 472325
rect 569876 465325 569918 465561
rect 570154 465325 570196 465561
rect 569876 458561 570196 465325
rect 569876 458325 569918 458561
rect 570154 458325 570196 458561
rect 569876 451561 570196 458325
rect 569876 451325 569918 451561
rect 570154 451325 570196 451561
rect 569876 444561 570196 451325
rect 569876 444325 569918 444561
rect 570154 444325 570196 444561
rect 569876 437561 570196 444325
rect 569876 437325 569918 437561
rect 570154 437325 570196 437561
rect 569876 430561 570196 437325
rect 569876 430325 569918 430561
rect 570154 430325 570196 430561
rect 569876 423561 570196 430325
rect 569876 423325 569918 423561
rect 570154 423325 570196 423561
rect 569876 416561 570196 423325
rect 569876 416325 569918 416561
rect 570154 416325 570196 416561
rect 569876 409561 570196 416325
rect 569876 409325 569918 409561
rect 570154 409325 570196 409561
rect 569876 402561 570196 409325
rect 569876 402325 569918 402561
rect 570154 402325 570196 402561
rect 569876 395561 570196 402325
rect 569876 395325 569918 395561
rect 570154 395325 570196 395561
rect 569876 388561 570196 395325
rect 569876 388325 569918 388561
rect 570154 388325 570196 388561
rect 569876 381561 570196 388325
rect 569876 381325 569918 381561
rect 570154 381325 570196 381561
rect 569876 374561 570196 381325
rect 569876 374325 569918 374561
rect 570154 374325 570196 374561
rect 569876 367561 570196 374325
rect 569876 367325 569918 367561
rect 570154 367325 570196 367561
rect 569876 360561 570196 367325
rect 569876 360325 569918 360561
rect 570154 360325 570196 360561
rect 569876 353561 570196 360325
rect 569876 353325 569918 353561
rect 570154 353325 570196 353561
rect 569876 346561 570196 353325
rect 569876 346325 569918 346561
rect 570154 346325 570196 346561
rect 569876 339561 570196 346325
rect 569876 339325 569918 339561
rect 570154 339325 570196 339561
rect 569876 332561 570196 339325
rect 569876 332325 569918 332561
rect 570154 332325 570196 332561
rect 569876 325561 570196 332325
rect 569876 325325 569918 325561
rect 570154 325325 570196 325561
rect 569876 318561 570196 325325
rect 569876 318325 569918 318561
rect 570154 318325 570196 318561
rect 569876 311561 570196 318325
rect 569876 311325 569918 311561
rect 570154 311325 570196 311561
rect 569876 304561 570196 311325
rect 569876 304325 569918 304561
rect 570154 304325 570196 304561
rect 569876 297561 570196 304325
rect 569876 297325 569918 297561
rect 570154 297325 570196 297561
rect 569876 290561 570196 297325
rect 569876 290325 569918 290561
rect 570154 290325 570196 290561
rect 569876 283561 570196 290325
rect 569876 283325 569918 283561
rect 570154 283325 570196 283561
rect 569876 276561 570196 283325
rect 569876 276325 569918 276561
rect 570154 276325 570196 276561
rect 569876 269561 570196 276325
rect 569876 269325 569918 269561
rect 570154 269325 570196 269561
rect 569876 262561 570196 269325
rect 569876 262325 569918 262561
rect 570154 262325 570196 262561
rect 569876 255561 570196 262325
rect 569876 255325 569918 255561
rect 570154 255325 570196 255561
rect 569876 248561 570196 255325
rect 569876 248325 569918 248561
rect 570154 248325 570196 248561
rect 569876 241561 570196 248325
rect 569876 241325 569918 241561
rect 570154 241325 570196 241561
rect 569876 234561 570196 241325
rect 569876 234325 569918 234561
rect 570154 234325 570196 234561
rect 569876 227561 570196 234325
rect 569876 227325 569918 227561
rect 570154 227325 570196 227561
rect 569876 220561 570196 227325
rect 569876 220325 569918 220561
rect 570154 220325 570196 220561
rect 569876 213561 570196 220325
rect 569876 213325 569918 213561
rect 570154 213325 570196 213561
rect 569876 206561 570196 213325
rect 569876 206325 569918 206561
rect 570154 206325 570196 206561
rect 569876 199561 570196 206325
rect 569876 199325 569918 199561
rect 570154 199325 570196 199561
rect 569876 192561 570196 199325
rect 569876 192325 569918 192561
rect 570154 192325 570196 192561
rect 569876 185561 570196 192325
rect 569876 185325 569918 185561
rect 570154 185325 570196 185561
rect 569876 178561 570196 185325
rect 569876 178325 569918 178561
rect 570154 178325 570196 178561
rect 569876 171561 570196 178325
rect 569876 171325 569918 171561
rect 570154 171325 570196 171561
rect 569876 164561 570196 171325
rect 569876 164325 569918 164561
rect 570154 164325 570196 164561
rect 569876 157561 570196 164325
rect 569876 157325 569918 157561
rect 570154 157325 570196 157561
rect 569876 150561 570196 157325
rect 569876 150325 569918 150561
rect 570154 150325 570196 150561
rect 569876 143561 570196 150325
rect 569876 143325 569918 143561
rect 570154 143325 570196 143561
rect 569876 136561 570196 143325
rect 569876 136325 569918 136561
rect 570154 136325 570196 136561
rect 569876 129561 570196 136325
rect 569876 129325 569918 129561
rect 570154 129325 570196 129561
rect 569876 122561 570196 129325
rect 569876 122325 569918 122561
rect 570154 122325 570196 122561
rect 569876 115561 570196 122325
rect 569876 115325 569918 115561
rect 570154 115325 570196 115561
rect 569876 108561 570196 115325
rect 569876 108325 569918 108561
rect 570154 108325 570196 108561
rect 569876 101561 570196 108325
rect 569876 101325 569918 101561
rect 570154 101325 570196 101561
rect 569876 94561 570196 101325
rect 569876 94325 569918 94561
rect 570154 94325 570196 94561
rect 569876 87561 570196 94325
rect 569876 87325 569918 87561
rect 570154 87325 570196 87561
rect 569876 80561 570196 87325
rect 569876 80325 569918 80561
rect 570154 80325 570196 80561
rect 569876 73561 570196 80325
rect 569876 73325 569918 73561
rect 570154 73325 570196 73561
rect 569876 66561 570196 73325
rect 569876 66325 569918 66561
rect 570154 66325 570196 66561
rect 569876 59561 570196 66325
rect 569876 59325 569918 59561
rect 570154 59325 570196 59561
rect 569876 52561 570196 59325
rect 569876 52325 569918 52561
rect 570154 52325 570196 52561
rect 569876 45561 570196 52325
rect 569876 45325 569918 45561
rect 570154 45325 570196 45561
rect 569876 38561 570196 45325
rect 569876 38325 569918 38561
rect 570154 38325 570196 38561
rect 569876 31561 570196 38325
rect 569876 31325 569918 31561
rect 570154 31325 570196 31561
rect 569876 24561 570196 31325
rect 569876 24325 569918 24561
rect 570154 24325 570196 24561
rect 569876 17561 570196 24325
rect 569876 17325 569918 17561
rect 570154 17325 570196 17561
rect 569876 10561 570196 17325
rect 569876 10325 569918 10561
rect 570154 10325 570196 10561
rect 569876 3561 570196 10325
rect 569876 3325 569918 3561
rect 570154 3325 570196 3561
rect 569876 -1706 570196 3325
rect 569876 -1942 569918 -1706
rect 570154 -1942 570196 -1706
rect 569876 -2026 570196 -1942
rect 569876 -2262 569918 -2026
rect 570154 -2262 570196 -2026
rect 569876 -2294 570196 -2262
rect 575144 705238 575464 706230
rect 575144 705002 575186 705238
rect 575422 705002 575464 705238
rect 575144 704918 575464 705002
rect 575144 704682 575186 704918
rect 575422 704682 575464 704918
rect 575144 695494 575464 704682
rect 575144 695258 575186 695494
rect 575422 695258 575464 695494
rect 575144 688494 575464 695258
rect 575144 688258 575186 688494
rect 575422 688258 575464 688494
rect 575144 681494 575464 688258
rect 575144 681258 575186 681494
rect 575422 681258 575464 681494
rect 575144 674494 575464 681258
rect 575144 674258 575186 674494
rect 575422 674258 575464 674494
rect 575144 667494 575464 674258
rect 575144 667258 575186 667494
rect 575422 667258 575464 667494
rect 575144 660494 575464 667258
rect 575144 660258 575186 660494
rect 575422 660258 575464 660494
rect 575144 653494 575464 660258
rect 575144 653258 575186 653494
rect 575422 653258 575464 653494
rect 575144 646494 575464 653258
rect 575144 646258 575186 646494
rect 575422 646258 575464 646494
rect 575144 639494 575464 646258
rect 575144 639258 575186 639494
rect 575422 639258 575464 639494
rect 575144 632494 575464 639258
rect 575144 632258 575186 632494
rect 575422 632258 575464 632494
rect 575144 625494 575464 632258
rect 575144 625258 575186 625494
rect 575422 625258 575464 625494
rect 575144 618494 575464 625258
rect 575144 618258 575186 618494
rect 575422 618258 575464 618494
rect 575144 611494 575464 618258
rect 575144 611258 575186 611494
rect 575422 611258 575464 611494
rect 575144 604494 575464 611258
rect 575144 604258 575186 604494
rect 575422 604258 575464 604494
rect 575144 597494 575464 604258
rect 575144 597258 575186 597494
rect 575422 597258 575464 597494
rect 575144 590494 575464 597258
rect 575144 590258 575186 590494
rect 575422 590258 575464 590494
rect 575144 583494 575464 590258
rect 575144 583258 575186 583494
rect 575422 583258 575464 583494
rect 575144 576494 575464 583258
rect 575144 576258 575186 576494
rect 575422 576258 575464 576494
rect 575144 569494 575464 576258
rect 575144 569258 575186 569494
rect 575422 569258 575464 569494
rect 575144 562494 575464 569258
rect 575144 562258 575186 562494
rect 575422 562258 575464 562494
rect 575144 555494 575464 562258
rect 575144 555258 575186 555494
rect 575422 555258 575464 555494
rect 575144 548494 575464 555258
rect 575144 548258 575186 548494
rect 575422 548258 575464 548494
rect 575144 541494 575464 548258
rect 575144 541258 575186 541494
rect 575422 541258 575464 541494
rect 575144 534494 575464 541258
rect 575144 534258 575186 534494
rect 575422 534258 575464 534494
rect 575144 527494 575464 534258
rect 575144 527258 575186 527494
rect 575422 527258 575464 527494
rect 575144 520494 575464 527258
rect 575144 520258 575186 520494
rect 575422 520258 575464 520494
rect 575144 513494 575464 520258
rect 575144 513258 575186 513494
rect 575422 513258 575464 513494
rect 575144 506494 575464 513258
rect 575144 506258 575186 506494
rect 575422 506258 575464 506494
rect 575144 499494 575464 506258
rect 575144 499258 575186 499494
rect 575422 499258 575464 499494
rect 575144 492494 575464 499258
rect 575144 492258 575186 492494
rect 575422 492258 575464 492494
rect 575144 485494 575464 492258
rect 575144 485258 575186 485494
rect 575422 485258 575464 485494
rect 575144 478494 575464 485258
rect 575144 478258 575186 478494
rect 575422 478258 575464 478494
rect 575144 471494 575464 478258
rect 575144 471258 575186 471494
rect 575422 471258 575464 471494
rect 575144 464494 575464 471258
rect 575144 464258 575186 464494
rect 575422 464258 575464 464494
rect 575144 457494 575464 464258
rect 575144 457258 575186 457494
rect 575422 457258 575464 457494
rect 575144 450494 575464 457258
rect 575144 450258 575186 450494
rect 575422 450258 575464 450494
rect 575144 443494 575464 450258
rect 575144 443258 575186 443494
rect 575422 443258 575464 443494
rect 575144 436494 575464 443258
rect 575144 436258 575186 436494
rect 575422 436258 575464 436494
rect 575144 429494 575464 436258
rect 575144 429258 575186 429494
rect 575422 429258 575464 429494
rect 575144 422494 575464 429258
rect 575144 422258 575186 422494
rect 575422 422258 575464 422494
rect 575144 415494 575464 422258
rect 575144 415258 575186 415494
rect 575422 415258 575464 415494
rect 575144 408494 575464 415258
rect 575144 408258 575186 408494
rect 575422 408258 575464 408494
rect 575144 401494 575464 408258
rect 575144 401258 575186 401494
rect 575422 401258 575464 401494
rect 575144 394494 575464 401258
rect 575144 394258 575186 394494
rect 575422 394258 575464 394494
rect 575144 387494 575464 394258
rect 575144 387258 575186 387494
rect 575422 387258 575464 387494
rect 575144 380494 575464 387258
rect 575144 380258 575186 380494
rect 575422 380258 575464 380494
rect 575144 373494 575464 380258
rect 575144 373258 575186 373494
rect 575422 373258 575464 373494
rect 575144 366494 575464 373258
rect 575144 366258 575186 366494
rect 575422 366258 575464 366494
rect 575144 359494 575464 366258
rect 575144 359258 575186 359494
rect 575422 359258 575464 359494
rect 575144 352494 575464 359258
rect 575144 352258 575186 352494
rect 575422 352258 575464 352494
rect 575144 345494 575464 352258
rect 575144 345258 575186 345494
rect 575422 345258 575464 345494
rect 575144 338494 575464 345258
rect 575144 338258 575186 338494
rect 575422 338258 575464 338494
rect 575144 331494 575464 338258
rect 575144 331258 575186 331494
rect 575422 331258 575464 331494
rect 575144 324494 575464 331258
rect 575144 324258 575186 324494
rect 575422 324258 575464 324494
rect 575144 317494 575464 324258
rect 575144 317258 575186 317494
rect 575422 317258 575464 317494
rect 575144 310494 575464 317258
rect 575144 310258 575186 310494
rect 575422 310258 575464 310494
rect 575144 303494 575464 310258
rect 575144 303258 575186 303494
rect 575422 303258 575464 303494
rect 575144 296494 575464 303258
rect 575144 296258 575186 296494
rect 575422 296258 575464 296494
rect 575144 289494 575464 296258
rect 575144 289258 575186 289494
rect 575422 289258 575464 289494
rect 575144 282494 575464 289258
rect 575144 282258 575186 282494
rect 575422 282258 575464 282494
rect 575144 275494 575464 282258
rect 575144 275258 575186 275494
rect 575422 275258 575464 275494
rect 575144 268494 575464 275258
rect 575144 268258 575186 268494
rect 575422 268258 575464 268494
rect 575144 261494 575464 268258
rect 575144 261258 575186 261494
rect 575422 261258 575464 261494
rect 575144 254494 575464 261258
rect 575144 254258 575186 254494
rect 575422 254258 575464 254494
rect 575144 247494 575464 254258
rect 575144 247258 575186 247494
rect 575422 247258 575464 247494
rect 575144 240494 575464 247258
rect 575144 240258 575186 240494
rect 575422 240258 575464 240494
rect 575144 233494 575464 240258
rect 575144 233258 575186 233494
rect 575422 233258 575464 233494
rect 575144 226494 575464 233258
rect 575144 226258 575186 226494
rect 575422 226258 575464 226494
rect 575144 219494 575464 226258
rect 575144 219258 575186 219494
rect 575422 219258 575464 219494
rect 575144 212494 575464 219258
rect 575144 212258 575186 212494
rect 575422 212258 575464 212494
rect 575144 205494 575464 212258
rect 575144 205258 575186 205494
rect 575422 205258 575464 205494
rect 575144 198494 575464 205258
rect 575144 198258 575186 198494
rect 575422 198258 575464 198494
rect 575144 191494 575464 198258
rect 575144 191258 575186 191494
rect 575422 191258 575464 191494
rect 575144 184494 575464 191258
rect 575144 184258 575186 184494
rect 575422 184258 575464 184494
rect 575144 177494 575464 184258
rect 575144 177258 575186 177494
rect 575422 177258 575464 177494
rect 575144 170494 575464 177258
rect 575144 170258 575186 170494
rect 575422 170258 575464 170494
rect 575144 163494 575464 170258
rect 575144 163258 575186 163494
rect 575422 163258 575464 163494
rect 575144 156494 575464 163258
rect 575144 156258 575186 156494
rect 575422 156258 575464 156494
rect 575144 149494 575464 156258
rect 575144 149258 575186 149494
rect 575422 149258 575464 149494
rect 575144 142494 575464 149258
rect 575144 142258 575186 142494
rect 575422 142258 575464 142494
rect 575144 135494 575464 142258
rect 575144 135258 575186 135494
rect 575422 135258 575464 135494
rect 575144 128494 575464 135258
rect 575144 128258 575186 128494
rect 575422 128258 575464 128494
rect 575144 121494 575464 128258
rect 575144 121258 575186 121494
rect 575422 121258 575464 121494
rect 575144 114494 575464 121258
rect 575144 114258 575186 114494
rect 575422 114258 575464 114494
rect 575144 107494 575464 114258
rect 575144 107258 575186 107494
rect 575422 107258 575464 107494
rect 575144 100494 575464 107258
rect 575144 100258 575186 100494
rect 575422 100258 575464 100494
rect 575144 93494 575464 100258
rect 575144 93258 575186 93494
rect 575422 93258 575464 93494
rect 575144 86494 575464 93258
rect 575144 86258 575186 86494
rect 575422 86258 575464 86494
rect 575144 79494 575464 86258
rect 575144 79258 575186 79494
rect 575422 79258 575464 79494
rect 575144 72494 575464 79258
rect 575144 72258 575186 72494
rect 575422 72258 575464 72494
rect 575144 65494 575464 72258
rect 575144 65258 575186 65494
rect 575422 65258 575464 65494
rect 575144 58494 575464 65258
rect 575144 58258 575186 58494
rect 575422 58258 575464 58494
rect 575144 51494 575464 58258
rect 575144 51258 575186 51494
rect 575422 51258 575464 51494
rect 575144 44494 575464 51258
rect 575144 44258 575186 44494
rect 575422 44258 575464 44494
rect 575144 37494 575464 44258
rect 575144 37258 575186 37494
rect 575422 37258 575464 37494
rect 575144 30494 575464 37258
rect 575144 30258 575186 30494
rect 575422 30258 575464 30494
rect 575144 23494 575464 30258
rect 575144 23258 575186 23494
rect 575422 23258 575464 23494
rect 575144 16494 575464 23258
rect 575144 16258 575186 16494
rect 575422 16258 575464 16494
rect 575144 9494 575464 16258
rect 575144 9258 575186 9494
rect 575422 9258 575464 9494
rect 575144 2494 575464 9258
rect 575144 2258 575186 2494
rect 575422 2258 575464 2494
rect 575144 -746 575464 2258
rect 575144 -982 575186 -746
rect 575422 -982 575464 -746
rect 575144 -1066 575464 -982
rect 575144 -1302 575186 -1066
rect 575422 -1302 575464 -1066
rect 575144 -2294 575464 -1302
rect 576876 706198 577196 706230
rect 576876 705962 576918 706198
rect 577154 705962 577196 706198
rect 576876 705878 577196 705962
rect 576876 705642 576918 705878
rect 577154 705642 577196 705878
rect 576876 696561 577196 705642
rect 576876 696325 576918 696561
rect 577154 696325 577196 696561
rect 576876 689561 577196 696325
rect 576876 689325 576918 689561
rect 577154 689325 577196 689561
rect 576876 682561 577196 689325
rect 576876 682325 576918 682561
rect 577154 682325 577196 682561
rect 576876 675561 577196 682325
rect 576876 675325 576918 675561
rect 577154 675325 577196 675561
rect 576876 668561 577196 675325
rect 576876 668325 576918 668561
rect 577154 668325 577196 668561
rect 576876 661561 577196 668325
rect 576876 661325 576918 661561
rect 577154 661325 577196 661561
rect 576876 654561 577196 661325
rect 576876 654325 576918 654561
rect 577154 654325 577196 654561
rect 576876 647561 577196 654325
rect 576876 647325 576918 647561
rect 577154 647325 577196 647561
rect 576876 640561 577196 647325
rect 576876 640325 576918 640561
rect 577154 640325 577196 640561
rect 576876 633561 577196 640325
rect 576876 633325 576918 633561
rect 577154 633325 577196 633561
rect 576876 626561 577196 633325
rect 576876 626325 576918 626561
rect 577154 626325 577196 626561
rect 576876 619561 577196 626325
rect 576876 619325 576918 619561
rect 577154 619325 577196 619561
rect 576876 612561 577196 619325
rect 576876 612325 576918 612561
rect 577154 612325 577196 612561
rect 576876 605561 577196 612325
rect 576876 605325 576918 605561
rect 577154 605325 577196 605561
rect 576876 598561 577196 605325
rect 576876 598325 576918 598561
rect 577154 598325 577196 598561
rect 576876 591561 577196 598325
rect 576876 591325 576918 591561
rect 577154 591325 577196 591561
rect 576876 584561 577196 591325
rect 576876 584325 576918 584561
rect 577154 584325 577196 584561
rect 576876 577561 577196 584325
rect 576876 577325 576918 577561
rect 577154 577325 577196 577561
rect 576876 570561 577196 577325
rect 576876 570325 576918 570561
rect 577154 570325 577196 570561
rect 576876 563561 577196 570325
rect 576876 563325 576918 563561
rect 577154 563325 577196 563561
rect 576876 556561 577196 563325
rect 576876 556325 576918 556561
rect 577154 556325 577196 556561
rect 576876 549561 577196 556325
rect 576876 549325 576918 549561
rect 577154 549325 577196 549561
rect 576876 542561 577196 549325
rect 576876 542325 576918 542561
rect 577154 542325 577196 542561
rect 576876 535561 577196 542325
rect 576876 535325 576918 535561
rect 577154 535325 577196 535561
rect 576876 528561 577196 535325
rect 576876 528325 576918 528561
rect 577154 528325 577196 528561
rect 576876 521561 577196 528325
rect 576876 521325 576918 521561
rect 577154 521325 577196 521561
rect 576876 514561 577196 521325
rect 576876 514325 576918 514561
rect 577154 514325 577196 514561
rect 576876 507561 577196 514325
rect 576876 507325 576918 507561
rect 577154 507325 577196 507561
rect 576876 500561 577196 507325
rect 576876 500325 576918 500561
rect 577154 500325 577196 500561
rect 576876 493561 577196 500325
rect 576876 493325 576918 493561
rect 577154 493325 577196 493561
rect 576876 486561 577196 493325
rect 576876 486325 576918 486561
rect 577154 486325 577196 486561
rect 576876 479561 577196 486325
rect 576876 479325 576918 479561
rect 577154 479325 577196 479561
rect 576876 472561 577196 479325
rect 576876 472325 576918 472561
rect 577154 472325 577196 472561
rect 576876 465561 577196 472325
rect 576876 465325 576918 465561
rect 577154 465325 577196 465561
rect 576876 458561 577196 465325
rect 576876 458325 576918 458561
rect 577154 458325 577196 458561
rect 576876 451561 577196 458325
rect 576876 451325 576918 451561
rect 577154 451325 577196 451561
rect 576876 444561 577196 451325
rect 576876 444325 576918 444561
rect 577154 444325 577196 444561
rect 576876 437561 577196 444325
rect 576876 437325 576918 437561
rect 577154 437325 577196 437561
rect 576876 430561 577196 437325
rect 576876 430325 576918 430561
rect 577154 430325 577196 430561
rect 576876 423561 577196 430325
rect 576876 423325 576918 423561
rect 577154 423325 577196 423561
rect 576876 416561 577196 423325
rect 576876 416325 576918 416561
rect 577154 416325 577196 416561
rect 576876 409561 577196 416325
rect 576876 409325 576918 409561
rect 577154 409325 577196 409561
rect 576876 402561 577196 409325
rect 576876 402325 576918 402561
rect 577154 402325 577196 402561
rect 576876 395561 577196 402325
rect 576876 395325 576918 395561
rect 577154 395325 577196 395561
rect 576876 388561 577196 395325
rect 576876 388325 576918 388561
rect 577154 388325 577196 388561
rect 576876 381561 577196 388325
rect 576876 381325 576918 381561
rect 577154 381325 577196 381561
rect 576876 374561 577196 381325
rect 576876 374325 576918 374561
rect 577154 374325 577196 374561
rect 576876 367561 577196 374325
rect 576876 367325 576918 367561
rect 577154 367325 577196 367561
rect 576876 360561 577196 367325
rect 576876 360325 576918 360561
rect 577154 360325 577196 360561
rect 576876 353561 577196 360325
rect 576876 353325 576918 353561
rect 577154 353325 577196 353561
rect 576876 346561 577196 353325
rect 576876 346325 576918 346561
rect 577154 346325 577196 346561
rect 576876 339561 577196 346325
rect 576876 339325 576918 339561
rect 577154 339325 577196 339561
rect 576876 332561 577196 339325
rect 576876 332325 576918 332561
rect 577154 332325 577196 332561
rect 576876 325561 577196 332325
rect 576876 325325 576918 325561
rect 577154 325325 577196 325561
rect 576876 318561 577196 325325
rect 576876 318325 576918 318561
rect 577154 318325 577196 318561
rect 576876 311561 577196 318325
rect 576876 311325 576918 311561
rect 577154 311325 577196 311561
rect 576876 304561 577196 311325
rect 576876 304325 576918 304561
rect 577154 304325 577196 304561
rect 576876 297561 577196 304325
rect 576876 297325 576918 297561
rect 577154 297325 577196 297561
rect 576876 290561 577196 297325
rect 576876 290325 576918 290561
rect 577154 290325 577196 290561
rect 576876 283561 577196 290325
rect 576876 283325 576918 283561
rect 577154 283325 577196 283561
rect 576876 276561 577196 283325
rect 576876 276325 576918 276561
rect 577154 276325 577196 276561
rect 576876 269561 577196 276325
rect 576876 269325 576918 269561
rect 577154 269325 577196 269561
rect 576876 262561 577196 269325
rect 576876 262325 576918 262561
rect 577154 262325 577196 262561
rect 576876 255561 577196 262325
rect 576876 255325 576918 255561
rect 577154 255325 577196 255561
rect 576876 248561 577196 255325
rect 576876 248325 576918 248561
rect 577154 248325 577196 248561
rect 576876 241561 577196 248325
rect 576876 241325 576918 241561
rect 577154 241325 577196 241561
rect 576876 234561 577196 241325
rect 576876 234325 576918 234561
rect 577154 234325 577196 234561
rect 576876 227561 577196 234325
rect 576876 227325 576918 227561
rect 577154 227325 577196 227561
rect 576876 220561 577196 227325
rect 576876 220325 576918 220561
rect 577154 220325 577196 220561
rect 576876 213561 577196 220325
rect 576876 213325 576918 213561
rect 577154 213325 577196 213561
rect 576876 206561 577196 213325
rect 576876 206325 576918 206561
rect 577154 206325 577196 206561
rect 576876 199561 577196 206325
rect 576876 199325 576918 199561
rect 577154 199325 577196 199561
rect 576876 192561 577196 199325
rect 576876 192325 576918 192561
rect 577154 192325 577196 192561
rect 576876 185561 577196 192325
rect 576876 185325 576918 185561
rect 577154 185325 577196 185561
rect 576876 178561 577196 185325
rect 576876 178325 576918 178561
rect 577154 178325 577196 178561
rect 576876 171561 577196 178325
rect 576876 171325 576918 171561
rect 577154 171325 577196 171561
rect 576876 164561 577196 171325
rect 576876 164325 576918 164561
rect 577154 164325 577196 164561
rect 576876 157561 577196 164325
rect 576876 157325 576918 157561
rect 577154 157325 577196 157561
rect 576876 150561 577196 157325
rect 576876 150325 576918 150561
rect 577154 150325 577196 150561
rect 576876 143561 577196 150325
rect 576876 143325 576918 143561
rect 577154 143325 577196 143561
rect 576876 136561 577196 143325
rect 576876 136325 576918 136561
rect 577154 136325 577196 136561
rect 576876 129561 577196 136325
rect 576876 129325 576918 129561
rect 577154 129325 577196 129561
rect 576876 122561 577196 129325
rect 576876 122325 576918 122561
rect 577154 122325 577196 122561
rect 576876 115561 577196 122325
rect 576876 115325 576918 115561
rect 577154 115325 577196 115561
rect 576876 108561 577196 115325
rect 576876 108325 576918 108561
rect 577154 108325 577196 108561
rect 576876 101561 577196 108325
rect 576876 101325 576918 101561
rect 577154 101325 577196 101561
rect 576876 94561 577196 101325
rect 576876 94325 576918 94561
rect 577154 94325 577196 94561
rect 576876 87561 577196 94325
rect 576876 87325 576918 87561
rect 577154 87325 577196 87561
rect 576876 80561 577196 87325
rect 576876 80325 576918 80561
rect 577154 80325 577196 80561
rect 576876 73561 577196 80325
rect 576876 73325 576918 73561
rect 577154 73325 577196 73561
rect 576876 66561 577196 73325
rect 576876 66325 576918 66561
rect 577154 66325 577196 66561
rect 576876 59561 577196 66325
rect 576876 59325 576918 59561
rect 577154 59325 577196 59561
rect 576876 52561 577196 59325
rect 576876 52325 576918 52561
rect 577154 52325 577196 52561
rect 576876 45561 577196 52325
rect 576876 45325 576918 45561
rect 577154 45325 577196 45561
rect 576876 38561 577196 45325
rect 576876 38325 576918 38561
rect 577154 38325 577196 38561
rect 576876 31561 577196 38325
rect 576876 31325 576918 31561
rect 577154 31325 577196 31561
rect 576876 24561 577196 31325
rect 576876 24325 576918 24561
rect 577154 24325 577196 24561
rect 576876 17561 577196 24325
rect 576876 17325 576918 17561
rect 577154 17325 577196 17561
rect 576876 10561 577196 17325
rect 576876 10325 576918 10561
rect 577154 10325 577196 10561
rect 576876 3561 577196 10325
rect 576876 3325 576918 3561
rect 577154 3325 577196 3561
rect 576876 -1706 577196 3325
rect 576876 -1942 576918 -1706
rect 577154 -1942 577196 -1706
rect 576876 -2026 577196 -1942
rect 576876 -2262 576918 -2026
rect 577154 -2262 577196 -2026
rect 576876 -2294 577196 -2262
rect 582144 705238 582464 706230
rect 582144 705002 582186 705238
rect 582422 705002 582464 705238
rect 582144 704918 582464 705002
rect 582144 704682 582186 704918
rect 582422 704682 582464 704918
rect 582144 695494 582464 704682
rect 582144 695258 582186 695494
rect 582422 695258 582464 695494
rect 582144 688494 582464 695258
rect 582144 688258 582186 688494
rect 582422 688258 582464 688494
rect 582144 681494 582464 688258
rect 582144 681258 582186 681494
rect 582422 681258 582464 681494
rect 582144 674494 582464 681258
rect 582144 674258 582186 674494
rect 582422 674258 582464 674494
rect 582144 667494 582464 674258
rect 582144 667258 582186 667494
rect 582422 667258 582464 667494
rect 582144 660494 582464 667258
rect 582144 660258 582186 660494
rect 582422 660258 582464 660494
rect 582144 653494 582464 660258
rect 582144 653258 582186 653494
rect 582422 653258 582464 653494
rect 582144 646494 582464 653258
rect 582144 646258 582186 646494
rect 582422 646258 582464 646494
rect 582144 639494 582464 646258
rect 582144 639258 582186 639494
rect 582422 639258 582464 639494
rect 582144 632494 582464 639258
rect 582144 632258 582186 632494
rect 582422 632258 582464 632494
rect 582144 625494 582464 632258
rect 582144 625258 582186 625494
rect 582422 625258 582464 625494
rect 582144 618494 582464 625258
rect 582144 618258 582186 618494
rect 582422 618258 582464 618494
rect 582144 611494 582464 618258
rect 582144 611258 582186 611494
rect 582422 611258 582464 611494
rect 582144 604494 582464 611258
rect 582144 604258 582186 604494
rect 582422 604258 582464 604494
rect 582144 597494 582464 604258
rect 582144 597258 582186 597494
rect 582422 597258 582464 597494
rect 582144 590494 582464 597258
rect 582144 590258 582186 590494
rect 582422 590258 582464 590494
rect 582144 583494 582464 590258
rect 582144 583258 582186 583494
rect 582422 583258 582464 583494
rect 582144 576494 582464 583258
rect 582144 576258 582186 576494
rect 582422 576258 582464 576494
rect 582144 569494 582464 576258
rect 582144 569258 582186 569494
rect 582422 569258 582464 569494
rect 582144 562494 582464 569258
rect 582144 562258 582186 562494
rect 582422 562258 582464 562494
rect 582144 555494 582464 562258
rect 582144 555258 582186 555494
rect 582422 555258 582464 555494
rect 582144 548494 582464 555258
rect 582144 548258 582186 548494
rect 582422 548258 582464 548494
rect 582144 541494 582464 548258
rect 582144 541258 582186 541494
rect 582422 541258 582464 541494
rect 582144 534494 582464 541258
rect 582144 534258 582186 534494
rect 582422 534258 582464 534494
rect 582144 527494 582464 534258
rect 582144 527258 582186 527494
rect 582422 527258 582464 527494
rect 582144 520494 582464 527258
rect 582144 520258 582186 520494
rect 582422 520258 582464 520494
rect 582144 513494 582464 520258
rect 582144 513258 582186 513494
rect 582422 513258 582464 513494
rect 582144 506494 582464 513258
rect 582144 506258 582186 506494
rect 582422 506258 582464 506494
rect 582144 499494 582464 506258
rect 582144 499258 582186 499494
rect 582422 499258 582464 499494
rect 582144 492494 582464 499258
rect 582144 492258 582186 492494
rect 582422 492258 582464 492494
rect 582144 485494 582464 492258
rect 582144 485258 582186 485494
rect 582422 485258 582464 485494
rect 582144 478494 582464 485258
rect 582144 478258 582186 478494
rect 582422 478258 582464 478494
rect 582144 471494 582464 478258
rect 582144 471258 582186 471494
rect 582422 471258 582464 471494
rect 582144 464494 582464 471258
rect 582144 464258 582186 464494
rect 582422 464258 582464 464494
rect 582144 457494 582464 464258
rect 582144 457258 582186 457494
rect 582422 457258 582464 457494
rect 582144 450494 582464 457258
rect 582144 450258 582186 450494
rect 582422 450258 582464 450494
rect 582144 443494 582464 450258
rect 582144 443258 582186 443494
rect 582422 443258 582464 443494
rect 582144 436494 582464 443258
rect 582144 436258 582186 436494
rect 582422 436258 582464 436494
rect 582144 429494 582464 436258
rect 582144 429258 582186 429494
rect 582422 429258 582464 429494
rect 582144 422494 582464 429258
rect 582144 422258 582186 422494
rect 582422 422258 582464 422494
rect 582144 415494 582464 422258
rect 582144 415258 582186 415494
rect 582422 415258 582464 415494
rect 582144 408494 582464 415258
rect 582144 408258 582186 408494
rect 582422 408258 582464 408494
rect 582144 401494 582464 408258
rect 582144 401258 582186 401494
rect 582422 401258 582464 401494
rect 582144 394494 582464 401258
rect 582144 394258 582186 394494
rect 582422 394258 582464 394494
rect 582144 387494 582464 394258
rect 582144 387258 582186 387494
rect 582422 387258 582464 387494
rect 582144 380494 582464 387258
rect 582144 380258 582186 380494
rect 582422 380258 582464 380494
rect 582144 373494 582464 380258
rect 582144 373258 582186 373494
rect 582422 373258 582464 373494
rect 582144 366494 582464 373258
rect 582144 366258 582186 366494
rect 582422 366258 582464 366494
rect 582144 359494 582464 366258
rect 582144 359258 582186 359494
rect 582422 359258 582464 359494
rect 582144 352494 582464 359258
rect 582144 352258 582186 352494
rect 582422 352258 582464 352494
rect 582144 345494 582464 352258
rect 582144 345258 582186 345494
rect 582422 345258 582464 345494
rect 582144 338494 582464 345258
rect 582144 338258 582186 338494
rect 582422 338258 582464 338494
rect 582144 331494 582464 338258
rect 582144 331258 582186 331494
rect 582422 331258 582464 331494
rect 582144 324494 582464 331258
rect 582144 324258 582186 324494
rect 582422 324258 582464 324494
rect 582144 317494 582464 324258
rect 582144 317258 582186 317494
rect 582422 317258 582464 317494
rect 582144 310494 582464 317258
rect 582144 310258 582186 310494
rect 582422 310258 582464 310494
rect 582144 303494 582464 310258
rect 582144 303258 582186 303494
rect 582422 303258 582464 303494
rect 582144 296494 582464 303258
rect 582144 296258 582186 296494
rect 582422 296258 582464 296494
rect 582144 289494 582464 296258
rect 582144 289258 582186 289494
rect 582422 289258 582464 289494
rect 582144 282494 582464 289258
rect 582144 282258 582186 282494
rect 582422 282258 582464 282494
rect 582144 275494 582464 282258
rect 582144 275258 582186 275494
rect 582422 275258 582464 275494
rect 582144 268494 582464 275258
rect 582144 268258 582186 268494
rect 582422 268258 582464 268494
rect 582144 261494 582464 268258
rect 582144 261258 582186 261494
rect 582422 261258 582464 261494
rect 582144 254494 582464 261258
rect 582144 254258 582186 254494
rect 582422 254258 582464 254494
rect 582144 247494 582464 254258
rect 582144 247258 582186 247494
rect 582422 247258 582464 247494
rect 582144 240494 582464 247258
rect 582144 240258 582186 240494
rect 582422 240258 582464 240494
rect 582144 233494 582464 240258
rect 582144 233258 582186 233494
rect 582422 233258 582464 233494
rect 582144 226494 582464 233258
rect 582144 226258 582186 226494
rect 582422 226258 582464 226494
rect 582144 219494 582464 226258
rect 582144 219258 582186 219494
rect 582422 219258 582464 219494
rect 582144 212494 582464 219258
rect 582144 212258 582186 212494
rect 582422 212258 582464 212494
rect 582144 205494 582464 212258
rect 582144 205258 582186 205494
rect 582422 205258 582464 205494
rect 582144 198494 582464 205258
rect 582144 198258 582186 198494
rect 582422 198258 582464 198494
rect 582144 191494 582464 198258
rect 582144 191258 582186 191494
rect 582422 191258 582464 191494
rect 582144 184494 582464 191258
rect 582144 184258 582186 184494
rect 582422 184258 582464 184494
rect 582144 177494 582464 184258
rect 582144 177258 582186 177494
rect 582422 177258 582464 177494
rect 582144 170494 582464 177258
rect 582144 170258 582186 170494
rect 582422 170258 582464 170494
rect 582144 163494 582464 170258
rect 582144 163258 582186 163494
rect 582422 163258 582464 163494
rect 582144 156494 582464 163258
rect 582144 156258 582186 156494
rect 582422 156258 582464 156494
rect 582144 149494 582464 156258
rect 582144 149258 582186 149494
rect 582422 149258 582464 149494
rect 582144 142494 582464 149258
rect 582144 142258 582186 142494
rect 582422 142258 582464 142494
rect 582144 135494 582464 142258
rect 582144 135258 582186 135494
rect 582422 135258 582464 135494
rect 582144 128494 582464 135258
rect 582144 128258 582186 128494
rect 582422 128258 582464 128494
rect 582144 121494 582464 128258
rect 582144 121258 582186 121494
rect 582422 121258 582464 121494
rect 582144 114494 582464 121258
rect 582144 114258 582186 114494
rect 582422 114258 582464 114494
rect 582144 107494 582464 114258
rect 582144 107258 582186 107494
rect 582422 107258 582464 107494
rect 582144 100494 582464 107258
rect 582144 100258 582186 100494
rect 582422 100258 582464 100494
rect 582144 93494 582464 100258
rect 582144 93258 582186 93494
rect 582422 93258 582464 93494
rect 582144 86494 582464 93258
rect 582144 86258 582186 86494
rect 582422 86258 582464 86494
rect 582144 79494 582464 86258
rect 582144 79258 582186 79494
rect 582422 79258 582464 79494
rect 582144 72494 582464 79258
rect 582144 72258 582186 72494
rect 582422 72258 582464 72494
rect 582144 65494 582464 72258
rect 582144 65258 582186 65494
rect 582422 65258 582464 65494
rect 582144 58494 582464 65258
rect 582144 58258 582186 58494
rect 582422 58258 582464 58494
rect 582144 51494 582464 58258
rect 582144 51258 582186 51494
rect 582422 51258 582464 51494
rect 582144 44494 582464 51258
rect 582144 44258 582186 44494
rect 582422 44258 582464 44494
rect 582144 37494 582464 44258
rect 582144 37258 582186 37494
rect 582422 37258 582464 37494
rect 582144 30494 582464 37258
rect 582144 30258 582186 30494
rect 582422 30258 582464 30494
rect 582144 23494 582464 30258
rect 582144 23258 582186 23494
rect 582422 23258 582464 23494
rect 582144 16494 582464 23258
rect 582144 16258 582186 16494
rect 582422 16258 582464 16494
rect 582144 9494 582464 16258
rect 582144 9258 582186 9494
rect 582422 9258 582464 9494
rect 582144 2494 582464 9258
rect 582144 2258 582186 2494
rect 582422 2258 582464 2494
rect 582144 -746 582464 2258
rect 582144 -982 582186 -746
rect 582422 -982 582464 -746
rect 582144 -1066 582464 -982
rect 582144 -1302 582186 -1066
rect 582422 -1302 582464 -1066
rect 582144 -2294 582464 -1302
rect 585710 705238 587122 706062
rect 585710 705002 585818 705238
rect 586054 705002 586138 705238
rect 586374 705002 586458 705238
rect 586694 705002 586778 705238
rect 587014 705002 587122 705238
rect 585710 704918 587122 705002
rect 585710 704682 585818 704918
rect 586054 704682 586138 704918
rect 586374 704682 586458 704918
rect 586694 704682 586778 704918
rect 587014 704682 587122 704918
rect 585710 695494 587122 704682
rect 585710 695258 585818 695494
rect 586054 695258 586138 695494
rect 586374 695258 586458 695494
rect 586694 695258 586778 695494
rect 587014 695258 587122 695494
rect 585710 688494 587122 695258
rect 585710 688258 585818 688494
rect 586054 688258 586138 688494
rect 586374 688258 586458 688494
rect 586694 688258 586778 688494
rect 587014 688258 587122 688494
rect 585710 681494 587122 688258
rect 585710 681258 585818 681494
rect 586054 681258 586138 681494
rect 586374 681258 586458 681494
rect 586694 681258 586778 681494
rect 587014 681258 587122 681494
rect 585710 674494 587122 681258
rect 585710 674258 585818 674494
rect 586054 674258 586138 674494
rect 586374 674258 586458 674494
rect 586694 674258 586778 674494
rect 587014 674258 587122 674494
rect 585710 667494 587122 674258
rect 585710 667258 585818 667494
rect 586054 667258 586138 667494
rect 586374 667258 586458 667494
rect 586694 667258 586778 667494
rect 587014 667258 587122 667494
rect 585710 660494 587122 667258
rect 585710 660258 585818 660494
rect 586054 660258 586138 660494
rect 586374 660258 586458 660494
rect 586694 660258 586778 660494
rect 587014 660258 587122 660494
rect 585710 653494 587122 660258
rect 585710 653258 585818 653494
rect 586054 653258 586138 653494
rect 586374 653258 586458 653494
rect 586694 653258 586778 653494
rect 587014 653258 587122 653494
rect 585710 646494 587122 653258
rect 585710 646258 585818 646494
rect 586054 646258 586138 646494
rect 586374 646258 586458 646494
rect 586694 646258 586778 646494
rect 587014 646258 587122 646494
rect 585710 639494 587122 646258
rect 585710 639258 585818 639494
rect 586054 639258 586138 639494
rect 586374 639258 586458 639494
rect 586694 639258 586778 639494
rect 587014 639258 587122 639494
rect 585710 632494 587122 639258
rect 585710 632258 585818 632494
rect 586054 632258 586138 632494
rect 586374 632258 586458 632494
rect 586694 632258 586778 632494
rect 587014 632258 587122 632494
rect 585710 625494 587122 632258
rect 585710 625258 585818 625494
rect 586054 625258 586138 625494
rect 586374 625258 586458 625494
rect 586694 625258 586778 625494
rect 587014 625258 587122 625494
rect 585710 618494 587122 625258
rect 585710 618258 585818 618494
rect 586054 618258 586138 618494
rect 586374 618258 586458 618494
rect 586694 618258 586778 618494
rect 587014 618258 587122 618494
rect 585710 611494 587122 618258
rect 585710 611258 585818 611494
rect 586054 611258 586138 611494
rect 586374 611258 586458 611494
rect 586694 611258 586778 611494
rect 587014 611258 587122 611494
rect 585710 604494 587122 611258
rect 585710 604258 585818 604494
rect 586054 604258 586138 604494
rect 586374 604258 586458 604494
rect 586694 604258 586778 604494
rect 587014 604258 587122 604494
rect 585710 597494 587122 604258
rect 585710 597258 585818 597494
rect 586054 597258 586138 597494
rect 586374 597258 586458 597494
rect 586694 597258 586778 597494
rect 587014 597258 587122 597494
rect 585710 590494 587122 597258
rect 585710 590258 585818 590494
rect 586054 590258 586138 590494
rect 586374 590258 586458 590494
rect 586694 590258 586778 590494
rect 587014 590258 587122 590494
rect 585710 583494 587122 590258
rect 585710 583258 585818 583494
rect 586054 583258 586138 583494
rect 586374 583258 586458 583494
rect 586694 583258 586778 583494
rect 587014 583258 587122 583494
rect 585710 576494 587122 583258
rect 585710 576258 585818 576494
rect 586054 576258 586138 576494
rect 586374 576258 586458 576494
rect 586694 576258 586778 576494
rect 587014 576258 587122 576494
rect 585710 569494 587122 576258
rect 585710 569258 585818 569494
rect 586054 569258 586138 569494
rect 586374 569258 586458 569494
rect 586694 569258 586778 569494
rect 587014 569258 587122 569494
rect 585710 562494 587122 569258
rect 585710 562258 585818 562494
rect 586054 562258 586138 562494
rect 586374 562258 586458 562494
rect 586694 562258 586778 562494
rect 587014 562258 587122 562494
rect 585710 555494 587122 562258
rect 585710 555258 585818 555494
rect 586054 555258 586138 555494
rect 586374 555258 586458 555494
rect 586694 555258 586778 555494
rect 587014 555258 587122 555494
rect 585710 548494 587122 555258
rect 585710 548258 585818 548494
rect 586054 548258 586138 548494
rect 586374 548258 586458 548494
rect 586694 548258 586778 548494
rect 587014 548258 587122 548494
rect 585710 541494 587122 548258
rect 585710 541258 585818 541494
rect 586054 541258 586138 541494
rect 586374 541258 586458 541494
rect 586694 541258 586778 541494
rect 587014 541258 587122 541494
rect 585710 534494 587122 541258
rect 585710 534258 585818 534494
rect 586054 534258 586138 534494
rect 586374 534258 586458 534494
rect 586694 534258 586778 534494
rect 587014 534258 587122 534494
rect 585710 527494 587122 534258
rect 585710 527258 585818 527494
rect 586054 527258 586138 527494
rect 586374 527258 586458 527494
rect 586694 527258 586778 527494
rect 587014 527258 587122 527494
rect 585710 520494 587122 527258
rect 585710 520258 585818 520494
rect 586054 520258 586138 520494
rect 586374 520258 586458 520494
rect 586694 520258 586778 520494
rect 587014 520258 587122 520494
rect 585710 513494 587122 520258
rect 585710 513258 585818 513494
rect 586054 513258 586138 513494
rect 586374 513258 586458 513494
rect 586694 513258 586778 513494
rect 587014 513258 587122 513494
rect 585710 506494 587122 513258
rect 585710 506258 585818 506494
rect 586054 506258 586138 506494
rect 586374 506258 586458 506494
rect 586694 506258 586778 506494
rect 587014 506258 587122 506494
rect 585710 499494 587122 506258
rect 585710 499258 585818 499494
rect 586054 499258 586138 499494
rect 586374 499258 586458 499494
rect 586694 499258 586778 499494
rect 587014 499258 587122 499494
rect 585710 492494 587122 499258
rect 585710 492258 585818 492494
rect 586054 492258 586138 492494
rect 586374 492258 586458 492494
rect 586694 492258 586778 492494
rect 587014 492258 587122 492494
rect 585710 485494 587122 492258
rect 585710 485258 585818 485494
rect 586054 485258 586138 485494
rect 586374 485258 586458 485494
rect 586694 485258 586778 485494
rect 587014 485258 587122 485494
rect 585710 478494 587122 485258
rect 585710 478258 585818 478494
rect 586054 478258 586138 478494
rect 586374 478258 586458 478494
rect 586694 478258 586778 478494
rect 587014 478258 587122 478494
rect 585710 471494 587122 478258
rect 585710 471258 585818 471494
rect 586054 471258 586138 471494
rect 586374 471258 586458 471494
rect 586694 471258 586778 471494
rect 587014 471258 587122 471494
rect 585710 464494 587122 471258
rect 585710 464258 585818 464494
rect 586054 464258 586138 464494
rect 586374 464258 586458 464494
rect 586694 464258 586778 464494
rect 587014 464258 587122 464494
rect 585710 457494 587122 464258
rect 585710 457258 585818 457494
rect 586054 457258 586138 457494
rect 586374 457258 586458 457494
rect 586694 457258 586778 457494
rect 587014 457258 587122 457494
rect 585710 450494 587122 457258
rect 585710 450258 585818 450494
rect 586054 450258 586138 450494
rect 586374 450258 586458 450494
rect 586694 450258 586778 450494
rect 587014 450258 587122 450494
rect 585710 443494 587122 450258
rect 585710 443258 585818 443494
rect 586054 443258 586138 443494
rect 586374 443258 586458 443494
rect 586694 443258 586778 443494
rect 587014 443258 587122 443494
rect 585710 436494 587122 443258
rect 585710 436258 585818 436494
rect 586054 436258 586138 436494
rect 586374 436258 586458 436494
rect 586694 436258 586778 436494
rect 587014 436258 587122 436494
rect 585710 429494 587122 436258
rect 585710 429258 585818 429494
rect 586054 429258 586138 429494
rect 586374 429258 586458 429494
rect 586694 429258 586778 429494
rect 587014 429258 587122 429494
rect 585710 422494 587122 429258
rect 585710 422258 585818 422494
rect 586054 422258 586138 422494
rect 586374 422258 586458 422494
rect 586694 422258 586778 422494
rect 587014 422258 587122 422494
rect 585710 415494 587122 422258
rect 585710 415258 585818 415494
rect 586054 415258 586138 415494
rect 586374 415258 586458 415494
rect 586694 415258 586778 415494
rect 587014 415258 587122 415494
rect 585710 408494 587122 415258
rect 585710 408258 585818 408494
rect 586054 408258 586138 408494
rect 586374 408258 586458 408494
rect 586694 408258 586778 408494
rect 587014 408258 587122 408494
rect 585710 401494 587122 408258
rect 585710 401258 585818 401494
rect 586054 401258 586138 401494
rect 586374 401258 586458 401494
rect 586694 401258 586778 401494
rect 587014 401258 587122 401494
rect 585710 394494 587122 401258
rect 585710 394258 585818 394494
rect 586054 394258 586138 394494
rect 586374 394258 586458 394494
rect 586694 394258 586778 394494
rect 587014 394258 587122 394494
rect 585710 387494 587122 394258
rect 585710 387258 585818 387494
rect 586054 387258 586138 387494
rect 586374 387258 586458 387494
rect 586694 387258 586778 387494
rect 587014 387258 587122 387494
rect 585710 380494 587122 387258
rect 585710 380258 585818 380494
rect 586054 380258 586138 380494
rect 586374 380258 586458 380494
rect 586694 380258 586778 380494
rect 587014 380258 587122 380494
rect 585710 373494 587122 380258
rect 585710 373258 585818 373494
rect 586054 373258 586138 373494
rect 586374 373258 586458 373494
rect 586694 373258 586778 373494
rect 587014 373258 587122 373494
rect 585710 366494 587122 373258
rect 585710 366258 585818 366494
rect 586054 366258 586138 366494
rect 586374 366258 586458 366494
rect 586694 366258 586778 366494
rect 587014 366258 587122 366494
rect 585710 359494 587122 366258
rect 585710 359258 585818 359494
rect 586054 359258 586138 359494
rect 586374 359258 586458 359494
rect 586694 359258 586778 359494
rect 587014 359258 587122 359494
rect 585710 352494 587122 359258
rect 585710 352258 585818 352494
rect 586054 352258 586138 352494
rect 586374 352258 586458 352494
rect 586694 352258 586778 352494
rect 587014 352258 587122 352494
rect 585710 345494 587122 352258
rect 585710 345258 585818 345494
rect 586054 345258 586138 345494
rect 586374 345258 586458 345494
rect 586694 345258 586778 345494
rect 587014 345258 587122 345494
rect 585710 338494 587122 345258
rect 585710 338258 585818 338494
rect 586054 338258 586138 338494
rect 586374 338258 586458 338494
rect 586694 338258 586778 338494
rect 587014 338258 587122 338494
rect 585710 331494 587122 338258
rect 585710 331258 585818 331494
rect 586054 331258 586138 331494
rect 586374 331258 586458 331494
rect 586694 331258 586778 331494
rect 587014 331258 587122 331494
rect 585710 324494 587122 331258
rect 585710 324258 585818 324494
rect 586054 324258 586138 324494
rect 586374 324258 586458 324494
rect 586694 324258 586778 324494
rect 587014 324258 587122 324494
rect 585710 317494 587122 324258
rect 585710 317258 585818 317494
rect 586054 317258 586138 317494
rect 586374 317258 586458 317494
rect 586694 317258 586778 317494
rect 587014 317258 587122 317494
rect 585710 310494 587122 317258
rect 585710 310258 585818 310494
rect 586054 310258 586138 310494
rect 586374 310258 586458 310494
rect 586694 310258 586778 310494
rect 587014 310258 587122 310494
rect 585710 303494 587122 310258
rect 585710 303258 585818 303494
rect 586054 303258 586138 303494
rect 586374 303258 586458 303494
rect 586694 303258 586778 303494
rect 587014 303258 587122 303494
rect 585710 296494 587122 303258
rect 585710 296258 585818 296494
rect 586054 296258 586138 296494
rect 586374 296258 586458 296494
rect 586694 296258 586778 296494
rect 587014 296258 587122 296494
rect 585710 289494 587122 296258
rect 585710 289258 585818 289494
rect 586054 289258 586138 289494
rect 586374 289258 586458 289494
rect 586694 289258 586778 289494
rect 587014 289258 587122 289494
rect 585710 282494 587122 289258
rect 585710 282258 585818 282494
rect 586054 282258 586138 282494
rect 586374 282258 586458 282494
rect 586694 282258 586778 282494
rect 587014 282258 587122 282494
rect 585710 275494 587122 282258
rect 585710 275258 585818 275494
rect 586054 275258 586138 275494
rect 586374 275258 586458 275494
rect 586694 275258 586778 275494
rect 587014 275258 587122 275494
rect 585710 268494 587122 275258
rect 585710 268258 585818 268494
rect 586054 268258 586138 268494
rect 586374 268258 586458 268494
rect 586694 268258 586778 268494
rect 587014 268258 587122 268494
rect 585710 261494 587122 268258
rect 585710 261258 585818 261494
rect 586054 261258 586138 261494
rect 586374 261258 586458 261494
rect 586694 261258 586778 261494
rect 587014 261258 587122 261494
rect 585710 254494 587122 261258
rect 585710 254258 585818 254494
rect 586054 254258 586138 254494
rect 586374 254258 586458 254494
rect 586694 254258 586778 254494
rect 587014 254258 587122 254494
rect 585710 247494 587122 254258
rect 585710 247258 585818 247494
rect 586054 247258 586138 247494
rect 586374 247258 586458 247494
rect 586694 247258 586778 247494
rect 587014 247258 587122 247494
rect 585710 240494 587122 247258
rect 585710 240258 585818 240494
rect 586054 240258 586138 240494
rect 586374 240258 586458 240494
rect 586694 240258 586778 240494
rect 587014 240258 587122 240494
rect 585710 233494 587122 240258
rect 585710 233258 585818 233494
rect 586054 233258 586138 233494
rect 586374 233258 586458 233494
rect 586694 233258 586778 233494
rect 587014 233258 587122 233494
rect 585710 226494 587122 233258
rect 585710 226258 585818 226494
rect 586054 226258 586138 226494
rect 586374 226258 586458 226494
rect 586694 226258 586778 226494
rect 587014 226258 587122 226494
rect 585710 219494 587122 226258
rect 585710 219258 585818 219494
rect 586054 219258 586138 219494
rect 586374 219258 586458 219494
rect 586694 219258 586778 219494
rect 587014 219258 587122 219494
rect 585710 212494 587122 219258
rect 585710 212258 585818 212494
rect 586054 212258 586138 212494
rect 586374 212258 586458 212494
rect 586694 212258 586778 212494
rect 587014 212258 587122 212494
rect 585710 205494 587122 212258
rect 585710 205258 585818 205494
rect 586054 205258 586138 205494
rect 586374 205258 586458 205494
rect 586694 205258 586778 205494
rect 587014 205258 587122 205494
rect 585710 198494 587122 205258
rect 585710 198258 585818 198494
rect 586054 198258 586138 198494
rect 586374 198258 586458 198494
rect 586694 198258 586778 198494
rect 587014 198258 587122 198494
rect 585710 191494 587122 198258
rect 585710 191258 585818 191494
rect 586054 191258 586138 191494
rect 586374 191258 586458 191494
rect 586694 191258 586778 191494
rect 587014 191258 587122 191494
rect 585710 184494 587122 191258
rect 585710 184258 585818 184494
rect 586054 184258 586138 184494
rect 586374 184258 586458 184494
rect 586694 184258 586778 184494
rect 587014 184258 587122 184494
rect 585710 177494 587122 184258
rect 585710 177258 585818 177494
rect 586054 177258 586138 177494
rect 586374 177258 586458 177494
rect 586694 177258 586778 177494
rect 587014 177258 587122 177494
rect 585710 170494 587122 177258
rect 585710 170258 585818 170494
rect 586054 170258 586138 170494
rect 586374 170258 586458 170494
rect 586694 170258 586778 170494
rect 587014 170258 587122 170494
rect 585710 163494 587122 170258
rect 585710 163258 585818 163494
rect 586054 163258 586138 163494
rect 586374 163258 586458 163494
rect 586694 163258 586778 163494
rect 587014 163258 587122 163494
rect 585710 156494 587122 163258
rect 585710 156258 585818 156494
rect 586054 156258 586138 156494
rect 586374 156258 586458 156494
rect 586694 156258 586778 156494
rect 587014 156258 587122 156494
rect 585710 149494 587122 156258
rect 585710 149258 585818 149494
rect 586054 149258 586138 149494
rect 586374 149258 586458 149494
rect 586694 149258 586778 149494
rect 587014 149258 587122 149494
rect 585710 142494 587122 149258
rect 585710 142258 585818 142494
rect 586054 142258 586138 142494
rect 586374 142258 586458 142494
rect 586694 142258 586778 142494
rect 587014 142258 587122 142494
rect 585710 135494 587122 142258
rect 585710 135258 585818 135494
rect 586054 135258 586138 135494
rect 586374 135258 586458 135494
rect 586694 135258 586778 135494
rect 587014 135258 587122 135494
rect 585710 128494 587122 135258
rect 585710 128258 585818 128494
rect 586054 128258 586138 128494
rect 586374 128258 586458 128494
rect 586694 128258 586778 128494
rect 587014 128258 587122 128494
rect 585710 121494 587122 128258
rect 585710 121258 585818 121494
rect 586054 121258 586138 121494
rect 586374 121258 586458 121494
rect 586694 121258 586778 121494
rect 587014 121258 587122 121494
rect 585710 114494 587122 121258
rect 585710 114258 585818 114494
rect 586054 114258 586138 114494
rect 586374 114258 586458 114494
rect 586694 114258 586778 114494
rect 587014 114258 587122 114494
rect 585710 107494 587122 114258
rect 585710 107258 585818 107494
rect 586054 107258 586138 107494
rect 586374 107258 586458 107494
rect 586694 107258 586778 107494
rect 587014 107258 587122 107494
rect 585710 100494 587122 107258
rect 585710 100258 585818 100494
rect 586054 100258 586138 100494
rect 586374 100258 586458 100494
rect 586694 100258 586778 100494
rect 587014 100258 587122 100494
rect 585710 93494 587122 100258
rect 585710 93258 585818 93494
rect 586054 93258 586138 93494
rect 586374 93258 586458 93494
rect 586694 93258 586778 93494
rect 587014 93258 587122 93494
rect 585710 86494 587122 93258
rect 585710 86258 585818 86494
rect 586054 86258 586138 86494
rect 586374 86258 586458 86494
rect 586694 86258 586778 86494
rect 587014 86258 587122 86494
rect 585710 79494 587122 86258
rect 585710 79258 585818 79494
rect 586054 79258 586138 79494
rect 586374 79258 586458 79494
rect 586694 79258 586778 79494
rect 587014 79258 587122 79494
rect 585710 72494 587122 79258
rect 585710 72258 585818 72494
rect 586054 72258 586138 72494
rect 586374 72258 586458 72494
rect 586694 72258 586778 72494
rect 587014 72258 587122 72494
rect 585710 65494 587122 72258
rect 585710 65258 585818 65494
rect 586054 65258 586138 65494
rect 586374 65258 586458 65494
rect 586694 65258 586778 65494
rect 587014 65258 587122 65494
rect 585710 58494 587122 65258
rect 585710 58258 585818 58494
rect 586054 58258 586138 58494
rect 586374 58258 586458 58494
rect 586694 58258 586778 58494
rect 587014 58258 587122 58494
rect 585710 51494 587122 58258
rect 585710 51258 585818 51494
rect 586054 51258 586138 51494
rect 586374 51258 586458 51494
rect 586694 51258 586778 51494
rect 587014 51258 587122 51494
rect 585710 44494 587122 51258
rect 585710 44258 585818 44494
rect 586054 44258 586138 44494
rect 586374 44258 586458 44494
rect 586694 44258 586778 44494
rect 587014 44258 587122 44494
rect 585710 37494 587122 44258
rect 585710 37258 585818 37494
rect 586054 37258 586138 37494
rect 586374 37258 586458 37494
rect 586694 37258 586778 37494
rect 587014 37258 587122 37494
rect 585710 30494 587122 37258
rect 585710 30258 585818 30494
rect 586054 30258 586138 30494
rect 586374 30258 586458 30494
rect 586694 30258 586778 30494
rect 587014 30258 587122 30494
rect 585710 23494 587122 30258
rect 585710 23258 585818 23494
rect 586054 23258 586138 23494
rect 586374 23258 586458 23494
rect 586694 23258 586778 23494
rect 587014 23258 587122 23494
rect 585710 16494 587122 23258
rect 585710 16258 585818 16494
rect 586054 16258 586138 16494
rect 586374 16258 586458 16494
rect 586694 16258 586778 16494
rect 587014 16258 587122 16494
rect 585710 9494 587122 16258
rect 585710 9258 585818 9494
rect 586054 9258 586138 9494
rect 586374 9258 586458 9494
rect 586694 9258 586778 9494
rect 587014 9258 587122 9494
rect 585710 2494 587122 9258
rect 585710 2258 585818 2494
rect 586054 2258 586138 2494
rect 586374 2258 586458 2494
rect 586694 2258 586778 2494
rect 587014 2258 587122 2494
rect 585710 -746 587122 2258
rect 585710 -982 585818 -746
rect 586054 -982 586138 -746
rect 586374 -982 586458 -746
rect 586694 -982 586778 -746
rect 587014 -982 587122 -746
rect 585710 -1066 587122 -982
rect 585710 -1302 585818 -1066
rect 586054 -1302 586138 -1066
rect 586374 -1302 586458 -1066
rect 586694 -1302 586778 -1066
rect 587014 -1302 587122 -1066
rect 585710 -2126 587122 -1302
rect 587462 696561 588874 707814
rect 587462 696325 587570 696561
rect 587806 696325 587890 696561
rect 588126 696325 588210 696561
rect 588446 696325 588530 696561
rect 588766 696325 588874 696561
rect 587462 689561 588874 696325
rect 587462 689325 587570 689561
rect 587806 689325 587890 689561
rect 588126 689325 588210 689561
rect 588446 689325 588530 689561
rect 588766 689325 588874 689561
rect 587462 682561 588874 689325
rect 587462 682325 587570 682561
rect 587806 682325 587890 682561
rect 588126 682325 588210 682561
rect 588446 682325 588530 682561
rect 588766 682325 588874 682561
rect 587462 675561 588874 682325
rect 587462 675325 587570 675561
rect 587806 675325 587890 675561
rect 588126 675325 588210 675561
rect 588446 675325 588530 675561
rect 588766 675325 588874 675561
rect 587462 668561 588874 675325
rect 587462 668325 587570 668561
rect 587806 668325 587890 668561
rect 588126 668325 588210 668561
rect 588446 668325 588530 668561
rect 588766 668325 588874 668561
rect 587462 661561 588874 668325
rect 587462 661325 587570 661561
rect 587806 661325 587890 661561
rect 588126 661325 588210 661561
rect 588446 661325 588530 661561
rect 588766 661325 588874 661561
rect 587462 654561 588874 661325
rect 587462 654325 587570 654561
rect 587806 654325 587890 654561
rect 588126 654325 588210 654561
rect 588446 654325 588530 654561
rect 588766 654325 588874 654561
rect 587462 647561 588874 654325
rect 587462 647325 587570 647561
rect 587806 647325 587890 647561
rect 588126 647325 588210 647561
rect 588446 647325 588530 647561
rect 588766 647325 588874 647561
rect 587462 640561 588874 647325
rect 587462 640325 587570 640561
rect 587806 640325 587890 640561
rect 588126 640325 588210 640561
rect 588446 640325 588530 640561
rect 588766 640325 588874 640561
rect 587462 633561 588874 640325
rect 587462 633325 587570 633561
rect 587806 633325 587890 633561
rect 588126 633325 588210 633561
rect 588446 633325 588530 633561
rect 588766 633325 588874 633561
rect 587462 626561 588874 633325
rect 587462 626325 587570 626561
rect 587806 626325 587890 626561
rect 588126 626325 588210 626561
rect 588446 626325 588530 626561
rect 588766 626325 588874 626561
rect 587462 619561 588874 626325
rect 587462 619325 587570 619561
rect 587806 619325 587890 619561
rect 588126 619325 588210 619561
rect 588446 619325 588530 619561
rect 588766 619325 588874 619561
rect 587462 612561 588874 619325
rect 587462 612325 587570 612561
rect 587806 612325 587890 612561
rect 588126 612325 588210 612561
rect 588446 612325 588530 612561
rect 588766 612325 588874 612561
rect 587462 605561 588874 612325
rect 587462 605325 587570 605561
rect 587806 605325 587890 605561
rect 588126 605325 588210 605561
rect 588446 605325 588530 605561
rect 588766 605325 588874 605561
rect 587462 598561 588874 605325
rect 587462 598325 587570 598561
rect 587806 598325 587890 598561
rect 588126 598325 588210 598561
rect 588446 598325 588530 598561
rect 588766 598325 588874 598561
rect 587462 591561 588874 598325
rect 587462 591325 587570 591561
rect 587806 591325 587890 591561
rect 588126 591325 588210 591561
rect 588446 591325 588530 591561
rect 588766 591325 588874 591561
rect 587462 584561 588874 591325
rect 587462 584325 587570 584561
rect 587806 584325 587890 584561
rect 588126 584325 588210 584561
rect 588446 584325 588530 584561
rect 588766 584325 588874 584561
rect 587462 577561 588874 584325
rect 587462 577325 587570 577561
rect 587806 577325 587890 577561
rect 588126 577325 588210 577561
rect 588446 577325 588530 577561
rect 588766 577325 588874 577561
rect 587462 570561 588874 577325
rect 587462 570325 587570 570561
rect 587806 570325 587890 570561
rect 588126 570325 588210 570561
rect 588446 570325 588530 570561
rect 588766 570325 588874 570561
rect 587462 563561 588874 570325
rect 587462 563325 587570 563561
rect 587806 563325 587890 563561
rect 588126 563325 588210 563561
rect 588446 563325 588530 563561
rect 588766 563325 588874 563561
rect 587462 556561 588874 563325
rect 587462 556325 587570 556561
rect 587806 556325 587890 556561
rect 588126 556325 588210 556561
rect 588446 556325 588530 556561
rect 588766 556325 588874 556561
rect 587462 549561 588874 556325
rect 587462 549325 587570 549561
rect 587806 549325 587890 549561
rect 588126 549325 588210 549561
rect 588446 549325 588530 549561
rect 588766 549325 588874 549561
rect 587462 542561 588874 549325
rect 587462 542325 587570 542561
rect 587806 542325 587890 542561
rect 588126 542325 588210 542561
rect 588446 542325 588530 542561
rect 588766 542325 588874 542561
rect 587462 535561 588874 542325
rect 587462 535325 587570 535561
rect 587806 535325 587890 535561
rect 588126 535325 588210 535561
rect 588446 535325 588530 535561
rect 588766 535325 588874 535561
rect 587462 528561 588874 535325
rect 587462 528325 587570 528561
rect 587806 528325 587890 528561
rect 588126 528325 588210 528561
rect 588446 528325 588530 528561
rect 588766 528325 588874 528561
rect 587462 521561 588874 528325
rect 587462 521325 587570 521561
rect 587806 521325 587890 521561
rect 588126 521325 588210 521561
rect 588446 521325 588530 521561
rect 588766 521325 588874 521561
rect 587462 514561 588874 521325
rect 587462 514325 587570 514561
rect 587806 514325 587890 514561
rect 588126 514325 588210 514561
rect 588446 514325 588530 514561
rect 588766 514325 588874 514561
rect 587462 507561 588874 514325
rect 587462 507325 587570 507561
rect 587806 507325 587890 507561
rect 588126 507325 588210 507561
rect 588446 507325 588530 507561
rect 588766 507325 588874 507561
rect 587462 500561 588874 507325
rect 587462 500325 587570 500561
rect 587806 500325 587890 500561
rect 588126 500325 588210 500561
rect 588446 500325 588530 500561
rect 588766 500325 588874 500561
rect 587462 493561 588874 500325
rect 587462 493325 587570 493561
rect 587806 493325 587890 493561
rect 588126 493325 588210 493561
rect 588446 493325 588530 493561
rect 588766 493325 588874 493561
rect 587462 486561 588874 493325
rect 587462 486325 587570 486561
rect 587806 486325 587890 486561
rect 588126 486325 588210 486561
rect 588446 486325 588530 486561
rect 588766 486325 588874 486561
rect 587462 479561 588874 486325
rect 587462 479325 587570 479561
rect 587806 479325 587890 479561
rect 588126 479325 588210 479561
rect 588446 479325 588530 479561
rect 588766 479325 588874 479561
rect 587462 472561 588874 479325
rect 587462 472325 587570 472561
rect 587806 472325 587890 472561
rect 588126 472325 588210 472561
rect 588446 472325 588530 472561
rect 588766 472325 588874 472561
rect 587462 465561 588874 472325
rect 587462 465325 587570 465561
rect 587806 465325 587890 465561
rect 588126 465325 588210 465561
rect 588446 465325 588530 465561
rect 588766 465325 588874 465561
rect 587462 458561 588874 465325
rect 587462 458325 587570 458561
rect 587806 458325 587890 458561
rect 588126 458325 588210 458561
rect 588446 458325 588530 458561
rect 588766 458325 588874 458561
rect 587462 451561 588874 458325
rect 587462 451325 587570 451561
rect 587806 451325 587890 451561
rect 588126 451325 588210 451561
rect 588446 451325 588530 451561
rect 588766 451325 588874 451561
rect 587462 444561 588874 451325
rect 587462 444325 587570 444561
rect 587806 444325 587890 444561
rect 588126 444325 588210 444561
rect 588446 444325 588530 444561
rect 588766 444325 588874 444561
rect 587462 437561 588874 444325
rect 587462 437325 587570 437561
rect 587806 437325 587890 437561
rect 588126 437325 588210 437561
rect 588446 437325 588530 437561
rect 588766 437325 588874 437561
rect 587462 430561 588874 437325
rect 587462 430325 587570 430561
rect 587806 430325 587890 430561
rect 588126 430325 588210 430561
rect 588446 430325 588530 430561
rect 588766 430325 588874 430561
rect 587462 423561 588874 430325
rect 587462 423325 587570 423561
rect 587806 423325 587890 423561
rect 588126 423325 588210 423561
rect 588446 423325 588530 423561
rect 588766 423325 588874 423561
rect 587462 416561 588874 423325
rect 587462 416325 587570 416561
rect 587806 416325 587890 416561
rect 588126 416325 588210 416561
rect 588446 416325 588530 416561
rect 588766 416325 588874 416561
rect 587462 409561 588874 416325
rect 587462 409325 587570 409561
rect 587806 409325 587890 409561
rect 588126 409325 588210 409561
rect 588446 409325 588530 409561
rect 588766 409325 588874 409561
rect 587462 402561 588874 409325
rect 587462 402325 587570 402561
rect 587806 402325 587890 402561
rect 588126 402325 588210 402561
rect 588446 402325 588530 402561
rect 588766 402325 588874 402561
rect 587462 395561 588874 402325
rect 587462 395325 587570 395561
rect 587806 395325 587890 395561
rect 588126 395325 588210 395561
rect 588446 395325 588530 395561
rect 588766 395325 588874 395561
rect 587462 388561 588874 395325
rect 587462 388325 587570 388561
rect 587806 388325 587890 388561
rect 588126 388325 588210 388561
rect 588446 388325 588530 388561
rect 588766 388325 588874 388561
rect 587462 381561 588874 388325
rect 587462 381325 587570 381561
rect 587806 381325 587890 381561
rect 588126 381325 588210 381561
rect 588446 381325 588530 381561
rect 588766 381325 588874 381561
rect 587462 374561 588874 381325
rect 587462 374325 587570 374561
rect 587806 374325 587890 374561
rect 588126 374325 588210 374561
rect 588446 374325 588530 374561
rect 588766 374325 588874 374561
rect 587462 367561 588874 374325
rect 587462 367325 587570 367561
rect 587806 367325 587890 367561
rect 588126 367325 588210 367561
rect 588446 367325 588530 367561
rect 588766 367325 588874 367561
rect 587462 360561 588874 367325
rect 587462 360325 587570 360561
rect 587806 360325 587890 360561
rect 588126 360325 588210 360561
rect 588446 360325 588530 360561
rect 588766 360325 588874 360561
rect 587462 353561 588874 360325
rect 587462 353325 587570 353561
rect 587806 353325 587890 353561
rect 588126 353325 588210 353561
rect 588446 353325 588530 353561
rect 588766 353325 588874 353561
rect 587462 346561 588874 353325
rect 587462 346325 587570 346561
rect 587806 346325 587890 346561
rect 588126 346325 588210 346561
rect 588446 346325 588530 346561
rect 588766 346325 588874 346561
rect 587462 339561 588874 346325
rect 587462 339325 587570 339561
rect 587806 339325 587890 339561
rect 588126 339325 588210 339561
rect 588446 339325 588530 339561
rect 588766 339325 588874 339561
rect 587462 332561 588874 339325
rect 587462 332325 587570 332561
rect 587806 332325 587890 332561
rect 588126 332325 588210 332561
rect 588446 332325 588530 332561
rect 588766 332325 588874 332561
rect 587462 325561 588874 332325
rect 587462 325325 587570 325561
rect 587806 325325 587890 325561
rect 588126 325325 588210 325561
rect 588446 325325 588530 325561
rect 588766 325325 588874 325561
rect 587462 318561 588874 325325
rect 587462 318325 587570 318561
rect 587806 318325 587890 318561
rect 588126 318325 588210 318561
rect 588446 318325 588530 318561
rect 588766 318325 588874 318561
rect 587462 311561 588874 318325
rect 587462 311325 587570 311561
rect 587806 311325 587890 311561
rect 588126 311325 588210 311561
rect 588446 311325 588530 311561
rect 588766 311325 588874 311561
rect 587462 304561 588874 311325
rect 587462 304325 587570 304561
rect 587806 304325 587890 304561
rect 588126 304325 588210 304561
rect 588446 304325 588530 304561
rect 588766 304325 588874 304561
rect 587462 297561 588874 304325
rect 587462 297325 587570 297561
rect 587806 297325 587890 297561
rect 588126 297325 588210 297561
rect 588446 297325 588530 297561
rect 588766 297325 588874 297561
rect 587462 290561 588874 297325
rect 587462 290325 587570 290561
rect 587806 290325 587890 290561
rect 588126 290325 588210 290561
rect 588446 290325 588530 290561
rect 588766 290325 588874 290561
rect 587462 283561 588874 290325
rect 587462 283325 587570 283561
rect 587806 283325 587890 283561
rect 588126 283325 588210 283561
rect 588446 283325 588530 283561
rect 588766 283325 588874 283561
rect 587462 276561 588874 283325
rect 587462 276325 587570 276561
rect 587806 276325 587890 276561
rect 588126 276325 588210 276561
rect 588446 276325 588530 276561
rect 588766 276325 588874 276561
rect 587462 269561 588874 276325
rect 587462 269325 587570 269561
rect 587806 269325 587890 269561
rect 588126 269325 588210 269561
rect 588446 269325 588530 269561
rect 588766 269325 588874 269561
rect 587462 262561 588874 269325
rect 587462 262325 587570 262561
rect 587806 262325 587890 262561
rect 588126 262325 588210 262561
rect 588446 262325 588530 262561
rect 588766 262325 588874 262561
rect 587462 255561 588874 262325
rect 587462 255325 587570 255561
rect 587806 255325 587890 255561
rect 588126 255325 588210 255561
rect 588446 255325 588530 255561
rect 588766 255325 588874 255561
rect 587462 248561 588874 255325
rect 587462 248325 587570 248561
rect 587806 248325 587890 248561
rect 588126 248325 588210 248561
rect 588446 248325 588530 248561
rect 588766 248325 588874 248561
rect 587462 241561 588874 248325
rect 587462 241325 587570 241561
rect 587806 241325 587890 241561
rect 588126 241325 588210 241561
rect 588446 241325 588530 241561
rect 588766 241325 588874 241561
rect 587462 234561 588874 241325
rect 587462 234325 587570 234561
rect 587806 234325 587890 234561
rect 588126 234325 588210 234561
rect 588446 234325 588530 234561
rect 588766 234325 588874 234561
rect 587462 227561 588874 234325
rect 587462 227325 587570 227561
rect 587806 227325 587890 227561
rect 588126 227325 588210 227561
rect 588446 227325 588530 227561
rect 588766 227325 588874 227561
rect 587462 220561 588874 227325
rect 587462 220325 587570 220561
rect 587806 220325 587890 220561
rect 588126 220325 588210 220561
rect 588446 220325 588530 220561
rect 588766 220325 588874 220561
rect 587462 213561 588874 220325
rect 587462 213325 587570 213561
rect 587806 213325 587890 213561
rect 588126 213325 588210 213561
rect 588446 213325 588530 213561
rect 588766 213325 588874 213561
rect 587462 206561 588874 213325
rect 587462 206325 587570 206561
rect 587806 206325 587890 206561
rect 588126 206325 588210 206561
rect 588446 206325 588530 206561
rect 588766 206325 588874 206561
rect 587462 199561 588874 206325
rect 587462 199325 587570 199561
rect 587806 199325 587890 199561
rect 588126 199325 588210 199561
rect 588446 199325 588530 199561
rect 588766 199325 588874 199561
rect 587462 192561 588874 199325
rect 587462 192325 587570 192561
rect 587806 192325 587890 192561
rect 588126 192325 588210 192561
rect 588446 192325 588530 192561
rect 588766 192325 588874 192561
rect 587462 185561 588874 192325
rect 587462 185325 587570 185561
rect 587806 185325 587890 185561
rect 588126 185325 588210 185561
rect 588446 185325 588530 185561
rect 588766 185325 588874 185561
rect 587462 178561 588874 185325
rect 587462 178325 587570 178561
rect 587806 178325 587890 178561
rect 588126 178325 588210 178561
rect 588446 178325 588530 178561
rect 588766 178325 588874 178561
rect 587462 171561 588874 178325
rect 587462 171325 587570 171561
rect 587806 171325 587890 171561
rect 588126 171325 588210 171561
rect 588446 171325 588530 171561
rect 588766 171325 588874 171561
rect 587462 164561 588874 171325
rect 587462 164325 587570 164561
rect 587806 164325 587890 164561
rect 588126 164325 588210 164561
rect 588446 164325 588530 164561
rect 588766 164325 588874 164561
rect 587462 157561 588874 164325
rect 587462 157325 587570 157561
rect 587806 157325 587890 157561
rect 588126 157325 588210 157561
rect 588446 157325 588530 157561
rect 588766 157325 588874 157561
rect 587462 150561 588874 157325
rect 587462 150325 587570 150561
rect 587806 150325 587890 150561
rect 588126 150325 588210 150561
rect 588446 150325 588530 150561
rect 588766 150325 588874 150561
rect 587462 143561 588874 150325
rect 587462 143325 587570 143561
rect 587806 143325 587890 143561
rect 588126 143325 588210 143561
rect 588446 143325 588530 143561
rect 588766 143325 588874 143561
rect 587462 136561 588874 143325
rect 587462 136325 587570 136561
rect 587806 136325 587890 136561
rect 588126 136325 588210 136561
rect 588446 136325 588530 136561
rect 588766 136325 588874 136561
rect 587462 129561 588874 136325
rect 587462 129325 587570 129561
rect 587806 129325 587890 129561
rect 588126 129325 588210 129561
rect 588446 129325 588530 129561
rect 588766 129325 588874 129561
rect 587462 122561 588874 129325
rect 587462 122325 587570 122561
rect 587806 122325 587890 122561
rect 588126 122325 588210 122561
rect 588446 122325 588530 122561
rect 588766 122325 588874 122561
rect 587462 115561 588874 122325
rect 587462 115325 587570 115561
rect 587806 115325 587890 115561
rect 588126 115325 588210 115561
rect 588446 115325 588530 115561
rect 588766 115325 588874 115561
rect 587462 108561 588874 115325
rect 587462 108325 587570 108561
rect 587806 108325 587890 108561
rect 588126 108325 588210 108561
rect 588446 108325 588530 108561
rect 588766 108325 588874 108561
rect 587462 101561 588874 108325
rect 587462 101325 587570 101561
rect 587806 101325 587890 101561
rect 588126 101325 588210 101561
rect 588446 101325 588530 101561
rect 588766 101325 588874 101561
rect 587462 94561 588874 101325
rect 587462 94325 587570 94561
rect 587806 94325 587890 94561
rect 588126 94325 588210 94561
rect 588446 94325 588530 94561
rect 588766 94325 588874 94561
rect 587462 87561 588874 94325
rect 587462 87325 587570 87561
rect 587806 87325 587890 87561
rect 588126 87325 588210 87561
rect 588446 87325 588530 87561
rect 588766 87325 588874 87561
rect 587462 80561 588874 87325
rect 587462 80325 587570 80561
rect 587806 80325 587890 80561
rect 588126 80325 588210 80561
rect 588446 80325 588530 80561
rect 588766 80325 588874 80561
rect 587462 73561 588874 80325
rect 587462 73325 587570 73561
rect 587806 73325 587890 73561
rect 588126 73325 588210 73561
rect 588446 73325 588530 73561
rect 588766 73325 588874 73561
rect 587462 66561 588874 73325
rect 587462 66325 587570 66561
rect 587806 66325 587890 66561
rect 588126 66325 588210 66561
rect 588446 66325 588530 66561
rect 588766 66325 588874 66561
rect 587462 59561 588874 66325
rect 587462 59325 587570 59561
rect 587806 59325 587890 59561
rect 588126 59325 588210 59561
rect 588446 59325 588530 59561
rect 588766 59325 588874 59561
rect 587462 52561 588874 59325
rect 587462 52325 587570 52561
rect 587806 52325 587890 52561
rect 588126 52325 588210 52561
rect 588446 52325 588530 52561
rect 588766 52325 588874 52561
rect 587462 45561 588874 52325
rect 587462 45325 587570 45561
rect 587806 45325 587890 45561
rect 588126 45325 588210 45561
rect 588446 45325 588530 45561
rect 588766 45325 588874 45561
rect 587462 38561 588874 45325
rect 587462 38325 587570 38561
rect 587806 38325 587890 38561
rect 588126 38325 588210 38561
rect 588446 38325 588530 38561
rect 588766 38325 588874 38561
rect 587462 31561 588874 38325
rect 587462 31325 587570 31561
rect 587806 31325 587890 31561
rect 588126 31325 588210 31561
rect 588446 31325 588530 31561
rect 588766 31325 588874 31561
rect 587462 24561 588874 31325
rect 587462 24325 587570 24561
rect 587806 24325 587890 24561
rect 588126 24325 588210 24561
rect 588446 24325 588530 24561
rect 588766 24325 588874 24561
rect 587462 17561 588874 24325
rect 587462 17325 587570 17561
rect 587806 17325 587890 17561
rect 588126 17325 588210 17561
rect 588446 17325 588530 17561
rect 588766 17325 588874 17561
rect 587462 10561 588874 17325
rect 587462 10325 587570 10561
rect 587806 10325 587890 10561
rect 588126 10325 588210 10561
rect 588446 10325 588530 10561
rect 588766 10325 588874 10561
rect 587462 3561 588874 10325
rect 587462 3325 587570 3561
rect 587806 3325 587890 3561
rect 588126 3325 588210 3561
rect 588446 3325 588530 3561
rect 588766 3325 588874 3561
rect 587462 -3878 588874 3325
<< via4 >>
rect -4842 696325 -4606 696561
rect -4522 696325 -4286 696561
rect -4202 696325 -3966 696561
rect -3882 696325 -3646 696561
rect -4842 689325 -4606 689561
rect -4522 689325 -4286 689561
rect -4202 689325 -3966 689561
rect -3882 689325 -3646 689561
rect -4842 682325 -4606 682561
rect -4522 682325 -4286 682561
rect -4202 682325 -3966 682561
rect -3882 682325 -3646 682561
rect -4842 675325 -4606 675561
rect -4522 675325 -4286 675561
rect -4202 675325 -3966 675561
rect -3882 675325 -3646 675561
rect -4842 668325 -4606 668561
rect -4522 668325 -4286 668561
rect -4202 668325 -3966 668561
rect -3882 668325 -3646 668561
rect -4842 661325 -4606 661561
rect -4522 661325 -4286 661561
rect -4202 661325 -3966 661561
rect -3882 661325 -3646 661561
rect -4842 654325 -4606 654561
rect -4522 654325 -4286 654561
rect -4202 654325 -3966 654561
rect -3882 654325 -3646 654561
rect -4842 647325 -4606 647561
rect -4522 647325 -4286 647561
rect -4202 647325 -3966 647561
rect -3882 647325 -3646 647561
rect -4842 640325 -4606 640561
rect -4522 640325 -4286 640561
rect -4202 640325 -3966 640561
rect -3882 640325 -3646 640561
rect -4842 633325 -4606 633561
rect -4522 633325 -4286 633561
rect -4202 633325 -3966 633561
rect -3882 633325 -3646 633561
rect -4842 626325 -4606 626561
rect -4522 626325 -4286 626561
rect -4202 626325 -3966 626561
rect -3882 626325 -3646 626561
rect -4842 619325 -4606 619561
rect -4522 619325 -4286 619561
rect -4202 619325 -3966 619561
rect -3882 619325 -3646 619561
rect -4842 612325 -4606 612561
rect -4522 612325 -4286 612561
rect -4202 612325 -3966 612561
rect -3882 612325 -3646 612561
rect -4842 605325 -4606 605561
rect -4522 605325 -4286 605561
rect -4202 605325 -3966 605561
rect -3882 605325 -3646 605561
rect -4842 598325 -4606 598561
rect -4522 598325 -4286 598561
rect -4202 598325 -3966 598561
rect -3882 598325 -3646 598561
rect -4842 591325 -4606 591561
rect -4522 591325 -4286 591561
rect -4202 591325 -3966 591561
rect -3882 591325 -3646 591561
rect -4842 584325 -4606 584561
rect -4522 584325 -4286 584561
rect -4202 584325 -3966 584561
rect -3882 584325 -3646 584561
rect -4842 577325 -4606 577561
rect -4522 577325 -4286 577561
rect -4202 577325 -3966 577561
rect -3882 577325 -3646 577561
rect -4842 570325 -4606 570561
rect -4522 570325 -4286 570561
rect -4202 570325 -3966 570561
rect -3882 570325 -3646 570561
rect -4842 563325 -4606 563561
rect -4522 563325 -4286 563561
rect -4202 563325 -3966 563561
rect -3882 563325 -3646 563561
rect -4842 556325 -4606 556561
rect -4522 556325 -4286 556561
rect -4202 556325 -3966 556561
rect -3882 556325 -3646 556561
rect -4842 549325 -4606 549561
rect -4522 549325 -4286 549561
rect -4202 549325 -3966 549561
rect -3882 549325 -3646 549561
rect -4842 542325 -4606 542561
rect -4522 542325 -4286 542561
rect -4202 542325 -3966 542561
rect -3882 542325 -3646 542561
rect -4842 535325 -4606 535561
rect -4522 535325 -4286 535561
rect -4202 535325 -3966 535561
rect -3882 535325 -3646 535561
rect -4842 528325 -4606 528561
rect -4522 528325 -4286 528561
rect -4202 528325 -3966 528561
rect -3882 528325 -3646 528561
rect -4842 521325 -4606 521561
rect -4522 521325 -4286 521561
rect -4202 521325 -3966 521561
rect -3882 521325 -3646 521561
rect -4842 514325 -4606 514561
rect -4522 514325 -4286 514561
rect -4202 514325 -3966 514561
rect -3882 514325 -3646 514561
rect -4842 507325 -4606 507561
rect -4522 507325 -4286 507561
rect -4202 507325 -3966 507561
rect -3882 507325 -3646 507561
rect -4842 500325 -4606 500561
rect -4522 500325 -4286 500561
rect -4202 500325 -3966 500561
rect -3882 500325 -3646 500561
rect -4842 493325 -4606 493561
rect -4522 493325 -4286 493561
rect -4202 493325 -3966 493561
rect -3882 493325 -3646 493561
rect -4842 486325 -4606 486561
rect -4522 486325 -4286 486561
rect -4202 486325 -3966 486561
rect -3882 486325 -3646 486561
rect -4842 479325 -4606 479561
rect -4522 479325 -4286 479561
rect -4202 479325 -3966 479561
rect -3882 479325 -3646 479561
rect -4842 472325 -4606 472561
rect -4522 472325 -4286 472561
rect -4202 472325 -3966 472561
rect -3882 472325 -3646 472561
rect -4842 465325 -4606 465561
rect -4522 465325 -4286 465561
rect -4202 465325 -3966 465561
rect -3882 465325 -3646 465561
rect -4842 458325 -4606 458561
rect -4522 458325 -4286 458561
rect -4202 458325 -3966 458561
rect -3882 458325 -3646 458561
rect -4842 451325 -4606 451561
rect -4522 451325 -4286 451561
rect -4202 451325 -3966 451561
rect -3882 451325 -3646 451561
rect -4842 444325 -4606 444561
rect -4522 444325 -4286 444561
rect -4202 444325 -3966 444561
rect -3882 444325 -3646 444561
rect -4842 437325 -4606 437561
rect -4522 437325 -4286 437561
rect -4202 437325 -3966 437561
rect -3882 437325 -3646 437561
rect -4842 430325 -4606 430561
rect -4522 430325 -4286 430561
rect -4202 430325 -3966 430561
rect -3882 430325 -3646 430561
rect -4842 423325 -4606 423561
rect -4522 423325 -4286 423561
rect -4202 423325 -3966 423561
rect -3882 423325 -3646 423561
rect -4842 416325 -4606 416561
rect -4522 416325 -4286 416561
rect -4202 416325 -3966 416561
rect -3882 416325 -3646 416561
rect -4842 409325 -4606 409561
rect -4522 409325 -4286 409561
rect -4202 409325 -3966 409561
rect -3882 409325 -3646 409561
rect -4842 402325 -4606 402561
rect -4522 402325 -4286 402561
rect -4202 402325 -3966 402561
rect -3882 402325 -3646 402561
rect -4842 395325 -4606 395561
rect -4522 395325 -4286 395561
rect -4202 395325 -3966 395561
rect -3882 395325 -3646 395561
rect -4842 388325 -4606 388561
rect -4522 388325 -4286 388561
rect -4202 388325 -3966 388561
rect -3882 388325 -3646 388561
rect -4842 381325 -4606 381561
rect -4522 381325 -4286 381561
rect -4202 381325 -3966 381561
rect -3882 381325 -3646 381561
rect -4842 374325 -4606 374561
rect -4522 374325 -4286 374561
rect -4202 374325 -3966 374561
rect -3882 374325 -3646 374561
rect -4842 367325 -4606 367561
rect -4522 367325 -4286 367561
rect -4202 367325 -3966 367561
rect -3882 367325 -3646 367561
rect -4842 360325 -4606 360561
rect -4522 360325 -4286 360561
rect -4202 360325 -3966 360561
rect -3882 360325 -3646 360561
rect -4842 353325 -4606 353561
rect -4522 353325 -4286 353561
rect -4202 353325 -3966 353561
rect -3882 353325 -3646 353561
rect -4842 346325 -4606 346561
rect -4522 346325 -4286 346561
rect -4202 346325 -3966 346561
rect -3882 346325 -3646 346561
rect -4842 339325 -4606 339561
rect -4522 339325 -4286 339561
rect -4202 339325 -3966 339561
rect -3882 339325 -3646 339561
rect -4842 332325 -4606 332561
rect -4522 332325 -4286 332561
rect -4202 332325 -3966 332561
rect -3882 332325 -3646 332561
rect -4842 325325 -4606 325561
rect -4522 325325 -4286 325561
rect -4202 325325 -3966 325561
rect -3882 325325 -3646 325561
rect -4842 318325 -4606 318561
rect -4522 318325 -4286 318561
rect -4202 318325 -3966 318561
rect -3882 318325 -3646 318561
rect -4842 311325 -4606 311561
rect -4522 311325 -4286 311561
rect -4202 311325 -3966 311561
rect -3882 311325 -3646 311561
rect -4842 304325 -4606 304561
rect -4522 304325 -4286 304561
rect -4202 304325 -3966 304561
rect -3882 304325 -3646 304561
rect -4842 297325 -4606 297561
rect -4522 297325 -4286 297561
rect -4202 297325 -3966 297561
rect -3882 297325 -3646 297561
rect -4842 290325 -4606 290561
rect -4522 290325 -4286 290561
rect -4202 290325 -3966 290561
rect -3882 290325 -3646 290561
rect -4842 283325 -4606 283561
rect -4522 283325 -4286 283561
rect -4202 283325 -3966 283561
rect -3882 283325 -3646 283561
rect -4842 276325 -4606 276561
rect -4522 276325 -4286 276561
rect -4202 276325 -3966 276561
rect -3882 276325 -3646 276561
rect -4842 269325 -4606 269561
rect -4522 269325 -4286 269561
rect -4202 269325 -3966 269561
rect -3882 269325 -3646 269561
rect -4842 262325 -4606 262561
rect -4522 262325 -4286 262561
rect -4202 262325 -3966 262561
rect -3882 262325 -3646 262561
rect -4842 255325 -4606 255561
rect -4522 255325 -4286 255561
rect -4202 255325 -3966 255561
rect -3882 255325 -3646 255561
rect -4842 248325 -4606 248561
rect -4522 248325 -4286 248561
rect -4202 248325 -3966 248561
rect -3882 248325 -3646 248561
rect -4842 241325 -4606 241561
rect -4522 241325 -4286 241561
rect -4202 241325 -3966 241561
rect -3882 241325 -3646 241561
rect -4842 234325 -4606 234561
rect -4522 234325 -4286 234561
rect -4202 234325 -3966 234561
rect -3882 234325 -3646 234561
rect -4842 227325 -4606 227561
rect -4522 227325 -4286 227561
rect -4202 227325 -3966 227561
rect -3882 227325 -3646 227561
rect -4842 220325 -4606 220561
rect -4522 220325 -4286 220561
rect -4202 220325 -3966 220561
rect -3882 220325 -3646 220561
rect -4842 213325 -4606 213561
rect -4522 213325 -4286 213561
rect -4202 213325 -3966 213561
rect -3882 213325 -3646 213561
rect -4842 206325 -4606 206561
rect -4522 206325 -4286 206561
rect -4202 206325 -3966 206561
rect -3882 206325 -3646 206561
rect -4842 199325 -4606 199561
rect -4522 199325 -4286 199561
rect -4202 199325 -3966 199561
rect -3882 199325 -3646 199561
rect -4842 192325 -4606 192561
rect -4522 192325 -4286 192561
rect -4202 192325 -3966 192561
rect -3882 192325 -3646 192561
rect -4842 185325 -4606 185561
rect -4522 185325 -4286 185561
rect -4202 185325 -3966 185561
rect -3882 185325 -3646 185561
rect -4842 178325 -4606 178561
rect -4522 178325 -4286 178561
rect -4202 178325 -3966 178561
rect -3882 178325 -3646 178561
rect -4842 171325 -4606 171561
rect -4522 171325 -4286 171561
rect -4202 171325 -3966 171561
rect -3882 171325 -3646 171561
rect -4842 164325 -4606 164561
rect -4522 164325 -4286 164561
rect -4202 164325 -3966 164561
rect -3882 164325 -3646 164561
rect -4842 157325 -4606 157561
rect -4522 157325 -4286 157561
rect -4202 157325 -3966 157561
rect -3882 157325 -3646 157561
rect -4842 150325 -4606 150561
rect -4522 150325 -4286 150561
rect -4202 150325 -3966 150561
rect -3882 150325 -3646 150561
rect -4842 143325 -4606 143561
rect -4522 143325 -4286 143561
rect -4202 143325 -3966 143561
rect -3882 143325 -3646 143561
rect -4842 136325 -4606 136561
rect -4522 136325 -4286 136561
rect -4202 136325 -3966 136561
rect -3882 136325 -3646 136561
rect -4842 129325 -4606 129561
rect -4522 129325 -4286 129561
rect -4202 129325 -3966 129561
rect -3882 129325 -3646 129561
rect -4842 122325 -4606 122561
rect -4522 122325 -4286 122561
rect -4202 122325 -3966 122561
rect -3882 122325 -3646 122561
rect -4842 115325 -4606 115561
rect -4522 115325 -4286 115561
rect -4202 115325 -3966 115561
rect -3882 115325 -3646 115561
rect -4842 108325 -4606 108561
rect -4522 108325 -4286 108561
rect -4202 108325 -3966 108561
rect -3882 108325 -3646 108561
rect -4842 101325 -4606 101561
rect -4522 101325 -4286 101561
rect -4202 101325 -3966 101561
rect -3882 101325 -3646 101561
rect -4842 94325 -4606 94561
rect -4522 94325 -4286 94561
rect -4202 94325 -3966 94561
rect -3882 94325 -3646 94561
rect -4842 87325 -4606 87561
rect -4522 87325 -4286 87561
rect -4202 87325 -3966 87561
rect -3882 87325 -3646 87561
rect -4842 80325 -4606 80561
rect -4522 80325 -4286 80561
rect -4202 80325 -3966 80561
rect -3882 80325 -3646 80561
rect -4842 73325 -4606 73561
rect -4522 73325 -4286 73561
rect -4202 73325 -3966 73561
rect -3882 73325 -3646 73561
rect -4842 66325 -4606 66561
rect -4522 66325 -4286 66561
rect -4202 66325 -3966 66561
rect -3882 66325 -3646 66561
rect -4842 59325 -4606 59561
rect -4522 59325 -4286 59561
rect -4202 59325 -3966 59561
rect -3882 59325 -3646 59561
rect -4842 52325 -4606 52561
rect -4522 52325 -4286 52561
rect -4202 52325 -3966 52561
rect -3882 52325 -3646 52561
rect -4842 45325 -4606 45561
rect -4522 45325 -4286 45561
rect -4202 45325 -3966 45561
rect -3882 45325 -3646 45561
rect -4842 38325 -4606 38561
rect -4522 38325 -4286 38561
rect -4202 38325 -3966 38561
rect -3882 38325 -3646 38561
rect -4842 31325 -4606 31561
rect -4522 31325 -4286 31561
rect -4202 31325 -3966 31561
rect -3882 31325 -3646 31561
rect -4842 24325 -4606 24561
rect -4522 24325 -4286 24561
rect -4202 24325 -3966 24561
rect -3882 24325 -3646 24561
rect -4842 17325 -4606 17561
rect -4522 17325 -4286 17561
rect -4202 17325 -3966 17561
rect -3882 17325 -3646 17561
rect -4842 10325 -4606 10561
rect -4522 10325 -4286 10561
rect -4202 10325 -3966 10561
rect -3882 10325 -3646 10561
rect -4842 3325 -4606 3561
rect -4522 3325 -4286 3561
rect -4202 3325 -3966 3561
rect -3882 3325 -3646 3561
rect -2374 705002 -2138 705238
rect -2054 705002 -1818 705238
rect -2374 704682 -2138 704918
rect -2054 704682 -1818 704918
rect -3090 695258 -2854 695494
rect -2770 695258 -2534 695494
rect -2450 695258 -2214 695494
rect -2130 695258 -1894 695494
rect -3090 688258 -2854 688494
rect -2770 688258 -2534 688494
rect -2450 688258 -2214 688494
rect -2130 688258 -1894 688494
rect -3090 681258 -2854 681494
rect -2770 681258 -2534 681494
rect -2450 681258 -2214 681494
rect -2130 681258 -1894 681494
rect -3090 674258 -2854 674494
rect -2770 674258 -2534 674494
rect -2450 674258 -2214 674494
rect -2130 674258 -1894 674494
rect -3090 667258 -2854 667494
rect -2770 667258 -2534 667494
rect -2450 667258 -2214 667494
rect -2130 667258 -1894 667494
rect -3090 660258 -2854 660494
rect -2770 660258 -2534 660494
rect -2450 660258 -2214 660494
rect -2130 660258 -1894 660494
rect -3090 653258 -2854 653494
rect -2770 653258 -2534 653494
rect -2450 653258 -2214 653494
rect -2130 653258 -1894 653494
rect -3090 646258 -2854 646494
rect -2770 646258 -2534 646494
rect -2450 646258 -2214 646494
rect -2130 646258 -1894 646494
rect -3090 639258 -2854 639494
rect -2770 639258 -2534 639494
rect -2450 639258 -2214 639494
rect -2130 639258 -1894 639494
rect -3090 632258 -2854 632494
rect -2770 632258 -2534 632494
rect -2450 632258 -2214 632494
rect -2130 632258 -1894 632494
rect -3090 625258 -2854 625494
rect -2770 625258 -2534 625494
rect -2450 625258 -2214 625494
rect -2130 625258 -1894 625494
rect -3090 618258 -2854 618494
rect -2770 618258 -2534 618494
rect -2450 618258 -2214 618494
rect -2130 618258 -1894 618494
rect -3090 611258 -2854 611494
rect -2770 611258 -2534 611494
rect -2450 611258 -2214 611494
rect -2130 611258 -1894 611494
rect -3090 604258 -2854 604494
rect -2770 604258 -2534 604494
rect -2450 604258 -2214 604494
rect -2130 604258 -1894 604494
rect -3090 597258 -2854 597494
rect -2770 597258 -2534 597494
rect -2450 597258 -2214 597494
rect -2130 597258 -1894 597494
rect -3090 590258 -2854 590494
rect -2770 590258 -2534 590494
rect -2450 590258 -2214 590494
rect -2130 590258 -1894 590494
rect -3090 583258 -2854 583494
rect -2770 583258 -2534 583494
rect -2450 583258 -2214 583494
rect -2130 583258 -1894 583494
rect -3090 576258 -2854 576494
rect -2770 576258 -2534 576494
rect -2450 576258 -2214 576494
rect -2130 576258 -1894 576494
rect -3090 569258 -2854 569494
rect -2770 569258 -2534 569494
rect -2450 569258 -2214 569494
rect -2130 569258 -1894 569494
rect -3090 562258 -2854 562494
rect -2770 562258 -2534 562494
rect -2450 562258 -2214 562494
rect -2130 562258 -1894 562494
rect -3090 555258 -2854 555494
rect -2770 555258 -2534 555494
rect -2450 555258 -2214 555494
rect -2130 555258 -1894 555494
rect -3090 548258 -2854 548494
rect -2770 548258 -2534 548494
rect -2450 548258 -2214 548494
rect -2130 548258 -1894 548494
rect -3090 541258 -2854 541494
rect -2770 541258 -2534 541494
rect -2450 541258 -2214 541494
rect -2130 541258 -1894 541494
rect -3090 534258 -2854 534494
rect -2770 534258 -2534 534494
rect -2450 534258 -2214 534494
rect -2130 534258 -1894 534494
rect -3090 527258 -2854 527494
rect -2770 527258 -2534 527494
rect -2450 527258 -2214 527494
rect -2130 527258 -1894 527494
rect -3090 520258 -2854 520494
rect -2770 520258 -2534 520494
rect -2450 520258 -2214 520494
rect -2130 520258 -1894 520494
rect -3090 513258 -2854 513494
rect -2770 513258 -2534 513494
rect -2450 513258 -2214 513494
rect -2130 513258 -1894 513494
rect -3090 506258 -2854 506494
rect -2770 506258 -2534 506494
rect -2450 506258 -2214 506494
rect -2130 506258 -1894 506494
rect -3090 499258 -2854 499494
rect -2770 499258 -2534 499494
rect -2450 499258 -2214 499494
rect -2130 499258 -1894 499494
rect -3090 492258 -2854 492494
rect -2770 492258 -2534 492494
rect -2450 492258 -2214 492494
rect -2130 492258 -1894 492494
rect -3090 485258 -2854 485494
rect -2770 485258 -2534 485494
rect -2450 485258 -2214 485494
rect -2130 485258 -1894 485494
rect -3090 478258 -2854 478494
rect -2770 478258 -2534 478494
rect -2450 478258 -2214 478494
rect -2130 478258 -1894 478494
rect -3090 471258 -2854 471494
rect -2770 471258 -2534 471494
rect -2450 471258 -2214 471494
rect -2130 471258 -1894 471494
rect -3090 464258 -2854 464494
rect -2770 464258 -2534 464494
rect -2450 464258 -2214 464494
rect -2130 464258 -1894 464494
rect -3090 457258 -2854 457494
rect -2770 457258 -2534 457494
rect -2450 457258 -2214 457494
rect -2130 457258 -1894 457494
rect -3090 450258 -2854 450494
rect -2770 450258 -2534 450494
rect -2450 450258 -2214 450494
rect -2130 450258 -1894 450494
rect -3090 443258 -2854 443494
rect -2770 443258 -2534 443494
rect -2450 443258 -2214 443494
rect -2130 443258 -1894 443494
rect -3090 436258 -2854 436494
rect -2770 436258 -2534 436494
rect -2450 436258 -2214 436494
rect -2130 436258 -1894 436494
rect -3090 429258 -2854 429494
rect -2770 429258 -2534 429494
rect -2450 429258 -2214 429494
rect -2130 429258 -1894 429494
rect -3090 422258 -2854 422494
rect -2770 422258 -2534 422494
rect -2450 422258 -2214 422494
rect -2130 422258 -1894 422494
rect -3090 415258 -2854 415494
rect -2770 415258 -2534 415494
rect -2450 415258 -2214 415494
rect -2130 415258 -1894 415494
rect -3090 408258 -2854 408494
rect -2770 408258 -2534 408494
rect -2450 408258 -2214 408494
rect -2130 408258 -1894 408494
rect -3090 401258 -2854 401494
rect -2770 401258 -2534 401494
rect -2450 401258 -2214 401494
rect -2130 401258 -1894 401494
rect -3090 394258 -2854 394494
rect -2770 394258 -2534 394494
rect -2450 394258 -2214 394494
rect -2130 394258 -1894 394494
rect -3090 387258 -2854 387494
rect -2770 387258 -2534 387494
rect -2450 387258 -2214 387494
rect -2130 387258 -1894 387494
rect -3090 380258 -2854 380494
rect -2770 380258 -2534 380494
rect -2450 380258 -2214 380494
rect -2130 380258 -1894 380494
rect -3090 373258 -2854 373494
rect -2770 373258 -2534 373494
rect -2450 373258 -2214 373494
rect -2130 373258 -1894 373494
rect -3090 366258 -2854 366494
rect -2770 366258 -2534 366494
rect -2450 366258 -2214 366494
rect -2130 366258 -1894 366494
rect -3090 359258 -2854 359494
rect -2770 359258 -2534 359494
rect -2450 359258 -2214 359494
rect -2130 359258 -1894 359494
rect -3090 352258 -2854 352494
rect -2770 352258 -2534 352494
rect -2450 352258 -2214 352494
rect -2130 352258 -1894 352494
rect -3090 345258 -2854 345494
rect -2770 345258 -2534 345494
rect -2450 345258 -2214 345494
rect -2130 345258 -1894 345494
rect -3090 338258 -2854 338494
rect -2770 338258 -2534 338494
rect -2450 338258 -2214 338494
rect -2130 338258 -1894 338494
rect -3090 331258 -2854 331494
rect -2770 331258 -2534 331494
rect -2450 331258 -2214 331494
rect -2130 331258 -1894 331494
rect -3090 324258 -2854 324494
rect -2770 324258 -2534 324494
rect -2450 324258 -2214 324494
rect -2130 324258 -1894 324494
rect -3090 317258 -2854 317494
rect -2770 317258 -2534 317494
rect -2450 317258 -2214 317494
rect -2130 317258 -1894 317494
rect -3090 310258 -2854 310494
rect -2770 310258 -2534 310494
rect -2450 310258 -2214 310494
rect -2130 310258 -1894 310494
rect -3090 303258 -2854 303494
rect -2770 303258 -2534 303494
rect -2450 303258 -2214 303494
rect -2130 303258 -1894 303494
rect -3090 296258 -2854 296494
rect -2770 296258 -2534 296494
rect -2450 296258 -2214 296494
rect -2130 296258 -1894 296494
rect -3090 289258 -2854 289494
rect -2770 289258 -2534 289494
rect -2450 289258 -2214 289494
rect -2130 289258 -1894 289494
rect -3090 282258 -2854 282494
rect -2770 282258 -2534 282494
rect -2450 282258 -2214 282494
rect -2130 282258 -1894 282494
rect -3090 275258 -2854 275494
rect -2770 275258 -2534 275494
rect -2450 275258 -2214 275494
rect -2130 275258 -1894 275494
rect -3090 268258 -2854 268494
rect -2770 268258 -2534 268494
rect -2450 268258 -2214 268494
rect -2130 268258 -1894 268494
rect -3090 261258 -2854 261494
rect -2770 261258 -2534 261494
rect -2450 261258 -2214 261494
rect -2130 261258 -1894 261494
rect -3090 254258 -2854 254494
rect -2770 254258 -2534 254494
rect -2450 254258 -2214 254494
rect -2130 254258 -1894 254494
rect -3090 247258 -2854 247494
rect -2770 247258 -2534 247494
rect -2450 247258 -2214 247494
rect -2130 247258 -1894 247494
rect -3090 240258 -2854 240494
rect -2770 240258 -2534 240494
rect -2450 240258 -2214 240494
rect -2130 240258 -1894 240494
rect -3090 233258 -2854 233494
rect -2770 233258 -2534 233494
rect -2450 233258 -2214 233494
rect -2130 233258 -1894 233494
rect -3090 226258 -2854 226494
rect -2770 226258 -2534 226494
rect -2450 226258 -2214 226494
rect -2130 226258 -1894 226494
rect -3090 219258 -2854 219494
rect -2770 219258 -2534 219494
rect -2450 219258 -2214 219494
rect -2130 219258 -1894 219494
rect -3090 212258 -2854 212494
rect -2770 212258 -2534 212494
rect -2450 212258 -2214 212494
rect -2130 212258 -1894 212494
rect -3090 205258 -2854 205494
rect -2770 205258 -2534 205494
rect -2450 205258 -2214 205494
rect -2130 205258 -1894 205494
rect -3090 198258 -2854 198494
rect -2770 198258 -2534 198494
rect -2450 198258 -2214 198494
rect -2130 198258 -1894 198494
rect -3090 191258 -2854 191494
rect -2770 191258 -2534 191494
rect -2450 191258 -2214 191494
rect -2130 191258 -1894 191494
rect -3090 184258 -2854 184494
rect -2770 184258 -2534 184494
rect -2450 184258 -2214 184494
rect -2130 184258 -1894 184494
rect -3090 177258 -2854 177494
rect -2770 177258 -2534 177494
rect -2450 177258 -2214 177494
rect -2130 177258 -1894 177494
rect -3090 170258 -2854 170494
rect -2770 170258 -2534 170494
rect -2450 170258 -2214 170494
rect -2130 170258 -1894 170494
rect -3090 163258 -2854 163494
rect -2770 163258 -2534 163494
rect -2450 163258 -2214 163494
rect -2130 163258 -1894 163494
rect -3090 156258 -2854 156494
rect -2770 156258 -2534 156494
rect -2450 156258 -2214 156494
rect -2130 156258 -1894 156494
rect -3090 149258 -2854 149494
rect -2770 149258 -2534 149494
rect -2450 149258 -2214 149494
rect -2130 149258 -1894 149494
rect -3090 142258 -2854 142494
rect -2770 142258 -2534 142494
rect -2450 142258 -2214 142494
rect -2130 142258 -1894 142494
rect -3090 135258 -2854 135494
rect -2770 135258 -2534 135494
rect -2450 135258 -2214 135494
rect -2130 135258 -1894 135494
rect -3090 128258 -2854 128494
rect -2770 128258 -2534 128494
rect -2450 128258 -2214 128494
rect -2130 128258 -1894 128494
rect -3090 121258 -2854 121494
rect -2770 121258 -2534 121494
rect -2450 121258 -2214 121494
rect -2130 121258 -1894 121494
rect -3090 114258 -2854 114494
rect -2770 114258 -2534 114494
rect -2450 114258 -2214 114494
rect -2130 114258 -1894 114494
rect -3090 107258 -2854 107494
rect -2770 107258 -2534 107494
rect -2450 107258 -2214 107494
rect -2130 107258 -1894 107494
rect -3090 100258 -2854 100494
rect -2770 100258 -2534 100494
rect -2450 100258 -2214 100494
rect -2130 100258 -1894 100494
rect -3090 93258 -2854 93494
rect -2770 93258 -2534 93494
rect -2450 93258 -2214 93494
rect -2130 93258 -1894 93494
rect -3090 86258 -2854 86494
rect -2770 86258 -2534 86494
rect -2450 86258 -2214 86494
rect -2130 86258 -1894 86494
rect -3090 79258 -2854 79494
rect -2770 79258 -2534 79494
rect -2450 79258 -2214 79494
rect -2130 79258 -1894 79494
rect -3090 72258 -2854 72494
rect -2770 72258 -2534 72494
rect -2450 72258 -2214 72494
rect -2130 72258 -1894 72494
rect -3090 65258 -2854 65494
rect -2770 65258 -2534 65494
rect -2450 65258 -2214 65494
rect -2130 65258 -1894 65494
rect -3090 58258 -2854 58494
rect -2770 58258 -2534 58494
rect -2450 58258 -2214 58494
rect -2130 58258 -1894 58494
rect -3090 51258 -2854 51494
rect -2770 51258 -2534 51494
rect -2450 51258 -2214 51494
rect -2130 51258 -1894 51494
rect -3090 44258 -2854 44494
rect -2770 44258 -2534 44494
rect -2450 44258 -2214 44494
rect -2130 44258 -1894 44494
rect -3090 37258 -2854 37494
rect -2770 37258 -2534 37494
rect -2450 37258 -2214 37494
rect -2130 37258 -1894 37494
rect -3090 30258 -2854 30494
rect -2770 30258 -2534 30494
rect -2450 30258 -2214 30494
rect -2130 30258 -1894 30494
rect -3090 23258 -2854 23494
rect -2770 23258 -2534 23494
rect -2450 23258 -2214 23494
rect -2130 23258 -1894 23494
rect -3090 16258 -2854 16494
rect -2770 16258 -2534 16494
rect -2450 16258 -2214 16494
rect -2130 16258 -1894 16494
rect -3090 9258 -2854 9494
rect -2770 9258 -2534 9494
rect -2450 9258 -2214 9494
rect -2130 9258 -1894 9494
rect -3090 2258 -2854 2494
rect -2770 2258 -2534 2494
rect -2450 2258 -2214 2494
rect -2130 2258 -1894 2494
rect -2374 -982 -2138 -746
rect -2054 -982 -1818 -746
rect -2374 -1302 -2138 -1066
rect -2054 -1302 -1818 -1066
rect 1186 705002 1422 705238
rect 1186 704682 1422 704918
rect 1186 695258 1422 695494
rect 1186 688258 1422 688494
rect 1186 681258 1422 681494
rect 1186 674258 1422 674494
rect 1186 667258 1422 667494
rect 1186 660258 1422 660494
rect 1186 653258 1422 653494
rect 1186 646258 1422 646494
rect 1186 639258 1422 639494
rect 1186 632258 1422 632494
rect 1186 625258 1422 625494
rect 1186 618258 1422 618494
rect 1186 611258 1422 611494
rect 1186 604258 1422 604494
rect 1186 597258 1422 597494
rect 1186 590258 1422 590494
rect 1186 583258 1422 583494
rect 1186 576258 1422 576494
rect 1186 569258 1422 569494
rect 1186 562258 1422 562494
rect 1186 555258 1422 555494
rect 1186 548258 1422 548494
rect 1186 541258 1422 541494
rect 1186 534258 1422 534494
rect 1186 527258 1422 527494
rect 1186 520258 1422 520494
rect 1186 513258 1422 513494
rect 1186 506258 1422 506494
rect 1186 499258 1422 499494
rect 1186 492258 1422 492494
rect 1186 485258 1422 485494
rect 1186 478258 1422 478494
rect 1186 471258 1422 471494
rect 1186 464258 1422 464494
rect 1186 457258 1422 457494
rect 1186 450258 1422 450494
rect 1186 443258 1422 443494
rect 1186 436258 1422 436494
rect 1186 429258 1422 429494
rect 1186 422258 1422 422494
rect 1186 415258 1422 415494
rect 1186 408258 1422 408494
rect 1186 401258 1422 401494
rect 1186 394258 1422 394494
rect 1186 387258 1422 387494
rect 1186 380258 1422 380494
rect 1186 373258 1422 373494
rect 1186 366258 1422 366494
rect 1186 359258 1422 359494
rect 1186 352258 1422 352494
rect 1186 345258 1422 345494
rect 1186 338258 1422 338494
rect 1186 331258 1422 331494
rect 1186 324258 1422 324494
rect 1186 317258 1422 317494
rect 1186 310258 1422 310494
rect 1186 303258 1422 303494
rect 1186 296258 1422 296494
rect 1186 289258 1422 289494
rect 1186 282258 1422 282494
rect 1186 275258 1422 275494
rect 1186 268258 1422 268494
rect 1186 261258 1422 261494
rect 1186 254258 1422 254494
rect 1186 247258 1422 247494
rect 1186 240258 1422 240494
rect 1186 233258 1422 233494
rect 1186 226258 1422 226494
rect 1186 219258 1422 219494
rect 1186 212258 1422 212494
rect 1186 205258 1422 205494
rect 1186 198258 1422 198494
rect 1186 191258 1422 191494
rect 1186 184258 1422 184494
rect 1186 177258 1422 177494
rect 1186 170258 1422 170494
rect 1186 163258 1422 163494
rect 1186 156258 1422 156494
rect 1186 149258 1422 149494
rect 1186 142258 1422 142494
rect 1186 135258 1422 135494
rect 1186 128258 1422 128494
rect 1186 121258 1422 121494
rect 1186 114258 1422 114494
rect 1186 107258 1422 107494
rect 1186 100258 1422 100494
rect 1186 93258 1422 93494
rect 1186 86258 1422 86494
rect 1186 79258 1422 79494
rect 1186 72258 1422 72494
rect 1186 65258 1422 65494
rect 1186 58258 1422 58494
rect 1186 51258 1422 51494
rect 1186 44258 1422 44494
rect 1186 37258 1422 37494
rect 1186 30258 1422 30494
rect 1186 23258 1422 23494
rect 1186 16258 1422 16494
rect 1186 9258 1422 9494
rect 1186 2258 1422 2494
rect 1186 -982 1422 -746
rect 1186 -1302 1422 -1066
rect 2918 705962 3154 706198
rect 2918 705642 3154 705878
rect 2918 696325 3154 696561
rect 2918 689325 3154 689561
rect 2918 682325 3154 682561
rect 2918 675325 3154 675561
rect 2918 668325 3154 668561
rect 2918 661325 3154 661561
rect 2918 654325 3154 654561
rect 2918 647325 3154 647561
rect 2918 640325 3154 640561
rect 2918 633325 3154 633561
rect 2918 626325 3154 626561
rect 2918 619325 3154 619561
rect 2918 612325 3154 612561
rect 2918 605325 3154 605561
rect 2918 598325 3154 598561
rect 2918 591325 3154 591561
rect 2918 584325 3154 584561
rect 2918 577325 3154 577561
rect 2918 570325 3154 570561
rect 2918 563325 3154 563561
rect 2918 556325 3154 556561
rect 2918 549325 3154 549561
rect 2918 542325 3154 542561
rect 2918 535325 3154 535561
rect 2918 528325 3154 528561
rect 2918 521325 3154 521561
rect 2918 514325 3154 514561
rect 2918 507325 3154 507561
rect 2918 500325 3154 500561
rect 2918 493325 3154 493561
rect 2918 486325 3154 486561
rect 2918 479325 3154 479561
rect 2918 472325 3154 472561
rect 2918 465325 3154 465561
rect 2918 458325 3154 458561
rect 2918 451325 3154 451561
rect 2918 444325 3154 444561
rect 2918 437325 3154 437561
rect 2918 430325 3154 430561
rect 2918 423325 3154 423561
rect 2918 416325 3154 416561
rect 2918 409325 3154 409561
rect 2918 402325 3154 402561
rect 2918 395325 3154 395561
rect 2918 388325 3154 388561
rect 2918 381325 3154 381561
rect 2918 374325 3154 374561
rect 2918 367325 3154 367561
rect 2918 360325 3154 360561
rect 2918 353325 3154 353561
rect 2918 346325 3154 346561
rect 2918 339325 3154 339561
rect 2918 332325 3154 332561
rect 2918 325325 3154 325561
rect 2918 318325 3154 318561
rect 2918 311325 3154 311561
rect 2918 304325 3154 304561
rect 2918 297325 3154 297561
rect 2918 290325 3154 290561
rect 2918 283325 3154 283561
rect 2918 276325 3154 276561
rect 2918 269325 3154 269561
rect 2918 262325 3154 262561
rect 2918 255325 3154 255561
rect 2918 248325 3154 248561
rect 2918 241325 3154 241561
rect 2918 234325 3154 234561
rect 2918 227325 3154 227561
rect 2918 220325 3154 220561
rect 2918 213325 3154 213561
rect 2918 206325 3154 206561
rect 2918 199325 3154 199561
rect 2918 192325 3154 192561
rect 2918 185325 3154 185561
rect 2918 178325 3154 178561
rect 2918 171325 3154 171561
rect 2918 164325 3154 164561
rect 2918 157325 3154 157561
rect 2918 150325 3154 150561
rect 2918 143325 3154 143561
rect 2918 136325 3154 136561
rect 2918 129325 3154 129561
rect 2918 122325 3154 122561
rect 2918 115325 3154 115561
rect 2918 108325 3154 108561
rect 2918 101325 3154 101561
rect 2918 94325 3154 94561
rect 2918 87325 3154 87561
rect 2918 80325 3154 80561
rect 2918 73325 3154 73561
rect 2918 66325 3154 66561
rect 2918 59325 3154 59561
rect 2918 52325 3154 52561
rect 2918 45325 3154 45561
rect 2918 38325 3154 38561
rect 2918 31325 3154 31561
rect 2918 24325 3154 24561
rect 2918 17325 3154 17561
rect 2918 10325 3154 10561
rect 2918 3325 3154 3561
rect 2918 -1942 3154 -1706
rect 2918 -2262 3154 -2026
rect 8186 705002 8422 705238
rect 8186 704682 8422 704918
rect 8186 695258 8422 695494
rect 8186 688258 8422 688494
rect 8186 681258 8422 681494
rect 8186 674258 8422 674494
rect 8186 667258 8422 667494
rect 8186 660258 8422 660494
rect 8186 653258 8422 653494
rect 8186 646258 8422 646494
rect 8186 639258 8422 639494
rect 8186 632258 8422 632494
rect 8186 625258 8422 625494
rect 8186 618258 8422 618494
rect 8186 611258 8422 611494
rect 8186 604258 8422 604494
rect 8186 597258 8422 597494
rect 8186 590258 8422 590494
rect 8186 583258 8422 583494
rect 8186 576258 8422 576494
rect 8186 569258 8422 569494
rect 8186 562258 8422 562494
rect 8186 555258 8422 555494
rect 8186 548258 8422 548494
rect 8186 541258 8422 541494
rect 8186 534258 8422 534494
rect 8186 527258 8422 527494
rect 8186 520258 8422 520494
rect 8186 513258 8422 513494
rect 8186 506258 8422 506494
rect 8186 499258 8422 499494
rect 8186 492258 8422 492494
rect 8186 485258 8422 485494
rect 8186 478258 8422 478494
rect 8186 471258 8422 471494
rect 8186 464258 8422 464494
rect 8186 457258 8422 457494
rect 8186 450258 8422 450494
rect 8186 443258 8422 443494
rect 8186 436258 8422 436494
rect 8186 429258 8422 429494
rect 8186 422258 8422 422494
rect 8186 415258 8422 415494
rect 8186 408258 8422 408494
rect 8186 401258 8422 401494
rect 8186 394258 8422 394494
rect 8186 387258 8422 387494
rect 8186 380258 8422 380494
rect 8186 373258 8422 373494
rect 8186 366258 8422 366494
rect 8186 359258 8422 359494
rect 8186 352258 8422 352494
rect 8186 345258 8422 345494
rect 8186 338258 8422 338494
rect 8186 331258 8422 331494
rect 8186 324258 8422 324494
rect 8186 317258 8422 317494
rect 8186 310258 8422 310494
rect 8186 303258 8422 303494
rect 8186 296258 8422 296494
rect 8186 289258 8422 289494
rect 8186 282258 8422 282494
rect 8186 275258 8422 275494
rect 8186 268258 8422 268494
rect 8186 261258 8422 261494
rect 8186 254258 8422 254494
rect 8186 247258 8422 247494
rect 8186 240258 8422 240494
rect 8186 233258 8422 233494
rect 8186 226258 8422 226494
rect 8186 219258 8422 219494
rect 8186 212258 8422 212494
rect 8186 205258 8422 205494
rect 8186 198258 8422 198494
rect 8186 191258 8422 191494
rect 8186 184258 8422 184494
rect 8186 177258 8422 177494
rect 8186 170258 8422 170494
rect 8186 163258 8422 163494
rect 8186 156258 8422 156494
rect 8186 149258 8422 149494
rect 8186 142258 8422 142494
rect 8186 135258 8422 135494
rect 8186 128258 8422 128494
rect 8186 121258 8422 121494
rect 8186 114258 8422 114494
rect 8186 107258 8422 107494
rect 8186 100258 8422 100494
rect 8186 93258 8422 93494
rect 8186 86258 8422 86494
rect 8186 79258 8422 79494
rect 8186 72258 8422 72494
rect 8186 65258 8422 65494
rect 8186 58258 8422 58494
rect 8186 51258 8422 51494
rect 8186 44258 8422 44494
rect 8186 37258 8422 37494
rect 8186 30258 8422 30494
rect 8186 23258 8422 23494
rect 8186 16258 8422 16494
rect 8186 9258 8422 9494
rect 8186 2258 8422 2494
rect 8186 -982 8422 -746
rect 8186 -1302 8422 -1066
rect 9918 705962 10154 706198
rect 9918 705642 10154 705878
rect 9918 696325 10154 696561
rect 9918 689325 10154 689561
rect 9918 682325 10154 682561
rect 9918 675325 10154 675561
rect 9918 668325 10154 668561
rect 9918 661325 10154 661561
rect 9918 654325 10154 654561
rect 9918 647325 10154 647561
rect 9918 640325 10154 640561
rect 9918 633325 10154 633561
rect 9918 626325 10154 626561
rect 9918 619325 10154 619561
rect 9918 612325 10154 612561
rect 9918 605325 10154 605561
rect 9918 598325 10154 598561
rect 9918 591325 10154 591561
rect 9918 584325 10154 584561
rect 9918 577325 10154 577561
rect 9918 570325 10154 570561
rect 9918 563325 10154 563561
rect 9918 556325 10154 556561
rect 9918 549325 10154 549561
rect 9918 542325 10154 542561
rect 9918 535325 10154 535561
rect 9918 528325 10154 528561
rect 9918 521325 10154 521561
rect 9918 514325 10154 514561
rect 9918 507325 10154 507561
rect 9918 500325 10154 500561
rect 9918 493325 10154 493561
rect 9918 486325 10154 486561
rect 9918 479325 10154 479561
rect 9918 472325 10154 472561
rect 9918 465325 10154 465561
rect 9918 458325 10154 458561
rect 9918 451325 10154 451561
rect 9918 444325 10154 444561
rect 9918 437325 10154 437561
rect 9918 430325 10154 430561
rect 9918 423325 10154 423561
rect 9918 416325 10154 416561
rect 9918 409325 10154 409561
rect 9918 402325 10154 402561
rect 9918 395325 10154 395561
rect 9918 388325 10154 388561
rect 9918 381325 10154 381561
rect 9918 374325 10154 374561
rect 9918 367325 10154 367561
rect 9918 360325 10154 360561
rect 9918 353325 10154 353561
rect 9918 346325 10154 346561
rect 9918 339325 10154 339561
rect 9918 332325 10154 332561
rect 9918 325325 10154 325561
rect 9918 318325 10154 318561
rect 9918 311325 10154 311561
rect 9918 304325 10154 304561
rect 9918 297325 10154 297561
rect 9918 290325 10154 290561
rect 9918 283325 10154 283561
rect 9918 276325 10154 276561
rect 9918 269325 10154 269561
rect 9918 262325 10154 262561
rect 9918 255325 10154 255561
rect 9918 248325 10154 248561
rect 9918 241325 10154 241561
rect 9918 234325 10154 234561
rect 9918 227325 10154 227561
rect 9918 220325 10154 220561
rect 9918 213325 10154 213561
rect 9918 206325 10154 206561
rect 9918 199325 10154 199561
rect 9918 192325 10154 192561
rect 9918 185325 10154 185561
rect 9918 178325 10154 178561
rect 9918 171325 10154 171561
rect 9918 164325 10154 164561
rect 9918 157325 10154 157561
rect 9918 150325 10154 150561
rect 9918 143325 10154 143561
rect 9918 136325 10154 136561
rect 9918 129325 10154 129561
rect 9918 122325 10154 122561
rect 9918 115325 10154 115561
rect 9918 108325 10154 108561
rect 9918 101325 10154 101561
rect 9918 94325 10154 94561
rect 9918 87325 10154 87561
rect 9918 80325 10154 80561
rect 9918 73325 10154 73561
rect 9918 66325 10154 66561
rect 9918 59325 10154 59561
rect 9918 52325 10154 52561
rect 9918 45325 10154 45561
rect 9918 38325 10154 38561
rect 9918 31325 10154 31561
rect 9918 24325 10154 24561
rect 9918 17325 10154 17561
rect 9918 10325 10154 10561
rect 9918 3325 10154 3561
rect 9918 -1942 10154 -1706
rect 9918 -2262 10154 -2026
rect 15186 705002 15422 705238
rect 15186 704682 15422 704918
rect 15186 695258 15422 695494
rect 15186 688258 15422 688494
rect 15186 681258 15422 681494
rect 15186 674258 15422 674494
rect 15186 667258 15422 667494
rect 15186 660258 15422 660494
rect 15186 653258 15422 653494
rect 15186 646258 15422 646494
rect 15186 639258 15422 639494
rect 15186 632258 15422 632494
rect 15186 625258 15422 625494
rect 15186 618258 15422 618494
rect 15186 611258 15422 611494
rect 15186 604258 15422 604494
rect 15186 597258 15422 597494
rect 15186 590258 15422 590494
rect 15186 583258 15422 583494
rect 15186 576258 15422 576494
rect 15186 569258 15422 569494
rect 15186 562258 15422 562494
rect 15186 555258 15422 555494
rect 15186 548258 15422 548494
rect 15186 541258 15422 541494
rect 15186 534258 15422 534494
rect 15186 527258 15422 527494
rect 15186 520258 15422 520494
rect 15186 513258 15422 513494
rect 15186 506258 15422 506494
rect 15186 499258 15422 499494
rect 15186 492258 15422 492494
rect 15186 485258 15422 485494
rect 15186 478258 15422 478494
rect 15186 471258 15422 471494
rect 15186 464258 15422 464494
rect 15186 457258 15422 457494
rect 15186 450258 15422 450494
rect 15186 443258 15422 443494
rect 15186 436258 15422 436494
rect 15186 429258 15422 429494
rect 15186 422258 15422 422494
rect 15186 415258 15422 415494
rect 15186 408258 15422 408494
rect 15186 401258 15422 401494
rect 15186 394258 15422 394494
rect 15186 387258 15422 387494
rect 15186 380258 15422 380494
rect 15186 373258 15422 373494
rect 15186 366258 15422 366494
rect 15186 359258 15422 359494
rect 15186 352258 15422 352494
rect 15186 345258 15422 345494
rect 15186 338258 15422 338494
rect 15186 331258 15422 331494
rect 15186 324258 15422 324494
rect 15186 317258 15422 317494
rect 15186 310258 15422 310494
rect 15186 303258 15422 303494
rect 15186 296258 15422 296494
rect 15186 289258 15422 289494
rect 15186 282258 15422 282494
rect 15186 275258 15422 275494
rect 15186 268258 15422 268494
rect 15186 261258 15422 261494
rect 15186 254258 15422 254494
rect 15186 247258 15422 247494
rect 15186 240258 15422 240494
rect 15186 233258 15422 233494
rect 15186 226258 15422 226494
rect 15186 219258 15422 219494
rect 15186 212258 15422 212494
rect 15186 205258 15422 205494
rect 15186 198258 15422 198494
rect 15186 191258 15422 191494
rect 15186 184258 15422 184494
rect 15186 177258 15422 177494
rect 15186 170258 15422 170494
rect 15186 163258 15422 163494
rect 15186 156258 15422 156494
rect 15186 149258 15422 149494
rect 15186 142258 15422 142494
rect 15186 135258 15422 135494
rect 15186 128258 15422 128494
rect 15186 121258 15422 121494
rect 15186 114258 15422 114494
rect 15186 107258 15422 107494
rect 15186 100258 15422 100494
rect 15186 93258 15422 93494
rect 15186 86258 15422 86494
rect 15186 79258 15422 79494
rect 15186 72258 15422 72494
rect 15186 65258 15422 65494
rect 15186 58258 15422 58494
rect 15186 51258 15422 51494
rect 15186 44258 15422 44494
rect 15186 37258 15422 37494
rect 15186 30258 15422 30494
rect 15186 23258 15422 23494
rect 15186 16258 15422 16494
rect 15186 9258 15422 9494
rect 15186 2258 15422 2494
rect 15186 -982 15422 -746
rect 15186 -1302 15422 -1066
rect 16918 705962 17154 706198
rect 16918 705642 17154 705878
rect 16918 696325 17154 696561
rect 16918 689325 17154 689561
rect 16918 682325 17154 682561
rect 16918 675325 17154 675561
rect 16918 668325 17154 668561
rect 16918 661325 17154 661561
rect 16918 654325 17154 654561
rect 16918 647325 17154 647561
rect 16918 640325 17154 640561
rect 16918 633325 17154 633561
rect 16918 626325 17154 626561
rect 16918 619325 17154 619561
rect 16918 612325 17154 612561
rect 16918 605325 17154 605561
rect 16918 598325 17154 598561
rect 16918 591325 17154 591561
rect 16918 584325 17154 584561
rect 16918 577325 17154 577561
rect 16918 570325 17154 570561
rect 16918 563325 17154 563561
rect 16918 556325 17154 556561
rect 16918 549325 17154 549561
rect 16918 542325 17154 542561
rect 16918 535325 17154 535561
rect 16918 528325 17154 528561
rect 16918 521325 17154 521561
rect 16918 514325 17154 514561
rect 16918 507325 17154 507561
rect 16918 500325 17154 500561
rect 16918 493325 17154 493561
rect 16918 486325 17154 486561
rect 16918 479325 17154 479561
rect 16918 472325 17154 472561
rect 16918 465325 17154 465561
rect 16918 458325 17154 458561
rect 16918 451325 17154 451561
rect 16918 444325 17154 444561
rect 16918 437325 17154 437561
rect 16918 430325 17154 430561
rect 16918 423325 17154 423561
rect 16918 416325 17154 416561
rect 16918 409325 17154 409561
rect 16918 402325 17154 402561
rect 16918 395325 17154 395561
rect 16918 388325 17154 388561
rect 16918 381325 17154 381561
rect 16918 374325 17154 374561
rect 16918 367325 17154 367561
rect 16918 360325 17154 360561
rect 16918 353325 17154 353561
rect 16918 346325 17154 346561
rect 16918 339325 17154 339561
rect 16918 332325 17154 332561
rect 16918 325325 17154 325561
rect 16918 318325 17154 318561
rect 16918 311325 17154 311561
rect 16918 304325 17154 304561
rect 16918 297325 17154 297561
rect 16918 290325 17154 290561
rect 16918 283325 17154 283561
rect 16918 276325 17154 276561
rect 16918 269325 17154 269561
rect 16918 262325 17154 262561
rect 16918 255325 17154 255561
rect 16918 248325 17154 248561
rect 16918 241325 17154 241561
rect 16918 234325 17154 234561
rect 16918 227325 17154 227561
rect 16918 220325 17154 220561
rect 16918 213325 17154 213561
rect 16918 206325 17154 206561
rect 16918 199325 17154 199561
rect 16918 192325 17154 192561
rect 16918 185325 17154 185561
rect 16918 178325 17154 178561
rect 16918 171325 17154 171561
rect 16918 164325 17154 164561
rect 16918 157325 17154 157561
rect 16918 150325 17154 150561
rect 16918 143325 17154 143561
rect 16918 136325 17154 136561
rect 16918 129325 17154 129561
rect 16918 122325 17154 122561
rect 16918 115325 17154 115561
rect 16918 108325 17154 108561
rect 16918 101325 17154 101561
rect 16918 94325 17154 94561
rect 16918 87325 17154 87561
rect 16918 80325 17154 80561
rect 16918 73325 17154 73561
rect 16918 66325 17154 66561
rect 16918 59325 17154 59561
rect 16918 52325 17154 52561
rect 16918 45325 17154 45561
rect 16918 38325 17154 38561
rect 16918 31325 17154 31561
rect 16918 24325 17154 24561
rect 16918 17325 17154 17561
rect 16918 10325 17154 10561
rect 16918 3325 17154 3561
rect 16918 -1942 17154 -1706
rect 16918 -2262 17154 -2026
rect 22186 705002 22422 705238
rect 22186 704682 22422 704918
rect 22186 695258 22422 695494
rect 22186 688258 22422 688494
rect 22186 681258 22422 681494
rect 22186 674258 22422 674494
rect 22186 667258 22422 667494
rect 22186 660258 22422 660494
rect 22186 653258 22422 653494
rect 22186 646258 22422 646494
rect 22186 639258 22422 639494
rect 22186 632258 22422 632494
rect 22186 625258 22422 625494
rect 22186 618258 22422 618494
rect 22186 611258 22422 611494
rect 22186 604258 22422 604494
rect 22186 597258 22422 597494
rect 22186 590258 22422 590494
rect 22186 583258 22422 583494
rect 22186 576258 22422 576494
rect 22186 569258 22422 569494
rect 22186 562258 22422 562494
rect 22186 555258 22422 555494
rect 22186 548258 22422 548494
rect 22186 541258 22422 541494
rect 22186 534258 22422 534494
rect 22186 527258 22422 527494
rect 22186 520258 22422 520494
rect 22186 513258 22422 513494
rect 22186 506258 22422 506494
rect 22186 499258 22422 499494
rect 22186 492258 22422 492494
rect 22186 485258 22422 485494
rect 22186 478258 22422 478494
rect 22186 471258 22422 471494
rect 22186 464258 22422 464494
rect 22186 457258 22422 457494
rect 22186 450258 22422 450494
rect 22186 443258 22422 443494
rect 22186 436258 22422 436494
rect 22186 429258 22422 429494
rect 22186 422258 22422 422494
rect 22186 415258 22422 415494
rect 22186 408258 22422 408494
rect 22186 401258 22422 401494
rect 22186 394258 22422 394494
rect 22186 387258 22422 387494
rect 22186 380258 22422 380494
rect 22186 373258 22422 373494
rect 22186 366258 22422 366494
rect 22186 359258 22422 359494
rect 22186 352258 22422 352494
rect 22186 345258 22422 345494
rect 22186 338258 22422 338494
rect 22186 331258 22422 331494
rect 22186 324258 22422 324494
rect 22186 317258 22422 317494
rect 22186 310258 22422 310494
rect 22186 303258 22422 303494
rect 22186 296258 22422 296494
rect 22186 289258 22422 289494
rect 22186 282258 22422 282494
rect 22186 275258 22422 275494
rect 22186 268258 22422 268494
rect 22186 261258 22422 261494
rect 22186 254258 22422 254494
rect 22186 247258 22422 247494
rect 22186 240258 22422 240494
rect 22186 233258 22422 233494
rect 22186 226258 22422 226494
rect 22186 219258 22422 219494
rect 22186 212258 22422 212494
rect 22186 205258 22422 205494
rect 22186 198258 22422 198494
rect 22186 191258 22422 191494
rect 22186 184258 22422 184494
rect 22186 177258 22422 177494
rect 22186 170258 22422 170494
rect 22186 163258 22422 163494
rect 22186 156258 22422 156494
rect 22186 149258 22422 149494
rect 22186 142258 22422 142494
rect 22186 135258 22422 135494
rect 22186 128258 22422 128494
rect 22186 121258 22422 121494
rect 22186 114258 22422 114494
rect 22186 107258 22422 107494
rect 22186 100258 22422 100494
rect 22186 93258 22422 93494
rect 22186 86258 22422 86494
rect 22186 79258 22422 79494
rect 22186 72258 22422 72494
rect 22186 65258 22422 65494
rect 22186 58258 22422 58494
rect 22186 51258 22422 51494
rect 22186 44258 22422 44494
rect 22186 37258 22422 37494
rect 22186 30258 22422 30494
rect 22186 23258 22422 23494
rect 22186 16258 22422 16494
rect 22186 9258 22422 9494
rect 22186 2258 22422 2494
rect 22186 -982 22422 -746
rect 22186 -1302 22422 -1066
rect 23918 705962 24154 706198
rect 23918 705642 24154 705878
rect 23918 696325 24154 696561
rect 23918 689325 24154 689561
rect 23918 682325 24154 682561
rect 23918 675325 24154 675561
rect 23918 668325 24154 668561
rect 23918 661325 24154 661561
rect 23918 654325 24154 654561
rect 23918 647325 24154 647561
rect 23918 640325 24154 640561
rect 23918 633325 24154 633561
rect 23918 626325 24154 626561
rect 23918 619325 24154 619561
rect 23918 612325 24154 612561
rect 23918 605325 24154 605561
rect 23918 598325 24154 598561
rect 23918 591325 24154 591561
rect 23918 584325 24154 584561
rect 23918 577325 24154 577561
rect 23918 570325 24154 570561
rect 23918 563325 24154 563561
rect 23918 556325 24154 556561
rect 23918 549325 24154 549561
rect 23918 542325 24154 542561
rect 23918 535325 24154 535561
rect 23918 528325 24154 528561
rect 23918 521325 24154 521561
rect 23918 514325 24154 514561
rect 23918 507325 24154 507561
rect 23918 500325 24154 500561
rect 23918 493325 24154 493561
rect 23918 486325 24154 486561
rect 23918 479325 24154 479561
rect 23918 472325 24154 472561
rect 23918 465325 24154 465561
rect 23918 458325 24154 458561
rect 23918 451325 24154 451561
rect 23918 444325 24154 444561
rect 23918 437325 24154 437561
rect 23918 430325 24154 430561
rect 23918 423325 24154 423561
rect 23918 416325 24154 416561
rect 23918 409325 24154 409561
rect 23918 402325 24154 402561
rect 23918 395325 24154 395561
rect 23918 388325 24154 388561
rect 23918 381325 24154 381561
rect 23918 374325 24154 374561
rect 23918 367325 24154 367561
rect 23918 360325 24154 360561
rect 23918 353325 24154 353561
rect 23918 346325 24154 346561
rect 23918 339325 24154 339561
rect 23918 332325 24154 332561
rect 23918 325325 24154 325561
rect 23918 318325 24154 318561
rect 23918 311325 24154 311561
rect 23918 304325 24154 304561
rect 23918 297325 24154 297561
rect 23918 290325 24154 290561
rect 23918 283325 24154 283561
rect 23918 276325 24154 276561
rect 23918 269325 24154 269561
rect 23918 262325 24154 262561
rect 23918 255325 24154 255561
rect 23918 248325 24154 248561
rect 23918 241325 24154 241561
rect 23918 234325 24154 234561
rect 23918 227325 24154 227561
rect 23918 220325 24154 220561
rect 23918 213325 24154 213561
rect 23918 206325 24154 206561
rect 23918 199325 24154 199561
rect 23918 192325 24154 192561
rect 23918 185325 24154 185561
rect 23918 178325 24154 178561
rect 23918 171325 24154 171561
rect 23918 164325 24154 164561
rect 23918 157325 24154 157561
rect 23918 150325 24154 150561
rect 23918 143325 24154 143561
rect 23918 136325 24154 136561
rect 23918 129325 24154 129561
rect 23918 122325 24154 122561
rect 23918 115325 24154 115561
rect 23918 108325 24154 108561
rect 23918 101325 24154 101561
rect 23918 94325 24154 94561
rect 23918 87325 24154 87561
rect 23918 80325 24154 80561
rect 23918 73325 24154 73561
rect 23918 66325 24154 66561
rect 23918 59325 24154 59561
rect 23918 52325 24154 52561
rect 23918 45325 24154 45561
rect 23918 38325 24154 38561
rect 23918 31325 24154 31561
rect 23918 24325 24154 24561
rect 23918 17325 24154 17561
rect 23918 10325 24154 10561
rect 23918 3325 24154 3561
rect 23918 -1942 24154 -1706
rect 23918 -2262 24154 -2026
rect 29186 705002 29422 705238
rect 29186 704682 29422 704918
rect 29186 695258 29422 695494
rect 29186 688258 29422 688494
rect 29186 681258 29422 681494
rect 29186 674258 29422 674494
rect 29186 667258 29422 667494
rect 29186 660258 29422 660494
rect 29186 653258 29422 653494
rect 29186 646258 29422 646494
rect 29186 639258 29422 639494
rect 29186 632258 29422 632494
rect 29186 625258 29422 625494
rect 29186 618258 29422 618494
rect 29186 611258 29422 611494
rect 29186 604258 29422 604494
rect 29186 597258 29422 597494
rect 29186 590258 29422 590494
rect 29186 583258 29422 583494
rect 29186 576258 29422 576494
rect 29186 569258 29422 569494
rect 29186 562258 29422 562494
rect 29186 555258 29422 555494
rect 29186 548258 29422 548494
rect 29186 541258 29422 541494
rect 29186 534258 29422 534494
rect 29186 527258 29422 527494
rect 29186 520258 29422 520494
rect 29186 513258 29422 513494
rect 29186 506258 29422 506494
rect 29186 499258 29422 499494
rect 29186 492258 29422 492494
rect 29186 485258 29422 485494
rect 29186 478258 29422 478494
rect 29186 471258 29422 471494
rect 29186 464258 29422 464494
rect 29186 457258 29422 457494
rect 29186 450258 29422 450494
rect 29186 443258 29422 443494
rect 29186 436258 29422 436494
rect 29186 429258 29422 429494
rect 29186 422258 29422 422494
rect 29186 415258 29422 415494
rect 29186 408258 29422 408494
rect 29186 401258 29422 401494
rect 29186 394258 29422 394494
rect 29186 387258 29422 387494
rect 29186 380258 29422 380494
rect 29186 373258 29422 373494
rect 29186 366258 29422 366494
rect 29186 359258 29422 359494
rect 29186 352258 29422 352494
rect 29186 345258 29422 345494
rect 29186 338258 29422 338494
rect 29186 331258 29422 331494
rect 29186 324258 29422 324494
rect 29186 317258 29422 317494
rect 29186 310258 29422 310494
rect 29186 303258 29422 303494
rect 29186 296258 29422 296494
rect 29186 289258 29422 289494
rect 29186 282258 29422 282494
rect 29186 275258 29422 275494
rect 29186 268258 29422 268494
rect 29186 261258 29422 261494
rect 29186 254258 29422 254494
rect 29186 247258 29422 247494
rect 29186 240258 29422 240494
rect 29186 233258 29422 233494
rect 29186 226258 29422 226494
rect 29186 219258 29422 219494
rect 29186 212258 29422 212494
rect 29186 205258 29422 205494
rect 29186 198258 29422 198494
rect 29186 191258 29422 191494
rect 29186 184258 29422 184494
rect 29186 177258 29422 177494
rect 29186 170258 29422 170494
rect 29186 163258 29422 163494
rect 29186 156258 29422 156494
rect 29186 149258 29422 149494
rect 29186 142258 29422 142494
rect 29186 135258 29422 135494
rect 29186 128258 29422 128494
rect 29186 121258 29422 121494
rect 29186 114258 29422 114494
rect 29186 107258 29422 107494
rect 29186 100258 29422 100494
rect 29186 93258 29422 93494
rect 29186 86258 29422 86494
rect 29186 79258 29422 79494
rect 29186 72258 29422 72494
rect 29186 65258 29422 65494
rect 29186 58258 29422 58494
rect 29186 51258 29422 51494
rect 29186 44258 29422 44494
rect 29186 37258 29422 37494
rect 29186 30258 29422 30494
rect 29186 23258 29422 23494
rect 29186 16258 29422 16494
rect 29186 9258 29422 9494
rect 29186 2258 29422 2494
rect 29186 -982 29422 -746
rect 29186 -1302 29422 -1066
rect 30918 705962 31154 706198
rect 30918 705642 31154 705878
rect 30918 696325 31154 696561
rect 30918 689325 31154 689561
rect 30918 682325 31154 682561
rect 30918 675325 31154 675561
rect 30918 668325 31154 668561
rect 30918 661325 31154 661561
rect 30918 654325 31154 654561
rect 30918 647325 31154 647561
rect 30918 640325 31154 640561
rect 30918 633325 31154 633561
rect 30918 626325 31154 626561
rect 30918 619325 31154 619561
rect 30918 612325 31154 612561
rect 30918 605325 31154 605561
rect 30918 598325 31154 598561
rect 30918 591325 31154 591561
rect 30918 584325 31154 584561
rect 30918 577325 31154 577561
rect 30918 570325 31154 570561
rect 30918 563325 31154 563561
rect 30918 556325 31154 556561
rect 30918 549325 31154 549561
rect 30918 542325 31154 542561
rect 30918 535325 31154 535561
rect 30918 528325 31154 528561
rect 30918 521325 31154 521561
rect 30918 514325 31154 514561
rect 30918 507325 31154 507561
rect 30918 500325 31154 500561
rect 30918 493325 31154 493561
rect 30918 486325 31154 486561
rect 30918 479325 31154 479561
rect 30918 472325 31154 472561
rect 30918 465325 31154 465561
rect 30918 458325 31154 458561
rect 30918 451325 31154 451561
rect 30918 444325 31154 444561
rect 30918 437325 31154 437561
rect 30918 430325 31154 430561
rect 30918 423325 31154 423561
rect 30918 416325 31154 416561
rect 30918 409325 31154 409561
rect 30918 402325 31154 402561
rect 30918 395325 31154 395561
rect 30918 388325 31154 388561
rect 30918 381325 31154 381561
rect 30918 374325 31154 374561
rect 30918 367325 31154 367561
rect 30918 360325 31154 360561
rect 30918 353325 31154 353561
rect 30918 346325 31154 346561
rect 30918 339325 31154 339561
rect 30918 332325 31154 332561
rect 30918 325325 31154 325561
rect 30918 318325 31154 318561
rect 30918 311325 31154 311561
rect 30918 304325 31154 304561
rect 30918 297325 31154 297561
rect 30918 290325 31154 290561
rect 30918 283325 31154 283561
rect 30918 276325 31154 276561
rect 30918 269325 31154 269561
rect 30918 262325 31154 262561
rect 30918 255325 31154 255561
rect 30918 248325 31154 248561
rect 30918 241325 31154 241561
rect 30918 234325 31154 234561
rect 30918 227325 31154 227561
rect 30918 220325 31154 220561
rect 30918 213325 31154 213561
rect 30918 206325 31154 206561
rect 30918 199325 31154 199561
rect 30918 192325 31154 192561
rect 30918 185325 31154 185561
rect 30918 178325 31154 178561
rect 30918 171325 31154 171561
rect 30918 164325 31154 164561
rect 30918 157325 31154 157561
rect 30918 150325 31154 150561
rect 30918 143325 31154 143561
rect 30918 136325 31154 136561
rect 30918 129325 31154 129561
rect 30918 122325 31154 122561
rect 30918 115325 31154 115561
rect 30918 108325 31154 108561
rect 30918 101325 31154 101561
rect 30918 94325 31154 94561
rect 30918 87325 31154 87561
rect 30918 80325 31154 80561
rect 30918 73325 31154 73561
rect 30918 66325 31154 66561
rect 30918 59325 31154 59561
rect 30918 52325 31154 52561
rect 30918 45325 31154 45561
rect 30918 38325 31154 38561
rect 30918 31325 31154 31561
rect 30918 24325 31154 24561
rect 30918 17325 31154 17561
rect 30918 10325 31154 10561
rect 30918 3325 31154 3561
rect 30918 -1942 31154 -1706
rect 30918 -2262 31154 -2026
rect 36186 705002 36422 705238
rect 36186 704682 36422 704918
rect 36186 695258 36422 695494
rect 36186 688258 36422 688494
rect 36186 681258 36422 681494
rect 36186 674258 36422 674494
rect 36186 667258 36422 667494
rect 36186 660258 36422 660494
rect 36186 653258 36422 653494
rect 36186 646258 36422 646494
rect 36186 639258 36422 639494
rect 36186 632258 36422 632494
rect 36186 625258 36422 625494
rect 36186 618258 36422 618494
rect 36186 611258 36422 611494
rect 36186 604258 36422 604494
rect 36186 597258 36422 597494
rect 36186 590258 36422 590494
rect 36186 583258 36422 583494
rect 36186 576258 36422 576494
rect 36186 569258 36422 569494
rect 36186 562258 36422 562494
rect 36186 555258 36422 555494
rect 36186 548258 36422 548494
rect 36186 541258 36422 541494
rect 36186 534258 36422 534494
rect 36186 527258 36422 527494
rect 36186 520258 36422 520494
rect 36186 513258 36422 513494
rect 36186 506258 36422 506494
rect 36186 499258 36422 499494
rect 36186 492258 36422 492494
rect 36186 485258 36422 485494
rect 36186 478258 36422 478494
rect 36186 471258 36422 471494
rect 36186 464258 36422 464494
rect 36186 457258 36422 457494
rect 36186 450258 36422 450494
rect 36186 443258 36422 443494
rect 36186 436258 36422 436494
rect 36186 429258 36422 429494
rect 36186 422258 36422 422494
rect 36186 415258 36422 415494
rect 36186 408258 36422 408494
rect 36186 401258 36422 401494
rect 36186 394258 36422 394494
rect 36186 387258 36422 387494
rect 36186 380258 36422 380494
rect 36186 373258 36422 373494
rect 36186 366258 36422 366494
rect 36186 359258 36422 359494
rect 36186 352258 36422 352494
rect 36186 345258 36422 345494
rect 36186 338258 36422 338494
rect 36186 331258 36422 331494
rect 36186 324258 36422 324494
rect 36186 317258 36422 317494
rect 36186 310258 36422 310494
rect 36186 303258 36422 303494
rect 36186 296258 36422 296494
rect 36186 289258 36422 289494
rect 36186 282258 36422 282494
rect 36186 275258 36422 275494
rect 36186 268258 36422 268494
rect 36186 261258 36422 261494
rect 36186 254258 36422 254494
rect 36186 247258 36422 247494
rect 36186 240258 36422 240494
rect 36186 233258 36422 233494
rect 36186 226258 36422 226494
rect 36186 219258 36422 219494
rect 36186 212258 36422 212494
rect 36186 205258 36422 205494
rect 36186 198258 36422 198494
rect 36186 191258 36422 191494
rect 36186 184258 36422 184494
rect 36186 177258 36422 177494
rect 36186 170258 36422 170494
rect 36186 163258 36422 163494
rect 36186 156258 36422 156494
rect 36186 149258 36422 149494
rect 36186 142258 36422 142494
rect 36186 135258 36422 135494
rect 36186 128258 36422 128494
rect 36186 121258 36422 121494
rect 36186 114258 36422 114494
rect 36186 107258 36422 107494
rect 36186 100258 36422 100494
rect 36186 93258 36422 93494
rect 36186 86258 36422 86494
rect 36186 79258 36422 79494
rect 36186 72258 36422 72494
rect 36186 65258 36422 65494
rect 36186 58258 36422 58494
rect 36186 51258 36422 51494
rect 36186 44258 36422 44494
rect 36186 37258 36422 37494
rect 36186 30258 36422 30494
rect 36186 23258 36422 23494
rect 36186 16258 36422 16494
rect 36186 9258 36422 9494
rect 36186 2258 36422 2494
rect 36186 -982 36422 -746
rect 36186 -1302 36422 -1066
rect 37918 705962 38154 706198
rect 37918 705642 38154 705878
rect 37918 696325 38154 696561
rect 37918 689325 38154 689561
rect 37918 682325 38154 682561
rect 37918 675325 38154 675561
rect 37918 668325 38154 668561
rect 37918 661325 38154 661561
rect 37918 654325 38154 654561
rect 37918 647325 38154 647561
rect 37918 640325 38154 640561
rect 37918 633325 38154 633561
rect 37918 626325 38154 626561
rect 37918 619325 38154 619561
rect 37918 612325 38154 612561
rect 37918 605325 38154 605561
rect 37918 598325 38154 598561
rect 37918 591325 38154 591561
rect 37918 584325 38154 584561
rect 37918 577325 38154 577561
rect 37918 570325 38154 570561
rect 37918 563325 38154 563561
rect 37918 556325 38154 556561
rect 37918 549325 38154 549561
rect 37918 542325 38154 542561
rect 37918 535325 38154 535561
rect 37918 528325 38154 528561
rect 37918 521325 38154 521561
rect 37918 514325 38154 514561
rect 37918 507325 38154 507561
rect 37918 500325 38154 500561
rect 37918 493325 38154 493561
rect 37918 486325 38154 486561
rect 37918 479325 38154 479561
rect 37918 472325 38154 472561
rect 37918 465325 38154 465561
rect 37918 458325 38154 458561
rect 37918 451325 38154 451561
rect 37918 444325 38154 444561
rect 37918 437325 38154 437561
rect 37918 430325 38154 430561
rect 37918 423325 38154 423561
rect 37918 416325 38154 416561
rect 37918 409325 38154 409561
rect 37918 402325 38154 402561
rect 37918 395325 38154 395561
rect 37918 388325 38154 388561
rect 37918 381325 38154 381561
rect 37918 374325 38154 374561
rect 37918 367325 38154 367561
rect 37918 360325 38154 360561
rect 37918 353325 38154 353561
rect 37918 346325 38154 346561
rect 37918 339325 38154 339561
rect 37918 332325 38154 332561
rect 37918 325325 38154 325561
rect 37918 318325 38154 318561
rect 37918 311325 38154 311561
rect 37918 304325 38154 304561
rect 37918 297325 38154 297561
rect 37918 290325 38154 290561
rect 37918 283325 38154 283561
rect 37918 276325 38154 276561
rect 37918 269325 38154 269561
rect 37918 262325 38154 262561
rect 37918 255325 38154 255561
rect 37918 248325 38154 248561
rect 37918 241325 38154 241561
rect 37918 234325 38154 234561
rect 37918 227325 38154 227561
rect 37918 220325 38154 220561
rect 37918 213325 38154 213561
rect 37918 206325 38154 206561
rect 37918 199325 38154 199561
rect 37918 192325 38154 192561
rect 37918 185325 38154 185561
rect 37918 178325 38154 178561
rect 37918 171325 38154 171561
rect 37918 164325 38154 164561
rect 37918 157325 38154 157561
rect 37918 150325 38154 150561
rect 37918 143325 38154 143561
rect 37918 136325 38154 136561
rect 37918 129325 38154 129561
rect 37918 122325 38154 122561
rect 37918 115325 38154 115561
rect 37918 108325 38154 108561
rect 37918 101325 38154 101561
rect 37918 94325 38154 94561
rect 37918 87325 38154 87561
rect 37918 80325 38154 80561
rect 37918 73325 38154 73561
rect 37918 66325 38154 66561
rect 37918 59325 38154 59561
rect 37918 52325 38154 52561
rect 37918 45325 38154 45561
rect 37918 38325 38154 38561
rect 37918 31325 38154 31561
rect 37918 24325 38154 24561
rect 37918 17325 38154 17561
rect 37918 10325 38154 10561
rect 37918 3325 38154 3561
rect 37918 -1942 38154 -1706
rect 37918 -2262 38154 -2026
rect 43186 705002 43422 705238
rect 43186 704682 43422 704918
rect 43186 695258 43422 695494
rect 43186 688258 43422 688494
rect 43186 681258 43422 681494
rect 43186 674258 43422 674494
rect 43186 667258 43422 667494
rect 43186 660258 43422 660494
rect 43186 653258 43422 653494
rect 43186 646258 43422 646494
rect 43186 639258 43422 639494
rect 43186 632258 43422 632494
rect 43186 625258 43422 625494
rect 43186 618258 43422 618494
rect 43186 611258 43422 611494
rect 43186 604258 43422 604494
rect 43186 597258 43422 597494
rect 43186 590258 43422 590494
rect 43186 583258 43422 583494
rect 43186 576258 43422 576494
rect 43186 569258 43422 569494
rect 43186 562258 43422 562494
rect 43186 555258 43422 555494
rect 43186 548258 43422 548494
rect 43186 541258 43422 541494
rect 43186 534258 43422 534494
rect 43186 527258 43422 527494
rect 43186 520258 43422 520494
rect 43186 513258 43422 513494
rect 43186 506258 43422 506494
rect 43186 499258 43422 499494
rect 43186 492258 43422 492494
rect 43186 485258 43422 485494
rect 43186 478258 43422 478494
rect 43186 471258 43422 471494
rect 43186 464258 43422 464494
rect 43186 457258 43422 457494
rect 43186 450258 43422 450494
rect 43186 443258 43422 443494
rect 43186 436258 43422 436494
rect 43186 429258 43422 429494
rect 43186 422258 43422 422494
rect 43186 415258 43422 415494
rect 43186 408258 43422 408494
rect 43186 401258 43422 401494
rect 43186 394258 43422 394494
rect 43186 387258 43422 387494
rect 43186 380258 43422 380494
rect 43186 373258 43422 373494
rect 43186 366258 43422 366494
rect 43186 359258 43422 359494
rect 43186 352258 43422 352494
rect 43186 345258 43422 345494
rect 43186 338258 43422 338494
rect 43186 331258 43422 331494
rect 43186 324258 43422 324494
rect 43186 317258 43422 317494
rect 43186 310258 43422 310494
rect 43186 303258 43422 303494
rect 43186 296258 43422 296494
rect 43186 289258 43422 289494
rect 43186 282258 43422 282494
rect 43186 275258 43422 275494
rect 43186 268258 43422 268494
rect 43186 261258 43422 261494
rect 43186 254258 43422 254494
rect 43186 247258 43422 247494
rect 43186 240258 43422 240494
rect 43186 233258 43422 233494
rect 43186 226258 43422 226494
rect 43186 219258 43422 219494
rect 43186 212258 43422 212494
rect 43186 205258 43422 205494
rect 43186 198258 43422 198494
rect 43186 191258 43422 191494
rect 43186 184258 43422 184494
rect 43186 177258 43422 177494
rect 43186 170258 43422 170494
rect 43186 163258 43422 163494
rect 43186 156258 43422 156494
rect 43186 149258 43422 149494
rect 43186 142258 43422 142494
rect 43186 135258 43422 135494
rect 43186 128258 43422 128494
rect 43186 121258 43422 121494
rect 43186 114258 43422 114494
rect 43186 107258 43422 107494
rect 43186 100258 43422 100494
rect 43186 93258 43422 93494
rect 43186 86258 43422 86494
rect 43186 79258 43422 79494
rect 43186 72258 43422 72494
rect 43186 65258 43422 65494
rect 43186 58258 43422 58494
rect 43186 51258 43422 51494
rect 43186 44258 43422 44494
rect 43186 37258 43422 37494
rect 43186 30258 43422 30494
rect 43186 23258 43422 23494
rect 43186 16258 43422 16494
rect 43186 9258 43422 9494
rect 43186 2258 43422 2494
rect 43186 -982 43422 -746
rect 43186 -1302 43422 -1066
rect 44918 705962 45154 706198
rect 44918 705642 45154 705878
rect 44918 696325 45154 696561
rect 44918 689325 45154 689561
rect 44918 682325 45154 682561
rect 44918 675325 45154 675561
rect 44918 668325 45154 668561
rect 44918 661325 45154 661561
rect 44918 654325 45154 654561
rect 44918 647325 45154 647561
rect 44918 640325 45154 640561
rect 44918 633325 45154 633561
rect 44918 626325 45154 626561
rect 44918 619325 45154 619561
rect 44918 612325 45154 612561
rect 44918 605325 45154 605561
rect 44918 598325 45154 598561
rect 44918 591325 45154 591561
rect 44918 584325 45154 584561
rect 44918 577325 45154 577561
rect 44918 570325 45154 570561
rect 44918 563325 45154 563561
rect 44918 556325 45154 556561
rect 44918 549325 45154 549561
rect 44918 542325 45154 542561
rect 44918 535325 45154 535561
rect 44918 528325 45154 528561
rect 44918 521325 45154 521561
rect 44918 514325 45154 514561
rect 44918 507325 45154 507561
rect 44918 500325 45154 500561
rect 44918 493325 45154 493561
rect 44918 486325 45154 486561
rect 44918 479325 45154 479561
rect 44918 472325 45154 472561
rect 44918 465325 45154 465561
rect 44918 458325 45154 458561
rect 44918 451325 45154 451561
rect 44918 444325 45154 444561
rect 44918 437325 45154 437561
rect 44918 430325 45154 430561
rect 44918 423325 45154 423561
rect 44918 416325 45154 416561
rect 44918 409325 45154 409561
rect 44918 402325 45154 402561
rect 44918 395325 45154 395561
rect 44918 388325 45154 388561
rect 44918 381325 45154 381561
rect 44918 374325 45154 374561
rect 44918 367325 45154 367561
rect 44918 360325 45154 360561
rect 44918 353325 45154 353561
rect 44918 346325 45154 346561
rect 44918 339325 45154 339561
rect 44918 332325 45154 332561
rect 44918 325325 45154 325561
rect 44918 318325 45154 318561
rect 44918 311325 45154 311561
rect 44918 304325 45154 304561
rect 44918 297325 45154 297561
rect 44918 290325 45154 290561
rect 44918 283325 45154 283561
rect 44918 276325 45154 276561
rect 44918 269325 45154 269561
rect 44918 262325 45154 262561
rect 44918 255325 45154 255561
rect 44918 248325 45154 248561
rect 44918 241325 45154 241561
rect 44918 234325 45154 234561
rect 44918 227325 45154 227561
rect 44918 220325 45154 220561
rect 44918 213325 45154 213561
rect 44918 206325 45154 206561
rect 44918 199325 45154 199561
rect 44918 192325 45154 192561
rect 44918 185325 45154 185561
rect 44918 178325 45154 178561
rect 44918 171325 45154 171561
rect 44918 164325 45154 164561
rect 44918 157325 45154 157561
rect 44918 150325 45154 150561
rect 44918 143325 45154 143561
rect 44918 136325 45154 136561
rect 44918 129325 45154 129561
rect 44918 122325 45154 122561
rect 44918 115325 45154 115561
rect 44918 108325 45154 108561
rect 44918 101325 45154 101561
rect 44918 94325 45154 94561
rect 44918 87325 45154 87561
rect 44918 80325 45154 80561
rect 44918 73325 45154 73561
rect 44918 66325 45154 66561
rect 44918 59325 45154 59561
rect 44918 52325 45154 52561
rect 44918 45325 45154 45561
rect 44918 38325 45154 38561
rect 44918 31325 45154 31561
rect 44918 24325 45154 24561
rect 44918 17325 45154 17561
rect 44918 10325 45154 10561
rect 44918 3325 45154 3561
rect 44918 -1942 45154 -1706
rect 44918 -2262 45154 -2026
rect 50186 705002 50422 705238
rect 50186 704682 50422 704918
rect 50186 695258 50422 695494
rect 50186 688258 50422 688494
rect 50186 681258 50422 681494
rect 50186 674258 50422 674494
rect 50186 667258 50422 667494
rect 50186 660258 50422 660494
rect 50186 653258 50422 653494
rect 50186 646258 50422 646494
rect 50186 639258 50422 639494
rect 50186 632258 50422 632494
rect 50186 625258 50422 625494
rect 50186 618258 50422 618494
rect 50186 611258 50422 611494
rect 50186 604258 50422 604494
rect 50186 597258 50422 597494
rect 50186 590258 50422 590494
rect 50186 583258 50422 583494
rect 50186 576258 50422 576494
rect 50186 569258 50422 569494
rect 50186 562258 50422 562494
rect 50186 555258 50422 555494
rect 50186 548258 50422 548494
rect 50186 541258 50422 541494
rect 50186 534258 50422 534494
rect 50186 527258 50422 527494
rect 50186 520258 50422 520494
rect 50186 513258 50422 513494
rect 50186 506258 50422 506494
rect 50186 499258 50422 499494
rect 50186 492258 50422 492494
rect 50186 485258 50422 485494
rect 50186 478258 50422 478494
rect 50186 471258 50422 471494
rect 50186 464258 50422 464494
rect 50186 457258 50422 457494
rect 50186 450258 50422 450494
rect 50186 443258 50422 443494
rect 50186 436258 50422 436494
rect 50186 429258 50422 429494
rect 50186 422258 50422 422494
rect 50186 415258 50422 415494
rect 50186 408258 50422 408494
rect 50186 401258 50422 401494
rect 50186 394258 50422 394494
rect 50186 387258 50422 387494
rect 50186 380258 50422 380494
rect 50186 373258 50422 373494
rect 50186 366258 50422 366494
rect 50186 359258 50422 359494
rect 50186 352258 50422 352494
rect 50186 345258 50422 345494
rect 50186 338258 50422 338494
rect 50186 331258 50422 331494
rect 50186 324258 50422 324494
rect 50186 317258 50422 317494
rect 50186 310258 50422 310494
rect 50186 303258 50422 303494
rect 50186 296258 50422 296494
rect 50186 289258 50422 289494
rect 50186 282258 50422 282494
rect 50186 275258 50422 275494
rect 50186 268258 50422 268494
rect 50186 261258 50422 261494
rect 50186 254258 50422 254494
rect 50186 247258 50422 247494
rect 50186 240258 50422 240494
rect 50186 233258 50422 233494
rect 50186 226258 50422 226494
rect 50186 219258 50422 219494
rect 50186 212258 50422 212494
rect 50186 205258 50422 205494
rect 50186 198258 50422 198494
rect 50186 191258 50422 191494
rect 50186 184258 50422 184494
rect 50186 177258 50422 177494
rect 50186 170258 50422 170494
rect 50186 163258 50422 163494
rect 50186 156258 50422 156494
rect 50186 149258 50422 149494
rect 50186 142258 50422 142494
rect 50186 135258 50422 135494
rect 50186 128258 50422 128494
rect 50186 121258 50422 121494
rect 50186 114258 50422 114494
rect 50186 107258 50422 107494
rect 50186 100258 50422 100494
rect 50186 93258 50422 93494
rect 50186 86258 50422 86494
rect 50186 79258 50422 79494
rect 50186 72258 50422 72494
rect 50186 65258 50422 65494
rect 50186 58258 50422 58494
rect 50186 51258 50422 51494
rect 50186 44258 50422 44494
rect 50186 37258 50422 37494
rect 50186 30258 50422 30494
rect 50186 23258 50422 23494
rect 50186 16258 50422 16494
rect 50186 9258 50422 9494
rect 50186 2258 50422 2494
rect 50186 -982 50422 -746
rect 50186 -1302 50422 -1066
rect 51918 705962 52154 706198
rect 51918 705642 52154 705878
rect 51918 696325 52154 696561
rect 51918 689325 52154 689561
rect 51918 682325 52154 682561
rect 51918 675325 52154 675561
rect 51918 668325 52154 668561
rect 51918 661325 52154 661561
rect 51918 654325 52154 654561
rect 51918 647325 52154 647561
rect 51918 640325 52154 640561
rect 51918 633325 52154 633561
rect 51918 626325 52154 626561
rect 51918 619325 52154 619561
rect 51918 612325 52154 612561
rect 51918 605325 52154 605561
rect 51918 598325 52154 598561
rect 51918 591325 52154 591561
rect 51918 584325 52154 584561
rect 51918 577325 52154 577561
rect 51918 570325 52154 570561
rect 51918 563325 52154 563561
rect 51918 556325 52154 556561
rect 51918 549325 52154 549561
rect 51918 542325 52154 542561
rect 51918 535325 52154 535561
rect 51918 528325 52154 528561
rect 51918 521325 52154 521561
rect 51918 514325 52154 514561
rect 51918 507325 52154 507561
rect 51918 500325 52154 500561
rect 51918 493325 52154 493561
rect 51918 486325 52154 486561
rect 51918 479325 52154 479561
rect 51918 472325 52154 472561
rect 51918 465325 52154 465561
rect 51918 458325 52154 458561
rect 51918 451325 52154 451561
rect 51918 444325 52154 444561
rect 51918 437325 52154 437561
rect 51918 430325 52154 430561
rect 51918 423325 52154 423561
rect 51918 416325 52154 416561
rect 51918 409325 52154 409561
rect 51918 402325 52154 402561
rect 51918 395325 52154 395561
rect 51918 388325 52154 388561
rect 51918 381325 52154 381561
rect 51918 374325 52154 374561
rect 51918 367325 52154 367561
rect 51918 360325 52154 360561
rect 51918 353325 52154 353561
rect 51918 346325 52154 346561
rect 51918 339325 52154 339561
rect 51918 332325 52154 332561
rect 51918 325325 52154 325561
rect 51918 318325 52154 318561
rect 51918 311325 52154 311561
rect 51918 304325 52154 304561
rect 51918 297325 52154 297561
rect 51918 290325 52154 290561
rect 51918 283325 52154 283561
rect 51918 276325 52154 276561
rect 51918 269325 52154 269561
rect 51918 262325 52154 262561
rect 51918 255325 52154 255561
rect 51918 248325 52154 248561
rect 51918 241325 52154 241561
rect 51918 234325 52154 234561
rect 51918 227325 52154 227561
rect 51918 220325 52154 220561
rect 51918 213325 52154 213561
rect 51918 206325 52154 206561
rect 51918 199325 52154 199561
rect 51918 192325 52154 192561
rect 51918 185325 52154 185561
rect 51918 178325 52154 178561
rect 51918 171325 52154 171561
rect 51918 164325 52154 164561
rect 51918 157325 52154 157561
rect 51918 150325 52154 150561
rect 51918 143325 52154 143561
rect 51918 136325 52154 136561
rect 51918 129325 52154 129561
rect 51918 122325 52154 122561
rect 51918 115325 52154 115561
rect 51918 108325 52154 108561
rect 51918 101325 52154 101561
rect 51918 94325 52154 94561
rect 51918 87325 52154 87561
rect 51918 80325 52154 80561
rect 51918 73325 52154 73561
rect 51918 66325 52154 66561
rect 51918 59325 52154 59561
rect 51918 52325 52154 52561
rect 51918 45325 52154 45561
rect 51918 38325 52154 38561
rect 51918 31325 52154 31561
rect 51918 24325 52154 24561
rect 51918 17325 52154 17561
rect 51918 10325 52154 10561
rect 51918 3325 52154 3561
rect 51918 -1942 52154 -1706
rect 51918 -2262 52154 -2026
rect 57186 705002 57422 705238
rect 57186 704682 57422 704918
rect 57186 695258 57422 695494
rect 57186 688258 57422 688494
rect 57186 681258 57422 681494
rect 57186 674258 57422 674494
rect 57186 667258 57422 667494
rect 57186 660258 57422 660494
rect 57186 653258 57422 653494
rect 57186 646258 57422 646494
rect 57186 639258 57422 639494
rect 57186 632258 57422 632494
rect 57186 625258 57422 625494
rect 57186 618258 57422 618494
rect 57186 611258 57422 611494
rect 57186 604258 57422 604494
rect 57186 597258 57422 597494
rect 57186 590258 57422 590494
rect 57186 583258 57422 583494
rect 57186 576258 57422 576494
rect 57186 569258 57422 569494
rect 57186 562258 57422 562494
rect 57186 555258 57422 555494
rect 57186 548258 57422 548494
rect 57186 541258 57422 541494
rect 57186 534258 57422 534494
rect 57186 527258 57422 527494
rect 57186 520258 57422 520494
rect 57186 513258 57422 513494
rect 57186 506258 57422 506494
rect 57186 499258 57422 499494
rect 57186 492258 57422 492494
rect 57186 485258 57422 485494
rect 57186 478258 57422 478494
rect 57186 471258 57422 471494
rect 57186 464258 57422 464494
rect 57186 457258 57422 457494
rect 57186 450258 57422 450494
rect 57186 443258 57422 443494
rect 57186 436258 57422 436494
rect 57186 429258 57422 429494
rect 57186 422258 57422 422494
rect 57186 415258 57422 415494
rect 57186 408258 57422 408494
rect 57186 401258 57422 401494
rect 57186 394258 57422 394494
rect 57186 387258 57422 387494
rect 57186 380258 57422 380494
rect 57186 373258 57422 373494
rect 57186 366258 57422 366494
rect 57186 359258 57422 359494
rect 57186 352258 57422 352494
rect 57186 345258 57422 345494
rect 57186 338258 57422 338494
rect 57186 331258 57422 331494
rect 57186 324258 57422 324494
rect 57186 317258 57422 317494
rect 57186 310258 57422 310494
rect 57186 303258 57422 303494
rect 57186 296258 57422 296494
rect 57186 289258 57422 289494
rect 57186 282258 57422 282494
rect 57186 275258 57422 275494
rect 57186 268258 57422 268494
rect 57186 261258 57422 261494
rect 57186 254258 57422 254494
rect 57186 247258 57422 247494
rect 57186 240258 57422 240494
rect 57186 233258 57422 233494
rect 57186 226258 57422 226494
rect 57186 219258 57422 219494
rect 57186 212258 57422 212494
rect 57186 205258 57422 205494
rect 57186 198258 57422 198494
rect 57186 191258 57422 191494
rect 57186 184258 57422 184494
rect 57186 177258 57422 177494
rect 57186 170258 57422 170494
rect 57186 163258 57422 163494
rect 57186 156258 57422 156494
rect 57186 149258 57422 149494
rect 57186 142258 57422 142494
rect 57186 135258 57422 135494
rect 57186 128258 57422 128494
rect 57186 121258 57422 121494
rect 57186 114258 57422 114494
rect 57186 107258 57422 107494
rect 57186 100258 57422 100494
rect 57186 93258 57422 93494
rect 57186 86258 57422 86494
rect 57186 79258 57422 79494
rect 57186 72258 57422 72494
rect 57186 65258 57422 65494
rect 57186 58258 57422 58494
rect 57186 51258 57422 51494
rect 57186 44258 57422 44494
rect 57186 37258 57422 37494
rect 57186 30258 57422 30494
rect 57186 23258 57422 23494
rect 57186 16258 57422 16494
rect 57186 9258 57422 9494
rect 57186 2258 57422 2494
rect 57186 -982 57422 -746
rect 57186 -1302 57422 -1066
rect 58918 705962 59154 706198
rect 58918 705642 59154 705878
rect 58918 696325 59154 696561
rect 58918 689325 59154 689561
rect 58918 682325 59154 682561
rect 58918 675325 59154 675561
rect 58918 668325 59154 668561
rect 58918 661325 59154 661561
rect 58918 654325 59154 654561
rect 58918 647325 59154 647561
rect 58918 640325 59154 640561
rect 58918 633325 59154 633561
rect 58918 626325 59154 626561
rect 58918 619325 59154 619561
rect 58918 612325 59154 612561
rect 58918 605325 59154 605561
rect 58918 598325 59154 598561
rect 58918 591325 59154 591561
rect 58918 584325 59154 584561
rect 58918 577325 59154 577561
rect 58918 570325 59154 570561
rect 58918 563325 59154 563561
rect 58918 556325 59154 556561
rect 58918 549325 59154 549561
rect 58918 542325 59154 542561
rect 58918 535325 59154 535561
rect 58918 528325 59154 528561
rect 58918 521325 59154 521561
rect 58918 514325 59154 514561
rect 58918 507325 59154 507561
rect 58918 500325 59154 500561
rect 58918 493325 59154 493561
rect 58918 486325 59154 486561
rect 58918 479325 59154 479561
rect 58918 472325 59154 472561
rect 58918 465325 59154 465561
rect 58918 458325 59154 458561
rect 58918 451325 59154 451561
rect 58918 444325 59154 444561
rect 58918 437325 59154 437561
rect 58918 430325 59154 430561
rect 58918 423325 59154 423561
rect 58918 416325 59154 416561
rect 58918 409325 59154 409561
rect 58918 402325 59154 402561
rect 58918 395325 59154 395561
rect 58918 388325 59154 388561
rect 58918 381325 59154 381561
rect 58918 374325 59154 374561
rect 58918 367325 59154 367561
rect 58918 360325 59154 360561
rect 58918 353325 59154 353561
rect 58918 346325 59154 346561
rect 58918 339325 59154 339561
rect 58918 332325 59154 332561
rect 58918 325325 59154 325561
rect 58918 318325 59154 318561
rect 58918 311325 59154 311561
rect 58918 304325 59154 304561
rect 58918 297325 59154 297561
rect 58918 290325 59154 290561
rect 58918 283325 59154 283561
rect 58918 276325 59154 276561
rect 58918 269325 59154 269561
rect 58918 262325 59154 262561
rect 58918 255325 59154 255561
rect 58918 248325 59154 248561
rect 58918 241325 59154 241561
rect 58918 234325 59154 234561
rect 58918 227325 59154 227561
rect 58918 220325 59154 220561
rect 58918 213325 59154 213561
rect 58918 206325 59154 206561
rect 58918 199325 59154 199561
rect 58918 192325 59154 192561
rect 58918 185325 59154 185561
rect 58918 178325 59154 178561
rect 58918 171325 59154 171561
rect 58918 164325 59154 164561
rect 58918 157325 59154 157561
rect 58918 150325 59154 150561
rect 58918 143325 59154 143561
rect 58918 136325 59154 136561
rect 58918 129325 59154 129561
rect 58918 122325 59154 122561
rect 58918 115325 59154 115561
rect 58918 108325 59154 108561
rect 58918 101325 59154 101561
rect 58918 94325 59154 94561
rect 58918 87325 59154 87561
rect 58918 80325 59154 80561
rect 58918 73325 59154 73561
rect 58918 66325 59154 66561
rect 58918 59325 59154 59561
rect 58918 52325 59154 52561
rect 58918 45325 59154 45561
rect 58918 38325 59154 38561
rect 58918 31325 59154 31561
rect 58918 24325 59154 24561
rect 58918 17325 59154 17561
rect 58918 10325 59154 10561
rect 58918 3325 59154 3561
rect 58918 -1942 59154 -1706
rect 58918 -2262 59154 -2026
rect 64186 705002 64422 705238
rect 64186 704682 64422 704918
rect 64186 695258 64422 695494
rect 64186 688258 64422 688494
rect 64186 681258 64422 681494
rect 64186 674258 64422 674494
rect 64186 667258 64422 667494
rect 64186 660258 64422 660494
rect 64186 653258 64422 653494
rect 64186 646258 64422 646494
rect 64186 639258 64422 639494
rect 64186 632258 64422 632494
rect 64186 625258 64422 625494
rect 64186 618258 64422 618494
rect 64186 611258 64422 611494
rect 64186 604258 64422 604494
rect 64186 597258 64422 597494
rect 64186 590258 64422 590494
rect 64186 583258 64422 583494
rect 64186 576258 64422 576494
rect 64186 569258 64422 569494
rect 64186 562258 64422 562494
rect 64186 555258 64422 555494
rect 64186 548258 64422 548494
rect 64186 541258 64422 541494
rect 64186 534258 64422 534494
rect 64186 527258 64422 527494
rect 64186 520258 64422 520494
rect 64186 513258 64422 513494
rect 64186 506258 64422 506494
rect 64186 499258 64422 499494
rect 64186 492258 64422 492494
rect 64186 485258 64422 485494
rect 64186 478258 64422 478494
rect 64186 471258 64422 471494
rect 64186 464258 64422 464494
rect 64186 457258 64422 457494
rect 64186 450258 64422 450494
rect 64186 443258 64422 443494
rect 64186 436258 64422 436494
rect 64186 429258 64422 429494
rect 64186 422258 64422 422494
rect 64186 415258 64422 415494
rect 64186 408258 64422 408494
rect 64186 401258 64422 401494
rect 64186 394258 64422 394494
rect 64186 387258 64422 387494
rect 64186 380258 64422 380494
rect 64186 373258 64422 373494
rect 64186 366258 64422 366494
rect 64186 359258 64422 359494
rect 64186 352258 64422 352494
rect 64186 345258 64422 345494
rect 64186 338258 64422 338494
rect 64186 331258 64422 331494
rect 64186 324258 64422 324494
rect 64186 317258 64422 317494
rect 64186 310258 64422 310494
rect 64186 303258 64422 303494
rect 64186 296258 64422 296494
rect 64186 289258 64422 289494
rect 64186 282258 64422 282494
rect 64186 275258 64422 275494
rect 64186 268258 64422 268494
rect 64186 261258 64422 261494
rect 64186 254258 64422 254494
rect 64186 247258 64422 247494
rect 64186 240258 64422 240494
rect 64186 233258 64422 233494
rect 64186 226258 64422 226494
rect 64186 219258 64422 219494
rect 64186 212258 64422 212494
rect 64186 205258 64422 205494
rect 64186 198258 64422 198494
rect 64186 191258 64422 191494
rect 64186 184258 64422 184494
rect 64186 177258 64422 177494
rect 64186 170258 64422 170494
rect 64186 163258 64422 163494
rect 64186 156258 64422 156494
rect 64186 149258 64422 149494
rect 64186 142258 64422 142494
rect 64186 135258 64422 135494
rect 64186 128258 64422 128494
rect 64186 121258 64422 121494
rect 64186 114258 64422 114494
rect 64186 107258 64422 107494
rect 64186 100258 64422 100494
rect 64186 93258 64422 93494
rect 64186 86258 64422 86494
rect 64186 79258 64422 79494
rect 64186 72258 64422 72494
rect 64186 65258 64422 65494
rect 64186 58258 64422 58494
rect 64186 51258 64422 51494
rect 64186 44258 64422 44494
rect 64186 37258 64422 37494
rect 64186 30258 64422 30494
rect 64186 23258 64422 23494
rect 64186 16258 64422 16494
rect 64186 9258 64422 9494
rect 64186 2258 64422 2494
rect 64186 -982 64422 -746
rect 64186 -1302 64422 -1066
rect 65918 705962 66154 706198
rect 65918 705642 66154 705878
rect 65918 696325 66154 696561
rect 65918 689325 66154 689561
rect 65918 682325 66154 682561
rect 65918 675325 66154 675561
rect 65918 668325 66154 668561
rect 65918 661325 66154 661561
rect 65918 654325 66154 654561
rect 65918 647325 66154 647561
rect 65918 640325 66154 640561
rect 65918 633325 66154 633561
rect 65918 626325 66154 626561
rect 65918 619325 66154 619561
rect 65918 612325 66154 612561
rect 65918 605325 66154 605561
rect 65918 598325 66154 598561
rect 65918 591325 66154 591561
rect 65918 584325 66154 584561
rect 65918 577325 66154 577561
rect 65918 570325 66154 570561
rect 65918 563325 66154 563561
rect 65918 556325 66154 556561
rect 65918 549325 66154 549561
rect 65918 542325 66154 542561
rect 65918 535325 66154 535561
rect 65918 528325 66154 528561
rect 65918 521325 66154 521561
rect 65918 514325 66154 514561
rect 65918 507325 66154 507561
rect 65918 500325 66154 500561
rect 65918 493325 66154 493561
rect 65918 486325 66154 486561
rect 65918 479325 66154 479561
rect 65918 472325 66154 472561
rect 65918 465325 66154 465561
rect 65918 458325 66154 458561
rect 65918 451325 66154 451561
rect 65918 444325 66154 444561
rect 65918 437325 66154 437561
rect 65918 430325 66154 430561
rect 65918 423325 66154 423561
rect 65918 416325 66154 416561
rect 65918 409325 66154 409561
rect 65918 402325 66154 402561
rect 65918 395325 66154 395561
rect 65918 388325 66154 388561
rect 65918 381325 66154 381561
rect 65918 374325 66154 374561
rect 65918 367325 66154 367561
rect 65918 360325 66154 360561
rect 65918 353325 66154 353561
rect 65918 346325 66154 346561
rect 65918 339325 66154 339561
rect 65918 332325 66154 332561
rect 65918 325325 66154 325561
rect 65918 318325 66154 318561
rect 65918 311325 66154 311561
rect 65918 304325 66154 304561
rect 65918 297325 66154 297561
rect 65918 290325 66154 290561
rect 65918 283325 66154 283561
rect 65918 276325 66154 276561
rect 65918 269325 66154 269561
rect 65918 262325 66154 262561
rect 65918 255325 66154 255561
rect 65918 248325 66154 248561
rect 65918 241325 66154 241561
rect 65918 234325 66154 234561
rect 65918 227325 66154 227561
rect 65918 220325 66154 220561
rect 65918 213325 66154 213561
rect 65918 206325 66154 206561
rect 65918 199325 66154 199561
rect 65918 192325 66154 192561
rect 65918 185325 66154 185561
rect 65918 178325 66154 178561
rect 65918 171325 66154 171561
rect 65918 164325 66154 164561
rect 65918 157325 66154 157561
rect 65918 150325 66154 150561
rect 65918 143325 66154 143561
rect 65918 136325 66154 136561
rect 65918 129325 66154 129561
rect 65918 122325 66154 122561
rect 65918 115325 66154 115561
rect 65918 108325 66154 108561
rect 65918 101325 66154 101561
rect 65918 94325 66154 94561
rect 65918 87325 66154 87561
rect 65918 80325 66154 80561
rect 65918 73325 66154 73561
rect 65918 66325 66154 66561
rect 65918 59325 66154 59561
rect 65918 52325 66154 52561
rect 65918 45325 66154 45561
rect 65918 38325 66154 38561
rect 65918 31325 66154 31561
rect 65918 24325 66154 24561
rect 65918 17325 66154 17561
rect 65918 10325 66154 10561
rect 65918 3325 66154 3561
rect 65918 -1942 66154 -1706
rect 65918 -2262 66154 -2026
rect 71186 705002 71422 705238
rect 71186 704682 71422 704918
rect 71186 695258 71422 695494
rect 71186 688258 71422 688494
rect 71186 681258 71422 681494
rect 71186 674258 71422 674494
rect 71186 667258 71422 667494
rect 71186 660258 71422 660494
rect 71186 653258 71422 653494
rect 71186 646258 71422 646494
rect 71186 639258 71422 639494
rect 71186 632258 71422 632494
rect 71186 625258 71422 625494
rect 71186 618258 71422 618494
rect 71186 611258 71422 611494
rect 71186 604258 71422 604494
rect 71186 597258 71422 597494
rect 71186 590258 71422 590494
rect 71186 583258 71422 583494
rect 71186 576258 71422 576494
rect 71186 569258 71422 569494
rect 71186 562258 71422 562494
rect 71186 555258 71422 555494
rect 71186 548258 71422 548494
rect 71186 541258 71422 541494
rect 71186 534258 71422 534494
rect 71186 527258 71422 527494
rect 71186 520258 71422 520494
rect 71186 513258 71422 513494
rect 71186 506258 71422 506494
rect 71186 499258 71422 499494
rect 71186 492258 71422 492494
rect 71186 485258 71422 485494
rect 71186 478258 71422 478494
rect 71186 471258 71422 471494
rect 71186 464258 71422 464494
rect 71186 457258 71422 457494
rect 71186 450258 71422 450494
rect 71186 443258 71422 443494
rect 71186 436258 71422 436494
rect 71186 429258 71422 429494
rect 71186 422258 71422 422494
rect 71186 415258 71422 415494
rect 71186 408258 71422 408494
rect 71186 401258 71422 401494
rect 71186 394258 71422 394494
rect 71186 387258 71422 387494
rect 71186 380258 71422 380494
rect 71186 373258 71422 373494
rect 71186 366258 71422 366494
rect 71186 359258 71422 359494
rect 71186 352258 71422 352494
rect 71186 345258 71422 345494
rect 71186 338258 71422 338494
rect 71186 331258 71422 331494
rect 71186 324258 71422 324494
rect 71186 317258 71422 317494
rect 71186 310258 71422 310494
rect 71186 303258 71422 303494
rect 71186 296258 71422 296494
rect 71186 289258 71422 289494
rect 71186 282258 71422 282494
rect 71186 275258 71422 275494
rect 71186 268258 71422 268494
rect 71186 261258 71422 261494
rect 71186 254258 71422 254494
rect 71186 247258 71422 247494
rect 71186 240258 71422 240494
rect 71186 233258 71422 233494
rect 71186 226258 71422 226494
rect 71186 219258 71422 219494
rect 71186 212258 71422 212494
rect 71186 205258 71422 205494
rect 71186 198258 71422 198494
rect 71186 191258 71422 191494
rect 71186 184258 71422 184494
rect 71186 177258 71422 177494
rect 71186 170258 71422 170494
rect 71186 163258 71422 163494
rect 71186 156258 71422 156494
rect 71186 149258 71422 149494
rect 71186 142258 71422 142494
rect 71186 135258 71422 135494
rect 71186 128258 71422 128494
rect 71186 121258 71422 121494
rect 71186 114258 71422 114494
rect 71186 107258 71422 107494
rect 71186 100258 71422 100494
rect 71186 93258 71422 93494
rect 71186 86258 71422 86494
rect 71186 79258 71422 79494
rect 71186 72258 71422 72494
rect 71186 65258 71422 65494
rect 71186 58258 71422 58494
rect 71186 51258 71422 51494
rect 71186 44258 71422 44494
rect 71186 37258 71422 37494
rect 71186 30258 71422 30494
rect 71186 23258 71422 23494
rect 71186 16258 71422 16494
rect 71186 9258 71422 9494
rect 71186 2258 71422 2494
rect 71186 -982 71422 -746
rect 71186 -1302 71422 -1066
rect 72918 705962 73154 706198
rect 72918 705642 73154 705878
rect 72918 696325 73154 696561
rect 72918 689325 73154 689561
rect 72918 682325 73154 682561
rect 72918 675325 73154 675561
rect 72918 668325 73154 668561
rect 72918 661325 73154 661561
rect 72918 654325 73154 654561
rect 72918 647325 73154 647561
rect 72918 640325 73154 640561
rect 72918 633325 73154 633561
rect 72918 626325 73154 626561
rect 72918 619325 73154 619561
rect 72918 612325 73154 612561
rect 72918 605325 73154 605561
rect 72918 598325 73154 598561
rect 72918 591325 73154 591561
rect 72918 584325 73154 584561
rect 72918 577325 73154 577561
rect 72918 570325 73154 570561
rect 72918 563325 73154 563561
rect 72918 556325 73154 556561
rect 72918 549325 73154 549561
rect 72918 542325 73154 542561
rect 72918 535325 73154 535561
rect 72918 528325 73154 528561
rect 72918 521325 73154 521561
rect 72918 514325 73154 514561
rect 72918 507325 73154 507561
rect 72918 500325 73154 500561
rect 72918 493325 73154 493561
rect 72918 486325 73154 486561
rect 72918 479325 73154 479561
rect 72918 472325 73154 472561
rect 72918 465325 73154 465561
rect 72918 458325 73154 458561
rect 72918 451325 73154 451561
rect 72918 444325 73154 444561
rect 72918 437325 73154 437561
rect 72918 430325 73154 430561
rect 72918 423325 73154 423561
rect 72918 416325 73154 416561
rect 72918 409325 73154 409561
rect 72918 402325 73154 402561
rect 72918 395325 73154 395561
rect 72918 388325 73154 388561
rect 72918 381325 73154 381561
rect 72918 374325 73154 374561
rect 72918 367325 73154 367561
rect 72918 360325 73154 360561
rect 72918 353325 73154 353561
rect 72918 346325 73154 346561
rect 72918 339325 73154 339561
rect 72918 332325 73154 332561
rect 72918 325325 73154 325561
rect 72918 318325 73154 318561
rect 72918 311325 73154 311561
rect 72918 304325 73154 304561
rect 72918 297325 73154 297561
rect 72918 290325 73154 290561
rect 72918 283325 73154 283561
rect 72918 276325 73154 276561
rect 72918 269325 73154 269561
rect 72918 262325 73154 262561
rect 72918 255325 73154 255561
rect 72918 248325 73154 248561
rect 72918 241325 73154 241561
rect 72918 234325 73154 234561
rect 72918 227325 73154 227561
rect 72918 220325 73154 220561
rect 72918 213325 73154 213561
rect 72918 206325 73154 206561
rect 72918 199325 73154 199561
rect 72918 192325 73154 192561
rect 72918 185325 73154 185561
rect 72918 178325 73154 178561
rect 72918 171325 73154 171561
rect 72918 164325 73154 164561
rect 72918 157325 73154 157561
rect 72918 150325 73154 150561
rect 72918 143325 73154 143561
rect 72918 136325 73154 136561
rect 72918 129325 73154 129561
rect 72918 122325 73154 122561
rect 72918 115325 73154 115561
rect 72918 108325 73154 108561
rect 72918 101325 73154 101561
rect 72918 94325 73154 94561
rect 72918 87325 73154 87561
rect 72918 80325 73154 80561
rect 72918 73325 73154 73561
rect 72918 66325 73154 66561
rect 72918 59325 73154 59561
rect 72918 52325 73154 52561
rect 72918 45325 73154 45561
rect 72918 38325 73154 38561
rect 72918 31325 73154 31561
rect 72918 24325 73154 24561
rect 72918 17325 73154 17561
rect 72918 10325 73154 10561
rect 72918 3325 73154 3561
rect 72918 -1942 73154 -1706
rect 72918 -2262 73154 -2026
rect 78186 705002 78422 705238
rect 78186 704682 78422 704918
rect 78186 695258 78422 695494
rect 78186 688258 78422 688494
rect 78186 681258 78422 681494
rect 78186 674258 78422 674494
rect 78186 667258 78422 667494
rect 78186 660258 78422 660494
rect 78186 653258 78422 653494
rect 78186 646258 78422 646494
rect 78186 639258 78422 639494
rect 78186 632258 78422 632494
rect 78186 625258 78422 625494
rect 78186 618258 78422 618494
rect 78186 611258 78422 611494
rect 78186 604258 78422 604494
rect 78186 597258 78422 597494
rect 78186 590258 78422 590494
rect 78186 583258 78422 583494
rect 78186 576258 78422 576494
rect 78186 569258 78422 569494
rect 78186 562258 78422 562494
rect 78186 555258 78422 555494
rect 78186 548258 78422 548494
rect 78186 541258 78422 541494
rect 78186 534258 78422 534494
rect 78186 527258 78422 527494
rect 78186 520258 78422 520494
rect 78186 513258 78422 513494
rect 78186 506258 78422 506494
rect 78186 499258 78422 499494
rect 78186 492258 78422 492494
rect 78186 485258 78422 485494
rect 78186 478258 78422 478494
rect 78186 471258 78422 471494
rect 78186 464258 78422 464494
rect 78186 457258 78422 457494
rect 78186 450258 78422 450494
rect 78186 443258 78422 443494
rect 78186 436258 78422 436494
rect 78186 429258 78422 429494
rect 78186 422258 78422 422494
rect 78186 415258 78422 415494
rect 78186 408258 78422 408494
rect 78186 401258 78422 401494
rect 78186 394258 78422 394494
rect 78186 387258 78422 387494
rect 78186 380258 78422 380494
rect 78186 373258 78422 373494
rect 78186 366258 78422 366494
rect 78186 359258 78422 359494
rect 78186 352258 78422 352494
rect 78186 345258 78422 345494
rect 78186 338258 78422 338494
rect 78186 331258 78422 331494
rect 78186 324258 78422 324494
rect 78186 317258 78422 317494
rect 78186 310258 78422 310494
rect 78186 303258 78422 303494
rect 78186 296258 78422 296494
rect 78186 289258 78422 289494
rect 78186 282258 78422 282494
rect 78186 275258 78422 275494
rect 78186 268258 78422 268494
rect 78186 261258 78422 261494
rect 78186 254258 78422 254494
rect 78186 247258 78422 247494
rect 78186 240258 78422 240494
rect 78186 233258 78422 233494
rect 78186 226258 78422 226494
rect 78186 219258 78422 219494
rect 78186 212258 78422 212494
rect 78186 205258 78422 205494
rect 78186 198258 78422 198494
rect 78186 191258 78422 191494
rect 78186 184258 78422 184494
rect 78186 177258 78422 177494
rect 78186 170258 78422 170494
rect 78186 163258 78422 163494
rect 78186 156258 78422 156494
rect 78186 149258 78422 149494
rect 78186 142258 78422 142494
rect 78186 135258 78422 135494
rect 78186 128258 78422 128494
rect 78186 121258 78422 121494
rect 78186 114258 78422 114494
rect 78186 107258 78422 107494
rect 78186 100258 78422 100494
rect 78186 93258 78422 93494
rect 78186 86258 78422 86494
rect 78186 79258 78422 79494
rect 78186 72258 78422 72494
rect 78186 65258 78422 65494
rect 78186 58258 78422 58494
rect 78186 51258 78422 51494
rect 78186 44258 78422 44494
rect 78186 37258 78422 37494
rect 78186 30258 78422 30494
rect 78186 23258 78422 23494
rect 78186 16258 78422 16494
rect 78186 9258 78422 9494
rect 78186 2258 78422 2494
rect 78186 -982 78422 -746
rect 78186 -1302 78422 -1066
rect 79918 705962 80154 706198
rect 79918 705642 80154 705878
rect 79918 696325 80154 696561
rect 79918 689325 80154 689561
rect 79918 682325 80154 682561
rect 79918 675325 80154 675561
rect 79918 668325 80154 668561
rect 79918 661325 80154 661561
rect 79918 654325 80154 654561
rect 79918 647325 80154 647561
rect 79918 640325 80154 640561
rect 79918 633325 80154 633561
rect 79918 626325 80154 626561
rect 79918 619325 80154 619561
rect 79918 612325 80154 612561
rect 79918 605325 80154 605561
rect 79918 598325 80154 598561
rect 79918 591325 80154 591561
rect 79918 584325 80154 584561
rect 79918 577325 80154 577561
rect 79918 570325 80154 570561
rect 79918 563325 80154 563561
rect 79918 556325 80154 556561
rect 79918 549325 80154 549561
rect 79918 542325 80154 542561
rect 79918 535325 80154 535561
rect 79918 528325 80154 528561
rect 79918 521325 80154 521561
rect 79918 514325 80154 514561
rect 79918 507325 80154 507561
rect 79918 500325 80154 500561
rect 79918 493325 80154 493561
rect 79918 486325 80154 486561
rect 79918 479325 80154 479561
rect 79918 472325 80154 472561
rect 79918 465325 80154 465561
rect 79918 458325 80154 458561
rect 79918 451325 80154 451561
rect 79918 444325 80154 444561
rect 79918 437325 80154 437561
rect 79918 430325 80154 430561
rect 79918 423325 80154 423561
rect 79918 416325 80154 416561
rect 79918 409325 80154 409561
rect 79918 402325 80154 402561
rect 79918 395325 80154 395561
rect 79918 388325 80154 388561
rect 79918 381325 80154 381561
rect 79918 374325 80154 374561
rect 79918 367325 80154 367561
rect 79918 360325 80154 360561
rect 79918 353325 80154 353561
rect 79918 346325 80154 346561
rect 79918 339325 80154 339561
rect 79918 332325 80154 332561
rect 79918 325325 80154 325561
rect 79918 318325 80154 318561
rect 79918 311325 80154 311561
rect 79918 304325 80154 304561
rect 79918 297325 80154 297561
rect 79918 290325 80154 290561
rect 79918 283325 80154 283561
rect 79918 276325 80154 276561
rect 79918 269325 80154 269561
rect 79918 262325 80154 262561
rect 79918 255325 80154 255561
rect 79918 248325 80154 248561
rect 79918 241325 80154 241561
rect 79918 234325 80154 234561
rect 79918 227325 80154 227561
rect 79918 220325 80154 220561
rect 79918 213325 80154 213561
rect 79918 206325 80154 206561
rect 79918 199325 80154 199561
rect 79918 192325 80154 192561
rect 79918 185325 80154 185561
rect 79918 178325 80154 178561
rect 79918 171325 80154 171561
rect 79918 164325 80154 164561
rect 79918 157325 80154 157561
rect 79918 150325 80154 150561
rect 79918 143325 80154 143561
rect 79918 136325 80154 136561
rect 79918 129325 80154 129561
rect 79918 122325 80154 122561
rect 79918 115325 80154 115561
rect 79918 108325 80154 108561
rect 79918 101325 80154 101561
rect 79918 94325 80154 94561
rect 79918 87325 80154 87561
rect 79918 80325 80154 80561
rect 79918 73325 80154 73561
rect 79918 66325 80154 66561
rect 79918 59325 80154 59561
rect 79918 52325 80154 52561
rect 79918 45325 80154 45561
rect 79918 38325 80154 38561
rect 79918 31325 80154 31561
rect 79918 24325 80154 24561
rect 79918 17325 80154 17561
rect 79918 10325 80154 10561
rect 79918 3325 80154 3561
rect 79918 -1942 80154 -1706
rect 79918 -2262 80154 -2026
rect 85186 705002 85422 705238
rect 85186 704682 85422 704918
rect 85186 695258 85422 695494
rect 85186 688258 85422 688494
rect 85186 681258 85422 681494
rect 85186 674258 85422 674494
rect 85186 667258 85422 667494
rect 85186 660258 85422 660494
rect 85186 653258 85422 653494
rect 85186 646258 85422 646494
rect 85186 639258 85422 639494
rect 85186 632258 85422 632494
rect 85186 625258 85422 625494
rect 85186 618258 85422 618494
rect 85186 611258 85422 611494
rect 85186 604258 85422 604494
rect 85186 597258 85422 597494
rect 85186 590258 85422 590494
rect 85186 583258 85422 583494
rect 85186 576258 85422 576494
rect 85186 569258 85422 569494
rect 85186 562258 85422 562494
rect 85186 555258 85422 555494
rect 85186 548258 85422 548494
rect 85186 541258 85422 541494
rect 85186 534258 85422 534494
rect 85186 527258 85422 527494
rect 85186 520258 85422 520494
rect 85186 513258 85422 513494
rect 85186 506258 85422 506494
rect 85186 499258 85422 499494
rect 85186 492258 85422 492494
rect 85186 485258 85422 485494
rect 85186 478258 85422 478494
rect 85186 471258 85422 471494
rect 85186 464258 85422 464494
rect 85186 457258 85422 457494
rect 85186 450258 85422 450494
rect 85186 443258 85422 443494
rect 85186 436258 85422 436494
rect 85186 429258 85422 429494
rect 85186 422258 85422 422494
rect 85186 415258 85422 415494
rect 85186 408258 85422 408494
rect 85186 401258 85422 401494
rect 85186 394258 85422 394494
rect 85186 387258 85422 387494
rect 85186 380258 85422 380494
rect 85186 373258 85422 373494
rect 85186 366258 85422 366494
rect 85186 359258 85422 359494
rect 85186 352258 85422 352494
rect 85186 345258 85422 345494
rect 85186 338258 85422 338494
rect 85186 331258 85422 331494
rect 85186 324258 85422 324494
rect 85186 317258 85422 317494
rect 85186 310258 85422 310494
rect 85186 303258 85422 303494
rect 85186 296258 85422 296494
rect 85186 289258 85422 289494
rect 85186 282258 85422 282494
rect 85186 275258 85422 275494
rect 85186 268258 85422 268494
rect 85186 261258 85422 261494
rect 85186 254258 85422 254494
rect 85186 247258 85422 247494
rect 85186 240258 85422 240494
rect 85186 233258 85422 233494
rect 85186 226258 85422 226494
rect 85186 219258 85422 219494
rect 85186 212258 85422 212494
rect 85186 205258 85422 205494
rect 85186 198258 85422 198494
rect 85186 191258 85422 191494
rect 85186 184258 85422 184494
rect 85186 177258 85422 177494
rect 85186 170258 85422 170494
rect 85186 163258 85422 163494
rect 85186 156258 85422 156494
rect 85186 149258 85422 149494
rect 85186 142258 85422 142494
rect 85186 135258 85422 135494
rect 85186 128258 85422 128494
rect 85186 121258 85422 121494
rect 85186 114258 85422 114494
rect 85186 107258 85422 107494
rect 85186 100258 85422 100494
rect 85186 93258 85422 93494
rect 85186 86258 85422 86494
rect 85186 79258 85422 79494
rect 85186 72258 85422 72494
rect 85186 65258 85422 65494
rect 85186 58258 85422 58494
rect 85186 51258 85422 51494
rect 85186 44258 85422 44494
rect 85186 37258 85422 37494
rect 85186 30258 85422 30494
rect 85186 23258 85422 23494
rect 85186 16258 85422 16494
rect 85186 9258 85422 9494
rect 85186 2258 85422 2494
rect 85186 -982 85422 -746
rect 85186 -1302 85422 -1066
rect 86918 705962 87154 706198
rect 86918 705642 87154 705878
rect 86918 696325 87154 696561
rect 86918 689325 87154 689561
rect 86918 682325 87154 682561
rect 86918 675325 87154 675561
rect 86918 668325 87154 668561
rect 86918 661325 87154 661561
rect 86918 654325 87154 654561
rect 86918 647325 87154 647561
rect 86918 640325 87154 640561
rect 86918 633325 87154 633561
rect 86918 626325 87154 626561
rect 86918 619325 87154 619561
rect 86918 612325 87154 612561
rect 86918 605325 87154 605561
rect 86918 598325 87154 598561
rect 86918 591325 87154 591561
rect 86918 584325 87154 584561
rect 86918 577325 87154 577561
rect 86918 570325 87154 570561
rect 86918 563325 87154 563561
rect 86918 556325 87154 556561
rect 86918 549325 87154 549561
rect 86918 542325 87154 542561
rect 86918 535325 87154 535561
rect 86918 528325 87154 528561
rect 86918 521325 87154 521561
rect 86918 514325 87154 514561
rect 86918 507325 87154 507561
rect 86918 500325 87154 500561
rect 86918 493325 87154 493561
rect 86918 486325 87154 486561
rect 86918 479325 87154 479561
rect 86918 472325 87154 472561
rect 86918 465325 87154 465561
rect 86918 458325 87154 458561
rect 86918 451325 87154 451561
rect 86918 444325 87154 444561
rect 86918 437325 87154 437561
rect 86918 430325 87154 430561
rect 86918 423325 87154 423561
rect 86918 416325 87154 416561
rect 86918 409325 87154 409561
rect 86918 402325 87154 402561
rect 86918 395325 87154 395561
rect 86918 388325 87154 388561
rect 86918 381325 87154 381561
rect 86918 374325 87154 374561
rect 86918 367325 87154 367561
rect 86918 360325 87154 360561
rect 86918 353325 87154 353561
rect 86918 346325 87154 346561
rect 86918 339325 87154 339561
rect 86918 332325 87154 332561
rect 86918 325325 87154 325561
rect 86918 318325 87154 318561
rect 86918 311325 87154 311561
rect 86918 304325 87154 304561
rect 86918 297325 87154 297561
rect 86918 290325 87154 290561
rect 86918 283325 87154 283561
rect 86918 276325 87154 276561
rect 86918 269325 87154 269561
rect 86918 262325 87154 262561
rect 86918 255325 87154 255561
rect 86918 248325 87154 248561
rect 86918 241325 87154 241561
rect 86918 234325 87154 234561
rect 86918 227325 87154 227561
rect 86918 220325 87154 220561
rect 86918 213325 87154 213561
rect 86918 206325 87154 206561
rect 86918 199325 87154 199561
rect 86918 192325 87154 192561
rect 86918 185325 87154 185561
rect 86918 178325 87154 178561
rect 86918 171325 87154 171561
rect 86918 164325 87154 164561
rect 86918 157325 87154 157561
rect 86918 150325 87154 150561
rect 86918 143325 87154 143561
rect 86918 136325 87154 136561
rect 86918 129325 87154 129561
rect 86918 122325 87154 122561
rect 86918 115325 87154 115561
rect 86918 108325 87154 108561
rect 86918 101325 87154 101561
rect 86918 94325 87154 94561
rect 86918 87325 87154 87561
rect 86918 80325 87154 80561
rect 86918 73325 87154 73561
rect 86918 66325 87154 66561
rect 86918 59325 87154 59561
rect 86918 52325 87154 52561
rect 86918 45325 87154 45561
rect 86918 38325 87154 38561
rect 86918 31325 87154 31561
rect 86918 24325 87154 24561
rect 86918 17325 87154 17561
rect 86918 10325 87154 10561
rect 86918 3325 87154 3561
rect 86918 -1942 87154 -1706
rect 86918 -2262 87154 -2026
rect 92186 705002 92422 705238
rect 92186 704682 92422 704918
rect 92186 695258 92422 695494
rect 92186 688258 92422 688494
rect 92186 681258 92422 681494
rect 92186 674258 92422 674494
rect 92186 667258 92422 667494
rect 92186 660258 92422 660494
rect 92186 653258 92422 653494
rect 92186 646258 92422 646494
rect 92186 639258 92422 639494
rect 92186 632258 92422 632494
rect 92186 625258 92422 625494
rect 92186 618258 92422 618494
rect 92186 611258 92422 611494
rect 92186 604258 92422 604494
rect 92186 597258 92422 597494
rect 92186 590258 92422 590494
rect 92186 583258 92422 583494
rect 92186 576258 92422 576494
rect 92186 569258 92422 569494
rect 92186 562258 92422 562494
rect 92186 555258 92422 555494
rect 92186 548258 92422 548494
rect 92186 541258 92422 541494
rect 92186 534258 92422 534494
rect 92186 527258 92422 527494
rect 92186 520258 92422 520494
rect 92186 513258 92422 513494
rect 92186 506258 92422 506494
rect 92186 499258 92422 499494
rect 92186 492258 92422 492494
rect 92186 485258 92422 485494
rect 92186 478258 92422 478494
rect 92186 471258 92422 471494
rect 92186 464258 92422 464494
rect 92186 457258 92422 457494
rect 92186 450258 92422 450494
rect 92186 443258 92422 443494
rect 92186 436258 92422 436494
rect 92186 429258 92422 429494
rect 92186 422258 92422 422494
rect 92186 415258 92422 415494
rect 92186 408258 92422 408494
rect 92186 401258 92422 401494
rect 92186 394258 92422 394494
rect 92186 387258 92422 387494
rect 92186 380258 92422 380494
rect 92186 373258 92422 373494
rect 92186 366258 92422 366494
rect 92186 359258 92422 359494
rect 92186 352258 92422 352494
rect 92186 345258 92422 345494
rect 92186 338258 92422 338494
rect 92186 331258 92422 331494
rect 92186 324258 92422 324494
rect 92186 317258 92422 317494
rect 92186 310258 92422 310494
rect 92186 303258 92422 303494
rect 92186 296258 92422 296494
rect 92186 289258 92422 289494
rect 92186 282258 92422 282494
rect 92186 275258 92422 275494
rect 92186 268258 92422 268494
rect 92186 261258 92422 261494
rect 92186 254258 92422 254494
rect 92186 247258 92422 247494
rect 92186 240258 92422 240494
rect 92186 233258 92422 233494
rect 92186 226258 92422 226494
rect 92186 219258 92422 219494
rect 92186 212258 92422 212494
rect 92186 205258 92422 205494
rect 92186 198258 92422 198494
rect 92186 191258 92422 191494
rect 92186 184258 92422 184494
rect 92186 177258 92422 177494
rect 92186 170258 92422 170494
rect 92186 163258 92422 163494
rect 92186 156258 92422 156494
rect 92186 149258 92422 149494
rect 92186 142258 92422 142494
rect 92186 135258 92422 135494
rect 92186 128258 92422 128494
rect 92186 121258 92422 121494
rect 92186 114258 92422 114494
rect 92186 107258 92422 107494
rect 92186 100258 92422 100494
rect 92186 93258 92422 93494
rect 92186 86258 92422 86494
rect 92186 79258 92422 79494
rect 92186 72258 92422 72494
rect 92186 65258 92422 65494
rect 92186 58258 92422 58494
rect 92186 51258 92422 51494
rect 92186 44258 92422 44494
rect 92186 37258 92422 37494
rect 92186 30258 92422 30494
rect 92186 23258 92422 23494
rect 92186 16258 92422 16494
rect 92186 9258 92422 9494
rect 92186 2258 92422 2494
rect 92186 -982 92422 -746
rect 92186 -1302 92422 -1066
rect 93918 705962 94154 706198
rect 93918 705642 94154 705878
rect 93918 696325 94154 696561
rect 93918 689325 94154 689561
rect 93918 682325 94154 682561
rect 93918 675325 94154 675561
rect 93918 668325 94154 668561
rect 93918 661325 94154 661561
rect 93918 654325 94154 654561
rect 93918 647325 94154 647561
rect 93918 640325 94154 640561
rect 93918 633325 94154 633561
rect 93918 626325 94154 626561
rect 93918 619325 94154 619561
rect 93918 612325 94154 612561
rect 93918 605325 94154 605561
rect 93918 598325 94154 598561
rect 93918 591325 94154 591561
rect 93918 584325 94154 584561
rect 93918 577325 94154 577561
rect 93918 570325 94154 570561
rect 93918 563325 94154 563561
rect 93918 556325 94154 556561
rect 93918 549325 94154 549561
rect 93918 542325 94154 542561
rect 93918 535325 94154 535561
rect 93918 528325 94154 528561
rect 93918 521325 94154 521561
rect 93918 514325 94154 514561
rect 93918 507325 94154 507561
rect 93918 500325 94154 500561
rect 93918 493325 94154 493561
rect 93918 486325 94154 486561
rect 93918 479325 94154 479561
rect 93918 472325 94154 472561
rect 93918 465325 94154 465561
rect 93918 458325 94154 458561
rect 93918 451325 94154 451561
rect 93918 444325 94154 444561
rect 93918 437325 94154 437561
rect 93918 430325 94154 430561
rect 93918 423325 94154 423561
rect 93918 416325 94154 416561
rect 93918 409325 94154 409561
rect 93918 402325 94154 402561
rect 93918 395325 94154 395561
rect 93918 388325 94154 388561
rect 93918 381325 94154 381561
rect 93918 374325 94154 374561
rect 93918 367325 94154 367561
rect 93918 360325 94154 360561
rect 93918 353325 94154 353561
rect 93918 346325 94154 346561
rect 93918 339325 94154 339561
rect 93918 332325 94154 332561
rect 93918 325325 94154 325561
rect 93918 318325 94154 318561
rect 93918 311325 94154 311561
rect 93918 304325 94154 304561
rect 93918 297325 94154 297561
rect 93918 290325 94154 290561
rect 93918 283325 94154 283561
rect 93918 276325 94154 276561
rect 93918 269325 94154 269561
rect 93918 262325 94154 262561
rect 93918 255325 94154 255561
rect 93918 248325 94154 248561
rect 93918 241325 94154 241561
rect 93918 234325 94154 234561
rect 93918 227325 94154 227561
rect 93918 220325 94154 220561
rect 93918 213325 94154 213561
rect 93918 206325 94154 206561
rect 93918 199325 94154 199561
rect 93918 192325 94154 192561
rect 93918 185325 94154 185561
rect 93918 178325 94154 178561
rect 93918 171325 94154 171561
rect 93918 164325 94154 164561
rect 93918 157325 94154 157561
rect 93918 150325 94154 150561
rect 93918 143325 94154 143561
rect 93918 136325 94154 136561
rect 93918 129325 94154 129561
rect 93918 122325 94154 122561
rect 93918 115325 94154 115561
rect 93918 108325 94154 108561
rect 93918 101325 94154 101561
rect 93918 94325 94154 94561
rect 93918 87325 94154 87561
rect 93918 80325 94154 80561
rect 93918 73325 94154 73561
rect 93918 66325 94154 66561
rect 93918 59325 94154 59561
rect 93918 52325 94154 52561
rect 93918 45325 94154 45561
rect 93918 38325 94154 38561
rect 93918 31325 94154 31561
rect 93918 24325 94154 24561
rect 93918 17325 94154 17561
rect 93918 10325 94154 10561
rect 93918 3325 94154 3561
rect 93918 -1942 94154 -1706
rect 93918 -2262 94154 -2026
rect 99186 705002 99422 705238
rect 99186 704682 99422 704918
rect 99186 695258 99422 695494
rect 99186 688258 99422 688494
rect 99186 681258 99422 681494
rect 99186 674258 99422 674494
rect 99186 667258 99422 667494
rect 99186 660258 99422 660494
rect 99186 653258 99422 653494
rect 99186 646258 99422 646494
rect 99186 639258 99422 639494
rect 99186 632258 99422 632494
rect 99186 625258 99422 625494
rect 99186 618258 99422 618494
rect 99186 611258 99422 611494
rect 99186 604258 99422 604494
rect 99186 597258 99422 597494
rect 99186 590258 99422 590494
rect 99186 583258 99422 583494
rect 99186 576258 99422 576494
rect 99186 569258 99422 569494
rect 99186 562258 99422 562494
rect 99186 555258 99422 555494
rect 99186 548258 99422 548494
rect 99186 541258 99422 541494
rect 99186 534258 99422 534494
rect 99186 527258 99422 527494
rect 99186 520258 99422 520494
rect 99186 513258 99422 513494
rect 99186 506258 99422 506494
rect 99186 499258 99422 499494
rect 99186 492258 99422 492494
rect 99186 485258 99422 485494
rect 99186 478258 99422 478494
rect 99186 471258 99422 471494
rect 99186 464258 99422 464494
rect 99186 457258 99422 457494
rect 99186 450258 99422 450494
rect 99186 443258 99422 443494
rect 99186 436258 99422 436494
rect 99186 429258 99422 429494
rect 99186 422258 99422 422494
rect 99186 415258 99422 415494
rect 99186 408258 99422 408494
rect 99186 401258 99422 401494
rect 99186 394258 99422 394494
rect 99186 387258 99422 387494
rect 99186 380258 99422 380494
rect 99186 373258 99422 373494
rect 99186 366258 99422 366494
rect 99186 359258 99422 359494
rect 99186 352258 99422 352494
rect 99186 345258 99422 345494
rect 99186 338258 99422 338494
rect 99186 331258 99422 331494
rect 99186 324258 99422 324494
rect 99186 317258 99422 317494
rect 99186 310258 99422 310494
rect 99186 303258 99422 303494
rect 99186 296258 99422 296494
rect 99186 289258 99422 289494
rect 99186 282258 99422 282494
rect 99186 275258 99422 275494
rect 99186 268258 99422 268494
rect 99186 261258 99422 261494
rect 99186 254258 99422 254494
rect 99186 247258 99422 247494
rect 99186 240258 99422 240494
rect 99186 233258 99422 233494
rect 99186 226258 99422 226494
rect 99186 219258 99422 219494
rect 99186 212258 99422 212494
rect 99186 205258 99422 205494
rect 99186 198258 99422 198494
rect 99186 191258 99422 191494
rect 99186 184258 99422 184494
rect 99186 177258 99422 177494
rect 99186 170258 99422 170494
rect 99186 163258 99422 163494
rect 99186 156258 99422 156494
rect 99186 149258 99422 149494
rect 99186 142258 99422 142494
rect 99186 135258 99422 135494
rect 99186 128258 99422 128494
rect 99186 121258 99422 121494
rect 99186 114258 99422 114494
rect 99186 107258 99422 107494
rect 99186 100258 99422 100494
rect 99186 93258 99422 93494
rect 99186 86258 99422 86494
rect 99186 79258 99422 79494
rect 99186 72258 99422 72494
rect 99186 65258 99422 65494
rect 99186 58258 99422 58494
rect 99186 51258 99422 51494
rect 99186 44258 99422 44494
rect 99186 37258 99422 37494
rect 99186 30258 99422 30494
rect 99186 23258 99422 23494
rect 99186 16258 99422 16494
rect 99186 9258 99422 9494
rect 99186 2258 99422 2494
rect 99186 -982 99422 -746
rect 99186 -1302 99422 -1066
rect 100918 705962 101154 706198
rect 100918 705642 101154 705878
rect 100918 696325 101154 696561
rect 100918 689325 101154 689561
rect 100918 682325 101154 682561
rect 100918 675325 101154 675561
rect 100918 668325 101154 668561
rect 100918 661325 101154 661561
rect 100918 654325 101154 654561
rect 100918 647325 101154 647561
rect 100918 640325 101154 640561
rect 100918 633325 101154 633561
rect 100918 626325 101154 626561
rect 100918 619325 101154 619561
rect 100918 612325 101154 612561
rect 100918 605325 101154 605561
rect 100918 598325 101154 598561
rect 100918 591325 101154 591561
rect 100918 584325 101154 584561
rect 100918 577325 101154 577561
rect 100918 570325 101154 570561
rect 100918 563325 101154 563561
rect 100918 556325 101154 556561
rect 100918 549325 101154 549561
rect 100918 542325 101154 542561
rect 100918 535325 101154 535561
rect 100918 528325 101154 528561
rect 100918 521325 101154 521561
rect 100918 514325 101154 514561
rect 100918 507325 101154 507561
rect 100918 500325 101154 500561
rect 100918 493325 101154 493561
rect 100918 486325 101154 486561
rect 100918 479325 101154 479561
rect 100918 472325 101154 472561
rect 100918 465325 101154 465561
rect 100918 458325 101154 458561
rect 100918 451325 101154 451561
rect 100918 444325 101154 444561
rect 100918 437325 101154 437561
rect 100918 430325 101154 430561
rect 100918 423325 101154 423561
rect 100918 416325 101154 416561
rect 100918 409325 101154 409561
rect 100918 402325 101154 402561
rect 100918 395325 101154 395561
rect 100918 388325 101154 388561
rect 100918 381325 101154 381561
rect 100918 374325 101154 374561
rect 100918 367325 101154 367561
rect 100918 360325 101154 360561
rect 100918 353325 101154 353561
rect 100918 346325 101154 346561
rect 100918 339325 101154 339561
rect 100918 332325 101154 332561
rect 100918 325325 101154 325561
rect 100918 318325 101154 318561
rect 100918 311325 101154 311561
rect 100918 304325 101154 304561
rect 100918 297325 101154 297561
rect 100918 290325 101154 290561
rect 100918 283325 101154 283561
rect 100918 276325 101154 276561
rect 100918 269325 101154 269561
rect 100918 262325 101154 262561
rect 100918 255325 101154 255561
rect 100918 248325 101154 248561
rect 100918 241325 101154 241561
rect 100918 234325 101154 234561
rect 100918 227325 101154 227561
rect 100918 220325 101154 220561
rect 100918 213325 101154 213561
rect 100918 206325 101154 206561
rect 100918 199325 101154 199561
rect 100918 192325 101154 192561
rect 100918 185325 101154 185561
rect 100918 178325 101154 178561
rect 100918 171325 101154 171561
rect 100918 164325 101154 164561
rect 100918 157325 101154 157561
rect 100918 150325 101154 150561
rect 100918 143325 101154 143561
rect 100918 136325 101154 136561
rect 100918 129325 101154 129561
rect 100918 122325 101154 122561
rect 100918 115325 101154 115561
rect 100918 108325 101154 108561
rect 100918 101325 101154 101561
rect 100918 94325 101154 94561
rect 100918 87325 101154 87561
rect 100918 80325 101154 80561
rect 100918 73325 101154 73561
rect 100918 66325 101154 66561
rect 100918 59325 101154 59561
rect 100918 52325 101154 52561
rect 100918 45325 101154 45561
rect 100918 38325 101154 38561
rect 100918 31325 101154 31561
rect 100918 24325 101154 24561
rect 100918 17325 101154 17561
rect 100918 10325 101154 10561
rect 100918 3325 101154 3561
rect 100918 -1942 101154 -1706
rect 100918 -2262 101154 -2026
rect 106186 705002 106422 705238
rect 106186 704682 106422 704918
rect 106186 695258 106422 695494
rect 106186 688258 106422 688494
rect 106186 681258 106422 681494
rect 106186 674258 106422 674494
rect 106186 667258 106422 667494
rect 106186 660258 106422 660494
rect 106186 653258 106422 653494
rect 106186 646258 106422 646494
rect 106186 639258 106422 639494
rect 106186 632258 106422 632494
rect 106186 625258 106422 625494
rect 106186 618258 106422 618494
rect 106186 611258 106422 611494
rect 106186 604258 106422 604494
rect 106186 597258 106422 597494
rect 106186 590258 106422 590494
rect 106186 583258 106422 583494
rect 106186 576258 106422 576494
rect 106186 569258 106422 569494
rect 106186 562258 106422 562494
rect 106186 555258 106422 555494
rect 106186 548258 106422 548494
rect 106186 541258 106422 541494
rect 106186 534258 106422 534494
rect 106186 527258 106422 527494
rect 106186 520258 106422 520494
rect 106186 513258 106422 513494
rect 106186 506258 106422 506494
rect 106186 499258 106422 499494
rect 106186 492258 106422 492494
rect 106186 485258 106422 485494
rect 106186 478258 106422 478494
rect 106186 471258 106422 471494
rect 106186 464258 106422 464494
rect 106186 457258 106422 457494
rect 106186 450258 106422 450494
rect 106186 443258 106422 443494
rect 106186 436258 106422 436494
rect 106186 429258 106422 429494
rect 106186 422258 106422 422494
rect 106186 415258 106422 415494
rect 106186 408258 106422 408494
rect 106186 401258 106422 401494
rect 106186 394258 106422 394494
rect 106186 387258 106422 387494
rect 106186 380258 106422 380494
rect 106186 373258 106422 373494
rect 106186 366258 106422 366494
rect 106186 359258 106422 359494
rect 106186 352258 106422 352494
rect 106186 345258 106422 345494
rect 106186 338258 106422 338494
rect 106186 331258 106422 331494
rect 106186 324258 106422 324494
rect 106186 317258 106422 317494
rect 106186 310258 106422 310494
rect 106186 303258 106422 303494
rect 106186 296258 106422 296494
rect 106186 289258 106422 289494
rect 106186 282258 106422 282494
rect 106186 275258 106422 275494
rect 106186 268258 106422 268494
rect 106186 261258 106422 261494
rect 106186 254258 106422 254494
rect 106186 247258 106422 247494
rect 106186 240258 106422 240494
rect 106186 233258 106422 233494
rect 106186 226258 106422 226494
rect 106186 219258 106422 219494
rect 106186 212258 106422 212494
rect 106186 205258 106422 205494
rect 106186 198258 106422 198494
rect 106186 191258 106422 191494
rect 106186 184258 106422 184494
rect 106186 177258 106422 177494
rect 106186 170258 106422 170494
rect 106186 163258 106422 163494
rect 106186 156258 106422 156494
rect 106186 149258 106422 149494
rect 106186 142258 106422 142494
rect 106186 135258 106422 135494
rect 106186 128258 106422 128494
rect 106186 121258 106422 121494
rect 106186 114258 106422 114494
rect 106186 107258 106422 107494
rect 106186 100258 106422 100494
rect 106186 93258 106422 93494
rect 106186 86258 106422 86494
rect 106186 79258 106422 79494
rect 106186 72258 106422 72494
rect 106186 65258 106422 65494
rect 106186 58258 106422 58494
rect 106186 51258 106422 51494
rect 106186 44258 106422 44494
rect 106186 37258 106422 37494
rect 106186 30258 106422 30494
rect 106186 23258 106422 23494
rect 106186 16258 106422 16494
rect 106186 9258 106422 9494
rect 106186 2258 106422 2494
rect 106186 -982 106422 -746
rect 106186 -1302 106422 -1066
rect 107918 705962 108154 706198
rect 107918 705642 108154 705878
rect 107918 696325 108154 696561
rect 107918 689325 108154 689561
rect 107918 682325 108154 682561
rect 107918 675325 108154 675561
rect 107918 668325 108154 668561
rect 107918 661325 108154 661561
rect 107918 654325 108154 654561
rect 107918 647325 108154 647561
rect 107918 640325 108154 640561
rect 107918 633325 108154 633561
rect 107918 626325 108154 626561
rect 107918 619325 108154 619561
rect 107918 612325 108154 612561
rect 107918 605325 108154 605561
rect 107918 598325 108154 598561
rect 107918 591325 108154 591561
rect 107918 584325 108154 584561
rect 107918 577325 108154 577561
rect 107918 570325 108154 570561
rect 107918 563325 108154 563561
rect 107918 556325 108154 556561
rect 107918 549325 108154 549561
rect 107918 542325 108154 542561
rect 107918 535325 108154 535561
rect 107918 528325 108154 528561
rect 107918 521325 108154 521561
rect 107918 514325 108154 514561
rect 107918 507325 108154 507561
rect 107918 500325 108154 500561
rect 107918 493325 108154 493561
rect 107918 486325 108154 486561
rect 107918 479325 108154 479561
rect 107918 472325 108154 472561
rect 107918 465325 108154 465561
rect 107918 458325 108154 458561
rect 107918 451325 108154 451561
rect 107918 444325 108154 444561
rect 107918 437325 108154 437561
rect 107918 430325 108154 430561
rect 107918 423325 108154 423561
rect 107918 416325 108154 416561
rect 107918 409325 108154 409561
rect 107918 402325 108154 402561
rect 107918 395325 108154 395561
rect 107918 388325 108154 388561
rect 107918 381325 108154 381561
rect 107918 374325 108154 374561
rect 107918 367325 108154 367561
rect 107918 360325 108154 360561
rect 107918 353325 108154 353561
rect 107918 346325 108154 346561
rect 107918 339325 108154 339561
rect 107918 332325 108154 332561
rect 107918 325325 108154 325561
rect 107918 318325 108154 318561
rect 107918 311325 108154 311561
rect 107918 304325 108154 304561
rect 107918 297325 108154 297561
rect 107918 290325 108154 290561
rect 107918 283325 108154 283561
rect 107918 276325 108154 276561
rect 107918 269325 108154 269561
rect 107918 262325 108154 262561
rect 107918 255325 108154 255561
rect 107918 248325 108154 248561
rect 107918 241325 108154 241561
rect 107918 234325 108154 234561
rect 107918 227325 108154 227561
rect 107918 220325 108154 220561
rect 107918 213325 108154 213561
rect 107918 206325 108154 206561
rect 107918 199325 108154 199561
rect 107918 192325 108154 192561
rect 107918 185325 108154 185561
rect 107918 178325 108154 178561
rect 107918 171325 108154 171561
rect 107918 164325 108154 164561
rect 107918 157325 108154 157561
rect 107918 150325 108154 150561
rect 107918 143325 108154 143561
rect 107918 136325 108154 136561
rect 107918 129325 108154 129561
rect 107918 122325 108154 122561
rect 107918 115325 108154 115561
rect 107918 108325 108154 108561
rect 107918 101325 108154 101561
rect 107918 94325 108154 94561
rect 107918 87325 108154 87561
rect 107918 80325 108154 80561
rect 107918 73325 108154 73561
rect 107918 66325 108154 66561
rect 107918 59325 108154 59561
rect 107918 52325 108154 52561
rect 107918 45325 108154 45561
rect 107918 38325 108154 38561
rect 107918 31325 108154 31561
rect 107918 24325 108154 24561
rect 107918 17325 108154 17561
rect 107918 10325 108154 10561
rect 107918 3325 108154 3561
rect 107918 -1942 108154 -1706
rect 107918 -2262 108154 -2026
rect 113186 705002 113422 705238
rect 113186 704682 113422 704918
rect 113186 695258 113422 695494
rect 113186 688258 113422 688494
rect 113186 681258 113422 681494
rect 113186 674258 113422 674494
rect 113186 667258 113422 667494
rect 113186 660258 113422 660494
rect 113186 653258 113422 653494
rect 113186 646258 113422 646494
rect 113186 639258 113422 639494
rect 113186 632258 113422 632494
rect 113186 625258 113422 625494
rect 113186 618258 113422 618494
rect 113186 611258 113422 611494
rect 113186 604258 113422 604494
rect 113186 597258 113422 597494
rect 113186 590258 113422 590494
rect 113186 583258 113422 583494
rect 113186 576258 113422 576494
rect 113186 569258 113422 569494
rect 113186 562258 113422 562494
rect 113186 555258 113422 555494
rect 113186 548258 113422 548494
rect 113186 541258 113422 541494
rect 113186 534258 113422 534494
rect 113186 527258 113422 527494
rect 113186 520258 113422 520494
rect 113186 513258 113422 513494
rect 113186 506258 113422 506494
rect 113186 499258 113422 499494
rect 113186 492258 113422 492494
rect 113186 485258 113422 485494
rect 113186 478258 113422 478494
rect 113186 471258 113422 471494
rect 113186 464258 113422 464494
rect 113186 457258 113422 457494
rect 113186 450258 113422 450494
rect 113186 443258 113422 443494
rect 113186 436258 113422 436494
rect 113186 429258 113422 429494
rect 113186 422258 113422 422494
rect 113186 415258 113422 415494
rect 113186 408258 113422 408494
rect 113186 401258 113422 401494
rect 113186 394258 113422 394494
rect 113186 387258 113422 387494
rect 113186 380258 113422 380494
rect 113186 373258 113422 373494
rect 113186 366258 113422 366494
rect 113186 359258 113422 359494
rect 113186 352258 113422 352494
rect 113186 345258 113422 345494
rect 113186 338258 113422 338494
rect 113186 331258 113422 331494
rect 113186 324258 113422 324494
rect 113186 317258 113422 317494
rect 113186 310258 113422 310494
rect 113186 303258 113422 303494
rect 113186 296258 113422 296494
rect 113186 289258 113422 289494
rect 113186 282258 113422 282494
rect 113186 275258 113422 275494
rect 113186 268258 113422 268494
rect 113186 261258 113422 261494
rect 113186 254258 113422 254494
rect 113186 247258 113422 247494
rect 113186 240258 113422 240494
rect 113186 233258 113422 233494
rect 113186 226258 113422 226494
rect 113186 219258 113422 219494
rect 113186 212258 113422 212494
rect 113186 205258 113422 205494
rect 113186 198258 113422 198494
rect 113186 191258 113422 191494
rect 113186 184258 113422 184494
rect 113186 177258 113422 177494
rect 113186 170258 113422 170494
rect 113186 163258 113422 163494
rect 113186 156258 113422 156494
rect 113186 149258 113422 149494
rect 113186 142258 113422 142494
rect 113186 135258 113422 135494
rect 113186 128258 113422 128494
rect 113186 121258 113422 121494
rect 113186 114258 113422 114494
rect 113186 107258 113422 107494
rect 113186 100258 113422 100494
rect 113186 93258 113422 93494
rect 113186 86258 113422 86494
rect 113186 79258 113422 79494
rect 113186 72258 113422 72494
rect 113186 65258 113422 65494
rect 113186 58258 113422 58494
rect 113186 51258 113422 51494
rect 113186 44258 113422 44494
rect 113186 37258 113422 37494
rect 113186 30258 113422 30494
rect 113186 23258 113422 23494
rect 113186 16258 113422 16494
rect 113186 9258 113422 9494
rect 113186 2258 113422 2494
rect 113186 -982 113422 -746
rect 113186 -1302 113422 -1066
rect 114918 705962 115154 706198
rect 114918 705642 115154 705878
rect 114918 696325 115154 696561
rect 114918 689325 115154 689561
rect 114918 682325 115154 682561
rect 114918 675325 115154 675561
rect 114918 668325 115154 668561
rect 114918 661325 115154 661561
rect 114918 654325 115154 654561
rect 114918 647325 115154 647561
rect 114918 640325 115154 640561
rect 114918 633325 115154 633561
rect 114918 626325 115154 626561
rect 114918 619325 115154 619561
rect 114918 612325 115154 612561
rect 114918 605325 115154 605561
rect 114918 598325 115154 598561
rect 114918 591325 115154 591561
rect 114918 584325 115154 584561
rect 114918 577325 115154 577561
rect 114918 570325 115154 570561
rect 114918 563325 115154 563561
rect 114918 556325 115154 556561
rect 114918 549325 115154 549561
rect 114918 542325 115154 542561
rect 114918 535325 115154 535561
rect 114918 528325 115154 528561
rect 114918 521325 115154 521561
rect 114918 514325 115154 514561
rect 114918 507325 115154 507561
rect 114918 500325 115154 500561
rect 114918 493325 115154 493561
rect 114918 486325 115154 486561
rect 114918 479325 115154 479561
rect 114918 472325 115154 472561
rect 114918 465325 115154 465561
rect 114918 458325 115154 458561
rect 114918 451325 115154 451561
rect 114918 444325 115154 444561
rect 114918 437325 115154 437561
rect 114918 430325 115154 430561
rect 114918 423325 115154 423561
rect 114918 416325 115154 416561
rect 114918 409325 115154 409561
rect 114918 402325 115154 402561
rect 114918 395325 115154 395561
rect 114918 388325 115154 388561
rect 114918 381325 115154 381561
rect 114918 374325 115154 374561
rect 114918 367325 115154 367561
rect 114918 360325 115154 360561
rect 114918 353325 115154 353561
rect 114918 346325 115154 346561
rect 114918 339325 115154 339561
rect 114918 332325 115154 332561
rect 114918 325325 115154 325561
rect 114918 318325 115154 318561
rect 114918 311325 115154 311561
rect 114918 304325 115154 304561
rect 114918 297325 115154 297561
rect 114918 290325 115154 290561
rect 114918 283325 115154 283561
rect 114918 276325 115154 276561
rect 114918 269325 115154 269561
rect 114918 262325 115154 262561
rect 114918 255325 115154 255561
rect 114918 248325 115154 248561
rect 114918 241325 115154 241561
rect 114918 234325 115154 234561
rect 114918 227325 115154 227561
rect 114918 220325 115154 220561
rect 114918 213325 115154 213561
rect 114918 206325 115154 206561
rect 114918 199325 115154 199561
rect 114918 192325 115154 192561
rect 114918 185325 115154 185561
rect 114918 178325 115154 178561
rect 114918 171325 115154 171561
rect 114918 164325 115154 164561
rect 114918 157325 115154 157561
rect 114918 150325 115154 150561
rect 114918 143325 115154 143561
rect 114918 136325 115154 136561
rect 114918 129325 115154 129561
rect 114918 122325 115154 122561
rect 114918 115325 115154 115561
rect 114918 108325 115154 108561
rect 114918 101325 115154 101561
rect 114918 94325 115154 94561
rect 114918 87325 115154 87561
rect 114918 80325 115154 80561
rect 114918 73325 115154 73561
rect 114918 66325 115154 66561
rect 114918 59325 115154 59561
rect 114918 52325 115154 52561
rect 114918 45325 115154 45561
rect 114918 38325 115154 38561
rect 114918 31325 115154 31561
rect 114918 24325 115154 24561
rect 114918 17325 115154 17561
rect 114918 10325 115154 10561
rect 114918 3325 115154 3561
rect 114918 -1942 115154 -1706
rect 114918 -2262 115154 -2026
rect 120186 705002 120422 705238
rect 120186 704682 120422 704918
rect 120186 695258 120422 695494
rect 120186 688258 120422 688494
rect 120186 681258 120422 681494
rect 120186 674258 120422 674494
rect 120186 667258 120422 667494
rect 120186 660258 120422 660494
rect 120186 653258 120422 653494
rect 120186 646258 120422 646494
rect 120186 639258 120422 639494
rect 120186 632258 120422 632494
rect 120186 625258 120422 625494
rect 120186 618258 120422 618494
rect 120186 611258 120422 611494
rect 120186 604258 120422 604494
rect 120186 597258 120422 597494
rect 120186 590258 120422 590494
rect 120186 583258 120422 583494
rect 120186 576258 120422 576494
rect 120186 569258 120422 569494
rect 120186 562258 120422 562494
rect 120186 555258 120422 555494
rect 120186 548258 120422 548494
rect 120186 541258 120422 541494
rect 120186 534258 120422 534494
rect 120186 527258 120422 527494
rect 120186 520258 120422 520494
rect 120186 513258 120422 513494
rect 120186 506258 120422 506494
rect 120186 499258 120422 499494
rect 120186 492258 120422 492494
rect 120186 485258 120422 485494
rect 120186 478258 120422 478494
rect 120186 471258 120422 471494
rect 120186 464258 120422 464494
rect 120186 457258 120422 457494
rect 120186 450258 120422 450494
rect 120186 443258 120422 443494
rect 120186 436258 120422 436494
rect 120186 429258 120422 429494
rect 120186 422258 120422 422494
rect 120186 415258 120422 415494
rect 120186 408258 120422 408494
rect 120186 401258 120422 401494
rect 120186 394258 120422 394494
rect 120186 387258 120422 387494
rect 120186 380258 120422 380494
rect 120186 373258 120422 373494
rect 120186 366258 120422 366494
rect 120186 359258 120422 359494
rect 120186 352258 120422 352494
rect 120186 345258 120422 345494
rect 120186 338258 120422 338494
rect 120186 331258 120422 331494
rect 120186 324258 120422 324494
rect 120186 317258 120422 317494
rect 120186 310258 120422 310494
rect 120186 303258 120422 303494
rect 120186 296258 120422 296494
rect 120186 289258 120422 289494
rect 120186 282258 120422 282494
rect 120186 275258 120422 275494
rect 120186 268258 120422 268494
rect 120186 261258 120422 261494
rect 120186 254258 120422 254494
rect 120186 247258 120422 247494
rect 120186 240258 120422 240494
rect 120186 233258 120422 233494
rect 120186 226258 120422 226494
rect 120186 219258 120422 219494
rect 120186 212258 120422 212494
rect 120186 205258 120422 205494
rect 120186 198258 120422 198494
rect 120186 191258 120422 191494
rect 120186 184258 120422 184494
rect 120186 177258 120422 177494
rect 120186 170258 120422 170494
rect 120186 163258 120422 163494
rect 120186 156258 120422 156494
rect 120186 149258 120422 149494
rect 120186 142258 120422 142494
rect 120186 135258 120422 135494
rect 120186 128258 120422 128494
rect 120186 121258 120422 121494
rect 120186 114258 120422 114494
rect 120186 107258 120422 107494
rect 120186 100258 120422 100494
rect 120186 93258 120422 93494
rect 120186 86258 120422 86494
rect 120186 79258 120422 79494
rect 120186 72258 120422 72494
rect 120186 65258 120422 65494
rect 120186 58258 120422 58494
rect 120186 51258 120422 51494
rect 120186 44258 120422 44494
rect 120186 37258 120422 37494
rect 120186 30258 120422 30494
rect 120186 23258 120422 23494
rect 120186 16258 120422 16494
rect 120186 9258 120422 9494
rect 120186 2258 120422 2494
rect 120186 -982 120422 -746
rect 120186 -1302 120422 -1066
rect 121918 705962 122154 706198
rect 121918 705642 122154 705878
rect 121918 696325 122154 696561
rect 121918 689325 122154 689561
rect 121918 682325 122154 682561
rect 121918 675325 122154 675561
rect 121918 668325 122154 668561
rect 121918 661325 122154 661561
rect 121918 654325 122154 654561
rect 121918 647325 122154 647561
rect 121918 640325 122154 640561
rect 121918 633325 122154 633561
rect 121918 626325 122154 626561
rect 121918 619325 122154 619561
rect 121918 612325 122154 612561
rect 121918 605325 122154 605561
rect 121918 598325 122154 598561
rect 121918 591325 122154 591561
rect 121918 584325 122154 584561
rect 121918 577325 122154 577561
rect 121918 570325 122154 570561
rect 121918 563325 122154 563561
rect 121918 556325 122154 556561
rect 121918 549325 122154 549561
rect 121918 542325 122154 542561
rect 121918 535325 122154 535561
rect 121918 528325 122154 528561
rect 121918 521325 122154 521561
rect 121918 514325 122154 514561
rect 121918 507325 122154 507561
rect 121918 500325 122154 500561
rect 121918 493325 122154 493561
rect 121918 486325 122154 486561
rect 121918 479325 122154 479561
rect 121918 472325 122154 472561
rect 121918 465325 122154 465561
rect 121918 458325 122154 458561
rect 121918 451325 122154 451561
rect 121918 444325 122154 444561
rect 121918 437325 122154 437561
rect 121918 430325 122154 430561
rect 121918 423325 122154 423561
rect 121918 416325 122154 416561
rect 121918 409325 122154 409561
rect 121918 402325 122154 402561
rect 121918 395325 122154 395561
rect 121918 388325 122154 388561
rect 121918 381325 122154 381561
rect 121918 374325 122154 374561
rect 121918 367325 122154 367561
rect 121918 360325 122154 360561
rect 121918 353325 122154 353561
rect 121918 346325 122154 346561
rect 121918 339325 122154 339561
rect 121918 332325 122154 332561
rect 121918 325325 122154 325561
rect 121918 318325 122154 318561
rect 121918 311325 122154 311561
rect 121918 304325 122154 304561
rect 121918 297325 122154 297561
rect 121918 290325 122154 290561
rect 121918 283325 122154 283561
rect 121918 276325 122154 276561
rect 121918 269325 122154 269561
rect 121918 262325 122154 262561
rect 121918 255325 122154 255561
rect 121918 248325 122154 248561
rect 121918 241325 122154 241561
rect 121918 234325 122154 234561
rect 121918 227325 122154 227561
rect 121918 220325 122154 220561
rect 121918 213325 122154 213561
rect 121918 206325 122154 206561
rect 121918 199325 122154 199561
rect 121918 192325 122154 192561
rect 121918 185325 122154 185561
rect 121918 178325 122154 178561
rect 121918 171325 122154 171561
rect 121918 164325 122154 164561
rect 121918 157325 122154 157561
rect 121918 150325 122154 150561
rect 121918 143325 122154 143561
rect 121918 136325 122154 136561
rect 121918 129325 122154 129561
rect 121918 122325 122154 122561
rect 121918 115325 122154 115561
rect 121918 108325 122154 108561
rect 121918 101325 122154 101561
rect 121918 94325 122154 94561
rect 121918 87325 122154 87561
rect 121918 80325 122154 80561
rect 121918 73325 122154 73561
rect 121918 66325 122154 66561
rect 121918 59325 122154 59561
rect 121918 52325 122154 52561
rect 121918 45325 122154 45561
rect 121918 38325 122154 38561
rect 121918 31325 122154 31561
rect 121918 24325 122154 24561
rect 121918 17325 122154 17561
rect 121918 10325 122154 10561
rect 121918 3325 122154 3561
rect 121918 -1942 122154 -1706
rect 121918 -2262 122154 -2026
rect 127186 705002 127422 705238
rect 127186 704682 127422 704918
rect 127186 695258 127422 695494
rect 127186 688258 127422 688494
rect 127186 681258 127422 681494
rect 127186 674258 127422 674494
rect 127186 667258 127422 667494
rect 127186 660258 127422 660494
rect 127186 653258 127422 653494
rect 127186 646258 127422 646494
rect 127186 639258 127422 639494
rect 127186 632258 127422 632494
rect 127186 625258 127422 625494
rect 127186 618258 127422 618494
rect 127186 611258 127422 611494
rect 127186 604258 127422 604494
rect 127186 597258 127422 597494
rect 127186 590258 127422 590494
rect 127186 583258 127422 583494
rect 127186 576258 127422 576494
rect 127186 569258 127422 569494
rect 127186 562258 127422 562494
rect 127186 555258 127422 555494
rect 127186 548258 127422 548494
rect 127186 541258 127422 541494
rect 127186 534258 127422 534494
rect 127186 527258 127422 527494
rect 127186 520258 127422 520494
rect 127186 513258 127422 513494
rect 127186 506258 127422 506494
rect 127186 499258 127422 499494
rect 127186 492258 127422 492494
rect 127186 485258 127422 485494
rect 127186 478258 127422 478494
rect 127186 471258 127422 471494
rect 127186 464258 127422 464494
rect 127186 457258 127422 457494
rect 127186 450258 127422 450494
rect 127186 443258 127422 443494
rect 127186 436258 127422 436494
rect 127186 429258 127422 429494
rect 127186 422258 127422 422494
rect 127186 415258 127422 415494
rect 127186 408258 127422 408494
rect 127186 401258 127422 401494
rect 127186 394258 127422 394494
rect 127186 387258 127422 387494
rect 127186 380258 127422 380494
rect 127186 373258 127422 373494
rect 127186 366258 127422 366494
rect 127186 359258 127422 359494
rect 127186 352258 127422 352494
rect 127186 345258 127422 345494
rect 127186 338258 127422 338494
rect 127186 331258 127422 331494
rect 127186 324258 127422 324494
rect 127186 317258 127422 317494
rect 127186 310258 127422 310494
rect 127186 303258 127422 303494
rect 127186 296258 127422 296494
rect 127186 289258 127422 289494
rect 127186 282258 127422 282494
rect 127186 275258 127422 275494
rect 127186 268258 127422 268494
rect 127186 261258 127422 261494
rect 127186 254258 127422 254494
rect 127186 247258 127422 247494
rect 127186 240258 127422 240494
rect 127186 233258 127422 233494
rect 127186 226258 127422 226494
rect 127186 219258 127422 219494
rect 127186 212258 127422 212494
rect 127186 205258 127422 205494
rect 127186 198258 127422 198494
rect 127186 191258 127422 191494
rect 127186 184258 127422 184494
rect 127186 177258 127422 177494
rect 127186 170258 127422 170494
rect 127186 163258 127422 163494
rect 127186 156258 127422 156494
rect 127186 149258 127422 149494
rect 127186 142258 127422 142494
rect 127186 135258 127422 135494
rect 127186 128258 127422 128494
rect 127186 121258 127422 121494
rect 127186 114258 127422 114494
rect 127186 107258 127422 107494
rect 127186 100258 127422 100494
rect 127186 93258 127422 93494
rect 127186 86258 127422 86494
rect 127186 79258 127422 79494
rect 127186 72258 127422 72494
rect 127186 65258 127422 65494
rect 127186 58258 127422 58494
rect 127186 51258 127422 51494
rect 127186 44258 127422 44494
rect 127186 37258 127422 37494
rect 127186 30258 127422 30494
rect 127186 23258 127422 23494
rect 127186 16258 127422 16494
rect 127186 9258 127422 9494
rect 127186 2258 127422 2494
rect 127186 -982 127422 -746
rect 127186 -1302 127422 -1066
rect 128918 705962 129154 706198
rect 128918 705642 129154 705878
rect 128918 696325 129154 696561
rect 128918 689325 129154 689561
rect 128918 682325 129154 682561
rect 128918 675325 129154 675561
rect 128918 668325 129154 668561
rect 128918 661325 129154 661561
rect 128918 654325 129154 654561
rect 128918 647325 129154 647561
rect 128918 640325 129154 640561
rect 128918 633325 129154 633561
rect 128918 626325 129154 626561
rect 128918 619325 129154 619561
rect 128918 612325 129154 612561
rect 128918 605325 129154 605561
rect 128918 598325 129154 598561
rect 128918 591325 129154 591561
rect 128918 584325 129154 584561
rect 128918 577325 129154 577561
rect 128918 570325 129154 570561
rect 128918 563325 129154 563561
rect 128918 556325 129154 556561
rect 128918 549325 129154 549561
rect 128918 542325 129154 542561
rect 128918 535325 129154 535561
rect 128918 528325 129154 528561
rect 128918 521325 129154 521561
rect 128918 514325 129154 514561
rect 128918 507325 129154 507561
rect 128918 500325 129154 500561
rect 128918 493325 129154 493561
rect 128918 486325 129154 486561
rect 128918 479325 129154 479561
rect 128918 472325 129154 472561
rect 128918 465325 129154 465561
rect 128918 458325 129154 458561
rect 128918 451325 129154 451561
rect 128918 444325 129154 444561
rect 128918 437325 129154 437561
rect 128918 430325 129154 430561
rect 128918 423325 129154 423561
rect 128918 416325 129154 416561
rect 128918 409325 129154 409561
rect 128918 402325 129154 402561
rect 128918 395325 129154 395561
rect 128918 388325 129154 388561
rect 128918 381325 129154 381561
rect 128918 374325 129154 374561
rect 128918 367325 129154 367561
rect 128918 360325 129154 360561
rect 128918 353325 129154 353561
rect 128918 346325 129154 346561
rect 128918 339325 129154 339561
rect 128918 332325 129154 332561
rect 128918 325325 129154 325561
rect 128918 318325 129154 318561
rect 128918 311325 129154 311561
rect 128918 304325 129154 304561
rect 128918 297325 129154 297561
rect 128918 290325 129154 290561
rect 128918 283325 129154 283561
rect 128918 276325 129154 276561
rect 128918 269325 129154 269561
rect 128918 262325 129154 262561
rect 128918 255325 129154 255561
rect 128918 248325 129154 248561
rect 128918 241325 129154 241561
rect 128918 234325 129154 234561
rect 128918 227325 129154 227561
rect 128918 220325 129154 220561
rect 128918 213325 129154 213561
rect 128918 206325 129154 206561
rect 128918 199325 129154 199561
rect 128918 192325 129154 192561
rect 128918 185325 129154 185561
rect 128918 178325 129154 178561
rect 128918 171325 129154 171561
rect 128918 164325 129154 164561
rect 128918 157325 129154 157561
rect 128918 150325 129154 150561
rect 128918 143325 129154 143561
rect 128918 136325 129154 136561
rect 128918 129325 129154 129561
rect 128918 122325 129154 122561
rect 128918 115325 129154 115561
rect 128918 108325 129154 108561
rect 128918 101325 129154 101561
rect 128918 94325 129154 94561
rect 128918 87325 129154 87561
rect 128918 80325 129154 80561
rect 128918 73325 129154 73561
rect 128918 66325 129154 66561
rect 128918 59325 129154 59561
rect 128918 52325 129154 52561
rect 128918 45325 129154 45561
rect 128918 38325 129154 38561
rect 128918 31325 129154 31561
rect 128918 24325 129154 24561
rect 128918 17325 129154 17561
rect 128918 10325 129154 10561
rect 128918 3325 129154 3561
rect 128918 -1942 129154 -1706
rect 128918 -2262 129154 -2026
rect 134186 705002 134422 705238
rect 134186 704682 134422 704918
rect 134186 695258 134422 695494
rect 134186 688258 134422 688494
rect 134186 681258 134422 681494
rect 134186 674258 134422 674494
rect 134186 667258 134422 667494
rect 134186 660258 134422 660494
rect 134186 653258 134422 653494
rect 134186 646258 134422 646494
rect 134186 639258 134422 639494
rect 134186 632258 134422 632494
rect 134186 625258 134422 625494
rect 134186 618258 134422 618494
rect 134186 611258 134422 611494
rect 134186 604258 134422 604494
rect 134186 597258 134422 597494
rect 134186 590258 134422 590494
rect 134186 583258 134422 583494
rect 134186 576258 134422 576494
rect 134186 569258 134422 569494
rect 134186 562258 134422 562494
rect 134186 555258 134422 555494
rect 134186 548258 134422 548494
rect 134186 541258 134422 541494
rect 134186 534258 134422 534494
rect 134186 527258 134422 527494
rect 134186 520258 134422 520494
rect 134186 513258 134422 513494
rect 134186 506258 134422 506494
rect 134186 499258 134422 499494
rect 134186 492258 134422 492494
rect 134186 485258 134422 485494
rect 134186 478258 134422 478494
rect 134186 471258 134422 471494
rect 134186 464258 134422 464494
rect 134186 457258 134422 457494
rect 134186 450258 134422 450494
rect 134186 443258 134422 443494
rect 134186 436258 134422 436494
rect 134186 429258 134422 429494
rect 134186 422258 134422 422494
rect 134186 415258 134422 415494
rect 134186 408258 134422 408494
rect 134186 401258 134422 401494
rect 134186 394258 134422 394494
rect 134186 387258 134422 387494
rect 134186 380258 134422 380494
rect 134186 373258 134422 373494
rect 134186 366258 134422 366494
rect 134186 359258 134422 359494
rect 134186 352258 134422 352494
rect 134186 345258 134422 345494
rect 134186 338258 134422 338494
rect 134186 331258 134422 331494
rect 134186 324258 134422 324494
rect 134186 317258 134422 317494
rect 134186 310258 134422 310494
rect 134186 303258 134422 303494
rect 134186 296258 134422 296494
rect 134186 289258 134422 289494
rect 134186 282258 134422 282494
rect 134186 275258 134422 275494
rect 134186 268258 134422 268494
rect 134186 261258 134422 261494
rect 134186 254258 134422 254494
rect 134186 247258 134422 247494
rect 134186 240258 134422 240494
rect 134186 233258 134422 233494
rect 134186 226258 134422 226494
rect 134186 219258 134422 219494
rect 134186 212258 134422 212494
rect 134186 205258 134422 205494
rect 134186 198258 134422 198494
rect 134186 191258 134422 191494
rect 134186 184258 134422 184494
rect 134186 177258 134422 177494
rect 134186 170258 134422 170494
rect 134186 163258 134422 163494
rect 134186 156258 134422 156494
rect 134186 149258 134422 149494
rect 134186 142258 134422 142494
rect 134186 135258 134422 135494
rect 134186 128258 134422 128494
rect 134186 121258 134422 121494
rect 134186 114258 134422 114494
rect 134186 107258 134422 107494
rect 134186 100258 134422 100494
rect 134186 93258 134422 93494
rect 134186 86258 134422 86494
rect 134186 79258 134422 79494
rect 134186 72258 134422 72494
rect 134186 65258 134422 65494
rect 134186 58258 134422 58494
rect 134186 51258 134422 51494
rect 134186 44258 134422 44494
rect 134186 37258 134422 37494
rect 134186 30258 134422 30494
rect 134186 23258 134422 23494
rect 134186 16258 134422 16494
rect 134186 9258 134422 9494
rect 134186 2258 134422 2494
rect 134186 -982 134422 -746
rect 134186 -1302 134422 -1066
rect 135918 705962 136154 706198
rect 135918 705642 136154 705878
rect 135918 696325 136154 696561
rect 135918 689325 136154 689561
rect 135918 682325 136154 682561
rect 135918 675325 136154 675561
rect 135918 668325 136154 668561
rect 135918 661325 136154 661561
rect 135918 654325 136154 654561
rect 135918 647325 136154 647561
rect 135918 640325 136154 640561
rect 135918 633325 136154 633561
rect 135918 626325 136154 626561
rect 135918 619325 136154 619561
rect 135918 612325 136154 612561
rect 135918 605325 136154 605561
rect 135918 598325 136154 598561
rect 135918 591325 136154 591561
rect 135918 584325 136154 584561
rect 135918 577325 136154 577561
rect 135918 570325 136154 570561
rect 135918 563325 136154 563561
rect 135918 556325 136154 556561
rect 135918 549325 136154 549561
rect 135918 542325 136154 542561
rect 135918 535325 136154 535561
rect 135918 528325 136154 528561
rect 135918 521325 136154 521561
rect 135918 514325 136154 514561
rect 135918 507325 136154 507561
rect 135918 500325 136154 500561
rect 135918 493325 136154 493561
rect 135918 486325 136154 486561
rect 135918 479325 136154 479561
rect 135918 472325 136154 472561
rect 135918 465325 136154 465561
rect 135918 458325 136154 458561
rect 135918 451325 136154 451561
rect 135918 444325 136154 444561
rect 135918 437325 136154 437561
rect 135918 430325 136154 430561
rect 135918 423325 136154 423561
rect 135918 416325 136154 416561
rect 135918 409325 136154 409561
rect 135918 402325 136154 402561
rect 135918 395325 136154 395561
rect 135918 388325 136154 388561
rect 135918 381325 136154 381561
rect 135918 374325 136154 374561
rect 135918 367325 136154 367561
rect 135918 360325 136154 360561
rect 135918 353325 136154 353561
rect 135918 346325 136154 346561
rect 135918 339325 136154 339561
rect 135918 332325 136154 332561
rect 135918 325325 136154 325561
rect 135918 318325 136154 318561
rect 135918 311325 136154 311561
rect 135918 304325 136154 304561
rect 135918 297325 136154 297561
rect 135918 290325 136154 290561
rect 135918 283325 136154 283561
rect 135918 276325 136154 276561
rect 135918 269325 136154 269561
rect 135918 262325 136154 262561
rect 135918 255325 136154 255561
rect 135918 248325 136154 248561
rect 135918 241325 136154 241561
rect 135918 234325 136154 234561
rect 135918 227325 136154 227561
rect 135918 220325 136154 220561
rect 135918 213325 136154 213561
rect 135918 206325 136154 206561
rect 135918 199325 136154 199561
rect 135918 192325 136154 192561
rect 135918 185325 136154 185561
rect 135918 178325 136154 178561
rect 135918 171325 136154 171561
rect 135918 164325 136154 164561
rect 135918 157325 136154 157561
rect 135918 150325 136154 150561
rect 135918 143325 136154 143561
rect 135918 136325 136154 136561
rect 135918 129325 136154 129561
rect 135918 122325 136154 122561
rect 135918 115325 136154 115561
rect 135918 108325 136154 108561
rect 135918 101325 136154 101561
rect 135918 94325 136154 94561
rect 135918 87325 136154 87561
rect 135918 80325 136154 80561
rect 135918 73325 136154 73561
rect 135918 66325 136154 66561
rect 135918 59325 136154 59561
rect 135918 52325 136154 52561
rect 135918 45325 136154 45561
rect 135918 38325 136154 38561
rect 135918 31325 136154 31561
rect 135918 24325 136154 24561
rect 135918 17325 136154 17561
rect 135918 10325 136154 10561
rect 135918 3325 136154 3561
rect 135918 -1942 136154 -1706
rect 135918 -2262 136154 -2026
rect 141186 705002 141422 705238
rect 141186 704682 141422 704918
rect 141186 695258 141422 695494
rect 141186 688258 141422 688494
rect 141186 681258 141422 681494
rect 141186 674258 141422 674494
rect 141186 667258 141422 667494
rect 141186 660258 141422 660494
rect 141186 653258 141422 653494
rect 141186 646258 141422 646494
rect 141186 639258 141422 639494
rect 141186 632258 141422 632494
rect 141186 625258 141422 625494
rect 141186 618258 141422 618494
rect 141186 611258 141422 611494
rect 141186 604258 141422 604494
rect 141186 597258 141422 597494
rect 141186 590258 141422 590494
rect 141186 583258 141422 583494
rect 141186 576258 141422 576494
rect 141186 569258 141422 569494
rect 141186 562258 141422 562494
rect 141186 555258 141422 555494
rect 141186 548258 141422 548494
rect 141186 541258 141422 541494
rect 141186 534258 141422 534494
rect 141186 527258 141422 527494
rect 141186 520258 141422 520494
rect 141186 513258 141422 513494
rect 141186 506258 141422 506494
rect 141186 499258 141422 499494
rect 141186 492258 141422 492494
rect 141186 485258 141422 485494
rect 141186 478258 141422 478494
rect 141186 471258 141422 471494
rect 141186 464258 141422 464494
rect 141186 457258 141422 457494
rect 141186 450258 141422 450494
rect 141186 443258 141422 443494
rect 141186 436258 141422 436494
rect 141186 429258 141422 429494
rect 141186 422258 141422 422494
rect 141186 415258 141422 415494
rect 141186 408258 141422 408494
rect 141186 401258 141422 401494
rect 141186 394258 141422 394494
rect 141186 387258 141422 387494
rect 141186 380258 141422 380494
rect 141186 373258 141422 373494
rect 141186 366258 141422 366494
rect 141186 359258 141422 359494
rect 141186 352258 141422 352494
rect 141186 345258 141422 345494
rect 141186 338258 141422 338494
rect 141186 331258 141422 331494
rect 141186 324258 141422 324494
rect 141186 317258 141422 317494
rect 141186 310258 141422 310494
rect 141186 303258 141422 303494
rect 141186 296258 141422 296494
rect 141186 289258 141422 289494
rect 141186 282258 141422 282494
rect 141186 275258 141422 275494
rect 141186 268258 141422 268494
rect 141186 261258 141422 261494
rect 141186 254258 141422 254494
rect 141186 247258 141422 247494
rect 141186 240258 141422 240494
rect 141186 233258 141422 233494
rect 141186 226258 141422 226494
rect 141186 219258 141422 219494
rect 141186 212258 141422 212494
rect 141186 205258 141422 205494
rect 141186 198258 141422 198494
rect 141186 191258 141422 191494
rect 141186 184258 141422 184494
rect 141186 177258 141422 177494
rect 141186 170258 141422 170494
rect 141186 163258 141422 163494
rect 141186 156258 141422 156494
rect 141186 149258 141422 149494
rect 141186 142258 141422 142494
rect 141186 135258 141422 135494
rect 141186 128258 141422 128494
rect 141186 121258 141422 121494
rect 141186 114258 141422 114494
rect 141186 107258 141422 107494
rect 141186 100258 141422 100494
rect 141186 93258 141422 93494
rect 141186 86258 141422 86494
rect 141186 79258 141422 79494
rect 141186 72258 141422 72494
rect 141186 65258 141422 65494
rect 141186 58258 141422 58494
rect 141186 51258 141422 51494
rect 141186 44258 141422 44494
rect 141186 37258 141422 37494
rect 141186 30258 141422 30494
rect 141186 23258 141422 23494
rect 141186 16258 141422 16494
rect 141186 9258 141422 9494
rect 141186 2258 141422 2494
rect 141186 -982 141422 -746
rect 141186 -1302 141422 -1066
rect 142918 705962 143154 706198
rect 142918 705642 143154 705878
rect 142918 696325 143154 696561
rect 142918 689325 143154 689561
rect 142918 682325 143154 682561
rect 142918 675325 143154 675561
rect 142918 668325 143154 668561
rect 142918 661325 143154 661561
rect 142918 654325 143154 654561
rect 142918 647325 143154 647561
rect 142918 640325 143154 640561
rect 142918 633325 143154 633561
rect 142918 626325 143154 626561
rect 142918 619325 143154 619561
rect 142918 612325 143154 612561
rect 142918 605325 143154 605561
rect 142918 598325 143154 598561
rect 142918 591325 143154 591561
rect 142918 584325 143154 584561
rect 142918 577325 143154 577561
rect 142918 570325 143154 570561
rect 142918 563325 143154 563561
rect 142918 556325 143154 556561
rect 142918 549325 143154 549561
rect 142918 542325 143154 542561
rect 142918 535325 143154 535561
rect 142918 528325 143154 528561
rect 142918 521325 143154 521561
rect 142918 514325 143154 514561
rect 142918 507325 143154 507561
rect 142918 500325 143154 500561
rect 142918 493325 143154 493561
rect 142918 486325 143154 486561
rect 142918 479325 143154 479561
rect 142918 472325 143154 472561
rect 142918 465325 143154 465561
rect 142918 458325 143154 458561
rect 142918 451325 143154 451561
rect 142918 444325 143154 444561
rect 142918 437325 143154 437561
rect 142918 430325 143154 430561
rect 142918 423325 143154 423561
rect 142918 416325 143154 416561
rect 142918 409325 143154 409561
rect 142918 402325 143154 402561
rect 142918 395325 143154 395561
rect 142918 388325 143154 388561
rect 142918 381325 143154 381561
rect 142918 374325 143154 374561
rect 142918 367325 143154 367561
rect 142918 360325 143154 360561
rect 142918 353325 143154 353561
rect 142918 346325 143154 346561
rect 142918 339325 143154 339561
rect 142918 332325 143154 332561
rect 142918 325325 143154 325561
rect 142918 318325 143154 318561
rect 142918 311325 143154 311561
rect 142918 304325 143154 304561
rect 142918 297325 143154 297561
rect 142918 290325 143154 290561
rect 142918 283325 143154 283561
rect 142918 276325 143154 276561
rect 142918 269325 143154 269561
rect 142918 262325 143154 262561
rect 142918 255325 143154 255561
rect 142918 248325 143154 248561
rect 142918 241325 143154 241561
rect 142918 234325 143154 234561
rect 142918 227325 143154 227561
rect 142918 220325 143154 220561
rect 142918 213325 143154 213561
rect 142918 206325 143154 206561
rect 142918 199325 143154 199561
rect 142918 192325 143154 192561
rect 142918 185325 143154 185561
rect 142918 178325 143154 178561
rect 142918 171325 143154 171561
rect 142918 164325 143154 164561
rect 142918 157325 143154 157561
rect 142918 150325 143154 150561
rect 142918 143325 143154 143561
rect 142918 136325 143154 136561
rect 142918 129325 143154 129561
rect 142918 122325 143154 122561
rect 142918 115325 143154 115561
rect 142918 108325 143154 108561
rect 142918 101325 143154 101561
rect 142918 94325 143154 94561
rect 142918 87325 143154 87561
rect 142918 80325 143154 80561
rect 142918 73325 143154 73561
rect 142918 66325 143154 66561
rect 142918 59325 143154 59561
rect 142918 52325 143154 52561
rect 142918 45325 143154 45561
rect 142918 38325 143154 38561
rect 142918 31325 143154 31561
rect 142918 24325 143154 24561
rect 142918 17325 143154 17561
rect 142918 10325 143154 10561
rect 142918 3325 143154 3561
rect 142918 -1942 143154 -1706
rect 142918 -2262 143154 -2026
rect 148186 705002 148422 705238
rect 148186 704682 148422 704918
rect 148186 695258 148422 695494
rect 148186 688258 148422 688494
rect 148186 681258 148422 681494
rect 148186 674258 148422 674494
rect 148186 667258 148422 667494
rect 148186 660258 148422 660494
rect 148186 653258 148422 653494
rect 148186 646258 148422 646494
rect 148186 639258 148422 639494
rect 148186 632258 148422 632494
rect 148186 625258 148422 625494
rect 148186 618258 148422 618494
rect 148186 611258 148422 611494
rect 148186 604258 148422 604494
rect 148186 597258 148422 597494
rect 148186 590258 148422 590494
rect 148186 583258 148422 583494
rect 148186 576258 148422 576494
rect 148186 569258 148422 569494
rect 148186 562258 148422 562494
rect 148186 555258 148422 555494
rect 148186 548258 148422 548494
rect 148186 541258 148422 541494
rect 148186 534258 148422 534494
rect 148186 527258 148422 527494
rect 148186 520258 148422 520494
rect 148186 513258 148422 513494
rect 148186 506258 148422 506494
rect 148186 499258 148422 499494
rect 148186 492258 148422 492494
rect 148186 485258 148422 485494
rect 148186 478258 148422 478494
rect 148186 471258 148422 471494
rect 148186 464258 148422 464494
rect 148186 457258 148422 457494
rect 148186 450258 148422 450494
rect 148186 443258 148422 443494
rect 148186 436258 148422 436494
rect 148186 429258 148422 429494
rect 148186 422258 148422 422494
rect 148186 415258 148422 415494
rect 148186 408258 148422 408494
rect 148186 401258 148422 401494
rect 148186 394258 148422 394494
rect 148186 387258 148422 387494
rect 148186 380258 148422 380494
rect 148186 373258 148422 373494
rect 148186 366258 148422 366494
rect 148186 359258 148422 359494
rect 148186 352258 148422 352494
rect 148186 345258 148422 345494
rect 148186 338258 148422 338494
rect 148186 331258 148422 331494
rect 148186 324258 148422 324494
rect 148186 317258 148422 317494
rect 148186 310258 148422 310494
rect 148186 303258 148422 303494
rect 148186 296258 148422 296494
rect 148186 289258 148422 289494
rect 148186 282258 148422 282494
rect 148186 275258 148422 275494
rect 148186 268258 148422 268494
rect 148186 261258 148422 261494
rect 148186 254258 148422 254494
rect 148186 247258 148422 247494
rect 148186 240258 148422 240494
rect 148186 233258 148422 233494
rect 148186 226258 148422 226494
rect 148186 219258 148422 219494
rect 148186 212258 148422 212494
rect 148186 205258 148422 205494
rect 148186 198258 148422 198494
rect 148186 191258 148422 191494
rect 148186 184258 148422 184494
rect 148186 177258 148422 177494
rect 148186 170258 148422 170494
rect 148186 163258 148422 163494
rect 148186 156258 148422 156494
rect 148186 149258 148422 149494
rect 148186 142258 148422 142494
rect 148186 135258 148422 135494
rect 148186 128258 148422 128494
rect 148186 121258 148422 121494
rect 148186 114258 148422 114494
rect 148186 107258 148422 107494
rect 148186 100258 148422 100494
rect 148186 93258 148422 93494
rect 148186 86258 148422 86494
rect 148186 79258 148422 79494
rect 148186 72258 148422 72494
rect 148186 65258 148422 65494
rect 148186 58258 148422 58494
rect 148186 51258 148422 51494
rect 148186 44258 148422 44494
rect 148186 37258 148422 37494
rect 148186 30258 148422 30494
rect 148186 23258 148422 23494
rect 148186 16258 148422 16494
rect 148186 9258 148422 9494
rect 148186 2258 148422 2494
rect 148186 -982 148422 -746
rect 148186 -1302 148422 -1066
rect 149918 705962 150154 706198
rect 149918 705642 150154 705878
rect 149918 696325 150154 696561
rect 149918 689325 150154 689561
rect 149918 682325 150154 682561
rect 149918 675325 150154 675561
rect 149918 668325 150154 668561
rect 149918 661325 150154 661561
rect 149918 654325 150154 654561
rect 149918 647325 150154 647561
rect 149918 640325 150154 640561
rect 149918 633325 150154 633561
rect 149918 626325 150154 626561
rect 149918 619325 150154 619561
rect 149918 612325 150154 612561
rect 149918 605325 150154 605561
rect 149918 598325 150154 598561
rect 149918 591325 150154 591561
rect 149918 584325 150154 584561
rect 149918 577325 150154 577561
rect 149918 570325 150154 570561
rect 149918 563325 150154 563561
rect 149918 556325 150154 556561
rect 149918 549325 150154 549561
rect 149918 542325 150154 542561
rect 149918 535325 150154 535561
rect 149918 528325 150154 528561
rect 149918 521325 150154 521561
rect 149918 514325 150154 514561
rect 149918 507325 150154 507561
rect 149918 500325 150154 500561
rect 149918 493325 150154 493561
rect 149918 486325 150154 486561
rect 149918 479325 150154 479561
rect 149918 472325 150154 472561
rect 149918 465325 150154 465561
rect 149918 458325 150154 458561
rect 149918 451325 150154 451561
rect 149918 444325 150154 444561
rect 149918 437325 150154 437561
rect 149918 430325 150154 430561
rect 149918 423325 150154 423561
rect 149918 416325 150154 416561
rect 149918 409325 150154 409561
rect 149918 402325 150154 402561
rect 149918 395325 150154 395561
rect 149918 388325 150154 388561
rect 149918 381325 150154 381561
rect 149918 374325 150154 374561
rect 149918 367325 150154 367561
rect 149918 360325 150154 360561
rect 149918 353325 150154 353561
rect 149918 346325 150154 346561
rect 149918 339325 150154 339561
rect 149918 332325 150154 332561
rect 149918 325325 150154 325561
rect 149918 318325 150154 318561
rect 149918 311325 150154 311561
rect 149918 304325 150154 304561
rect 149918 297325 150154 297561
rect 149918 290325 150154 290561
rect 149918 283325 150154 283561
rect 149918 276325 150154 276561
rect 149918 269325 150154 269561
rect 149918 262325 150154 262561
rect 149918 255325 150154 255561
rect 149918 248325 150154 248561
rect 149918 241325 150154 241561
rect 149918 234325 150154 234561
rect 149918 227325 150154 227561
rect 149918 220325 150154 220561
rect 149918 213325 150154 213561
rect 149918 206325 150154 206561
rect 149918 199325 150154 199561
rect 149918 192325 150154 192561
rect 149918 185325 150154 185561
rect 149918 178325 150154 178561
rect 149918 171325 150154 171561
rect 149918 164325 150154 164561
rect 149918 157325 150154 157561
rect 149918 150325 150154 150561
rect 149918 143325 150154 143561
rect 149918 136325 150154 136561
rect 149918 129325 150154 129561
rect 149918 122325 150154 122561
rect 149918 115325 150154 115561
rect 149918 108325 150154 108561
rect 149918 101325 150154 101561
rect 149918 94325 150154 94561
rect 149918 87325 150154 87561
rect 149918 80325 150154 80561
rect 149918 73325 150154 73561
rect 149918 66325 150154 66561
rect 149918 59325 150154 59561
rect 149918 52325 150154 52561
rect 149918 45325 150154 45561
rect 149918 38325 150154 38561
rect 149918 31325 150154 31561
rect 149918 24325 150154 24561
rect 149918 17325 150154 17561
rect 149918 10325 150154 10561
rect 149918 3325 150154 3561
rect 149918 -1942 150154 -1706
rect 149918 -2262 150154 -2026
rect 155186 705002 155422 705238
rect 155186 704682 155422 704918
rect 155186 695258 155422 695494
rect 155186 688258 155422 688494
rect 155186 681258 155422 681494
rect 155186 674258 155422 674494
rect 155186 667258 155422 667494
rect 155186 660258 155422 660494
rect 155186 653258 155422 653494
rect 155186 646258 155422 646494
rect 155186 639258 155422 639494
rect 155186 632258 155422 632494
rect 155186 625258 155422 625494
rect 155186 618258 155422 618494
rect 155186 611258 155422 611494
rect 155186 604258 155422 604494
rect 155186 597258 155422 597494
rect 155186 590258 155422 590494
rect 155186 583258 155422 583494
rect 155186 576258 155422 576494
rect 155186 569258 155422 569494
rect 155186 562258 155422 562494
rect 155186 555258 155422 555494
rect 155186 548258 155422 548494
rect 155186 541258 155422 541494
rect 155186 534258 155422 534494
rect 155186 527258 155422 527494
rect 155186 520258 155422 520494
rect 155186 513258 155422 513494
rect 155186 506258 155422 506494
rect 155186 499258 155422 499494
rect 155186 492258 155422 492494
rect 155186 485258 155422 485494
rect 155186 478258 155422 478494
rect 155186 471258 155422 471494
rect 155186 464258 155422 464494
rect 155186 457258 155422 457494
rect 155186 450258 155422 450494
rect 155186 443258 155422 443494
rect 155186 436258 155422 436494
rect 155186 429258 155422 429494
rect 155186 422258 155422 422494
rect 155186 415258 155422 415494
rect 155186 408258 155422 408494
rect 155186 401258 155422 401494
rect 155186 394258 155422 394494
rect 155186 387258 155422 387494
rect 155186 380258 155422 380494
rect 155186 373258 155422 373494
rect 155186 366258 155422 366494
rect 155186 359258 155422 359494
rect 155186 352258 155422 352494
rect 155186 345258 155422 345494
rect 155186 338258 155422 338494
rect 155186 331258 155422 331494
rect 155186 324258 155422 324494
rect 155186 317258 155422 317494
rect 155186 310258 155422 310494
rect 155186 303258 155422 303494
rect 155186 296258 155422 296494
rect 155186 289258 155422 289494
rect 155186 282258 155422 282494
rect 155186 275258 155422 275494
rect 155186 268258 155422 268494
rect 155186 261258 155422 261494
rect 155186 254258 155422 254494
rect 155186 247258 155422 247494
rect 155186 240258 155422 240494
rect 155186 233258 155422 233494
rect 155186 226258 155422 226494
rect 155186 219258 155422 219494
rect 155186 212258 155422 212494
rect 155186 205258 155422 205494
rect 155186 198258 155422 198494
rect 155186 191258 155422 191494
rect 155186 184258 155422 184494
rect 155186 177258 155422 177494
rect 155186 170258 155422 170494
rect 155186 163258 155422 163494
rect 155186 156258 155422 156494
rect 155186 149258 155422 149494
rect 155186 142258 155422 142494
rect 155186 135258 155422 135494
rect 155186 128258 155422 128494
rect 155186 121258 155422 121494
rect 155186 114258 155422 114494
rect 155186 107258 155422 107494
rect 155186 100258 155422 100494
rect 155186 93258 155422 93494
rect 155186 86258 155422 86494
rect 155186 79258 155422 79494
rect 155186 72258 155422 72494
rect 155186 65258 155422 65494
rect 155186 58258 155422 58494
rect 155186 51258 155422 51494
rect 155186 44258 155422 44494
rect 155186 37258 155422 37494
rect 155186 30258 155422 30494
rect 155186 23258 155422 23494
rect 155186 16258 155422 16494
rect 155186 9258 155422 9494
rect 155186 2258 155422 2494
rect 155186 -982 155422 -746
rect 155186 -1302 155422 -1066
rect 156918 705962 157154 706198
rect 156918 705642 157154 705878
rect 156918 696325 157154 696561
rect 156918 689325 157154 689561
rect 156918 682325 157154 682561
rect 156918 675325 157154 675561
rect 156918 668325 157154 668561
rect 156918 661325 157154 661561
rect 156918 654325 157154 654561
rect 156918 647325 157154 647561
rect 156918 640325 157154 640561
rect 156918 633325 157154 633561
rect 156918 626325 157154 626561
rect 156918 619325 157154 619561
rect 156918 612325 157154 612561
rect 156918 605325 157154 605561
rect 156918 598325 157154 598561
rect 156918 591325 157154 591561
rect 156918 584325 157154 584561
rect 156918 577325 157154 577561
rect 156918 570325 157154 570561
rect 156918 563325 157154 563561
rect 156918 556325 157154 556561
rect 156918 549325 157154 549561
rect 156918 542325 157154 542561
rect 156918 535325 157154 535561
rect 156918 528325 157154 528561
rect 156918 521325 157154 521561
rect 156918 514325 157154 514561
rect 156918 507325 157154 507561
rect 156918 500325 157154 500561
rect 156918 493325 157154 493561
rect 156918 486325 157154 486561
rect 156918 479325 157154 479561
rect 156918 472325 157154 472561
rect 156918 465325 157154 465561
rect 156918 458325 157154 458561
rect 156918 451325 157154 451561
rect 156918 444325 157154 444561
rect 156918 437325 157154 437561
rect 156918 430325 157154 430561
rect 156918 423325 157154 423561
rect 156918 416325 157154 416561
rect 156918 409325 157154 409561
rect 156918 402325 157154 402561
rect 156918 395325 157154 395561
rect 156918 388325 157154 388561
rect 156918 381325 157154 381561
rect 156918 374325 157154 374561
rect 156918 367325 157154 367561
rect 156918 360325 157154 360561
rect 156918 353325 157154 353561
rect 156918 346325 157154 346561
rect 156918 339325 157154 339561
rect 156918 332325 157154 332561
rect 156918 325325 157154 325561
rect 156918 318325 157154 318561
rect 156918 311325 157154 311561
rect 156918 304325 157154 304561
rect 156918 297325 157154 297561
rect 156918 290325 157154 290561
rect 156918 283325 157154 283561
rect 156918 276325 157154 276561
rect 156918 269325 157154 269561
rect 156918 262325 157154 262561
rect 156918 255325 157154 255561
rect 156918 248325 157154 248561
rect 156918 241325 157154 241561
rect 156918 234325 157154 234561
rect 156918 227325 157154 227561
rect 156918 220325 157154 220561
rect 156918 213325 157154 213561
rect 156918 206325 157154 206561
rect 156918 199325 157154 199561
rect 156918 192325 157154 192561
rect 156918 185325 157154 185561
rect 156918 178325 157154 178561
rect 156918 171325 157154 171561
rect 156918 164325 157154 164561
rect 156918 157325 157154 157561
rect 156918 150325 157154 150561
rect 156918 143325 157154 143561
rect 156918 136325 157154 136561
rect 156918 129325 157154 129561
rect 156918 122325 157154 122561
rect 156918 115325 157154 115561
rect 156918 108325 157154 108561
rect 156918 101325 157154 101561
rect 156918 94325 157154 94561
rect 156918 87325 157154 87561
rect 156918 80325 157154 80561
rect 156918 73325 157154 73561
rect 156918 66325 157154 66561
rect 156918 59325 157154 59561
rect 156918 52325 157154 52561
rect 156918 45325 157154 45561
rect 156918 38325 157154 38561
rect 156918 31325 157154 31561
rect 156918 24325 157154 24561
rect 156918 17325 157154 17561
rect 156918 10325 157154 10561
rect 156918 3325 157154 3561
rect 156918 -1942 157154 -1706
rect 156918 -2262 157154 -2026
rect 162186 705002 162422 705238
rect 162186 704682 162422 704918
rect 162186 695258 162422 695494
rect 162186 688258 162422 688494
rect 162186 681258 162422 681494
rect 162186 674258 162422 674494
rect 162186 667258 162422 667494
rect 162186 660258 162422 660494
rect 162186 653258 162422 653494
rect 162186 646258 162422 646494
rect 162186 639258 162422 639494
rect 162186 632258 162422 632494
rect 162186 625258 162422 625494
rect 162186 618258 162422 618494
rect 162186 611258 162422 611494
rect 162186 604258 162422 604494
rect 162186 597258 162422 597494
rect 162186 590258 162422 590494
rect 162186 583258 162422 583494
rect 162186 576258 162422 576494
rect 162186 569258 162422 569494
rect 162186 562258 162422 562494
rect 162186 555258 162422 555494
rect 162186 548258 162422 548494
rect 162186 541258 162422 541494
rect 162186 534258 162422 534494
rect 162186 527258 162422 527494
rect 162186 520258 162422 520494
rect 162186 513258 162422 513494
rect 162186 506258 162422 506494
rect 162186 499258 162422 499494
rect 162186 492258 162422 492494
rect 162186 485258 162422 485494
rect 162186 478258 162422 478494
rect 162186 471258 162422 471494
rect 162186 464258 162422 464494
rect 162186 457258 162422 457494
rect 162186 450258 162422 450494
rect 162186 443258 162422 443494
rect 162186 436258 162422 436494
rect 162186 429258 162422 429494
rect 162186 422258 162422 422494
rect 162186 415258 162422 415494
rect 162186 408258 162422 408494
rect 162186 401258 162422 401494
rect 162186 394258 162422 394494
rect 162186 387258 162422 387494
rect 162186 380258 162422 380494
rect 162186 373258 162422 373494
rect 162186 366258 162422 366494
rect 162186 359258 162422 359494
rect 162186 352258 162422 352494
rect 162186 345258 162422 345494
rect 162186 338258 162422 338494
rect 162186 331258 162422 331494
rect 162186 324258 162422 324494
rect 162186 317258 162422 317494
rect 162186 310258 162422 310494
rect 162186 303258 162422 303494
rect 162186 296258 162422 296494
rect 162186 289258 162422 289494
rect 162186 282258 162422 282494
rect 162186 275258 162422 275494
rect 162186 268258 162422 268494
rect 162186 261258 162422 261494
rect 162186 254258 162422 254494
rect 162186 247258 162422 247494
rect 162186 240258 162422 240494
rect 162186 233258 162422 233494
rect 162186 226258 162422 226494
rect 162186 219258 162422 219494
rect 162186 212258 162422 212494
rect 162186 205258 162422 205494
rect 162186 198258 162422 198494
rect 162186 191258 162422 191494
rect 162186 184258 162422 184494
rect 162186 177258 162422 177494
rect 162186 170258 162422 170494
rect 162186 163258 162422 163494
rect 162186 156258 162422 156494
rect 162186 149258 162422 149494
rect 162186 142258 162422 142494
rect 162186 135258 162422 135494
rect 162186 128258 162422 128494
rect 162186 121258 162422 121494
rect 162186 114258 162422 114494
rect 162186 107258 162422 107494
rect 162186 100258 162422 100494
rect 162186 93258 162422 93494
rect 162186 86258 162422 86494
rect 162186 79258 162422 79494
rect 162186 72258 162422 72494
rect 162186 65258 162422 65494
rect 162186 58258 162422 58494
rect 162186 51258 162422 51494
rect 162186 44258 162422 44494
rect 162186 37258 162422 37494
rect 162186 30258 162422 30494
rect 162186 23258 162422 23494
rect 162186 16258 162422 16494
rect 162186 9258 162422 9494
rect 162186 2258 162422 2494
rect 162186 -982 162422 -746
rect 162186 -1302 162422 -1066
rect 163918 705962 164154 706198
rect 163918 705642 164154 705878
rect 163918 696325 164154 696561
rect 163918 689325 164154 689561
rect 163918 682325 164154 682561
rect 163918 675325 164154 675561
rect 163918 668325 164154 668561
rect 163918 661325 164154 661561
rect 163918 654325 164154 654561
rect 163918 647325 164154 647561
rect 163918 640325 164154 640561
rect 163918 633325 164154 633561
rect 163918 626325 164154 626561
rect 163918 619325 164154 619561
rect 163918 612325 164154 612561
rect 163918 605325 164154 605561
rect 163918 598325 164154 598561
rect 163918 591325 164154 591561
rect 163918 584325 164154 584561
rect 163918 577325 164154 577561
rect 163918 570325 164154 570561
rect 163918 563325 164154 563561
rect 163918 556325 164154 556561
rect 163918 549325 164154 549561
rect 163918 542325 164154 542561
rect 163918 535325 164154 535561
rect 163918 528325 164154 528561
rect 163918 521325 164154 521561
rect 163918 514325 164154 514561
rect 163918 507325 164154 507561
rect 163918 500325 164154 500561
rect 163918 493325 164154 493561
rect 163918 486325 164154 486561
rect 163918 479325 164154 479561
rect 163918 472325 164154 472561
rect 163918 465325 164154 465561
rect 163918 458325 164154 458561
rect 163918 451325 164154 451561
rect 163918 444325 164154 444561
rect 163918 437325 164154 437561
rect 163918 430325 164154 430561
rect 163918 423325 164154 423561
rect 163918 416325 164154 416561
rect 163918 409325 164154 409561
rect 163918 402325 164154 402561
rect 163918 395325 164154 395561
rect 163918 388325 164154 388561
rect 163918 381325 164154 381561
rect 163918 374325 164154 374561
rect 163918 367325 164154 367561
rect 163918 360325 164154 360561
rect 163918 353325 164154 353561
rect 163918 346325 164154 346561
rect 163918 339325 164154 339561
rect 163918 332325 164154 332561
rect 163918 325325 164154 325561
rect 163918 318325 164154 318561
rect 163918 311325 164154 311561
rect 163918 304325 164154 304561
rect 163918 297325 164154 297561
rect 163918 290325 164154 290561
rect 163918 283325 164154 283561
rect 163918 276325 164154 276561
rect 163918 269325 164154 269561
rect 163918 262325 164154 262561
rect 163918 255325 164154 255561
rect 163918 248325 164154 248561
rect 163918 241325 164154 241561
rect 163918 234325 164154 234561
rect 163918 227325 164154 227561
rect 163918 220325 164154 220561
rect 163918 213325 164154 213561
rect 163918 206325 164154 206561
rect 163918 199325 164154 199561
rect 163918 192325 164154 192561
rect 163918 185325 164154 185561
rect 163918 178325 164154 178561
rect 163918 171325 164154 171561
rect 163918 164325 164154 164561
rect 163918 157325 164154 157561
rect 163918 150325 164154 150561
rect 163918 143325 164154 143561
rect 163918 136325 164154 136561
rect 163918 129325 164154 129561
rect 163918 122325 164154 122561
rect 163918 115325 164154 115561
rect 163918 108325 164154 108561
rect 163918 101325 164154 101561
rect 163918 94325 164154 94561
rect 163918 87325 164154 87561
rect 163918 80325 164154 80561
rect 163918 73325 164154 73561
rect 163918 66325 164154 66561
rect 163918 59325 164154 59561
rect 163918 52325 164154 52561
rect 163918 45325 164154 45561
rect 163918 38325 164154 38561
rect 163918 31325 164154 31561
rect 163918 24325 164154 24561
rect 163918 17325 164154 17561
rect 163918 10325 164154 10561
rect 163918 3325 164154 3561
rect 163918 -1942 164154 -1706
rect 163918 -2262 164154 -2026
rect 169186 705002 169422 705238
rect 169186 704682 169422 704918
rect 169186 695258 169422 695494
rect 169186 688258 169422 688494
rect 169186 681258 169422 681494
rect 169186 674258 169422 674494
rect 169186 667258 169422 667494
rect 169186 660258 169422 660494
rect 169186 653258 169422 653494
rect 169186 646258 169422 646494
rect 169186 639258 169422 639494
rect 169186 632258 169422 632494
rect 169186 625258 169422 625494
rect 169186 618258 169422 618494
rect 169186 611258 169422 611494
rect 169186 604258 169422 604494
rect 169186 597258 169422 597494
rect 169186 590258 169422 590494
rect 169186 583258 169422 583494
rect 169186 576258 169422 576494
rect 169186 569258 169422 569494
rect 169186 562258 169422 562494
rect 169186 555258 169422 555494
rect 169186 548258 169422 548494
rect 169186 541258 169422 541494
rect 169186 534258 169422 534494
rect 169186 527258 169422 527494
rect 169186 520258 169422 520494
rect 169186 513258 169422 513494
rect 169186 506258 169422 506494
rect 169186 499258 169422 499494
rect 169186 492258 169422 492494
rect 169186 485258 169422 485494
rect 169186 478258 169422 478494
rect 169186 471258 169422 471494
rect 169186 464258 169422 464494
rect 169186 457258 169422 457494
rect 169186 450258 169422 450494
rect 169186 443258 169422 443494
rect 169186 436258 169422 436494
rect 169186 429258 169422 429494
rect 169186 422258 169422 422494
rect 169186 415258 169422 415494
rect 169186 408258 169422 408494
rect 169186 401258 169422 401494
rect 169186 394258 169422 394494
rect 169186 387258 169422 387494
rect 169186 380258 169422 380494
rect 169186 373258 169422 373494
rect 169186 366258 169422 366494
rect 169186 359258 169422 359494
rect 169186 352258 169422 352494
rect 169186 345258 169422 345494
rect 169186 338258 169422 338494
rect 169186 331258 169422 331494
rect 169186 324258 169422 324494
rect 169186 317258 169422 317494
rect 169186 310258 169422 310494
rect 169186 303258 169422 303494
rect 169186 296258 169422 296494
rect 169186 289258 169422 289494
rect 169186 282258 169422 282494
rect 169186 275258 169422 275494
rect 169186 268258 169422 268494
rect 169186 261258 169422 261494
rect 169186 254258 169422 254494
rect 169186 247258 169422 247494
rect 169186 240258 169422 240494
rect 169186 233258 169422 233494
rect 169186 226258 169422 226494
rect 169186 219258 169422 219494
rect 169186 212258 169422 212494
rect 169186 205258 169422 205494
rect 169186 198258 169422 198494
rect 169186 191258 169422 191494
rect 169186 184258 169422 184494
rect 169186 177258 169422 177494
rect 169186 170258 169422 170494
rect 169186 163258 169422 163494
rect 169186 156258 169422 156494
rect 169186 149258 169422 149494
rect 169186 142258 169422 142494
rect 169186 135258 169422 135494
rect 169186 128258 169422 128494
rect 169186 121258 169422 121494
rect 169186 114258 169422 114494
rect 169186 107258 169422 107494
rect 169186 100258 169422 100494
rect 169186 93258 169422 93494
rect 169186 86258 169422 86494
rect 169186 79258 169422 79494
rect 169186 72258 169422 72494
rect 169186 65258 169422 65494
rect 169186 58258 169422 58494
rect 169186 51258 169422 51494
rect 169186 44258 169422 44494
rect 169186 37258 169422 37494
rect 169186 30258 169422 30494
rect 169186 23258 169422 23494
rect 169186 16258 169422 16494
rect 169186 9258 169422 9494
rect 169186 2258 169422 2494
rect 169186 -982 169422 -746
rect 169186 -1302 169422 -1066
rect 170918 705962 171154 706198
rect 170918 705642 171154 705878
rect 170918 696325 171154 696561
rect 170918 689325 171154 689561
rect 170918 682325 171154 682561
rect 170918 675325 171154 675561
rect 170918 668325 171154 668561
rect 170918 661325 171154 661561
rect 170918 654325 171154 654561
rect 170918 647325 171154 647561
rect 170918 640325 171154 640561
rect 170918 633325 171154 633561
rect 170918 626325 171154 626561
rect 170918 619325 171154 619561
rect 170918 612325 171154 612561
rect 170918 605325 171154 605561
rect 170918 598325 171154 598561
rect 170918 591325 171154 591561
rect 170918 584325 171154 584561
rect 170918 577325 171154 577561
rect 170918 570325 171154 570561
rect 170918 563325 171154 563561
rect 170918 556325 171154 556561
rect 170918 549325 171154 549561
rect 170918 542325 171154 542561
rect 170918 535325 171154 535561
rect 170918 528325 171154 528561
rect 170918 521325 171154 521561
rect 170918 514325 171154 514561
rect 170918 507325 171154 507561
rect 170918 500325 171154 500561
rect 170918 493325 171154 493561
rect 170918 486325 171154 486561
rect 170918 479325 171154 479561
rect 170918 472325 171154 472561
rect 170918 465325 171154 465561
rect 170918 458325 171154 458561
rect 170918 451325 171154 451561
rect 170918 444325 171154 444561
rect 170918 437325 171154 437561
rect 170918 430325 171154 430561
rect 170918 423325 171154 423561
rect 170918 416325 171154 416561
rect 170918 409325 171154 409561
rect 170918 402325 171154 402561
rect 170918 395325 171154 395561
rect 170918 388325 171154 388561
rect 170918 381325 171154 381561
rect 170918 374325 171154 374561
rect 170918 367325 171154 367561
rect 170918 360325 171154 360561
rect 170918 353325 171154 353561
rect 170918 346325 171154 346561
rect 170918 339325 171154 339561
rect 170918 332325 171154 332561
rect 170918 325325 171154 325561
rect 170918 318325 171154 318561
rect 170918 311325 171154 311561
rect 170918 304325 171154 304561
rect 170918 297325 171154 297561
rect 170918 290325 171154 290561
rect 170918 283325 171154 283561
rect 170918 276325 171154 276561
rect 170918 269325 171154 269561
rect 170918 262325 171154 262561
rect 170918 255325 171154 255561
rect 170918 248325 171154 248561
rect 170918 241325 171154 241561
rect 170918 234325 171154 234561
rect 170918 227325 171154 227561
rect 170918 220325 171154 220561
rect 170918 213325 171154 213561
rect 170918 206325 171154 206561
rect 170918 199325 171154 199561
rect 170918 192325 171154 192561
rect 170918 185325 171154 185561
rect 170918 178325 171154 178561
rect 170918 171325 171154 171561
rect 170918 164325 171154 164561
rect 170918 157325 171154 157561
rect 170918 150325 171154 150561
rect 170918 143325 171154 143561
rect 170918 136325 171154 136561
rect 170918 129325 171154 129561
rect 170918 122325 171154 122561
rect 170918 115325 171154 115561
rect 170918 108325 171154 108561
rect 170918 101325 171154 101561
rect 170918 94325 171154 94561
rect 170918 87325 171154 87561
rect 170918 80325 171154 80561
rect 170918 73325 171154 73561
rect 170918 66325 171154 66561
rect 170918 59325 171154 59561
rect 170918 52325 171154 52561
rect 170918 45325 171154 45561
rect 170918 38325 171154 38561
rect 170918 31325 171154 31561
rect 170918 24325 171154 24561
rect 170918 17325 171154 17561
rect 170918 10325 171154 10561
rect 170918 3325 171154 3561
rect 170918 -1942 171154 -1706
rect 170918 -2262 171154 -2026
rect 176186 705002 176422 705238
rect 176186 704682 176422 704918
rect 176186 695258 176422 695494
rect 176186 688258 176422 688494
rect 176186 681258 176422 681494
rect 176186 674258 176422 674494
rect 176186 667258 176422 667494
rect 176186 660258 176422 660494
rect 176186 653258 176422 653494
rect 176186 646258 176422 646494
rect 176186 639258 176422 639494
rect 176186 632258 176422 632494
rect 176186 625258 176422 625494
rect 176186 618258 176422 618494
rect 176186 611258 176422 611494
rect 176186 604258 176422 604494
rect 176186 597258 176422 597494
rect 176186 590258 176422 590494
rect 176186 583258 176422 583494
rect 176186 576258 176422 576494
rect 176186 569258 176422 569494
rect 176186 562258 176422 562494
rect 176186 555258 176422 555494
rect 176186 548258 176422 548494
rect 176186 541258 176422 541494
rect 176186 534258 176422 534494
rect 176186 527258 176422 527494
rect 176186 520258 176422 520494
rect 176186 513258 176422 513494
rect 176186 506258 176422 506494
rect 176186 499258 176422 499494
rect 176186 492258 176422 492494
rect 176186 485258 176422 485494
rect 176186 478258 176422 478494
rect 176186 471258 176422 471494
rect 176186 464258 176422 464494
rect 176186 457258 176422 457494
rect 176186 450258 176422 450494
rect 176186 443258 176422 443494
rect 176186 436258 176422 436494
rect 176186 429258 176422 429494
rect 176186 422258 176422 422494
rect 176186 415258 176422 415494
rect 176186 408258 176422 408494
rect 176186 401258 176422 401494
rect 176186 394258 176422 394494
rect 176186 387258 176422 387494
rect 176186 380258 176422 380494
rect 176186 373258 176422 373494
rect 176186 366258 176422 366494
rect 176186 359258 176422 359494
rect 176186 352258 176422 352494
rect 176186 345258 176422 345494
rect 176186 338258 176422 338494
rect 176186 331258 176422 331494
rect 176186 324258 176422 324494
rect 176186 317258 176422 317494
rect 176186 310258 176422 310494
rect 176186 303258 176422 303494
rect 176186 296258 176422 296494
rect 176186 289258 176422 289494
rect 176186 282258 176422 282494
rect 176186 275258 176422 275494
rect 176186 268258 176422 268494
rect 176186 261258 176422 261494
rect 176186 254258 176422 254494
rect 176186 247258 176422 247494
rect 176186 240258 176422 240494
rect 176186 233258 176422 233494
rect 176186 226258 176422 226494
rect 176186 219258 176422 219494
rect 176186 212258 176422 212494
rect 176186 205258 176422 205494
rect 176186 198258 176422 198494
rect 176186 191258 176422 191494
rect 176186 184258 176422 184494
rect 176186 177258 176422 177494
rect 176186 170258 176422 170494
rect 176186 163258 176422 163494
rect 176186 156258 176422 156494
rect 176186 149258 176422 149494
rect 176186 142258 176422 142494
rect 176186 135258 176422 135494
rect 176186 128258 176422 128494
rect 176186 121258 176422 121494
rect 176186 114258 176422 114494
rect 176186 107258 176422 107494
rect 176186 100258 176422 100494
rect 176186 93258 176422 93494
rect 176186 86258 176422 86494
rect 176186 79258 176422 79494
rect 176186 72258 176422 72494
rect 176186 65258 176422 65494
rect 176186 58258 176422 58494
rect 176186 51258 176422 51494
rect 176186 44258 176422 44494
rect 176186 37258 176422 37494
rect 176186 30258 176422 30494
rect 176186 23258 176422 23494
rect 176186 16258 176422 16494
rect 176186 9258 176422 9494
rect 176186 2258 176422 2494
rect 176186 -982 176422 -746
rect 176186 -1302 176422 -1066
rect 177918 705962 178154 706198
rect 177918 705642 178154 705878
rect 177918 696325 178154 696561
rect 177918 689325 178154 689561
rect 177918 682325 178154 682561
rect 177918 675325 178154 675561
rect 177918 668325 178154 668561
rect 177918 661325 178154 661561
rect 177918 654325 178154 654561
rect 177918 647325 178154 647561
rect 177918 640325 178154 640561
rect 177918 633325 178154 633561
rect 177918 626325 178154 626561
rect 177918 619325 178154 619561
rect 177918 612325 178154 612561
rect 177918 605325 178154 605561
rect 177918 598325 178154 598561
rect 177918 591325 178154 591561
rect 177918 584325 178154 584561
rect 177918 577325 178154 577561
rect 177918 570325 178154 570561
rect 177918 563325 178154 563561
rect 177918 556325 178154 556561
rect 177918 549325 178154 549561
rect 177918 542325 178154 542561
rect 177918 535325 178154 535561
rect 177918 528325 178154 528561
rect 177918 521325 178154 521561
rect 177918 514325 178154 514561
rect 177918 507325 178154 507561
rect 177918 500325 178154 500561
rect 177918 493325 178154 493561
rect 177918 486325 178154 486561
rect 177918 479325 178154 479561
rect 177918 472325 178154 472561
rect 177918 465325 178154 465561
rect 177918 458325 178154 458561
rect 177918 451325 178154 451561
rect 177918 444325 178154 444561
rect 177918 437325 178154 437561
rect 177918 430325 178154 430561
rect 177918 423325 178154 423561
rect 177918 416325 178154 416561
rect 177918 409325 178154 409561
rect 177918 402325 178154 402561
rect 177918 395325 178154 395561
rect 177918 388325 178154 388561
rect 177918 381325 178154 381561
rect 177918 374325 178154 374561
rect 177918 367325 178154 367561
rect 177918 360325 178154 360561
rect 177918 353325 178154 353561
rect 177918 346325 178154 346561
rect 177918 339325 178154 339561
rect 177918 332325 178154 332561
rect 177918 325325 178154 325561
rect 177918 318325 178154 318561
rect 177918 311325 178154 311561
rect 177918 304325 178154 304561
rect 177918 297325 178154 297561
rect 177918 290325 178154 290561
rect 177918 283325 178154 283561
rect 177918 276325 178154 276561
rect 177918 269325 178154 269561
rect 177918 262325 178154 262561
rect 177918 255325 178154 255561
rect 177918 248325 178154 248561
rect 177918 241325 178154 241561
rect 177918 234325 178154 234561
rect 177918 227325 178154 227561
rect 177918 220325 178154 220561
rect 177918 213325 178154 213561
rect 177918 206325 178154 206561
rect 177918 199325 178154 199561
rect 177918 192325 178154 192561
rect 177918 185325 178154 185561
rect 177918 178325 178154 178561
rect 177918 171325 178154 171561
rect 177918 164325 178154 164561
rect 177918 157325 178154 157561
rect 177918 150325 178154 150561
rect 177918 143325 178154 143561
rect 177918 136325 178154 136561
rect 177918 129325 178154 129561
rect 177918 122325 178154 122561
rect 177918 115325 178154 115561
rect 177918 108325 178154 108561
rect 177918 101325 178154 101561
rect 177918 94325 178154 94561
rect 177918 87325 178154 87561
rect 177918 80325 178154 80561
rect 177918 73325 178154 73561
rect 177918 66325 178154 66561
rect 177918 59325 178154 59561
rect 177918 52325 178154 52561
rect 177918 45325 178154 45561
rect 177918 38325 178154 38561
rect 177918 31325 178154 31561
rect 177918 24325 178154 24561
rect 177918 17325 178154 17561
rect 177918 10325 178154 10561
rect 177918 3325 178154 3561
rect 177918 -1942 178154 -1706
rect 177918 -2262 178154 -2026
rect 183186 705002 183422 705238
rect 183186 704682 183422 704918
rect 183186 695258 183422 695494
rect 183186 688258 183422 688494
rect 183186 681258 183422 681494
rect 183186 674258 183422 674494
rect 183186 667258 183422 667494
rect 183186 660258 183422 660494
rect 183186 653258 183422 653494
rect 183186 646258 183422 646494
rect 183186 639258 183422 639494
rect 183186 632258 183422 632494
rect 183186 625258 183422 625494
rect 183186 618258 183422 618494
rect 183186 611258 183422 611494
rect 183186 604258 183422 604494
rect 183186 597258 183422 597494
rect 183186 590258 183422 590494
rect 183186 583258 183422 583494
rect 183186 576258 183422 576494
rect 183186 569258 183422 569494
rect 183186 562258 183422 562494
rect 183186 555258 183422 555494
rect 183186 548258 183422 548494
rect 183186 541258 183422 541494
rect 183186 534258 183422 534494
rect 183186 527258 183422 527494
rect 183186 520258 183422 520494
rect 183186 513258 183422 513494
rect 183186 506258 183422 506494
rect 183186 499258 183422 499494
rect 183186 492258 183422 492494
rect 183186 485258 183422 485494
rect 183186 478258 183422 478494
rect 183186 471258 183422 471494
rect 183186 464258 183422 464494
rect 183186 457258 183422 457494
rect 183186 450258 183422 450494
rect 183186 443258 183422 443494
rect 183186 436258 183422 436494
rect 183186 429258 183422 429494
rect 183186 422258 183422 422494
rect 183186 415258 183422 415494
rect 183186 408258 183422 408494
rect 183186 401258 183422 401494
rect 183186 394258 183422 394494
rect 183186 387258 183422 387494
rect 183186 380258 183422 380494
rect 183186 373258 183422 373494
rect 183186 366258 183422 366494
rect 183186 359258 183422 359494
rect 183186 352258 183422 352494
rect 183186 345258 183422 345494
rect 183186 338258 183422 338494
rect 183186 331258 183422 331494
rect 183186 324258 183422 324494
rect 183186 317258 183422 317494
rect 183186 310258 183422 310494
rect 183186 303258 183422 303494
rect 183186 296258 183422 296494
rect 183186 289258 183422 289494
rect 183186 282258 183422 282494
rect 183186 275258 183422 275494
rect 183186 268258 183422 268494
rect 183186 261258 183422 261494
rect 183186 254258 183422 254494
rect 183186 247258 183422 247494
rect 183186 240258 183422 240494
rect 183186 233258 183422 233494
rect 183186 226258 183422 226494
rect 183186 219258 183422 219494
rect 183186 212258 183422 212494
rect 183186 205258 183422 205494
rect 183186 198258 183422 198494
rect 183186 191258 183422 191494
rect 183186 184258 183422 184494
rect 183186 177258 183422 177494
rect 183186 170258 183422 170494
rect 183186 163258 183422 163494
rect 183186 156258 183422 156494
rect 183186 149258 183422 149494
rect 183186 142258 183422 142494
rect 183186 135258 183422 135494
rect 183186 128258 183422 128494
rect 183186 121258 183422 121494
rect 183186 114258 183422 114494
rect 183186 107258 183422 107494
rect 183186 100258 183422 100494
rect 183186 93258 183422 93494
rect 183186 86258 183422 86494
rect 183186 79258 183422 79494
rect 183186 72258 183422 72494
rect 183186 65258 183422 65494
rect 183186 58258 183422 58494
rect 183186 51258 183422 51494
rect 183186 44258 183422 44494
rect 183186 37258 183422 37494
rect 183186 30258 183422 30494
rect 183186 23258 183422 23494
rect 183186 16258 183422 16494
rect 183186 9258 183422 9494
rect 183186 2258 183422 2494
rect 183186 -982 183422 -746
rect 183186 -1302 183422 -1066
rect 184918 705962 185154 706198
rect 184918 705642 185154 705878
rect 184918 696325 185154 696561
rect 184918 689325 185154 689561
rect 184918 682325 185154 682561
rect 184918 675325 185154 675561
rect 184918 668325 185154 668561
rect 184918 661325 185154 661561
rect 184918 654325 185154 654561
rect 184918 647325 185154 647561
rect 184918 640325 185154 640561
rect 184918 633325 185154 633561
rect 184918 626325 185154 626561
rect 184918 619325 185154 619561
rect 184918 612325 185154 612561
rect 184918 605325 185154 605561
rect 184918 598325 185154 598561
rect 184918 591325 185154 591561
rect 184918 584325 185154 584561
rect 184918 577325 185154 577561
rect 184918 570325 185154 570561
rect 184918 563325 185154 563561
rect 184918 556325 185154 556561
rect 184918 549325 185154 549561
rect 184918 542325 185154 542561
rect 184918 535325 185154 535561
rect 184918 528325 185154 528561
rect 184918 521325 185154 521561
rect 184918 514325 185154 514561
rect 184918 507325 185154 507561
rect 184918 500325 185154 500561
rect 184918 493325 185154 493561
rect 184918 486325 185154 486561
rect 184918 479325 185154 479561
rect 184918 472325 185154 472561
rect 184918 465325 185154 465561
rect 184918 458325 185154 458561
rect 184918 451325 185154 451561
rect 184918 444325 185154 444561
rect 184918 437325 185154 437561
rect 184918 430325 185154 430561
rect 184918 423325 185154 423561
rect 184918 416325 185154 416561
rect 184918 409325 185154 409561
rect 184918 402325 185154 402561
rect 184918 395325 185154 395561
rect 184918 388325 185154 388561
rect 184918 381325 185154 381561
rect 184918 374325 185154 374561
rect 184918 367325 185154 367561
rect 184918 360325 185154 360561
rect 184918 353325 185154 353561
rect 184918 346325 185154 346561
rect 184918 339325 185154 339561
rect 184918 332325 185154 332561
rect 184918 325325 185154 325561
rect 184918 318325 185154 318561
rect 184918 311325 185154 311561
rect 184918 304325 185154 304561
rect 184918 297325 185154 297561
rect 184918 290325 185154 290561
rect 184918 283325 185154 283561
rect 184918 276325 185154 276561
rect 184918 269325 185154 269561
rect 184918 262325 185154 262561
rect 184918 255325 185154 255561
rect 184918 248325 185154 248561
rect 184918 241325 185154 241561
rect 184918 234325 185154 234561
rect 184918 227325 185154 227561
rect 184918 220325 185154 220561
rect 184918 213325 185154 213561
rect 184918 206325 185154 206561
rect 184918 199325 185154 199561
rect 184918 192325 185154 192561
rect 184918 185325 185154 185561
rect 184918 178325 185154 178561
rect 184918 171325 185154 171561
rect 184918 164325 185154 164561
rect 184918 157325 185154 157561
rect 184918 150325 185154 150561
rect 184918 143325 185154 143561
rect 184918 136325 185154 136561
rect 184918 129325 185154 129561
rect 184918 122325 185154 122561
rect 184918 115325 185154 115561
rect 184918 108325 185154 108561
rect 184918 101325 185154 101561
rect 184918 94325 185154 94561
rect 184918 87325 185154 87561
rect 184918 80325 185154 80561
rect 184918 73325 185154 73561
rect 184918 66325 185154 66561
rect 184918 59325 185154 59561
rect 184918 52325 185154 52561
rect 184918 45325 185154 45561
rect 184918 38325 185154 38561
rect 184918 31325 185154 31561
rect 184918 24325 185154 24561
rect 184918 17325 185154 17561
rect 184918 10325 185154 10561
rect 184918 3325 185154 3561
rect 184918 -1942 185154 -1706
rect 184918 -2262 185154 -2026
rect 190186 705002 190422 705238
rect 190186 704682 190422 704918
rect 190186 695258 190422 695494
rect 190186 688258 190422 688494
rect 190186 681258 190422 681494
rect 190186 674258 190422 674494
rect 190186 667258 190422 667494
rect 190186 660258 190422 660494
rect 190186 653258 190422 653494
rect 190186 646258 190422 646494
rect 190186 639258 190422 639494
rect 190186 632258 190422 632494
rect 190186 625258 190422 625494
rect 190186 618258 190422 618494
rect 190186 611258 190422 611494
rect 190186 604258 190422 604494
rect 190186 597258 190422 597494
rect 190186 590258 190422 590494
rect 190186 583258 190422 583494
rect 190186 576258 190422 576494
rect 190186 569258 190422 569494
rect 190186 562258 190422 562494
rect 190186 555258 190422 555494
rect 190186 548258 190422 548494
rect 190186 541258 190422 541494
rect 190186 534258 190422 534494
rect 190186 527258 190422 527494
rect 190186 520258 190422 520494
rect 190186 513258 190422 513494
rect 190186 506258 190422 506494
rect 190186 499258 190422 499494
rect 190186 492258 190422 492494
rect 190186 485258 190422 485494
rect 190186 478258 190422 478494
rect 190186 471258 190422 471494
rect 190186 464258 190422 464494
rect 190186 457258 190422 457494
rect 190186 450258 190422 450494
rect 190186 443258 190422 443494
rect 190186 436258 190422 436494
rect 190186 429258 190422 429494
rect 190186 422258 190422 422494
rect 190186 415258 190422 415494
rect 190186 408258 190422 408494
rect 190186 401258 190422 401494
rect 190186 394258 190422 394494
rect 190186 387258 190422 387494
rect 190186 380258 190422 380494
rect 190186 373258 190422 373494
rect 190186 366258 190422 366494
rect 190186 359258 190422 359494
rect 190186 352258 190422 352494
rect 190186 345258 190422 345494
rect 190186 338258 190422 338494
rect 190186 331258 190422 331494
rect 190186 324258 190422 324494
rect 190186 317258 190422 317494
rect 190186 310258 190422 310494
rect 190186 303258 190422 303494
rect 190186 296258 190422 296494
rect 190186 289258 190422 289494
rect 190186 282258 190422 282494
rect 190186 275258 190422 275494
rect 190186 268258 190422 268494
rect 190186 261258 190422 261494
rect 190186 254258 190422 254494
rect 190186 247258 190422 247494
rect 190186 240258 190422 240494
rect 190186 233258 190422 233494
rect 190186 226258 190422 226494
rect 190186 219258 190422 219494
rect 190186 212258 190422 212494
rect 190186 205258 190422 205494
rect 190186 198258 190422 198494
rect 190186 191258 190422 191494
rect 190186 184258 190422 184494
rect 190186 177258 190422 177494
rect 190186 170258 190422 170494
rect 190186 163258 190422 163494
rect 190186 156258 190422 156494
rect 190186 149258 190422 149494
rect 190186 142258 190422 142494
rect 190186 135258 190422 135494
rect 190186 128258 190422 128494
rect 190186 121258 190422 121494
rect 190186 114258 190422 114494
rect 190186 107258 190422 107494
rect 190186 100258 190422 100494
rect 190186 93258 190422 93494
rect 190186 86258 190422 86494
rect 190186 79258 190422 79494
rect 190186 72258 190422 72494
rect 190186 65258 190422 65494
rect 190186 58258 190422 58494
rect 190186 51258 190422 51494
rect 190186 44258 190422 44494
rect 190186 37258 190422 37494
rect 190186 30258 190422 30494
rect 190186 23258 190422 23494
rect 190186 16258 190422 16494
rect 190186 9258 190422 9494
rect 190186 2258 190422 2494
rect 190186 -982 190422 -746
rect 190186 -1302 190422 -1066
rect 191918 705962 192154 706198
rect 191918 705642 192154 705878
rect 191918 696325 192154 696561
rect 191918 689325 192154 689561
rect 191918 682325 192154 682561
rect 191918 675325 192154 675561
rect 191918 668325 192154 668561
rect 191918 661325 192154 661561
rect 191918 654325 192154 654561
rect 191918 647325 192154 647561
rect 191918 640325 192154 640561
rect 191918 633325 192154 633561
rect 191918 626325 192154 626561
rect 191918 619325 192154 619561
rect 191918 612325 192154 612561
rect 191918 605325 192154 605561
rect 191918 598325 192154 598561
rect 191918 591325 192154 591561
rect 191918 584325 192154 584561
rect 191918 577325 192154 577561
rect 191918 570325 192154 570561
rect 191918 563325 192154 563561
rect 191918 556325 192154 556561
rect 191918 549325 192154 549561
rect 191918 542325 192154 542561
rect 191918 535325 192154 535561
rect 191918 528325 192154 528561
rect 191918 521325 192154 521561
rect 191918 514325 192154 514561
rect 191918 507325 192154 507561
rect 191918 500325 192154 500561
rect 191918 493325 192154 493561
rect 191918 486325 192154 486561
rect 191918 479325 192154 479561
rect 191918 472325 192154 472561
rect 191918 465325 192154 465561
rect 191918 458325 192154 458561
rect 191918 451325 192154 451561
rect 191918 444325 192154 444561
rect 191918 437325 192154 437561
rect 191918 430325 192154 430561
rect 191918 423325 192154 423561
rect 191918 416325 192154 416561
rect 191918 409325 192154 409561
rect 191918 402325 192154 402561
rect 191918 395325 192154 395561
rect 191918 388325 192154 388561
rect 191918 381325 192154 381561
rect 191918 374325 192154 374561
rect 191918 367325 192154 367561
rect 191918 360325 192154 360561
rect 191918 353325 192154 353561
rect 191918 346325 192154 346561
rect 191918 339325 192154 339561
rect 191918 332325 192154 332561
rect 191918 325325 192154 325561
rect 191918 318325 192154 318561
rect 191918 311325 192154 311561
rect 191918 304325 192154 304561
rect 191918 297325 192154 297561
rect 191918 290325 192154 290561
rect 191918 283325 192154 283561
rect 191918 276325 192154 276561
rect 191918 269325 192154 269561
rect 191918 262325 192154 262561
rect 191918 255325 192154 255561
rect 191918 248325 192154 248561
rect 191918 241325 192154 241561
rect 191918 234325 192154 234561
rect 191918 227325 192154 227561
rect 191918 220325 192154 220561
rect 191918 213325 192154 213561
rect 191918 206325 192154 206561
rect 191918 199325 192154 199561
rect 191918 192325 192154 192561
rect 191918 185325 192154 185561
rect 191918 178325 192154 178561
rect 191918 171325 192154 171561
rect 191918 164325 192154 164561
rect 191918 157325 192154 157561
rect 191918 150325 192154 150561
rect 191918 143325 192154 143561
rect 191918 136325 192154 136561
rect 191918 129325 192154 129561
rect 191918 122325 192154 122561
rect 191918 115325 192154 115561
rect 191918 108325 192154 108561
rect 191918 101325 192154 101561
rect 191918 94325 192154 94561
rect 191918 87325 192154 87561
rect 191918 80325 192154 80561
rect 191918 73325 192154 73561
rect 191918 66325 192154 66561
rect 191918 59325 192154 59561
rect 191918 52325 192154 52561
rect 191918 45325 192154 45561
rect 191918 38325 192154 38561
rect 191918 31325 192154 31561
rect 191918 24325 192154 24561
rect 191918 17325 192154 17561
rect 191918 10325 192154 10561
rect 191918 3325 192154 3561
rect 191918 -1942 192154 -1706
rect 191918 -2262 192154 -2026
rect 197186 705002 197422 705238
rect 197186 704682 197422 704918
rect 197186 695258 197422 695494
rect 197186 688258 197422 688494
rect 197186 681258 197422 681494
rect 197186 674258 197422 674494
rect 197186 667258 197422 667494
rect 197186 660258 197422 660494
rect 197186 653258 197422 653494
rect 197186 646258 197422 646494
rect 197186 639258 197422 639494
rect 197186 632258 197422 632494
rect 197186 625258 197422 625494
rect 197186 618258 197422 618494
rect 197186 611258 197422 611494
rect 197186 604258 197422 604494
rect 197186 597258 197422 597494
rect 197186 590258 197422 590494
rect 197186 583258 197422 583494
rect 197186 576258 197422 576494
rect 197186 569258 197422 569494
rect 197186 562258 197422 562494
rect 197186 555258 197422 555494
rect 197186 548258 197422 548494
rect 197186 541258 197422 541494
rect 197186 534258 197422 534494
rect 197186 527258 197422 527494
rect 197186 520258 197422 520494
rect 197186 513258 197422 513494
rect 197186 506258 197422 506494
rect 197186 499258 197422 499494
rect 197186 492258 197422 492494
rect 197186 485258 197422 485494
rect 197186 478258 197422 478494
rect 197186 471258 197422 471494
rect 197186 464258 197422 464494
rect 197186 457258 197422 457494
rect 197186 450258 197422 450494
rect 197186 443258 197422 443494
rect 197186 436258 197422 436494
rect 197186 429258 197422 429494
rect 197186 422258 197422 422494
rect 197186 415258 197422 415494
rect 197186 408258 197422 408494
rect 197186 401258 197422 401494
rect 197186 394258 197422 394494
rect 197186 387258 197422 387494
rect 197186 380258 197422 380494
rect 197186 373258 197422 373494
rect 197186 366258 197422 366494
rect 197186 359258 197422 359494
rect 197186 352258 197422 352494
rect 197186 345258 197422 345494
rect 197186 338258 197422 338494
rect 197186 331258 197422 331494
rect 197186 324258 197422 324494
rect 197186 317258 197422 317494
rect 197186 310258 197422 310494
rect 197186 303258 197422 303494
rect 197186 296258 197422 296494
rect 197186 289258 197422 289494
rect 197186 282258 197422 282494
rect 197186 275258 197422 275494
rect 197186 268258 197422 268494
rect 197186 261258 197422 261494
rect 197186 254258 197422 254494
rect 197186 247258 197422 247494
rect 197186 240258 197422 240494
rect 197186 233258 197422 233494
rect 197186 226258 197422 226494
rect 197186 219258 197422 219494
rect 197186 212258 197422 212494
rect 197186 205258 197422 205494
rect 197186 198258 197422 198494
rect 197186 191258 197422 191494
rect 197186 184258 197422 184494
rect 197186 177258 197422 177494
rect 197186 170258 197422 170494
rect 197186 163258 197422 163494
rect 197186 156258 197422 156494
rect 197186 149258 197422 149494
rect 197186 142258 197422 142494
rect 197186 135258 197422 135494
rect 197186 128258 197422 128494
rect 197186 121258 197422 121494
rect 197186 114258 197422 114494
rect 197186 107258 197422 107494
rect 197186 100258 197422 100494
rect 197186 93258 197422 93494
rect 197186 86258 197422 86494
rect 197186 79258 197422 79494
rect 197186 72258 197422 72494
rect 197186 65258 197422 65494
rect 197186 58258 197422 58494
rect 197186 51258 197422 51494
rect 197186 44258 197422 44494
rect 197186 37258 197422 37494
rect 197186 30258 197422 30494
rect 197186 23258 197422 23494
rect 197186 16258 197422 16494
rect 197186 9258 197422 9494
rect 197186 2258 197422 2494
rect 197186 -982 197422 -746
rect 197186 -1302 197422 -1066
rect 198918 705962 199154 706198
rect 198918 705642 199154 705878
rect 198918 696325 199154 696561
rect 198918 689325 199154 689561
rect 198918 682325 199154 682561
rect 198918 675325 199154 675561
rect 198918 668325 199154 668561
rect 198918 661325 199154 661561
rect 198918 654325 199154 654561
rect 198918 647325 199154 647561
rect 198918 640325 199154 640561
rect 198918 633325 199154 633561
rect 198918 626325 199154 626561
rect 198918 619325 199154 619561
rect 198918 612325 199154 612561
rect 198918 605325 199154 605561
rect 198918 598325 199154 598561
rect 198918 591325 199154 591561
rect 198918 584325 199154 584561
rect 198918 577325 199154 577561
rect 198918 570325 199154 570561
rect 198918 563325 199154 563561
rect 198918 556325 199154 556561
rect 198918 549325 199154 549561
rect 198918 542325 199154 542561
rect 198918 535325 199154 535561
rect 198918 528325 199154 528561
rect 198918 521325 199154 521561
rect 198918 514325 199154 514561
rect 198918 507325 199154 507561
rect 198918 500325 199154 500561
rect 198918 493325 199154 493561
rect 198918 486325 199154 486561
rect 198918 479325 199154 479561
rect 198918 472325 199154 472561
rect 198918 465325 199154 465561
rect 198918 458325 199154 458561
rect 198918 451325 199154 451561
rect 198918 444325 199154 444561
rect 198918 437325 199154 437561
rect 198918 430325 199154 430561
rect 198918 423325 199154 423561
rect 198918 416325 199154 416561
rect 198918 409325 199154 409561
rect 198918 402325 199154 402561
rect 198918 395325 199154 395561
rect 198918 388325 199154 388561
rect 198918 381325 199154 381561
rect 198918 374325 199154 374561
rect 198918 367325 199154 367561
rect 198918 360325 199154 360561
rect 198918 353325 199154 353561
rect 198918 346325 199154 346561
rect 198918 339325 199154 339561
rect 198918 332325 199154 332561
rect 198918 325325 199154 325561
rect 198918 318325 199154 318561
rect 198918 311325 199154 311561
rect 198918 304325 199154 304561
rect 198918 297325 199154 297561
rect 198918 290325 199154 290561
rect 198918 283325 199154 283561
rect 198918 276325 199154 276561
rect 198918 269325 199154 269561
rect 198918 262325 199154 262561
rect 198918 255325 199154 255561
rect 198918 248325 199154 248561
rect 198918 241325 199154 241561
rect 198918 234325 199154 234561
rect 198918 227325 199154 227561
rect 198918 220325 199154 220561
rect 198918 213325 199154 213561
rect 198918 206325 199154 206561
rect 198918 199325 199154 199561
rect 198918 192325 199154 192561
rect 198918 185325 199154 185561
rect 198918 178325 199154 178561
rect 198918 171325 199154 171561
rect 198918 164325 199154 164561
rect 198918 157325 199154 157561
rect 198918 150325 199154 150561
rect 198918 143325 199154 143561
rect 198918 136325 199154 136561
rect 198918 129325 199154 129561
rect 198918 122325 199154 122561
rect 198918 115325 199154 115561
rect 198918 108325 199154 108561
rect 198918 101325 199154 101561
rect 198918 94325 199154 94561
rect 198918 87325 199154 87561
rect 198918 80325 199154 80561
rect 198918 73325 199154 73561
rect 198918 66325 199154 66561
rect 198918 59325 199154 59561
rect 198918 52325 199154 52561
rect 198918 45325 199154 45561
rect 198918 38325 199154 38561
rect 198918 31325 199154 31561
rect 198918 24325 199154 24561
rect 198918 17325 199154 17561
rect 198918 10325 199154 10561
rect 198918 3325 199154 3561
rect 198918 -1942 199154 -1706
rect 198918 -2262 199154 -2026
rect 204186 705002 204422 705238
rect 204186 704682 204422 704918
rect 204186 695258 204422 695494
rect 204186 688258 204422 688494
rect 204186 681258 204422 681494
rect 204186 674258 204422 674494
rect 204186 667258 204422 667494
rect 204186 660258 204422 660494
rect 204186 653258 204422 653494
rect 204186 646258 204422 646494
rect 204186 639258 204422 639494
rect 204186 632258 204422 632494
rect 204186 625258 204422 625494
rect 204186 618258 204422 618494
rect 204186 611258 204422 611494
rect 204186 604258 204422 604494
rect 204186 597258 204422 597494
rect 204186 590258 204422 590494
rect 204186 583258 204422 583494
rect 204186 576258 204422 576494
rect 204186 569258 204422 569494
rect 204186 562258 204422 562494
rect 204186 555258 204422 555494
rect 204186 548258 204422 548494
rect 204186 541258 204422 541494
rect 204186 534258 204422 534494
rect 204186 527258 204422 527494
rect 204186 520258 204422 520494
rect 204186 513258 204422 513494
rect 204186 506258 204422 506494
rect 204186 499258 204422 499494
rect 204186 492258 204422 492494
rect 204186 485258 204422 485494
rect 204186 478258 204422 478494
rect 204186 471258 204422 471494
rect 204186 464258 204422 464494
rect 204186 457258 204422 457494
rect 204186 450258 204422 450494
rect 204186 443258 204422 443494
rect 204186 436258 204422 436494
rect 204186 429258 204422 429494
rect 204186 422258 204422 422494
rect 204186 415258 204422 415494
rect 204186 408258 204422 408494
rect 204186 401258 204422 401494
rect 204186 394258 204422 394494
rect 204186 387258 204422 387494
rect 204186 380258 204422 380494
rect 204186 373258 204422 373494
rect 204186 366258 204422 366494
rect 204186 359258 204422 359494
rect 204186 352258 204422 352494
rect 204186 345258 204422 345494
rect 204186 338258 204422 338494
rect 204186 331258 204422 331494
rect 204186 324258 204422 324494
rect 204186 317258 204422 317494
rect 204186 310258 204422 310494
rect 204186 303258 204422 303494
rect 204186 296258 204422 296494
rect 204186 289258 204422 289494
rect 204186 282258 204422 282494
rect 204186 275258 204422 275494
rect 204186 268258 204422 268494
rect 204186 261258 204422 261494
rect 204186 254258 204422 254494
rect 204186 247258 204422 247494
rect 204186 240258 204422 240494
rect 204186 233258 204422 233494
rect 204186 226258 204422 226494
rect 204186 219258 204422 219494
rect 204186 212258 204422 212494
rect 204186 205258 204422 205494
rect 204186 198258 204422 198494
rect 204186 191258 204422 191494
rect 204186 184258 204422 184494
rect 204186 177258 204422 177494
rect 204186 170258 204422 170494
rect 204186 163258 204422 163494
rect 204186 156258 204422 156494
rect 204186 149258 204422 149494
rect 204186 142258 204422 142494
rect 204186 135258 204422 135494
rect 204186 128258 204422 128494
rect 204186 121258 204422 121494
rect 204186 114258 204422 114494
rect 204186 107258 204422 107494
rect 204186 100258 204422 100494
rect 204186 93258 204422 93494
rect 204186 86258 204422 86494
rect 204186 79258 204422 79494
rect 204186 72258 204422 72494
rect 204186 65258 204422 65494
rect 204186 58258 204422 58494
rect 204186 51258 204422 51494
rect 204186 44258 204422 44494
rect 204186 37258 204422 37494
rect 204186 30258 204422 30494
rect 204186 23258 204422 23494
rect 204186 16258 204422 16494
rect 204186 9258 204422 9494
rect 204186 2258 204422 2494
rect 204186 -982 204422 -746
rect 204186 -1302 204422 -1066
rect 205918 705962 206154 706198
rect 205918 705642 206154 705878
rect 205918 696325 206154 696561
rect 205918 689325 206154 689561
rect 205918 682325 206154 682561
rect 205918 675325 206154 675561
rect 205918 668325 206154 668561
rect 205918 661325 206154 661561
rect 205918 654325 206154 654561
rect 205918 647325 206154 647561
rect 205918 640325 206154 640561
rect 205918 633325 206154 633561
rect 205918 626325 206154 626561
rect 205918 619325 206154 619561
rect 205918 612325 206154 612561
rect 205918 605325 206154 605561
rect 205918 598325 206154 598561
rect 205918 591325 206154 591561
rect 205918 584325 206154 584561
rect 205918 577325 206154 577561
rect 205918 570325 206154 570561
rect 205918 563325 206154 563561
rect 205918 556325 206154 556561
rect 205918 549325 206154 549561
rect 205918 542325 206154 542561
rect 205918 535325 206154 535561
rect 205918 528325 206154 528561
rect 205918 521325 206154 521561
rect 205918 514325 206154 514561
rect 205918 507325 206154 507561
rect 205918 500325 206154 500561
rect 205918 493325 206154 493561
rect 205918 486325 206154 486561
rect 205918 479325 206154 479561
rect 205918 472325 206154 472561
rect 205918 465325 206154 465561
rect 205918 458325 206154 458561
rect 205918 451325 206154 451561
rect 205918 444325 206154 444561
rect 205918 437325 206154 437561
rect 205918 430325 206154 430561
rect 205918 423325 206154 423561
rect 205918 416325 206154 416561
rect 205918 409325 206154 409561
rect 205918 402325 206154 402561
rect 205918 395325 206154 395561
rect 205918 388325 206154 388561
rect 205918 381325 206154 381561
rect 205918 374325 206154 374561
rect 205918 367325 206154 367561
rect 205918 360325 206154 360561
rect 205918 353325 206154 353561
rect 205918 346325 206154 346561
rect 205918 339325 206154 339561
rect 205918 332325 206154 332561
rect 205918 325325 206154 325561
rect 205918 318325 206154 318561
rect 205918 311325 206154 311561
rect 205918 304325 206154 304561
rect 205918 297325 206154 297561
rect 205918 290325 206154 290561
rect 205918 283325 206154 283561
rect 205918 276325 206154 276561
rect 205918 269325 206154 269561
rect 205918 262325 206154 262561
rect 205918 255325 206154 255561
rect 205918 248325 206154 248561
rect 205918 241325 206154 241561
rect 205918 234325 206154 234561
rect 205918 227325 206154 227561
rect 205918 220325 206154 220561
rect 205918 213325 206154 213561
rect 205918 206325 206154 206561
rect 205918 199325 206154 199561
rect 205918 192325 206154 192561
rect 205918 185325 206154 185561
rect 205918 178325 206154 178561
rect 205918 171325 206154 171561
rect 205918 164325 206154 164561
rect 205918 157325 206154 157561
rect 205918 150325 206154 150561
rect 205918 143325 206154 143561
rect 205918 136325 206154 136561
rect 205918 129325 206154 129561
rect 205918 122325 206154 122561
rect 205918 115325 206154 115561
rect 205918 108325 206154 108561
rect 205918 101325 206154 101561
rect 205918 94325 206154 94561
rect 205918 87325 206154 87561
rect 205918 80325 206154 80561
rect 205918 73325 206154 73561
rect 205918 66325 206154 66561
rect 205918 59325 206154 59561
rect 205918 52325 206154 52561
rect 205918 45325 206154 45561
rect 205918 38325 206154 38561
rect 205918 31325 206154 31561
rect 205918 24325 206154 24561
rect 205918 17325 206154 17561
rect 205918 10325 206154 10561
rect 205918 3325 206154 3561
rect 205918 -1942 206154 -1706
rect 205918 -2262 206154 -2026
rect 211186 705002 211422 705238
rect 211186 704682 211422 704918
rect 211186 695258 211422 695494
rect 211186 688258 211422 688494
rect 211186 681258 211422 681494
rect 211186 674258 211422 674494
rect 211186 667258 211422 667494
rect 211186 660258 211422 660494
rect 211186 653258 211422 653494
rect 211186 646258 211422 646494
rect 211186 639258 211422 639494
rect 211186 632258 211422 632494
rect 211186 625258 211422 625494
rect 211186 618258 211422 618494
rect 211186 611258 211422 611494
rect 211186 604258 211422 604494
rect 211186 597258 211422 597494
rect 211186 590258 211422 590494
rect 211186 583258 211422 583494
rect 211186 576258 211422 576494
rect 211186 569258 211422 569494
rect 211186 562258 211422 562494
rect 211186 555258 211422 555494
rect 211186 548258 211422 548494
rect 211186 541258 211422 541494
rect 211186 534258 211422 534494
rect 211186 527258 211422 527494
rect 211186 520258 211422 520494
rect 211186 513258 211422 513494
rect 211186 506258 211422 506494
rect 211186 499258 211422 499494
rect 211186 492258 211422 492494
rect 211186 485258 211422 485494
rect 211186 478258 211422 478494
rect 211186 471258 211422 471494
rect 211186 464258 211422 464494
rect 211186 457258 211422 457494
rect 211186 450258 211422 450494
rect 211186 443258 211422 443494
rect 211186 436258 211422 436494
rect 211186 429258 211422 429494
rect 211186 422258 211422 422494
rect 211186 415258 211422 415494
rect 211186 408258 211422 408494
rect 211186 401258 211422 401494
rect 211186 394258 211422 394494
rect 211186 387258 211422 387494
rect 211186 380258 211422 380494
rect 211186 373258 211422 373494
rect 211186 366258 211422 366494
rect 211186 359258 211422 359494
rect 211186 352258 211422 352494
rect 211186 345258 211422 345494
rect 211186 338258 211422 338494
rect 211186 331258 211422 331494
rect 211186 324258 211422 324494
rect 211186 317258 211422 317494
rect 211186 310258 211422 310494
rect 211186 303258 211422 303494
rect 211186 296258 211422 296494
rect 211186 289258 211422 289494
rect 211186 282258 211422 282494
rect 211186 275258 211422 275494
rect 211186 268258 211422 268494
rect 211186 261258 211422 261494
rect 211186 254258 211422 254494
rect 211186 247258 211422 247494
rect 211186 240258 211422 240494
rect 211186 233258 211422 233494
rect 211186 226258 211422 226494
rect 211186 219258 211422 219494
rect 211186 212258 211422 212494
rect 211186 205258 211422 205494
rect 211186 198258 211422 198494
rect 211186 191258 211422 191494
rect 211186 184258 211422 184494
rect 211186 177258 211422 177494
rect 211186 170258 211422 170494
rect 211186 163258 211422 163494
rect 211186 156258 211422 156494
rect 211186 149258 211422 149494
rect 211186 142258 211422 142494
rect 211186 135258 211422 135494
rect 211186 128258 211422 128494
rect 211186 121258 211422 121494
rect 211186 114258 211422 114494
rect 211186 107258 211422 107494
rect 211186 100258 211422 100494
rect 211186 93258 211422 93494
rect 211186 86258 211422 86494
rect 211186 79258 211422 79494
rect 211186 72258 211422 72494
rect 211186 65258 211422 65494
rect 211186 58258 211422 58494
rect 211186 51258 211422 51494
rect 211186 44258 211422 44494
rect 211186 37258 211422 37494
rect 211186 30258 211422 30494
rect 211186 23258 211422 23494
rect 211186 16258 211422 16494
rect 211186 9258 211422 9494
rect 211186 2258 211422 2494
rect 211186 -982 211422 -746
rect 211186 -1302 211422 -1066
rect 212918 705962 213154 706198
rect 212918 705642 213154 705878
rect 212918 696325 213154 696561
rect 212918 689325 213154 689561
rect 212918 682325 213154 682561
rect 212918 675325 213154 675561
rect 212918 668325 213154 668561
rect 212918 661325 213154 661561
rect 212918 654325 213154 654561
rect 212918 647325 213154 647561
rect 212918 640325 213154 640561
rect 212918 633325 213154 633561
rect 212918 626325 213154 626561
rect 212918 619325 213154 619561
rect 212918 612325 213154 612561
rect 212918 605325 213154 605561
rect 212918 598325 213154 598561
rect 212918 591325 213154 591561
rect 212918 584325 213154 584561
rect 212918 577325 213154 577561
rect 212918 570325 213154 570561
rect 212918 563325 213154 563561
rect 212918 556325 213154 556561
rect 212918 549325 213154 549561
rect 212918 542325 213154 542561
rect 212918 535325 213154 535561
rect 212918 528325 213154 528561
rect 212918 521325 213154 521561
rect 212918 514325 213154 514561
rect 212918 507325 213154 507561
rect 212918 500325 213154 500561
rect 212918 493325 213154 493561
rect 212918 486325 213154 486561
rect 212918 479325 213154 479561
rect 212918 472325 213154 472561
rect 212918 465325 213154 465561
rect 212918 458325 213154 458561
rect 212918 451325 213154 451561
rect 212918 444325 213154 444561
rect 212918 437325 213154 437561
rect 212918 430325 213154 430561
rect 212918 423325 213154 423561
rect 212918 416325 213154 416561
rect 212918 409325 213154 409561
rect 212918 402325 213154 402561
rect 212918 395325 213154 395561
rect 212918 388325 213154 388561
rect 212918 381325 213154 381561
rect 212918 374325 213154 374561
rect 212918 367325 213154 367561
rect 212918 360325 213154 360561
rect 212918 353325 213154 353561
rect 212918 346325 213154 346561
rect 212918 339325 213154 339561
rect 212918 332325 213154 332561
rect 212918 325325 213154 325561
rect 212918 318325 213154 318561
rect 212918 311325 213154 311561
rect 212918 304325 213154 304561
rect 212918 297325 213154 297561
rect 212918 290325 213154 290561
rect 212918 283325 213154 283561
rect 212918 276325 213154 276561
rect 212918 269325 213154 269561
rect 212918 262325 213154 262561
rect 212918 255325 213154 255561
rect 212918 248325 213154 248561
rect 212918 241325 213154 241561
rect 212918 234325 213154 234561
rect 212918 227325 213154 227561
rect 212918 220325 213154 220561
rect 212918 213325 213154 213561
rect 212918 206325 213154 206561
rect 212918 199325 213154 199561
rect 212918 192325 213154 192561
rect 212918 185325 213154 185561
rect 212918 178325 213154 178561
rect 212918 171325 213154 171561
rect 212918 164325 213154 164561
rect 212918 157325 213154 157561
rect 212918 150325 213154 150561
rect 212918 143325 213154 143561
rect 212918 136325 213154 136561
rect 212918 129325 213154 129561
rect 212918 122325 213154 122561
rect 212918 115325 213154 115561
rect 212918 108325 213154 108561
rect 212918 101325 213154 101561
rect 212918 94325 213154 94561
rect 212918 87325 213154 87561
rect 212918 80325 213154 80561
rect 212918 73325 213154 73561
rect 212918 66325 213154 66561
rect 212918 59325 213154 59561
rect 212918 52325 213154 52561
rect 212918 45325 213154 45561
rect 212918 38325 213154 38561
rect 212918 31325 213154 31561
rect 212918 24325 213154 24561
rect 212918 17325 213154 17561
rect 212918 10325 213154 10561
rect 212918 3325 213154 3561
rect 212918 -1942 213154 -1706
rect 212918 -2262 213154 -2026
rect 218186 705002 218422 705238
rect 218186 704682 218422 704918
rect 218186 695258 218422 695494
rect 218186 688258 218422 688494
rect 218186 681258 218422 681494
rect 218186 674258 218422 674494
rect 218186 667258 218422 667494
rect 218186 660258 218422 660494
rect 218186 653258 218422 653494
rect 218186 646258 218422 646494
rect 218186 639258 218422 639494
rect 218186 632258 218422 632494
rect 218186 625258 218422 625494
rect 218186 618258 218422 618494
rect 218186 611258 218422 611494
rect 218186 604258 218422 604494
rect 218186 597258 218422 597494
rect 218186 590258 218422 590494
rect 218186 583258 218422 583494
rect 218186 576258 218422 576494
rect 218186 569258 218422 569494
rect 218186 562258 218422 562494
rect 218186 555258 218422 555494
rect 218186 548258 218422 548494
rect 218186 541258 218422 541494
rect 218186 534258 218422 534494
rect 218186 527258 218422 527494
rect 218186 520258 218422 520494
rect 218186 513258 218422 513494
rect 218186 506258 218422 506494
rect 218186 499258 218422 499494
rect 218186 492258 218422 492494
rect 218186 485258 218422 485494
rect 218186 478258 218422 478494
rect 218186 471258 218422 471494
rect 218186 464258 218422 464494
rect 218186 457258 218422 457494
rect 218186 450258 218422 450494
rect 218186 443258 218422 443494
rect 218186 436258 218422 436494
rect 218186 429258 218422 429494
rect 218186 422258 218422 422494
rect 218186 415258 218422 415494
rect 218186 408258 218422 408494
rect 218186 401258 218422 401494
rect 218186 394258 218422 394494
rect 218186 387258 218422 387494
rect 218186 380258 218422 380494
rect 218186 373258 218422 373494
rect 218186 366258 218422 366494
rect 218186 359258 218422 359494
rect 218186 352258 218422 352494
rect 218186 345258 218422 345494
rect 218186 338258 218422 338494
rect 218186 331258 218422 331494
rect 218186 324258 218422 324494
rect 218186 317258 218422 317494
rect 218186 310258 218422 310494
rect 218186 303258 218422 303494
rect 218186 296258 218422 296494
rect 218186 289258 218422 289494
rect 218186 282258 218422 282494
rect 218186 275258 218422 275494
rect 218186 268258 218422 268494
rect 218186 261258 218422 261494
rect 218186 254258 218422 254494
rect 218186 247258 218422 247494
rect 218186 240258 218422 240494
rect 218186 233258 218422 233494
rect 218186 226258 218422 226494
rect 218186 219258 218422 219494
rect 218186 212258 218422 212494
rect 218186 205258 218422 205494
rect 218186 198258 218422 198494
rect 218186 191258 218422 191494
rect 218186 184258 218422 184494
rect 218186 177258 218422 177494
rect 218186 170258 218422 170494
rect 218186 163258 218422 163494
rect 218186 156258 218422 156494
rect 218186 149258 218422 149494
rect 218186 142258 218422 142494
rect 218186 135258 218422 135494
rect 218186 128258 218422 128494
rect 218186 121258 218422 121494
rect 218186 114258 218422 114494
rect 218186 107258 218422 107494
rect 218186 100258 218422 100494
rect 218186 93258 218422 93494
rect 218186 86258 218422 86494
rect 218186 79258 218422 79494
rect 218186 72258 218422 72494
rect 218186 65258 218422 65494
rect 218186 58258 218422 58494
rect 218186 51258 218422 51494
rect 218186 44258 218422 44494
rect 218186 37258 218422 37494
rect 218186 30258 218422 30494
rect 218186 23258 218422 23494
rect 218186 16258 218422 16494
rect 218186 9258 218422 9494
rect 218186 2258 218422 2494
rect 218186 -982 218422 -746
rect 218186 -1302 218422 -1066
rect 219918 705962 220154 706198
rect 219918 705642 220154 705878
rect 219918 696325 220154 696561
rect 219918 689325 220154 689561
rect 219918 682325 220154 682561
rect 219918 675325 220154 675561
rect 219918 668325 220154 668561
rect 219918 661325 220154 661561
rect 219918 654325 220154 654561
rect 219918 647325 220154 647561
rect 219918 640325 220154 640561
rect 219918 633325 220154 633561
rect 219918 626325 220154 626561
rect 219918 619325 220154 619561
rect 219918 612325 220154 612561
rect 219918 605325 220154 605561
rect 219918 598325 220154 598561
rect 219918 591325 220154 591561
rect 219918 584325 220154 584561
rect 219918 577325 220154 577561
rect 219918 570325 220154 570561
rect 219918 563325 220154 563561
rect 219918 556325 220154 556561
rect 219918 549325 220154 549561
rect 219918 542325 220154 542561
rect 219918 535325 220154 535561
rect 219918 528325 220154 528561
rect 219918 521325 220154 521561
rect 219918 514325 220154 514561
rect 219918 507325 220154 507561
rect 219918 500325 220154 500561
rect 219918 493325 220154 493561
rect 219918 486325 220154 486561
rect 219918 479325 220154 479561
rect 219918 472325 220154 472561
rect 219918 465325 220154 465561
rect 219918 458325 220154 458561
rect 219918 451325 220154 451561
rect 219918 444325 220154 444561
rect 219918 437325 220154 437561
rect 219918 430325 220154 430561
rect 219918 423325 220154 423561
rect 219918 416325 220154 416561
rect 219918 409325 220154 409561
rect 219918 402325 220154 402561
rect 219918 395325 220154 395561
rect 219918 388325 220154 388561
rect 219918 381325 220154 381561
rect 219918 374325 220154 374561
rect 219918 367325 220154 367561
rect 219918 360325 220154 360561
rect 219918 353325 220154 353561
rect 219918 346325 220154 346561
rect 219918 339325 220154 339561
rect 219918 332325 220154 332561
rect 219918 325325 220154 325561
rect 219918 318325 220154 318561
rect 219918 311325 220154 311561
rect 219918 304325 220154 304561
rect 219918 297325 220154 297561
rect 219918 290325 220154 290561
rect 219918 283325 220154 283561
rect 219918 276325 220154 276561
rect 219918 269325 220154 269561
rect 219918 262325 220154 262561
rect 219918 255325 220154 255561
rect 219918 248325 220154 248561
rect 219918 241325 220154 241561
rect 219918 234325 220154 234561
rect 219918 227325 220154 227561
rect 219918 220325 220154 220561
rect 219918 213325 220154 213561
rect 219918 206325 220154 206561
rect 219918 199325 220154 199561
rect 219918 192325 220154 192561
rect 219918 185325 220154 185561
rect 219918 178325 220154 178561
rect 219918 171325 220154 171561
rect 219918 164325 220154 164561
rect 219918 157325 220154 157561
rect 219918 150325 220154 150561
rect 219918 143325 220154 143561
rect 219918 136325 220154 136561
rect 219918 129325 220154 129561
rect 219918 122325 220154 122561
rect 219918 115325 220154 115561
rect 219918 108325 220154 108561
rect 219918 101325 220154 101561
rect 219918 94325 220154 94561
rect 219918 87325 220154 87561
rect 219918 80325 220154 80561
rect 219918 73325 220154 73561
rect 219918 66325 220154 66561
rect 219918 59325 220154 59561
rect 219918 52325 220154 52561
rect 219918 45325 220154 45561
rect 219918 38325 220154 38561
rect 219918 31325 220154 31561
rect 219918 24325 220154 24561
rect 219918 17325 220154 17561
rect 219918 10325 220154 10561
rect 219918 3325 220154 3561
rect 219918 -1942 220154 -1706
rect 219918 -2262 220154 -2026
rect 225186 705002 225422 705238
rect 225186 704682 225422 704918
rect 225186 695258 225422 695494
rect 225186 688258 225422 688494
rect 225186 681258 225422 681494
rect 225186 674258 225422 674494
rect 225186 667258 225422 667494
rect 225186 660258 225422 660494
rect 225186 653258 225422 653494
rect 225186 646258 225422 646494
rect 225186 639258 225422 639494
rect 225186 632258 225422 632494
rect 225186 625258 225422 625494
rect 225186 618258 225422 618494
rect 225186 611258 225422 611494
rect 225186 604258 225422 604494
rect 225186 597258 225422 597494
rect 225186 590258 225422 590494
rect 225186 583258 225422 583494
rect 225186 576258 225422 576494
rect 225186 569258 225422 569494
rect 225186 562258 225422 562494
rect 225186 555258 225422 555494
rect 225186 548258 225422 548494
rect 225186 541258 225422 541494
rect 225186 534258 225422 534494
rect 225186 527258 225422 527494
rect 225186 520258 225422 520494
rect 225186 513258 225422 513494
rect 225186 506258 225422 506494
rect 225186 499258 225422 499494
rect 225186 492258 225422 492494
rect 225186 485258 225422 485494
rect 225186 478258 225422 478494
rect 225186 471258 225422 471494
rect 225186 464258 225422 464494
rect 225186 457258 225422 457494
rect 225186 450258 225422 450494
rect 225186 443258 225422 443494
rect 225186 436258 225422 436494
rect 225186 429258 225422 429494
rect 225186 422258 225422 422494
rect 225186 415258 225422 415494
rect 225186 408258 225422 408494
rect 225186 401258 225422 401494
rect 225186 394258 225422 394494
rect 225186 387258 225422 387494
rect 225186 380258 225422 380494
rect 225186 373258 225422 373494
rect 225186 366258 225422 366494
rect 225186 359258 225422 359494
rect 225186 352258 225422 352494
rect 225186 345258 225422 345494
rect 225186 338258 225422 338494
rect 225186 331258 225422 331494
rect 225186 324258 225422 324494
rect 225186 317258 225422 317494
rect 225186 310258 225422 310494
rect 225186 303258 225422 303494
rect 225186 296258 225422 296494
rect 225186 289258 225422 289494
rect 225186 282258 225422 282494
rect 225186 275258 225422 275494
rect 225186 268258 225422 268494
rect 225186 261258 225422 261494
rect 225186 254258 225422 254494
rect 225186 247258 225422 247494
rect 225186 240258 225422 240494
rect 225186 233258 225422 233494
rect 225186 226258 225422 226494
rect 225186 219258 225422 219494
rect 225186 212258 225422 212494
rect 225186 205258 225422 205494
rect 225186 198258 225422 198494
rect 225186 191258 225422 191494
rect 225186 184258 225422 184494
rect 225186 177258 225422 177494
rect 225186 170258 225422 170494
rect 225186 163258 225422 163494
rect 225186 156258 225422 156494
rect 225186 149258 225422 149494
rect 225186 142258 225422 142494
rect 225186 135258 225422 135494
rect 225186 128258 225422 128494
rect 225186 121258 225422 121494
rect 225186 114258 225422 114494
rect 225186 107258 225422 107494
rect 225186 100258 225422 100494
rect 225186 93258 225422 93494
rect 225186 86258 225422 86494
rect 225186 79258 225422 79494
rect 225186 72258 225422 72494
rect 225186 65258 225422 65494
rect 225186 58258 225422 58494
rect 225186 51258 225422 51494
rect 225186 44258 225422 44494
rect 225186 37258 225422 37494
rect 225186 30258 225422 30494
rect 225186 23258 225422 23494
rect 225186 16258 225422 16494
rect 225186 9258 225422 9494
rect 225186 2258 225422 2494
rect 225186 -982 225422 -746
rect 225186 -1302 225422 -1066
rect 226918 705962 227154 706198
rect 226918 705642 227154 705878
rect 226918 696325 227154 696561
rect 226918 689325 227154 689561
rect 226918 682325 227154 682561
rect 226918 675325 227154 675561
rect 226918 668325 227154 668561
rect 226918 661325 227154 661561
rect 226918 654325 227154 654561
rect 226918 647325 227154 647561
rect 226918 640325 227154 640561
rect 226918 633325 227154 633561
rect 226918 626325 227154 626561
rect 226918 619325 227154 619561
rect 226918 612325 227154 612561
rect 226918 605325 227154 605561
rect 226918 598325 227154 598561
rect 226918 591325 227154 591561
rect 226918 584325 227154 584561
rect 226918 577325 227154 577561
rect 226918 570325 227154 570561
rect 226918 563325 227154 563561
rect 226918 556325 227154 556561
rect 226918 549325 227154 549561
rect 226918 542325 227154 542561
rect 226918 535325 227154 535561
rect 226918 528325 227154 528561
rect 226918 521325 227154 521561
rect 226918 514325 227154 514561
rect 226918 507325 227154 507561
rect 226918 500325 227154 500561
rect 226918 493325 227154 493561
rect 226918 486325 227154 486561
rect 226918 479325 227154 479561
rect 226918 472325 227154 472561
rect 226918 465325 227154 465561
rect 226918 458325 227154 458561
rect 226918 451325 227154 451561
rect 226918 444325 227154 444561
rect 226918 437325 227154 437561
rect 226918 430325 227154 430561
rect 226918 423325 227154 423561
rect 226918 416325 227154 416561
rect 226918 409325 227154 409561
rect 226918 402325 227154 402561
rect 226918 395325 227154 395561
rect 226918 388325 227154 388561
rect 226918 381325 227154 381561
rect 226918 374325 227154 374561
rect 226918 367325 227154 367561
rect 226918 360325 227154 360561
rect 226918 353325 227154 353561
rect 226918 346325 227154 346561
rect 226918 339325 227154 339561
rect 226918 332325 227154 332561
rect 226918 325325 227154 325561
rect 226918 318325 227154 318561
rect 226918 311325 227154 311561
rect 226918 304325 227154 304561
rect 226918 297325 227154 297561
rect 226918 290325 227154 290561
rect 226918 283325 227154 283561
rect 226918 276325 227154 276561
rect 226918 269325 227154 269561
rect 226918 262325 227154 262561
rect 226918 255325 227154 255561
rect 226918 248325 227154 248561
rect 226918 241325 227154 241561
rect 226918 234325 227154 234561
rect 226918 227325 227154 227561
rect 226918 220325 227154 220561
rect 226918 213325 227154 213561
rect 226918 206325 227154 206561
rect 226918 199325 227154 199561
rect 226918 192325 227154 192561
rect 226918 185325 227154 185561
rect 226918 178325 227154 178561
rect 226918 171325 227154 171561
rect 226918 164325 227154 164561
rect 226918 157325 227154 157561
rect 226918 150325 227154 150561
rect 226918 143325 227154 143561
rect 226918 136325 227154 136561
rect 226918 129325 227154 129561
rect 226918 122325 227154 122561
rect 226918 115325 227154 115561
rect 226918 108325 227154 108561
rect 226918 101325 227154 101561
rect 226918 94325 227154 94561
rect 226918 87325 227154 87561
rect 226918 80325 227154 80561
rect 226918 73325 227154 73561
rect 226918 66325 227154 66561
rect 226918 59325 227154 59561
rect 226918 52325 227154 52561
rect 226918 45325 227154 45561
rect 226918 38325 227154 38561
rect 226918 31325 227154 31561
rect 226918 24325 227154 24561
rect 226918 17325 227154 17561
rect 226918 10325 227154 10561
rect 226918 3325 227154 3561
rect 226918 -1942 227154 -1706
rect 226918 -2262 227154 -2026
rect 232186 705002 232422 705238
rect 232186 704682 232422 704918
rect 232186 695258 232422 695494
rect 232186 688258 232422 688494
rect 232186 681258 232422 681494
rect 232186 674258 232422 674494
rect 232186 667258 232422 667494
rect 232186 660258 232422 660494
rect 232186 653258 232422 653494
rect 232186 646258 232422 646494
rect 232186 639258 232422 639494
rect 232186 632258 232422 632494
rect 232186 625258 232422 625494
rect 232186 618258 232422 618494
rect 232186 611258 232422 611494
rect 232186 604258 232422 604494
rect 232186 597258 232422 597494
rect 232186 590258 232422 590494
rect 232186 583258 232422 583494
rect 232186 576258 232422 576494
rect 232186 569258 232422 569494
rect 232186 562258 232422 562494
rect 232186 555258 232422 555494
rect 232186 548258 232422 548494
rect 232186 541258 232422 541494
rect 232186 534258 232422 534494
rect 232186 527258 232422 527494
rect 232186 520258 232422 520494
rect 232186 513258 232422 513494
rect 232186 506258 232422 506494
rect 232186 499258 232422 499494
rect 232186 492258 232422 492494
rect 232186 485258 232422 485494
rect 232186 478258 232422 478494
rect 232186 471258 232422 471494
rect 232186 464258 232422 464494
rect 232186 457258 232422 457494
rect 232186 450258 232422 450494
rect 232186 443258 232422 443494
rect 232186 436258 232422 436494
rect 232186 429258 232422 429494
rect 232186 422258 232422 422494
rect 232186 415258 232422 415494
rect 232186 408258 232422 408494
rect 232186 401258 232422 401494
rect 232186 394258 232422 394494
rect 232186 387258 232422 387494
rect 232186 380258 232422 380494
rect 232186 373258 232422 373494
rect 232186 366258 232422 366494
rect 232186 359258 232422 359494
rect 232186 352258 232422 352494
rect 232186 345258 232422 345494
rect 232186 338258 232422 338494
rect 232186 331258 232422 331494
rect 232186 324258 232422 324494
rect 232186 317258 232422 317494
rect 232186 310258 232422 310494
rect 232186 303258 232422 303494
rect 232186 296258 232422 296494
rect 232186 289258 232422 289494
rect 232186 282258 232422 282494
rect 232186 275258 232422 275494
rect 232186 268258 232422 268494
rect 232186 261258 232422 261494
rect 232186 254258 232422 254494
rect 232186 247258 232422 247494
rect 232186 240258 232422 240494
rect 232186 233258 232422 233494
rect 232186 226258 232422 226494
rect 232186 219258 232422 219494
rect 232186 212258 232422 212494
rect 232186 205258 232422 205494
rect 232186 198258 232422 198494
rect 232186 191258 232422 191494
rect 232186 184258 232422 184494
rect 232186 177258 232422 177494
rect 232186 170258 232422 170494
rect 232186 163258 232422 163494
rect 232186 156258 232422 156494
rect 232186 149258 232422 149494
rect 232186 142258 232422 142494
rect 232186 135258 232422 135494
rect 232186 128258 232422 128494
rect 232186 121258 232422 121494
rect 232186 114258 232422 114494
rect 232186 107258 232422 107494
rect 232186 100258 232422 100494
rect 232186 93258 232422 93494
rect 232186 86258 232422 86494
rect 232186 79258 232422 79494
rect 232186 72258 232422 72494
rect 232186 65258 232422 65494
rect 232186 58258 232422 58494
rect 232186 51258 232422 51494
rect 232186 44258 232422 44494
rect 232186 37258 232422 37494
rect 232186 30258 232422 30494
rect 232186 23258 232422 23494
rect 232186 16258 232422 16494
rect 232186 9258 232422 9494
rect 232186 2258 232422 2494
rect 232186 -982 232422 -746
rect 232186 -1302 232422 -1066
rect 233918 705962 234154 706198
rect 233918 705642 234154 705878
rect 233918 696325 234154 696561
rect 233918 689325 234154 689561
rect 233918 682325 234154 682561
rect 233918 675325 234154 675561
rect 233918 668325 234154 668561
rect 233918 661325 234154 661561
rect 233918 654325 234154 654561
rect 233918 647325 234154 647561
rect 233918 640325 234154 640561
rect 233918 633325 234154 633561
rect 233918 626325 234154 626561
rect 233918 619325 234154 619561
rect 233918 612325 234154 612561
rect 233918 605325 234154 605561
rect 233918 598325 234154 598561
rect 233918 591325 234154 591561
rect 233918 584325 234154 584561
rect 233918 577325 234154 577561
rect 233918 570325 234154 570561
rect 233918 563325 234154 563561
rect 233918 556325 234154 556561
rect 233918 549325 234154 549561
rect 233918 542325 234154 542561
rect 233918 535325 234154 535561
rect 233918 528325 234154 528561
rect 233918 521325 234154 521561
rect 233918 514325 234154 514561
rect 233918 507325 234154 507561
rect 233918 500325 234154 500561
rect 233918 493325 234154 493561
rect 233918 486325 234154 486561
rect 233918 479325 234154 479561
rect 233918 472325 234154 472561
rect 233918 465325 234154 465561
rect 233918 458325 234154 458561
rect 233918 451325 234154 451561
rect 233918 444325 234154 444561
rect 233918 437325 234154 437561
rect 233918 430325 234154 430561
rect 233918 423325 234154 423561
rect 233918 416325 234154 416561
rect 233918 409325 234154 409561
rect 233918 402325 234154 402561
rect 233918 395325 234154 395561
rect 233918 388325 234154 388561
rect 233918 381325 234154 381561
rect 233918 374325 234154 374561
rect 233918 367325 234154 367561
rect 233918 360325 234154 360561
rect 233918 353325 234154 353561
rect 233918 346325 234154 346561
rect 233918 339325 234154 339561
rect 233918 332325 234154 332561
rect 233918 325325 234154 325561
rect 233918 318325 234154 318561
rect 233918 311325 234154 311561
rect 233918 304325 234154 304561
rect 233918 297325 234154 297561
rect 233918 290325 234154 290561
rect 233918 283325 234154 283561
rect 233918 276325 234154 276561
rect 233918 269325 234154 269561
rect 233918 262325 234154 262561
rect 233918 255325 234154 255561
rect 233918 248325 234154 248561
rect 233918 241325 234154 241561
rect 233918 234325 234154 234561
rect 233918 227325 234154 227561
rect 233918 220325 234154 220561
rect 233918 213325 234154 213561
rect 233918 206325 234154 206561
rect 233918 199325 234154 199561
rect 233918 192325 234154 192561
rect 233918 185325 234154 185561
rect 233918 178325 234154 178561
rect 233918 171325 234154 171561
rect 233918 164325 234154 164561
rect 233918 157325 234154 157561
rect 233918 150325 234154 150561
rect 233918 143325 234154 143561
rect 233918 136325 234154 136561
rect 233918 129325 234154 129561
rect 233918 122325 234154 122561
rect 233918 115325 234154 115561
rect 233918 108325 234154 108561
rect 233918 101325 234154 101561
rect 233918 94325 234154 94561
rect 233918 87325 234154 87561
rect 233918 80325 234154 80561
rect 233918 73325 234154 73561
rect 233918 66325 234154 66561
rect 233918 59325 234154 59561
rect 233918 52325 234154 52561
rect 233918 45325 234154 45561
rect 233918 38325 234154 38561
rect 233918 31325 234154 31561
rect 233918 24325 234154 24561
rect 233918 17325 234154 17561
rect 233918 10325 234154 10561
rect 233918 3325 234154 3561
rect 233918 -1942 234154 -1706
rect 233918 -2262 234154 -2026
rect 239186 705002 239422 705238
rect 239186 704682 239422 704918
rect 239186 695258 239422 695494
rect 239186 688258 239422 688494
rect 239186 681258 239422 681494
rect 239186 674258 239422 674494
rect 239186 667258 239422 667494
rect 239186 660258 239422 660494
rect 239186 653258 239422 653494
rect 239186 646258 239422 646494
rect 239186 639258 239422 639494
rect 239186 632258 239422 632494
rect 239186 625258 239422 625494
rect 239186 618258 239422 618494
rect 239186 611258 239422 611494
rect 239186 604258 239422 604494
rect 239186 597258 239422 597494
rect 239186 590258 239422 590494
rect 239186 583258 239422 583494
rect 239186 576258 239422 576494
rect 239186 569258 239422 569494
rect 239186 562258 239422 562494
rect 239186 555258 239422 555494
rect 239186 548258 239422 548494
rect 239186 541258 239422 541494
rect 239186 534258 239422 534494
rect 239186 527258 239422 527494
rect 239186 520258 239422 520494
rect 239186 513258 239422 513494
rect 239186 506258 239422 506494
rect 239186 499258 239422 499494
rect 239186 492258 239422 492494
rect 239186 485258 239422 485494
rect 239186 478258 239422 478494
rect 239186 471258 239422 471494
rect 239186 464258 239422 464494
rect 239186 457258 239422 457494
rect 239186 450258 239422 450494
rect 239186 443258 239422 443494
rect 239186 436258 239422 436494
rect 239186 429258 239422 429494
rect 239186 422258 239422 422494
rect 239186 415258 239422 415494
rect 239186 408258 239422 408494
rect 239186 401258 239422 401494
rect 239186 394258 239422 394494
rect 239186 387258 239422 387494
rect 239186 380258 239422 380494
rect 239186 373258 239422 373494
rect 239186 366258 239422 366494
rect 239186 359258 239422 359494
rect 239186 352258 239422 352494
rect 239186 345258 239422 345494
rect 239186 338258 239422 338494
rect 239186 331258 239422 331494
rect 239186 324258 239422 324494
rect 239186 317258 239422 317494
rect 239186 310258 239422 310494
rect 239186 303258 239422 303494
rect 239186 296258 239422 296494
rect 239186 289258 239422 289494
rect 239186 282258 239422 282494
rect 239186 275258 239422 275494
rect 239186 268258 239422 268494
rect 239186 261258 239422 261494
rect 239186 254258 239422 254494
rect 239186 247258 239422 247494
rect 239186 240258 239422 240494
rect 239186 233258 239422 233494
rect 239186 226258 239422 226494
rect 239186 219258 239422 219494
rect 239186 212258 239422 212494
rect 239186 205258 239422 205494
rect 239186 198258 239422 198494
rect 239186 191258 239422 191494
rect 239186 184258 239422 184494
rect 239186 177258 239422 177494
rect 239186 170258 239422 170494
rect 239186 163258 239422 163494
rect 239186 156258 239422 156494
rect 239186 149258 239422 149494
rect 239186 142258 239422 142494
rect 239186 135258 239422 135494
rect 239186 128258 239422 128494
rect 239186 121258 239422 121494
rect 239186 114258 239422 114494
rect 239186 107258 239422 107494
rect 239186 100258 239422 100494
rect 239186 93258 239422 93494
rect 239186 86258 239422 86494
rect 239186 79258 239422 79494
rect 239186 72258 239422 72494
rect 239186 65258 239422 65494
rect 239186 58258 239422 58494
rect 239186 51258 239422 51494
rect 239186 44258 239422 44494
rect 239186 37258 239422 37494
rect 239186 30258 239422 30494
rect 239186 23258 239422 23494
rect 239186 16258 239422 16494
rect 239186 9258 239422 9494
rect 239186 2258 239422 2494
rect 239186 -982 239422 -746
rect 239186 -1302 239422 -1066
rect 240918 705962 241154 706198
rect 240918 705642 241154 705878
rect 240918 696325 241154 696561
rect 240918 689325 241154 689561
rect 240918 682325 241154 682561
rect 240918 675325 241154 675561
rect 240918 668325 241154 668561
rect 240918 661325 241154 661561
rect 240918 654325 241154 654561
rect 240918 647325 241154 647561
rect 240918 640325 241154 640561
rect 240918 633325 241154 633561
rect 240918 626325 241154 626561
rect 240918 619325 241154 619561
rect 240918 612325 241154 612561
rect 240918 605325 241154 605561
rect 240918 598325 241154 598561
rect 240918 591325 241154 591561
rect 240918 584325 241154 584561
rect 240918 577325 241154 577561
rect 240918 570325 241154 570561
rect 240918 563325 241154 563561
rect 240918 556325 241154 556561
rect 240918 549325 241154 549561
rect 240918 542325 241154 542561
rect 240918 535325 241154 535561
rect 240918 528325 241154 528561
rect 240918 521325 241154 521561
rect 240918 514325 241154 514561
rect 240918 507325 241154 507561
rect 240918 500325 241154 500561
rect 240918 493325 241154 493561
rect 240918 486325 241154 486561
rect 240918 479325 241154 479561
rect 240918 472325 241154 472561
rect 240918 465325 241154 465561
rect 240918 458325 241154 458561
rect 240918 451325 241154 451561
rect 240918 444325 241154 444561
rect 240918 437325 241154 437561
rect 240918 430325 241154 430561
rect 240918 423325 241154 423561
rect 240918 416325 241154 416561
rect 240918 409325 241154 409561
rect 240918 402325 241154 402561
rect 240918 395325 241154 395561
rect 240918 388325 241154 388561
rect 240918 381325 241154 381561
rect 240918 374325 241154 374561
rect 240918 367325 241154 367561
rect 240918 360325 241154 360561
rect 240918 353325 241154 353561
rect 240918 346325 241154 346561
rect 240918 339325 241154 339561
rect 240918 332325 241154 332561
rect 240918 325325 241154 325561
rect 240918 318325 241154 318561
rect 240918 311325 241154 311561
rect 240918 304325 241154 304561
rect 240918 297325 241154 297561
rect 240918 290325 241154 290561
rect 240918 283325 241154 283561
rect 240918 276325 241154 276561
rect 240918 269325 241154 269561
rect 240918 262325 241154 262561
rect 240918 255325 241154 255561
rect 240918 248325 241154 248561
rect 240918 241325 241154 241561
rect 240918 234325 241154 234561
rect 240918 227325 241154 227561
rect 240918 220325 241154 220561
rect 240918 213325 241154 213561
rect 240918 206325 241154 206561
rect 240918 199325 241154 199561
rect 240918 192325 241154 192561
rect 240918 185325 241154 185561
rect 240918 178325 241154 178561
rect 240918 171325 241154 171561
rect 240918 164325 241154 164561
rect 240918 157325 241154 157561
rect 240918 150325 241154 150561
rect 240918 143325 241154 143561
rect 240918 136325 241154 136561
rect 240918 129325 241154 129561
rect 240918 122325 241154 122561
rect 240918 115325 241154 115561
rect 240918 108325 241154 108561
rect 240918 101325 241154 101561
rect 240918 94325 241154 94561
rect 240918 87325 241154 87561
rect 240918 80325 241154 80561
rect 240918 73325 241154 73561
rect 240918 66325 241154 66561
rect 240918 59325 241154 59561
rect 240918 52325 241154 52561
rect 240918 45325 241154 45561
rect 240918 38325 241154 38561
rect 240918 31325 241154 31561
rect 240918 24325 241154 24561
rect 240918 17325 241154 17561
rect 240918 10325 241154 10561
rect 240918 3325 241154 3561
rect 240918 -1942 241154 -1706
rect 240918 -2262 241154 -2026
rect 246186 705002 246422 705238
rect 246186 704682 246422 704918
rect 246186 695258 246422 695494
rect 246186 688258 246422 688494
rect 246186 681258 246422 681494
rect 246186 674258 246422 674494
rect 246186 667258 246422 667494
rect 246186 660258 246422 660494
rect 246186 653258 246422 653494
rect 246186 646258 246422 646494
rect 246186 639258 246422 639494
rect 246186 632258 246422 632494
rect 246186 625258 246422 625494
rect 246186 618258 246422 618494
rect 246186 611258 246422 611494
rect 246186 604258 246422 604494
rect 246186 597258 246422 597494
rect 246186 590258 246422 590494
rect 246186 583258 246422 583494
rect 246186 576258 246422 576494
rect 246186 569258 246422 569494
rect 246186 562258 246422 562494
rect 246186 555258 246422 555494
rect 246186 548258 246422 548494
rect 246186 541258 246422 541494
rect 246186 534258 246422 534494
rect 246186 527258 246422 527494
rect 246186 520258 246422 520494
rect 246186 513258 246422 513494
rect 246186 506258 246422 506494
rect 246186 499258 246422 499494
rect 246186 492258 246422 492494
rect 246186 485258 246422 485494
rect 246186 478258 246422 478494
rect 246186 471258 246422 471494
rect 246186 464258 246422 464494
rect 246186 457258 246422 457494
rect 246186 450258 246422 450494
rect 246186 443258 246422 443494
rect 246186 436258 246422 436494
rect 246186 429258 246422 429494
rect 246186 422258 246422 422494
rect 246186 415258 246422 415494
rect 246186 408258 246422 408494
rect 246186 401258 246422 401494
rect 246186 394258 246422 394494
rect 246186 387258 246422 387494
rect 246186 380258 246422 380494
rect 246186 373258 246422 373494
rect 246186 366258 246422 366494
rect 246186 359258 246422 359494
rect 246186 352258 246422 352494
rect 246186 345258 246422 345494
rect 246186 338258 246422 338494
rect 246186 331258 246422 331494
rect 246186 324258 246422 324494
rect 246186 317258 246422 317494
rect 246186 310258 246422 310494
rect 246186 303258 246422 303494
rect 246186 296258 246422 296494
rect 246186 289258 246422 289494
rect 246186 282258 246422 282494
rect 246186 275258 246422 275494
rect 246186 268258 246422 268494
rect 246186 261258 246422 261494
rect 246186 254258 246422 254494
rect 246186 247258 246422 247494
rect 246186 240258 246422 240494
rect 246186 233258 246422 233494
rect 246186 226258 246422 226494
rect 246186 219258 246422 219494
rect 246186 212258 246422 212494
rect 246186 205258 246422 205494
rect 246186 198258 246422 198494
rect 246186 191258 246422 191494
rect 246186 184258 246422 184494
rect 246186 177258 246422 177494
rect 246186 170258 246422 170494
rect 246186 163258 246422 163494
rect 246186 156258 246422 156494
rect 246186 149258 246422 149494
rect 246186 142258 246422 142494
rect 246186 135258 246422 135494
rect 246186 128258 246422 128494
rect 246186 121258 246422 121494
rect 246186 114258 246422 114494
rect 246186 107258 246422 107494
rect 246186 100258 246422 100494
rect 246186 93258 246422 93494
rect 246186 86258 246422 86494
rect 246186 79258 246422 79494
rect 246186 72258 246422 72494
rect 246186 65258 246422 65494
rect 246186 58258 246422 58494
rect 246186 51258 246422 51494
rect 246186 44258 246422 44494
rect 246186 37258 246422 37494
rect 246186 30258 246422 30494
rect 246186 23258 246422 23494
rect 246186 16258 246422 16494
rect 246186 9258 246422 9494
rect 246186 2258 246422 2494
rect 246186 -982 246422 -746
rect 246186 -1302 246422 -1066
rect 247918 705962 248154 706198
rect 247918 705642 248154 705878
rect 247918 696325 248154 696561
rect 247918 689325 248154 689561
rect 247918 682325 248154 682561
rect 247918 675325 248154 675561
rect 247918 668325 248154 668561
rect 247918 661325 248154 661561
rect 247918 654325 248154 654561
rect 247918 647325 248154 647561
rect 247918 640325 248154 640561
rect 247918 633325 248154 633561
rect 247918 626325 248154 626561
rect 247918 619325 248154 619561
rect 247918 612325 248154 612561
rect 247918 605325 248154 605561
rect 247918 598325 248154 598561
rect 247918 591325 248154 591561
rect 247918 584325 248154 584561
rect 247918 577325 248154 577561
rect 247918 570325 248154 570561
rect 247918 563325 248154 563561
rect 247918 556325 248154 556561
rect 247918 549325 248154 549561
rect 247918 542325 248154 542561
rect 247918 535325 248154 535561
rect 247918 528325 248154 528561
rect 247918 521325 248154 521561
rect 247918 514325 248154 514561
rect 247918 507325 248154 507561
rect 247918 500325 248154 500561
rect 247918 493325 248154 493561
rect 247918 486325 248154 486561
rect 247918 479325 248154 479561
rect 247918 472325 248154 472561
rect 247918 465325 248154 465561
rect 247918 458325 248154 458561
rect 247918 451325 248154 451561
rect 247918 444325 248154 444561
rect 247918 437325 248154 437561
rect 247918 430325 248154 430561
rect 247918 423325 248154 423561
rect 247918 416325 248154 416561
rect 247918 409325 248154 409561
rect 247918 402325 248154 402561
rect 247918 395325 248154 395561
rect 247918 388325 248154 388561
rect 247918 381325 248154 381561
rect 247918 374325 248154 374561
rect 247918 367325 248154 367561
rect 247918 360325 248154 360561
rect 247918 353325 248154 353561
rect 247918 346325 248154 346561
rect 247918 339325 248154 339561
rect 247918 332325 248154 332561
rect 247918 325325 248154 325561
rect 247918 318325 248154 318561
rect 247918 311325 248154 311561
rect 247918 304325 248154 304561
rect 247918 297325 248154 297561
rect 247918 290325 248154 290561
rect 247918 283325 248154 283561
rect 247918 276325 248154 276561
rect 247918 269325 248154 269561
rect 247918 262325 248154 262561
rect 247918 255325 248154 255561
rect 247918 248325 248154 248561
rect 247918 241325 248154 241561
rect 247918 234325 248154 234561
rect 247918 227325 248154 227561
rect 247918 220325 248154 220561
rect 247918 213325 248154 213561
rect 247918 206325 248154 206561
rect 247918 199325 248154 199561
rect 247918 192325 248154 192561
rect 247918 185325 248154 185561
rect 247918 178325 248154 178561
rect 247918 171325 248154 171561
rect 247918 164325 248154 164561
rect 247918 157325 248154 157561
rect 247918 150325 248154 150561
rect 247918 143325 248154 143561
rect 247918 136325 248154 136561
rect 247918 129325 248154 129561
rect 247918 122325 248154 122561
rect 247918 115325 248154 115561
rect 247918 108325 248154 108561
rect 247918 101325 248154 101561
rect 247918 94325 248154 94561
rect 247918 87325 248154 87561
rect 247918 80325 248154 80561
rect 247918 73325 248154 73561
rect 247918 66325 248154 66561
rect 247918 59325 248154 59561
rect 247918 52325 248154 52561
rect 247918 45325 248154 45561
rect 247918 38325 248154 38561
rect 247918 31325 248154 31561
rect 247918 24325 248154 24561
rect 247918 17325 248154 17561
rect 247918 10325 248154 10561
rect 247918 3325 248154 3561
rect 247918 -1942 248154 -1706
rect 247918 -2262 248154 -2026
rect 253186 705002 253422 705238
rect 253186 704682 253422 704918
rect 253186 695258 253422 695494
rect 253186 688258 253422 688494
rect 253186 681258 253422 681494
rect 253186 674258 253422 674494
rect 253186 667258 253422 667494
rect 253186 660258 253422 660494
rect 253186 653258 253422 653494
rect 253186 646258 253422 646494
rect 253186 639258 253422 639494
rect 253186 632258 253422 632494
rect 253186 625258 253422 625494
rect 253186 618258 253422 618494
rect 253186 611258 253422 611494
rect 253186 604258 253422 604494
rect 253186 597258 253422 597494
rect 253186 590258 253422 590494
rect 253186 583258 253422 583494
rect 253186 576258 253422 576494
rect 253186 569258 253422 569494
rect 253186 562258 253422 562494
rect 253186 555258 253422 555494
rect 253186 548258 253422 548494
rect 253186 541258 253422 541494
rect 253186 534258 253422 534494
rect 253186 527258 253422 527494
rect 253186 520258 253422 520494
rect 253186 513258 253422 513494
rect 253186 506258 253422 506494
rect 253186 499258 253422 499494
rect 253186 492258 253422 492494
rect 253186 485258 253422 485494
rect 253186 478258 253422 478494
rect 253186 471258 253422 471494
rect 253186 464258 253422 464494
rect 253186 457258 253422 457494
rect 253186 450258 253422 450494
rect 253186 443258 253422 443494
rect 253186 436258 253422 436494
rect 253186 429258 253422 429494
rect 253186 422258 253422 422494
rect 253186 415258 253422 415494
rect 253186 408258 253422 408494
rect 253186 401258 253422 401494
rect 253186 394258 253422 394494
rect 253186 387258 253422 387494
rect 253186 380258 253422 380494
rect 253186 373258 253422 373494
rect 253186 366258 253422 366494
rect 253186 359258 253422 359494
rect 253186 352258 253422 352494
rect 253186 345258 253422 345494
rect 253186 338258 253422 338494
rect 253186 331258 253422 331494
rect 253186 324258 253422 324494
rect 253186 317258 253422 317494
rect 253186 310258 253422 310494
rect 253186 303258 253422 303494
rect 253186 296258 253422 296494
rect 253186 289258 253422 289494
rect 253186 282258 253422 282494
rect 253186 275258 253422 275494
rect 253186 268258 253422 268494
rect 253186 261258 253422 261494
rect 253186 254258 253422 254494
rect 253186 247258 253422 247494
rect 253186 240258 253422 240494
rect 253186 233258 253422 233494
rect 253186 226258 253422 226494
rect 253186 219258 253422 219494
rect 253186 212258 253422 212494
rect 253186 205258 253422 205494
rect 253186 198258 253422 198494
rect 253186 191258 253422 191494
rect 253186 184258 253422 184494
rect 253186 177258 253422 177494
rect 253186 170258 253422 170494
rect 253186 163258 253422 163494
rect 253186 156258 253422 156494
rect 253186 149258 253422 149494
rect 253186 142258 253422 142494
rect 253186 135258 253422 135494
rect 253186 128258 253422 128494
rect 253186 121258 253422 121494
rect 253186 114258 253422 114494
rect 253186 107258 253422 107494
rect 253186 100258 253422 100494
rect 253186 93258 253422 93494
rect 253186 86258 253422 86494
rect 253186 79258 253422 79494
rect 253186 72258 253422 72494
rect 253186 65258 253422 65494
rect 253186 58258 253422 58494
rect 253186 51258 253422 51494
rect 253186 44258 253422 44494
rect 253186 37258 253422 37494
rect 253186 30258 253422 30494
rect 253186 23258 253422 23494
rect 253186 16258 253422 16494
rect 253186 9258 253422 9494
rect 253186 2258 253422 2494
rect 253186 -982 253422 -746
rect 253186 -1302 253422 -1066
rect 254918 705962 255154 706198
rect 254918 705642 255154 705878
rect 254918 696325 255154 696561
rect 254918 689325 255154 689561
rect 254918 682325 255154 682561
rect 254918 675325 255154 675561
rect 254918 668325 255154 668561
rect 254918 661325 255154 661561
rect 254918 654325 255154 654561
rect 254918 647325 255154 647561
rect 254918 640325 255154 640561
rect 254918 633325 255154 633561
rect 254918 626325 255154 626561
rect 254918 619325 255154 619561
rect 254918 612325 255154 612561
rect 254918 605325 255154 605561
rect 254918 598325 255154 598561
rect 254918 591325 255154 591561
rect 254918 584325 255154 584561
rect 254918 577325 255154 577561
rect 254918 570325 255154 570561
rect 254918 563325 255154 563561
rect 254918 556325 255154 556561
rect 254918 549325 255154 549561
rect 254918 542325 255154 542561
rect 254918 535325 255154 535561
rect 254918 528325 255154 528561
rect 254918 521325 255154 521561
rect 254918 514325 255154 514561
rect 254918 507325 255154 507561
rect 254918 500325 255154 500561
rect 254918 493325 255154 493561
rect 254918 486325 255154 486561
rect 254918 479325 255154 479561
rect 254918 472325 255154 472561
rect 254918 465325 255154 465561
rect 254918 458325 255154 458561
rect 254918 451325 255154 451561
rect 254918 444325 255154 444561
rect 254918 437325 255154 437561
rect 254918 430325 255154 430561
rect 254918 423325 255154 423561
rect 254918 416325 255154 416561
rect 254918 409325 255154 409561
rect 254918 402325 255154 402561
rect 254918 395325 255154 395561
rect 254918 388325 255154 388561
rect 254918 381325 255154 381561
rect 254918 374325 255154 374561
rect 254918 367325 255154 367561
rect 254918 360325 255154 360561
rect 254918 353325 255154 353561
rect 254918 346325 255154 346561
rect 254918 339325 255154 339561
rect 254918 332325 255154 332561
rect 254918 325325 255154 325561
rect 254918 318325 255154 318561
rect 254918 311325 255154 311561
rect 254918 304325 255154 304561
rect 254918 297325 255154 297561
rect 254918 290325 255154 290561
rect 254918 283325 255154 283561
rect 254918 276325 255154 276561
rect 254918 269325 255154 269561
rect 254918 262325 255154 262561
rect 254918 255325 255154 255561
rect 254918 248325 255154 248561
rect 254918 241325 255154 241561
rect 254918 234325 255154 234561
rect 254918 227325 255154 227561
rect 254918 220325 255154 220561
rect 254918 213325 255154 213561
rect 254918 206325 255154 206561
rect 254918 199325 255154 199561
rect 254918 192325 255154 192561
rect 254918 185325 255154 185561
rect 254918 178325 255154 178561
rect 254918 171325 255154 171561
rect 254918 164325 255154 164561
rect 254918 157325 255154 157561
rect 254918 150325 255154 150561
rect 254918 143325 255154 143561
rect 254918 136325 255154 136561
rect 254918 129325 255154 129561
rect 254918 122325 255154 122561
rect 254918 115325 255154 115561
rect 254918 108325 255154 108561
rect 254918 101325 255154 101561
rect 254918 94325 255154 94561
rect 254918 87325 255154 87561
rect 254918 80325 255154 80561
rect 254918 73325 255154 73561
rect 254918 66325 255154 66561
rect 254918 59325 255154 59561
rect 254918 52325 255154 52561
rect 254918 45325 255154 45561
rect 254918 38325 255154 38561
rect 254918 31325 255154 31561
rect 254918 24325 255154 24561
rect 254918 17325 255154 17561
rect 254918 10325 255154 10561
rect 254918 3325 255154 3561
rect 254918 -1942 255154 -1706
rect 254918 -2262 255154 -2026
rect 260186 705002 260422 705238
rect 260186 704682 260422 704918
rect 260186 695258 260422 695494
rect 260186 688258 260422 688494
rect 260186 681258 260422 681494
rect 260186 674258 260422 674494
rect 260186 667258 260422 667494
rect 260186 660258 260422 660494
rect 260186 653258 260422 653494
rect 260186 646258 260422 646494
rect 260186 639258 260422 639494
rect 260186 632258 260422 632494
rect 260186 625258 260422 625494
rect 260186 618258 260422 618494
rect 260186 611258 260422 611494
rect 260186 604258 260422 604494
rect 260186 597258 260422 597494
rect 260186 590258 260422 590494
rect 260186 583258 260422 583494
rect 260186 576258 260422 576494
rect 260186 569258 260422 569494
rect 260186 562258 260422 562494
rect 260186 555258 260422 555494
rect 260186 548258 260422 548494
rect 260186 541258 260422 541494
rect 260186 534258 260422 534494
rect 260186 527258 260422 527494
rect 260186 520258 260422 520494
rect 260186 513258 260422 513494
rect 260186 506258 260422 506494
rect 260186 499258 260422 499494
rect 260186 492258 260422 492494
rect 260186 485258 260422 485494
rect 260186 478258 260422 478494
rect 260186 471258 260422 471494
rect 260186 464258 260422 464494
rect 260186 457258 260422 457494
rect 260186 450258 260422 450494
rect 260186 443258 260422 443494
rect 260186 436258 260422 436494
rect 260186 429258 260422 429494
rect 260186 422258 260422 422494
rect 260186 415258 260422 415494
rect 260186 408258 260422 408494
rect 260186 401258 260422 401494
rect 260186 394258 260422 394494
rect 260186 387258 260422 387494
rect 260186 380258 260422 380494
rect 260186 373258 260422 373494
rect 260186 366258 260422 366494
rect 260186 359258 260422 359494
rect 260186 352258 260422 352494
rect 260186 345258 260422 345494
rect 260186 338258 260422 338494
rect 260186 331258 260422 331494
rect 260186 324258 260422 324494
rect 260186 317258 260422 317494
rect 260186 310258 260422 310494
rect 260186 303258 260422 303494
rect 260186 296258 260422 296494
rect 260186 289258 260422 289494
rect 260186 282258 260422 282494
rect 260186 275258 260422 275494
rect 260186 268258 260422 268494
rect 260186 261258 260422 261494
rect 260186 254258 260422 254494
rect 260186 247258 260422 247494
rect 260186 240258 260422 240494
rect 260186 233258 260422 233494
rect 260186 226258 260422 226494
rect 260186 219258 260422 219494
rect 260186 212258 260422 212494
rect 260186 205258 260422 205494
rect 260186 198258 260422 198494
rect 260186 191258 260422 191494
rect 260186 184258 260422 184494
rect 260186 177258 260422 177494
rect 260186 170258 260422 170494
rect 260186 163258 260422 163494
rect 260186 156258 260422 156494
rect 260186 149258 260422 149494
rect 260186 142258 260422 142494
rect 260186 135258 260422 135494
rect 260186 128258 260422 128494
rect 260186 121258 260422 121494
rect 260186 114258 260422 114494
rect 260186 107258 260422 107494
rect 260186 100258 260422 100494
rect 260186 93258 260422 93494
rect 260186 86258 260422 86494
rect 260186 79258 260422 79494
rect 260186 72258 260422 72494
rect 260186 65258 260422 65494
rect 260186 58258 260422 58494
rect 260186 51258 260422 51494
rect 260186 44258 260422 44494
rect 260186 37258 260422 37494
rect 260186 30258 260422 30494
rect 260186 23258 260422 23494
rect 260186 16258 260422 16494
rect 260186 9258 260422 9494
rect 260186 2258 260422 2494
rect 260186 -982 260422 -746
rect 260186 -1302 260422 -1066
rect 261918 705962 262154 706198
rect 261918 705642 262154 705878
rect 261918 696325 262154 696561
rect 261918 689325 262154 689561
rect 261918 682325 262154 682561
rect 261918 675325 262154 675561
rect 261918 668325 262154 668561
rect 261918 661325 262154 661561
rect 261918 654325 262154 654561
rect 261918 647325 262154 647561
rect 261918 640325 262154 640561
rect 261918 633325 262154 633561
rect 261918 626325 262154 626561
rect 261918 619325 262154 619561
rect 261918 612325 262154 612561
rect 261918 605325 262154 605561
rect 261918 598325 262154 598561
rect 261918 591325 262154 591561
rect 261918 584325 262154 584561
rect 261918 577325 262154 577561
rect 261918 570325 262154 570561
rect 261918 563325 262154 563561
rect 261918 556325 262154 556561
rect 261918 549325 262154 549561
rect 261918 542325 262154 542561
rect 261918 535325 262154 535561
rect 261918 528325 262154 528561
rect 261918 521325 262154 521561
rect 261918 514325 262154 514561
rect 261918 507325 262154 507561
rect 261918 500325 262154 500561
rect 261918 493325 262154 493561
rect 261918 486325 262154 486561
rect 261918 479325 262154 479561
rect 261918 472325 262154 472561
rect 261918 465325 262154 465561
rect 261918 458325 262154 458561
rect 261918 451325 262154 451561
rect 261918 444325 262154 444561
rect 261918 437325 262154 437561
rect 261918 430325 262154 430561
rect 261918 423325 262154 423561
rect 261918 416325 262154 416561
rect 261918 409325 262154 409561
rect 261918 402325 262154 402561
rect 261918 395325 262154 395561
rect 261918 388325 262154 388561
rect 261918 381325 262154 381561
rect 261918 374325 262154 374561
rect 261918 367325 262154 367561
rect 261918 360325 262154 360561
rect 261918 353325 262154 353561
rect 261918 346325 262154 346561
rect 261918 339325 262154 339561
rect 261918 332325 262154 332561
rect 261918 325325 262154 325561
rect 261918 318325 262154 318561
rect 261918 311325 262154 311561
rect 261918 304325 262154 304561
rect 261918 297325 262154 297561
rect 261918 290325 262154 290561
rect 261918 283325 262154 283561
rect 261918 276325 262154 276561
rect 261918 269325 262154 269561
rect 261918 262325 262154 262561
rect 261918 255325 262154 255561
rect 261918 248325 262154 248561
rect 261918 241325 262154 241561
rect 261918 234325 262154 234561
rect 261918 227325 262154 227561
rect 261918 220325 262154 220561
rect 261918 213325 262154 213561
rect 261918 206325 262154 206561
rect 261918 199325 262154 199561
rect 261918 192325 262154 192561
rect 261918 185325 262154 185561
rect 261918 178325 262154 178561
rect 261918 171325 262154 171561
rect 261918 164325 262154 164561
rect 261918 157325 262154 157561
rect 261918 150325 262154 150561
rect 261918 143325 262154 143561
rect 261918 136325 262154 136561
rect 261918 129325 262154 129561
rect 261918 122325 262154 122561
rect 261918 115325 262154 115561
rect 261918 108325 262154 108561
rect 261918 101325 262154 101561
rect 261918 94325 262154 94561
rect 261918 87325 262154 87561
rect 261918 80325 262154 80561
rect 261918 73325 262154 73561
rect 261918 66325 262154 66561
rect 261918 59325 262154 59561
rect 261918 52325 262154 52561
rect 261918 45325 262154 45561
rect 261918 38325 262154 38561
rect 261918 31325 262154 31561
rect 261918 24325 262154 24561
rect 261918 17325 262154 17561
rect 261918 10325 262154 10561
rect 261918 3325 262154 3561
rect 261918 -1942 262154 -1706
rect 261918 -2262 262154 -2026
rect 267186 705002 267422 705238
rect 267186 704682 267422 704918
rect 267186 695258 267422 695494
rect 267186 688258 267422 688494
rect 267186 681258 267422 681494
rect 267186 674258 267422 674494
rect 267186 667258 267422 667494
rect 267186 660258 267422 660494
rect 267186 653258 267422 653494
rect 267186 646258 267422 646494
rect 267186 639258 267422 639494
rect 267186 632258 267422 632494
rect 267186 625258 267422 625494
rect 267186 618258 267422 618494
rect 267186 611258 267422 611494
rect 267186 604258 267422 604494
rect 267186 597258 267422 597494
rect 267186 590258 267422 590494
rect 267186 583258 267422 583494
rect 267186 576258 267422 576494
rect 267186 569258 267422 569494
rect 267186 562258 267422 562494
rect 267186 555258 267422 555494
rect 267186 548258 267422 548494
rect 267186 541258 267422 541494
rect 267186 534258 267422 534494
rect 267186 527258 267422 527494
rect 267186 520258 267422 520494
rect 267186 513258 267422 513494
rect 267186 506258 267422 506494
rect 267186 499258 267422 499494
rect 267186 492258 267422 492494
rect 267186 485258 267422 485494
rect 267186 478258 267422 478494
rect 267186 471258 267422 471494
rect 267186 464258 267422 464494
rect 267186 457258 267422 457494
rect 267186 450258 267422 450494
rect 267186 443258 267422 443494
rect 267186 436258 267422 436494
rect 267186 429258 267422 429494
rect 267186 422258 267422 422494
rect 267186 415258 267422 415494
rect 267186 408258 267422 408494
rect 267186 401258 267422 401494
rect 267186 394258 267422 394494
rect 267186 387258 267422 387494
rect 267186 380258 267422 380494
rect 267186 373258 267422 373494
rect 267186 366258 267422 366494
rect 267186 359258 267422 359494
rect 267186 352258 267422 352494
rect 267186 345258 267422 345494
rect 267186 338258 267422 338494
rect 267186 331258 267422 331494
rect 267186 324258 267422 324494
rect 267186 317258 267422 317494
rect 267186 310258 267422 310494
rect 267186 303258 267422 303494
rect 267186 296258 267422 296494
rect 267186 289258 267422 289494
rect 267186 282258 267422 282494
rect 267186 275258 267422 275494
rect 267186 268258 267422 268494
rect 267186 261258 267422 261494
rect 267186 254258 267422 254494
rect 267186 247258 267422 247494
rect 267186 240258 267422 240494
rect 267186 233258 267422 233494
rect 267186 226258 267422 226494
rect 267186 219258 267422 219494
rect 267186 212258 267422 212494
rect 267186 205258 267422 205494
rect 267186 198258 267422 198494
rect 267186 191258 267422 191494
rect 267186 184258 267422 184494
rect 267186 177258 267422 177494
rect 267186 170258 267422 170494
rect 267186 163258 267422 163494
rect 267186 156258 267422 156494
rect 267186 149258 267422 149494
rect 267186 142258 267422 142494
rect 267186 135258 267422 135494
rect 267186 128258 267422 128494
rect 267186 121258 267422 121494
rect 267186 114258 267422 114494
rect 267186 107258 267422 107494
rect 267186 100258 267422 100494
rect 267186 93258 267422 93494
rect 267186 86258 267422 86494
rect 267186 79258 267422 79494
rect 267186 72258 267422 72494
rect 267186 65258 267422 65494
rect 267186 58258 267422 58494
rect 267186 51258 267422 51494
rect 267186 44258 267422 44494
rect 267186 37258 267422 37494
rect 267186 30258 267422 30494
rect 267186 23258 267422 23494
rect 267186 16258 267422 16494
rect 267186 9258 267422 9494
rect 267186 2258 267422 2494
rect 267186 -982 267422 -746
rect 267186 -1302 267422 -1066
rect 268918 705962 269154 706198
rect 268918 705642 269154 705878
rect 268918 696325 269154 696561
rect 268918 689325 269154 689561
rect 268918 682325 269154 682561
rect 268918 675325 269154 675561
rect 268918 668325 269154 668561
rect 268918 661325 269154 661561
rect 268918 654325 269154 654561
rect 268918 647325 269154 647561
rect 268918 640325 269154 640561
rect 268918 633325 269154 633561
rect 268918 626325 269154 626561
rect 268918 619325 269154 619561
rect 268918 612325 269154 612561
rect 268918 605325 269154 605561
rect 268918 598325 269154 598561
rect 268918 591325 269154 591561
rect 268918 584325 269154 584561
rect 268918 577325 269154 577561
rect 268918 570325 269154 570561
rect 268918 563325 269154 563561
rect 268918 556325 269154 556561
rect 268918 549325 269154 549561
rect 268918 542325 269154 542561
rect 268918 535325 269154 535561
rect 268918 528325 269154 528561
rect 268918 521325 269154 521561
rect 268918 514325 269154 514561
rect 268918 507325 269154 507561
rect 268918 500325 269154 500561
rect 268918 493325 269154 493561
rect 268918 486325 269154 486561
rect 268918 479325 269154 479561
rect 268918 472325 269154 472561
rect 268918 465325 269154 465561
rect 268918 458325 269154 458561
rect 268918 451325 269154 451561
rect 268918 444325 269154 444561
rect 268918 437325 269154 437561
rect 268918 430325 269154 430561
rect 268918 423325 269154 423561
rect 268918 416325 269154 416561
rect 268918 409325 269154 409561
rect 268918 402325 269154 402561
rect 268918 395325 269154 395561
rect 268918 388325 269154 388561
rect 268918 381325 269154 381561
rect 268918 374325 269154 374561
rect 268918 367325 269154 367561
rect 268918 360325 269154 360561
rect 268918 353325 269154 353561
rect 268918 346325 269154 346561
rect 268918 339325 269154 339561
rect 268918 332325 269154 332561
rect 268918 325325 269154 325561
rect 268918 318325 269154 318561
rect 268918 311325 269154 311561
rect 268918 304325 269154 304561
rect 268918 297325 269154 297561
rect 268918 290325 269154 290561
rect 268918 283325 269154 283561
rect 268918 276325 269154 276561
rect 268918 269325 269154 269561
rect 268918 262325 269154 262561
rect 268918 255325 269154 255561
rect 268918 248325 269154 248561
rect 268918 241325 269154 241561
rect 268918 234325 269154 234561
rect 268918 227325 269154 227561
rect 268918 220325 269154 220561
rect 268918 213325 269154 213561
rect 268918 206325 269154 206561
rect 268918 199325 269154 199561
rect 268918 192325 269154 192561
rect 268918 185325 269154 185561
rect 268918 178325 269154 178561
rect 268918 171325 269154 171561
rect 268918 164325 269154 164561
rect 268918 157325 269154 157561
rect 268918 150325 269154 150561
rect 268918 143325 269154 143561
rect 268918 136325 269154 136561
rect 268918 129325 269154 129561
rect 268918 122325 269154 122561
rect 268918 115325 269154 115561
rect 268918 108325 269154 108561
rect 268918 101325 269154 101561
rect 268918 94325 269154 94561
rect 268918 87325 269154 87561
rect 268918 80325 269154 80561
rect 268918 73325 269154 73561
rect 268918 66325 269154 66561
rect 268918 59325 269154 59561
rect 268918 52325 269154 52561
rect 268918 45325 269154 45561
rect 268918 38325 269154 38561
rect 268918 31325 269154 31561
rect 268918 24325 269154 24561
rect 268918 17325 269154 17561
rect 268918 10325 269154 10561
rect 268918 3325 269154 3561
rect 268918 -1942 269154 -1706
rect 268918 -2262 269154 -2026
rect 274186 705002 274422 705238
rect 274186 704682 274422 704918
rect 274186 695258 274422 695494
rect 274186 688258 274422 688494
rect 274186 681258 274422 681494
rect 274186 674258 274422 674494
rect 274186 667258 274422 667494
rect 274186 660258 274422 660494
rect 274186 653258 274422 653494
rect 274186 646258 274422 646494
rect 274186 639258 274422 639494
rect 274186 632258 274422 632494
rect 274186 625258 274422 625494
rect 274186 618258 274422 618494
rect 274186 611258 274422 611494
rect 274186 604258 274422 604494
rect 274186 597258 274422 597494
rect 274186 590258 274422 590494
rect 274186 583258 274422 583494
rect 274186 576258 274422 576494
rect 274186 569258 274422 569494
rect 274186 562258 274422 562494
rect 274186 555258 274422 555494
rect 274186 548258 274422 548494
rect 274186 541258 274422 541494
rect 274186 534258 274422 534494
rect 274186 527258 274422 527494
rect 274186 520258 274422 520494
rect 274186 513258 274422 513494
rect 274186 506258 274422 506494
rect 274186 499258 274422 499494
rect 274186 492258 274422 492494
rect 274186 485258 274422 485494
rect 274186 478258 274422 478494
rect 274186 471258 274422 471494
rect 274186 464258 274422 464494
rect 274186 457258 274422 457494
rect 274186 450258 274422 450494
rect 274186 443258 274422 443494
rect 274186 436258 274422 436494
rect 274186 429258 274422 429494
rect 274186 422258 274422 422494
rect 274186 415258 274422 415494
rect 274186 408258 274422 408494
rect 274186 401258 274422 401494
rect 274186 394258 274422 394494
rect 274186 387258 274422 387494
rect 274186 380258 274422 380494
rect 274186 373258 274422 373494
rect 274186 366258 274422 366494
rect 274186 359258 274422 359494
rect 274186 352258 274422 352494
rect 274186 345258 274422 345494
rect 274186 338258 274422 338494
rect 274186 331258 274422 331494
rect 274186 324258 274422 324494
rect 274186 317258 274422 317494
rect 274186 310258 274422 310494
rect 274186 303258 274422 303494
rect 274186 296258 274422 296494
rect 274186 289258 274422 289494
rect 274186 282258 274422 282494
rect 274186 275258 274422 275494
rect 274186 268258 274422 268494
rect 274186 261258 274422 261494
rect 274186 254258 274422 254494
rect 274186 247258 274422 247494
rect 274186 240258 274422 240494
rect 274186 233258 274422 233494
rect 274186 226258 274422 226494
rect 274186 219258 274422 219494
rect 274186 212258 274422 212494
rect 274186 205258 274422 205494
rect 274186 198258 274422 198494
rect 274186 191258 274422 191494
rect 274186 184258 274422 184494
rect 274186 177258 274422 177494
rect 274186 170258 274422 170494
rect 274186 163258 274422 163494
rect 274186 156258 274422 156494
rect 274186 149258 274422 149494
rect 274186 142258 274422 142494
rect 274186 135258 274422 135494
rect 274186 128258 274422 128494
rect 274186 121258 274422 121494
rect 274186 114258 274422 114494
rect 274186 107258 274422 107494
rect 274186 100258 274422 100494
rect 274186 93258 274422 93494
rect 274186 86258 274422 86494
rect 274186 79258 274422 79494
rect 274186 72258 274422 72494
rect 274186 65258 274422 65494
rect 274186 58258 274422 58494
rect 274186 51258 274422 51494
rect 274186 44258 274422 44494
rect 274186 37258 274422 37494
rect 274186 30258 274422 30494
rect 274186 23258 274422 23494
rect 274186 16258 274422 16494
rect 274186 9258 274422 9494
rect 274186 2258 274422 2494
rect 274186 -982 274422 -746
rect 274186 -1302 274422 -1066
rect 275918 705962 276154 706198
rect 275918 705642 276154 705878
rect 275918 696325 276154 696561
rect 275918 689325 276154 689561
rect 275918 682325 276154 682561
rect 275918 675325 276154 675561
rect 275918 668325 276154 668561
rect 275918 661325 276154 661561
rect 275918 654325 276154 654561
rect 275918 647325 276154 647561
rect 275918 640325 276154 640561
rect 275918 633325 276154 633561
rect 275918 626325 276154 626561
rect 275918 619325 276154 619561
rect 275918 612325 276154 612561
rect 275918 605325 276154 605561
rect 275918 598325 276154 598561
rect 275918 591325 276154 591561
rect 275918 584325 276154 584561
rect 275918 577325 276154 577561
rect 275918 570325 276154 570561
rect 275918 563325 276154 563561
rect 275918 556325 276154 556561
rect 275918 549325 276154 549561
rect 275918 542325 276154 542561
rect 275918 535325 276154 535561
rect 275918 528325 276154 528561
rect 275918 521325 276154 521561
rect 275918 514325 276154 514561
rect 275918 507325 276154 507561
rect 275918 500325 276154 500561
rect 275918 493325 276154 493561
rect 275918 486325 276154 486561
rect 275918 479325 276154 479561
rect 275918 472325 276154 472561
rect 275918 465325 276154 465561
rect 275918 458325 276154 458561
rect 275918 451325 276154 451561
rect 275918 444325 276154 444561
rect 275918 437325 276154 437561
rect 275918 430325 276154 430561
rect 275918 423325 276154 423561
rect 275918 416325 276154 416561
rect 275918 409325 276154 409561
rect 275918 402325 276154 402561
rect 275918 395325 276154 395561
rect 275918 388325 276154 388561
rect 275918 381325 276154 381561
rect 275918 374325 276154 374561
rect 275918 367325 276154 367561
rect 275918 360325 276154 360561
rect 275918 353325 276154 353561
rect 275918 346325 276154 346561
rect 275918 339325 276154 339561
rect 275918 332325 276154 332561
rect 275918 325325 276154 325561
rect 275918 318325 276154 318561
rect 275918 311325 276154 311561
rect 275918 304325 276154 304561
rect 275918 297325 276154 297561
rect 275918 290325 276154 290561
rect 275918 283325 276154 283561
rect 275918 276325 276154 276561
rect 275918 269325 276154 269561
rect 275918 262325 276154 262561
rect 275918 255325 276154 255561
rect 275918 248325 276154 248561
rect 275918 241325 276154 241561
rect 275918 234325 276154 234561
rect 275918 227325 276154 227561
rect 275918 220325 276154 220561
rect 275918 213325 276154 213561
rect 275918 206325 276154 206561
rect 275918 199325 276154 199561
rect 275918 192325 276154 192561
rect 275918 185325 276154 185561
rect 275918 178325 276154 178561
rect 275918 171325 276154 171561
rect 275918 164325 276154 164561
rect 275918 157325 276154 157561
rect 275918 150325 276154 150561
rect 275918 143325 276154 143561
rect 275918 136325 276154 136561
rect 275918 129325 276154 129561
rect 275918 122325 276154 122561
rect 275918 115325 276154 115561
rect 275918 108325 276154 108561
rect 275918 101325 276154 101561
rect 275918 94325 276154 94561
rect 275918 87325 276154 87561
rect 275918 80325 276154 80561
rect 275918 73325 276154 73561
rect 275918 66325 276154 66561
rect 275918 59325 276154 59561
rect 275918 52325 276154 52561
rect 275918 45325 276154 45561
rect 275918 38325 276154 38561
rect 275918 31325 276154 31561
rect 275918 24325 276154 24561
rect 275918 17325 276154 17561
rect 275918 10325 276154 10561
rect 275918 3325 276154 3561
rect 275918 -1942 276154 -1706
rect 275918 -2262 276154 -2026
rect 281186 705002 281422 705238
rect 281186 704682 281422 704918
rect 281186 695258 281422 695494
rect 281186 688258 281422 688494
rect 281186 681258 281422 681494
rect 281186 674258 281422 674494
rect 281186 667258 281422 667494
rect 281186 660258 281422 660494
rect 281186 653258 281422 653494
rect 281186 646258 281422 646494
rect 281186 639258 281422 639494
rect 281186 632258 281422 632494
rect 281186 625258 281422 625494
rect 281186 618258 281422 618494
rect 281186 611258 281422 611494
rect 281186 604258 281422 604494
rect 281186 597258 281422 597494
rect 281186 590258 281422 590494
rect 281186 583258 281422 583494
rect 281186 576258 281422 576494
rect 281186 569258 281422 569494
rect 281186 562258 281422 562494
rect 281186 555258 281422 555494
rect 281186 548258 281422 548494
rect 281186 541258 281422 541494
rect 281186 534258 281422 534494
rect 281186 527258 281422 527494
rect 281186 520258 281422 520494
rect 281186 513258 281422 513494
rect 281186 506258 281422 506494
rect 281186 499258 281422 499494
rect 281186 492258 281422 492494
rect 281186 485258 281422 485494
rect 281186 478258 281422 478494
rect 281186 471258 281422 471494
rect 281186 464258 281422 464494
rect 281186 457258 281422 457494
rect 281186 450258 281422 450494
rect 281186 443258 281422 443494
rect 281186 436258 281422 436494
rect 281186 429258 281422 429494
rect 281186 422258 281422 422494
rect 281186 415258 281422 415494
rect 281186 408258 281422 408494
rect 281186 401258 281422 401494
rect 281186 394258 281422 394494
rect 281186 387258 281422 387494
rect 281186 380258 281422 380494
rect 281186 373258 281422 373494
rect 281186 366258 281422 366494
rect 281186 359258 281422 359494
rect 281186 352258 281422 352494
rect 281186 345258 281422 345494
rect 281186 338258 281422 338494
rect 281186 331258 281422 331494
rect 281186 324258 281422 324494
rect 281186 317258 281422 317494
rect 281186 310258 281422 310494
rect 281186 303258 281422 303494
rect 281186 296258 281422 296494
rect 281186 289258 281422 289494
rect 281186 282258 281422 282494
rect 281186 275258 281422 275494
rect 281186 268258 281422 268494
rect 281186 261258 281422 261494
rect 281186 254258 281422 254494
rect 281186 247258 281422 247494
rect 281186 240258 281422 240494
rect 281186 233258 281422 233494
rect 281186 226258 281422 226494
rect 281186 219258 281422 219494
rect 281186 212258 281422 212494
rect 281186 205258 281422 205494
rect 281186 198258 281422 198494
rect 281186 191258 281422 191494
rect 281186 184258 281422 184494
rect 281186 177258 281422 177494
rect 281186 170258 281422 170494
rect 281186 163258 281422 163494
rect 281186 156258 281422 156494
rect 281186 149258 281422 149494
rect 281186 142258 281422 142494
rect 281186 135258 281422 135494
rect 281186 128258 281422 128494
rect 281186 121258 281422 121494
rect 281186 114258 281422 114494
rect 281186 107258 281422 107494
rect 281186 100258 281422 100494
rect 281186 93258 281422 93494
rect 281186 86258 281422 86494
rect 281186 79258 281422 79494
rect 281186 72258 281422 72494
rect 281186 65258 281422 65494
rect 281186 58258 281422 58494
rect 281186 51258 281422 51494
rect 281186 44258 281422 44494
rect 281186 37258 281422 37494
rect 281186 30258 281422 30494
rect 281186 23258 281422 23494
rect 281186 16258 281422 16494
rect 281186 9258 281422 9494
rect 281186 2258 281422 2494
rect 281186 -982 281422 -746
rect 281186 -1302 281422 -1066
rect 282918 705962 283154 706198
rect 282918 705642 283154 705878
rect 282918 696325 283154 696561
rect 282918 689325 283154 689561
rect 282918 682325 283154 682561
rect 282918 675325 283154 675561
rect 282918 668325 283154 668561
rect 282918 661325 283154 661561
rect 282918 654325 283154 654561
rect 282918 647325 283154 647561
rect 282918 640325 283154 640561
rect 282918 633325 283154 633561
rect 282918 626325 283154 626561
rect 282918 619325 283154 619561
rect 282918 612325 283154 612561
rect 282918 605325 283154 605561
rect 282918 598325 283154 598561
rect 282918 591325 283154 591561
rect 282918 584325 283154 584561
rect 282918 577325 283154 577561
rect 282918 570325 283154 570561
rect 282918 563325 283154 563561
rect 282918 556325 283154 556561
rect 282918 549325 283154 549561
rect 282918 542325 283154 542561
rect 282918 535325 283154 535561
rect 282918 528325 283154 528561
rect 282918 521325 283154 521561
rect 282918 514325 283154 514561
rect 282918 507325 283154 507561
rect 282918 500325 283154 500561
rect 282918 493325 283154 493561
rect 282918 486325 283154 486561
rect 282918 479325 283154 479561
rect 282918 472325 283154 472561
rect 282918 465325 283154 465561
rect 282918 458325 283154 458561
rect 282918 451325 283154 451561
rect 282918 444325 283154 444561
rect 282918 437325 283154 437561
rect 282918 430325 283154 430561
rect 282918 423325 283154 423561
rect 282918 416325 283154 416561
rect 282918 409325 283154 409561
rect 282918 402325 283154 402561
rect 282918 395325 283154 395561
rect 282918 388325 283154 388561
rect 282918 381325 283154 381561
rect 282918 374325 283154 374561
rect 282918 367325 283154 367561
rect 282918 360325 283154 360561
rect 282918 353325 283154 353561
rect 282918 346325 283154 346561
rect 282918 339325 283154 339561
rect 282918 332325 283154 332561
rect 282918 325325 283154 325561
rect 282918 318325 283154 318561
rect 282918 311325 283154 311561
rect 282918 304325 283154 304561
rect 282918 297325 283154 297561
rect 282918 290325 283154 290561
rect 282918 283325 283154 283561
rect 282918 276325 283154 276561
rect 282918 269325 283154 269561
rect 282918 262325 283154 262561
rect 282918 255325 283154 255561
rect 282918 248325 283154 248561
rect 282918 241325 283154 241561
rect 282918 234325 283154 234561
rect 282918 227325 283154 227561
rect 282918 220325 283154 220561
rect 282918 213325 283154 213561
rect 282918 206325 283154 206561
rect 282918 199325 283154 199561
rect 282918 192325 283154 192561
rect 282918 185325 283154 185561
rect 282918 178325 283154 178561
rect 282918 171325 283154 171561
rect 282918 164325 283154 164561
rect 282918 157325 283154 157561
rect 282918 150325 283154 150561
rect 282918 143325 283154 143561
rect 282918 136325 283154 136561
rect 282918 129325 283154 129561
rect 282918 122325 283154 122561
rect 282918 115325 283154 115561
rect 282918 108325 283154 108561
rect 282918 101325 283154 101561
rect 282918 94325 283154 94561
rect 282918 87325 283154 87561
rect 282918 80325 283154 80561
rect 282918 73325 283154 73561
rect 282918 66325 283154 66561
rect 282918 59325 283154 59561
rect 282918 52325 283154 52561
rect 282918 45325 283154 45561
rect 282918 38325 283154 38561
rect 282918 31325 283154 31561
rect 282918 24325 283154 24561
rect 282918 17325 283154 17561
rect 282918 10325 283154 10561
rect 282918 3325 283154 3561
rect 282918 -1942 283154 -1706
rect 282918 -2262 283154 -2026
rect 288186 705002 288422 705238
rect 288186 704682 288422 704918
rect 288186 695258 288422 695494
rect 288186 688258 288422 688494
rect 288186 681258 288422 681494
rect 288186 674258 288422 674494
rect 288186 667258 288422 667494
rect 288186 660258 288422 660494
rect 288186 653258 288422 653494
rect 288186 646258 288422 646494
rect 288186 639258 288422 639494
rect 288186 632258 288422 632494
rect 288186 625258 288422 625494
rect 288186 618258 288422 618494
rect 288186 611258 288422 611494
rect 288186 604258 288422 604494
rect 288186 597258 288422 597494
rect 288186 590258 288422 590494
rect 288186 583258 288422 583494
rect 288186 576258 288422 576494
rect 288186 569258 288422 569494
rect 288186 562258 288422 562494
rect 288186 555258 288422 555494
rect 288186 548258 288422 548494
rect 288186 541258 288422 541494
rect 288186 534258 288422 534494
rect 288186 527258 288422 527494
rect 288186 520258 288422 520494
rect 288186 513258 288422 513494
rect 288186 506258 288422 506494
rect 288186 499258 288422 499494
rect 288186 492258 288422 492494
rect 288186 485258 288422 485494
rect 288186 478258 288422 478494
rect 288186 471258 288422 471494
rect 288186 464258 288422 464494
rect 288186 457258 288422 457494
rect 288186 450258 288422 450494
rect 288186 443258 288422 443494
rect 288186 436258 288422 436494
rect 288186 429258 288422 429494
rect 288186 422258 288422 422494
rect 288186 415258 288422 415494
rect 288186 408258 288422 408494
rect 288186 401258 288422 401494
rect 288186 394258 288422 394494
rect 288186 387258 288422 387494
rect 288186 380258 288422 380494
rect 288186 373258 288422 373494
rect 288186 366258 288422 366494
rect 288186 359258 288422 359494
rect 288186 352258 288422 352494
rect 288186 345258 288422 345494
rect 288186 338258 288422 338494
rect 288186 331258 288422 331494
rect 288186 324258 288422 324494
rect 288186 317258 288422 317494
rect 288186 310258 288422 310494
rect 288186 303258 288422 303494
rect 288186 296258 288422 296494
rect 288186 289258 288422 289494
rect 288186 282258 288422 282494
rect 288186 275258 288422 275494
rect 288186 268258 288422 268494
rect 288186 261258 288422 261494
rect 288186 254258 288422 254494
rect 288186 247258 288422 247494
rect 288186 240258 288422 240494
rect 288186 233258 288422 233494
rect 288186 226258 288422 226494
rect 288186 219258 288422 219494
rect 288186 212258 288422 212494
rect 288186 205258 288422 205494
rect 288186 198258 288422 198494
rect 288186 191258 288422 191494
rect 288186 184258 288422 184494
rect 288186 177258 288422 177494
rect 288186 170258 288422 170494
rect 288186 163258 288422 163494
rect 288186 156258 288422 156494
rect 288186 149258 288422 149494
rect 288186 142258 288422 142494
rect 288186 135258 288422 135494
rect 288186 128258 288422 128494
rect 288186 121258 288422 121494
rect 288186 114258 288422 114494
rect 288186 107258 288422 107494
rect 288186 100258 288422 100494
rect 288186 93258 288422 93494
rect 288186 86258 288422 86494
rect 288186 79258 288422 79494
rect 288186 72258 288422 72494
rect 288186 65258 288422 65494
rect 288186 58258 288422 58494
rect 288186 51258 288422 51494
rect 288186 44258 288422 44494
rect 288186 37258 288422 37494
rect 288186 30258 288422 30494
rect 288186 23258 288422 23494
rect 288186 16258 288422 16494
rect 288186 9258 288422 9494
rect 288186 2258 288422 2494
rect 288186 -982 288422 -746
rect 288186 -1302 288422 -1066
rect 289918 705962 290154 706198
rect 289918 705642 290154 705878
rect 289918 696325 290154 696561
rect 289918 689325 290154 689561
rect 289918 682325 290154 682561
rect 289918 675325 290154 675561
rect 289918 668325 290154 668561
rect 289918 661325 290154 661561
rect 289918 654325 290154 654561
rect 289918 647325 290154 647561
rect 289918 640325 290154 640561
rect 289918 633325 290154 633561
rect 289918 626325 290154 626561
rect 289918 619325 290154 619561
rect 289918 612325 290154 612561
rect 289918 605325 290154 605561
rect 289918 598325 290154 598561
rect 289918 591325 290154 591561
rect 289918 584325 290154 584561
rect 289918 577325 290154 577561
rect 289918 570325 290154 570561
rect 289918 563325 290154 563561
rect 289918 556325 290154 556561
rect 289918 549325 290154 549561
rect 289918 542325 290154 542561
rect 289918 535325 290154 535561
rect 289918 528325 290154 528561
rect 289918 521325 290154 521561
rect 289918 514325 290154 514561
rect 289918 507325 290154 507561
rect 289918 500325 290154 500561
rect 289918 493325 290154 493561
rect 289918 486325 290154 486561
rect 289918 479325 290154 479561
rect 289918 472325 290154 472561
rect 289918 465325 290154 465561
rect 289918 458325 290154 458561
rect 289918 451325 290154 451561
rect 289918 444325 290154 444561
rect 289918 437325 290154 437561
rect 289918 430325 290154 430561
rect 289918 423325 290154 423561
rect 289918 416325 290154 416561
rect 289918 409325 290154 409561
rect 289918 402325 290154 402561
rect 289918 395325 290154 395561
rect 289918 388325 290154 388561
rect 289918 381325 290154 381561
rect 289918 374325 290154 374561
rect 295186 705002 295422 705238
rect 295186 704682 295422 704918
rect 295186 695258 295422 695494
rect 295186 688258 295422 688494
rect 295186 681258 295422 681494
rect 295186 674258 295422 674494
rect 295186 667258 295422 667494
rect 295186 660258 295422 660494
rect 295186 653258 295422 653494
rect 295186 646258 295422 646494
rect 295186 639258 295422 639494
rect 295186 632258 295422 632494
rect 295186 625258 295422 625494
rect 295186 618258 295422 618494
rect 295186 611258 295422 611494
rect 295186 604258 295422 604494
rect 295186 597258 295422 597494
rect 295186 590258 295422 590494
rect 295186 583258 295422 583494
rect 295186 576258 295422 576494
rect 295186 569258 295422 569494
rect 295186 562258 295422 562494
rect 295186 555258 295422 555494
rect 295186 548258 295422 548494
rect 295186 541258 295422 541494
rect 295186 534258 295422 534494
rect 295186 527258 295422 527494
rect 295186 520258 295422 520494
rect 295186 513258 295422 513494
rect 295186 506258 295422 506494
rect 295186 499258 295422 499494
rect 295186 492258 295422 492494
rect 295186 485258 295422 485494
rect 295186 478258 295422 478494
rect 295186 471258 295422 471494
rect 295186 464258 295422 464494
rect 295186 457258 295422 457494
rect 295186 450258 295422 450494
rect 295186 443258 295422 443494
rect 295186 436258 295422 436494
rect 295186 429258 295422 429494
rect 295186 422258 295422 422494
rect 295186 415258 295422 415494
rect 295186 408258 295422 408494
rect 295186 401258 295422 401494
rect 295186 394258 295422 394494
rect 295186 387258 295422 387494
rect 295186 380258 295422 380494
rect 295186 373258 295422 373494
rect 296918 705962 297154 706198
rect 296918 705642 297154 705878
rect 296918 696325 297154 696561
rect 296918 689325 297154 689561
rect 296918 682325 297154 682561
rect 296918 675325 297154 675561
rect 296918 668325 297154 668561
rect 296918 661325 297154 661561
rect 296918 654325 297154 654561
rect 296918 647325 297154 647561
rect 296918 640325 297154 640561
rect 296918 633325 297154 633561
rect 296918 626325 297154 626561
rect 296918 619325 297154 619561
rect 296918 612325 297154 612561
rect 296918 605325 297154 605561
rect 296918 598325 297154 598561
rect 296918 591325 297154 591561
rect 296918 584325 297154 584561
rect 296918 577325 297154 577561
rect 296918 570325 297154 570561
rect 296918 563325 297154 563561
rect 296918 556325 297154 556561
rect 296918 549325 297154 549561
rect 296918 542325 297154 542561
rect 296918 535325 297154 535561
rect 296918 528325 297154 528561
rect 296918 521325 297154 521561
rect 296918 514325 297154 514561
rect 296918 507325 297154 507561
rect 296918 500325 297154 500561
rect 296918 493325 297154 493561
rect 296918 486325 297154 486561
rect 296918 479325 297154 479561
rect 296918 472325 297154 472561
rect 296918 465325 297154 465561
rect 296918 458325 297154 458561
rect 296918 451514 296948 451561
rect 296948 451514 296964 451561
rect 296964 451514 297028 451561
rect 297028 451514 297044 451561
rect 297044 451514 297108 451561
rect 297108 451514 297124 451561
rect 297124 451514 297154 451561
rect 296918 451498 297154 451514
rect 296918 451434 296948 451498
rect 296948 451434 296964 451498
rect 296964 451434 297028 451498
rect 297028 451434 297044 451498
rect 297044 451434 297108 451498
rect 297108 451434 297124 451498
rect 297124 451434 297154 451498
rect 296918 451418 297154 451434
rect 296918 451354 296948 451418
rect 296948 451354 296964 451418
rect 296964 451354 297028 451418
rect 297028 451354 297044 451418
rect 297044 451354 297108 451418
rect 297108 451354 297124 451418
rect 297124 451354 297154 451418
rect 296918 451338 297154 451354
rect 296918 451325 296948 451338
rect 296948 451325 296964 451338
rect 296964 451325 297028 451338
rect 297028 451325 297044 451338
rect 297044 451325 297108 451338
rect 297108 451325 297124 451338
rect 297124 451325 297154 451338
rect 296918 444325 297154 444561
rect 296918 437325 297154 437561
rect 296918 430325 297154 430561
rect 296918 423325 297154 423561
rect 296918 416325 297154 416561
rect 296918 409325 297154 409561
rect 296918 402325 297154 402561
rect 296918 395325 297154 395561
rect 296918 388325 297154 388561
rect 296918 381325 297154 381561
rect 296918 374325 297154 374561
rect 302186 705002 302422 705238
rect 302186 704682 302422 704918
rect 302186 695258 302422 695494
rect 302186 688258 302422 688494
rect 302186 681258 302422 681494
rect 302186 674258 302422 674494
rect 302186 667258 302422 667494
rect 302186 660258 302422 660494
rect 302186 653258 302422 653494
rect 302186 646258 302422 646494
rect 302186 639258 302422 639494
rect 302186 632258 302422 632494
rect 302186 625258 302422 625494
rect 302186 618258 302422 618494
rect 302186 611258 302422 611494
rect 302186 604258 302422 604494
rect 302186 597258 302422 597494
rect 302186 590258 302422 590494
rect 302186 583258 302422 583494
rect 302186 576258 302422 576494
rect 302186 569258 302422 569494
rect 302186 562258 302422 562494
rect 302186 555258 302422 555494
rect 302186 548258 302422 548494
rect 302186 541258 302422 541494
rect 302186 534258 302422 534494
rect 302186 527258 302422 527494
rect 302186 520258 302422 520494
rect 302186 513258 302422 513494
rect 302186 506258 302422 506494
rect 302186 499258 302422 499494
rect 302186 492258 302422 492494
rect 302186 485258 302422 485494
rect 302186 478258 302422 478494
rect 302186 471258 302422 471494
rect 302186 464258 302422 464494
rect 302186 457258 302422 457494
rect 302186 450258 302422 450494
rect 302186 443258 302422 443494
rect 302186 436258 302422 436494
rect 302186 429258 302422 429494
rect 302186 422258 302422 422494
rect 302186 415258 302422 415494
rect 302186 408258 302422 408494
rect 302186 401258 302422 401494
rect 302186 394258 302422 394494
rect 302186 387258 302422 387494
rect 302186 380258 302422 380494
rect 302186 373258 302422 373494
rect 303918 705962 304154 706198
rect 303918 705642 304154 705878
rect 303918 696325 304154 696561
rect 303918 689325 304154 689561
rect 303918 682325 304154 682561
rect 303918 675325 304154 675561
rect 303918 668325 304154 668561
rect 303918 661325 304154 661561
rect 303918 654325 304154 654561
rect 303918 647325 304154 647561
rect 303918 640325 304154 640561
rect 303918 633325 304154 633561
rect 303918 626325 304154 626561
rect 303918 619325 304154 619561
rect 303918 612325 304154 612561
rect 303918 605325 304154 605561
rect 303918 598325 304154 598561
rect 303918 591325 304154 591561
rect 303918 584325 304154 584561
rect 303918 577325 304154 577561
rect 303918 570325 304154 570561
rect 303918 563325 304154 563561
rect 303918 556325 304154 556561
rect 303918 549325 304154 549561
rect 303918 542325 304154 542561
rect 303918 535325 304154 535561
rect 303918 528325 304154 528561
rect 303918 521325 304154 521561
rect 303918 514325 304154 514561
rect 303918 507325 304154 507561
rect 303918 500325 304154 500561
rect 303918 493325 304154 493561
rect 303918 486325 304154 486561
rect 303918 479325 304154 479561
rect 303918 472325 304154 472561
rect 303918 465325 304154 465561
rect 303918 458325 304154 458561
rect 303918 451514 303948 451561
rect 303948 451514 303964 451561
rect 303964 451514 304028 451561
rect 304028 451514 304044 451561
rect 304044 451514 304108 451561
rect 304108 451514 304124 451561
rect 304124 451514 304154 451561
rect 303918 451498 304154 451514
rect 303918 451434 303948 451498
rect 303948 451434 303964 451498
rect 303964 451434 304028 451498
rect 304028 451434 304044 451498
rect 304044 451434 304108 451498
rect 304108 451434 304124 451498
rect 304124 451434 304154 451498
rect 303918 451418 304154 451434
rect 303918 451354 303948 451418
rect 303948 451354 303964 451418
rect 303964 451354 304028 451418
rect 304028 451354 304044 451418
rect 304044 451354 304108 451418
rect 304108 451354 304124 451418
rect 304124 451354 304154 451418
rect 303918 451338 304154 451354
rect 303918 451325 303948 451338
rect 303948 451325 303964 451338
rect 303964 451325 304028 451338
rect 304028 451325 304044 451338
rect 304044 451325 304108 451338
rect 304108 451325 304124 451338
rect 304124 451325 304154 451338
rect 303918 444325 304154 444561
rect 303918 437325 304154 437561
rect 303918 430325 304154 430561
rect 303918 423325 304154 423561
rect 303918 416325 304154 416561
rect 303918 409325 304154 409561
rect 303918 402325 304154 402561
rect 303918 395325 304154 395561
rect 303918 388325 304154 388561
rect 303918 381325 304154 381561
rect 303918 374325 304154 374561
rect 309186 705002 309422 705238
rect 309186 704682 309422 704918
rect 309186 695258 309422 695494
rect 309186 688258 309422 688494
rect 309186 681258 309422 681494
rect 309186 674258 309422 674494
rect 309186 667258 309422 667494
rect 309186 660258 309422 660494
rect 309186 653258 309422 653494
rect 309186 646258 309422 646494
rect 309186 639258 309422 639494
rect 309186 632258 309422 632494
rect 309186 625258 309422 625494
rect 309186 618258 309422 618494
rect 309186 611258 309422 611494
rect 309186 604258 309422 604494
rect 309186 597258 309422 597494
rect 309186 590258 309422 590494
rect 309186 583258 309422 583494
rect 309186 576258 309422 576494
rect 309186 569258 309422 569494
rect 309186 562258 309422 562494
rect 309186 555258 309422 555494
rect 309186 548258 309422 548494
rect 309186 541258 309422 541494
rect 309186 534258 309422 534494
rect 309186 527258 309422 527494
rect 309186 520258 309422 520494
rect 309186 513258 309422 513494
rect 309186 506258 309422 506494
rect 309186 499258 309422 499494
rect 309186 492258 309422 492494
rect 309186 485258 309422 485494
rect 309186 478258 309422 478494
rect 309186 471258 309422 471494
rect 309186 464258 309422 464494
rect 309186 457258 309422 457494
rect 309186 450258 309422 450494
rect 309186 443258 309422 443494
rect 309186 436258 309422 436494
rect 309186 429258 309422 429494
rect 309186 422258 309422 422494
rect 309186 415258 309422 415494
rect 309186 408258 309422 408494
rect 309186 401258 309422 401494
rect 309186 394258 309422 394494
rect 309186 387258 309422 387494
rect 309186 380258 309422 380494
rect 309186 373258 309422 373494
rect 310918 705962 311154 706198
rect 310918 705642 311154 705878
rect 310918 696325 311154 696561
rect 310918 689325 311154 689561
rect 310918 682325 311154 682561
rect 310918 675325 311154 675561
rect 310918 668325 311154 668561
rect 310918 661325 311154 661561
rect 310918 654325 311154 654561
rect 310918 647325 311154 647561
rect 310918 640325 311154 640561
rect 310918 633325 311154 633561
rect 310918 626325 311154 626561
rect 310918 619325 311154 619561
rect 310918 612325 311154 612561
rect 310918 605325 311154 605561
rect 310918 598325 311154 598561
rect 310918 591325 311154 591561
rect 310918 584325 311154 584561
rect 310918 577325 311154 577561
rect 310918 570325 311154 570561
rect 310918 563325 311154 563561
rect 310918 556325 311154 556561
rect 310918 549325 311154 549561
rect 310918 542325 311154 542561
rect 310918 535325 311154 535561
rect 310918 528325 311154 528561
rect 310918 521325 311154 521561
rect 310918 514325 311154 514561
rect 310918 507325 311154 507561
rect 310918 500325 311154 500561
rect 310918 493325 311154 493561
rect 310918 486325 311154 486561
rect 310918 479325 311154 479561
rect 310918 472325 311154 472561
rect 310918 465325 311154 465561
rect 310918 458325 311154 458561
rect 310918 451514 310979 451561
rect 310979 451514 310995 451561
rect 310995 451514 311059 451561
rect 311059 451514 311154 451561
rect 310918 451498 311154 451514
rect 310918 451434 310979 451498
rect 310979 451434 310995 451498
rect 310995 451434 311059 451498
rect 311059 451434 311154 451498
rect 310918 451418 311154 451434
rect 310918 451354 310979 451418
rect 310979 451354 310995 451418
rect 310995 451354 311059 451418
rect 311059 451354 311154 451418
rect 310918 451338 311154 451354
rect 310918 451325 310979 451338
rect 310979 451325 310995 451338
rect 310995 451325 311059 451338
rect 311059 451325 311154 451338
rect 310918 444325 311154 444561
rect 310918 437325 311154 437561
rect 310918 430325 311154 430561
rect 310918 423325 311154 423561
rect 310918 416325 311154 416561
rect 310918 409325 311154 409561
rect 310918 402325 311154 402561
rect 310918 395325 311154 395561
rect 310918 388325 311154 388561
rect 310918 381325 311154 381561
rect 310918 374325 311154 374561
rect 316186 705002 316422 705238
rect 316186 704682 316422 704918
rect 316186 695258 316422 695494
rect 316186 688258 316422 688494
rect 316186 681258 316422 681494
rect 316186 674258 316422 674494
rect 316186 667258 316422 667494
rect 316186 660258 316422 660494
rect 316186 653258 316422 653494
rect 316186 646258 316422 646494
rect 316186 639258 316422 639494
rect 316186 632258 316422 632494
rect 316186 625258 316422 625494
rect 316186 618258 316422 618494
rect 316186 611258 316422 611494
rect 316186 604258 316422 604494
rect 316186 597258 316422 597494
rect 316186 590258 316422 590494
rect 316186 583258 316422 583494
rect 316186 576258 316422 576494
rect 316186 569258 316422 569494
rect 316186 562258 316422 562494
rect 316186 555258 316422 555494
rect 316186 548258 316422 548494
rect 316186 541258 316422 541494
rect 316186 534258 316422 534494
rect 316186 527258 316422 527494
rect 316186 520258 316422 520494
rect 316186 513258 316422 513494
rect 316186 506258 316422 506494
rect 316186 499258 316422 499494
rect 316186 492258 316422 492494
rect 316186 485258 316422 485494
rect 316186 478258 316422 478494
rect 316186 471258 316422 471494
rect 316186 464258 316422 464494
rect 316186 457258 316422 457494
rect 316186 450258 316422 450494
rect 316186 443258 316422 443494
rect 316186 436258 316422 436494
rect 316186 429258 316422 429494
rect 316186 422258 316422 422494
rect 316186 415258 316422 415494
rect 316186 408258 316422 408494
rect 316186 401258 316422 401494
rect 316186 394258 316422 394494
rect 316186 387258 316422 387494
rect 316186 380258 316422 380494
rect 316186 373258 316422 373494
rect 289918 367325 290154 367561
rect 316186 366258 316422 366494
rect 289918 360325 290154 360561
rect 289918 353325 290154 353561
rect 289918 346325 290154 346561
rect 289918 339325 290154 339561
rect 289918 332325 290154 332561
rect 289918 325325 290154 325561
rect 289918 318325 290154 318561
rect 289918 311325 290154 311561
rect 289918 304325 290154 304561
rect 289918 297325 290154 297561
rect 289918 290325 290154 290561
rect 289918 283325 290154 283561
rect 289918 276325 290154 276561
rect 289918 269325 290154 269561
rect 289918 262325 290154 262561
rect 289918 255325 290154 255561
rect 289918 248325 290154 248561
rect 289918 241325 290154 241561
rect 289918 234325 290154 234561
rect 289918 227325 290154 227561
rect 289918 220325 290154 220561
rect 289918 213325 290154 213561
rect 289918 206325 290154 206561
rect 295186 359258 295422 359494
rect 295186 352258 295422 352494
rect 295186 345258 295422 345494
rect 295186 338258 295422 338494
rect 295186 331258 295422 331494
rect 295186 324258 295422 324494
rect 295186 317258 295422 317494
rect 295186 310258 295422 310494
rect 295186 303258 295422 303494
rect 295186 296258 295422 296494
rect 295186 289258 295422 289494
rect 295186 282258 295422 282494
rect 295186 275258 295422 275494
rect 295186 268258 295422 268494
rect 295186 261258 295422 261494
rect 295186 254258 295422 254494
rect 295186 247258 295422 247494
rect 295186 240258 295422 240494
rect 295186 233258 295422 233494
rect 295186 226258 295422 226494
rect 295186 219258 295422 219494
rect 295186 212258 295422 212494
rect 295186 205258 295422 205494
rect 296918 360325 297154 360561
rect 296918 353325 297154 353561
rect 296918 346325 297154 346561
rect 296918 339325 297154 339561
rect 296918 332325 297154 332561
rect 296918 325325 297154 325561
rect 296918 318325 297154 318561
rect 296918 311325 297154 311561
rect 296918 304325 297154 304561
rect 296918 297325 297154 297561
rect 296918 290325 297154 290561
rect 296918 283325 297154 283561
rect 296918 276325 297154 276561
rect 296918 269325 297154 269561
rect 296918 262325 297154 262561
rect 296918 255325 297154 255561
rect 296918 248325 297154 248561
rect 296918 241325 297154 241561
rect 296918 234325 297154 234561
rect 296918 227325 297154 227561
rect 296918 220325 297154 220561
rect 296918 213325 297154 213561
rect 296918 206325 297154 206561
rect 302186 359258 302422 359494
rect 302186 352258 302422 352494
rect 302186 345258 302422 345494
rect 302186 338258 302422 338494
rect 302186 331258 302422 331494
rect 302186 324258 302422 324494
rect 302186 317258 302422 317494
rect 302186 310258 302422 310494
rect 302186 303258 302422 303494
rect 302186 296258 302422 296494
rect 302186 289258 302422 289494
rect 302186 282258 302422 282494
rect 302186 275258 302422 275494
rect 302186 268258 302422 268494
rect 302186 261258 302422 261494
rect 302186 254258 302422 254494
rect 302186 247258 302422 247494
rect 302186 240258 302422 240494
rect 302186 233258 302422 233494
rect 302186 226258 302422 226494
rect 302186 219258 302422 219494
rect 302186 212258 302422 212494
rect 302186 205258 302422 205494
rect 303918 360325 304154 360561
rect 303918 353325 304154 353561
rect 303918 346325 304154 346561
rect 303918 339325 304154 339561
rect 303918 332325 304154 332561
rect 303918 325325 304154 325561
rect 303918 318325 304154 318561
rect 303918 311325 304154 311561
rect 303918 304325 304154 304561
rect 303918 297325 304154 297561
rect 303918 290325 304154 290561
rect 303918 283325 304154 283561
rect 303918 276325 304154 276561
rect 303918 269325 304154 269561
rect 303918 262325 304154 262561
rect 303918 255325 304154 255561
rect 303918 248325 304154 248561
rect 303918 241325 304154 241561
rect 303918 234325 304154 234561
rect 303918 227325 304154 227561
rect 303918 220325 304154 220561
rect 303918 213325 304154 213561
rect 303918 206325 304154 206561
rect 309186 359258 309422 359494
rect 309186 352258 309422 352494
rect 309186 345258 309422 345494
rect 309186 338258 309422 338494
rect 309186 331258 309422 331494
rect 309186 324258 309422 324494
rect 309186 317258 309422 317494
rect 309186 310258 309422 310494
rect 309186 303258 309422 303494
rect 309186 296258 309422 296494
rect 309186 289258 309422 289494
rect 309186 282258 309422 282494
rect 309186 275258 309422 275494
rect 309186 268258 309422 268494
rect 309186 261258 309422 261494
rect 309186 254258 309422 254494
rect 309186 247258 309422 247494
rect 309186 240258 309422 240494
rect 309186 233258 309422 233494
rect 309186 226258 309422 226494
rect 309186 219258 309422 219494
rect 309186 212258 309422 212494
rect 309186 205258 309422 205494
rect 310918 360325 311154 360561
rect 310918 353325 311154 353561
rect 310918 346325 311154 346561
rect 310918 339325 311154 339561
rect 310918 332325 311154 332561
rect 310918 325325 311154 325561
rect 310918 318325 311154 318561
rect 310918 311325 311154 311561
rect 310918 304325 311154 304561
rect 310918 297325 311154 297561
rect 310918 290325 311154 290561
rect 310918 283325 311154 283561
rect 310918 276325 311154 276561
rect 310918 269325 311154 269561
rect 310918 262325 311154 262561
rect 310918 255325 311154 255561
rect 310918 248325 311154 248561
rect 310918 241325 311154 241561
rect 310918 234325 311154 234561
rect 310918 227325 311154 227561
rect 310918 220325 311154 220561
rect 310918 213325 311154 213561
rect 310918 206325 311154 206561
rect 316186 359258 316422 359494
rect 316186 352258 316422 352494
rect 316186 345258 316422 345494
rect 316186 338258 316422 338494
rect 316186 331258 316422 331494
rect 316186 324258 316422 324494
rect 316186 317258 316422 317494
rect 316186 310258 316422 310494
rect 316186 303258 316422 303494
rect 316186 296258 316422 296494
rect 316186 289258 316422 289494
rect 316186 282258 316422 282494
rect 316186 275258 316422 275494
rect 316186 268258 316422 268494
rect 316186 261258 316422 261494
rect 316186 254258 316422 254494
rect 316186 247258 316422 247494
rect 316186 240258 316422 240494
rect 316186 233258 316422 233494
rect 316186 226258 316422 226494
rect 316186 219258 316422 219494
rect 316186 212258 316422 212494
rect 316186 205258 316422 205494
rect 289918 199325 290154 199561
rect 316186 198258 316422 198494
rect 289918 192325 290154 192561
rect 289918 185325 290154 185561
rect 289918 178325 290154 178561
rect 289918 171325 290154 171561
rect 289918 164325 290154 164561
rect 289918 157325 290154 157561
rect 289918 150325 290154 150561
rect 289918 143325 290154 143561
rect 289918 136325 290154 136561
rect 289918 129325 290154 129561
rect 289918 122325 290154 122561
rect 289918 115325 290154 115561
rect 289918 108325 290154 108561
rect 289918 101325 290154 101561
rect 289918 94325 290154 94561
rect 289918 87325 290154 87561
rect 289918 80325 290154 80561
rect 289918 73325 290154 73561
rect 289918 66325 290154 66561
rect 289918 59325 290154 59561
rect 289918 52325 290154 52561
rect 289918 45325 290154 45561
rect 289918 38325 290154 38561
rect 289918 31325 290154 31561
rect 289918 24325 290154 24561
rect 289918 17325 290154 17561
rect 289918 10325 290154 10561
rect 289918 3325 290154 3561
rect 289918 -1942 290154 -1706
rect 289918 -2262 290154 -2026
rect 295186 191258 295422 191494
rect 295186 184258 295422 184494
rect 295186 177258 295422 177494
rect 295186 170258 295422 170494
rect 295186 163258 295422 163494
rect 295186 156258 295422 156494
rect 295186 149258 295422 149494
rect 295186 142258 295422 142494
rect 295186 135258 295422 135494
rect 295186 128258 295422 128494
rect 295186 121258 295422 121494
rect 295186 114258 295422 114494
rect 295186 107258 295422 107494
rect 295186 100258 295422 100494
rect 295186 93258 295422 93494
rect 295186 86258 295422 86494
rect 295186 79258 295422 79494
rect 295186 72258 295422 72494
rect 295186 65258 295422 65494
rect 295186 58258 295422 58494
rect 295186 51258 295422 51494
rect 295186 44258 295422 44494
rect 295186 37258 295422 37494
rect 295186 30258 295422 30494
rect 295186 23258 295422 23494
rect 295186 16258 295422 16494
rect 295186 9258 295422 9494
rect 295186 2258 295422 2494
rect 295186 -982 295422 -746
rect 295186 -1302 295422 -1066
rect 296918 192325 297154 192561
rect 296918 185325 297154 185561
rect 296918 178325 297154 178561
rect 296918 171325 297154 171561
rect 296918 164325 297154 164561
rect 296918 157325 297154 157561
rect 296918 150325 297154 150561
rect 296918 143325 297154 143561
rect 296918 136325 297154 136561
rect 296918 129325 297154 129561
rect 296918 122325 297154 122561
rect 296918 115325 297154 115561
rect 296918 108325 297154 108561
rect 296918 101325 297154 101561
rect 296918 94325 297154 94561
rect 296918 87325 297154 87561
rect 296918 80325 297154 80561
rect 296918 73325 297154 73561
rect 296918 66325 297154 66561
rect 296918 59325 297154 59561
rect 296918 52325 297154 52561
rect 296918 45325 297154 45561
rect 296918 38325 297154 38561
rect 296918 31325 297154 31561
rect 296918 24325 297154 24561
rect 296918 17325 297154 17561
rect 296918 10325 297154 10561
rect 296918 3325 297154 3561
rect 296918 -1942 297154 -1706
rect 296918 -2262 297154 -2026
rect 302186 191258 302422 191494
rect 302186 184258 302422 184494
rect 302186 177258 302422 177494
rect 302186 170258 302422 170494
rect 302186 163258 302422 163494
rect 302186 156258 302422 156494
rect 302186 149258 302422 149494
rect 302186 142258 302422 142494
rect 302186 135258 302422 135494
rect 302186 128258 302422 128494
rect 302186 121258 302422 121494
rect 302186 114258 302422 114494
rect 302186 107258 302422 107494
rect 302186 100258 302422 100494
rect 302186 93258 302422 93494
rect 302186 86258 302422 86494
rect 302186 79258 302422 79494
rect 302186 72258 302422 72494
rect 302186 65258 302422 65494
rect 302186 58258 302422 58494
rect 302186 51258 302422 51494
rect 302186 44258 302422 44494
rect 302186 37258 302422 37494
rect 302186 30258 302422 30494
rect 302186 23258 302422 23494
rect 302186 16258 302422 16494
rect 302186 9258 302422 9494
rect 302186 2258 302422 2494
rect 302186 -982 302422 -746
rect 302186 -1302 302422 -1066
rect 303918 192325 304154 192561
rect 303918 185325 304154 185561
rect 303918 178325 304154 178561
rect 303918 171325 304154 171561
rect 303918 164325 304154 164561
rect 303918 157325 304154 157561
rect 303918 150325 304154 150561
rect 303918 143325 304154 143561
rect 303918 136325 304154 136561
rect 303918 129325 304154 129561
rect 303918 122325 304154 122561
rect 303918 115325 304154 115561
rect 303918 108325 304154 108561
rect 303918 101325 304154 101561
rect 303918 94325 304154 94561
rect 303918 87325 304154 87561
rect 303918 80325 304154 80561
rect 303918 73325 304154 73561
rect 303918 66325 304154 66561
rect 303918 59325 304154 59561
rect 303918 52325 304154 52561
rect 303918 45325 304154 45561
rect 303918 38325 304154 38561
rect 303918 31325 304154 31561
rect 303918 24325 304154 24561
rect 303918 17325 304154 17561
rect 303918 10325 304154 10561
rect 303918 3325 304154 3561
rect 303918 -1942 304154 -1706
rect 303918 -2262 304154 -2026
rect 309186 191258 309422 191494
rect 309186 184258 309422 184494
rect 309186 177258 309422 177494
rect 309186 170258 309422 170494
rect 309186 163258 309422 163494
rect 309186 156258 309422 156494
rect 309186 149258 309422 149494
rect 309186 142258 309422 142494
rect 309186 135258 309422 135494
rect 309186 128258 309422 128494
rect 309186 121258 309422 121494
rect 309186 114258 309422 114494
rect 309186 107258 309422 107494
rect 309186 100258 309422 100494
rect 309186 93258 309422 93494
rect 309186 86258 309422 86494
rect 309186 79258 309422 79494
rect 309186 72258 309422 72494
rect 309186 65258 309422 65494
rect 309186 58258 309422 58494
rect 309186 51258 309422 51494
rect 309186 44258 309422 44494
rect 309186 37258 309422 37494
rect 309186 30258 309422 30494
rect 309186 23258 309422 23494
rect 309186 16258 309422 16494
rect 309186 9258 309422 9494
rect 309186 2258 309422 2494
rect 309186 -982 309422 -746
rect 309186 -1302 309422 -1066
rect 310918 192325 311154 192561
rect 310918 185325 311154 185561
rect 310918 178325 311154 178561
rect 310918 171325 311154 171561
rect 310918 164325 311154 164561
rect 310918 157325 311154 157561
rect 310918 150325 311154 150561
rect 310918 143325 311154 143561
rect 310918 136325 311154 136561
rect 310918 129325 311154 129561
rect 310918 122325 311154 122561
rect 310918 115325 311154 115561
rect 310918 108325 311154 108561
rect 310918 101325 311154 101561
rect 310918 94325 311154 94561
rect 310918 87325 311154 87561
rect 310918 80325 311154 80561
rect 310918 73325 311154 73561
rect 310918 66325 311154 66561
rect 310918 59325 311154 59561
rect 310918 52325 311154 52561
rect 310918 45325 311154 45561
rect 310918 38325 311154 38561
rect 310918 31325 311154 31561
rect 310918 24325 311154 24561
rect 310918 17325 311154 17561
rect 310918 10325 311154 10561
rect 310918 3325 311154 3561
rect 310918 -1942 311154 -1706
rect 310918 -2262 311154 -2026
rect 316186 191258 316422 191494
rect 316186 184258 316422 184494
rect 316186 177258 316422 177494
rect 316186 170258 316422 170494
rect 316186 163258 316422 163494
rect 316186 156258 316422 156494
rect 316186 149258 316422 149494
rect 316186 142258 316422 142494
rect 316186 135258 316422 135494
rect 316186 128258 316422 128494
rect 316186 121258 316422 121494
rect 316186 114258 316422 114494
rect 316186 107258 316422 107494
rect 316186 100258 316422 100494
rect 316186 93258 316422 93494
rect 316186 86258 316422 86494
rect 316186 79258 316422 79494
rect 316186 72258 316422 72494
rect 316186 65258 316422 65494
rect 316186 58258 316422 58494
rect 316186 51258 316422 51494
rect 316186 44258 316422 44494
rect 316186 37258 316422 37494
rect 316186 30258 316422 30494
rect 316186 23258 316422 23494
rect 316186 16258 316422 16494
rect 316186 9258 316422 9494
rect 316186 2258 316422 2494
rect 316186 -982 316422 -746
rect 316186 -1302 316422 -1066
rect 317918 705962 318154 706198
rect 317918 705642 318154 705878
rect 317918 696325 318154 696561
rect 317918 689325 318154 689561
rect 317918 682325 318154 682561
rect 317918 675325 318154 675561
rect 317918 668325 318154 668561
rect 317918 661325 318154 661561
rect 317918 654325 318154 654561
rect 317918 647325 318154 647561
rect 317918 640325 318154 640561
rect 317918 633325 318154 633561
rect 317918 626325 318154 626561
rect 317918 619325 318154 619561
rect 317918 612325 318154 612561
rect 317918 605325 318154 605561
rect 317918 598325 318154 598561
rect 317918 591325 318154 591561
rect 317918 584325 318154 584561
rect 317918 577325 318154 577561
rect 317918 570325 318154 570561
rect 317918 563325 318154 563561
rect 317918 556325 318154 556561
rect 317918 549325 318154 549561
rect 317918 542325 318154 542561
rect 317918 535325 318154 535561
rect 317918 528325 318154 528561
rect 317918 521325 318154 521561
rect 317918 514325 318154 514561
rect 317918 507325 318154 507561
rect 317918 500325 318154 500561
rect 317918 493325 318154 493561
rect 317918 486325 318154 486561
rect 317918 479325 318154 479561
rect 317918 472325 318154 472561
rect 317918 465325 318154 465561
rect 317918 458325 318154 458561
rect 317918 451325 318154 451561
rect 317918 444325 318154 444561
rect 317918 437325 318154 437561
rect 317918 430325 318154 430561
rect 317918 423325 318154 423561
rect 317918 416325 318154 416561
rect 317918 409325 318154 409561
rect 317918 402325 318154 402561
rect 317918 395325 318154 395561
rect 317918 388325 318154 388561
rect 317918 381325 318154 381561
rect 317918 374325 318154 374561
rect 317918 367325 318154 367561
rect 317918 360325 318154 360561
rect 317918 353325 318154 353561
rect 317918 346325 318154 346561
rect 317918 339325 318154 339561
rect 317918 332325 318154 332561
rect 317918 325325 318154 325561
rect 317918 318325 318154 318561
rect 317918 311325 318154 311561
rect 317918 304325 318154 304561
rect 317918 297325 318154 297561
rect 317918 290325 318154 290561
rect 317918 283325 318154 283561
rect 317918 276325 318154 276561
rect 317918 269325 318154 269561
rect 317918 262325 318154 262561
rect 317918 255325 318154 255561
rect 317918 248325 318154 248561
rect 317918 241325 318154 241561
rect 317918 234325 318154 234561
rect 317918 227325 318154 227561
rect 317918 220325 318154 220561
rect 317918 213325 318154 213561
rect 317918 206325 318154 206561
rect 317918 199325 318154 199561
rect 317918 192325 318154 192561
rect 317918 185325 318154 185561
rect 317918 178325 318154 178561
rect 317918 171325 318154 171561
rect 317918 164325 318154 164561
rect 317918 157325 318154 157561
rect 317918 150325 318154 150561
rect 317918 143325 318154 143561
rect 317918 136325 318154 136561
rect 317918 129325 318154 129561
rect 317918 122325 318154 122561
rect 317918 115325 318154 115561
rect 317918 108325 318154 108561
rect 317918 101325 318154 101561
rect 317918 94325 318154 94561
rect 317918 87325 318154 87561
rect 317918 80325 318154 80561
rect 317918 73325 318154 73561
rect 317918 66325 318154 66561
rect 317918 59325 318154 59561
rect 317918 52325 318154 52561
rect 317918 45325 318154 45561
rect 317918 38325 318154 38561
rect 317918 31325 318154 31561
rect 317918 24325 318154 24561
rect 317918 17325 318154 17561
rect 317918 10325 318154 10561
rect 317918 3325 318154 3561
rect 317918 -1942 318154 -1706
rect 317918 -2262 318154 -2026
rect 323186 705002 323422 705238
rect 323186 704682 323422 704918
rect 323186 695258 323422 695494
rect 323186 688258 323422 688494
rect 323186 681258 323422 681494
rect 323186 674258 323422 674494
rect 323186 667258 323422 667494
rect 323186 660258 323422 660494
rect 323186 653258 323422 653494
rect 323186 646258 323422 646494
rect 323186 639258 323422 639494
rect 323186 632258 323422 632494
rect 323186 625258 323422 625494
rect 323186 618258 323422 618494
rect 323186 611258 323422 611494
rect 323186 604258 323422 604494
rect 323186 597258 323422 597494
rect 323186 590258 323422 590494
rect 323186 583258 323422 583494
rect 323186 576258 323422 576494
rect 323186 569258 323422 569494
rect 323186 562258 323422 562494
rect 323186 555258 323422 555494
rect 323186 548258 323422 548494
rect 323186 541258 323422 541494
rect 323186 534258 323422 534494
rect 323186 527258 323422 527494
rect 323186 520258 323422 520494
rect 323186 513258 323422 513494
rect 323186 506258 323422 506494
rect 323186 499258 323422 499494
rect 323186 492258 323422 492494
rect 323186 485258 323422 485494
rect 323186 478258 323422 478494
rect 323186 471258 323422 471494
rect 323186 464258 323422 464494
rect 323186 457258 323422 457494
rect 323186 450258 323422 450494
rect 323186 443258 323422 443494
rect 323186 436258 323422 436494
rect 323186 429258 323422 429494
rect 323186 422258 323422 422494
rect 323186 415258 323422 415494
rect 323186 408258 323422 408494
rect 323186 401258 323422 401494
rect 323186 394258 323422 394494
rect 323186 387258 323422 387494
rect 323186 380258 323422 380494
rect 323186 373258 323422 373494
rect 323186 366258 323422 366494
rect 323186 359258 323422 359494
rect 323186 352258 323422 352494
rect 323186 345258 323422 345494
rect 323186 338258 323422 338494
rect 323186 331258 323422 331494
rect 323186 324258 323422 324494
rect 323186 317258 323422 317494
rect 323186 310258 323422 310494
rect 323186 303258 323422 303494
rect 323186 296258 323422 296494
rect 323186 289258 323422 289494
rect 323186 282258 323422 282494
rect 323186 275258 323422 275494
rect 323186 268258 323422 268494
rect 323186 261258 323422 261494
rect 323186 254258 323422 254494
rect 323186 247258 323422 247494
rect 323186 240258 323422 240494
rect 323186 233258 323422 233494
rect 323186 226258 323422 226494
rect 323186 219258 323422 219494
rect 323186 212258 323422 212494
rect 323186 205258 323422 205494
rect 323186 198258 323422 198494
rect 323186 191258 323422 191494
rect 323186 184258 323422 184494
rect 323186 177258 323422 177494
rect 323186 170258 323422 170494
rect 323186 163258 323422 163494
rect 323186 156258 323422 156494
rect 323186 149258 323422 149494
rect 323186 142258 323422 142494
rect 323186 135258 323422 135494
rect 323186 128258 323422 128494
rect 323186 121258 323422 121494
rect 323186 114258 323422 114494
rect 323186 107258 323422 107494
rect 323186 100258 323422 100494
rect 323186 93258 323422 93494
rect 323186 86258 323422 86494
rect 323186 79258 323422 79494
rect 323186 72258 323422 72494
rect 323186 65258 323422 65494
rect 323186 58258 323422 58494
rect 323186 51258 323422 51494
rect 323186 44258 323422 44494
rect 323186 37258 323422 37494
rect 323186 30258 323422 30494
rect 323186 23258 323422 23494
rect 323186 16258 323422 16494
rect 323186 9258 323422 9494
rect 323186 2258 323422 2494
rect 323186 -982 323422 -746
rect 323186 -1302 323422 -1066
rect 324918 705962 325154 706198
rect 324918 705642 325154 705878
rect 324918 696325 325154 696561
rect 324918 689325 325154 689561
rect 324918 682325 325154 682561
rect 324918 675325 325154 675561
rect 324918 668325 325154 668561
rect 324918 661325 325154 661561
rect 324918 654325 325154 654561
rect 324918 647325 325154 647561
rect 324918 640325 325154 640561
rect 324918 633325 325154 633561
rect 324918 626325 325154 626561
rect 324918 619325 325154 619561
rect 324918 612325 325154 612561
rect 324918 605325 325154 605561
rect 324918 598325 325154 598561
rect 324918 591325 325154 591561
rect 324918 584325 325154 584561
rect 324918 577325 325154 577561
rect 324918 570325 325154 570561
rect 324918 563325 325154 563561
rect 324918 556325 325154 556561
rect 324918 549325 325154 549561
rect 324918 542325 325154 542561
rect 324918 535325 325154 535561
rect 324918 528325 325154 528561
rect 324918 521325 325154 521561
rect 324918 514325 325154 514561
rect 324918 507325 325154 507561
rect 324918 500325 325154 500561
rect 324918 493325 325154 493561
rect 324918 486325 325154 486561
rect 324918 479325 325154 479561
rect 324918 472325 325154 472561
rect 324918 465325 325154 465561
rect 324918 458325 325154 458561
rect 324918 451325 325154 451561
rect 324918 444325 325154 444561
rect 324918 437325 325154 437561
rect 324918 430325 325154 430561
rect 324918 423325 325154 423561
rect 324918 416325 325154 416561
rect 324918 409325 325154 409561
rect 324918 402325 325154 402561
rect 324918 395325 325154 395561
rect 324918 388325 325154 388561
rect 324918 381325 325154 381561
rect 324918 374325 325154 374561
rect 324918 367325 325154 367561
rect 324918 360325 325154 360561
rect 324918 353325 325154 353561
rect 324918 346325 325154 346561
rect 324918 339325 325154 339561
rect 324918 332325 325154 332561
rect 324918 325325 325154 325561
rect 324918 318325 325154 318561
rect 324918 311325 325154 311561
rect 324918 304325 325154 304561
rect 324918 297325 325154 297561
rect 324918 290325 325154 290561
rect 324918 283325 325154 283561
rect 324918 276325 325154 276561
rect 324918 269325 325154 269561
rect 324918 262325 325154 262561
rect 324918 255325 325154 255561
rect 324918 248325 325154 248561
rect 324918 241325 325154 241561
rect 324918 234325 325154 234561
rect 324918 227325 325154 227561
rect 324918 220325 325154 220561
rect 324918 213325 325154 213561
rect 324918 206325 325154 206561
rect 324918 199325 325154 199561
rect 324918 192325 325154 192561
rect 324918 185325 325154 185561
rect 324918 178325 325154 178561
rect 324918 171325 325154 171561
rect 324918 164325 325154 164561
rect 324918 157325 325154 157561
rect 324918 150325 325154 150561
rect 324918 143325 325154 143561
rect 324918 136325 325154 136561
rect 324918 129325 325154 129561
rect 324918 122325 325154 122561
rect 324918 115325 325154 115561
rect 324918 108325 325154 108561
rect 324918 101325 325154 101561
rect 324918 94325 325154 94561
rect 324918 87325 325154 87561
rect 324918 80325 325154 80561
rect 324918 73325 325154 73561
rect 324918 66325 325154 66561
rect 324918 59325 325154 59561
rect 324918 52325 325154 52561
rect 324918 45325 325154 45561
rect 324918 38325 325154 38561
rect 324918 31325 325154 31561
rect 324918 24325 325154 24561
rect 324918 17325 325154 17561
rect 324918 10325 325154 10561
rect 324918 3325 325154 3561
rect 324918 -1942 325154 -1706
rect 324918 -2262 325154 -2026
rect 330186 705002 330422 705238
rect 330186 704682 330422 704918
rect 330186 695258 330422 695494
rect 330186 688258 330422 688494
rect 330186 681258 330422 681494
rect 330186 674258 330422 674494
rect 330186 667258 330422 667494
rect 330186 660258 330422 660494
rect 330186 653258 330422 653494
rect 330186 646258 330422 646494
rect 330186 639258 330422 639494
rect 330186 632258 330422 632494
rect 330186 625258 330422 625494
rect 330186 618258 330422 618494
rect 330186 611258 330422 611494
rect 330186 604258 330422 604494
rect 330186 597258 330422 597494
rect 330186 590258 330422 590494
rect 330186 583258 330422 583494
rect 330186 576258 330422 576494
rect 330186 569258 330422 569494
rect 330186 562258 330422 562494
rect 330186 555258 330422 555494
rect 330186 548258 330422 548494
rect 330186 541258 330422 541494
rect 330186 534258 330422 534494
rect 330186 527258 330422 527494
rect 330186 520258 330422 520494
rect 330186 513258 330422 513494
rect 330186 506258 330422 506494
rect 330186 499258 330422 499494
rect 330186 492258 330422 492494
rect 330186 485258 330422 485494
rect 330186 478258 330422 478494
rect 330186 471258 330422 471494
rect 330186 464258 330422 464494
rect 330186 457258 330422 457494
rect 330186 450258 330422 450494
rect 330186 443258 330422 443494
rect 330186 436258 330422 436494
rect 330186 429258 330422 429494
rect 330186 422258 330422 422494
rect 330186 415258 330422 415494
rect 330186 408258 330422 408494
rect 330186 401258 330422 401494
rect 330186 394258 330422 394494
rect 330186 387258 330422 387494
rect 330186 380258 330422 380494
rect 330186 373258 330422 373494
rect 330186 366258 330422 366494
rect 330186 359258 330422 359494
rect 330186 352258 330422 352494
rect 330186 345258 330422 345494
rect 330186 338258 330422 338494
rect 330186 331258 330422 331494
rect 330186 324258 330422 324494
rect 330186 317258 330422 317494
rect 330186 310258 330422 310494
rect 330186 303258 330422 303494
rect 330186 296258 330422 296494
rect 330186 289258 330422 289494
rect 330186 282258 330422 282494
rect 330186 275258 330422 275494
rect 330186 268258 330422 268494
rect 330186 261258 330422 261494
rect 330186 254258 330422 254494
rect 330186 247258 330422 247494
rect 330186 240258 330422 240494
rect 330186 233258 330422 233494
rect 330186 226258 330422 226494
rect 330186 219258 330422 219494
rect 330186 212258 330422 212494
rect 330186 205258 330422 205494
rect 330186 198258 330422 198494
rect 330186 191258 330422 191494
rect 330186 184258 330422 184494
rect 330186 177258 330422 177494
rect 330186 170258 330422 170494
rect 330186 163258 330422 163494
rect 330186 156258 330422 156494
rect 330186 149258 330422 149494
rect 330186 142258 330422 142494
rect 330186 135258 330422 135494
rect 330186 128258 330422 128494
rect 330186 121258 330422 121494
rect 330186 114258 330422 114494
rect 330186 107258 330422 107494
rect 330186 100258 330422 100494
rect 330186 93258 330422 93494
rect 330186 86258 330422 86494
rect 330186 79258 330422 79494
rect 330186 72258 330422 72494
rect 330186 65258 330422 65494
rect 330186 58258 330422 58494
rect 330186 51258 330422 51494
rect 330186 44258 330422 44494
rect 330186 37258 330422 37494
rect 330186 30258 330422 30494
rect 330186 23258 330422 23494
rect 330186 16258 330422 16494
rect 330186 9258 330422 9494
rect 330186 2258 330422 2494
rect 330186 -982 330422 -746
rect 330186 -1302 330422 -1066
rect 331918 705962 332154 706198
rect 331918 705642 332154 705878
rect 331918 696325 332154 696561
rect 331918 689325 332154 689561
rect 331918 682325 332154 682561
rect 331918 675325 332154 675561
rect 331918 668325 332154 668561
rect 331918 661325 332154 661561
rect 331918 654325 332154 654561
rect 331918 647325 332154 647561
rect 331918 640325 332154 640561
rect 331918 633325 332154 633561
rect 331918 626325 332154 626561
rect 331918 619325 332154 619561
rect 331918 612325 332154 612561
rect 331918 605325 332154 605561
rect 331918 598325 332154 598561
rect 331918 591325 332154 591561
rect 331918 584325 332154 584561
rect 331918 577325 332154 577561
rect 331918 570325 332154 570561
rect 331918 563325 332154 563561
rect 331918 556325 332154 556561
rect 331918 549325 332154 549561
rect 331918 542325 332154 542561
rect 331918 535325 332154 535561
rect 331918 528325 332154 528561
rect 331918 521325 332154 521561
rect 331918 514325 332154 514561
rect 331918 507325 332154 507561
rect 331918 500325 332154 500561
rect 331918 493325 332154 493561
rect 331918 486325 332154 486561
rect 331918 479325 332154 479561
rect 331918 472325 332154 472561
rect 331918 465325 332154 465561
rect 331918 458325 332154 458561
rect 331918 451325 332154 451561
rect 331918 444325 332154 444561
rect 331918 437325 332154 437561
rect 331918 430325 332154 430561
rect 331918 423325 332154 423561
rect 331918 416325 332154 416561
rect 331918 409325 332154 409561
rect 331918 402325 332154 402561
rect 331918 395325 332154 395561
rect 331918 388325 332154 388561
rect 331918 381325 332154 381561
rect 331918 374325 332154 374561
rect 331918 367325 332154 367561
rect 331918 360325 332154 360561
rect 331918 353325 332154 353561
rect 331918 346325 332154 346561
rect 331918 339325 332154 339561
rect 331918 332325 332154 332561
rect 331918 325325 332154 325561
rect 331918 318325 332154 318561
rect 331918 311325 332154 311561
rect 331918 304325 332154 304561
rect 331918 297325 332154 297561
rect 331918 290325 332154 290561
rect 331918 283325 332154 283561
rect 331918 276325 332154 276561
rect 331918 269325 332154 269561
rect 331918 262325 332154 262561
rect 331918 255325 332154 255561
rect 331918 248325 332154 248561
rect 331918 241325 332154 241561
rect 331918 234325 332154 234561
rect 331918 227325 332154 227561
rect 331918 220325 332154 220561
rect 331918 213325 332154 213561
rect 331918 206325 332154 206561
rect 331918 199325 332154 199561
rect 331918 192325 332154 192561
rect 331918 185325 332154 185561
rect 331918 178325 332154 178561
rect 331918 171325 332154 171561
rect 331918 164325 332154 164561
rect 331918 157325 332154 157561
rect 331918 150325 332154 150561
rect 331918 143325 332154 143561
rect 331918 136325 332154 136561
rect 331918 129325 332154 129561
rect 331918 122325 332154 122561
rect 331918 115325 332154 115561
rect 331918 108325 332154 108561
rect 331918 101325 332154 101561
rect 331918 94325 332154 94561
rect 331918 87325 332154 87561
rect 331918 80325 332154 80561
rect 331918 73325 332154 73561
rect 331918 66325 332154 66561
rect 331918 59325 332154 59561
rect 331918 52325 332154 52561
rect 331918 45325 332154 45561
rect 331918 38325 332154 38561
rect 331918 31325 332154 31561
rect 331918 24325 332154 24561
rect 331918 17325 332154 17561
rect 331918 10325 332154 10561
rect 331918 3325 332154 3561
rect 331918 -1942 332154 -1706
rect 331918 -2262 332154 -2026
rect 337186 705002 337422 705238
rect 337186 704682 337422 704918
rect 337186 695258 337422 695494
rect 337186 688258 337422 688494
rect 337186 681258 337422 681494
rect 337186 674258 337422 674494
rect 337186 667258 337422 667494
rect 337186 660258 337422 660494
rect 337186 653258 337422 653494
rect 337186 646258 337422 646494
rect 337186 639258 337422 639494
rect 337186 632258 337422 632494
rect 337186 625258 337422 625494
rect 337186 618258 337422 618494
rect 337186 611258 337422 611494
rect 337186 604258 337422 604494
rect 337186 597258 337422 597494
rect 337186 590258 337422 590494
rect 337186 583258 337422 583494
rect 337186 576258 337422 576494
rect 337186 569258 337422 569494
rect 337186 562258 337422 562494
rect 337186 555258 337422 555494
rect 337186 548258 337422 548494
rect 337186 541258 337422 541494
rect 337186 534258 337422 534494
rect 337186 527258 337422 527494
rect 337186 520258 337422 520494
rect 337186 513258 337422 513494
rect 337186 506258 337422 506494
rect 337186 499258 337422 499494
rect 337186 492258 337422 492494
rect 337186 485258 337422 485494
rect 337186 478258 337422 478494
rect 337186 471258 337422 471494
rect 337186 464258 337422 464494
rect 337186 457258 337422 457494
rect 337186 450258 337422 450494
rect 337186 443258 337422 443494
rect 337186 436258 337422 436494
rect 337186 429258 337422 429494
rect 337186 422258 337422 422494
rect 337186 415258 337422 415494
rect 337186 408258 337422 408494
rect 337186 401258 337422 401494
rect 337186 394258 337422 394494
rect 337186 387258 337422 387494
rect 337186 380258 337422 380494
rect 337186 373258 337422 373494
rect 337186 366258 337422 366494
rect 337186 359258 337422 359494
rect 337186 352258 337422 352494
rect 337186 345258 337422 345494
rect 337186 338258 337422 338494
rect 337186 331258 337422 331494
rect 337186 324258 337422 324494
rect 337186 317258 337422 317494
rect 337186 310258 337422 310494
rect 337186 303258 337422 303494
rect 337186 296258 337422 296494
rect 337186 289258 337422 289494
rect 337186 282258 337422 282494
rect 337186 275258 337422 275494
rect 337186 268258 337422 268494
rect 337186 261258 337422 261494
rect 337186 254258 337422 254494
rect 337186 247258 337422 247494
rect 337186 240258 337422 240494
rect 337186 233258 337422 233494
rect 337186 226258 337422 226494
rect 337186 219258 337422 219494
rect 337186 212258 337422 212494
rect 337186 205258 337422 205494
rect 337186 198258 337422 198494
rect 337186 191258 337422 191494
rect 337186 184258 337422 184494
rect 337186 177258 337422 177494
rect 337186 170258 337422 170494
rect 337186 163258 337422 163494
rect 337186 156258 337422 156494
rect 337186 149258 337422 149494
rect 337186 142258 337422 142494
rect 337186 135258 337422 135494
rect 337186 128258 337422 128494
rect 337186 121258 337422 121494
rect 337186 114258 337422 114494
rect 337186 107258 337422 107494
rect 337186 100258 337422 100494
rect 337186 93258 337422 93494
rect 337186 86258 337422 86494
rect 337186 79258 337422 79494
rect 337186 72258 337422 72494
rect 337186 65258 337422 65494
rect 337186 58258 337422 58494
rect 337186 51258 337422 51494
rect 337186 44258 337422 44494
rect 337186 37258 337422 37494
rect 337186 30258 337422 30494
rect 337186 23258 337422 23494
rect 337186 16258 337422 16494
rect 337186 9258 337422 9494
rect 337186 2258 337422 2494
rect 337186 -982 337422 -746
rect 337186 -1302 337422 -1066
rect 338918 705962 339154 706198
rect 338918 705642 339154 705878
rect 338918 696325 339154 696561
rect 338918 689325 339154 689561
rect 338918 682325 339154 682561
rect 338918 675325 339154 675561
rect 338918 668325 339154 668561
rect 338918 661325 339154 661561
rect 338918 654325 339154 654561
rect 338918 647325 339154 647561
rect 338918 640325 339154 640561
rect 338918 633325 339154 633561
rect 338918 626325 339154 626561
rect 338918 619325 339154 619561
rect 338918 612325 339154 612561
rect 338918 605325 339154 605561
rect 338918 598325 339154 598561
rect 338918 591325 339154 591561
rect 338918 584325 339154 584561
rect 338918 577325 339154 577561
rect 338918 570325 339154 570561
rect 338918 563325 339154 563561
rect 338918 556325 339154 556561
rect 338918 549325 339154 549561
rect 338918 542325 339154 542561
rect 338918 535325 339154 535561
rect 338918 528325 339154 528561
rect 338918 521325 339154 521561
rect 338918 514325 339154 514561
rect 338918 507325 339154 507561
rect 338918 500325 339154 500561
rect 338918 493325 339154 493561
rect 338918 486325 339154 486561
rect 338918 479325 339154 479561
rect 338918 472325 339154 472561
rect 338918 465325 339154 465561
rect 338918 458325 339154 458561
rect 338918 451325 339154 451561
rect 338918 444325 339154 444561
rect 338918 437325 339154 437561
rect 338918 430325 339154 430561
rect 338918 423325 339154 423561
rect 338918 416325 339154 416561
rect 338918 409325 339154 409561
rect 338918 402325 339154 402561
rect 338918 395325 339154 395561
rect 338918 388325 339154 388561
rect 338918 381325 339154 381561
rect 338918 374325 339154 374561
rect 338918 367325 339154 367561
rect 338918 360325 339154 360561
rect 338918 353325 339154 353561
rect 338918 346325 339154 346561
rect 338918 339325 339154 339561
rect 338918 332325 339154 332561
rect 338918 325325 339154 325561
rect 338918 318325 339154 318561
rect 338918 311325 339154 311561
rect 338918 304325 339154 304561
rect 338918 297325 339154 297561
rect 338918 290325 339154 290561
rect 338918 283325 339154 283561
rect 338918 276325 339154 276561
rect 338918 269325 339154 269561
rect 338918 262325 339154 262561
rect 338918 255325 339154 255561
rect 338918 248325 339154 248561
rect 338918 241325 339154 241561
rect 338918 234325 339154 234561
rect 338918 227325 339154 227561
rect 338918 220325 339154 220561
rect 338918 213325 339154 213561
rect 338918 206325 339154 206561
rect 338918 199325 339154 199561
rect 338918 192325 339154 192561
rect 338918 185325 339154 185561
rect 338918 178325 339154 178561
rect 338918 171325 339154 171561
rect 338918 164325 339154 164561
rect 338918 157325 339154 157561
rect 338918 150325 339154 150561
rect 338918 143325 339154 143561
rect 338918 136325 339154 136561
rect 338918 129325 339154 129561
rect 338918 122325 339154 122561
rect 338918 115325 339154 115561
rect 338918 108325 339154 108561
rect 338918 101325 339154 101561
rect 338918 94325 339154 94561
rect 338918 87325 339154 87561
rect 338918 80325 339154 80561
rect 338918 73325 339154 73561
rect 338918 66325 339154 66561
rect 338918 59325 339154 59561
rect 338918 52325 339154 52561
rect 338918 45325 339154 45561
rect 338918 38325 339154 38561
rect 338918 31325 339154 31561
rect 338918 24325 339154 24561
rect 338918 17325 339154 17561
rect 338918 10325 339154 10561
rect 338918 3325 339154 3561
rect 338918 -1942 339154 -1706
rect 338918 -2262 339154 -2026
rect 344186 705002 344422 705238
rect 344186 704682 344422 704918
rect 344186 695258 344422 695494
rect 344186 688258 344422 688494
rect 344186 681258 344422 681494
rect 344186 674258 344422 674494
rect 344186 667258 344422 667494
rect 344186 660258 344422 660494
rect 344186 653258 344422 653494
rect 344186 646258 344422 646494
rect 344186 639258 344422 639494
rect 344186 632258 344422 632494
rect 344186 625258 344422 625494
rect 344186 618258 344422 618494
rect 344186 611258 344422 611494
rect 344186 604258 344422 604494
rect 344186 597258 344422 597494
rect 344186 590258 344422 590494
rect 344186 583258 344422 583494
rect 344186 576258 344422 576494
rect 344186 569258 344422 569494
rect 344186 562258 344422 562494
rect 344186 555258 344422 555494
rect 344186 548258 344422 548494
rect 344186 541258 344422 541494
rect 344186 534258 344422 534494
rect 344186 527258 344422 527494
rect 344186 520258 344422 520494
rect 344186 513258 344422 513494
rect 344186 506258 344422 506494
rect 344186 499258 344422 499494
rect 344186 492258 344422 492494
rect 344186 485258 344422 485494
rect 344186 478258 344422 478494
rect 344186 471258 344422 471494
rect 344186 464258 344422 464494
rect 344186 457258 344422 457494
rect 344186 450258 344422 450494
rect 344186 443258 344422 443494
rect 344186 436258 344422 436494
rect 344186 429258 344422 429494
rect 344186 422258 344422 422494
rect 344186 415258 344422 415494
rect 344186 408258 344422 408494
rect 344186 401258 344422 401494
rect 344186 394258 344422 394494
rect 344186 387258 344422 387494
rect 344186 380258 344422 380494
rect 344186 373258 344422 373494
rect 344186 366258 344422 366494
rect 344186 359258 344422 359494
rect 344186 352258 344422 352494
rect 344186 345258 344422 345494
rect 344186 338258 344422 338494
rect 344186 331258 344422 331494
rect 344186 324258 344422 324494
rect 344186 317258 344422 317494
rect 344186 310258 344422 310494
rect 344186 303258 344422 303494
rect 344186 296258 344422 296494
rect 344186 289258 344422 289494
rect 344186 282258 344422 282494
rect 344186 275258 344422 275494
rect 344186 268258 344422 268494
rect 344186 261258 344422 261494
rect 344186 254258 344422 254494
rect 344186 247258 344422 247494
rect 344186 240258 344422 240494
rect 344186 233258 344422 233494
rect 344186 226258 344422 226494
rect 344186 219258 344422 219494
rect 344186 212258 344422 212494
rect 344186 205258 344422 205494
rect 344186 198258 344422 198494
rect 344186 191258 344422 191494
rect 344186 184258 344422 184494
rect 344186 177258 344422 177494
rect 344186 170258 344422 170494
rect 344186 163258 344422 163494
rect 344186 156258 344422 156494
rect 344186 149258 344422 149494
rect 344186 142258 344422 142494
rect 344186 135258 344422 135494
rect 344186 128258 344422 128494
rect 344186 121258 344422 121494
rect 344186 114258 344422 114494
rect 344186 107258 344422 107494
rect 344186 100258 344422 100494
rect 344186 93258 344422 93494
rect 344186 86258 344422 86494
rect 344186 79258 344422 79494
rect 344186 72258 344422 72494
rect 344186 65258 344422 65494
rect 344186 58258 344422 58494
rect 344186 51258 344422 51494
rect 344186 44258 344422 44494
rect 344186 37258 344422 37494
rect 344186 30258 344422 30494
rect 344186 23258 344422 23494
rect 344186 16258 344422 16494
rect 344186 9258 344422 9494
rect 344186 2258 344422 2494
rect 344186 -982 344422 -746
rect 344186 -1302 344422 -1066
rect 345918 705962 346154 706198
rect 345918 705642 346154 705878
rect 345918 696325 346154 696561
rect 345918 689325 346154 689561
rect 345918 682325 346154 682561
rect 345918 675325 346154 675561
rect 345918 668325 346154 668561
rect 345918 661325 346154 661561
rect 345918 654325 346154 654561
rect 345918 647325 346154 647561
rect 345918 640325 346154 640561
rect 345918 633325 346154 633561
rect 345918 626325 346154 626561
rect 345918 619325 346154 619561
rect 345918 612325 346154 612561
rect 345918 605325 346154 605561
rect 345918 598325 346154 598561
rect 345918 591325 346154 591561
rect 345918 584325 346154 584561
rect 345918 577325 346154 577561
rect 345918 570325 346154 570561
rect 345918 563325 346154 563561
rect 345918 556325 346154 556561
rect 345918 549325 346154 549561
rect 345918 542325 346154 542561
rect 345918 535325 346154 535561
rect 345918 528325 346154 528561
rect 345918 521325 346154 521561
rect 345918 514325 346154 514561
rect 345918 507325 346154 507561
rect 345918 500325 346154 500561
rect 345918 493325 346154 493561
rect 345918 486325 346154 486561
rect 345918 479325 346154 479561
rect 345918 472325 346154 472561
rect 345918 465325 346154 465561
rect 345918 458325 346154 458561
rect 345918 451325 346154 451561
rect 345918 444325 346154 444561
rect 345918 437325 346154 437561
rect 345918 430325 346154 430561
rect 345918 423325 346154 423561
rect 345918 416325 346154 416561
rect 345918 409325 346154 409561
rect 345918 402325 346154 402561
rect 345918 395325 346154 395561
rect 345918 388325 346154 388561
rect 345918 381325 346154 381561
rect 345918 374325 346154 374561
rect 345918 367325 346154 367561
rect 345918 360325 346154 360561
rect 345918 353325 346154 353561
rect 345918 346325 346154 346561
rect 345918 339325 346154 339561
rect 345918 332325 346154 332561
rect 345918 325325 346154 325561
rect 345918 318325 346154 318561
rect 345918 311325 346154 311561
rect 345918 304325 346154 304561
rect 345918 297325 346154 297561
rect 345918 290325 346154 290561
rect 345918 283325 346154 283561
rect 345918 276325 346154 276561
rect 345918 269325 346154 269561
rect 345918 262325 346154 262561
rect 345918 255325 346154 255561
rect 345918 248325 346154 248561
rect 345918 241325 346154 241561
rect 345918 234325 346154 234561
rect 345918 227325 346154 227561
rect 345918 220325 346154 220561
rect 345918 213325 346154 213561
rect 345918 206325 346154 206561
rect 345918 199325 346154 199561
rect 345918 192325 346154 192561
rect 345918 185325 346154 185561
rect 345918 178325 346154 178561
rect 345918 171325 346154 171561
rect 345918 164325 346154 164561
rect 345918 157325 346154 157561
rect 345918 150325 346154 150561
rect 345918 143325 346154 143561
rect 345918 136325 346154 136561
rect 345918 129325 346154 129561
rect 345918 122325 346154 122561
rect 345918 115325 346154 115561
rect 345918 108325 346154 108561
rect 345918 101325 346154 101561
rect 345918 94325 346154 94561
rect 345918 87325 346154 87561
rect 345918 80325 346154 80561
rect 345918 73325 346154 73561
rect 345918 66325 346154 66561
rect 345918 59325 346154 59561
rect 345918 52325 346154 52561
rect 345918 45325 346154 45561
rect 345918 38325 346154 38561
rect 345918 31325 346154 31561
rect 345918 24325 346154 24561
rect 345918 17325 346154 17561
rect 345918 10325 346154 10561
rect 345918 3325 346154 3561
rect 345918 -1942 346154 -1706
rect 345918 -2262 346154 -2026
rect 351186 705002 351422 705238
rect 351186 704682 351422 704918
rect 351186 695258 351422 695494
rect 351186 688258 351422 688494
rect 351186 681258 351422 681494
rect 351186 674258 351422 674494
rect 351186 667258 351422 667494
rect 351186 660258 351422 660494
rect 351186 653258 351422 653494
rect 351186 646258 351422 646494
rect 351186 639258 351422 639494
rect 351186 632258 351422 632494
rect 351186 625258 351422 625494
rect 351186 618258 351422 618494
rect 351186 611258 351422 611494
rect 351186 604258 351422 604494
rect 351186 597258 351422 597494
rect 351186 590258 351422 590494
rect 351186 583258 351422 583494
rect 351186 576258 351422 576494
rect 351186 569258 351422 569494
rect 351186 562258 351422 562494
rect 351186 555258 351422 555494
rect 351186 548258 351422 548494
rect 351186 541258 351422 541494
rect 351186 534258 351422 534494
rect 351186 527258 351422 527494
rect 351186 520258 351422 520494
rect 351186 513258 351422 513494
rect 351186 506258 351422 506494
rect 351186 499258 351422 499494
rect 351186 492258 351422 492494
rect 351186 485258 351422 485494
rect 351186 478258 351422 478494
rect 351186 471258 351422 471494
rect 351186 464258 351422 464494
rect 351186 457258 351422 457494
rect 351186 450258 351422 450494
rect 351186 443258 351422 443494
rect 351186 436258 351422 436494
rect 351186 429258 351422 429494
rect 351186 422258 351422 422494
rect 351186 415258 351422 415494
rect 351186 408258 351422 408494
rect 351186 401258 351422 401494
rect 351186 394258 351422 394494
rect 351186 387258 351422 387494
rect 351186 380258 351422 380494
rect 351186 373258 351422 373494
rect 351186 366258 351422 366494
rect 351186 359258 351422 359494
rect 351186 352258 351422 352494
rect 351186 345258 351422 345494
rect 351186 338258 351422 338494
rect 351186 331258 351422 331494
rect 351186 324258 351422 324494
rect 351186 317258 351422 317494
rect 351186 310258 351422 310494
rect 351186 303258 351422 303494
rect 351186 296258 351422 296494
rect 351186 289258 351422 289494
rect 351186 282258 351422 282494
rect 351186 275258 351422 275494
rect 351186 268258 351422 268494
rect 351186 261258 351422 261494
rect 351186 254258 351422 254494
rect 351186 247258 351422 247494
rect 351186 240258 351422 240494
rect 351186 233258 351422 233494
rect 351186 226258 351422 226494
rect 351186 219258 351422 219494
rect 351186 212258 351422 212494
rect 351186 205258 351422 205494
rect 351186 198258 351422 198494
rect 351186 191258 351422 191494
rect 351186 184258 351422 184494
rect 351186 177258 351422 177494
rect 351186 170258 351422 170494
rect 351186 163258 351422 163494
rect 351186 156258 351422 156494
rect 351186 149258 351422 149494
rect 351186 142258 351422 142494
rect 351186 135258 351422 135494
rect 351186 128258 351422 128494
rect 351186 121258 351422 121494
rect 351186 114258 351422 114494
rect 351186 107258 351422 107494
rect 351186 100258 351422 100494
rect 351186 93258 351422 93494
rect 351186 86258 351422 86494
rect 351186 79258 351422 79494
rect 351186 72258 351422 72494
rect 351186 65258 351422 65494
rect 351186 58258 351422 58494
rect 351186 51258 351422 51494
rect 351186 44258 351422 44494
rect 351186 37258 351422 37494
rect 351186 30258 351422 30494
rect 351186 23258 351422 23494
rect 351186 16258 351422 16494
rect 351186 9258 351422 9494
rect 351186 2258 351422 2494
rect 351186 -982 351422 -746
rect 351186 -1302 351422 -1066
rect 352918 705962 353154 706198
rect 352918 705642 353154 705878
rect 352918 696325 353154 696561
rect 352918 689325 353154 689561
rect 352918 682325 353154 682561
rect 352918 675325 353154 675561
rect 352918 668325 353154 668561
rect 352918 661325 353154 661561
rect 352918 654325 353154 654561
rect 352918 647325 353154 647561
rect 352918 640325 353154 640561
rect 352918 633325 353154 633561
rect 352918 626325 353154 626561
rect 352918 619325 353154 619561
rect 352918 612325 353154 612561
rect 352918 605325 353154 605561
rect 352918 598325 353154 598561
rect 352918 591325 353154 591561
rect 352918 584325 353154 584561
rect 352918 577325 353154 577561
rect 352918 570325 353154 570561
rect 352918 563325 353154 563561
rect 352918 556325 353154 556561
rect 352918 549325 353154 549561
rect 352918 542325 353154 542561
rect 352918 535325 353154 535561
rect 352918 528325 353154 528561
rect 352918 521325 353154 521561
rect 352918 514325 353154 514561
rect 352918 507325 353154 507561
rect 352918 500325 353154 500561
rect 352918 493325 353154 493561
rect 352918 486325 353154 486561
rect 352918 479325 353154 479561
rect 352918 472325 353154 472561
rect 352918 465325 353154 465561
rect 352918 458325 353154 458561
rect 352918 451325 353154 451561
rect 352918 444325 353154 444561
rect 352918 437325 353154 437561
rect 352918 430325 353154 430561
rect 352918 423325 353154 423561
rect 352918 416325 353154 416561
rect 352918 409325 353154 409561
rect 352918 402325 353154 402561
rect 352918 395325 353154 395561
rect 352918 388325 353154 388561
rect 352918 381325 353154 381561
rect 352918 374325 353154 374561
rect 352918 367325 353154 367561
rect 352918 360325 353154 360561
rect 352918 353325 353154 353561
rect 352918 346325 353154 346561
rect 352918 339325 353154 339561
rect 352918 332325 353154 332561
rect 352918 325325 353154 325561
rect 352918 318325 353154 318561
rect 352918 311325 353154 311561
rect 352918 304325 353154 304561
rect 352918 297325 353154 297561
rect 352918 290325 353154 290561
rect 352918 283325 353154 283561
rect 352918 276325 353154 276561
rect 352918 269325 353154 269561
rect 352918 262325 353154 262561
rect 352918 255325 353154 255561
rect 352918 248325 353154 248561
rect 352918 241325 353154 241561
rect 352918 234325 353154 234561
rect 352918 227325 353154 227561
rect 352918 220325 353154 220561
rect 352918 213325 353154 213561
rect 352918 206325 353154 206561
rect 352918 199325 353154 199561
rect 352918 192325 353154 192561
rect 352918 185325 353154 185561
rect 352918 178325 353154 178561
rect 352918 171325 353154 171561
rect 352918 164325 353154 164561
rect 352918 157325 353154 157561
rect 352918 150325 353154 150561
rect 352918 143325 353154 143561
rect 352918 136325 353154 136561
rect 352918 129325 353154 129561
rect 352918 122325 353154 122561
rect 352918 115325 353154 115561
rect 352918 108325 353154 108561
rect 352918 101325 353154 101561
rect 352918 94325 353154 94561
rect 352918 87325 353154 87561
rect 352918 80325 353154 80561
rect 352918 73325 353154 73561
rect 352918 66325 353154 66561
rect 352918 59325 353154 59561
rect 352918 52325 353154 52561
rect 352918 45325 353154 45561
rect 352918 38325 353154 38561
rect 352918 31325 353154 31561
rect 352918 24325 353154 24561
rect 352918 17325 353154 17561
rect 352918 10325 353154 10561
rect 352918 3325 353154 3561
rect 352918 -1942 353154 -1706
rect 352918 -2262 353154 -2026
rect 358186 705002 358422 705238
rect 358186 704682 358422 704918
rect 358186 695258 358422 695494
rect 358186 688258 358422 688494
rect 358186 681258 358422 681494
rect 358186 674258 358422 674494
rect 358186 667258 358422 667494
rect 358186 660258 358422 660494
rect 358186 653258 358422 653494
rect 358186 646258 358422 646494
rect 358186 639258 358422 639494
rect 358186 632258 358422 632494
rect 358186 625258 358422 625494
rect 358186 618258 358422 618494
rect 358186 611258 358422 611494
rect 358186 604258 358422 604494
rect 358186 597258 358422 597494
rect 358186 590258 358422 590494
rect 358186 583258 358422 583494
rect 358186 576258 358422 576494
rect 358186 569258 358422 569494
rect 358186 562258 358422 562494
rect 358186 555258 358422 555494
rect 358186 548258 358422 548494
rect 358186 541258 358422 541494
rect 358186 534258 358422 534494
rect 358186 527258 358422 527494
rect 358186 520258 358422 520494
rect 358186 513258 358422 513494
rect 358186 506258 358422 506494
rect 358186 499258 358422 499494
rect 358186 492258 358422 492494
rect 358186 485258 358422 485494
rect 358186 478258 358422 478494
rect 358186 471258 358422 471494
rect 358186 464258 358422 464494
rect 358186 457258 358422 457494
rect 358186 450258 358422 450494
rect 358186 443258 358422 443494
rect 358186 436258 358422 436494
rect 358186 429258 358422 429494
rect 358186 422258 358422 422494
rect 358186 415258 358422 415494
rect 358186 408258 358422 408494
rect 358186 401258 358422 401494
rect 358186 394258 358422 394494
rect 358186 387258 358422 387494
rect 358186 380258 358422 380494
rect 358186 373258 358422 373494
rect 358186 366258 358422 366494
rect 358186 359258 358422 359494
rect 358186 352258 358422 352494
rect 358186 345258 358422 345494
rect 358186 338258 358422 338494
rect 358186 331258 358422 331494
rect 358186 324258 358422 324494
rect 358186 317258 358422 317494
rect 358186 310258 358422 310494
rect 358186 303258 358422 303494
rect 358186 296258 358422 296494
rect 358186 289258 358422 289494
rect 358186 282258 358422 282494
rect 358186 275258 358422 275494
rect 358186 268258 358422 268494
rect 358186 261258 358422 261494
rect 358186 254258 358422 254494
rect 358186 247258 358422 247494
rect 358186 240258 358422 240494
rect 358186 233258 358422 233494
rect 358186 226258 358422 226494
rect 358186 219258 358422 219494
rect 358186 212258 358422 212494
rect 358186 205258 358422 205494
rect 358186 198258 358422 198494
rect 358186 191258 358422 191494
rect 358186 184258 358422 184494
rect 358186 177258 358422 177494
rect 358186 170258 358422 170494
rect 358186 163258 358422 163494
rect 358186 156258 358422 156494
rect 358186 149258 358422 149494
rect 358186 142258 358422 142494
rect 358186 135258 358422 135494
rect 358186 128258 358422 128494
rect 358186 121258 358422 121494
rect 358186 114258 358422 114494
rect 358186 107258 358422 107494
rect 358186 100258 358422 100494
rect 358186 93258 358422 93494
rect 358186 86258 358422 86494
rect 358186 79258 358422 79494
rect 358186 72258 358422 72494
rect 358186 65258 358422 65494
rect 358186 58258 358422 58494
rect 358186 51258 358422 51494
rect 358186 44258 358422 44494
rect 358186 37258 358422 37494
rect 358186 30258 358422 30494
rect 358186 23258 358422 23494
rect 358186 16258 358422 16494
rect 358186 9258 358422 9494
rect 358186 2258 358422 2494
rect 358186 -982 358422 -746
rect 358186 -1302 358422 -1066
rect 359918 705962 360154 706198
rect 359918 705642 360154 705878
rect 359918 696325 360154 696561
rect 359918 689325 360154 689561
rect 359918 682325 360154 682561
rect 359918 675325 360154 675561
rect 359918 668325 360154 668561
rect 359918 661325 360154 661561
rect 359918 654325 360154 654561
rect 359918 647325 360154 647561
rect 359918 640325 360154 640561
rect 359918 633325 360154 633561
rect 359918 626325 360154 626561
rect 359918 619325 360154 619561
rect 359918 612325 360154 612561
rect 359918 605325 360154 605561
rect 359918 598325 360154 598561
rect 359918 591325 360154 591561
rect 359918 584325 360154 584561
rect 359918 577325 360154 577561
rect 359918 570325 360154 570561
rect 359918 563325 360154 563561
rect 359918 556325 360154 556561
rect 359918 549325 360154 549561
rect 359918 542325 360154 542561
rect 359918 535325 360154 535561
rect 359918 528325 360154 528561
rect 359918 521325 360154 521561
rect 359918 514325 360154 514561
rect 359918 507325 360154 507561
rect 359918 500325 360154 500561
rect 359918 493325 360154 493561
rect 359918 486325 360154 486561
rect 359918 479325 360154 479561
rect 359918 472325 360154 472561
rect 359918 465325 360154 465561
rect 359918 458325 360154 458561
rect 359918 451325 360154 451561
rect 359918 444325 360154 444561
rect 359918 437325 360154 437561
rect 359918 430325 360154 430561
rect 359918 423325 360154 423561
rect 359918 416325 360154 416561
rect 359918 409325 360154 409561
rect 359918 402325 360154 402561
rect 359918 395325 360154 395561
rect 359918 388325 360154 388561
rect 359918 381325 360154 381561
rect 359918 374325 360154 374561
rect 359918 367325 360154 367561
rect 359918 360325 360154 360561
rect 359918 353325 360154 353561
rect 359918 346325 360154 346561
rect 359918 339325 360154 339561
rect 359918 332325 360154 332561
rect 359918 325325 360154 325561
rect 359918 318325 360154 318561
rect 359918 311325 360154 311561
rect 359918 304325 360154 304561
rect 359918 297325 360154 297561
rect 359918 290325 360154 290561
rect 359918 283325 360154 283561
rect 359918 276325 360154 276561
rect 359918 269325 360154 269561
rect 359918 262325 360154 262561
rect 359918 255325 360154 255561
rect 359918 248325 360154 248561
rect 359918 241325 360154 241561
rect 359918 234325 360154 234561
rect 359918 227325 360154 227561
rect 359918 220325 360154 220561
rect 359918 213325 360154 213561
rect 359918 206325 360154 206561
rect 359918 199325 360154 199561
rect 359918 192325 360154 192561
rect 359918 185325 360154 185561
rect 359918 178325 360154 178561
rect 359918 171325 360154 171561
rect 359918 164325 360154 164561
rect 359918 157325 360154 157561
rect 359918 150325 360154 150561
rect 359918 143325 360154 143561
rect 359918 136325 360154 136561
rect 359918 129325 360154 129561
rect 359918 122325 360154 122561
rect 359918 115325 360154 115561
rect 359918 108325 360154 108561
rect 359918 101325 360154 101561
rect 359918 94325 360154 94561
rect 359918 87325 360154 87561
rect 359918 80325 360154 80561
rect 359918 73325 360154 73561
rect 359918 66325 360154 66561
rect 359918 59325 360154 59561
rect 359918 52325 360154 52561
rect 359918 45325 360154 45561
rect 359918 38325 360154 38561
rect 359918 31325 360154 31561
rect 359918 24325 360154 24561
rect 359918 17325 360154 17561
rect 359918 10325 360154 10561
rect 359918 3325 360154 3561
rect 359918 -1942 360154 -1706
rect 359918 -2262 360154 -2026
rect 365186 705002 365422 705238
rect 365186 704682 365422 704918
rect 365186 695258 365422 695494
rect 365186 688258 365422 688494
rect 365186 681258 365422 681494
rect 365186 674258 365422 674494
rect 365186 667258 365422 667494
rect 365186 660258 365422 660494
rect 365186 653258 365422 653494
rect 365186 646258 365422 646494
rect 365186 639258 365422 639494
rect 365186 632258 365422 632494
rect 365186 625258 365422 625494
rect 365186 618258 365422 618494
rect 365186 611258 365422 611494
rect 365186 604258 365422 604494
rect 365186 597258 365422 597494
rect 365186 590258 365422 590494
rect 365186 583258 365422 583494
rect 365186 576258 365422 576494
rect 365186 569258 365422 569494
rect 365186 562258 365422 562494
rect 365186 555258 365422 555494
rect 365186 548258 365422 548494
rect 365186 541258 365422 541494
rect 365186 534258 365422 534494
rect 365186 527258 365422 527494
rect 365186 520258 365422 520494
rect 365186 513258 365422 513494
rect 365186 506258 365422 506494
rect 365186 499258 365422 499494
rect 365186 492258 365422 492494
rect 365186 485258 365422 485494
rect 365186 478258 365422 478494
rect 365186 471258 365422 471494
rect 365186 464258 365422 464494
rect 365186 457258 365422 457494
rect 365186 450258 365422 450494
rect 365186 443258 365422 443494
rect 365186 436258 365422 436494
rect 365186 429258 365422 429494
rect 365186 422258 365422 422494
rect 365186 415258 365422 415494
rect 365186 408258 365422 408494
rect 365186 401258 365422 401494
rect 365186 394258 365422 394494
rect 365186 387258 365422 387494
rect 365186 380258 365422 380494
rect 365186 373258 365422 373494
rect 365186 366258 365422 366494
rect 365186 359258 365422 359494
rect 365186 352258 365422 352494
rect 365186 345258 365422 345494
rect 365186 338258 365422 338494
rect 365186 331258 365422 331494
rect 365186 324258 365422 324494
rect 365186 317258 365422 317494
rect 365186 310258 365422 310494
rect 365186 303258 365422 303494
rect 365186 296258 365422 296494
rect 365186 289258 365422 289494
rect 365186 282258 365422 282494
rect 365186 275258 365422 275494
rect 365186 268258 365422 268494
rect 365186 261258 365422 261494
rect 365186 254258 365422 254494
rect 365186 247258 365422 247494
rect 365186 240258 365422 240494
rect 365186 233258 365422 233494
rect 365186 226258 365422 226494
rect 365186 219258 365422 219494
rect 365186 212258 365422 212494
rect 365186 205258 365422 205494
rect 365186 198258 365422 198494
rect 365186 191258 365422 191494
rect 365186 184258 365422 184494
rect 365186 177258 365422 177494
rect 365186 170258 365422 170494
rect 365186 163258 365422 163494
rect 365186 156258 365422 156494
rect 365186 149258 365422 149494
rect 365186 142258 365422 142494
rect 365186 135258 365422 135494
rect 365186 128258 365422 128494
rect 365186 121258 365422 121494
rect 365186 114258 365422 114494
rect 365186 107258 365422 107494
rect 365186 100258 365422 100494
rect 365186 93258 365422 93494
rect 365186 86258 365422 86494
rect 365186 79258 365422 79494
rect 365186 72258 365422 72494
rect 365186 65258 365422 65494
rect 365186 58258 365422 58494
rect 365186 51258 365422 51494
rect 365186 44258 365422 44494
rect 365186 37258 365422 37494
rect 365186 30258 365422 30494
rect 365186 23258 365422 23494
rect 365186 16258 365422 16494
rect 365186 9258 365422 9494
rect 365186 2258 365422 2494
rect 365186 -982 365422 -746
rect 365186 -1302 365422 -1066
rect 366918 705962 367154 706198
rect 366918 705642 367154 705878
rect 366918 696325 367154 696561
rect 366918 689325 367154 689561
rect 366918 682325 367154 682561
rect 366918 675325 367154 675561
rect 366918 668325 367154 668561
rect 366918 661325 367154 661561
rect 366918 654325 367154 654561
rect 366918 647325 367154 647561
rect 366918 640325 367154 640561
rect 366918 633325 367154 633561
rect 366918 626325 367154 626561
rect 366918 619325 367154 619561
rect 366918 612325 367154 612561
rect 366918 605325 367154 605561
rect 366918 598325 367154 598561
rect 366918 591325 367154 591561
rect 366918 584325 367154 584561
rect 366918 577325 367154 577561
rect 366918 570325 367154 570561
rect 366918 563325 367154 563561
rect 366918 556325 367154 556561
rect 366918 549325 367154 549561
rect 366918 542325 367154 542561
rect 366918 535325 367154 535561
rect 366918 528325 367154 528561
rect 366918 521325 367154 521561
rect 366918 514325 367154 514561
rect 366918 507325 367154 507561
rect 366918 500325 367154 500561
rect 366918 493325 367154 493561
rect 366918 486325 367154 486561
rect 366918 479325 367154 479561
rect 366918 472325 367154 472561
rect 366918 465325 367154 465561
rect 366918 458325 367154 458561
rect 366918 451325 367154 451561
rect 366918 444325 367154 444561
rect 366918 437325 367154 437561
rect 366918 430325 367154 430561
rect 366918 423325 367154 423561
rect 366918 416325 367154 416561
rect 366918 409325 367154 409561
rect 366918 402325 367154 402561
rect 366918 395325 367154 395561
rect 366918 388325 367154 388561
rect 366918 381325 367154 381561
rect 366918 374325 367154 374561
rect 366918 367325 367154 367561
rect 366918 360325 367154 360561
rect 366918 353325 367154 353561
rect 366918 346325 367154 346561
rect 366918 339325 367154 339561
rect 366918 332325 367154 332561
rect 366918 325325 367154 325561
rect 366918 318325 367154 318561
rect 366918 311325 367154 311561
rect 366918 304325 367154 304561
rect 366918 297325 367154 297561
rect 366918 290325 367154 290561
rect 366918 283325 367154 283561
rect 366918 276325 367154 276561
rect 366918 269325 367154 269561
rect 366918 262325 367154 262561
rect 366918 255325 367154 255561
rect 366918 248325 367154 248561
rect 366918 241325 367154 241561
rect 366918 234325 367154 234561
rect 366918 227325 367154 227561
rect 366918 220325 367154 220561
rect 366918 213325 367154 213561
rect 366918 206325 367154 206561
rect 366918 199325 367154 199561
rect 366918 192325 367154 192561
rect 366918 185325 367154 185561
rect 366918 178325 367154 178561
rect 366918 171325 367154 171561
rect 366918 164325 367154 164561
rect 366918 157325 367154 157561
rect 366918 150325 367154 150561
rect 366918 143325 367154 143561
rect 366918 136325 367154 136561
rect 366918 129325 367154 129561
rect 366918 122325 367154 122561
rect 366918 115325 367154 115561
rect 366918 108325 367154 108561
rect 366918 101325 367154 101561
rect 366918 94325 367154 94561
rect 366918 87325 367154 87561
rect 366918 80325 367154 80561
rect 366918 73325 367154 73561
rect 366918 66325 367154 66561
rect 366918 59325 367154 59561
rect 366918 52325 367154 52561
rect 366918 45325 367154 45561
rect 366918 38325 367154 38561
rect 366918 31325 367154 31561
rect 366918 24325 367154 24561
rect 366918 17325 367154 17561
rect 366918 10325 367154 10561
rect 366918 3325 367154 3561
rect 366918 -1942 367154 -1706
rect 366918 -2262 367154 -2026
rect 372186 705002 372422 705238
rect 372186 704682 372422 704918
rect 372186 695258 372422 695494
rect 372186 688258 372422 688494
rect 372186 681258 372422 681494
rect 372186 674258 372422 674494
rect 372186 667258 372422 667494
rect 372186 660258 372422 660494
rect 372186 653258 372422 653494
rect 372186 646258 372422 646494
rect 372186 639258 372422 639494
rect 372186 632258 372422 632494
rect 372186 625258 372422 625494
rect 372186 618258 372422 618494
rect 372186 611258 372422 611494
rect 372186 604258 372422 604494
rect 372186 597258 372422 597494
rect 372186 590258 372422 590494
rect 372186 583258 372422 583494
rect 372186 576258 372422 576494
rect 372186 569258 372422 569494
rect 372186 562258 372422 562494
rect 372186 555258 372422 555494
rect 372186 548258 372422 548494
rect 372186 541258 372422 541494
rect 372186 534258 372422 534494
rect 372186 527258 372422 527494
rect 372186 520258 372422 520494
rect 372186 513258 372422 513494
rect 372186 506258 372422 506494
rect 372186 499258 372422 499494
rect 372186 492258 372422 492494
rect 372186 485258 372422 485494
rect 372186 478258 372422 478494
rect 372186 471258 372422 471494
rect 372186 464258 372422 464494
rect 372186 457258 372422 457494
rect 372186 450258 372422 450494
rect 372186 443258 372422 443494
rect 372186 436258 372422 436494
rect 372186 429258 372422 429494
rect 372186 422258 372422 422494
rect 372186 415258 372422 415494
rect 372186 408258 372422 408494
rect 372186 401258 372422 401494
rect 372186 394258 372422 394494
rect 372186 387258 372422 387494
rect 372186 380258 372422 380494
rect 372186 373258 372422 373494
rect 372186 366258 372422 366494
rect 372186 359258 372422 359494
rect 372186 352258 372422 352494
rect 372186 345258 372422 345494
rect 372186 338258 372422 338494
rect 372186 331258 372422 331494
rect 372186 324258 372422 324494
rect 372186 317258 372422 317494
rect 372186 310258 372422 310494
rect 372186 303258 372422 303494
rect 372186 296258 372422 296494
rect 372186 289258 372422 289494
rect 372186 282258 372422 282494
rect 372186 275258 372422 275494
rect 372186 268258 372422 268494
rect 372186 261258 372422 261494
rect 372186 254258 372422 254494
rect 372186 247258 372422 247494
rect 372186 240258 372422 240494
rect 372186 233258 372422 233494
rect 372186 226258 372422 226494
rect 372186 219258 372422 219494
rect 372186 212258 372422 212494
rect 372186 205258 372422 205494
rect 372186 198258 372422 198494
rect 372186 191258 372422 191494
rect 372186 184258 372422 184494
rect 372186 177258 372422 177494
rect 372186 170258 372422 170494
rect 372186 163258 372422 163494
rect 372186 156258 372422 156494
rect 372186 149258 372422 149494
rect 372186 142258 372422 142494
rect 372186 135258 372422 135494
rect 372186 128258 372422 128494
rect 372186 121258 372422 121494
rect 372186 114258 372422 114494
rect 372186 107258 372422 107494
rect 372186 100258 372422 100494
rect 372186 93258 372422 93494
rect 372186 86258 372422 86494
rect 372186 79258 372422 79494
rect 372186 72258 372422 72494
rect 372186 65258 372422 65494
rect 372186 58258 372422 58494
rect 372186 51258 372422 51494
rect 372186 44258 372422 44494
rect 372186 37258 372422 37494
rect 372186 30258 372422 30494
rect 372186 23258 372422 23494
rect 372186 16258 372422 16494
rect 372186 9258 372422 9494
rect 372186 2258 372422 2494
rect 372186 -982 372422 -746
rect 372186 -1302 372422 -1066
rect 373918 705962 374154 706198
rect 373918 705642 374154 705878
rect 373918 696325 374154 696561
rect 373918 689325 374154 689561
rect 373918 682325 374154 682561
rect 373918 675325 374154 675561
rect 373918 668325 374154 668561
rect 373918 661325 374154 661561
rect 373918 654325 374154 654561
rect 373918 647325 374154 647561
rect 373918 640325 374154 640561
rect 373918 633325 374154 633561
rect 373918 626325 374154 626561
rect 373918 619325 374154 619561
rect 373918 612325 374154 612561
rect 373918 605325 374154 605561
rect 373918 598325 374154 598561
rect 373918 591325 374154 591561
rect 373918 584325 374154 584561
rect 373918 577325 374154 577561
rect 373918 570325 374154 570561
rect 373918 563325 374154 563561
rect 373918 556325 374154 556561
rect 373918 549325 374154 549561
rect 373918 542325 374154 542561
rect 373918 535325 374154 535561
rect 373918 528325 374154 528561
rect 373918 521325 374154 521561
rect 373918 514325 374154 514561
rect 373918 507325 374154 507561
rect 373918 500325 374154 500561
rect 373918 493325 374154 493561
rect 373918 486325 374154 486561
rect 373918 479325 374154 479561
rect 373918 472325 374154 472561
rect 373918 465325 374154 465561
rect 373918 458325 374154 458561
rect 373918 451325 374154 451561
rect 373918 444325 374154 444561
rect 373918 437325 374154 437561
rect 373918 430325 374154 430561
rect 373918 423325 374154 423561
rect 373918 416325 374154 416561
rect 373918 409325 374154 409561
rect 373918 402325 374154 402561
rect 373918 395325 374154 395561
rect 373918 388325 374154 388561
rect 373918 381325 374154 381561
rect 373918 374325 374154 374561
rect 373918 367325 374154 367561
rect 373918 360325 374154 360561
rect 373918 353325 374154 353561
rect 373918 346325 374154 346561
rect 373918 339325 374154 339561
rect 373918 332325 374154 332561
rect 373918 325325 374154 325561
rect 373918 318325 374154 318561
rect 373918 311325 374154 311561
rect 373918 304325 374154 304561
rect 373918 297325 374154 297561
rect 373918 290325 374154 290561
rect 373918 283325 374154 283561
rect 373918 276325 374154 276561
rect 373918 269325 374154 269561
rect 373918 262325 374154 262561
rect 373918 255325 374154 255561
rect 373918 248325 374154 248561
rect 373918 241325 374154 241561
rect 373918 234325 374154 234561
rect 373918 227325 374154 227561
rect 373918 220325 374154 220561
rect 373918 213325 374154 213561
rect 373918 206325 374154 206561
rect 373918 199325 374154 199561
rect 373918 192325 374154 192561
rect 373918 185325 374154 185561
rect 373918 178325 374154 178561
rect 373918 171325 374154 171561
rect 373918 164325 374154 164561
rect 373918 157325 374154 157561
rect 373918 150325 374154 150561
rect 373918 143325 374154 143561
rect 373918 136325 374154 136561
rect 373918 129325 374154 129561
rect 373918 122325 374154 122561
rect 373918 115325 374154 115561
rect 373918 108325 374154 108561
rect 373918 101325 374154 101561
rect 373918 94325 374154 94561
rect 373918 87325 374154 87561
rect 373918 80325 374154 80561
rect 373918 73325 374154 73561
rect 373918 66325 374154 66561
rect 373918 59325 374154 59561
rect 373918 52325 374154 52561
rect 373918 45325 374154 45561
rect 373918 38325 374154 38561
rect 373918 31325 374154 31561
rect 373918 24325 374154 24561
rect 373918 17325 374154 17561
rect 373918 10325 374154 10561
rect 373918 3325 374154 3561
rect 373918 -1942 374154 -1706
rect 373918 -2262 374154 -2026
rect 379186 705002 379422 705238
rect 379186 704682 379422 704918
rect 379186 695258 379422 695494
rect 379186 688258 379422 688494
rect 379186 681258 379422 681494
rect 379186 674258 379422 674494
rect 379186 667258 379422 667494
rect 379186 660258 379422 660494
rect 379186 653258 379422 653494
rect 379186 646258 379422 646494
rect 379186 639258 379422 639494
rect 379186 632258 379422 632494
rect 379186 625258 379422 625494
rect 379186 618258 379422 618494
rect 379186 611258 379422 611494
rect 379186 604258 379422 604494
rect 379186 597258 379422 597494
rect 379186 590258 379422 590494
rect 379186 583258 379422 583494
rect 379186 576258 379422 576494
rect 379186 569258 379422 569494
rect 379186 562258 379422 562494
rect 379186 555258 379422 555494
rect 379186 548258 379422 548494
rect 379186 541258 379422 541494
rect 379186 534258 379422 534494
rect 379186 527258 379422 527494
rect 379186 520258 379422 520494
rect 379186 513258 379422 513494
rect 379186 506258 379422 506494
rect 379186 499258 379422 499494
rect 379186 492258 379422 492494
rect 379186 485258 379422 485494
rect 379186 478258 379422 478494
rect 379186 471258 379422 471494
rect 379186 464258 379422 464494
rect 379186 457258 379422 457494
rect 379186 450258 379422 450494
rect 379186 443258 379422 443494
rect 379186 436258 379422 436494
rect 379186 429258 379422 429494
rect 379186 422258 379422 422494
rect 379186 415258 379422 415494
rect 379186 408258 379422 408494
rect 379186 401258 379422 401494
rect 379186 394258 379422 394494
rect 379186 387258 379422 387494
rect 379186 380258 379422 380494
rect 379186 373258 379422 373494
rect 379186 366258 379422 366494
rect 379186 359258 379422 359494
rect 379186 352258 379422 352494
rect 379186 345258 379422 345494
rect 379186 338258 379422 338494
rect 379186 331258 379422 331494
rect 379186 324258 379422 324494
rect 379186 317258 379422 317494
rect 379186 310258 379422 310494
rect 379186 303258 379422 303494
rect 379186 296258 379422 296494
rect 379186 289258 379422 289494
rect 379186 282258 379422 282494
rect 379186 275258 379422 275494
rect 379186 268258 379422 268494
rect 379186 261258 379422 261494
rect 379186 254258 379422 254494
rect 379186 247258 379422 247494
rect 379186 240258 379422 240494
rect 379186 233258 379422 233494
rect 379186 226258 379422 226494
rect 379186 219258 379422 219494
rect 379186 212258 379422 212494
rect 379186 205258 379422 205494
rect 379186 198258 379422 198494
rect 379186 191258 379422 191494
rect 379186 184258 379422 184494
rect 379186 177258 379422 177494
rect 379186 170258 379422 170494
rect 379186 163258 379422 163494
rect 379186 156258 379422 156494
rect 379186 149258 379422 149494
rect 379186 142258 379422 142494
rect 379186 135258 379422 135494
rect 379186 128258 379422 128494
rect 379186 121258 379422 121494
rect 379186 114258 379422 114494
rect 379186 107258 379422 107494
rect 379186 100258 379422 100494
rect 379186 93258 379422 93494
rect 379186 86258 379422 86494
rect 379186 79258 379422 79494
rect 379186 72258 379422 72494
rect 379186 65258 379422 65494
rect 379186 58258 379422 58494
rect 379186 51258 379422 51494
rect 379186 44258 379422 44494
rect 379186 37258 379422 37494
rect 379186 30258 379422 30494
rect 379186 23258 379422 23494
rect 379186 16258 379422 16494
rect 379186 9258 379422 9494
rect 379186 2258 379422 2494
rect 379186 -982 379422 -746
rect 379186 -1302 379422 -1066
rect 380918 705962 381154 706198
rect 380918 705642 381154 705878
rect 380918 696325 381154 696561
rect 380918 689325 381154 689561
rect 380918 682325 381154 682561
rect 380918 675325 381154 675561
rect 380918 668325 381154 668561
rect 380918 661325 381154 661561
rect 380918 654325 381154 654561
rect 380918 647325 381154 647561
rect 380918 640325 381154 640561
rect 380918 633325 381154 633561
rect 380918 626325 381154 626561
rect 380918 619325 381154 619561
rect 380918 612325 381154 612561
rect 380918 605325 381154 605561
rect 380918 598325 381154 598561
rect 380918 591325 381154 591561
rect 380918 584325 381154 584561
rect 380918 577325 381154 577561
rect 380918 570325 381154 570561
rect 380918 563325 381154 563561
rect 380918 556325 381154 556561
rect 380918 549325 381154 549561
rect 380918 542325 381154 542561
rect 380918 535325 381154 535561
rect 380918 528325 381154 528561
rect 380918 521325 381154 521561
rect 380918 514325 381154 514561
rect 380918 507325 381154 507561
rect 380918 500325 381154 500561
rect 380918 493325 381154 493561
rect 380918 486325 381154 486561
rect 380918 479325 381154 479561
rect 380918 472325 381154 472561
rect 380918 465325 381154 465561
rect 380918 458325 381154 458561
rect 380918 451325 381154 451561
rect 380918 444325 381154 444561
rect 380918 437325 381154 437561
rect 380918 430325 381154 430561
rect 380918 423325 381154 423561
rect 380918 416325 381154 416561
rect 380918 409325 381154 409561
rect 380918 402325 381154 402561
rect 380918 395325 381154 395561
rect 380918 388325 381154 388561
rect 380918 381325 381154 381561
rect 380918 374325 381154 374561
rect 380918 367325 381154 367561
rect 380918 360325 381154 360561
rect 380918 353325 381154 353561
rect 380918 346325 381154 346561
rect 380918 339325 381154 339561
rect 380918 332325 381154 332561
rect 380918 325325 381154 325561
rect 380918 318325 381154 318561
rect 380918 311325 381154 311561
rect 380918 304325 381154 304561
rect 380918 297325 381154 297561
rect 380918 290325 381154 290561
rect 380918 283325 381154 283561
rect 380918 276325 381154 276561
rect 380918 269325 381154 269561
rect 380918 262325 381154 262561
rect 380918 255325 381154 255561
rect 380918 248325 381154 248561
rect 380918 241325 381154 241561
rect 380918 234325 381154 234561
rect 380918 227325 381154 227561
rect 380918 220325 381154 220561
rect 380918 213325 381154 213561
rect 380918 206325 381154 206561
rect 380918 199325 381154 199561
rect 380918 192325 381154 192561
rect 380918 185325 381154 185561
rect 380918 178325 381154 178561
rect 380918 171325 381154 171561
rect 380918 164325 381154 164561
rect 380918 157325 381154 157561
rect 380918 150325 381154 150561
rect 380918 143325 381154 143561
rect 380918 136325 381154 136561
rect 380918 129325 381154 129561
rect 380918 122325 381154 122561
rect 380918 115325 381154 115561
rect 380918 108325 381154 108561
rect 380918 101325 381154 101561
rect 380918 94325 381154 94561
rect 380918 87325 381154 87561
rect 380918 80325 381154 80561
rect 380918 73325 381154 73561
rect 380918 66325 381154 66561
rect 380918 59325 381154 59561
rect 380918 52325 381154 52561
rect 380918 45325 381154 45561
rect 380918 38325 381154 38561
rect 380918 31325 381154 31561
rect 380918 24325 381154 24561
rect 380918 17325 381154 17561
rect 380918 10325 381154 10561
rect 380918 3325 381154 3561
rect 380918 -1942 381154 -1706
rect 380918 -2262 381154 -2026
rect 386186 705002 386422 705238
rect 386186 704682 386422 704918
rect 386186 695258 386422 695494
rect 386186 688258 386422 688494
rect 386186 681258 386422 681494
rect 386186 674258 386422 674494
rect 386186 667258 386422 667494
rect 386186 660258 386422 660494
rect 386186 653258 386422 653494
rect 386186 646258 386422 646494
rect 386186 639258 386422 639494
rect 386186 632258 386422 632494
rect 386186 625258 386422 625494
rect 386186 618258 386422 618494
rect 386186 611258 386422 611494
rect 386186 604258 386422 604494
rect 386186 597258 386422 597494
rect 386186 590258 386422 590494
rect 386186 583258 386422 583494
rect 386186 576258 386422 576494
rect 386186 569258 386422 569494
rect 386186 562258 386422 562494
rect 386186 555258 386422 555494
rect 386186 548258 386422 548494
rect 386186 541258 386422 541494
rect 386186 534258 386422 534494
rect 386186 527258 386422 527494
rect 386186 520258 386422 520494
rect 386186 513258 386422 513494
rect 386186 506258 386422 506494
rect 386186 499258 386422 499494
rect 386186 492258 386422 492494
rect 386186 485258 386422 485494
rect 386186 478258 386422 478494
rect 386186 471258 386422 471494
rect 386186 464258 386422 464494
rect 386186 457258 386422 457494
rect 386186 450258 386422 450494
rect 386186 443258 386422 443494
rect 386186 436258 386422 436494
rect 386186 429258 386422 429494
rect 386186 422258 386422 422494
rect 386186 415258 386422 415494
rect 386186 408258 386422 408494
rect 386186 401258 386422 401494
rect 386186 394258 386422 394494
rect 386186 387258 386422 387494
rect 386186 380258 386422 380494
rect 386186 373258 386422 373494
rect 386186 366258 386422 366494
rect 386186 359258 386422 359494
rect 386186 352258 386422 352494
rect 386186 345258 386422 345494
rect 386186 338258 386422 338494
rect 386186 331258 386422 331494
rect 386186 324258 386422 324494
rect 386186 317258 386422 317494
rect 386186 310258 386422 310494
rect 386186 303258 386422 303494
rect 386186 296258 386422 296494
rect 386186 289258 386422 289494
rect 386186 282258 386422 282494
rect 386186 275258 386422 275494
rect 386186 268258 386422 268494
rect 386186 261258 386422 261494
rect 386186 254258 386422 254494
rect 386186 247258 386422 247494
rect 386186 240258 386422 240494
rect 386186 233258 386422 233494
rect 386186 226258 386422 226494
rect 386186 219258 386422 219494
rect 386186 212258 386422 212494
rect 386186 205258 386422 205494
rect 386186 198258 386422 198494
rect 386186 191258 386422 191494
rect 386186 184258 386422 184494
rect 386186 177258 386422 177494
rect 386186 170258 386422 170494
rect 386186 163258 386422 163494
rect 386186 156258 386422 156494
rect 386186 149258 386422 149494
rect 386186 142258 386422 142494
rect 386186 135258 386422 135494
rect 386186 128258 386422 128494
rect 386186 121258 386422 121494
rect 386186 114258 386422 114494
rect 386186 107258 386422 107494
rect 386186 100258 386422 100494
rect 386186 93258 386422 93494
rect 386186 86258 386422 86494
rect 386186 79258 386422 79494
rect 386186 72258 386422 72494
rect 386186 65258 386422 65494
rect 386186 58258 386422 58494
rect 386186 51258 386422 51494
rect 386186 44258 386422 44494
rect 386186 37258 386422 37494
rect 386186 30258 386422 30494
rect 386186 23258 386422 23494
rect 386186 16258 386422 16494
rect 386186 9258 386422 9494
rect 386186 2258 386422 2494
rect 386186 -982 386422 -746
rect 386186 -1302 386422 -1066
rect 387918 705962 388154 706198
rect 387918 705642 388154 705878
rect 387918 696325 388154 696561
rect 387918 689325 388154 689561
rect 387918 682325 388154 682561
rect 387918 675325 388154 675561
rect 387918 668325 388154 668561
rect 387918 661325 388154 661561
rect 387918 654325 388154 654561
rect 387918 647325 388154 647561
rect 387918 640325 388154 640561
rect 387918 633325 388154 633561
rect 387918 626325 388154 626561
rect 387918 619325 388154 619561
rect 387918 612325 388154 612561
rect 387918 605325 388154 605561
rect 387918 598325 388154 598561
rect 387918 591325 388154 591561
rect 387918 584325 388154 584561
rect 387918 577325 388154 577561
rect 387918 570325 388154 570561
rect 387918 563325 388154 563561
rect 387918 556325 388154 556561
rect 387918 549325 388154 549561
rect 387918 542325 388154 542561
rect 387918 535325 388154 535561
rect 387918 528325 388154 528561
rect 387918 521325 388154 521561
rect 387918 514325 388154 514561
rect 387918 507325 388154 507561
rect 387918 500325 388154 500561
rect 387918 493325 388154 493561
rect 387918 486325 388154 486561
rect 387918 479325 388154 479561
rect 387918 472325 388154 472561
rect 387918 465325 388154 465561
rect 387918 458325 388154 458561
rect 387918 451325 388154 451561
rect 387918 444325 388154 444561
rect 387918 437325 388154 437561
rect 387918 430325 388154 430561
rect 387918 423325 388154 423561
rect 387918 416325 388154 416561
rect 387918 409325 388154 409561
rect 387918 402325 388154 402561
rect 387918 395325 388154 395561
rect 387918 388325 388154 388561
rect 387918 381325 388154 381561
rect 387918 374325 388154 374561
rect 387918 367325 388154 367561
rect 387918 360325 388154 360561
rect 387918 353325 388154 353561
rect 387918 346325 388154 346561
rect 387918 339325 388154 339561
rect 387918 332325 388154 332561
rect 387918 325325 388154 325561
rect 387918 318325 388154 318561
rect 387918 311325 388154 311561
rect 387918 304325 388154 304561
rect 387918 297325 388154 297561
rect 387918 290325 388154 290561
rect 387918 283325 388154 283561
rect 387918 276325 388154 276561
rect 387918 269325 388154 269561
rect 387918 262325 388154 262561
rect 387918 255325 388154 255561
rect 387918 248325 388154 248561
rect 387918 241325 388154 241561
rect 387918 234325 388154 234561
rect 387918 227325 388154 227561
rect 387918 220325 388154 220561
rect 387918 213325 388154 213561
rect 387918 206325 388154 206561
rect 387918 199325 388154 199561
rect 387918 192325 388154 192561
rect 387918 185325 388154 185561
rect 387918 178325 388154 178561
rect 387918 171325 388154 171561
rect 387918 164325 388154 164561
rect 387918 157325 388154 157561
rect 387918 150325 388154 150561
rect 387918 143325 388154 143561
rect 387918 136325 388154 136561
rect 387918 129325 388154 129561
rect 387918 122325 388154 122561
rect 387918 115325 388154 115561
rect 387918 108325 388154 108561
rect 387918 101325 388154 101561
rect 387918 94325 388154 94561
rect 387918 87325 388154 87561
rect 387918 80325 388154 80561
rect 387918 73325 388154 73561
rect 387918 66325 388154 66561
rect 387918 59325 388154 59561
rect 387918 52325 388154 52561
rect 387918 45325 388154 45561
rect 387918 38325 388154 38561
rect 387918 31325 388154 31561
rect 387918 24325 388154 24561
rect 387918 17325 388154 17561
rect 387918 10325 388154 10561
rect 387918 3325 388154 3561
rect 387918 -1942 388154 -1706
rect 387918 -2262 388154 -2026
rect 393186 705002 393422 705238
rect 393186 704682 393422 704918
rect 393186 695258 393422 695494
rect 393186 688258 393422 688494
rect 393186 681258 393422 681494
rect 393186 674258 393422 674494
rect 393186 667258 393422 667494
rect 393186 660258 393422 660494
rect 393186 653258 393422 653494
rect 393186 646258 393422 646494
rect 393186 639258 393422 639494
rect 393186 632258 393422 632494
rect 393186 625258 393422 625494
rect 393186 618258 393422 618494
rect 393186 611258 393422 611494
rect 393186 604258 393422 604494
rect 393186 597258 393422 597494
rect 393186 590258 393422 590494
rect 393186 583258 393422 583494
rect 393186 576258 393422 576494
rect 393186 569258 393422 569494
rect 393186 562258 393422 562494
rect 393186 555258 393422 555494
rect 393186 548258 393422 548494
rect 393186 541258 393422 541494
rect 393186 534258 393422 534494
rect 393186 527258 393422 527494
rect 393186 520258 393422 520494
rect 393186 513258 393422 513494
rect 393186 506258 393422 506494
rect 393186 499258 393422 499494
rect 393186 492258 393422 492494
rect 393186 485258 393422 485494
rect 393186 478258 393422 478494
rect 393186 471258 393422 471494
rect 393186 464258 393422 464494
rect 393186 457258 393422 457494
rect 393186 450258 393422 450494
rect 393186 443258 393422 443494
rect 393186 436258 393422 436494
rect 393186 429258 393422 429494
rect 393186 422258 393422 422494
rect 393186 415258 393422 415494
rect 393186 408258 393422 408494
rect 393186 401258 393422 401494
rect 393186 394258 393422 394494
rect 393186 387258 393422 387494
rect 393186 380258 393422 380494
rect 393186 373258 393422 373494
rect 393186 366258 393422 366494
rect 393186 359258 393422 359494
rect 393186 352258 393422 352494
rect 393186 345258 393422 345494
rect 393186 338258 393422 338494
rect 393186 331258 393422 331494
rect 393186 324258 393422 324494
rect 393186 317258 393422 317494
rect 393186 310258 393422 310494
rect 393186 303258 393422 303494
rect 393186 296258 393422 296494
rect 393186 289258 393422 289494
rect 393186 282258 393422 282494
rect 393186 275258 393422 275494
rect 393186 268258 393422 268494
rect 393186 261258 393422 261494
rect 393186 254258 393422 254494
rect 393186 247258 393422 247494
rect 393186 240258 393422 240494
rect 393186 233258 393422 233494
rect 393186 226258 393422 226494
rect 393186 219258 393422 219494
rect 393186 212258 393422 212494
rect 393186 205258 393422 205494
rect 393186 198258 393422 198494
rect 393186 191258 393422 191494
rect 393186 184258 393422 184494
rect 393186 177258 393422 177494
rect 393186 170258 393422 170494
rect 393186 163258 393422 163494
rect 393186 156258 393422 156494
rect 393186 149258 393422 149494
rect 393186 142258 393422 142494
rect 393186 135258 393422 135494
rect 393186 128258 393422 128494
rect 393186 121258 393422 121494
rect 393186 114258 393422 114494
rect 393186 107258 393422 107494
rect 393186 100258 393422 100494
rect 393186 93258 393422 93494
rect 393186 86258 393422 86494
rect 393186 79258 393422 79494
rect 393186 72258 393422 72494
rect 393186 65258 393422 65494
rect 393186 58258 393422 58494
rect 393186 51258 393422 51494
rect 393186 44258 393422 44494
rect 393186 37258 393422 37494
rect 393186 30258 393422 30494
rect 393186 23258 393422 23494
rect 393186 16258 393422 16494
rect 393186 9258 393422 9494
rect 393186 2258 393422 2494
rect 393186 -982 393422 -746
rect 393186 -1302 393422 -1066
rect 394918 705962 395154 706198
rect 394918 705642 395154 705878
rect 394918 696325 395154 696561
rect 394918 689325 395154 689561
rect 394918 682325 395154 682561
rect 394918 675325 395154 675561
rect 394918 668325 395154 668561
rect 394918 661325 395154 661561
rect 394918 654325 395154 654561
rect 394918 647325 395154 647561
rect 394918 640325 395154 640561
rect 394918 633325 395154 633561
rect 394918 626325 395154 626561
rect 394918 619325 395154 619561
rect 394918 612325 395154 612561
rect 394918 605325 395154 605561
rect 394918 598325 395154 598561
rect 394918 591325 395154 591561
rect 394918 584325 395154 584561
rect 394918 577325 395154 577561
rect 394918 570325 395154 570561
rect 394918 563325 395154 563561
rect 394918 556325 395154 556561
rect 394918 549325 395154 549561
rect 394918 542325 395154 542561
rect 394918 535325 395154 535561
rect 394918 528325 395154 528561
rect 394918 521325 395154 521561
rect 394918 514325 395154 514561
rect 394918 507325 395154 507561
rect 394918 500325 395154 500561
rect 394918 493325 395154 493561
rect 394918 486325 395154 486561
rect 394918 479325 395154 479561
rect 394918 472325 395154 472561
rect 394918 465325 395154 465561
rect 394918 458325 395154 458561
rect 394918 451325 395154 451561
rect 394918 444325 395154 444561
rect 394918 437325 395154 437561
rect 394918 430325 395154 430561
rect 394918 423325 395154 423561
rect 394918 416325 395154 416561
rect 394918 409325 395154 409561
rect 394918 402325 395154 402561
rect 394918 395325 395154 395561
rect 394918 388325 395154 388561
rect 394918 381325 395154 381561
rect 394918 374325 395154 374561
rect 394918 367325 395154 367561
rect 394918 360325 395154 360561
rect 394918 353325 395154 353561
rect 394918 346325 395154 346561
rect 394918 339325 395154 339561
rect 394918 332325 395154 332561
rect 394918 325325 395154 325561
rect 394918 318325 395154 318561
rect 394918 311325 395154 311561
rect 394918 304325 395154 304561
rect 394918 297325 395154 297561
rect 394918 290325 395154 290561
rect 394918 283325 395154 283561
rect 394918 276325 395154 276561
rect 394918 269325 395154 269561
rect 394918 262325 395154 262561
rect 394918 255325 395154 255561
rect 394918 248325 395154 248561
rect 394918 241325 395154 241561
rect 394918 234325 395154 234561
rect 394918 227325 395154 227561
rect 394918 220325 395154 220561
rect 394918 213325 395154 213561
rect 394918 206325 395154 206561
rect 394918 199325 395154 199561
rect 394918 192325 395154 192561
rect 394918 185325 395154 185561
rect 394918 178325 395154 178561
rect 394918 171325 395154 171561
rect 394918 164325 395154 164561
rect 394918 157325 395154 157561
rect 394918 150325 395154 150561
rect 394918 143325 395154 143561
rect 394918 136325 395154 136561
rect 394918 129325 395154 129561
rect 394918 122325 395154 122561
rect 394918 115325 395154 115561
rect 394918 108325 395154 108561
rect 394918 101325 395154 101561
rect 394918 94325 395154 94561
rect 394918 87325 395154 87561
rect 394918 80325 395154 80561
rect 394918 73325 395154 73561
rect 394918 66325 395154 66561
rect 394918 59325 395154 59561
rect 394918 52325 395154 52561
rect 394918 45325 395154 45561
rect 394918 38325 395154 38561
rect 394918 31325 395154 31561
rect 394918 24325 395154 24561
rect 394918 17325 395154 17561
rect 394918 10325 395154 10561
rect 394918 3325 395154 3561
rect 394918 -1942 395154 -1706
rect 394918 -2262 395154 -2026
rect 400186 705002 400422 705238
rect 400186 704682 400422 704918
rect 400186 695258 400422 695494
rect 400186 688258 400422 688494
rect 400186 681258 400422 681494
rect 400186 674258 400422 674494
rect 400186 667258 400422 667494
rect 400186 660258 400422 660494
rect 400186 653258 400422 653494
rect 400186 646258 400422 646494
rect 400186 639258 400422 639494
rect 400186 632258 400422 632494
rect 400186 625258 400422 625494
rect 400186 618258 400422 618494
rect 400186 611258 400422 611494
rect 400186 604258 400422 604494
rect 400186 597258 400422 597494
rect 400186 590258 400422 590494
rect 400186 583258 400422 583494
rect 400186 576258 400422 576494
rect 400186 569258 400422 569494
rect 400186 562258 400422 562494
rect 400186 555258 400422 555494
rect 400186 548258 400422 548494
rect 400186 541258 400422 541494
rect 400186 534258 400422 534494
rect 400186 527258 400422 527494
rect 400186 520258 400422 520494
rect 400186 513258 400422 513494
rect 400186 506258 400422 506494
rect 400186 499258 400422 499494
rect 400186 492258 400422 492494
rect 400186 485258 400422 485494
rect 400186 478258 400422 478494
rect 400186 471258 400422 471494
rect 400186 464258 400422 464494
rect 400186 457258 400422 457494
rect 400186 450258 400422 450494
rect 400186 443258 400422 443494
rect 400186 436258 400422 436494
rect 400186 429258 400422 429494
rect 400186 422258 400422 422494
rect 400186 415258 400422 415494
rect 400186 408258 400422 408494
rect 400186 401258 400422 401494
rect 400186 394258 400422 394494
rect 400186 387258 400422 387494
rect 400186 380258 400422 380494
rect 400186 373258 400422 373494
rect 400186 366258 400422 366494
rect 400186 359258 400422 359494
rect 400186 352258 400422 352494
rect 400186 345258 400422 345494
rect 400186 338258 400422 338494
rect 400186 331258 400422 331494
rect 400186 324258 400422 324494
rect 400186 317258 400422 317494
rect 400186 310258 400422 310494
rect 400186 303258 400422 303494
rect 400186 296258 400422 296494
rect 400186 289258 400422 289494
rect 400186 282258 400422 282494
rect 400186 275258 400422 275494
rect 400186 268258 400422 268494
rect 400186 261258 400422 261494
rect 400186 254258 400422 254494
rect 400186 247258 400422 247494
rect 400186 240258 400422 240494
rect 400186 233258 400422 233494
rect 400186 226258 400422 226494
rect 400186 219258 400422 219494
rect 400186 212258 400422 212494
rect 400186 205258 400422 205494
rect 400186 198258 400422 198494
rect 400186 191258 400422 191494
rect 400186 184258 400422 184494
rect 400186 177258 400422 177494
rect 400186 170258 400422 170494
rect 400186 163258 400422 163494
rect 400186 156258 400422 156494
rect 400186 149258 400422 149494
rect 400186 142258 400422 142494
rect 400186 135258 400422 135494
rect 400186 128258 400422 128494
rect 400186 121258 400422 121494
rect 400186 114258 400422 114494
rect 400186 107258 400422 107494
rect 400186 100258 400422 100494
rect 400186 93258 400422 93494
rect 400186 86258 400422 86494
rect 400186 79258 400422 79494
rect 400186 72258 400422 72494
rect 400186 65258 400422 65494
rect 400186 58258 400422 58494
rect 400186 51258 400422 51494
rect 400186 44258 400422 44494
rect 400186 37258 400422 37494
rect 400186 30258 400422 30494
rect 400186 23258 400422 23494
rect 400186 16258 400422 16494
rect 400186 9258 400422 9494
rect 400186 2258 400422 2494
rect 400186 -982 400422 -746
rect 400186 -1302 400422 -1066
rect 401918 705962 402154 706198
rect 401918 705642 402154 705878
rect 401918 696325 402154 696561
rect 401918 689325 402154 689561
rect 401918 682325 402154 682561
rect 401918 675325 402154 675561
rect 401918 668325 402154 668561
rect 401918 661325 402154 661561
rect 401918 654325 402154 654561
rect 401918 647325 402154 647561
rect 401918 640325 402154 640561
rect 401918 633325 402154 633561
rect 401918 626325 402154 626561
rect 401918 619325 402154 619561
rect 401918 612325 402154 612561
rect 401918 605325 402154 605561
rect 401918 598325 402154 598561
rect 401918 591325 402154 591561
rect 401918 584325 402154 584561
rect 401918 577325 402154 577561
rect 401918 570325 402154 570561
rect 401918 563325 402154 563561
rect 401918 556325 402154 556561
rect 401918 549325 402154 549561
rect 401918 542325 402154 542561
rect 401918 535325 402154 535561
rect 401918 528325 402154 528561
rect 401918 521325 402154 521561
rect 401918 514325 402154 514561
rect 401918 507325 402154 507561
rect 401918 500325 402154 500561
rect 401918 493325 402154 493561
rect 401918 486325 402154 486561
rect 401918 479325 402154 479561
rect 401918 472325 402154 472561
rect 401918 465325 402154 465561
rect 401918 458325 402154 458561
rect 401918 451325 402154 451561
rect 401918 444325 402154 444561
rect 401918 437325 402154 437561
rect 401918 430325 402154 430561
rect 401918 423325 402154 423561
rect 401918 416325 402154 416561
rect 401918 409325 402154 409561
rect 401918 402325 402154 402561
rect 401918 395325 402154 395561
rect 401918 388325 402154 388561
rect 401918 381325 402154 381561
rect 401918 374325 402154 374561
rect 401918 367325 402154 367561
rect 401918 360325 402154 360561
rect 401918 353325 402154 353561
rect 401918 346325 402154 346561
rect 401918 339325 402154 339561
rect 401918 332325 402154 332561
rect 401918 325325 402154 325561
rect 401918 318325 402154 318561
rect 401918 311325 402154 311561
rect 401918 304325 402154 304561
rect 401918 297325 402154 297561
rect 401918 290325 402154 290561
rect 401918 283325 402154 283561
rect 401918 276325 402154 276561
rect 401918 269325 402154 269561
rect 401918 262325 402154 262561
rect 401918 255325 402154 255561
rect 401918 248325 402154 248561
rect 401918 241325 402154 241561
rect 401918 234325 402154 234561
rect 401918 227325 402154 227561
rect 401918 220325 402154 220561
rect 401918 213325 402154 213561
rect 401918 206325 402154 206561
rect 401918 199325 402154 199561
rect 401918 192325 402154 192561
rect 401918 185325 402154 185561
rect 401918 178325 402154 178561
rect 401918 171325 402154 171561
rect 401918 164325 402154 164561
rect 401918 157325 402154 157561
rect 401918 150325 402154 150561
rect 401918 143325 402154 143561
rect 401918 136325 402154 136561
rect 401918 129325 402154 129561
rect 401918 122325 402154 122561
rect 401918 115325 402154 115561
rect 401918 108325 402154 108561
rect 401918 101325 402154 101561
rect 401918 94325 402154 94561
rect 401918 87325 402154 87561
rect 401918 80325 402154 80561
rect 401918 73325 402154 73561
rect 401918 66325 402154 66561
rect 401918 59325 402154 59561
rect 401918 52325 402154 52561
rect 401918 45325 402154 45561
rect 401918 38325 402154 38561
rect 401918 31325 402154 31561
rect 401918 24325 402154 24561
rect 401918 17325 402154 17561
rect 401918 10325 402154 10561
rect 401918 3325 402154 3561
rect 401918 -1942 402154 -1706
rect 401918 -2262 402154 -2026
rect 407186 705002 407422 705238
rect 407186 704682 407422 704918
rect 407186 695258 407422 695494
rect 407186 688258 407422 688494
rect 407186 681258 407422 681494
rect 407186 674258 407422 674494
rect 407186 667258 407422 667494
rect 407186 660258 407422 660494
rect 407186 653258 407422 653494
rect 407186 646258 407422 646494
rect 407186 639258 407422 639494
rect 407186 632258 407422 632494
rect 407186 625258 407422 625494
rect 407186 618258 407422 618494
rect 407186 611258 407422 611494
rect 407186 604258 407422 604494
rect 407186 597258 407422 597494
rect 407186 590258 407422 590494
rect 407186 583258 407422 583494
rect 407186 576258 407422 576494
rect 407186 569258 407422 569494
rect 407186 562258 407422 562494
rect 407186 555258 407422 555494
rect 407186 548258 407422 548494
rect 407186 541258 407422 541494
rect 407186 534258 407422 534494
rect 407186 527258 407422 527494
rect 407186 520258 407422 520494
rect 407186 513258 407422 513494
rect 407186 506258 407422 506494
rect 407186 499258 407422 499494
rect 407186 492258 407422 492494
rect 407186 485258 407422 485494
rect 407186 478258 407422 478494
rect 407186 471258 407422 471494
rect 407186 464258 407422 464494
rect 407186 457258 407422 457494
rect 407186 450258 407422 450494
rect 407186 443258 407422 443494
rect 407186 436258 407422 436494
rect 407186 429258 407422 429494
rect 407186 422258 407422 422494
rect 407186 415258 407422 415494
rect 407186 408258 407422 408494
rect 407186 401258 407422 401494
rect 407186 394258 407422 394494
rect 407186 387258 407422 387494
rect 407186 380258 407422 380494
rect 407186 373258 407422 373494
rect 407186 366258 407422 366494
rect 407186 359258 407422 359494
rect 407186 352258 407422 352494
rect 407186 345258 407422 345494
rect 407186 338258 407422 338494
rect 407186 331258 407422 331494
rect 407186 324258 407422 324494
rect 407186 317258 407422 317494
rect 407186 310258 407422 310494
rect 407186 303258 407422 303494
rect 407186 296258 407422 296494
rect 407186 289258 407422 289494
rect 407186 282258 407422 282494
rect 407186 275258 407422 275494
rect 407186 268258 407422 268494
rect 407186 261258 407422 261494
rect 407186 254258 407422 254494
rect 407186 247258 407422 247494
rect 407186 240258 407422 240494
rect 407186 233258 407422 233494
rect 407186 226258 407422 226494
rect 407186 219258 407422 219494
rect 407186 212258 407422 212494
rect 407186 205258 407422 205494
rect 407186 198258 407422 198494
rect 407186 191258 407422 191494
rect 407186 184258 407422 184494
rect 407186 177258 407422 177494
rect 407186 170258 407422 170494
rect 407186 163258 407422 163494
rect 407186 156258 407422 156494
rect 407186 149258 407422 149494
rect 407186 142258 407422 142494
rect 407186 135258 407422 135494
rect 407186 128258 407422 128494
rect 407186 121258 407422 121494
rect 407186 114258 407422 114494
rect 407186 107258 407422 107494
rect 407186 100258 407422 100494
rect 407186 93258 407422 93494
rect 407186 86258 407422 86494
rect 407186 79258 407422 79494
rect 407186 72258 407422 72494
rect 407186 65258 407422 65494
rect 407186 58258 407422 58494
rect 407186 51258 407422 51494
rect 407186 44258 407422 44494
rect 407186 37258 407422 37494
rect 407186 30258 407422 30494
rect 407186 23258 407422 23494
rect 407186 16258 407422 16494
rect 407186 9258 407422 9494
rect 407186 2258 407422 2494
rect 407186 -982 407422 -746
rect 407186 -1302 407422 -1066
rect 408918 705962 409154 706198
rect 408918 705642 409154 705878
rect 408918 696325 409154 696561
rect 408918 689325 409154 689561
rect 408918 682325 409154 682561
rect 408918 675325 409154 675561
rect 408918 668325 409154 668561
rect 408918 661325 409154 661561
rect 408918 654325 409154 654561
rect 408918 647325 409154 647561
rect 408918 640325 409154 640561
rect 408918 633325 409154 633561
rect 408918 626325 409154 626561
rect 408918 619325 409154 619561
rect 408918 612325 409154 612561
rect 408918 605325 409154 605561
rect 408918 598325 409154 598561
rect 408918 591325 409154 591561
rect 408918 584325 409154 584561
rect 408918 577325 409154 577561
rect 408918 570325 409154 570561
rect 408918 563325 409154 563561
rect 408918 556325 409154 556561
rect 408918 549325 409154 549561
rect 408918 542325 409154 542561
rect 408918 535325 409154 535561
rect 408918 528325 409154 528561
rect 408918 521325 409154 521561
rect 408918 514325 409154 514561
rect 408918 507325 409154 507561
rect 408918 500325 409154 500561
rect 408918 493325 409154 493561
rect 408918 486325 409154 486561
rect 408918 479325 409154 479561
rect 408918 472325 409154 472561
rect 408918 465325 409154 465561
rect 408918 458325 409154 458561
rect 408918 451325 409154 451561
rect 408918 444325 409154 444561
rect 408918 437325 409154 437561
rect 408918 430325 409154 430561
rect 408918 423325 409154 423561
rect 408918 416325 409154 416561
rect 408918 409325 409154 409561
rect 408918 402325 409154 402561
rect 408918 395325 409154 395561
rect 408918 388325 409154 388561
rect 408918 381325 409154 381561
rect 408918 374325 409154 374561
rect 408918 367325 409154 367561
rect 408918 360325 409154 360561
rect 408918 353325 409154 353561
rect 408918 346325 409154 346561
rect 408918 339325 409154 339561
rect 408918 332325 409154 332561
rect 408918 325325 409154 325561
rect 408918 318325 409154 318561
rect 408918 311325 409154 311561
rect 408918 304325 409154 304561
rect 408918 297325 409154 297561
rect 408918 290325 409154 290561
rect 408918 283325 409154 283561
rect 408918 276325 409154 276561
rect 408918 269325 409154 269561
rect 408918 262325 409154 262561
rect 408918 255325 409154 255561
rect 408918 248325 409154 248561
rect 408918 241325 409154 241561
rect 408918 234325 409154 234561
rect 408918 227325 409154 227561
rect 408918 220325 409154 220561
rect 408918 213325 409154 213561
rect 408918 206325 409154 206561
rect 408918 199325 409154 199561
rect 408918 192325 409154 192561
rect 408918 185325 409154 185561
rect 408918 178325 409154 178561
rect 408918 171325 409154 171561
rect 408918 164325 409154 164561
rect 408918 157325 409154 157561
rect 408918 150325 409154 150561
rect 408918 143325 409154 143561
rect 408918 136325 409154 136561
rect 408918 129325 409154 129561
rect 408918 122325 409154 122561
rect 408918 115325 409154 115561
rect 408918 108325 409154 108561
rect 408918 101325 409154 101561
rect 408918 94325 409154 94561
rect 408918 87325 409154 87561
rect 408918 80325 409154 80561
rect 408918 73325 409154 73561
rect 408918 66325 409154 66561
rect 408918 59325 409154 59561
rect 408918 52325 409154 52561
rect 408918 45325 409154 45561
rect 408918 38325 409154 38561
rect 408918 31325 409154 31561
rect 408918 24325 409154 24561
rect 408918 17325 409154 17561
rect 408918 10325 409154 10561
rect 408918 3325 409154 3561
rect 408918 -1942 409154 -1706
rect 408918 -2262 409154 -2026
rect 414186 705002 414422 705238
rect 414186 704682 414422 704918
rect 414186 695258 414422 695494
rect 414186 688258 414422 688494
rect 414186 681258 414422 681494
rect 414186 674258 414422 674494
rect 414186 667258 414422 667494
rect 414186 660258 414422 660494
rect 414186 653258 414422 653494
rect 414186 646258 414422 646494
rect 414186 639258 414422 639494
rect 414186 632258 414422 632494
rect 414186 625258 414422 625494
rect 414186 618258 414422 618494
rect 414186 611258 414422 611494
rect 414186 604258 414422 604494
rect 414186 597258 414422 597494
rect 414186 590258 414422 590494
rect 414186 583258 414422 583494
rect 414186 576258 414422 576494
rect 414186 569258 414422 569494
rect 414186 562258 414422 562494
rect 414186 555258 414422 555494
rect 414186 548258 414422 548494
rect 414186 541258 414422 541494
rect 414186 534258 414422 534494
rect 414186 527258 414422 527494
rect 414186 520258 414422 520494
rect 414186 513258 414422 513494
rect 414186 506258 414422 506494
rect 414186 499258 414422 499494
rect 414186 492258 414422 492494
rect 414186 485258 414422 485494
rect 414186 478258 414422 478494
rect 414186 471258 414422 471494
rect 414186 464258 414422 464494
rect 414186 457258 414422 457494
rect 414186 450258 414422 450494
rect 414186 443258 414422 443494
rect 414186 436258 414422 436494
rect 414186 429258 414422 429494
rect 414186 422258 414422 422494
rect 414186 415258 414422 415494
rect 414186 408258 414422 408494
rect 414186 401258 414422 401494
rect 414186 394258 414422 394494
rect 414186 387258 414422 387494
rect 414186 380258 414422 380494
rect 414186 373258 414422 373494
rect 414186 366258 414422 366494
rect 414186 359258 414422 359494
rect 414186 352258 414422 352494
rect 414186 345258 414422 345494
rect 414186 338258 414422 338494
rect 414186 331258 414422 331494
rect 414186 324258 414422 324494
rect 414186 317258 414422 317494
rect 414186 310258 414422 310494
rect 414186 303258 414422 303494
rect 414186 296258 414422 296494
rect 414186 289258 414422 289494
rect 414186 282258 414422 282494
rect 414186 275258 414422 275494
rect 414186 268258 414422 268494
rect 414186 261258 414422 261494
rect 414186 254258 414422 254494
rect 414186 247258 414422 247494
rect 414186 240258 414422 240494
rect 414186 233258 414422 233494
rect 414186 226258 414422 226494
rect 414186 219258 414422 219494
rect 414186 212258 414422 212494
rect 414186 205258 414422 205494
rect 414186 198258 414422 198494
rect 414186 191258 414422 191494
rect 414186 184258 414422 184494
rect 414186 177258 414422 177494
rect 414186 170258 414422 170494
rect 414186 163258 414422 163494
rect 414186 156258 414422 156494
rect 414186 149258 414422 149494
rect 414186 142258 414422 142494
rect 414186 135258 414422 135494
rect 414186 128258 414422 128494
rect 414186 121258 414422 121494
rect 414186 114258 414422 114494
rect 414186 107258 414422 107494
rect 414186 100258 414422 100494
rect 414186 93258 414422 93494
rect 414186 86258 414422 86494
rect 414186 79258 414422 79494
rect 414186 72258 414422 72494
rect 414186 65258 414422 65494
rect 414186 58258 414422 58494
rect 414186 51258 414422 51494
rect 414186 44258 414422 44494
rect 414186 37258 414422 37494
rect 414186 30258 414422 30494
rect 414186 23258 414422 23494
rect 414186 16258 414422 16494
rect 414186 9258 414422 9494
rect 414186 2258 414422 2494
rect 414186 -982 414422 -746
rect 414186 -1302 414422 -1066
rect 415918 705962 416154 706198
rect 415918 705642 416154 705878
rect 415918 696325 416154 696561
rect 415918 689325 416154 689561
rect 415918 682325 416154 682561
rect 415918 675325 416154 675561
rect 415918 668325 416154 668561
rect 415918 661325 416154 661561
rect 415918 654325 416154 654561
rect 415918 647325 416154 647561
rect 415918 640325 416154 640561
rect 415918 633325 416154 633561
rect 415918 626325 416154 626561
rect 415918 619325 416154 619561
rect 415918 612325 416154 612561
rect 415918 605325 416154 605561
rect 415918 598325 416154 598561
rect 415918 591325 416154 591561
rect 415918 584325 416154 584561
rect 415918 577325 416154 577561
rect 415918 570325 416154 570561
rect 415918 563325 416154 563561
rect 415918 556325 416154 556561
rect 415918 549325 416154 549561
rect 415918 542325 416154 542561
rect 415918 535325 416154 535561
rect 415918 528325 416154 528561
rect 415918 521325 416154 521561
rect 415918 514325 416154 514561
rect 415918 507325 416154 507561
rect 415918 500325 416154 500561
rect 415918 493325 416154 493561
rect 415918 486325 416154 486561
rect 415918 479325 416154 479561
rect 415918 472325 416154 472561
rect 415918 465325 416154 465561
rect 415918 458325 416154 458561
rect 415918 451325 416154 451561
rect 415918 444325 416154 444561
rect 415918 437325 416154 437561
rect 415918 430325 416154 430561
rect 415918 423325 416154 423561
rect 415918 416325 416154 416561
rect 415918 409325 416154 409561
rect 415918 402325 416154 402561
rect 415918 395325 416154 395561
rect 415918 388325 416154 388561
rect 415918 381325 416154 381561
rect 415918 374325 416154 374561
rect 415918 367325 416154 367561
rect 415918 360325 416154 360561
rect 415918 353325 416154 353561
rect 415918 346325 416154 346561
rect 415918 339325 416154 339561
rect 415918 332325 416154 332561
rect 415918 325325 416154 325561
rect 415918 318325 416154 318561
rect 415918 311325 416154 311561
rect 415918 304325 416154 304561
rect 415918 297325 416154 297561
rect 415918 290325 416154 290561
rect 415918 283325 416154 283561
rect 415918 276325 416154 276561
rect 415918 269325 416154 269561
rect 415918 262325 416154 262561
rect 415918 255325 416154 255561
rect 415918 248325 416154 248561
rect 415918 241325 416154 241561
rect 415918 234325 416154 234561
rect 415918 227325 416154 227561
rect 415918 220325 416154 220561
rect 415918 213325 416154 213561
rect 415918 206325 416154 206561
rect 415918 199325 416154 199561
rect 415918 192325 416154 192561
rect 415918 185325 416154 185561
rect 415918 178325 416154 178561
rect 415918 171325 416154 171561
rect 415918 164325 416154 164561
rect 415918 157325 416154 157561
rect 415918 150325 416154 150561
rect 415918 143325 416154 143561
rect 415918 136325 416154 136561
rect 415918 129325 416154 129561
rect 415918 122325 416154 122561
rect 415918 115325 416154 115561
rect 415918 108325 416154 108561
rect 415918 101325 416154 101561
rect 415918 94325 416154 94561
rect 415918 87325 416154 87561
rect 415918 80325 416154 80561
rect 415918 73325 416154 73561
rect 415918 66325 416154 66561
rect 415918 59325 416154 59561
rect 415918 52325 416154 52561
rect 415918 45325 416154 45561
rect 415918 38325 416154 38561
rect 415918 31325 416154 31561
rect 415918 24325 416154 24561
rect 415918 17325 416154 17561
rect 415918 10325 416154 10561
rect 415918 3325 416154 3561
rect 415918 -1942 416154 -1706
rect 415918 -2262 416154 -2026
rect 421186 705002 421422 705238
rect 421186 704682 421422 704918
rect 421186 695258 421422 695494
rect 421186 688258 421422 688494
rect 421186 681258 421422 681494
rect 421186 674258 421422 674494
rect 421186 667258 421422 667494
rect 421186 660258 421422 660494
rect 421186 653258 421422 653494
rect 421186 646258 421422 646494
rect 421186 639258 421422 639494
rect 421186 632258 421422 632494
rect 421186 625258 421422 625494
rect 421186 618258 421422 618494
rect 421186 611258 421422 611494
rect 421186 604258 421422 604494
rect 421186 597258 421422 597494
rect 421186 590258 421422 590494
rect 421186 583258 421422 583494
rect 421186 576258 421422 576494
rect 421186 569258 421422 569494
rect 421186 562258 421422 562494
rect 421186 555258 421422 555494
rect 421186 548258 421422 548494
rect 421186 541258 421422 541494
rect 421186 534258 421422 534494
rect 421186 527258 421422 527494
rect 421186 520258 421422 520494
rect 421186 513258 421422 513494
rect 421186 506258 421422 506494
rect 421186 499258 421422 499494
rect 421186 492258 421422 492494
rect 421186 485258 421422 485494
rect 421186 478258 421422 478494
rect 421186 471258 421422 471494
rect 421186 464258 421422 464494
rect 421186 457258 421422 457494
rect 421186 450258 421422 450494
rect 421186 443258 421422 443494
rect 421186 436258 421422 436494
rect 421186 429258 421422 429494
rect 421186 422258 421422 422494
rect 421186 415258 421422 415494
rect 421186 408258 421422 408494
rect 421186 401258 421422 401494
rect 421186 394258 421422 394494
rect 421186 387258 421422 387494
rect 421186 380258 421422 380494
rect 421186 373258 421422 373494
rect 421186 366258 421422 366494
rect 421186 359258 421422 359494
rect 421186 352258 421422 352494
rect 421186 345258 421422 345494
rect 421186 338258 421422 338494
rect 421186 331258 421422 331494
rect 421186 324258 421422 324494
rect 421186 317258 421422 317494
rect 421186 310258 421422 310494
rect 421186 303258 421422 303494
rect 421186 296258 421422 296494
rect 421186 289258 421422 289494
rect 421186 282258 421422 282494
rect 421186 275258 421422 275494
rect 421186 268258 421422 268494
rect 421186 261258 421422 261494
rect 421186 254258 421422 254494
rect 421186 247258 421422 247494
rect 421186 240258 421422 240494
rect 421186 233258 421422 233494
rect 421186 226258 421422 226494
rect 421186 219258 421422 219494
rect 421186 212258 421422 212494
rect 421186 205258 421422 205494
rect 421186 198258 421422 198494
rect 421186 191258 421422 191494
rect 421186 184258 421422 184494
rect 421186 177258 421422 177494
rect 421186 170258 421422 170494
rect 421186 163258 421422 163494
rect 421186 156258 421422 156494
rect 421186 149258 421422 149494
rect 421186 142258 421422 142494
rect 421186 135258 421422 135494
rect 421186 128258 421422 128494
rect 421186 121258 421422 121494
rect 421186 114258 421422 114494
rect 421186 107258 421422 107494
rect 421186 100258 421422 100494
rect 421186 93258 421422 93494
rect 421186 86258 421422 86494
rect 421186 79258 421422 79494
rect 421186 72258 421422 72494
rect 421186 65258 421422 65494
rect 421186 58258 421422 58494
rect 421186 51258 421422 51494
rect 421186 44258 421422 44494
rect 421186 37258 421422 37494
rect 421186 30258 421422 30494
rect 421186 23258 421422 23494
rect 421186 16258 421422 16494
rect 421186 9258 421422 9494
rect 421186 2258 421422 2494
rect 421186 -982 421422 -746
rect 421186 -1302 421422 -1066
rect 422918 705962 423154 706198
rect 422918 705642 423154 705878
rect 422918 696325 423154 696561
rect 422918 689325 423154 689561
rect 422918 682325 423154 682561
rect 422918 675325 423154 675561
rect 422918 668325 423154 668561
rect 422918 661325 423154 661561
rect 422918 654325 423154 654561
rect 422918 647325 423154 647561
rect 422918 640325 423154 640561
rect 422918 633325 423154 633561
rect 422918 626325 423154 626561
rect 422918 619325 423154 619561
rect 422918 612325 423154 612561
rect 422918 605325 423154 605561
rect 422918 598325 423154 598561
rect 422918 591325 423154 591561
rect 422918 584325 423154 584561
rect 422918 577325 423154 577561
rect 422918 570325 423154 570561
rect 422918 563325 423154 563561
rect 422918 556325 423154 556561
rect 422918 549325 423154 549561
rect 422918 542325 423154 542561
rect 422918 535325 423154 535561
rect 422918 528325 423154 528561
rect 422918 521325 423154 521561
rect 422918 514325 423154 514561
rect 422918 507325 423154 507561
rect 422918 500325 423154 500561
rect 422918 493325 423154 493561
rect 422918 486325 423154 486561
rect 422918 479325 423154 479561
rect 422918 472325 423154 472561
rect 422918 465325 423154 465561
rect 422918 458325 423154 458561
rect 422918 451325 423154 451561
rect 422918 444325 423154 444561
rect 422918 437325 423154 437561
rect 422918 430325 423154 430561
rect 422918 423325 423154 423561
rect 422918 416325 423154 416561
rect 422918 409325 423154 409561
rect 422918 402325 423154 402561
rect 422918 395325 423154 395561
rect 422918 388325 423154 388561
rect 422918 381325 423154 381561
rect 422918 374325 423154 374561
rect 422918 367325 423154 367561
rect 422918 360325 423154 360561
rect 422918 353325 423154 353561
rect 422918 346325 423154 346561
rect 422918 339325 423154 339561
rect 422918 332325 423154 332561
rect 422918 325325 423154 325561
rect 422918 318325 423154 318561
rect 422918 311325 423154 311561
rect 422918 304325 423154 304561
rect 422918 297325 423154 297561
rect 422918 290325 423154 290561
rect 422918 283325 423154 283561
rect 422918 276325 423154 276561
rect 422918 269325 423154 269561
rect 422918 262325 423154 262561
rect 422918 255325 423154 255561
rect 422918 248325 423154 248561
rect 422918 241325 423154 241561
rect 422918 234325 423154 234561
rect 422918 227325 423154 227561
rect 422918 220325 423154 220561
rect 422918 213325 423154 213561
rect 422918 206325 423154 206561
rect 422918 199325 423154 199561
rect 422918 192325 423154 192561
rect 422918 185325 423154 185561
rect 422918 178325 423154 178561
rect 422918 171325 423154 171561
rect 422918 164325 423154 164561
rect 422918 157325 423154 157561
rect 422918 150325 423154 150561
rect 422918 143325 423154 143561
rect 422918 136325 423154 136561
rect 422918 129325 423154 129561
rect 422918 122325 423154 122561
rect 422918 115325 423154 115561
rect 422918 108325 423154 108561
rect 422918 101325 423154 101561
rect 422918 94325 423154 94561
rect 422918 87325 423154 87561
rect 422918 80325 423154 80561
rect 422918 73325 423154 73561
rect 422918 66325 423154 66561
rect 422918 59325 423154 59561
rect 422918 52325 423154 52561
rect 422918 45325 423154 45561
rect 422918 38325 423154 38561
rect 422918 31325 423154 31561
rect 422918 24325 423154 24561
rect 422918 17325 423154 17561
rect 422918 10325 423154 10561
rect 422918 3325 423154 3561
rect 422918 -1942 423154 -1706
rect 422918 -2262 423154 -2026
rect 428186 705002 428422 705238
rect 428186 704682 428422 704918
rect 428186 695258 428422 695494
rect 428186 688258 428422 688494
rect 428186 681258 428422 681494
rect 428186 674258 428422 674494
rect 428186 667258 428422 667494
rect 428186 660258 428422 660494
rect 428186 653258 428422 653494
rect 428186 646258 428422 646494
rect 428186 639258 428422 639494
rect 428186 632258 428422 632494
rect 428186 625258 428422 625494
rect 428186 618258 428422 618494
rect 428186 611258 428422 611494
rect 428186 604258 428422 604494
rect 428186 597258 428422 597494
rect 428186 590258 428422 590494
rect 428186 583258 428422 583494
rect 428186 576258 428422 576494
rect 428186 569258 428422 569494
rect 428186 562258 428422 562494
rect 428186 555258 428422 555494
rect 428186 548258 428422 548494
rect 428186 541258 428422 541494
rect 428186 534258 428422 534494
rect 428186 527258 428422 527494
rect 428186 520258 428422 520494
rect 428186 513258 428422 513494
rect 428186 506258 428422 506494
rect 428186 499258 428422 499494
rect 428186 492258 428422 492494
rect 428186 485258 428422 485494
rect 428186 478258 428422 478494
rect 428186 471258 428422 471494
rect 428186 464258 428422 464494
rect 428186 457258 428422 457494
rect 428186 450258 428422 450494
rect 428186 443258 428422 443494
rect 428186 436258 428422 436494
rect 428186 429258 428422 429494
rect 428186 422258 428422 422494
rect 428186 415258 428422 415494
rect 428186 408258 428422 408494
rect 428186 401258 428422 401494
rect 428186 394258 428422 394494
rect 428186 387258 428422 387494
rect 428186 380258 428422 380494
rect 428186 373258 428422 373494
rect 428186 366258 428422 366494
rect 428186 359258 428422 359494
rect 428186 352258 428422 352494
rect 428186 345258 428422 345494
rect 428186 338258 428422 338494
rect 428186 331258 428422 331494
rect 428186 324258 428422 324494
rect 428186 317258 428422 317494
rect 428186 310258 428422 310494
rect 428186 303258 428422 303494
rect 428186 296258 428422 296494
rect 428186 289258 428422 289494
rect 428186 282258 428422 282494
rect 428186 275258 428422 275494
rect 428186 268258 428422 268494
rect 428186 261258 428422 261494
rect 428186 254258 428422 254494
rect 428186 247258 428422 247494
rect 428186 240258 428422 240494
rect 428186 233258 428422 233494
rect 428186 226258 428422 226494
rect 428186 219258 428422 219494
rect 428186 212258 428422 212494
rect 428186 205258 428422 205494
rect 428186 198258 428422 198494
rect 428186 191258 428422 191494
rect 428186 184258 428422 184494
rect 428186 177258 428422 177494
rect 428186 170258 428422 170494
rect 428186 163258 428422 163494
rect 428186 156258 428422 156494
rect 428186 149258 428422 149494
rect 428186 142258 428422 142494
rect 428186 135258 428422 135494
rect 428186 128258 428422 128494
rect 428186 121258 428422 121494
rect 428186 114258 428422 114494
rect 428186 107258 428422 107494
rect 428186 100258 428422 100494
rect 428186 93258 428422 93494
rect 428186 86258 428422 86494
rect 428186 79258 428422 79494
rect 428186 72258 428422 72494
rect 428186 65258 428422 65494
rect 428186 58258 428422 58494
rect 428186 51258 428422 51494
rect 428186 44258 428422 44494
rect 428186 37258 428422 37494
rect 428186 30258 428422 30494
rect 428186 23258 428422 23494
rect 428186 16258 428422 16494
rect 428186 9258 428422 9494
rect 428186 2258 428422 2494
rect 428186 -982 428422 -746
rect 428186 -1302 428422 -1066
rect 429918 705962 430154 706198
rect 429918 705642 430154 705878
rect 429918 696325 430154 696561
rect 429918 689325 430154 689561
rect 429918 682325 430154 682561
rect 429918 675325 430154 675561
rect 429918 668325 430154 668561
rect 429918 661325 430154 661561
rect 429918 654325 430154 654561
rect 429918 647325 430154 647561
rect 429918 640325 430154 640561
rect 429918 633325 430154 633561
rect 429918 626325 430154 626561
rect 429918 619325 430154 619561
rect 429918 612325 430154 612561
rect 429918 605325 430154 605561
rect 429918 598325 430154 598561
rect 429918 591325 430154 591561
rect 429918 584325 430154 584561
rect 429918 577325 430154 577561
rect 429918 570325 430154 570561
rect 429918 563325 430154 563561
rect 429918 556325 430154 556561
rect 429918 549325 430154 549561
rect 429918 542325 430154 542561
rect 429918 535325 430154 535561
rect 429918 528325 430154 528561
rect 429918 521325 430154 521561
rect 429918 514325 430154 514561
rect 429918 507325 430154 507561
rect 429918 500325 430154 500561
rect 429918 493325 430154 493561
rect 429918 486325 430154 486561
rect 429918 479325 430154 479561
rect 429918 472325 430154 472561
rect 429918 465325 430154 465561
rect 429918 458325 430154 458561
rect 429918 451325 430154 451561
rect 429918 444325 430154 444561
rect 429918 437325 430154 437561
rect 429918 430325 430154 430561
rect 429918 423325 430154 423561
rect 429918 416325 430154 416561
rect 429918 409325 430154 409561
rect 429918 402325 430154 402561
rect 429918 395325 430154 395561
rect 429918 388325 430154 388561
rect 429918 381325 430154 381561
rect 429918 374325 430154 374561
rect 429918 367325 430154 367561
rect 429918 360325 430154 360561
rect 429918 353325 430154 353561
rect 429918 346325 430154 346561
rect 429918 339325 430154 339561
rect 429918 332325 430154 332561
rect 429918 325325 430154 325561
rect 429918 318325 430154 318561
rect 429918 311325 430154 311561
rect 429918 304325 430154 304561
rect 429918 297325 430154 297561
rect 429918 290325 430154 290561
rect 429918 283325 430154 283561
rect 429918 276325 430154 276561
rect 429918 269325 430154 269561
rect 429918 262325 430154 262561
rect 429918 255325 430154 255561
rect 429918 248325 430154 248561
rect 429918 241325 430154 241561
rect 429918 234325 430154 234561
rect 429918 227325 430154 227561
rect 429918 220325 430154 220561
rect 429918 213325 430154 213561
rect 429918 206325 430154 206561
rect 429918 199325 430154 199561
rect 429918 192325 430154 192561
rect 429918 185325 430154 185561
rect 429918 178325 430154 178561
rect 429918 171325 430154 171561
rect 429918 164325 430154 164561
rect 429918 157325 430154 157561
rect 429918 150325 430154 150561
rect 429918 143325 430154 143561
rect 429918 136325 430154 136561
rect 429918 129325 430154 129561
rect 429918 122325 430154 122561
rect 429918 115325 430154 115561
rect 429918 108325 430154 108561
rect 429918 101325 430154 101561
rect 429918 94325 430154 94561
rect 429918 87325 430154 87561
rect 429918 80325 430154 80561
rect 429918 73325 430154 73561
rect 429918 66325 430154 66561
rect 429918 59325 430154 59561
rect 429918 52325 430154 52561
rect 429918 45325 430154 45561
rect 429918 38325 430154 38561
rect 429918 31325 430154 31561
rect 429918 24325 430154 24561
rect 429918 17325 430154 17561
rect 429918 10325 430154 10561
rect 429918 3325 430154 3561
rect 429918 -1942 430154 -1706
rect 429918 -2262 430154 -2026
rect 435186 705002 435422 705238
rect 435186 704682 435422 704918
rect 435186 695258 435422 695494
rect 435186 688258 435422 688494
rect 435186 681258 435422 681494
rect 435186 674258 435422 674494
rect 435186 667258 435422 667494
rect 435186 660258 435422 660494
rect 435186 653258 435422 653494
rect 435186 646258 435422 646494
rect 435186 639258 435422 639494
rect 435186 632258 435422 632494
rect 435186 625258 435422 625494
rect 435186 618258 435422 618494
rect 435186 611258 435422 611494
rect 435186 604258 435422 604494
rect 435186 597258 435422 597494
rect 435186 590258 435422 590494
rect 435186 583258 435422 583494
rect 435186 576258 435422 576494
rect 435186 569258 435422 569494
rect 435186 562258 435422 562494
rect 435186 555258 435422 555494
rect 435186 548258 435422 548494
rect 435186 541258 435422 541494
rect 435186 534258 435422 534494
rect 435186 527258 435422 527494
rect 435186 520258 435422 520494
rect 435186 513258 435422 513494
rect 435186 506258 435422 506494
rect 435186 499258 435422 499494
rect 435186 492258 435422 492494
rect 435186 485258 435422 485494
rect 435186 478258 435422 478494
rect 435186 471258 435422 471494
rect 435186 464258 435422 464494
rect 435186 457258 435422 457494
rect 435186 450258 435422 450494
rect 435186 443258 435422 443494
rect 435186 436258 435422 436494
rect 435186 429258 435422 429494
rect 435186 422258 435422 422494
rect 435186 415258 435422 415494
rect 435186 408258 435422 408494
rect 435186 401258 435422 401494
rect 435186 394258 435422 394494
rect 435186 387258 435422 387494
rect 435186 380258 435422 380494
rect 435186 373258 435422 373494
rect 435186 366258 435422 366494
rect 435186 359258 435422 359494
rect 435186 352258 435422 352494
rect 435186 345258 435422 345494
rect 435186 338258 435422 338494
rect 435186 331258 435422 331494
rect 435186 324258 435422 324494
rect 435186 317258 435422 317494
rect 435186 310258 435422 310494
rect 435186 303258 435422 303494
rect 435186 296258 435422 296494
rect 435186 289258 435422 289494
rect 435186 282258 435422 282494
rect 435186 275258 435422 275494
rect 435186 268258 435422 268494
rect 435186 261258 435422 261494
rect 435186 254258 435422 254494
rect 435186 247258 435422 247494
rect 435186 240258 435422 240494
rect 435186 233258 435422 233494
rect 435186 226258 435422 226494
rect 435186 219258 435422 219494
rect 435186 212258 435422 212494
rect 435186 205258 435422 205494
rect 435186 198258 435422 198494
rect 435186 191258 435422 191494
rect 435186 184258 435422 184494
rect 435186 177258 435422 177494
rect 435186 170258 435422 170494
rect 435186 163258 435422 163494
rect 435186 156258 435422 156494
rect 435186 149258 435422 149494
rect 435186 142258 435422 142494
rect 435186 135258 435422 135494
rect 435186 128258 435422 128494
rect 435186 121258 435422 121494
rect 435186 114258 435422 114494
rect 435186 107258 435422 107494
rect 435186 100258 435422 100494
rect 435186 93258 435422 93494
rect 435186 86258 435422 86494
rect 435186 79258 435422 79494
rect 435186 72258 435422 72494
rect 435186 65258 435422 65494
rect 435186 58258 435422 58494
rect 435186 51258 435422 51494
rect 435186 44258 435422 44494
rect 435186 37258 435422 37494
rect 435186 30258 435422 30494
rect 435186 23258 435422 23494
rect 435186 16258 435422 16494
rect 435186 9258 435422 9494
rect 435186 2258 435422 2494
rect 435186 -982 435422 -746
rect 435186 -1302 435422 -1066
rect 436918 705962 437154 706198
rect 436918 705642 437154 705878
rect 436918 696325 437154 696561
rect 436918 689325 437154 689561
rect 436918 682325 437154 682561
rect 436918 675325 437154 675561
rect 436918 668325 437154 668561
rect 436918 661325 437154 661561
rect 436918 654325 437154 654561
rect 436918 647325 437154 647561
rect 436918 640325 437154 640561
rect 436918 633325 437154 633561
rect 436918 626325 437154 626561
rect 436918 619325 437154 619561
rect 436918 612325 437154 612561
rect 436918 605325 437154 605561
rect 436918 598325 437154 598561
rect 436918 591325 437154 591561
rect 436918 584325 437154 584561
rect 436918 577325 437154 577561
rect 436918 570325 437154 570561
rect 436918 563325 437154 563561
rect 436918 556325 437154 556561
rect 436918 549325 437154 549561
rect 436918 542325 437154 542561
rect 436918 535325 437154 535561
rect 436918 528325 437154 528561
rect 436918 521325 437154 521561
rect 436918 514325 437154 514561
rect 436918 507325 437154 507561
rect 436918 500325 437154 500561
rect 436918 493325 437154 493561
rect 436918 486325 437154 486561
rect 436918 479325 437154 479561
rect 436918 472325 437154 472561
rect 436918 465325 437154 465561
rect 436918 458325 437154 458561
rect 436918 451325 437154 451561
rect 436918 444325 437154 444561
rect 436918 437325 437154 437561
rect 436918 430325 437154 430561
rect 436918 423325 437154 423561
rect 436918 416325 437154 416561
rect 436918 409325 437154 409561
rect 436918 402325 437154 402561
rect 436918 395325 437154 395561
rect 436918 388325 437154 388561
rect 436918 381325 437154 381561
rect 436918 374325 437154 374561
rect 436918 367325 437154 367561
rect 436918 360325 437154 360561
rect 436918 353325 437154 353561
rect 436918 346325 437154 346561
rect 436918 339325 437154 339561
rect 436918 332325 437154 332561
rect 436918 325325 437154 325561
rect 436918 318325 437154 318561
rect 436918 311325 437154 311561
rect 436918 304325 437154 304561
rect 436918 297325 437154 297561
rect 436918 290325 437154 290561
rect 436918 283325 437154 283561
rect 436918 276325 437154 276561
rect 436918 269325 437154 269561
rect 436918 262325 437154 262561
rect 436918 255325 437154 255561
rect 436918 248325 437154 248561
rect 436918 241325 437154 241561
rect 436918 234325 437154 234561
rect 436918 227325 437154 227561
rect 436918 220325 437154 220561
rect 436918 213325 437154 213561
rect 436918 206325 437154 206561
rect 436918 199325 437154 199561
rect 436918 192325 437154 192561
rect 436918 185325 437154 185561
rect 436918 178325 437154 178561
rect 436918 171325 437154 171561
rect 436918 164325 437154 164561
rect 436918 157325 437154 157561
rect 436918 150325 437154 150561
rect 436918 143325 437154 143561
rect 436918 136325 437154 136561
rect 436918 129325 437154 129561
rect 436918 122325 437154 122561
rect 436918 115325 437154 115561
rect 436918 108325 437154 108561
rect 436918 101325 437154 101561
rect 436918 94325 437154 94561
rect 436918 87325 437154 87561
rect 436918 80325 437154 80561
rect 436918 73325 437154 73561
rect 436918 66325 437154 66561
rect 436918 59325 437154 59561
rect 436918 52325 437154 52561
rect 436918 45325 437154 45561
rect 436918 38325 437154 38561
rect 436918 31325 437154 31561
rect 436918 24325 437154 24561
rect 436918 17325 437154 17561
rect 436918 10325 437154 10561
rect 436918 3325 437154 3561
rect 436918 -1942 437154 -1706
rect 436918 -2262 437154 -2026
rect 442186 705002 442422 705238
rect 442186 704682 442422 704918
rect 442186 695258 442422 695494
rect 442186 688258 442422 688494
rect 442186 681258 442422 681494
rect 442186 674258 442422 674494
rect 442186 667258 442422 667494
rect 442186 660258 442422 660494
rect 442186 653258 442422 653494
rect 442186 646258 442422 646494
rect 442186 639258 442422 639494
rect 442186 632258 442422 632494
rect 442186 625258 442422 625494
rect 442186 618258 442422 618494
rect 442186 611258 442422 611494
rect 442186 604258 442422 604494
rect 442186 597258 442422 597494
rect 442186 590258 442422 590494
rect 442186 583258 442422 583494
rect 442186 576258 442422 576494
rect 442186 569258 442422 569494
rect 442186 562258 442422 562494
rect 442186 555258 442422 555494
rect 442186 548258 442422 548494
rect 442186 541258 442422 541494
rect 442186 534258 442422 534494
rect 442186 527258 442422 527494
rect 442186 520258 442422 520494
rect 442186 513258 442422 513494
rect 442186 506258 442422 506494
rect 442186 499258 442422 499494
rect 442186 492258 442422 492494
rect 442186 485258 442422 485494
rect 442186 478258 442422 478494
rect 442186 471258 442422 471494
rect 442186 464258 442422 464494
rect 442186 457258 442422 457494
rect 442186 450258 442422 450494
rect 442186 443258 442422 443494
rect 442186 436258 442422 436494
rect 442186 429258 442422 429494
rect 442186 422258 442422 422494
rect 442186 415258 442422 415494
rect 442186 408258 442422 408494
rect 442186 401258 442422 401494
rect 442186 394258 442422 394494
rect 442186 387258 442422 387494
rect 442186 380258 442422 380494
rect 442186 373258 442422 373494
rect 442186 366258 442422 366494
rect 442186 359258 442422 359494
rect 442186 352258 442422 352494
rect 442186 345258 442422 345494
rect 442186 338258 442422 338494
rect 442186 331258 442422 331494
rect 442186 324258 442422 324494
rect 442186 317258 442422 317494
rect 442186 310258 442422 310494
rect 442186 303258 442422 303494
rect 442186 296258 442422 296494
rect 442186 289258 442422 289494
rect 442186 282258 442422 282494
rect 442186 275258 442422 275494
rect 442186 268258 442422 268494
rect 442186 261258 442422 261494
rect 442186 254258 442422 254494
rect 442186 247258 442422 247494
rect 442186 240258 442422 240494
rect 442186 233258 442422 233494
rect 442186 226258 442422 226494
rect 442186 219258 442422 219494
rect 442186 212258 442422 212494
rect 442186 205258 442422 205494
rect 442186 198258 442422 198494
rect 442186 191258 442422 191494
rect 442186 184258 442422 184494
rect 442186 177258 442422 177494
rect 442186 170258 442422 170494
rect 442186 163258 442422 163494
rect 442186 156258 442422 156494
rect 442186 149258 442422 149494
rect 442186 142258 442422 142494
rect 442186 135258 442422 135494
rect 442186 128258 442422 128494
rect 442186 121258 442422 121494
rect 442186 114258 442422 114494
rect 442186 107258 442422 107494
rect 442186 100258 442422 100494
rect 442186 93258 442422 93494
rect 442186 86258 442422 86494
rect 442186 79258 442422 79494
rect 442186 72258 442422 72494
rect 442186 65258 442422 65494
rect 442186 58258 442422 58494
rect 442186 51258 442422 51494
rect 442186 44258 442422 44494
rect 442186 37258 442422 37494
rect 442186 30258 442422 30494
rect 442186 23258 442422 23494
rect 442186 16258 442422 16494
rect 442186 9258 442422 9494
rect 442186 2258 442422 2494
rect 442186 -982 442422 -746
rect 442186 -1302 442422 -1066
rect 443918 705962 444154 706198
rect 443918 705642 444154 705878
rect 443918 696325 444154 696561
rect 443918 689325 444154 689561
rect 443918 682325 444154 682561
rect 443918 675325 444154 675561
rect 443918 668325 444154 668561
rect 443918 661325 444154 661561
rect 443918 654325 444154 654561
rect 443918 647325 444154 647561
rect 443918 640325 444154 640561
rect 443918 633325 444154 633561
rect 443918 626325 444154 626561
rect 443918 619325 444154 619561
rect 443918 612325 444154 612561
rect 443918 605325 444154 605561
rect 443918 598325 444154 598561
rect 443918 591325 444154 591561
rect 443918 584325 444154 584561
rect 443918 577325 444154 577561
rect 443918 570325 444154 570561
rect 443918 563325 444154 563561
rect 443918 556325 444154 556561
rect 443918 549325 444154 549561
rect 443918 542325 444154 542561
rect 443918 535325 444154 535561
rect 443918 528325 444154 528561
rect 443918 521325 444154 521561
rect 443918 514325 444154 514561
rect 443918 507325 444154 507561
rect 443918 500325 444154 500561
rect 443918 493325 444154 493561
rect 443918 486325 444154 486561
rect 443918 479325 444154 479561
rect 443918 472325 444154 472561
rect 443918 465325 444154 465561
rect 443918 458325 444154 458561
rect 443918 451325 444154 451561
rect 443918 444325 444154 444561
rect 443918 437325 444154 437561
rect 443918 430325 444154 430561
rect 443918 423325 444154 423561
rect 443918 416325 444154 416561
rect 443918 409325 444154 409561
rect 443918 402325 444154 402561
rect 443918 395325 444154 395561
rect 443918 388325 444154 388561
rect 443918 381325 444154 381561
rect 443918 374325 444154 374561
rect 443918 367325 444154 367561
rect 443918 360325 444154 360561
rect 443918 353325 444154 353561
rect 443918 346325 444154 346561
rect 443918 339325 444154 339561
rect 443918 332325 444154 332561
rect 443918 325325 444154 325561
rect 443918 318325 444154 318561
rect 443918 311325 444154 311561
rect 443918 304325 444154 304561
rect 443918 297325 444154 297561
rect 443918 290325 444154 290561
rect 443918 283325 444154 283561
rect 443918 276325 444154 276561
rect 443918 269325 444154 269561
rect 443918 262325 444154 262561
rect 443918 255325 444154 255561
rect 443918 248325 444154 248561
rect 443918 241325 444154 241561
rect 443918 234325 444154 234561
rect 443918 227325 444154 227561
rect 443918 220325 444154 220561
rect 443918 213325 444154 213561
rect 443918 206325 444154 206561
rect 443918 199325 444154 199561
rect 443918 192325 444154 192561
rect 443918 185325 444154 185561
rect 443918 178325 444154 178561
rect 443918 171325 444154 171561
rect 443918 164325 444154 164561
rect 443918 157325 444154 157561
rect 443918 150325 444154 150561
rect 443918 143325 444154 143561
rect 443918 136325 444154 136561
rect 443918 129325 444154 129561
rect 443918 122325 444154 122561
rect 443918 115325 444154 115561
rect 443918 108325 444154 108561
rect 443918 101325 444154 101561
rect 443918 94325 444154 94561
rect 443918 87325 444154 87561
rect 443918 80325 444154 80561
rect 443918 73325 444154 73561
rect 443918 66325 444154 66561
rect 443918 59325 444154 59561
rect 443918 52325 444154 52561
rect 443918 45325 444154 45561
rect 443918 38325 444154 38561
rect 443918 31325 444154 31561
rect 443918 24325 444154 24561
rect 443918 17325 444154 17561
rect 443918 10325 444154 10561
rect 443918 3325 444154 3561
rect 443918 -1942 444154 -1706
rect 443918 -2262 444154 -2026
rect 449186 705002 449422 705238
rect 449186 704682 449422 704918
rect 449186 695258 449422 695494
rect 449186 688258 449422 688494
rect 449186 681258 449422 681494
rect 449186 674258 449422 674494
rect 449186 667258 449422 667494
rect 449186 660258 449422 660494
rect 449186 653258 449422 653494
rect 449186 646258 449422 646494
rect 449186 639258 449422 639494
rect 449186 632258 449422 632494
rect 449186 625258 449422 625494
rect 449186 618258 449422 618494
rect 449186 611258 449422 611494
rect 449186 604258 449422 604494
rect 449186 597258 449422 597494
rect 449186 590258 449422 590494
rect 449186 583258 449422 583494
rect 449186 576258 449422 576494
rect 449186 569258 449422 569494
rect 449186 562258 449422 562494
rect 449186 555258 449422 555494
rect 449186 548258 449422 548494
rect 449186 541258 449422 541494
rect 449186 534258 449422 534494
rect 449186 527258 449422 527494
rect 449186 520258 449422 520494
rect 449186 513258 449422 513494
rect 449186 506258 449422 506494
rect 449186 499258 449422 499494
rect 449186 492258 449422 492494
rect 449186 485258 449422 485494
rect 449186 478258 449422 478494
rect 449186 471258 449422 471494
rect 449186 464258 449422 464494
rect 449186 457258 449422 457494
rect 449186 450258 449422 450494
rect 449186 443258 449422 443494
rect 449186 436258 449422 436494
rect 449186 429258 449422 429494
rect 449186 422258 449422 422494
rect 449186 415258 449422 415494
rect 449186 408258 449422 408494
rect 449186 401258 449422 401494
rect 449186 394258 449422 394494
rect 449186 387258 449422 387494
rect 449186 380258 449422 380494
rect 449186 373258 449422 373494
rect 449186 366258 449422 366494
rect 449186 359258 449422 359494
rect 449186 352258 449422 352494
rect 449186 345258 449422 345494
rect 449186 338258 449422 338494
rect 449186 331258 449422 331494
rect 449186 324258 449422 324494
rect 449186 317258 449422 317494
rect 449186 310258 449422 310494
rect 449186 303258 449422 303494
rect 449186 296258 449422 296494
rect 449186 289258 449422 289494
rect 449186 282258 449422 282494
rect 449186 275258 449422 275494
rect 449186 268258 449422 268494
rect 449186 261258 449422 261494
rect 449186 254258 449422 254494
rect 449186 247258 449422 247494
rect 449186 240258 449422 240494
rect 449186 233258 449422 233494
rect 449186 226258 449422 226494
rect 449186 219258 449422 219494
rect 449186 212258 449422 212494
rect 449186 205258 449422 205494
rect 449186 198258 449422 198494
rect 449186 191258 449422 191494
rect 449186 184258 449422 184494
rect 449186 177258 449422 177494
rect 449186 170258 449422 170494
rect 449186 163258 449422 163494
rect 449186 156258 449422 156494
rect 449186 149258 449422 149494
rect 449186 142258 449422 142494
rect 449186 135258 449422 135494
rect 449186 128258 449422 128494
rect 449186 121258 449422 121494
rect 449186 114258 449422 114494
rect 449186 107258 449422 107494
rect 449186 100258 449422 100494
rect 449186 93258 449422 93494
rect 449186 86258 449422 86494
rect 449186 79258 449422 79494
rect 449186 72258 449422 72494
rect 449186 65258 449422 65494
rect 449186 58258 449422 58494
rect 449186 51258 449422 51494
rect 449186 44258 449422 44494
rect 449186 37258 449422 37494
rect 449186 30258 449422 30494
rect 449186 23258 449422 23494
rect 449186 16258 449422 16494
rect 449186 9258 449422 9494
rect 449186 2258 449422 2494
rect 449186 -982 449422 -746
rect 449186 -1302 449422 -1066
rect 450918 705962 451154 706198
rect 450918 705642 451154 705878
rect 450918 696325 451154 696561
rect 450918 689325 451154 689561
rect 450918 682325 451154 682561
rect 450918 675325 451154 675561
rect 450918 668325 451154 668561
rect 450918 661325 451154 661561
rect 450918 654325 451154 654561
rect 450918 647325 451154 647561
rect 450918 640325 451154 640561
rect 450918 633325 451154 633561
rect 450918 626325 451154 626561
rect 450918 619325 451154 619561
rect 450918 612325 451154 612561
rect 450918 605325 451154 605561
rect 450918 598325 451154 598561
rect 450918 591325 451154 591561
rect 450918 584325 451154 584561
rect 450918 577325 451154 577561
rect 450918 570325 451154 570561
rect 450918 563325 451154 563561
rect 450918 556325 451154 556561
rect 450918 549325 451154 549561
rect 450918 542325 451154 542561
rect 450918 535325 451154 535561
rect 450918 528325 451154 528561
rect 450918 521325 451154 521561
rect 450918 514325 451154 514561
rect 450918 507325 451154 507561
rect 450918 500325 451154 500561
rect 450918 493325 451154 493561
rect 450918 486325 451154 486561
rect 450918 479325 451154 479561
rect 450918 472325 451154 472561
rect 450918 465325 451154 465561
rect 450918 458325 451154 458561
rect 450918 451325 451154 451561
rect 450918 444325 451154 444561
rect 450918 437325 451154 437561
rect 450918 430325 451154 430561
rect 450918 423325 451154 423561
rect 450918 416325 451154 416561
rect 450918 409325 451154 409561
rect 450918 402325 451154 402561
rect 450918 395325 451154 395561
rect 450918 388325 451154 388561
rect 450918 381325 451154 381561
rect 450918 374325 451154 374561
rect 450918 367325 451154 367561
rect 450918 360325 451154 360561
rect 450918 353325 451154 353561
rect 450918 346325 451154 346561
rect 450918 339325 451154 339561
rect 450918 332325 451154 332561
rect 450918 325325 451154 325561
rect 450918 318325 451154 318561
rect 450918 311325 451154 311561
rect 450918 304325 451154 304561
rect 450918 297325 451154 297561
rect 450918 290325 451154 290561
rect 450918 283325 451154 283561
rect 450918 276325 451154 276561
rect 450918 269325 451154 269561
rect 450918 262325 451154 262561
rect 450918 255325 451154 255561
rect 450918 248325 451154 248561
rect 450918 241325 451154 241561
rect 450918 234325 451154 234561
rect 450918 227325 451154 227561
rect 450918 220325 451154 220561
rect 450918 213325 451154 213561
rect 450918 206325 451154 206561
rect 450918 199325 451154 199561
rect 450918 192325 451154 192561
rect 450918 185325 451154 185561
rect 450918 178325 451154 178561
rect 450918 171325 451154 171561
rect 450918 164325 451154 164561
rect 450918 157325 451154 157561
rect 450918 150325 451154 150561
rect 450918 143325 451154 143561
rect 450918 136325 451154 136561
rect 450918 129325 451154 129561
rect 450918 122325 451154 122561
rect 450918 115325 451154 115561
rect 450918 108325 451154 108561
rect 450918 101325 451154 101561
rect 450918 94325 451154 94561
rect 450918 87325 451154 87561
rect 450918 80325 451154 80561
rect 450918 73325 451154 73561
rect 450918 66325 451154 66561
rect 450918 59325 451154 59561
rect 450918 52325 451154 52561
rect 450918 45325 451154 45561
rect 450918 38325 451154 38561
rect 450918 31325 451154 31561
rect 450918 24325 451154 24561
rect 450918 17325 451154 17561
rect 450918 10325 451154 10561
rect 450918 3325 451154 3561
rect 450918 -1942 451154 -1706
rect 450918 -2262 451154 -2026
rect 456186 705002 456422 705238
rect 456186 704682 456422 704918
rect 456186 695258 456422 695494
rect 456186 688258 456422 688494
rect 456186 681258 456422 681494
rect 456186 674258 456422 674494
rect 456186 667258 456422 667494
rect 456186 660258 456422 660494
rect 456186 653258 456422 653494
rect 456186 646258 456422 646494
rect 456186 639258 456422 639494
rect 456186 632258 456422 632494
rect 456186 625258 456422 625494
rect 456186 618258 456422 618494
rect 456186 611258 456422 611494
rect 456186 604258 456422 604494
rect 456186 597258 456422 597494
rect 456186 590258 456422 590494
rect 456186 583258 456422 583494
rect 456186 576258 456422 576494
rect 456186 569258 456422 569494
rect 456186 562258 456422 562494
rect 456186 555258 456422 555494
rect 456186 548258 456422 548494
rect 456186 541258 456422 541494
rect 456186 534258 456422 534494
rect 456186 527258 456422 527494
rect 456186 520258 456422 520494
rect 456186 513258 456422 513494
rect 456186 506258 456422 506494
rect 456186 499258 456422 499494
rect 456186 492258 456422 492494
rect 456186 485258 456422 485494
rect 456186 478258 456422 478494
rect 456186 471258 456422 471494
rect 456186 464258 456422 464494
rect 456186 457258 456422 457494
rect 456186 450258 456422 450494
rect 456186 443258 456422 443494
rect 456186 436258 456422 436494
rect 456186 429258 456422 429494
rect 456186 422258 456422 422494
rect 456186 415258 456422 415494
rect 456186 408258 456422 408494
rect 456186 401258 456422 401494
rect 456186 394258 456422 394494
rect 456186 387258 456422 387494
rect 456186 380258 456422 380494
rect 456186 373258 456422 373494
rect 456186 366258 456422 366494
rect 456186 359258 456422 359494
rect 456186 352258 456422 352494
rect 456186 345258 456422 345494
rect 456186 338258 456422 338494
rect 456186 331258 456422 331494
rect 456186 324258 456422 324494
rect 456186 317258 456422 317494
rect 456186 310258 456422 310494
rect 456186 303258 456422 303494
rect 456186 296258 456422 296494
rect 456186 289258 456422 289494
rect 456186 282258 456422 282494
rect 456186 275258 456422 275494
rect 456186 268258 456422 268494
rect 456186 261258 456422 261494
rect 456186 254258 456422 254494
rect 456186 247258 456422 247494
rect 456186 240258 456422 240494
rect 456186 233258 456422 233494
rect 456186 226258 456422 226494
rect 456186 219258 456422 219494
rect 456186 212258 456422 212494
rect 456186 205258 456422 205494
rect 456186 198258 456422 198494
rect 456186 191258 456422 191494
rect 456186 184258 456422 184494
rect 456186 177258 456422 177494
rect 456186 170258 456422 170494
rect 456186 163258 456422 163494
rect 456186 156258 456422 156494
rect 456186 149258 456422 149494
rect 456186 142258 456422 142494
rect 456186 135258 456422 135494
rect 456186 128258 456422 128494
rect 456186 121258 456422 121494
rect 456186 114258 456422 114494
rect 456186 107258 456422 107494
rect 456186 100258 456422 100494
rect 456186 93258 456422 93494
rect 456186 86258 456422 86494
rect 456186 79258 456422 79494
rect 456186 72258 456422 72494
rect 456186 65258 456422 65494
rect 456186 58258 456422 58494
rect 456186 51258 456422 51494
rect 456186 44258 456422 44494
rect 456186 37258 456422 37494
rect 456186 30258 456422 30494
rect 456186 23258 456422 23494
rect 456186 16258 456422 16494
rect 456186 9258 456422 9494
rect 456186 2258 456422 2494
rect 456186 -982 456422 -746
rect 456186 -1302 456422 -1066
rect 457918 705962 458154 706198
rect 457918 705642 458154 705878
rect 457918 696325 458154 696561
rect 457918 689325 458154 689561
rect 457918 682325 458154 682561
rect 457918 675325 458154 675561
rect 457918 668325 458154 668561
rect 457918 661325 458154 661561
rect 457918 654325 458154 654561
rect 457918 647325 458154 647561
rect 457918 640325 458154 640561
rect 457918 633325 458154 633561
rect 457918 626325 458154 626561
rect 457918 619325 458154 619561
rect 457918 612325 458154 612561
rect 457918 605325 458154 605561
rect 457918 598325 458154 598561
rect 457918 591325 458154 591561
rect 457918 584325 458154 584561
rect 457918 577325 458154 577561
rect 457918 570325 458154 570561
rect 457918 563325 458154 563561
rect 457918 556325 458154 556561
rect 457918 549325 458154 549561
rect 457918 542325 458154 542561
rect 457918 535325 458154 535561
rect 457918 528325 458154 528561
rect 457918 521325 458154 521561
rect 457918 514325 458154 514561
rect 457918 507325 458154 507561
rect 457918 500325 458154 500561
rect 457918 493325 458154 493561
rect 457918 486325 458154 486561
rect 457918 479325 458154 479561
rect 457918 472325 458154 472561
rect 457918 465325 458154 465561
rect 457918 458325 458154 458561
rect 457918 451325 458154 451561
rect 457918 444325 458154 444561
rect 457918 437325 458154 437561
rect 457918 430325 458154 430561
rect 457918 423325 458154 423561
rect 457918 416325 458154 416561
rect 457918 409325 458154 409561
rect 457918 402325 458154 402561
rect 457918 395325 458154 395561
rect 457918 388325 458154 388561
rect 457918 381325 458154 381561
rect 457918 374325 458154 374561
rect 457918 367325 458154 367561
rect 457918 360325 458154 360561
rect 457918 353325 458154 353561
rect 457918 346325 458154 346561
rect 457918 339325 458154 339561
rect 457918 332325 458154 332561
rect 457918 325325 458154 325561
rect 457918 318325 458154 318561
rect 457918 311325 458154 311561
rect 457918 304325 458154 304561
rect 457918 297325 458154 297561
rect 457918 290325 458154 290561
rect 457918 283325 458154 283561
rect 457918 276325 458154 276561
rect 457918 269325 458154 269561
rect 457918 262325 458154 262561
rect 457918 255325 458154 255561
rect 457918 248325 458154 248561
rect 457918 241325 458154 241561
rect 457918 234325 458154 234561
rect 457918 227325 458154 227561
rect 457918 220325 458154 220561
rect 457918 213325 458154 213561
rect 457918 206325 458154 206561
rect 457918 199325 458154 199561
rect 457918 192325 458154 192561
rect 457918 185325 458154 185561
rect 457918 178325 458154 178561
rect 457918 171325 458154 171561
rect 457918 164325 458154 164561
rect 457918 157325 458154 157561
rect 457918 150325 458154 150561
rect 457918 143325 458154 143561
rect 457918 136325 458154 136561
rect 457918 129325 458154 129561
rect 457918 122325 458154 122561
rect 457918 115325 458154 115561
rect 457918 108325 458154 108561
rect 457918 101325 458154 101561
rect 457918 94325 458154 94561
rect 457918 87325 458154 87561
rect 457918 80325 458154 80561
rect 457918 73325 458154 73561
rect 457918 66325 458154 66561
rect 457918 59325 458154 59561
rect 457918 52325 458154 52561
rect 457918 45325 458154 45561
rect 457918 38325 458154 38561
rect 457918 31325 458154 31561
rect 457918 24325 458154 24561
rect 457918 17325 458154 17561
rect 457918 10325 458154 10561
rect 457918 3325 458154 3561
rect 457918 -1942 458154 -1706
rect 457918 -2262 458154 -2026
rect 463186 705002 463422 705238
rect 463186 704682 463422 704918
rect 463186 695258 463422 695494
rect 463186 688258 463422 688494
rect 463186 681258 463422 681494
rect 463186 674258 463422 674494
rect 463186 667258 463422 667494
rect 463186 660258 463422 660494
rect 463186 653258 463422 653494
rect 463186 646258 463422 646494
rect 463186 639258 463422 639494
rect 463186 632258 463422 632494
rect 463186 625258 463422 625494
rect 463186 618258 463422 618494
rect 463186 611258 463422 611494
rect 463186 604258 463422 604494
rect 463186 597258 463422 597494
rect 463186 590258 463422 590494
rect 463186 583258 463422 583494
rect 463186 576258 463422 576494
rect 463186 569258 463422 569494
rect 463186 562258 463422 562494
rect 463186 555258 463422 555494
rect 463186 548258 463422 548494
rect 463186 541258 463422 541494
rect 463186 534258 463422 534494
rect 463186 527258 463422 527494
rect 463186 520258 463422 520494
rect 463186 513258 463422 513494
rect 463186 506258 463422 506494
rect 463186 499258 463422 499494
rect 463186 492258 463422 492494
rect 463186 485258 463422 485494
rect 463186 478258 463422 478494
rect 463186 471258 463422 471494
rect 463186 464258 463422 464494
rect 463186 457258 463422 457494
rect 463186 450258 463422 450494
rect 463186 443258 463422 443494
rect 463186 436258 463422 436494
rect 463186 429258 463422 429494
rect 463186 422258 463422 422494
rect 463186 415258 463422 415494
rect 463186 408258 463422 408494
rect 463186 401258 463422 401494
rect 463186 394258 463422 394494
rect 463186 387258 463422 387494
rect 463186 380258 463422 380494
rect 463186 373258 463422 373494
rect 463186 366258 463422 366494
rect 463186 359258 463422 359494
rect 463186 352258 463422 352494
rect 463186 345258 463422 345494
rect 463186 338258 463422 338494
rect 463186 331258 463422 331494
rect 463186 324258 463422 324494
rect 463186 317258 463422 317494
rect 463186 310258 463422 310494
rect 463186 303258 463422 303494
rect 463186 296258 463422 296494
rect 463186 289258 463422 289494
rect 463186 282258 463422 282494
rect 463186 275258 463422 275494
rect 463186 268258 463422 268494
rect 463186 261258 463422 261494
rect 463186 254258 463422 254494
rect 463186 247258 463422 247494
rect 463186 240258 463422 240494
rect 463186 233258 463422 233494
rect 463186 226258 463422 226494
rect 463186 219258 463422 219494
rect 463186 212258 463422 212494
rect 463186 205258 463422 205494
rect 463186 198258 463422 198494
rect 463186 191258 463422 191494
rect 463186 184258 463422 184494
rect 463186 177258 463422 177494
rect 463186 170258 463422 170494
rect 463186 163258 463422 163494
rect 463186 156258 463422 156494
rect 463186 149258 463422 149494
rect 463186 142258 463422 142494
rect 463186 135258 463422 135494
rect 463186 128258 463422 128494
rect 463186 121258 463422 121494
rect 463186 114258 463422 114494
rect 463186 107258 463422 107494
rect 463186 100258 463422 100494
rect 463186 93258 463422 93494
rect 463186 86258 463422 86494
rect 463186 79258 463422 79494
rect 463186 72258 463422 72494
rect 463186 65258 463422 65494
rect 463186 58258 463422 58494
rect 463186 51258 463422 51494
rect 463186 44258 463422 44494
rect 463186 37258 463422 37494
rect 463186 30258 463422 30494
rect 463186 23258 463422 23494
rect 463186 16258 463422 16494
rect 463186 9258 463422 9494
rect 463186 2258 463422 2494
rect 463186 -982 463422 -746
rect 463186 -1302 463422 -1066
rect 464918 705962 465154 706198
rect 464918 705642 465154 705878
rect 464918 696325 465154 696561
rect 464918 689325 465154 689561
rect 464918 682325 465154 682561
rect 464918 675325 465154 675561
rect 464918 668325 465154 668561
rect 464918 661325 465154 661561
rect 464918 654325 465154 654561
rect 464918 647325 465154 647561
rect 464918 640325 465154 640561
rect 464918 633325 465154 633561
rect 464918 626325 465154 626561
rect 464918 619325 465154 619561
rect 464918 612325 465154 612561
rect 464918 605325 465154 605561
rect 464918 598325 465154 598561
rect 464918 591325 465154 591561
rect 464918 584325 465154 584561
rect 464918 577325 465154 577561
rect 464918 570325 465154 570561
rect 464918 563325 465154 563561
rect 464918 556325 465154 556561
rect 464918 549325 465154 549561
rect 464918 542325 465154 542561
rect 464918 535325 465154 535561
rect 464918 528325 465154 528561
rect 464918 521325 465154 521561
rect 464918 514325 465154 514561
rect 464918 507325 465154 507561
rect 464918 500325 465154 500561
rect 464918 493325 465154 493561
rect 464918 486325 465154 486561
rect 464918 479325 465154 479561
rect 464918 472325 465154 472561
rect 464918 465325 465154 465561
rect 464918 458325 465154 458561
rect 464918 451325 465154 451561
rect 464918 444325 465154 444561
rect 464918 437325 465154 437561
rect 464918 430325 465154 430561
rect 464918 423325 465154 423561
rect 464918 416325 465154 416561
rect 464918 409325 465154 409561
rect 464918 402325 465154 402561
rect 464918 395325 465154 395561
rect 464918 388325 465154 388561
rect 464918 381325 465154 381561
rect 464918 374325 465154 374561
rect 464918 367325 465154 367561
rect 464918 360325 465154 360561
rect 464918 353325 465154 353561
rect 464918 346325 465154 346561
rect 464918 339325 465154 339561
rect 464918 332325 465154 332561
rect 464918 325325 465154 325561
rect 464918 318325 465154 318561
rect 464918 311325 465154 311561
rect 464918 304325 465154 304561
rect 464918 297325 465154 297561
rect 464918 290325 465154 290561
rect 464918 283325 465154 283561
rect 464918 276325 465154 276561
rect 464918 269325 465154 269561
rect 464918 262325 465154 262561
rect 464918 255325 465154 255561
rect 464918 248325 465154 248561
rect 464918 241325 465154 241561
rect 464918 234325 465154 234561
rect 464918 227325 465154 227561
rect 464918 220325 465154 220561
rect 464918 213325 465154 213561
rect 464918 206325 465154 206561
rect 464918 199325 465154 199561
rect 464918 192325 465154 192561
rect 464918 185325 465154 185561
rect 464918 178325 465154 178561
rect 464918 171325 465154 171561
rect 464918 164325 465154 164561
rect 464918 157325 465154 157561
rect 464918 150325 465154 150561
rect 464918 143325 465154 143561
rect 464918 136325 465154 136561
rect 464918 129325 465154 129561
rect 464918 122325 465154 122561
rect 464918 115325 465154 115561
rect 464918 108325 465154 108561
rect 464918 101325 465154 101561
rect 464918 94325 465154 94561
rect 464918 87325 465154 87561
rect 464918 80325 465154 80561
rect 464918 73325 465154 73561
rect 464918 66325 465154 66561
rect 464918 59325 465154 59561
rect 464918 52325 465154 52561
rect 464918 45325 465154 45561
rect 464918 38325 465154 38561
rect 464918 31325 465154 31561
rect 464918 24325 465154 24561
rect 464918 17325 465154 17561
rect 464918 10325 465154 10561
rect 464918 3325 465154 3561
rect 464918 -1942 465154 -1706
rect 464918 -2262 465154 -2026
rect 470186 705002 470422 705238
rect 470186 704682 470422 704918
rect 470186 695258 470422 695494
rect 470186 688258 470422 688494
rect 470186 681258 470422 681494
rect 470186 674258 470422 674494
rect 470186 667258 470422 667494
rect 470186 660258 470422 660494
rect 470186 653258 470422 653494
rect 470186 646258 470422 646494
rect 470186 639258 470422 639494
rect 470186 632258 470422 632494
rect 470186 625258 470422 625494
rect 470186 618258 470422 618494
rect 470186 611258 470422 611494
rect 470186 604258 470422 604494
rect 470186 597258 470422 597494
rect 470186 590258 470422 590494
rect 470186 583258 470422 583494
rect 470186 576258 470422 576494
rect 470186 569258 470422 569494
rect 470186 562258 470422 562494
rect 470186 555258 470422 555494
rect 470186 548258 470422 548494
rect 470186 541258 470422 541494
rect 470186 534258 470422 534494
rect 470186 527258 470422 527494
rect 470186 520258 470422 520494
rect 470186 513258 470422 513494
rect 470186 506258 470422 506494
rect 470186 499258 470422 499494
rect 470186 492258 470422 492494
rect 470186 485258 470422 485494
rect 470186 478258 470422 478494
rect 470186 471258 470422 471494
rect 470186 464258 470422 464494
rect 470186 457258 470422 457494
rect 470186 450258 470422 450494
rect 470186 443258 470422 443494
rect 470186 436258 470422 436494
rect 470186 429258 470422 429494
rect 470186 422258 470422 422494
rect 470186 415258 470422 415494
rect 470186 408258 470422 408494
rect 470186 401258 470422 401494
rect 470186 394258 470422 394494
rect 470186 387258 470422 387494
rect 470186 380258 470422 380494
rect 470186 373258 470422 373494
rect 470186 366258 470422 366494
rect 470186 359258 470422 359494
rect 470186 352258 470422 352494
rect 470186 345258 470422 345494
rect 470186 338258 470422 338494
rect 470186 331258 470422 331494
rect 470186 324258 470422 324494
rect 470186 317258 470422 317494
rect 470186 310258 470422 310494
rect 470186 303258 470422 303494
rect 470186 296258 470422 296494
rect 470186 289258 470422 289494
rect 470186 282258 470422 282494
rect 470186 275258 470422 275494
rect 470186 268258 470422 268494
rect 470186 261258 470422 261494
rect 470186 254258 470422 254494
rect 470186 247258 470422 247494
rect 470186 240258 470422 240494
rect 470186 233258 470422 233494
rect 470186 226258 470422 226494
rect 470186 219258 470422 219494
rect 470186 212258 470422 212494
rect 470186 205258 470422 205494
rect 470186 198258 470422 198494
rect 470186 191258 470422 191494
rect 470186 184258 470422 184494
rect 470186 177258 470422 177494
rect 470186 170258 470422 170494
rect 470186 163258 470422 163494
rect 470186 156258 470422 156494
rect 470186 149258 470422 149494
rect 470186 142258 470422 142494
rect 470186 135258 470422 135494
rect 470186 128258 470422 128494
rect 470186 121258 470422 121494
rect 470186 114258 470422 114494
rect 470186 107258 470422 107494
rect 470186 100258 470422 100494
rect 470186 93258 470422 93494
rect 470186 86258 470422 86494
rect 470186 79258 470422 79494
rect 470186 72258 470422 72494
rect 470186 65258 470422 65494
rect 470186 58258 470422 58494
rect 470186 51258 470422 51494
rect 470186 44258 470422 44494
rect 470186 37258 470422 37494
rect 470186 30258 470422 30494
rect 470186 23258 470422 23494
rect 470186 16258 470422 16494
rect 470186 9258 470422 9494
rect 470186 2258 470422 2494
rect 470186 -982 470422 -746
rect 470186 -1302 470422 -1066
rect 471918 705962 472154 706198
rect 471918 705642 472154 705878
rect 471918 696325 472154 696561
rect 471918 689325 472154 689561
rect 471918 682325 472154 682561
rect 471918 675325 472154 675561
rect 471918 668325 472154 668561
rect 471918 661325 472154 661561
rect 471918 654325 472154 654561
rect 471918 647325 472154 647561
rect 471918 640325 472154 640561
rect 471918 633325 472154 633561
rect 471918 626325 472154 626561
rect 471918 619325 472154 619561
rect 471918 612325 472154 612561
rect 471918 605325 472154 605561
rect 471918 598325 472154 598561
rect 471918 591325 472154 591561
rect 471918 584325 472154 584561
rect 471918 577325 472154 577561
rect 471918 570325 472154 570561
rect 471918 563325 472154 563561
rect 471918 556325 472154 556561
rect 471918 549325 472154 549561
rect 471918 542325 472154 542561
rect 471918 535325 472154 535561
rect 471918 528325 472154 528561
rect 471918 521325 472154 521561
rect 471918 514325 472154 514561
rect 471918 507325 472154 507561
rect 471918 500325 472154 500561
rect 471918 493325 472154 493561
rect 471918 486325 472154 486561
rect 471918 479325 472154 479561
rect 471918 472325 472154 472561
rect 471918 465325 472154 465561
rect 471918 458325 472154 458561
rect 471918 451325 472154 451561
rect 471918 444325 472154 444561
rect 471918 437325 472154 437561
rect 471918 430325 472154 430561
rect 471918 423325 472154 423561
rect 471918 416325 472154 416561
rect 471918 409325 472154 409561
rect 471918 402325 472154 402561
rect 471918 395325 472154 395561
rect 471918 388325 472154 388561
rect 471918 381325 472154 381561
rect 471918 374325 472154 374561
rect 471918 367325 472154 367561
rect 471918 360325 472154 360561
rect 471918 353325 472154 353561
rect 471918 346325 472154 346561
rect 471918 339325 472154 339561
rect 471918 332325 472154 332561
rect 471918 325325 472154 325561
rect 471918 318325 472154 318561
rect 471918 311325 472154 311561
rect 471918 304325 472154 304561
rect 471918 297325 472154 297561
rect 471918 290325 472154 290561
rect 471918 283325 472154 283561
rect 471918 276325 472154 276561
rect 471918 269325 472154 269561
rect 471918 262325 472154 262561
rect 471918 255325 472154 255561
rect 471918 248325 472154 248561
rect 471918 241325 472154 241561
rect 471918 234325 472154 234561
rect 471918 227325 472154 227561
rect 471918 220325 472154 220561
rect 471918 213325 472154 213561
rect 471918 206325 472154 206561
rect 471918 199325 472154 199561
rect 471918 192325 472154 192561
rect 471918 185325 472154 185561
rect 471918 178325 472154 178561
rect 471918 171325 472154 171561
rect 471918 164325 472154 164561
rect 471918 157325 472154 157561
rect 471918 150325 472154 150561
rect 471918 143325 472154 143561
rect 471918 136325 472154 136561
rect 471918 129325 472154 129561
rect 471918 122325 472154 122561
rect 471918 115325 472154 115561
rect 471918 108325 472154 108561
rect 471918 101325 472154 101561
rect 471918 94325 472154 94561
rect 471918 87325 472154 87561
rect 471918 80325 472154 80561
rect 471918 73325 472154 73561
rect 471918 66325 472154 66561
rect 471918 59325 472154 59561
rect 471918 52325 472154 52561
rect 471918 45325 472154 45561
rect 471918 38325 472154 38561
rect 471918 31325 472154 31561
rect 471918 24325 472154 24561
rect 471918 17325 472154 17561
rect 471918 10325 472154 10561
rect 471918 3325 472154 3561
rect 471918 -1942 472154 -1706
rect 471918 -2262 472154 -2026
rect 477186 705002 477422 705238
rect 477186 704682 477422 704918
rect 477186 695258 477422 695494
rect 477186 688258 477422 688494
rect 477186 681258 477422 681494
rect 477186 674258 477422 674494
rect 477186 667258 477422 667494
rect 477186 660258 477422 660494
rect 477186 653258 477422 653494
rect 477186 646258 477422 646494
rect 477186 639258 477422 639494
rect 477186 632258 477422 632494
rect 477186 625258 477422 625494
rect 477186 618258 477422 618494
rect 477186 611258 477422 611494
rect 477186 604258 477422 604494
rect 477186 597258 477422 597494
rect 477186 590258 477422 590494
rect 477186 583258 477422 583494
rect 477186 576258 477422 576494
rect 477186 569258 477422 569494
rect 477186 562258 477422 562494
rect 477186 555258 477422 555494
rect 477186 548258 477422 548494
rect 477186 541258 477422 541494
rect 477186 534258 477422 534494
rect 477186 527258 477422 527494
rect 477186 520258 477422 520494
rect 477186 513258 477422 513494
rect 477186 506258 477422 506494
rect 477186 499258 477422 499494
rect 477186 492258 477422 492494
rect 477186 485258 477422 485494
rect 477186 478258 477422 478494
rect 477186 471258 477422 471494
rect 477186 464258 477422 464494
rect 477186 457258 477422 457494
rect 477186 450258 477422 450494
rect 477186 443258 477422 443494
rect 477186 436258 477422 436494
rect 477186 429258 477422 429494
rect 477186 422258 477422 422494
rect 477186 415258 477422 415494
rect 477186 408258 477422 408494
rect 477186 401258 477422 401494
rect 477186 394258 477422 394494
rect 477186 387258 477422 387494
rect 477186 380258 477422 380494
rect 477186 373258 477422 373494
rect 477186 366258 477422 366494
rect 477186 359258 477422 359494
rect 477186 352258 477422 352494
rect 477186 345258 477422 345494
rect 477186 338258 477422 338494
rect 477186 331258 477422 331494
rect 477186 324258 477422 324494
rect 477186 317258 477422 317494
rect 477186 310258 477422 310494
rect 477186 303258 477422 303494
rect 477186 296258 477422 296494
rect 477186 289258 477422 289494
rect 477186 282258 477422 282494
rect 477186 275258 477422 275494
rect 477186 268258 477422 268494
rect 477186 261258 477422 261494
rect 477186 254258 477422 254494
rect 477186 247258 477422 247494
rect 477186 240258 477422 240494
rect 477186 233258 477422 233494
rect 477186 226258 477422 226494
rect 477186 219258 477422 219494
rect 477186 212258 477422 212494
rect 477186 205258 477422 205494
rect 477186 198258 477422 198494
rect 477186 191258 477422 191494
rect 477186 184258 477422 184494
rect 477186 177258 477422 177494
rect 477186 170258 477422 170494
rect 477186 163258 477422 163494
rect 477186 156258 477422 156494
rect 477186 149258 477422 149494
rect 477186 142258 477422 142494
rect 477186 135258 477422 135494
rect 477186 128258 477422 128494
rect 477186 121258 477422 121494
rect 477186 114258 477422 114494
rect 477186 107258 477422 107494
rect 477186 100258 477422 100494
rect 477186 93258 477422 93494
rect 477186 86258 477422 86494
rect 477186 79258 477422 79494
rect 477186 72258 477422 72494
rect 477186 65258 477422 65494
rect 477186 58258 477422 58494
rect 477186 51258 477422 51494
rect 477186 44258 477422 44494
rect 477186 37258 477422 37494
rect 477186 30258 477422 30494
rect 477186 23258 477422 23494
rect 477186 16258 477422 16494
rect 477186 9258 477422 9494
rect 477186 2258 477422 2494
rect 477186 -982 477422 -746
rect 477186 -1302 477422 -1066
rect 478918 705962 479154 706198
rect 478918 705642 479154 705878
rect 478918 696325 479154 696561
rect 478918 689325 479154 689561
rect 478918 682325 479154 682561
rect 478918 675325 479154 675561
rect 478918 668325 479154 668561
rect 478918 661325 479154 661561
rect 478918 654325 479154 654561
rect 478918 647325 479154 647561
rect 478918 640325 479154 640561
rect 478918 633325 479154 633561
rect 478918 626325 479154 626561
rect 478918 619325 479154 619561
rect 478918 612325 479154 612561
rect 478918 605325 479154 605561
rect 478918 598325 479154 598561
rect 478918 591325 479154 591561
rect 478918 584325 479154 584561
rect 478918 577325 479154 577561
rect 478918 570325 479154 570561
rect 478918 563325 479154 563561
rect 478918 556325 479154 556561
rect 478918 549325 479154 549561
rect 478918 542325 479154 542561
rect 478918 535325 479154 535561
rect 478918 528325 479154 528561
rect 478918 521325 479154 521561
rect 478918 514325 479154 514561
rect 478918 507325 479154 507561
rect 478918 500325 479154 500561
rect 478918 493325 479154 493561
rect 478918 486325 479154 486561
rect 478918 479325 479154 479561
rect 478918 472325 479154 472561
rect 478918 465325 479154 465561
rect 478918 458325 479154 458561
rect 478918 451325 479154 451561
rect 478918 444325 479154 444561
rect 478918 437325 479154 437561
rect 478918 430325 479154 430561
rect 478918 423325 479154 423561
rect 478918 416325 479154 416561
rect 478918 409325 479154 409561
rect 478918 402325 479154 402561
rect 478918 395325 479154 395561
rect 478918 388325 479154 388561
rect 478918 381325 479154 381561
rect 478918 374325 479154 374561
rect 478918 367325 479154 367561
rect 478918 360325 479154 360561
rect 478918 353325 479154 353561
rect 478918 346325 479154 346561
rect 478918 339325 479154 339561
rect 478918 332325 479154 332561
rect 478918 325325 479154 325561
rect 478918 318325 479154 318561
rect 478918 311325 479154 311561
rect 478918 304325 479154 304561
rect 478918 297325 479154 297561
rect 478918 290325 479154 290561
rect 478918 283325 479154 283561
rect 478918 276325 479154 276561
rect 478918 269325 479154 269561
rect 478918 262325 479154 262561
rect 478918 255325 479154 255561
rect 478918 248325 479154 248561
rect 478918 241325 479154 241561
rect 478918 234325 479154 234561
rect 478918 227325 479154 227561
rect 478918 220325 479154 220561
rect 478918 213325 479154 213561
rect 478918 206325 479154 206561
rect 478918 199325 479154 199561
rect 478918 192325 479154 192561
rect 478918 185325 479154 185561
rect 478918 178325 479154 178561
rect 478918 171325 479154 171561
rect 478918 164325 479154 164561
rect 478918 157325 479154 157561
rect 478918 150325 479154 150561
rect 478918 143325 479154 143561
rect 478918 136325 479154 136561
rect 478918 129325 479154 129561
rect 478918 122325 479154 122561
rect 478918 115325 479154 115561
rect 478918 108325 479154 108561
rect 478918 101325 479154 101561
rect 478918 94325 479154 94561
rect 478918 87325 479154 87561
rect 478918 80325 479154 80561
rect 478918 73325 479154 73561
rect 478918 66325 479154 66561
rect 478918 59325 479154 59561
rect 478918 52325 479154 52561
rect 478918 45325 479154 45561
rect 478918 38325 479154 38561
rect 478918 31325 479154 31561
rect 478918 24325 479154 24561
rect 478918 17325 479154 17561
rect 478918 10325 479154 10561
rect 478918 3325 479154 3561
rect 478918 -1942 479154 -1706
rect 478918 -2262 479154 -2026
rect 484186 705002 484422 705238
rect 484186 704682 484422 704918
rect 484186 695258 484422 695494
rect 484186 688258 484422 688494
rect 484186 681258 484422 681494
rect 484186 674258 484422 674494
rect 484186 667258 484422 667494
rect 484186 660258 484422 660494
rect 484186 653258 484422 653494
rect 484186 646258 484422 646494
rect 484186 639258 484422 639494
rect 484186 632258 484422 632494
rect 484186 625258 484422 625494
rect 484186 618258 484422 618494
rect 484186 611258 484422 611494
rect 484186 604258 484422 604494
rect 484186 597258 484422 597494
rect 484186 590258 484422 590494
rect 484186 583258 484422 583494
rect 484186 576258 484422 576494
rect 484186 569258 484422 569494
rect 484186 562258 484422 562494
rect 484186 555258 484422 555494
rect 484186 548258 484422 548494
rect 484186 541258 484422 541494
rect 484186 534258 484422 534494
rect 484186 527258 484422 527494
rect 484186 520258 484422 520494
rect 484186 513258 484422 513494
rect 484186 506258 484422 506494
rect 484186 499258 484422 499494
rect 484186 492258 484422 492494
rect 484186 485258 484422 485494
rect 484186 478258 484422 478494
rect 484186 471258 484422 471494
rect 484186 464258 484422 464494
rect 484186 457258 484422 457494
rect 484186 450258 484422 450494
rect 484186 443258 484422 443494
rect 484186 436258 484422 436494
rect 484186 429258 484422 429494
rect 484186 422258 484422 422494
rect 484186 415258 484422 415494
rect 484186 408258 484422 408494
rect 484186 401258 484422 401494
rect 484186 394258 484422 394494
rect 484186 387258 484422 387494
rect 484186 380258 484422 380494
rect 484186 373258 484422 373494
rect 484186 366258 484422 366494
rect 484186 359258 484422 359494
rect 484186 352258 484422 352494
rect 484186 345258 484422 345494
rect 484186 338258 484422 338494
rect 484186 331258 484422 331494
rect 484186 324258 484422 324494
rect 484186 317258 484422 317494
rect 484186 310258 484422 310494
rect 484186 303258 484422 303494
rect 484186 296258 484422 296494
rect 484186 289258 484422 289494
rect 484186 282258 484422 282494
rect 484186 275258 484422 275494
rect 484186 268258 484422 268494
rect 484186 261258 484422 261494
rect 484186 254258 484422 254494
rect 484186 247258 484422 247494
rect 484186 240258 484422 240494
rect 484186 233258 484422 233494
rect 484186 226258 484422 226494
rect 484186 219258 484422 219494
rect 484186 212258 484422 212494
rect 484186 205258 484422 205494
rect 484186 198258 484422 198494
rect 484186 191258 484422 191494
rect 484186 184258 484422 184494
rect 484186 177258 484422 177494
rect 484186 170258 484422 170494
rect 484186 163258 484422 163494
rect 484186 156258 484422 156494
rect 484186 149258 484422 149494
rect 484186 142258 484422 142494
rect 484186 135258 484422 135494
rect 484186 128258 484422 128494
rect 484186 121258 484422 121494
rect 484186 114258 484422 114494
rect 484186 107258 484422 107494
rect 484186 100258 484422 100494
rect 484186 93258 484422 93494
rect 484186 86258 484422 86494
rect 484186 79258 484422 79494
rect 484186 72258 484422 72494
rect 484186 65258 484422 65494
rect 484186 58258 484422 58494
rect 484186 51258 484422 51494
rect 484186 44258 484422 44494
rect 484186 37258 484422 37494
rect 484186 30258 484422 30494
rect 484186 23258 484422 23494
rect 484186 16258 484422 16494
rect 484186 9258 484422 9494
rect 484186 2258 484422 2494
rect 484186 -982 484422 -746
rect 484186 -1302 484422 -1066
rect 485918 705962 486154 706198
rect 485918 705642 486154 705878
rect 485918 696325 486154 696561
rect 485918 689325 486154 689561
rect 485918 682325 486154 682561
rect 485918 675325 486154 675561
rect 485918 668325 486154 668561
rect 485918 661325 486154 661561
rect 485918 654325 486154 654561
rect 485918 647325 486154 647561
rect 485918 640325 486154 640561
rect 485918 633325 486154 633561
rect 485918 626325 486154 626561
rect 485918 619325 486154 619561
rect 485918 612325 486154 612561
rect 485918 605325 486154 605561
rect 485918 598325 486154 598561
rect 485918 591325 486154 591561
rect 485918 584325 486154 584561
rect 485918 577325 486154 577561
rect 485918 570325 486154 570561
rect 485918 563325 486154 563561
rect 485918 556325 486154 556561
rect 485918 549325 486154 549561
rect 485918 542325 486154 542561
rect 485918 535325 486154 535561
rect 485918 528325 486154 528561
rect 485918 521325 486154 521561
rect 485918 514325 486154 514561
rect 485918 507325 486154 507561
rect 485918 500325 486154 500561
rect 485918 493325 486154 493561
rect 485918 486325 486154 486561
rect 485918 479325 486154 479561
rect 485918 472325 486154 472561
rect 485918 465325 486154 465561
rect 485918 458325 486154 458561
rect 485918 451325 486154 451561
rect 485918 444325 486154 444561
rect 485918 437325 486154 437561
rect 485918 430325 486154 430561
rect 485918 423325 486154 423561
rect 485918 416325 486154 416561
rect 485918 409325 486154 409561
rect 485918 402325 486154 402561
rect 485918 395325 486154 395561
rect 485918 388325 486154 388561
rect 485918 381325 486154 381561
rect 485918 374325 486154 374561
rect 485918 367325 486154 367561
rect 485918 360325 486154 360561
rect 485918 353325 486154 353561
rect 485918 346325 486154 346561
rect 485918 339325 486154 339561
rect 485918 332325 486154 332561
rect 485918 325325 486154 325561
rect 485918 318325 486154 318561
rect 485918 311325 486154 311561
rect 485918 304325 486154 304561
rect 485918 297325 486154 297561
rect 485918 290325 486154 290561
rect 485918 283325 486154 283561
rect 485918 276325 486154 276561
rect 485918 269325 486154 269561
rect 485918 262325 486154 262561
rect 485918 255325 486154 255561
rect 485918 248325 486154 248561
rect 485918 241325 486154 241561
rect 485918 234325 486154 234561
rect 485918 227325 486154 227561
rect 485918 220325 486154 220561
rect 485918 213325 486154 213561
rect 485918 206325 486154 206561
rect 485918 199325 486154 199561
rect 485918 192325 486154 192561
rect 485918 185325 486154 185561
rect 485918 178325 486154 178561
rect 485918 171325 486154 171561
rect 485918 164325 486154 164561
rect 485918 157325 486154 157561
rect 485918 150325 486154 150561
rect 485918 143325 486154 143561
rect 485918 136325 486154 136561
rect 485918 129325 486154 129561
rect 485918 122325 486154 122561
rect 485918 115325 486154 115561
rect 485918 108325 486154 108561
rect 485918 101325 486154 101561
rect 485918 94325 486154 94561
rect 485918 87325 486154 87561
rect 485918 80325 486154 80561
rect 485918 73325 486154 73561
rect 485918 66325 486154 66561
rect 485918 59325 486154 59561
rect 485918 52325 486154 52561
rect 485918 45325 486154 45561
rect 485918 38325 486154 38561
rect 485918 31325 486154 31561
rect 485918 24325 486154 24561
rect 485918 17325 486154 17561
rect 485918 10325 486154 10561
rect 485918 3325 486154 3561
rect 485918 -1942 486154 -1706
rect 485918 -2262 486154 -2026
rect 491186 705002 491422 705238
rect 491186 704682 491422 704918
rect 491186 695258 491422 695494
rect 491186 688258 491422 688494
rect 491186 681258 491422 681494
rect 491186 674258 491422 674494
rect 491186 667258 491422 667494
rect 491186 660258 491422 660494
rect 491186 653258 491422 653494
rect 491186 646258 491422 646494
rect 491186 639258 491422 639494
rect 491186 632258 491422 632494
rect 491186 625258 491422 625494
rect 491186 618258 491422 618494
rect 491186 611258 491422 611494
rect 491186 604258 491422 604494
rect 491186 597258 491422 597494
rect 491186 590258 491422 590494
rect 491186 583258 491422 583494
rect 491186 576258 491422 576494
rect 491186 569258 491422 569494
rect 491186 562258 491422 562494
rect 491186 555258 491422 555494
rect 491186 548258 491422 548494
rect 491186 541258 491422 541494
rect 491186 534258 491422 534494
rect 491186 527258 491422 527494
rect 491186 520258 491422 520494
rect 491186 513258 491422 513494
rect 491186 506258 491422 506494
rect 491186 499258 491422 499494
rect 491186 492258 491422 492494
rect 491186 485258 491422 485494
rect 491186 478258 491422 478494
rect 491186 471258 491422 471494
rect 491186 464258 491422 464494
rect 491186 457258 491422 457494
rect 491186 450258 491422 450494
rect 491186 443258 491422 443494
rect 491186 436258 491422 436494
rect 491186 429258 491422 429494
rect 491186 422258 491422 422494
rect 491186 415258 491422 415494
rect 491186 408258 491422 408494
rect 491186 401258 491422 401494
rect 491186 394258 491422 394494
rect 491186 387258 491422 387494
rect 491186 380258 491422 380494
rect 491186 373258 491422 373494
rect 491186 366258 491422 366494
rect 491186 359258 491422 359494
rect 491186 352258 491422 352494
rect 491186 345258 491422 345494
rect 491186 338258 491422 338494
rect 491186 331258 491422 331494
rect 491186 324258 491422 324494
rect 491186 317258 491422 317494
rect 491186 310258 491422 310494
rect 491186 303258 491422 303494
rect 491186 296258 491422 296494
rect 491186 289258 491422 289494
rect 491186 282258 491422 282494
rect 491186 275258 491422 275494
rect 491186 268258 491422 268494
rect 491186 261258 491422 261494
rect 491186 254258 491422 254494
rect 491186 247258 491422 247494
rect 491186 240258 491422 240494
rect 491186 233258 491422 233494
rect 491186 226258 491422 226494
rect 491186 219258 491422 219494
rect 491186 212258 491422 212494
rect 491186 205258 491422 205494
rect 491186 198258 491422 198494
rect 491186 191258 491422 191494
rect 491186 184258 491422 184494
rect 491186 177258 491422 177494
rect 491186 170258 491422 170494
rect 491186 163258 491422 163494
rect 491186 156258 491422 156494
rect 491186 149258 491422 149494
rect 491186 142258 491422 142494
rect 491186 135258 491422 135494
rect 491186 128258 491422 128494
rect 491186 121258 491422 121494
rect 491186 114258 491422 114494
rect 491186 107258 491422 107494
rect 491186 100258 491422 100494
rect 491186 93258 491422 93494
rect 491186 86258 491422 86494
rect 491186 79258 491422 79494
rect 491186 72258 491422 72494
rect 491186 65258 491422 65494
rect 491186 58258 491422 58494
rect 491186 51258 491422 51494
rect 491186 44258 491422 44494
rect 491186 37258 491422 37494
rect 491186 30258 491422 30494
rect 491186 23258 491422 23494
rect 491186 16258 491422 16494
rect 491186 9258 491422 9494
rect 491186 2258 491422 2494
rect 491186 -982 491422 -746
rect 491186 -1302 491422 -1066
rect 492918 705962 493154 706198
rect 492918 705642 493154 705878
rect 492918 696325 493154 696561
rect 492918 689325 493154 689561
rect 492918 682325 493154 682561
rect 492918 675325 493154 675561
rect 492918 668325 493154 668561
rect 492918 661325 493154 661561
rect 492918 654325 493154 654561
rect 492918 647325 493154 647561
rect 492918 640325 493154 640561
rect 492918 633325 493154 633561
rect 492918 626325 493154 626561
rect 492918 619325 493154 619561
rect 492918 612325 493154 612561
rect 492918 605325 493154 605561
rect 492918 598325 493154 598561
rect 492918 591325 493154 591561
rect 492918 584325 493154 584561
rect 492918 577325 493154 577561
rect 492918 570325 493154 570561
rect 492918 563325 493154 563561
rect 492918 556325 493154 556561
rect 492918 549325 493154 549561
rect 492918 542325 493154 542561
rect 492918 535325 493154 535561
rect 492918 528325 493154 528561
rect 492918 521325 493154 521561
rect 492918 514325 493154 514561
rect 492918 507325 493154 507561
rect 492918 500325 493154 500561
rect 492918 493325 493154 493561
rect 492918 486325 493154 486561
rect 492918 479325 493154 479561
rect 492918 472325 493154 472561
rect 492918 465325 493154 465561
rect 492918 458325 493154 458561
rect 492918 451325 493154 451561
rect 492918 444325 493154 444561
rect 492918 437325 493154 437561
rect 492918 430325 493154 430561
rect 492918 423325 493154 423561
rect 492918 416325 493154 416561
rect 492918 409325 493154 409561
rect 492918 402325 493154 402561
rect 492918 395325 493154 395561
rect 492918 388325 493154 388561
rect 492918 381325 493154 381561
rect 492918 374325 493154 374561
rect 492918 367325 493154 367561
rect 492918 360325 493154 360561
rect 492918 353325 493154 353561
rect 492918 346325 493154 346561
rect 492918 339325 493154 339561
rect 492918 332325 493154 332561
rect 492918 325325 493154 325561
rect 492918 318325 493154 318561
rect 492918 311325 493154 311561
rect 492918 304325 493154 304561
rect 492918 297325 493154 297561
rect 492918 290325 493154 290561
rect 492918 283325 493154 283561
rect 492918 276325 493154 276561
rect 492918 269325 493154 269561
rect 492918 262325 493154 262561
rect 492918 255325 493154 255561
rect 492918 248325 493154 248561
rect 492918 241325 493154 241561
rect 492918 234325 493154 234561
rect 492918 227325 493154 227561
rect 492918 220325 493154 220561
rect 492918 213325 493154 213561
rect 492918 206325 493154 206561
rect 492918 199325 493154 199561
rect 492918 192325 493154 192561
rect 492918 185325 493154 185561
rect 492918 178325 493154 178561
rect 492918 171325 493154 171561
rect 492918 164325 493154 164561
rect 492918 157325 493154 157561
rect 492918 150325 493154 150561
rect 492918 143325 493154 143561
rect 492918 136325 493154 136561
rect 492918 129325 493154 129561
rect 492918 122325 493154 122561
rect 492918 115325 493154 115561
rect 492918 108325 493154 108561
rect 492918 101325 493154 101561
rect 492918 94325 493154 94561
rect 492918 87325 493154 87561
rect 492918 80325 493154 80561
rect 492918 73325 493154 73561
rect 492918 66325 493154 66561
rect 492918 59325 493154 59561
rect 492918 52325 493154 52561
rect 492918 45325 493154 45561
rect 492918 38325 493154 38561
rect 492918 31325 493154 31561
rect 492918 24325 493154 24561
rect 492918 17325 493154 17561
rect 492918 10325 493154 10561
rect 492918 3325 493154 3561
rect 492918 -1942 493154 -1706
rect 492918 -2262 493154 -2026
rect 498186 705002 498422 705238
rect 498186 704682 498422 704918
rect 498186 695258 498422 695494
rect 498186 688258 498422 688494
rect 498186 681258 498422 681494
rect 498186 674258 498422 674494
rect 498186 667258 498422 667494
rect 498186 660258 498422 660494
rect 498186 653258 498422 653494
rect 498186 646258 498422 646494
rect 498186 639258 498422 639494
rect 498186 632258 498422 632494
rect 498186 625258 498422 625494
rect 498186 618258 498422 618494
rect 498186 611258 498422 611494
rect 498186 604258 498422 604494
rect 498186 597258 498422 597494
rect 498186 590258 498422 590494
rect 498186 583258 498422 583494
rect 498186 576258 498422 576494
rect 498186 569258 498422 569494
rect 498186 562258 498422 562494
rect 498186 555258 498422 555494
rect 498186 548258 498422 548494
rect 498186 541258 498422 541494
rect 498186 534258 498422 534494
rect 498186 527258 498422 527494
rect 498186 520258 498422 520494
rect 498186 513258 498422 513494
rect 498186 506258 498422 506494
rect 498186 499258 498422 499494
rect 498186 492258 498422 492494
rect 498186 485258 498422 485494
rect 498186 478258 498422 478494
rect 498186 471258 498422 471494
rect 498186 464258 498422 464494
rect 498186 457258 498422 457494
rect 498186 450258 498422 450494
rect 498186 443258 498422 443494
rect 498186 436258 498422 436494
rect 498186 429258 498422 429494
rect 498186 422258 498422 422494
rect 498186 415258 498422 415494
rect 498186 408258 498422 408494
rect 498186 401258 498422 401494
rect 498186 394258 498422 394494
rect 498186 387258 498422 387494
rect 498186 380258 498422 380494
rect 498186 373258 498422 373494
rect 498186 366258 498422 366494
rect 498186 359258 498422 359494
rect 498186 352258 498422 352494
rect 498186 345258 498422 345494
rect 498186 338258 498422 338494
rect 498186 331258 498422 331494
rect 498186 324258 498422 324494
rect 498186 317258 498422 317494
rect 498186 310258 498422 310494
rect 498186 303258 498422 303494
rect 498186 296258 498422 296494
rect 498186 289258 498422 289494
rect 498186 282258 498422 282494
rect 498186 275258 498422 275494
rect 498186 268258 498422 268494
rect 498186 261258 498422 261494
rect 498186 254258 498422 254494
rect 498186 247258 498422 247494
rect 498186 240258 498422 240494
rect 498186 233258 498422 233494
rect 498186 226258 498422 226494
rect 498186 219258 498422 219494
rect 498186 212258 498422 212494
rect 498186 205258 498422 205494
rect 498186 198258 498422 198494
rect 498186 191258 498422 191494
rect 498186 184258 498422 184494
rect 498186 177258 498422 177494
rect 498186 170258 498422 170494
rect 498186 163258 498422 163494
rect 498186 156258 498422 156494
rect 498186 149258 498422 149494
rect 498186 142258 498422 142494
rect 498186 135258 498422 135494
rect 498186 128258 498422 128494
rect 498186 121258 498422 121494
rect 498186 114258 498422 114494
rect 498186 107258 498422 107494
rect 498186 100258 498422 100494
rect 498186 93258 498422 93494
rect 498186 86258 498422 86494
rect 498186 79258 498422 79494
rect 498186 72258 498422 72494
rect 498186 65258 498422 65494
rect 498186 58258 498422 58494
rect 498186 51258 498422 51494
rect 498186 44258 498422 44494
rect 498186 37258 498422 37494
rect 498186 30258 498422 30494
rect 498186 23258 498422 23494
rect 498186 16258 498422 16494
rect 498186 9258 498422 9494
rect 498186 2258 498422 2494
rect 498186 -982 498422 -746
rect 498186 -1302 498422 -1066
rect 499918 705962 500154 706198
rect 499918 705642 500154 705878
rect 499918 696325 500154 696561
rect 499918 689325 500154 689561
rect 499918 682325 500154 682561
rect 499918 675325 500154 675561
rect 499918 668325 500154 668561
rect 499918 661325 500154 661561
rect 499918 654325 500154 654561
rect 499918 647325 500154 647561
rect 499918 640325 500154 640561
rect 499918 633325 500154 633561
rect 499918 626325 500154 626561
rect 499918 619325 500154 619561
rect 499918 612325 500154 612561
rect 499918 605325 500154 605561
rect 499918 598325 500154 598561
rect 499918 591325 500154 591561
rect 499918 584325 500154 584561
rect 499918 577325 500154 577561
rect 499918 570325 500154 570561
rect 499918 563325 500154 563561
rect 499918 556325 500154 556561
rect 499918 549325 500154 549561
rect 499918 542325 500154 542561
rect 499918 535325 500154 535561
rect 499918 528325 500154 528561
rect 499918 521325 500154 521561
rect 499918 514325 500154 514561
rect 499918 507325 500154 507561
rect 499918 500325 500154 500561
rect 499918 493325 500154 493561
rect 499918 486325 500154 486561
rect 499918 479325 500154 479561
rect 499918 472325 500154 472561
rect 499918 465325 500154 465561
rect 499918 458325 500154 458561
rect 499918 451325 500154 451561
rect 499918 444325 500154 444561
rect 499918 437325 500154 437561
rect 499918 430325 500154 430561
rect 499918 423325 500154 423561
rect 499918 416325 500154 416561
rect 499918 409325 500154 409561
rect 499918 402325 500154 402561
rect 499918 395325 500154 395561
rect 499918 388325 500154 388561
rect 499918 381325 500154 381561
rect 499918 374325 500154 374561
rect 499918 367325 500154 367561
rect 499918 360325 500154 360561
rect 499918 353325 500154 353561
rect 499918 346325 500154 346561
rect 499918 339325 500154 339561
rect 499918 332325 500154 332561
rect 499918 325325 500154 325561
rect 499918 318325 500154 318561
rect 499918 311325 500154 311561
rect 499918 304325 500154 304561
rect 499918 297325 500154 297561
rect 499918 290325 500154 290561
rect 499918 283325 500154 283561
rect 499918 276325 500154 276561
rect 499918 269325 500154 269561
rect 499918 262325 500154 262561
rect 499918 255325 500154 255561
rect 499918 248325 500154 248561
rect 499918 241325 500154 241561
rect 499918 234325 500154 234561
rect 499918 227325 500154 227561
rect 499918 220325 500154 220561
rect 499918 213325 500154 213561
rect 499918 206325 500154 206561
rect 499918 199325 500154 199561
rect 499918 192325 500154 192561
rect 499918 185325 500154 185561
rect 499918 178325 500154 178561
rect 499918 171325 500154 171561
rect 499918 164325 500154 164561
rect 499918 157325 500154 157561
rect 499918 150325 500154 150561
rect 499918 143325 500154 143561
rect 499918 136325 500154 136561
rect 499918 129325 500154 129561
rect 499918 122325 500154 122561
rect 499918 115325 500154 115561
rect 499918 108325 500154 108561
rect 499918 101325 500154 101561
rect 499918 94325 500154 94561
rect 499918 87325 500154 87561
rect 499918 80325 500154 80561
rect 499918 73325 500154 73561
rect 499918 66325 500154 66561
rect 499918 59325 500154 59561
rect 499918 52325 500154 52561
rect 499918 45325 500154 45561
rect 499918 38325 500154 38561
rect 499918 31325 500154 31561
rect 499918 24325 500154 24561
rect 499918 17325 500154 17561
rect 499918 10325 500154 10561
rect 499918 3325 500154 3561
rect 499918 -1942 500154 -1706
rect 499918 -2262 500154 -2026
rect 505186 705002 505422 705238
rect 505186 704682 505422 704918
rect 505186 695258 505422 695494
rect 505186 688258 505422 688494
rect 505186 681258 505422 681494
rect 505186 674258 505422 674494
rect 505186 667258 505422 667494
rect 505186 660258 505422 660494
rect 505186 653258 505422 653494
rect 505186 646258 505422 646494
rect 505186 639258 505422 639494
rect 505186 632258 505422 632494
rect 505186 625258 505422 625494
rect 505186 618258 505422 618494
rect 505186 611258 505422 611494
rect 505186 604258 505422 604494
rect 505186 597258 505422 597494
rect 505186 590258 505422 590494
rect 505186 583258 505422 583494
rect 505186 576258 505422 576494
rect 505186 569258 505422 569494
rect 505186 562258 505422 562494
rect 505186 555258 505422 555494
rect 505186 548258 505422 548494
rect 505186 541258 505422 541494
rect 505186 534258 505422 534494
rect 505186 527258 505422 527494
rect 505186 520258 505422 520494
rect 505186 513258 505422 513494
rect 505186 506258 505422 506494
rect 505186 499258 505422 499494
rect 505186 492258 505422 492494
rect 505186 485258 505422 485494
rect 505186 478258 505422 478494
rect 505186 471258 505422 471494
rect 505186 464258 505422 464494
rect 505186 457258 505422 457494
rect 505186 450258 505422 450494
rect 505186 443258 505422 443494
rect 505186 436258 505422 436494
rect 505186 429258 505422 429494
rect 505186 422258 505422 422494
rect 505186 415258 505422 415494
rect 505186 408258 505422 408494
rect 505186 401258 505422 401494
rect 505186 394258 505422 394494
rect 505186 387258 505422 387494
rect 505186 380258 505422 380494
rect 505186 373258 505422 373494
rect 505186 366258 505422 366494
rect 505186 359258 505422 359494
rect 505186 352258 505422 352494
rect 505186 345258 505422 345494
rect 505186 338258 505422 338494
rect 505186 331258 505422 331494
rect 505186 324258 505422 324494
rect 505186 317258 505422 317494
rect 505186 310258 505422 310494
rect 505186 303258 505422 303494
rect 505186 296258 505422 296494
rect 505186 289258 505422 289494
rect 505186 282258 505422 282494
rect 505186 275258 505422 275494
rect 505186 268258 505422 268494
rect 505186 261258 505422 261494
rect 505186 254258 505422 254494
rect 505186 247258 505422 247494
rect 505186 240258 505422 240494
rect 505186 233258 505422 233494
rect 505186 226258 505422 226494
rect 505186 219258 505422 219494
rect 505186 212258 505422 212494
rect 505186 205258 505422 205494
rect 505186 198258 505422 198494
rect 505186 191258 505422 191494
rect 505186 184258 505422 184494
rect 505186 177258 505422 177494
rect 505186 170258 505422 170494
rect 505186 163258 505422 163494
rect 505186 156258 505422 156494
rect 505186 149258 505422 149494
rect 505186 142258 505422 142494
rect 505186 135258 505422 135494
rect 505186 128258 505422 128494
rect 505186 121258 505422 121494
rect 505186 114258 505422 114494
rect 505186 107258 505422 107494
rect 505186 100258 505422 100494
rect 505186 93258 505422 93494
rect 505186 86258 505422 86494
rect 505186 79258 505422 79494
rect 505186 72258 505422 72494
rect 505186 65258 505422 65494
rect 505186 58258 505422 58494
rect 505186 51258 505422 51494
rect 505186 44258 505422 44494
rect 505186 37258 505422 37494
rect 505186 30258 505422 30494
rect 505186 23258 505422 23494
rect 505186 16258 505422 16494
rect 505186 9258 505422 9494
rect 505186 2258 505422 2494
rect 505186 -982 505422 -746
rect 505186 -1302 505422 -1066
rect 506918 705962 507154 706198
rect 506918 705642 507154 705878
rect 506918 696325 507154 696561
rect 506918 689325 507154 689561
rect 506918 682325 507154 682561
rect 506918 675325 507154 675561
rect 506918 668325 507154 668561
rect 506918 661325 507154 661561
rect 506918 654325 507154 654561
rect 506918 647325 507154 647561
rect 506918 640325 507154 640561
rect 506918 633325 507154 633561
rect 506918 626325 507154 626561
rect 506918 619325 507154 619561
rect 506918 612325 507154 612561
rect 506918 605325 507154 605561
rect 506918 598325 507154 598561
rect 506918 591325 507154 591561
rect 506918 584325 507154 584561
rect 506918 577325 507154 577561
rect 506918 570325 507154 570561
rect 506918 563325 507154 563561
rect 506918 556325 507154 556561
rect 506918 549325 507154 549561
rect 506918 542325 507154 542561
rect 506918 535325 507154 535561
rect 506918 528325 507154 528561
rect 506918 521325 507154 521561
rect 506918 514325 507154 514561
rect 506918 507325 507154 507561
rect 506918 500325 507154 500561
rect 506918 493325 507154 493561
rect 506918 486325 507154 486561
rect 506918 479325 507154 479561
rect 506918 472325 507154 472561
rect 506918 465325 507154 465561
rect 506918 458325 507154 458561
rect 506918 451325 507154 451561
rect 506918 444325 507154 444561
rect 506918 437325 507154 437561
rect 506918 430325 507154 430561
rect 506918 423325 507154 423561
rect 506918 416325 507154 416561
rect 506918 409325 507154 409561
rect 506918 402325 507154 402561
rect 506918 395325 507154 395561
rect 506918 388325 507154 388561
rect 506918 381325 507154 381561
rect 506918 374325 507154 374561
rect 506918 367325 507154 367561
rect 506918 360325 507154 360561
rect 506918 353325 507154 353561
rect 506918 346325 507154 346561
rect 506918 339325 507154 339561
rect 506918 332325 507154 332561
rect 506918 325325 507154 325561
rect 506918 318325 507154 318561
rect 506918 311325 507154 311561
rect 506918 304325 507154 304561
rect 506918 297325 507154 297561
rect 506918 290325 507154 290561
rect 506918 283325 507154 283561
rect 506918 276325 507154 276561
rect 506918 269325 507154 269561
rect 506918 262325 507154 262561
rect 506918 255325 507154 255561
rect 506918 248325 507154 248561
rect 506918 241325 507154 241561
rect 506918 234325 507154 234561
rect 506918 227325 507154 227561
rect 506918 220325 507154 220561
rect 506918 213325 507154 213561
rect 506918 206325 507154 206561
rect 506918 199325 507154 199561
rect 506918 192325 507154 192561
rect 506918 185325 507154 185561
rect 506918 178325 507154 178561
rect 506918 171325 507154 171561
rect 506918 164325 507154 164561
rect 506918 157325 507154 157561
rect 506918 150325 507154 150561
rect 506918 143325 507154 143561
rect 506918 136325 507154 136561
rect 506918 129325 507154 129561
rect 506918 122325 507154 122561
rect 506918 115325 507154 115561
rect 506918 108325 507154 108561
rect 506918 101325 507154 101561
rect 506918 94325 507154 94561
rect 506918 87325 507154 87561
rect 506918 80325 507154 80561
rect 506918 73325 507154 73561
rect 506918 66325 507154 66561
rect 506918 59325 507154 59561
rect 506918 52325 507154 52561
rect 506918 45325 507154 45561
rect 506918 38325 507154 38561
rect 506918 31325 507154 31561
rect 506918 24325 507154 24561
rect 506918 17325 507154 17561
rect 506918 10325 507154 10561
rect 506918 3325 507154 3561
rect 506918 -1942 507154 -1706
rect 506918 -2262 507154 -2026
rect 512186 705002 512422 705238
rect 512186 704682 512422 704918
rect 512186 695258 512422 695494
rect 512186 688258 512422 688494
rect 512186 681258 512422 681494
rect 512186 674258 512422 674494
rect 512186 667258 512422 667494
rect 512186 660258 512422 660494
rect 512186 653258 512422 653494
rect 512186 646258 512422 646494
rect 512186 639258 512422 639494
rect 512186 632258 512422 632494
rect 512186 625258 512422 625494
rect 512186 618258 512422 618494
rect 512186 611258 512422 611494
rect 512186 604258 512422 604494
rect 512186 597258 512422 597494
rect 512186 590258 512422 590494
rect 512186 583258 512422 583494
rect 512186 576258 512422 576494
rect 512186 569258 512422 569494
rect 512186 562258 512422 562494
rect 512186 555258 512422 555494
rect 512186 548258 512422 548494
rect 512186 541258 512422 541494
rect 512186 534258 512422 534494
rect 512186 527258 512422 527494
rect 512186 520258 512422 520494
rect 512186 513258 512422 513494
rect 512186 506258 512422 506494
rect 512186 499258 512422 499494
rect 512186 492258 512422 492494
rect 512186 485258 512422 485494
rect 512186 478258 512422 478494
rect 512186 471258 512422 471494
rect 512186 464258 512422 464494
rect 512186 457258 512422 457494
rect 512186 450258 512422 450494
rect 512186 443258 512422 443494
rect 512186 436258 512422 436494
rect 512186 429258 512422 429494
rect 512186 422258 512422 422494
rect 512186 415258 512422 415494
rect 512186 408258 512422 408494
rect 512186 401258 512422 401494
rect 512186 394258 512422 394494
rect 512186 387258 512422 387494
rect 512186 380258 512422 380494
rect 512186 373258 512422 373494
rect 512186 366258 512422 366494
rect 512186 359258 512422 359494
rect 512186 352258 512422 352494
rect 512186 345258 512422 345494
rect 512186 338258 512422 338494
rect 512186 331258 512422 331494
rect 512186 324258 512422 324494
rect 512186 317258 512422 317494
rect 512186 310258 512422 310494
rect 512186 303258 512422 303494
rect 512186 296258 512422 296494
rect 512186 289258 512422 289494
rect 512186 282258 512422 282494
rect 512186 275258 512422 275494
rect 512186 268258 512422 268494
rect 512186 261258 512422 261494
rect 512186 254258 512422 254494
rect 512186 247258 512422 247494
rect 512186 240258 512422 240494
rect 512186 233258 512422 233494
rect 512186 226258 512422 226494
rect 512186 219258 512422 219494
rect 512186 212258 512422 212494
rect 512186 205258 512422 205494
rect 512186 198258 512422 198494
rect 512186 191258 512422 191494
rect 512186 184258 512422 184494
rect 512186 177258 512422 177494
rect 512186 170258 512422 170494
rect 512186 163258 512422 163494
rect 512186 156258 512422 156494
rect 512186 149258 512422 149494
rect 512186 142258 512422 142494
rect 512186 135258 512422 135494
rect 512186 128258 512422 128494
rect 512186 121258 512422 121494
rect 512186 114258 512422 114494
rect 512186 107258 512422 107494
rect 512186 100258 512422 100494
rect 512186 93258 512422 93494
rect 512186 86258 512422 86494
rect 512186 79258 512422 79494
rect 512186 72258 512422 72494
rect 512186 65258 512422 65494
rect 512186 58258 512422 58494
rect 512186 51258 512422 51494
rect 512186 44258 512422 44494
rect 512186 37258 512422 37494
rect 512186 30258 512422 30494
rect 512186 23258 512422 23494
rect 512186 16258 512422 16494
rect 512186 9258 512422 9494
rect 512186 2258 512422 2494
rect 512186 -982 512422 -746
rect 512186 -1302 512422 -1066
rect 513918 705962 514154 706198
rect 513918 705642 514154 705878
rect 513918 696325 514154 696561
rect 513918 689325 514154 689561
rect 513918 682325 514154 682561
rect 513918 675325 514154 675561
rect 513918 668325 514154 668561
rect 513918 661325 514154 661561
rect 513918 654325 514154 654561
rect 513918 647325 514154 647561
rect 513918 640325 514154 640561
rect 513918 633325 514154 633561
rect 513918 626325 514154 626561
rect 513918 619325 514154 619561
rect 513918 612325 514154 612561
rect 513918 605325 514154 605561
rect 513918 598325 514154 598561
rect 513918 591325 514154 591561
rect 513918 584325 514154 584561
rect 513918 577325 514154 577561
rect 513918 570325 514154 570561
rect 513918 563325 514154 563561
rect 513918 556325 514154 556561
rect 513918 549325 514154 549561
rect 513918 542325 514154 542561
rect 513918 535325 514154 535561
rect 513918 528325 514154 528561
rect 513918 521325 514154 521561
rect 513918 514325 514154 514561
rect 513918 507325 514154 507561
rect 513918 500325 514154 500561
rect 513918 493325 514154 493561
rect 513918 486325 514154 486561
rect 513918 479325 514154 479561
rect 513918 472325 514154 472561
rect 513918 465325 514154 465561
rect 513918 458325 514154 458561
rect 513918 451325 514154 451561
rect 513918 444325 514154 444561
rect 513918 437325 514154 437561
rect 513918 430325 514154 430561
rect 513918 423325 514154 423561
rect 513918 416325 514154 416561
rect 513918 409325 514154 409561
rect 513918 402325 514154 402561
rect 513918 395325 514154 395561
rect 513918 388325 514154 388561
rect 513918 381325 514154 381561
rect 513918 374325 514154 374561
rect 513918 367325 514154 367561
rect 513918 360325 514154 360561
rect 513918 353325 514154 353561
rect 513918 346325 514154 346561
rect 513918 339325 514154 339561
rect 513918 332325 514154 332561
rect 513918 325325 514154 325561
rect 513918 318325 514154 318561
rect 513918 311325 514154 311561
rect 513918 304325 514154 304561
rect 513918 297325 514154 297561
rect 513918 290325 514154 290561
rect 513918 283325 514154 283561
rect 513918 276325 514154 276561
rect 513918 269325 514154 269561
rect 513918 262325 514154 262561
rect 513918 255325 514154 255561
rect 513918 248325 514154 248561
rect 513918 241325 514154 241561
rect 513918 234325 514154 234561
rect 513918 227325 514154 227561
rect 513918 220325 514154 220561
rect 513918 213325 514154 213561
rect 513918 206325 514154 206561
rect 513918 199325 514154 199561
rect 513918 192325 514154 192561
rect 513918 185325 514154 185561
rect 513918 178325 514154 178561
rect 513918 171325 514154 171561
rect 513918 164325 514154 164561
rect 513918 157325 514154 157561
rect 513918 150325 514154 150561
rect 513918 143325 514154 143561
rect 513918 136325 514154 136561
rect 513918 129325 514154 129561
rect 513918 122325 514154 122561
rect 513918 115325 514154 115561
rect 513918 108325 514154 108561
rect 513918 101325 514154 101561
rect 513918 94325 514154 94561
rect 513918 87325 514154 87561
rect 513918 80325 514154 80561
rect 513918 73325 514154 73561
rect 513918 66325 514154 66561
rect 513918 59325 514154 59561
rect 513918 52325 514154 52561
rect 513918 45325 514154 45561
rect 513918 38325 514154 38561
rect 513918 31325 514154 31561
rect 513918 24325 514154 24561
rect 513918 17325 514154 17561
rect 513918 10325 514154 10561
rect 513918 3325 514154 3561
rect 513918 -1942 514154 -1706
rect 513918 -2262 514154 -2026
rect 519186 705002 519422 705238
rect 519186 704682 519422 704918
rect 519186 695258 519422 695494
rect 519186 688258 519422 688494
rect 519186 681258 519422 681494
rect 519186 674258 519422 674494
rect 519186 667258 519422 667494
rect 519186 660258 519422 660494
rect 519186 653258 519422 653494
rect 519186 646258 519422 646494
rect 519186 639258 519422 639494
rect 519186 632258 519422 632494
rect 519186 625258 519422 625494
rect 519186 618258 519422 618494
rect 519186 611258 519422 611494
rect 519186 604258 519422 604494
rect 519186 597258 519422 597494
rect 519186 590258 519422 590494
rect 519186 583258 519422 583494
rect 519186 576258 519422 576494
rect 519186 569258 519422 569494
rect 519186 562258 519422 562494
rect 519186 555258 519422 555494
rect 519186 548258 519422 548494
rect 519186 541258 519422 541494
rect 519186 534258 519422 534494
rect 519186 527258 519422 527494
rect 519186 520258 519422 520494
rect 519186 513258 519422 513494
rect 519186 506258 519422 506494
rect 519186 499258 519422 499494
rect 519186 492258 519422 492494
rect 519186 485258 519422 485494
rect 519186 478258 519422 478494
rect 519186 471258 519422 471494
rect 519186 464258 519422 464494
rect 519186 457258 519422 457494
rect 519186 450258 519422 450494
rect 519186 443258 519422 443494
rect 519186 436258 519422 436494
rect 519186 429258 519422 429494
rect 519186 422258 519422 422494
rect 520918 705962 521154 706198
rect 520918 705642 521154 705878
rect 520918 696325 521154 696561
rect 520918 689325 521154 689561
rect 520918 682325 521154 682561
rect 520918 675325 521154 675561
rect 520918 668325 521154 668561
rect 520918 661325 521154 661561
rect 520918 654325 521154 654561
rect 520918 647325 521154 647561
rect 520918 640325 521154 640561
rect 520918 633325 521154 633561
rect 520918 626325 521154 626561
rect 520918 619325 521154 619561
rect 520918 612325 521154 612561
rect 520918 605325 521154 605561
rect 520918 598325 521154 598561
rect 520918 591325 521154 591561
rect 520918 584325 521154 584561
rect 520918 577325 521154 577561
rect 520918 570325 521154 570561
rect 520918 563325 521154 563561
rect 520918 556325 521154 556561
rect 520918 549325 521154 549561
rect 520918 542325 521154 542561
rect 520918 535325 521154 535561
rect 520918 528325 521154 528561
rect 520918 521325 521154 521561
rect 520918 514325 521154 514561
rect 520918 507325 521154 507561
rect 520918 500325 521154 500561
rect 520918 493325 521154 493561
rect 520918 486325 521154 486561
rect 520918 479325 521154 479561
rect 520918 472325 521154 472561
rect 520918 465325 521154 465561
rect 520918 458325 521154 458561
rect 520918 451325 521154 451561
rect 520918 444325 521154 444561
rect 520918 437325 521154 437561
rect 520918 430325 521154 430561
rect 520918 423325 521154 423561
rect 526186 705002 526422 705238
rect 526186 704682 526422 704918
rect 526186 695258 526422 695494
rect 526186 688258 526422 688494
rect 526186 681258 526422 681494
rect 526186 674258 526422 674494
rect 526186 667258 526422 667494
rect 526186 660258 526422 660494
rect 526186 653258 526422 653494
rect 526186 646258 526422 646494
rect 526186 639258 526422 639494
rect 526186 632258 526422 632494
rect 526186 625258 526422 625494
rect 526186 618258 526422 618494
rect 526186 611258 526422 611494
rect 526186 604258 526422 604494
rect 526186 597258 526422 597494
rect 526186 590258 526422 590494
rect 526186 583258 526422 583494
rect 526186 576258 526422 576494
rect 526186 569258 526422 569494
rect 526186 562258 526422 562494
rect 526186 555258 526422 555494
rect 526186 548258 526422 548494
rect 526186 541258 526422 541494
rect 526186 534258 526422 534494
rect 526186 527258 526422 527494
rect 526186 520258 526422 520494
rect 526186 513258 526422 513494
rect 526186 506258 526422 506494
rect 526186 499258 526422 499494
rect 526186 492258 526422 492494
rect 526186 485258 526422 485494
rect 526186 478258 526422 478494
rect 526186 471258 526422 471494
rect 526186 464258 526422 464494
rect 526186 457258 526422 457494
rect 526186 450258 526422 450494
rect 526186 443258 526422 443494
rect 526186 436258 526422 436494
rect 526186 429258 526422 429494
rect 526186 422258 526422 422494
rect 527918 705962 528154 706198
rect 527918 705642 528154 705878
rect 527918 696325 528154 696561
rect 527918 689325 528154 689561
rect 527918 682325 528154 682561
rect 527918 675325 528154 675561
rect 527918 668325 528154 668561
rect 527918 661325 528154 661561
rect 527918 654325 528154 654561
rect 527918 647325 528154 647561
rect 527918 640325 528154 640561
rect 527918 633325 528154 633561
rect 527918 626325 528154 626561
rect 527918 619325 528154 619561
rect 527918 612325 528154 612561
rect 527918 605325 528154 605561
rect 527918 598325 528154 598561
rect 527918 591325 528154 591561
rect 527918 584325 528154 584561
rect 527918 577325 528154 577561
rect 527918 570325 528154 570561
rect 527918 563325 528154 563561
rect 527918 556325 528154 556561
rect 527918 549325 528154 549561
rect 527918 542325 528154 542561
rect 527918 535325 528154 535561
rect 527918 528325 528154 528561
rect 527918 521325 528154 521561
rect 527918 514325 528154 514561
rect 527918 507325 528154 507561
rect 527918 500325 528154 500561
rect 527918 493325 528154 493561
rect 527918 486325 528154 486561
rect 527918 479325 528154 479561
rect 527918 472325 528154 472561
rect 527918 465325 528154 465561
rect 527918 458325 528154 458561
rect 527918 451325 528154 451561
rect 527918 444325 528154 444561
rect 527918 437325 528154 437561
rect 527918 430325 528154 430561
rect 527918 423325 528154 423561
rect 520918 416325 521154 416561
rect 522850 416325 523086 416561
rect 524782 416325 525018 416561
rect 526714 416325 526950 416561
rect 527918 416325 528154 416561
rect 519186 415258 519422 415494
rect 519952 415258 520188 415494
rect 521884 415258 522120 415494
rect 523816 415258 524052 415494
rect 525748 415258 525984 415494
rect 520918 409325 521154 409561
rect 522850 409325 523086 409561
rect 524782 409325 525018 409561
rect 526714 409325 526950 409561
rect 527918 409325 528154 409561
rect 519186 408258 519422 408494
rect 519952 408258 520188 408494
rect 521884 408258 522120 408494
rect 523816 408258 524052 408494
rect 525748 408258 525984 408494
rect 520918 402325 521154 402561
rect 522850 402325 523086 402561
rect 524782 402325 525018 402561
rect 526714 402325 526950 402561
rect 527918 402325 528154 402561
rect 519186 401258 519422 401494
rect 519186 394258 519422 394494
rect 519186 387258 519422 387494
rect 520918 395325 521154 395561
rect 520918 388325 521154 388561
rect 526186 394258 526422 394494
rect 526186 387258 526422 387494
rect 527918 395325 528154 395561
rect 527918 388325 528154 388561
rect 519186 380258 519422 380494
rect 527918 381325 528154 381561
rect 520918 374325 521154 374561
rect 522850 374325 523086 374561
rect 524782 374325 525018 374561
rect 526714 374325 526950 374561
rect 527918 374325 528154 374561
rect 519186 373258 519422 373494
rect 519952 373258 520188 373494
rect 521884 373258 522120 373494
rect 523816 373258 524052 373494
rect 525748 373258 525984 373494
rect 520918 367325 521154 367561
rect 522850 367325 523086 367561
rect 524782 367325 525018 367561
rect 526714 367325 526950 367561
rect 527918 367325 528154 367561
rect 519186 366258 519422 366494
rect 519952 366258 520188 366494
rect 521884 366258 522120 366494
rect 523816 366258 524052 366494
rect 525748 366258 525984 366494
rect 527918 360325 528154 360561
rect 519186 359258 519422 359494
rect 519186 352258 519422 352494
rect 519186 345258 519422 345494
rect 520918 353325 521154 353561
rect 520918 346325 521154 346561
rect 526186 359258 526422 359494
rect 526186 352258 526422 352494
rect 526186 345258 526422 345494
rect 527918 353325 528154 353561
rect 527918 346325 528154 346561
rect 520918 339325 521154 339561
rect 522850 339325 523086 339561
rect 524782 339325 525018 339561
rect 526714 339325 526950 339561
rect 527918 339325 528154 339561
rect 519186 338258 519422 338494
rect 519952 338258 520188 338494
rect 521884 338258 522120 338494
rect 523816 338258 524052 338494
rect 525748 338258 525984 338494
rect 520918 332325 521154 332561
rect 522850 332325 523086 332561
rect 524782 332325 525018 332561
rect 526714 332325 526950 332561
rect 527918 332325 528154 332561
rect 519186 331258 519422 331494
rect 519952 331258 520188 331494
rect 521884 331258 522120 331494
rect 523816 331258 524052 331494
rect 525748 331258 525984 331494
rect 520918 325325 521154 325561
rect 522850 325325 523086 325561
rect 524782 325325 525018 325561
rect 526714 325325 526950 325561
rect 527918 325325 528154 325561
rect 519186 324258 519422 324494
rect 519952 324258 520188 324494
rect 521884 324258 522120 324494
rect 523816 324258 524052 324494
rect 525748 324258 525984 324494
rect 519186 317258 519422 317494
rect 519186 310258 519422 310494
rect 519186 303258 519422 303494
rect 520918 318325 521154 318561
rect 520918 311325 521154 311561
rect 520918 304325 521154 304561
rect 526186 317258 526422 317494
rect 526186 310258 526422 310494
rect 526186 303258 526422 303494
rect 527918 318325 528154 318561
rect 527918 311325 528154 311561
rect 527918 304325 528154 304561
rect 520918 297325 521154 297561
rect 522850 297325 523086 297561
rect 524782 297325 525018 297561
rect 526714 297325 526950 297561
rect 527918 297325 528154 297561
rect 519186 296258 519422 296494
rect 519952 296258 520188 296494
rect 521884 296258 522120 296494
rect 523816 296258 524052 296494
rect 525748 296258 525984 296494
rect 520918 290325 521154 290561
rect 522850 290325 523086 290561
rect 524782 290325 525018 290561
rect 526714 290325 526950 290561
rect 527918 290325 528154 290561
rect 519186 289258 519422 289494
rect 519952 289258 520188 289494
rect 521884 289258 522120 289494
rect 523816 289258 524052 289494
rect 525748 289258 525984 289494
rect 520918 283325 521154 283561
rect 522850 283325 523086 283561
rect 524782 283325 525018 283561
rect 526714 283325 526950 283561
rect 527918 283325 528154 283561
rect 519186 282258 519422 282494
rect 519952 282258 520188 282494
rect 521884 282258 522120 282494
rect 523816 282258 524052 282494
rect 525748 282258 525984 282494
rect 519186 275258 519422 275494
rect 519186 268258 519422 268494
rect 520918 276325 521154 276561
rect 520918 269325 521154 269561
rect 520918 262325 521154 262561
rect 526186 275258 526422 275494
rect 526186 268258 526422 268494
rect 527918 276325 528154 276561
rect 527918 269325 528154 269561
rect 527918 262325 528154 262561
rect 519186 261258 519422 261494
rect 520918 255325 521154 255561
rect 522850 255325 523086 255561
rect 524782 255325 525018 255561
rect 526714 255325 526950 255561
rect 527918 255325 528154 255561
rect 519186 254258 519422 254494
rect 519952 254258 520188 254494
rect 521884 254258 522120 254494
rect 523816 254258 524052 254494
rect 525748 254258 525984 254494
rect 520918 248325 521154 248561
rect 522850 248325 523086 248561
rect 524782 248325 525018 248561
rect 526714 248325 526950 248561
rect 527918 248325 528154 248561
rect 519186 247258 519422 247494
rect 519952 247258 520188 247494
rect 521884 247258 522120 247494
rect 523816 247258 524052 247494
rect 525748 247258 525984 247494
rect 519186 240258 519422 240494
rect 527918 241325 528154 241561
rect 519186 233258 519422 233494
rect 519186 226258 519422 226494
rect 519186 219258 519422 219494
rect 519186 212258 519422 212494
rect 519186 205258 519422 205494
rect 519186 198258 519422 198494
rect 519186 191258 519422 191494
rect 519186 184258 519422 184494
rect 519186 177258 519422 177494
rect 519186 170258 519422 170494
rect 519186 163258 519422 163494
rect 519186 156258 519422 156494
rect 519186 149258 519422 149494
rect 519186 142258 519422 142494
rect 519186 135258 519422 135494
rect 519186 128258 519422 128494
rect 519186 121258 519422 121494
rect 519186 114258 519422 114494
rect 519186 107258 519422 107494
rect 519186 100258 519422 100494
rect 519186 93258 519422 93494
rect 519186 86258 519422 86494
rect 519186 79258 519422 79494
rect 519186 72258 519422 72494
rect 519186 65258 519422 65494
rect 519186 58258 519422 58494
rect 519186 51258 519422 51494
rect 519186 44258 519422 44494
rect 519186 37258 519422 37494
rect 519186 30258 519422 30494
rect 519186 23258 519422 23494
rect 519186 16258 519422 16494
rect 519186 9258 519422 9494
rect 519186 2258 519422 2494
rect 519186 -982 519422 -746
rect 519186 -1302 519422 -1066
rect 520918 234325 521154 234561
rect 520918 227325 521154 227561
rect 520918 220325 521154 220561
rect 520918 213325 521154 213561
rect 520918 206325 521154 206561
rect 520918 199325 521154 199561
rect 520918 192325 521154 192561
rect 520918 185325 521154 185561
rect 520918 178325 521154 178561
rect 520918 171325 521154 171561
rect 520918 164325 521154 164561
rect 520918 157325 521154 157561
rect 520918 150325 521154 150561
rect 520918 143325 521154 143561
rect 520918 136325 521154 136561
rect 520918 129325 521154 129561
rect 520918 122325 521154 122561
rect 520918 115325 521154 115561
rect 520918 108325 521154 108561
rect 520918 101325 521154 101561
rect 520918 94325 521154 94561
rect 520918 87325 521154 87561
rect 520918 80325 521154 80561
rect 520918 73325 521154 73561
rect 520918 66325 521154 66561
rect 520918 59325 521154 59561
rect 520918 52325 521154 52561
rect 520918 45325 521154 45561
rect 520918 38325 521154 38561
rect 520918 31325 521154 31561
rect 520918 24325 521154 24561
rect 520918 17325 521154 17561
rect 520918 10325 521154 10561
rect 520918 3325 521154 3561
rect 520918 -1942 521154 -1706
rect 520918 -2262 521154 -2026
rect 526186 233258 526422 233494
rect 526186 226258 526422 226494
rect 526186 219258 526422 219494
rect 526186 212258 526422 212494
rect 526186 205258 526422 205494
rect 526186 198258 526422 198494
rect 526186 191258 526422 191494
rect 526186 184258 526422 184494
rect 526186 177258 526422 177494
rect 526186 170258 526422 170494
rect 526186 163258 526422 163494
rect 526186 156258 526422 156494
rect 526186 149258 526422 149494
rect 526186 142258 526422 142494
rect 526186 135258 526422 135494
rect 526186 128258 526422 128494
rect 526186 121258 526422 121494
rect 526186 114258 526422 114494
rect 526186 107258 526422 107494
rect 526186 100258 526422 100494
rect 526186 93258 526422 93494
rect 526186 86258 526422 86494
rect 526186 79258 526422 79494
rect 526186 72258 526422 72494
rect 526186 65258 526422 65494
rect 526186 58258 526422 58494
rect 526186 51258 526422 51494
rect 526186 44258 526422 44494
rect 526186 37258 526422 37494
rect 526186 30258 526422 30494
rect 526186 23258 526422 23494
rect 526186 16258 526422 16494
rect 526186 9258 526422 9494
rect 526186 2258 526422 2494
rect 526186 -982 526422 -746
rect 526186 -1302 526422 -1066
rect 527918 234325 528154 234561
rect 527918 227325 528154 227561
rect 527918 220325 528154 220561
rect 527918 213325 528154 213561
rect 527918 206325 528154 206561
rect 527918 199325 528154 199561
rect 527918 192325 528154 192561
rect 527918 185325 528154 185561
rect 527918 178325 528154 178561
rect 527918 171325 528154 171561
rect 527918 164325 528154 164561
rect 527918 157325 528154 157561
rect 527918 150325 528154 150561
rect 527918 143325 528154 143561
rect 527918 136325 528154 136561
rect 527918 129325 528154 129561
rect 527918 122325 528154 122561
rect 527918 115325 528154 115561
rect 527918 108325 528154 108561
rect 527918 101325 528154 101561
rect 527918 94325 528154 94561
rect 527918 87325 528154 87561
rect 527918 80325 528154 80561
rect 527918 73325 528154 73561
rect 527918 66325 528154 66561
rect 527918 59325 528154 59561
rect 527918 52325 528154 52561
rect 527918 45325 528154 45561
rect 527918 38325 528154 38561
rect 527918 31325 528154 31561
rect 527918 24325 528154 24561
rect 527918 17325 528154 17561
rect 527918 10325 528154 10561
rect 527918 3325 528154 3561
rect 527918 -1942 528154 -1706
rect 527918 -2262 528154 -2026
rect 533186 705002 533422 705238
rect 533186 704682 533422 704918
rect 533186 695258 533422 695494
rect 533186 688258 533422 688494
rect 533186 681258 533422 681494
rect 533186 674258 533422 674494
rect 533186 667258 533422 667494
rect 533186 660258 533422 660494
rect 533186 653258 533422 653494
rect 533186 646258 533422 646494
rect 533186 639258 533422 639494
rect 533186 632258 533422 632494
rect 533186 625258 533422 625494
rect 533186 618258 533422 618494
rect 533186 611258 533422 611494
rect 533186 604258 533422 604494
rect 533186 597258 533422 597494
rect 533186 590258 533422 590494
rect 533186 583258 533422 583494
rect 533186 576258 533422 576494
rect 533186 569258 533422 569494
rect 533186 562258 533422 562494
rect 533186 555258 533422 555494
rect 533186 548258 533422 548494
rect 533186 541258 533422 541494
rect 533186 534258 533422 534494
rect 533186 527258 533422 527494
rect 533186 520258 533422 520494
rect 533186 513258 533422 513494
rect 533186 506258 533422 506494
rect 533186 499258 533422 499494
rect 533186 492258 533422 492494
rect 533186 485258 533422 485494
rect 533186 478258 533422 478494
rect 533186 471258 533422 471494
rect 533186 464258 533422 464494
rect 533186 457258 533422 457494
rect 533186 450258 533422 450494
rect 533186 443258 533422 443494
rect 533186 436258 533422 436494
rect 533186 429258 533422 429494
rect 533186 422258 533422 422494
rect 533186 415258 533422 415494
rect 533186 408258 533422 408494
rect 533186 401258 533422 401494
rect 533186 394258 533422 394494
rect 533186 387258 533422 387494
rect 533186 380258 533422 380494
rect 533186 373258 533422 373494
rect 533186 366258 533422 366494
rect 533186 359258 533422 359494
rect 533186 352258 533422 352494
rect 533186 345258 533422 345494
rect 533186 338258 533422 338494
rect 533186 331258 533422 331494
rect 533186 324258 533422 324494
rect 533186 317258 533422 317494
rect 533186 310258 533422 310494
rect 533186 303258 533422 303494
rect 533186 296258 533422 296494
rect 533186 289258 533422 289494
rect 533186 282258 533422 282494
rect 533186 275258 533422 275494
rect 533186 268258 533422 268494
rect 533186 261258 533422 261494
rect 533186 254258 533422 254494
rect 533186 247258 533422 247494
rect 533186 240258 533422 240494
rect 533186 233258 533422 233494
rect 533186 226258 533422 226494
rect 533186 219258 533422 219494
rect 533186 212258 533422 212494
rect 533186 205258 533422 205494
rect 533186 198258 533422 198494
rect 533186 191258 533422 191494
rect 533186 184258 533422 184494
rect 533186 177258 533422 177494
rect 533186 170258 533422 170494
rect 533186 163258 533422 163494
rect 533186 156258 533422 156494
rect 533186 149258 533422 149494
rect 533186 142258 533422 142494
rect 533186 135258 533422 135494
rect 533186 128258 533422 128494
rect 533186 121258 533422 121494
rect 533186 114258 533422 114494
rect 533186 107258 533422 107494
rect 533186 100258 533422 100494
rect 533186 93258 533422 93494
rect 533186 86258 533422 86494
rect 533186 79258 533422 79494
rect 533186 72258 533422 72494
rect 533186 65258 533422 65494
rect 533186 58258 533422 58494
rect 533186 51258 533422 51494
rect 533186 44258 533422 44494
rect 533186 37258 533422 37494
rect 533186 30258 533422 30494
rect 533186 23258 533422 23494
rect 533186 16258 533422 16494
rect 533186 9258 533422 9494
rect 533186 2258 533422 2494
rect 533186 -982 533422 -746
rect 533186 -1302 533422 -1066
rect 534918 705962 535154 706198
rect 534918 705642 535154 705878
rect 534918 696325 535154 696561
rect 534918 689325 535154 689561
rect 534918 682325 535154 682561
rect 534918 675325 535154 675561
rect 534918 668325 535154 668561
rect 534918 661325 535154 661561
rect 534918 654325 535154 654561
rect 534918 647325 535154 647561
rect 534918 640325 535154 640561
rect 534918 633325 535154 633561
rect 534918 626325 535154 626561
rect 534918 619325 535154 619561
rect 534918 612325 535154 612561
rect 534918 605325 535154 605561
rect 534918 598325 535154 598561
rect 534918 591325 535154 591561
rect 534918 584325 535154 584561
rect 534918 577325 535154 577561
rect 534918 570325 535154 570561
rect 534918 563325 535154 563561
rect 534918 556325 535154 556561
rect 534918 549325 535154 549561
rect 534918 542325 535154 542561
rect 534918 535325 535154 535561
rect 534918 528325 535154 528561
rect 534918 521325 535154 521561
rect 534918 514325 535154 514561
rect 534918 507325 535154 507561
rect 534918 500325 535154 500561
rect 534918 493325 535154 493561
rect 534918 486325 535154 486561
rect 534918 479325 535154 479561
rect 534918 472325 535154 472561
rect 534918 465325 535154 465561
rect 534918 458325 535154 458561
rect 534918 451325 535154 451561
rect 534918 444325 535154 444561
rect 534918 437325 535154 437561
rect 534918 430325 535154 430561
rect 534918 423325 535154 423561
rect 534918 416325 535154 416561
rect 534918 409325 535154 409561
rect 534918 402325 535154 402561
rect 534918 395325 535154 395561
rect 534918 388325 535154 388561
rect 534918 381325 535154 381561
rect 534918 374325 535154 374561
rect 534918 367325 535154 367561
rect 534918 360325 535154 360561
rect 534918 353325 535154 353561
rect 534918 346325 535154 346561
rect 534918 339325 535154 339561
rect 534918 332325 535154 332561
rect 534918 325325 535154 325561
rect 534918 318325 535154 318561
rect 534918 311325 535154 311561
rect 534918 304325 535154 304561
rect 534918 297325 535154 297561
rect 534918 290325 535154 290561
rect 534918 283325 535154 283561
rect 534918 276325 535154 276561
rect 534918 269325 535154 269561
rect 534918 262325 535154 262561
rect 534918 255325 535154 255561
rect 534918 248325 535154 248561
rect 534918 241325 535154 241561
rect 534918 234325 535154 234561
rect 534918 227325 535154 227561
rect 534918 220325 535154 220561
rect 534918 213325 535154 213561
rect 534918 206325 535154 206561
rect 534918 199325 535154 199561
rect 534918 192325 535154 192561
rect 534918 185325 535154 185561
rect 534918 178325 535154 178561
rect 534918 171325 535154 171561
rect 534918 164325 535154 164561
rect 534918 157325 535154 157561
rect 534918 150325 535154 150561
rect 534918 143325 535154 143561
rect 534918 136325 535154 136561
rect 534918 129325 535154 129561
rect 534918 122325 535154 122561
rect 534918 115325 535154 115561
rect 534918 108325 535154 108561
rect 534918 101325 535154 101561
rect 534918 94325 535154 94561
rect 534918 87325 535154 87561
rect 534918 80325 535154 80561
rect 534918 73325 535154 73561
rect 534918 66325 535154 66561
rect 534918 59325 535154 59561
rect 534918 52325 535154 52561
rect 534918 45325 535154 45561
rect 534918 38325 535154 38561
rect 534918 31325 535154 31561
rect 534918 24325 535154 24561
rect 534918 17325 535154 17561
rect 534918 10325 535154 10561
rect 534918 3325 535154 3561
rect 534918 -1942 535154 -1706
rect 534918 -2262 535154 -2026
rect 540186 705002 540422 705238
rect 540186 704682 540422 704918
rect 540186 695258 540422 695494
rect 540186 688258 540422 688494
rect 540186 681258 540422 681494
rect 540186 674258 540422 674494
rect 540186 667258 540422 667494
rect 540186 660258 540422 660494
rect 540186 653258 540422 653494
rect 540186 646258 540422 646494
rect 540186 639258 540422 639494
rect 540186 632258 540422 632494
rect 540186 625258 540422 625494
rect 540186 618258 540422 618494
rect 540186 611258 540422 611494
rect 540186 604258 540422 604494
rect 540186 597258 540422 597494
rect 540186 590258 540422 590494
rect 540186 583258 540422 583494
rect 540186 576258 540422 576494
rect 540186 569258 540422 569494
rect 540186 562258 540422 562494
rect 540186 555258 540422 555494
rect 540186 548258 540422 548494
rect 540186 541258 540422 541494
rect 540186 534258 540422 534494
rect 540186 527258 540422 527494
rect 540186 520258 540422 520494
rect 540186 513258 540422 513494
rect 540186 506258 540422 506494
rect 540186 499258 540422 499494
rect 540186 492258 540422 492494
rect 540186 485258 540422 485494
rect 540186 478258 540422 478494
rect 540186 471258 540422 471494
rect 540186 464258 540422 464494
rect 540186 457258 540422 457494
rect 540186 450258 540422 450494
rect 540186 443258 540422 443494
rect 540186 436258 540422 436494
rect 540186 429258 540422 429494
rect 540186 422258 540422 422494
rect 540186 415258 540422 415494
rect 540186 408258 540422 408494
rect 540186 401258 540422 401494
rect 540186 394258 540422 394494
rect 540186 387258 540422 387494
rect 540186 380258 540422 380494
rect 540186 373258 540422 373494
rect 540186 366258 540422 366494
rect 540186 359258 540422 359494
rect 540186 352258 540422 352494
rect 540186 345258 540422 345494
rect 540186 338258 540422 338494
rect 540186 331258 540422 331494
rect 540186 324258 540422 324494
rect 540186 317258 540422 317494
rect 540186 310258 540422 310494
rect 540186 303258 540422 303494
rect 540186 296258 540422 296494
rect 540186 289258 540422 289494
rect 540186 282258 540422 282494
rect 540186 275258 540422 275494
rect 540186 268258 540422 268494
rect 540186 261258 540422 261494
rect 540186 254258 540422 254494
rect 540186 247258 540422 247494
rect 540186 240258 540422 240494
rect 540186 233258 540422 233494
rect 540186 226258 540422 226494
rect 540186 219258 540422 219494
rect 540186 212258 540422 212494
rect 540186 205258 540422 205494
rect 540186 198258 540422 198494
rect 540186 191258 540422 191494
rect 540186 184258 540422 184494
rect 540186 177258 540422 177494
rect 540186 170258 540422 170494
rect 540186 163258 540422 163494
rect 540186 156258 540422 156494
rect 540186 149258 540422 149494
rect 540186 142258 540422 142494
rect 540186 135258 540422 135494
rect 540186 128258 540422 128494
rect 540186 121258 540422 121494
rect 540186 114258 540422 114494
rect 540186 107258 540422 107494
rect 540186 100258 540422 100494
rect 540186 93258 540422 93494
rect 540186 86258 540422 86494
rect 540186 79258 540422 79494
rect 540186 72258 540422 72494
rect 540186 65258 540422 65494
rect 540186 58258 540422 58494
rect 540186 51258 540422 51494
rect 540186 44258 540422 44494
rect 540186 37258 540422 37494
rect 540186 30258 540422 30494
rect 540186 23258 540422 23494
rect 540186 16258 540422 16494
rect 540186 9258 540422 9494
rect 540186 2258 540422 2494
rect 540186 -982 540422 -746
rect 540186 -1302 540422 -1066
rect 541918 705962 542154 706198
rect 541918 705642 542154 705878
rect 541918 696325 542154 696561
rect 541918 689325 542154 689561
rect 541918 682325 542154 682561
rect 541918 675325 542154 675561
rect 541918 668325 542154 668561
rect 541918 661325 542154 661561
rect 541918 654325 542154 654561
rect 541918 647325 542154 647561
rect 541918 640325 542154 640561
rect 541918 633325 542154 633561
rect 541918 626325 542154 626561
rect 541918 619325 542154 619561
rect 541918 612325 542154 612561
rect 541918 605325 542154 605561
rect 541918 598325 542154 598561
rect 541918 591325 542154 591561
rect 541918 584325 542154 584561
rect 541918 577325 542154 577561
rect 541918 570325 542154 570561
rect 541918 563325 542154 563561
rect 541918 556325 542154 556561
rect 541918 549325 542154 549561
rect 541918 542325 542154 542561
rect 541918 535325 542154 535561
rect 541918 528325 542154 528561
rect 541918 521325 542154 521561
rect 541918 514325 542154 514561
rect 541918 507325 542154 507561
rect 541918 500325 542154 500561
rect 541918 493325 542154 493561
rect 541918 486325 542154 486561
rect 541918 479325 542154 479561
rect 541918 472325 542154 472561
rect 541918 465325 542154 465561
rect 541918 458325 542154 458561
rect 541918 451325 542154 451561
rect 541918 444325 542154 444561
rect 541918 437325 542154 437561
rect 541918 430325 542154 430561
rect 541918 423325 542154 423561
rect 541918 416325 542154 416561
rect 541918 409325 542154 409561
rect 541918 402325 542154 402561
rect 541918 395325 542154 395561
rect 541918 388325 542154 388561
rect 541918 381325 542154 381561
rect 541918 374325 542154 374561
rect 541918 367325 542154 367561
rect 541918 360325 542154 360561
rect 541918 353325 542154 353561
rect 541918 346325 542154 346561
rect 541918 339325 542154 339561
rect 541918 332325 542154 332561
rect 541918 325325 542154 325561
rect 541918 318325 542154 318561
rect 541918 311325 542154 311561
rect 541918 304325 542154 304561
rect 541918 297325 542154 297561
rect 541918 290325 542154 290561
rect 541918 283325 542154 283561
rect 541918 276325 542154 276561
rect 541918 269325 542154 269561
rect 541918 262325 542154 262561
rect 541918 255325 542154 255561
rect 541918 248325 542154 248561
rect 541918 241325 542154 241561
rect 541918 234325 542154 234561
rect 541918 227325 542154 227561
rect 541918 220325 542154 220561
rect 541918 213325 542154 213561
rect 541918 206325 542154 206561
rect 541918 199325 542154 199561
rect 541918 192325 542154 192561
rect 541918 185325 542154 185561
rect 541918 178325 542154 178561
rect 541918 171325 542154 171561
rect 541918 164325 542154 164561
rect 541918 157325 542154 157561
rect 541918 150325 542154 150561
rect 541918 143325 542154 143561
rect 541918 136325 542154 136561
rect 541918 129325 542154 129561
rect 541918 122325 542154 122561
rect 541918 115325 542154 115561
rect 541918 108325 542154 108561
rect 541918 101325 542154 101561
rect 541918 94325 542154 94561
rect 541918 87325 542154 87561
rect 541918 80325 542154 80561
rect 541918 73325 542154 73561
rect 541918 66325 542154 66561
rect 541918 59325 542154 59561
rect 541918 52325 542154 52561
rect 541918 45325 542154 45561
rect 541918 38325 542154 38561
rect 541918 31325 542154 31561
rect 541918 24325 542154 24561
rect 541918 17325 542154 17561
rect 541918 10325 542154 10561
rect 541918 3325 542154 3561
rect 541918 -1942 542154 -1706
rect 541918 -2262 542154 -2026
rect 547186 705002 547422 705238
rect 547186 704682 547422 704918
rect 547186 695258 547422 695494
rect 547186 688258 547422 688494
rect 547186 681258 547422 681494
rect 547186 674258 547422 674494
rect 547186 667258 547422 667494
rect 547186 660258 547422 660494
rect 547186 653258 547422 653494
rect 547186 646258 547422 646494
rect 547186 639258 547422 639494
rect 547186 632258 547422 632494
rect 547186 625258 547422 625494
rect 547186 618258 547422 618494
rect 547186 611258 547422 611494
rect 547186 604258 547422 604494
rect 547186 597258 547422 597494
rect 547186 590258 547422 590494
rect 547186 583258 547422 583494
rect 547186 576258 547422 576494
rect 547186 569258 547422 569494
rect 547186 562258 547422 562494
rect 547186 555258 547422 555494
rect 547186 548258 547422 548494
rect 547186 541258 547422 541494
rect 547186 534258 547422 534494
rect 547186 527258 547422 527494
rect 547186 520258 547422 520494
rect 547186 513258 547422 513494
rect 547186 506258 547422 506494
rect 547186 499258 547422 499494
rect 547186 492258 547422 492494
rect 547186 485258 547422 485494
rect 547186 478258 547422 478494
rect 547186 471258 547422 471494
rect 547186 464258 547422 464494
rect 547186 457258 547422 457494
rect 547186 450258 547422 450494
rect 547186 443258 547422 443494
rect 547186 436258 547422 436494
rect 547186 429258 547422 429494
rect 547186 422258 547422 422494
rect 547186 415258 547422 415494
rect 547186 408258 547422 408494
rect 547186 401258 547422 401494
rect 547186 394258 547422 394494
rect 547186 387258 547422 387494
rect 547186 380258 547422 380494
rect 547186 373258 547422 373494
rect 547186 366258 547422 366494
rect 547186 359258 547422 359494
rect 547186 352258 547422 352494
rect 547186 345258 547422 345494
rect 547186 338258 547422 338494
rect 547186 331258 547422 331494
rect 547186 324258 547422 324494
rect 547186 317258 547422 317494
rect 547186 310258 547422 310494
rect 547186 303258 547422 303494
rect 547186 296258 547422 296494
rect 547186 289258 547422 289494
rect 547186 282258 547422 282494
rect 547186 275258 547422 275494
rect 547186 268258 547422 268494
rect 547186 261258 547422 261494
rect 547186 254258 547422 254494
rect 547186 247258 547422 247494
rect 547186 240258 547422 240494
rect 547186 233258 547422 233494
rect 547186 226258 547422 226494
rect 547186 219258 547422 219494
rect 547186 212258 547422 212494
rect 547186 205258 547422 205494
rect 547186 198258 547422 198494
rect 547186 191258 547422 191494
rect 547186 184258 547422 184494
rect 547186 177258 547422 177494
rect 547186 170258 547422 170494
rect 547186 163258 547422 163494
rect 547186 156258 547422 156494
rect 547186 149258 547422 149494
rect 547186 142258 547422 142494
rect 547186 135258 547422 135494
rect 547186 128258 547422 128494
rect 547186 121258 547422 121494
rect 547186 114258 547422 114494
rect 547186 107258 547422 107494
rect 547186 100258 547422 100494
rect 547186 93258 547422 93494
rect 547186 86258 547422 86494
rect 547186 79258 547422 79494
rect 547186 72258 547422 72494
rect 547186 65258 547422 65494
rect 547186 58258 547422 58494
rect 547186 51258 547422 51494
rect 547186 44258 547422 44494
rect 547186 37258 547422 37494
rect 547186 30258 547422 30494
rect 547186 23258 547422 23494
rect 547186 16258 547422 16494
rect 547186 9258 547422 9494
rect 547186 2258 547422 2494
rect 547186 -982 547422 -746
rect 547186 -1302 547422 -1066
rect 548918 705962 549154 706198
rect 548918 705642 549154 705878
rect 548918 696325 549154 696561
rect 548918 689325 549154 689561
rect 548918 682325 549154 682561
rect 548918 675325 549154 675561
rect 548918 668325 549154 668561
rect 548918 661325 549154 661561
rect 548918 654325 549154 654561
rect 548918 647325 549154 647561
rect 548918 640325 549154 640561
rect 548918 633325 549154 633561
rect 548918 626325 549154 626561
rect 548918 619325 549154 619561
rect 548918 612325 549154 612561
rect 548918 605325 549154 605561
rect 548918 598325 549154 598561
rect 548918 591325 549154 591561
rect 548918 584325 549154 584561
rect 548918 577325 549154 577561
rect 548918 570325 549154 570561
rect 548918 563325 549154 563561
rect 548918 556325 549154 556561
rect 548918 549325 549154 549561
rect 548918 542325 549154 542561
rect 548918 535325 549154 535561
rect 548918 528325 549154 528561
rect 548918 521325 549154 521561
rect 548918 514325 549154 514561
rect 548918 507325 549154 507561
rect 548918 500325 549154 500561
rect 548918 493325 549154 493561
rect 548918 486325 549154 486561
rect 548918 479325 549154 479561
rect 548918 472325 549154 472561
rect 548918 465325 549154 465561
rect 548918 458325 549154 458561
rect 548918 451325 549154 451561
rect 548918 444325 549154 444561
rect 548918 437325 549154 437561
rect 548918 430325 549154 430561
rect 548918 423325 549154 423561
rect 548918 416325 549154 416561
rect 548918 409325 549154 409561
rect 548918 402325 549154 402561
rect 548918 395325 549154 395561
rect 548918 388325 549154 388561
rect 548918 381325 549154 381561
rect 548918 374325 549154 374561
rect 548918 367325 549154 367561
rect 548918 360325 549154 360561
rect 548918 353325 549154 353561
rect 548918 346325 549154 346561
rect 548918 339325 549154 339561
rect 548918 332325 549154 332561
rect 548918 325325 549154 325561
rect 548918 318325 549154 318561
rect 548918 311325 549154 311561
rect 548918 304325 549154 304561
rect 548918 297325 549154 297561
rect 548918 290325 549154 290561
rect 548918 283325 549154 283561
rect 548918 276325 549154 276561
rect 548918 269325 549154 269561
rect 548918 262325 549154 262561
rect 548918 255325 549154 255561
rect 548918 248325 549154 248561
rect 548918 241325 549154 241561
rect 548918 234325 549154 234561
rect 548918 227325 549154 227561
rect 548918 220325 549154 220561
rect 548918 213325 549154 213561
rect 548918 206325 549154 206561
rect 548918 199325 549154 199561
rect 548918 192325 549154 192561
rect 548918 185325 549154 185561
rect 548918 178325 549154 178561
rect 548918 171325 549154 171561
rect 548918 164325 549154 164561
rect 548918 157325 549154 157561
rect 548918 150325 549154 150561
rect 548918 143325 549154 143561
rect 548918 136325 549154 136561
rect 548918 129325 549154 129561
rect 548918 122325 549154 122561
rect 548918 115325 549154 115561
rect 548918 108325 549154 108561
rect 548918 101325 549154 101561
rect 548918 94325 549154 94561
rect 548918 87325 549154 87561
rect 548918 80325 549154 80561
rect 548918 73325 549154 73561
rect 548918 66325 549154 66561
rect 548918 59325 549154 59561
rect 548918 52325 549154 52561
rect 548918 45325 549154 45561
rect 548918 38325 549154 38561
rect 548918 31325 549154 31561
rect 548918 24325 549154 24561
rect 548918 17325 549154 17561
rect 548918 10325 549154 10561
rect 548918 3325 549154 3561
rect 548918 -1942 549154 -1706
rect 548918 -2262 549154 -2026
rect 554186 705002 554422 705238
rect 554186 704682 554422 704918
rect 554186 695258 554422 695494
rect 554186 688258 554422 688494
rect 554186 681258 554422 681494
rect 554186 674258 554422 674494
rect 554186 667258 554422 667494
rect 554186 660258 554422 660494
rect 554186 653258 554422 653494
rect 554186 646258 554422 646494
rect 554186 639258 554422 639494
rect 554186 632258 554422 632494
rect 554186 625258 554422 625494
rect 554186 618258 554422 618494
rect 554186 611258 554422 611494
rect 554186 604258 554422 604494
rect 554186 597258 554422 597494
rect 554186 590258 554422 590494
rect 554186 583258 554422 583494
rect 554186 576258 554422 576494
rect 554186 569258 554422 569494
rect 554186 562258 554422 562494
rect 554186 555258 554422 555494
rect 554186 548258 554422 548494
rect 554186 541258 554422 541494
rect 554186 534258 554422 534494
rect 554186 527258 554422 527494
rect 554186 520258 554422 520494
rect 554186 513258 554422 513494
rect 554186 506258 554422 506494
rect 554186 499258 554422 499494
rect 554186 492258 554422 492494
rect 554186 485258 554422 485494
rect 554186 478258 554422 478494
rect 554186 471258 554422 471494
rect 554186 464258 554422 464494
rect 554186 457258 554422 457494
rect 554186 450258 554422 450494
rect 554186 443258 554422 443494
rect 554186 436258 554422 436494
rect 554186 429258 554422 429494
rect 554186 422258 554422 422494
rect 554186 415258 554422 415494
rect 554186 408258 554422 408494
rect 554186 401258 554422 401494
rect 554186 394258 554422 394494
rect 554186 387258 554422 387494
rect 554186 380258 554422 380494
rect 554186 373258 554422 373494
rect 554186 366258 554422 366494
rect 554186 359258 554422 359494
rect 554186 352258 554422 352494
rect 554186 345258 554422 345494
rect 554186 338258 554422 338494
rect 554186 331258 554422 331494
rect 554186 324258 554422 324494
rect 554186 317258 554422 317494
rect 554186 310258 554422 310494
rect 554186 303258 554422 303494
rect 554186 296258 554422 296494
rect 554186 289258 554422 289494
rect 554186 282258 554422 282494
rect 554186 275258 554422 275494
rect 554186 268258 554422 268494
rect 554186 261258 554422 261494
rect 554186 254258 554422 254494
rect 554186 247258 554422 247494
rect 554186 240258 554422 240494
rect 554186 233258 554422 233494
rect 554186 226258 554422 226494
rect 554186 219258 554422 219494
rect 554186 212258 554422 212494
rect 554186 205258 554422 205494
rect 554186 198258 554422 198494
rect 554186 191258 554422 191494
rect 554186 184258 554422 184494
rect 554186 177258 554422 177494
rect 554186 170258 554422 170494
rect 554186 163258 554422 163494
rect 554186 156258 554422 156494
rect 554186 149258 554422 149494
rect 554186 142258 554422 142494
rect 554186 135258 554422 135494
rect 554186 128258 554422 128494
rect 554186 121258 554422 121494
rect 554186 114258 554422 114494
rect 554186 107258 554422 107494
rect 554186 100258 554422 100494
rect 554186 93258 554422 93494
rect 554186 86258 554422 86494
rect 554186 79258 554422 79494
rect 554186 72258 554422 72494
rect 554186 65258 554422 65494
rect 554186 58258 554422 58494
rect 554186 51258 554422 51494
rect 554186 44258 554422 44494
rect 554186 37258 554422 37494
rect 554186 30258 554422 30494
rect 554186 23258 554422 23494
rect 554186 16258 554422 16494
rect 554186 9258 554422 9494
rect 554186 2258 554422 2494
rect 554186 -982 554422 -746
rect 554186 -1302 554422 -1066
rect 555918 705962 556154 706198
rect 555918 705642 556154 705878
rect 555918 696325 556154 696561
rect 555918 689325 556154 689561
rect 555918 682325 556154 682561
rect 555918 675325 556154 675561
rect 555918 668325 556154 668561
rect 555918 661325 556154 661561
rect 555918 654325 556154 654561
rect 555918 647325 556154 647561
rect 555918 640325 556154 640561
rect 555918 633325 556154 633561
rect 555918 626325 556154 626561
rect 555918 619325 556154 619561
rect 555918 612325 556154 612561
rect 555918 605325 556154 605561
rect 555918 598325 556154 598561
rect 555918 591325 556154 591561
rect 555918 584325 556154 584561
rect 555918 577325 556154 577561
rect 555918 570325 556154 570561
rect 555918 563325 556154 563561
rect 555918 556325 556154 556561
rect 555918 549325 556154 549561
rect 555918 542325 556154 542561
rect 555918 535325 556154 535561
rect 555918 528325 556154 528561
rect 555918 521325 556154 521561
rect 555918 514325 556154 514561
rect 555918 507325 556154 507561
rect 555918 500325 556154 500561
rect 555918 493325 556154 493561
rect 555918 486325 556154 486561
rect 555918 479325 556154 479561
rect 555918 472325 556154 472561
rect 555918 465325 556154 465561
rect 555918 458325 556154 458561
rect 555918 451325 556154 451561
rect 555918 444325 556154 444561
rect 555918 437325 556154 437561
rect 555918 430325 556154 430561
rect 555918 423325 556154 423561
rect 555918 416325 556154 416561
rect 555918 409325 556154 409561
rect 555918 402325 556154 402561
rect 555918 395325 556154 395561
rect 555918 388325 556154 388561
rect 555918 381325 556154 381561
rect 555918 374325 556154 374561
rect 555918 367325 556154 367561
rect 555918 360325 556154 360561
rect 555918 353325 556154 353561
rect 555918 346325 556154 346561
rect 555918 339325 556154 339561
rect 555918 332325 556154 332561
rect 555918 325325 556154 325561
rect 555918 318325 556154 318561
rect 555918 311325 556154 311561
rect 555918 304325 556154 304561
rect 555918 297325 556154 297561
rect 555918 290325 556154 290561
rect 555918 283325 556154 283561
rect 555918 276325 556154 276561
rect 555918 269325 556154 269561
rect 555918 262325 556154 262561
rect 555918 255325 556154 255561
rect 555918 248325 556154 248561
rect 555918 241325 556154 241561
rect 555918 234325 556154 234561
rect 555918 227325 556154 227561
rect 555918 220325 556154 220561
rect 555918 213325 556154 213561
rect 555918 206325 556154 206561
rect 555918 199325 556154 199561
rect 555918 192325 556154 192561
rect 555918 185325 556154 185561
rect 555918 178325 556154 178561
rect 555918 171325 556154 171561
rect 555918 164325 556154 164561
rect 555918 157325 556154 157561
rect 555918 150325 556154 150561
rect 555918 143325 556154 143561
rect 555918 136325 556154 136561
rect 555918 129325 556154 129561
rect 555918 122325 556154 122561
rect 555918 115325 556154 115561
rect 555918 108325 556154 108561
rect 555918 101325 556154 101561
rect 555918 94325 556154 94561
rect 555918 87325 556154 87561
rect 555918 80325 556154 80561
rect 555918 73325 556154 73561
rect 555918 66325 556154 66561
rect 555918 59325 556154 59561
rect 555918 52325 556154 52561
rect 555918 45325 556154 45561
rect 555918 38325 556154 38561
rect 555918 31325 556154 31561
rect 555918 24325 556154 24561
rect 555918 17325 556154 17561
rect 555918 10325 556154 10561
rect 555918 3325 556154 3561
rect 555918 -1942 556154 -1706
rect 555918 -2262 556154 -2026
rect 561186 705002 561422 705238
rect 561186 704682 561422 704918
rect 561186 695258 561422 695494
rect 561186 688258 561422 688494
rect 561186 681258 561422 681494
rect 561186 674258 561422 674494
rect 561186 667258 561422 667494
rect 561186 660258 561422 660494
rect 561186 653258 561422 653494
rect 561186 646258 561422 646494
rect 561186 639258 561422 639494
rect 561186 632258 561422 632494
rect 561186 625258 561422 625494
rect 561186 618258 561422 618494
rect 561186 611258 561422 611494
rect 561186 604258 561422 604494
rect 561186 597258 561422 597494
rect 561186 590258 561422 590494
rect 561186 583258 561422 583494
rect 561186 576258 561422 576494
rect 561186 569258 561422 569494
rect 561186 562258 561422 562494
rect 561186 555258 561422 555494
rect 561186 548258 561422 548494
rect 561186 541258 561422 541494
rect 561186 534258 561422 534494
rect 561186 527258 561422 527494
rect 561186 520258 561422 520494
rect 561186 513258 561422 513494
rect 561186 506258 561422 506494
rect 561186 499258 561422 499494
rect 561186 492258 561422 492494
rect 561186 485258 561422 485494
rect 561186 478258 561422 478494
rect 561186 471258 561422 471494
rect 561186 464258 561422 464494
rect 561186 457258 561422 457494
rect 561186 450258 561422 450494
rect 561186 443258 561422 443494
rect 561186 436258 561422 436494
rect 561186 429258 561422 429494
rect 561186 422258 561422 422494
rect 561186 415258 561422 415494
rect 561186 408258 561422 408494
rect 561186 401258 561422 401494
rect 561186 394258 561422 394494
rect 561186 387258 561422 387494
rect 561186 380258 561422 380494
rect 561186 373258 561422 373494
rect 561186 366258 561422 366494
rect 561186 359258 561422 359494
rect 561186 352258 561422 352494
rect 561186 345258 561422 345494
rect 561186 338258 561422 338494
rect 561186 331258 561422 331494
rect 561186 324258 561422 324494
rect 561186 317258 561422 317494
rect 561186 310258 561422 310494
rect 561186 303258 561422 303494
rect 561186 296258 561422 296494
rect 561186 289258 561422 289494
rect 561186 282258 561422 282494
rect 561186 275258 561422 275494
rect 561186 268258 561422 268494
rect 561186 261258 561422 261494
rect 561186 254258 561422 254494
rect 561186 247258 561422 247494
rect 561186 240258 561422 240494
rect 561186 233258 561422 233494
rect 561186 226258 561422 226494
rect 561186 219258 561422 219494
rect 561186 212258 561422 212494
rect 561186 205258 561422 205494
rect 561186 198258 561422 198494
rect 561186 191258 561422 191494
rect 561186 184258 561422 184494
rect 561186 177258 561422 177494
rect 561186 170258 561422 170494
rect 561186 163258 561422 163494
rect 561186 156258 561422 156494
rect 561186 149258 561422 149494
rect 561186 142258 561422 142494
rect 561186 135258 561422 135494
rect 561186 128258 561422 128494
rect 561186 121258 561422 121494
rect 561186 114258 561422 114494
rect 561186 107258 561422 107494
rect 561186 100258 561422 100494
rect 561186 93258 561422 93494
rect 561186 86258 561422 86494
rect 561186 79258 561422 79494
rect 561186 72258 561422 72494
rect 561186 65258 561422 65494
rect 561186 58258 561422 58494
rect 561186 51258 561422 51494
rect 561186 44258 561422 44494
rect 561186 37258 561422 37494
rect 561186 30258 561422 30494
rect 561186 23258 561422 23494
rect 561186 16258 561422 16494
rect 561186 9258 561422 9494
rect 561186 2258 561422 2494
rect 561186 -982 561422 -746
rect 561186 -1302 561422 -1066
rect 562918 705962 563154 706198
rect 562918 705642 563154 705878
rect 562918 696325 563154 696561
rect 562918 689325 563154 689561
rect 562918 682325 563154 682561
rect 562918 675325 563154 675561
rect 562918 668325 563154 668561
rect 562918 661325 563154 661561
rect 562918 654325 563154 654561
rect 562918 647325 563154 647561
rect 562918 640325 563154 640561
rect 562918 633325 563154 633561
rect 562918 626325 563154 626561
rect 562918 619325 563154 619561
rect 562918 612325 563154 612561
rect 562918 605325 563154 605561
rect 562918 598325 563154 598561
rect 562918 591325 563154 591561
rect 562918 584325 563154 584561
rect 562918 577325 563154 577561
rect 562918 570325 563154 570561
rect 562918 563325 563154 563561
rect 562918 556325 563154 556561
rect 562918 549325 563154 549561
rect 562918 542325 563154 542561
rect 562918 535325 563154 535561
rect 562918 528325 563154 528561
rect 562918 521325 563154 521561
rect 562918 514325 563154 514561
rect 562918 507325 563154 507561
rect 562918 500325 563154 500561
rect 562918 493325 563154 493561
rect 562918 486325 563154 486561
rect 562918 479325 563154 479561
rect 562918 472325 563154 472561
rect 562918 465325 563154 465561
rect 562918 458325 563154 458561
rect 562918 451325 563154 451561
rect 562918 444325 563154 444561
rect 562918 437325 563154 437561
rect 562918 430325 563154 430561
rect 562918 423325 563154 423561
rect 562918 416325 563154 416561
rect 562918 409325 563154 409561
rect 562918 402325 563154 402561
rect 562918 395325 563154 395561
rect 562918 388325 563154 388561
rect 562918 381325 563154 381561
rect 562918 374325 563154 374561
rect 562918 367325 563154 367561
rect 562918 360325 563154 360561
rect 562918 353325 563154 353561
rect 562918 346325 563154 346561
rect 562918 339325 563154 339561
rect 562918 332325 563154 332561
rect 562918 325325 563154 325561
rect 562918 318325 563154 318561
rect 562918 311325 563154 311561
rect 562918 304325 563154 304561
rect 562918 297325 563154 297561
rect 562918 290325 563154 290561
rect 562918 283325 563154 283561
rect 562918 276325 563154 276561
rect 562918 269325 563154 269561
rect 562918 262325 563154 262561
rect 562918 255325 563154 255561
rect 562918 248325 563154 248561
rect 562918 241325 563154 241561
rect 562918 234325 563154 234561
rect 562918 227325 563154 227561
rect 562918 220325 563154 220561
rect 562918 213325 563154 213561
rect 562918 206325 563154 206561
rect 562918 199325 563154 199561
rect 562918 192325 563154 192561
rect 562918 185325 563154 185561
rect 562918 178325 563154 178561
rect 562918 171325 563154 171561
rect 562918 164325 563154 164561
rect 562918 157325 563154 157561
rect 562918 150325 563154 150561
rect 562918 143325 563154 143561
rect 562918 136325 563154 136561
rect 562918 129325 563154 129561
rect 562918 122325 563154 122561
rect 562918 115325 563154 115561
rect 562918 108325 563154 108561
rect 562918 101325 563154 101561
rect 562918 94325 563154 94561
rect 562918 87325 563154 87561
rect 562918 80325 563154 80561
rect 562918 73325 563154 73561
rect 562918 66325 563154 66561
rect 562918 59325 563154 59561
rect 562918 52325 563154 52561
rect 562918 45325 563154 45561
rect 562918 38325 563154 38561
rect 562918 31325 563154 31561
rect 562918 24325 563154 24561
rect 562918 17325 563154 17561
rect 562918 10325 563154 10561
rect 562918 3325 563154 3561
rect 562918 -1942 563154 -1706
rect 562918 -2262 563154 -2026
rect 568186 705002 568422 705238
rect 568186 704682 568422 704918
rect 568186 695258 568422 695494
rect 568186 688258 568422 688494
rect 568186 681258 568422 681494
rect 568186 674258 568422 674494
rect 568186 667258 568422 667494
rect 568186 660258 568422 660494
rect 568186 653258 568422 653494
rect 568186 646258 568422 646494
rect 568186 639258 568422 639494
rect 568186 632258 568422 632494
rect 568186 625258 568422 625494
rect 568186 618258 568422 618494
rect 568186 611258 568422 611494
rect 568186 604258 568422 604494
rect 568186 597258 568422 597494
rect 568186 590258 568422 590494
rect 568186 583258 568422 583494
rect 568186 576258 568422 576494
rect 568186 569258 568422 569494
rect 568186 562258 568422 562494
rect 568186 555258 568422 555494
rect 568186 548258 568422 548494
rect 568186 541258 568422 541494
rect 568186 534258 568422 534494
rect 568186 527258 568422 527494
rect 568186 520258 568422 520494
rect 568186 513258 568422 513494
rect 568186 506258 568422 506494
rect 568186 499258 568422 499494
rect 568186 492258 568422 492494
rect 568186 485258 568422 485494
rect 568186 478258 568422 478494
rect 568186 471258 568422 471494
rect 568186 464258 568422 464494
rect 568186 457258 568422 457494
rect 568186 450258 568422 450494
rect 568186 443258 568422 443494
rect 568186 436258 568422 436494
rect 568186 429258 568422 429494
rect 568186 422258 568422 422494
rect 568186 415258 568422 415494
rect 568186 408258 568422 408494
rect 568186 401258 568422 401494
rect 568186 394258 568422 394494
rect 568186 387258 568422 387494
rect 568186 380258 568422 380494
rect 568186 373258 568422 373494
rect 568186 366258 568422 366494
rect 568186 359258 568422 359494
rect 568186 352258 568422 352494
rect 568186 345258 568422 345494
rect 568186 338258 568422 338494
rect 568186 331258 568422 331494
rect 568186 324258 568422 324494
rect 568186 317258 568422 317494
rect 568186 310258 568422 310494
rect 568186 303258 568422 303494
rect 568186 296258 568422 296494
rect 568186 289258 568422 289494
rect 568186 282258 568422 282494
rect 568186 275258 568422 275494
rect 568186 268258 568422 268494
rect 568186 261258 568422 261494
rect 568186 254258 568422 254494
rect 568186 247258 568422 247494
rect 568186 240258 568422 240494
rect 568186 233258 568422 233494
rect 568186 226258 568422 226494
rect 568186 219258 568422 219494
rect 568186 212258 568422 212494
rect 568186 205258 568422 205494
rect 568186 198258 568422 198494
rect 568186 191258 568422 191494
rect 568186 184258 568422 184494
rect 568186 177258 568422 177494
rect 568186 170258 568422 170494
rect 568186 163258 568422 163494
rect 568186 156258 568422 156494
rect 568186 149258 568422 149494
rect 568186 142258 568422 142494
rect 568186 135258 568422 135494
rect 568186 128258 568422 128494
rect 568186 121258 568422 121494
rect 568186 114258 568422 114494
rect 568186 107258 568422 107494
rect 568186 100258 568422 100494
rect 568186 93258 568422 93494
rect 568186 86258 568422 86494
rect 568186 79258 568422 79494
rect 568186 72258 568422 72494
rect 568186 65258 568422 65494
rect 568186 58258 568422 58494
rect 568186 51258 568422 51494
rect 568186 44258 568422 44494
rect 568186 37258 568422 37494
rect 568186 30258 568422 30494
rect 568186 23258 568422 23494
rect 568186 16258 568422 16494
rect 568186 9258 568422 9494
rect 568186 2258 568422 2494
rect 568186 -982 568422 -746
rect 568186 -1302 568422 -1066
rect 569918 705962 570154 706198
rect 569918 705642 570154 705878
rect 569918 696325 570154 696561
rect 569918 689325 570154 689561
rect 569918 682325 570154 682561
rect 569918 675325 570154 675561
rect 569918 668325 570154 668561
rect 569918 661325 570154 661561
rect 569918 654325 570154 654561
rect 569918 647325 570154 647561
rect 569918 640325 570154 640561
rect 569918 633325 570154 633561
rect 569918 626325 570154 626561
rect 569918 619325 570154 619561
rect 569918 612325 570154 612561
rect 569918 605325 570154 605561
rect 569918 598325 570154 598561
rect 569918 591325 570154 591561
rect 569918 584325 570154 584561
rect 569918 577325 570154 577561
rect 569918 570325 570154 570561
rect 569918 563325 570154 563561
rect 569918 556325 570154 556561
rect 569918 549325 570154 549561
rect 569918 542325 570154 542561
rect 569918 535325 570154 535561
rect 569918 528325 570154 528561
rect 569918 521325 570154 521561
rect 569918 514325 570154 514561
rect 569918 507325 570154 507561
rect 569918 500325 570154 500561
rect 569918 493325 570154 493561
rect 569918 486325 570154 486561
rect 569918 479325 570154 479561
rect 569918 472325 570154 472561
rect 569918 465325 570154 465561
rect 569918 458325 570154 458561
rect 569918 451325 570154 451561
rect 569918 444325 570154 444561
rect 569918 437325 570154 437561
rect 569918 430325 570154 430561
rect 569918 423325 570154 423561
rect 569918 416325 570154 416561
rect 569918 409325 570154 409561
rect 569918 402325 570154 402561
rect 569918 395325 570154 395561
rect 569918 388325 570154 388561
rect 569918 381325 570154 381561
rect 569918 374325 570154 374561
rect 569918 367325 570154 367561
rect 569918 360325 570154 360561
rect 569918 353325 570154 353561
rect 569918 346325 570154 346561
rect 569918 339325 570154 339561
rect 569918 332325 570154 332561
rect 569918 325325 570154 325561
rect 569918 318325 570154 318561
rect 569918 311325 570154 311561
rect 569918 304325 570154 304561
rect 569918 297325 570154 297561
rect 569918 290325 570154 290561
rect 569918 283325 570154 283561
rect 569918 276325 570154 276561
rect 569918 269325 570154 269561
rect 569918 262325 570154 262561
rect 569918 255325 570154 255561
rect 569918 248325 570154 248561
rect 569918 241325 570154 241561
rect 569918 234325 570154 234561
rect 569918 227325 570154 227561
rect 569918 220325 570154 220561
rect 569918 213325 570154 213561
rect 569918 206325 570154 206561
rect 569918 199325 570154 199561
rect 569918 192325 570154 192561
rect 569918 185325 570154 185561
rect 569918 178325 570154 178561
rect 569918 171325 570154 171561
rect 569918 164325 570154 164561
rect 569918 157325 570154 157561
rect 569918 150325 570154 150561
rect 569918 143325 570154 143561
rect 569918 136325 570154 136561
rect 569918 129325 570154 129561
rect 569918 122325 570154 122561
rect 569918 115325 570154 115561
rect 569918 108325 570154 108561
rect 569918 101325 570154 101561
rect 569918 94325 570154 94561
rect 569918 87325 570154 87561
rect 569918 80325 570154 80561
rect 569918 73325 570154 73561
rect 569918 66325 570154 66561
rect 569918 59325 570154 59561
rect 569918 52325 570154 52561
rect 569918 45325 570154 45561
rect 569918 38325 570154 38561
rect 569918 31325 570154 31561
rect 569918 24325 570154 24561
rect 569918 17325 570154 17561
rect 569918 10325 570154 10561
rect 569918 3325 570154 3561
rect 569918 -1942 570154 -1706
rect 569918 -2262 570154 -2026
rect 575186 705002 575422 705238
rect 575186 704682 575422 704918
rect 575186 695258 575422 695494
rect 575186 688258 575422 688494
rect 575186 681258 575422 681494
rect 575186 674258 575422 674494
rect 575186 667258 575422 667494
rect 575186 660258 575422 660494
rect 575186 653258 575422 653494
rect 575186 646258 575422 646494
rect 575186 639258 575422 639494
rect 575186 632258 575422 632494
rect 575186 625258 575422 625494
rect 575186 618258 575422 618494
rect 575186 611258 575422 611494
rect 575186 604258 575422 604494
rect 575186 597258 575422 597494
rect 575186 590258 575422 590494
rect 575186 583258 575422 583494
rect 575186 576258 575422 576494
rect 575186 569258 575422 569494
rect 575186 562258 575422 562494
rect 575186 555258 575422 555494
rect 575186 548258 575422 548494
rect 575186 541258 575422 541494
rect 575186 534258 575422 534494
rect 575186 527258 575422 527494
rect 575186 520258 575422 520494
rect 575186 513258 575422 513494
rect 575186 506258 575422 506494
rect 575186 499258 575422 499494
rect 575186 492258 575422 492494
rect 575186 485258 575422 485494
rect 575186 478258 575422 478494
rect 575186 471258 575422 471494
rect 575186 464258 575422 464494
rect 575186 457258 575422 457494
rect 575186 450258 575422 450494
rect 575186 443258 575422 443494
rect 575186 436258 575422 436494
rect 575186 429258 575422 429494
rect 575186 422258 575422 422494
rect 575186 415258 575422 415494
rect 575186 408258 575422 408494
rect 575186 401258 575422 401494
rect 575186 394258 575422 394494
rect 575186 387258 575422 387494
rect 575186 380258 575422 380494
rect 575186 373258 575422 373494
rect 575186 366258 575422 366494
rect 575186 359258 575422 359494
rect 575186 352258 575422 352494
rect 575186 345258 575422 345494
rect 575186 338258 575422 338494
rect 575186 331258 575422 331494
rect 575186 324258 575422 324494
rect 575186 317258 575422 317494
rect 575186 310258 575422 310494
rect 575186 303258 575422 303494
rect 575186 296258 575422 296494
rect 575186 289258 575422 289494
rect 575186 282258 575422 282494
rect 575186 275258 575422 275494
rect 575186 268258 575422 268494
rect 575186 261258 575422 261494
rect 575186 254258 575422 254494
rect 575186 247258 575422 247494
rect 575186 240258 575422 240494
rect 575186 233258 575422 233494
rect 575186 226258 575422 226494
rect 575186 219258 575422 219494
rect 575186 212258 575422 212494
rect 575186 205258 575422 205494
rect 575186 198258 575422 198494
rect 575186 191258 575422 191494
rect 575186 184258 575422 184494
rect 575186 177258 575422 177494
rect 575186 170258 575422 170494
rect 575186 163258 575422 163494
rect 575186 156258 575422 156494
rect 575186 149258 575422 149494
rect 575186 142258 575422 142494
rect 575186 135258 575422 135494
rect 575186 128258 575422 128494
rect 575186 121258 575422 121494
rect 575186 114258 575422 114494
rect 575186 107258 575422 107494
rect 575186 100258 575422 100494
rect 575186 93258 575422 93494
rect 575186 86258 575422 86494
rect 575186 79258 575422 79494
rect 575186 72258 575422 72494
rect 575186 65258 575422 65494
rect 575186 58258 575422 58494
rect 575186 51258 575422 51494
rect 575186 44258 575422 44494
rect 575186 37258 575422 37494
rect 575186 30258 575422 30494
rect 575186 23258 575422 23494
rect 575186 16258 575422 16494
rect 575186 9258 575422 9494
rect 575186 2258 575422 2494
rect 575186 -982 575422 -746
rect 575186 -1302 575422 -1066
rect 576918 705962 577154 706198
rect 576918 705642 577154 705878
rect 576918 696325 577154 696561
rect 576918 689325 577154 689561
rect 576918 682325 577154 682561
rect 576918 675325 577154 675561
rect 576918 668325 577154 668561
rect 576918 661325 577154 661561
rect 576918 654325 577154 654561
rect 576918 647325 577154 647561
rect 576918 640325 577154 640561
rect 576918 633325 577154 633561
rect 576918 626325 577154 626561
rect 576918 619325 577154 619561
rect 576918 612325 577154 612561
rect 576918 605325 577154 605561
rect 576918 598325 577154 598561
rect 576918 591325 577154 591561
rect 576918 584325 577154 584561
rect 576918 577325 577154 577561
rect 576918 570325 577154 570561
rect 576918 563325 577154 563561
rect 576918 556325 577154 556561
rect 576918 549325 577154 549561
rect 576918 542325 577154 542561
rect 576918 535325 577154 535561
rect 576918 528325 577154 528561
rect 576918 521325 577154 521561
rect 576918 514325 577154 514561
rect 576918 507325 577154 507561
rect 576918 500325 577154 500561
rect 576918 493325 577154 493561
rect 576918 486325 577154 486561
rect 576918 479325 577154 479561
rect 576918 472325 577154 472561
rect 576918 465325 577154 465561
rect 576918 458325 577154 458561
rect 576918 451325 577154 451561
rect 576918 444325 577154 444561
rect 576918 437325 577154 437561
rect 576918 430325 577154 430561
rect 576918 423325 577154 423561
rect 576918 416325 577154 416561
rect 576918 409325 577154 409561
rect 576918 402325 577154 402561
rect 576918 395325 577154 395561
rect 576918 388325 577154 388561
rect 576918 381325 577154 381561
rect 576918 374325 577154 374561
rect 576918 367325 577154 367561
rect 576918 360325 577154 360561
rect 576918 353325 577154 353561
rect 576918 346325 577154 346561
rect 576918 339325 577154 339561
rect 576918 332325 577154 332561
rect 576918 325325 577154 325561
rect 576918 318325 577154 318561
rect 576918 311325 577154 311561
rect 576918 304325 577154 304561
rect 576918 297325 577154 297561
rect 576918 290325 577154 290561
rect 576918 283325 577154 283561
rect 576918 276325 577154 276561
rect 576918 269325 577154 269561
rect 576918 262325 577154 262561
rect 576918 255325 577154 255561
rect 576918 248325 577154 248561
rect 576918 241325 577154 241561
rect 576918 234325 577154 234561
rect 576918 227325 577154 227561
rect 576918 220325 577154 220561
rect 576918 213325 577154 213561
rect 576918 206325 577154 206561
rect 576918 199325 577154 199561
rect 576918 192325 577154 192561
rect 576918 185325 577154 185561
rect 576918 178325 577154 178561
rect 576918 171325 577154 171561
rect 576918 164325 577154 164561
rect 576918 157325 577154 157561
rect 576918 150325 577154 150561
rect 576918 143325 577154 143561
rect 576918 136325 577154 136561
rect 576918 129325 577154 129561
rect 576918 122325 577154 122561
rect 576918 115325 577154 115561
rect 576918 108325 577154 108561
rect 576918 101325 577154 101561
rect 576918 94325 577154 94561
rect 576918 87325 577154 87561
rect 576918 80325 577154 80561
rect 576918 73325 577154 73561
rect 576918 66325 577154 66561
rect 576918 59325 577154 59561
rect 576918 52325 577154 52561
rect 576918 45325 577154 45561
rect 576918 38325 577154 38561
rect 576918 31325 577154 31561
rect 576918 24325 577154 24561
rect 576918 17325 577154 17561
rect 576918 10325 577154 10561
rect 576918 3325 577154 3561
rect 576918 -1942 577154 -1706
rect 576918 -2262 577154 -2026
rect 582186 705002 582422 705238
rect 582186 704682 582422 704918
rect 582186 695258 582422 695494
rect 582186 688258 582422 688494
rect 582186 681258 582422 681494
rect 582186 674258 582422 674494
rect 582186 667258 582422 667494
rect 582186 660258 582422 660494
rect 582186 653258 582422 653494
rect 582186 646258 582422 646494
rect 582186 639258 582422 639494
rect 582186 632258 582422 632494
rect 582186 625258 582422 625494
rect 582186 618258 582422 618494
rect 582186 611258 582422 611494
rect 582186 604258 582422 604494
rect 582186 597258 582422 597494
rect 582186 590258 582422 590494
rect 582186 583258 582422 583494
rect 582186 576258 582422 576494
rect 582186 569258 582422 569494
rect 582186 562258 582422 562494
rect 582186 555258 582422 555494
rect 582186 548258 582422 548494
rect 582186 541258 582422 541494
rect 582186 534258 582422 534494
rect 582186 527258 582422 527494
rect 582186 520258 582422 520494
rect 582186 513258 582422 513494
rect 582186 506258 582422 506494
rect 582186 499258 582422 499494
rect 582186 492258 582422 492494
rect 582186 485258 582422 485494
rect 582186 478258 582422 478494
rect 582186 471258 582422 471494
rect 582186 464258 582422 464494
rect 582186 457258 582422 457494
rect 582186 450258 582422 450494
rect 582186 443258 582422 443494
rect 582186 436258 582422 436494
rect 582186 429258 582422 429494
rect 582186 422258 582422 422494
rect 582186 415258 582422 415494
rect 582186 408258 582422 408494
rect 582186 401258 582422 401494
rect 582186 394258 582422 394494
rect 582186 387258 582422 387494
rect 582186 380258 582422 380494
rect 582186 373258 582422 373494
rect 582186 366258 582422 366494
rect 582186 359258 582422 359494
rect 582186 352258 582422 352494
rect 582186 345258 582422 345494
rect 582186 338258 582422 338494
rect 582186 331258 582422 331494
rect 582186 324258 582422 324494
rect 582186 317258 582422 317494
rect 582186 310258 582422 310494
rect 582186 303258 582422 303494
rect 582186 296258 582422 296494
rect 582186 289258 582422 289494
rect 582186 282258 582422 282494
rect 582186 275258 582422 275494
rect 582186 268258 582422 268494
rect 582186 261258 582422 261494
rect 582186 254258 582422 254494
rect 582186 247258 582422 247494
rect 582186 240258 582422 240494
rect 582186 233258 582422 233494
rect 582186 226258 582422 226494
rect 582186 219258 582422 219494
rect 582186 212258 582422 212494
rect 582186 205258 582422 205494
rect 582186 198258 582422 198494
rect 582186 191258 582422 191494
rect 582186 184258 582422 184494
rect 582186 177258 582422 177494
rect 582186 170258 582422 170494
rect 582186 163258 582422 163494
rect 582186 156258 582422 156494
rect 582186 149258 582422 149494
rect 582186 142258 582422 142494
rect 582186 135258 582422 135494
rect 582186 128258 582422 128494
rect 582186 121258 582422 121494
rect 582186 114258 582422 114494
rect 582186 107258 582422 107494
rect 582186 100258 582422 100494
rect 582186 93258 582422 93494
rect 582186 86258 582422 86494
rect 582186 79258 582422 79494
rect 582186 72258 582422 72494
rect 582186 65258 582422 65494
rect 582186 58258 582422 58494
rect 582186 51258 582422 51494
rect 582186 44258 582422 44494
rect 582186 37258 582422 37494
rect 582186 30258 582422 30494
rect 582186 23258 582422 23494
rect 582186 16258 582422 16494
rect 582186 9258 582422 9494
rect 582186 2258 582422 2494
rect 582186 -982 582422 -746
rect 582186 -1302 582422 -1066
rect 585818 705002 586054 705238
rect 586138 705002 586374 705238
rect 586458 705002 586694 705238
rect 586778 705002 587014 705238
rect 585818 704682 586054 704918
rect 586138 704682 586374 704918
rect 586458 704682 586694 704918
rect 586778 704682 587014 704918
rect 585818 695258 586054 695494
rect 586138 695258 586374 695494
rect 586458 695258 586694 695494
rect 586778 695258 587014 695494
rect 585818 688258 586054 688494
rect 586138 688258 586374 688494
rect 586458 688258 586694 688494
rect 586778 688258 587014 688494
rect 585818 681258 586054 681494
rect 586138 681258 586374 681494
rect 586458 681258 586694 681494
rect 586778 681258 587014 681494
rect 585818 674258 586054 674494
rect 586138 674258 586374 674494
rect 586458 674258 586694 674494
rect 586778 674258 587014 674494
rect 585818 667258 586054 667494
rect 586138 667258 586374 667494
rect 586458 667258 586694 667494
rect 586778 667258 587014 667494
rect 585818 660258 586054 660494
rect 586138 660258 586374 660494
rect 586458 660258 586694 660494
rect 586778 660258 587014 660494
rect 585818 653258 586054 653494
rect 586138 653258 586374 653494
rect 586458 653258 586694 653494
rect 586778 653258 587014 653494
rect 585818 646258 586054 646494
rect 586138 646258 586374 646494
rect 586458 646258 586694 646494
rect 586778 646258 587014 646494
rect 585818 639258 586054 639494
rect 586138 639258 586374 639494
rect 586458 639258 586694 639494
rect 586778 639258 587014 639494
rect 585818 632258 586054 632494
rect 586138 632258 586374 632494
rect 586458 632258 586694 632494
rect 586778 632258 587014 632494
rect 585818 625258 586054 625494
rect 586138 625258 586374 625494
rect 586458 625258 586694 625494
rect 586778 625258 587014 625494
rect 585818 618258 586054 618494
rect 586138 618258 586374 618494
rect 586458 618258 586694 618494
rect 586778 618258 587014 618494
rect 585818 611258 586054 611494
rect 586138 611258 586374 611494
rect 586458 611258 586694 611494
rect 586778 611258 587014 611494
rect 585818 604258 586054 604494
rect 586138 604258 586374 604494
rect 586458 604258 586694 604494
rect 586778 604258 587014 604494
rect 585818 597258 586054 597494
rect 586138 597258 586374 597494
rect 586458 597258 586694 597494
rect 586778 597258 587014 597494
rect 585818 590258 586054 590494
rect 586138 590258 586374 590494
rect 586458 590258 586694 590494
rect 586778 590258 587014 590494
rect 585818 583258 586054 583494
rect 586138 583258 586374 583494
rect 586458 583258 586694 583494
rect 586778 583258 587014 583494
rect 585818 576258 586054 576494
rect 586138 576258 586374 576494
rect 586458 576258 586694 576494
rect 586778 576258 587014 576494
rect 585818 569258 586054 569494
rect 586138 569258 586374 569494
rect 586458 569258 586694 569494
rect 586778 569258 587014 569494
rect 585818 562258 586054 562494
rect 586138 562258 586374 562494
rect 586458 562258 586694 562494
rect 586778 562258 587014 562494
rect 585818 555258 586054 555494
rect 586138 555258 586374 555494
rect 586458 555258 586694 555494
rect 586778 555258 587014 555494
rect 585818 548258 586054 548494
rect 586138 548258 586374 548494
rect 586458 548258 586694 548494
rect 586778 548258 587014 548494
rect 585818 541258 586054 541494
rect 586138 541258 586374 541494
rect 586458 541258 586694 541494
rect 586778 541258 587014 541494
rect 585818 534258 586054 534494
rect 586138 534258 586374 534494
rect 586458 534258 586694 534494
rect 586778 534258 587014 534494
rect 585818 527258 586054 527494
rect 586138 527258 586374 527494
rect 586458 527258 586694 527494
rect 586778 527258 587014 527494
rect 585818 520258 586054 520494
rect 586138 520258 586374 520494
rect 586458 520258 586694 520494
rect 586778 520258 587014 520494
rect 585818 513258 586054 513494
rect 586138 513258 586374 513494
rect 586458 513258 586694 513494
rect 586778 513258 587014 513494
rect 585818 506258 586054 506494
rect 586138 506258 586374 506494
rect 586458 506258 586694 506494
rect 586778 506258 587014 506494
rect 585818 499258 586054 499494
rect 586138 499258 586374 499494
rect 586458 499258 586694 499494
rect 586778 499258 587014 499494
rect 585818 492258 586054 492494
rect 586138 492258 586374 492494
rect 586458 492258 586694 492494
rect 586778 492258 587014 492494
rect 585818 485258 586054 485494
rect 586138 485258 586374 485494
rect 586458 485258 586694 485494
rect 586778 485258 587014 485494
rect 585818 478258 586054 478494
rect 586138 478258 586374 478494
rect 586458 478258 586694 478494
rect 586778 478258 587014 478494
rect 585818 471258 586054 471494
rect 586138 471258 586374 471494
rect 586458 471258 586694 471494
rect 586778 471258 587014 471494
rect 585818 464258 586054 464494
rect 586138 464258 586374 464494
rect 586458 464258 586694 464494
rect 586778 464258 587014 464494
rect 585818 457258 586054 457494
rect 586138 457258 586374 457494
rect 586458 457258 586694 457494
rect 586778 457258 587014 457494
rect 585818 450258 586054 450494
rect 586138 450258 586374 450494
rect 586458 450258 586694 450494
rect 586778 450258 587014 450494
rect 585818 443258 586054 443494
rect 586138 443258 586374 443494
rect 586458 443258 586694 443494
rect 586778 443258 587014 443494
rect 585818 436258 586054 436494
rect 586138 436258 586374 436494
rect 586458 436258 586694 436494
rect 586778 436258 587014 436494
rect 585818 429258 586054 429494
rect 586138 429258 586374 429494
rect 586458 429258 586694 429494
rect 586778 429258 587014 429494
rect 585818 422258 586054 422494
rect 586138 422258 586374 422494
rect 586458 422258 586694 422494
rect 586778 422258 587014 422494
rect 585818 415258 586054 415494
rect 586138 415258 586374 415494
rect 586458 415258 586694 415494
rect 586778 415258 587014 415494
rect 585818 408258 586054 408494
rect 586138 408258 586374 408494
rect 586458 408258 586694 408494
rect 586778 408258 587014 408494
rect 585818 401258 586054 401494
rect 586138 401258 586374 401494
rect 586458 401258 586694 401494
rect 586778 401258 587014 401494
rect 585818 394258 586054 394494
rect 586138 394258 586374 394494
rect 586458 394258 586694 394494
rect 586778 394258 587014 394494
rect 585818 387258 586054 387494
rect 586138 387258 586374 387494
rect 586458 387258 586694 387494
rect 586778 387258 587014 387494
rect 585818 380258 586054 380494
rect 586138 380258 586374 380494
rect 586458 380258 586694 380494
rect 586778 380258 587014 380494
rect 585818 373258 586054 373494
rect 586138 373258 586374 373494
rect 586458 373258 586694 373494
rect 586778 373258 587014 373494
rect 585818 366258 586054 366494
rect 586138 366258 586374 366494
rect 586458 366258 586694 366494
rect 586778 366258 587014 366494
rect 585818 359258 586054 359494
rect 586138 359258 586374 359494
rect 586458 359258 586694 359494
rect 586778 359258 587014 359494
rect 585818 352258 586054 352494
rect 586138 352258 586374 352494
rect 586458 352258 586694 352494
rect 586778 352258 587014 352494
rect 585818 345258 586054 345494
rect 586138 345258 586374 345494
rect 586458 345258 586694 345494
rect 586778 345258 587014 345494
rect 585818 338258 586054 338494
rect 586138 338258 586374 338494
rect 586458 338258 586694 338494
rect 586778 338258 587014 338494
rect 585818 331258 586054 331494
rect 586138 331258 586374 331494
rect 586458 331258 586694 331494
rect 586778 331258 587014 331494
rect 585818 324258 586054 324494
rect 586138 324258 586374 324494
rect 586458 324258 586694 324494
rect 586778 324258 587014 324494
rect 585818 317258 586054 317494
rect 586138 317258 586374 317494
rect 586458 317258 586694 317494
rect 586778 317258 587014 317494
rect 585818 310258 586054 310494
rect 586138 310258 586374 310494
rect 586458 310258 586694 310494
rect 586778 310258 587014 310494
rect 585818 303258 586054 303494
rect 586138 303258 586374 303494
rect 586458 303258 586694 303494
rect 586778 303258 587014 303494
rect 585818 296258 586054 296494
rect 586138 296258 586374 296494
rect 586458 296258 586694 296494
rect 586778 296258 587014 296494
rect 585818 289258 586054 289494
rect 586138 289258 586374 289494
rect 586458 289258 586694 289494
rect 586778 289258 587014 289494
rect 585818 282258 586054 282494
rect 586138 282258 586374 282494
rect 586458 282258 586694 282494
rect 586778 282258 587014 282494
rect 585818 275258 586054 275494
rect 586138 275258 586374 275494
rect 586458 275258 586694 275494
rect 586778 275258 587014 275494
rect 585818 268258 586054 268494
rect 586138 268258 586374 268494
rect 586458 268258 586694 268494
rect 586778 268258 587014 268494
rect 585818 261258 586054 261494
rect 586138 261258 586374 261494
rect 586458 261258 586694 261494
rect 586778 261258 587014 261494
rect 585818 254258 586054 254494
rect 586138 254258 586374 254494
rect 586458 254258 586694 254494
rect 586778 254258 587014 254494
rect 585818 247258 586054 247494
rect 586138 247258 586374 247494
rect 586458 247258 586694 247494
rect 586778 247258 587014 247494
rect 585818 240258 586054 240494
rect 586138 240258 586374 240494
rect 586458 240258 586694 240494
rect 586778 240258 587014 240494
rect 585818 233258 586054 233494
rect 586138 233258 586374 233494
rect 586458 233258 586694 233494
rect 586778 233258 587014 233494
rect 585818 226258 586054 226494
rect 586138 226258 586374 226494
rect 586458 226258 586694 226494
rect 586778 226258 587014 226494
rect 585818 219258 586054 219494
rect 586138 219258 586374 219494
rect 586458 219258 586694 219494
rect 586778 219258 587014 219494
rect 585818 212258 586054 212494
rect 586138 212258 586374 212494
rect 586458 212258 586694 212494
rect 586778 212258 587014 212494
rect 585818 205258 586054 205494
rect 586138 205258 586374 205494
rect 586458 205258 586694 205494
rect 586778 205258 587014 205494
rect 585818 198258 586054 198494
rect 586138 198258 586374 198494
rect 586458 198258 586694 198494
rect 586778 198258 587014 198494
rect 585818 191258 586054 191494
rect 586138 191258 586374 191494
rect 586458 191258 586694 191494
rect 586778 191258 587014 191494
rect 585818 184258 586054 184494
rect 586138 184258 586374 184494
rect 586458 184258 586694 184494
rect 586778 184258 587014 184494
rect 585818 177258 586054 177494
rect 586138 177258 586374 177494
rect 586458 177258 586694 177494
rect 586778 177258 587014 177494
rect 585818 170258 586054 170494
rect 586138 170258 586374 170494
rect 586458 170258 586694 170494
rect 586778 170258 587014 170494
rect 585818 163258 586054 163494
rect 586138 163258 586374 163494
rect 586458 163258 586694 163494
rect 586778 163258 587014 163494
rect 585818 156258 586054 156494
rect 586138 156258 586374 156494
rect 586458 156258 586694 156494
rect 586778 156258 587014 156494
rect 585818 149258 586054 149494
rect 586138 149258 586374 149494
rect 586458 149258 586694 149494
rect 586778 149258 587014 149494
rect 585818 142258 586054 142494
rect 586138 142258 586374 142494
rect 586458 142258 586694 142494
rect 586778 142258 587014 142494
rect 585818 135258 586054 135494
rect 586138 135258 586374 135494
rect 586458 135258 586694 135494
rect 586778 135258 587014 135494
rect 585818 128258 586054 128494
rect 586138 128258 586374 128494
rect 586458 128258 586694 128494
rect 586778 128258 587014 128494
rect 585818 121258 586054 121494
rect 586138 121258 586374 121494
rect 586458 121258 586694 121494
rect 586778 121258 587014 121494
rect 585818 114258 586054 114494
rect 586138 114258 586374 114494
rect 586458 114258 586694 114494
rect 586778 114258 587014 114494
rect 585818 107258 586054 107494
rect 586138 107258 586374 107494
rect 586458 107258 586694 107494
rect 586778 107258 587014 107494
rect 585818 100258 586054 100494
rect 586138 100258 586374 100494
rect 586458 100258 586694 100494
rect 586778 100258 587014 100494
rect 585818 93258 586054 93494
rect 586138 93258 586374 93494
rect 586458 93258 586694 93494
rect 586778 93258 587014 93494
rect 585818 86258 586054 86494
rect 586138 86258 586374 86494
rect 586458 86258 586694 86494
rect 586778 86258 587014 86494
rect 585818 79258 586054 79494
rect 586138 79258 586374 79494
rect 586458 79258 586694 79494
rect 586778 79258 587014 79494
rect 585818 72258 586054 72494
rect 586138 72258 586374 72494
rect 586458 72258 586694 72494
rect 586778 72258 587014 72494
rect 585818 65258 586054 65494
rect 586138 65258 586374 65494
rect 586458 65258 586694 65494
rect 586778 65258 587014 65494
rect 585818 58258 586054 58494
rect 586138 58258 586374 58494
rect 586458 58258 586694 58494
rect 586778 58258 587014 58494
rect 585818 51258 586054 51494
rect 586138 51258 586374 51494
rect 586458 51258 586694 51494
rect 586778 51258 587014 51494
rect 585818 44258 586054 44494
rect 586138 44258 586374 44494
rect 586458 44258 586694 44494
rect 586778 44258 587014 44494
rect 585818 37258 586054 37494
rect 586138 37258 586374 37494
rect 586458 37258 586694 37494
rect 586778 37258 587014 37494
rect 585818 30258 586054 30494
rect 586138 30258 586374 30494
rect 586458 30258 586694 30494
rect 586778 30258 587014 30494
rect 585818 23258 586054 23494
rect 586138 23258 586374 23494
rect 586458 23258 586694 23494
rect 586778 23258 587014 23494
rect 585818 16258 586054 16494
rect 586138 16258 586374 16494
rect 586458 16258 586694 16494
rect 586778 16258 587014 16494
rect 585818 9258 586054 9494
rect 586138 9258 586374 9494
rect 586458 9258 586694 9494
rect 586778 9258 587014 9494
rect 585818 2258 586054 2494
rect 586138 2258 586374 2494
rect 586458 2258 586694 2494
rect 586778 2258 587014 2494
rect 585818 -982 586054 -746
rect 586138 -982 586374 -746
rect 586458 -982 586694 -746
rect 586778 -982 587014 -746
rect 585818 -1302 586054 -1066
rect 586138 -1302 586374 -1066
rect 586458 -1302 586694 -1066
rect 586778 -1302 587014 -1066
rect 587570 696325 587806 696561
rect 587890 696325 588126 696561
rect 588210 696325 588446 696561
rect 588530 696325 588766 696561
rect 587570 689325 587806 689561
rect 587890 689325 588126 689561
rect 588210 689325 588446 689561
rect 588530 689325 588766 689561
rect 587570 682325 587806 682561
rect 587890 682325 588126 682561
rect 588210 682325 588446 682561
rect 588530 682325 588766 682561
rect 587570 675325 587806 675561
rect 587890 675325 588126 675561
rect 588210 675325 588446 675561
rect 588530 675325 588766 675561
rect 587570 668325 587806 668561
rect 587890 668325 588126 668561
rect 588210 668325 588446 668561
rect 588530 668325 588766 668561
rect 587570 661325 587806 661561
rect 587890 661325 588126 661561
rect 588210 661325 588446 661561
rect 588530 661325 588766 661561
rect 587570 654325 587806 654561
rect 587890 654325 588126 654561
rect 588210 654325 588446 654561
rect 588530 654325 588766 654561
rect 587570 647325 587806 647561
rect 587890 647325 588126 647561
rect 588210 647325 588446 647561
rect 588530 647325 588766 647561
rect 587570 640325 587806 640561
rect 587890 640325 588126 640561
rect 588210 640325 588446 640561
rect 588530 640325 588766 640561
rect 587570 633325 587806 633561
rect 587890 633325 588126 633561
rect 588210 633325 588446 633561
rect 588530 633325 588766 633561
rect 587570 626325 587806 626561
rect 587890 626325 588126 626561
rect 588210 626325 588446 626561
rect 588530 626325 588766 626561
rect 587570 619325 587806 619561
rect 587890 619325 588126 619561
rect 588210 619325 588446 619561
rect 588530 619325 588766 619561
rect 587570 612325 587806 612561
rect 587890 612325 588126 612561
rect 588210 612325 588446 612561
rect 588530 612325 588766 612561
rect 587570 605325 587806 605561
rect 587890 605325 588126 605561
rect 588210 605325 588446 605561
rect 588530 605325 588766 605561
rect 587570 598325 587806 598561
rect 587890 598325 588126 598561
rect 588210 598325 588446 598561
rect 588530 598325 588766 598561
rect 587570 591325 587806 591561
rect 587890 591325 588126 591561
rect 588210 591325 588446 591561
rect 588530 591325 588766 591561
rect 587570 584325 587806 584561
rect 587890 584325 588126 584561
rect 588210 584325 588446 584561
rect 588530 584325 588766 584561
rect 587570 577325 587806 577561
rect 587890 577325 588126 577561
rect 588210 577325 588446 577561
rect 588530 577325 588766 577561
rect 587570 570325 587806 570561
rect 587890 570325 588126 570561
rect 588210 570325 588446 570561
rect 588530 570325 588766 570561
rect 587570 563325 587806 563561
rect 587890 563325 588126 563561
rect 588210 563325 588446 563561
rect 588530 563325 588766 563561
rect 587570 556325 587806 556561
rect 587890 556325 588126 556561
rect 588210 556325 588446 556561
rect 588530 556325 588766 556561
rect 587570 549325 587806 549561
rect 587890 549325 588126 549561
rect 588210 549325 588446 549561
rect 588530 549325 588766 549561
rect 587570 542325 587806 542561
rect 587890 542325 588126 542561
rect 588210 542325 588446 542561
rect 588530 542325 588766 542561
rect 587570 535325 587806 535561
rect 587890 535325 588126 535561
rect 588210 535325 588446 535561
rect 588530 535325 588766 535561
rect 587570 528325 587806 528561
rect 587890 528325 588126 528561
rect 588210 528325 588446 528561
rect 588530 528325 588766 528561
rect 587570 521325 587806 521561
rect 587890 521325 588126 521561
rect 588210 521325 588446 521561
rect 588530 521325 588766 521561
rect 587570 514325 587806 514561
rect 587890 514325 588126 514561
rect 588210 514325 588446 514561
rect 588530 514325 588766 514561
rect 587570 507325 587806 507561
rect 587890 507325 588126 507561
rect 588210 507325 588446 507561
rect 588530 507325 588766 507561
rect 587570 500325 587806 500561
rect 587890 500325 588126 500561
rect 588210 500325 588446 500561
rect 588530 500325 588766 500561
rect 587570 493325 587806 493561
rect 587890 493325 588126 493561
rect 588210 493325 588446 493561
rect 588530 493325 588766 493561
rect 587570 486325 587806 486561
rect 587890 486325 588126 486561
rect 588210 486325 588446 486561
rect 588530 486325 588766 486561
rect 587570 479325 587806 479561
rect 587890 479325 588126 479561
rect 588210 479325 588446 479561
rect 588530 479325 588766 479561
rect 587570 472325 587806 472561
rect 587890 472325 588126 472561
rect 588210 472325 588446 472561
rect 588530 472325 588766 472561
rect 587570 465325 587806 465561
rect 587890 465325 588126 465561
rect 588210 465325 588446 465561
rect 588530 465325 588766 465561
rect 587570 458325 587806 458561
rect 587890 458325 588126 458561
rect 588210 458325 588446 458561
rect 588530 458325 588766 458561
rect 587570 451325 587806 451561
rect 587890 451325 588126 451561
rect 588210 451325 588446 451561
rect 588530 451325 588766 451561
rect 587570 444325 587806 444561
rect 587890 444325 588126 444561
rect 588210 444325 588446 444561
rect 588530 444325 588766 444561
rect 587570 437325 587806 437561
rect 587890 437325 588126 437561
rect 588210 437325 588446 437561
rect 588530 437325 588766 437561
rect 587570 430325 587806 430561
rect 587890 430325 588126 430561
rect 588210 430325 588446 430561
rect 588530 430325 588766 430561
rect 587570 423325 587806 423561
rect 587890 423325 588126 423561
rect 588210 423325 588446 423561
rect 588530 423325 588766 423561
rect 587570 416325 587806 416561
rect 587890 416325 588126 416561
rect 588210 416325 588446 416561
rect 588530 416325 588766 416561
rect 587570 409325 587806 409561
rect 587890 409325 588126 409561
rect 588210 409325 588446 409561
rect 588530 409325 588766 409561
rect 587570 402325 587806 402561
rect 587890 402325 588126 402561
rect 588210 402325 588446 402561
rect 588530 402325 588766 402561
rect 587570 395325 587806 395561
rect 587890 395325 588126 395561
rect 588210 395325 588446 395561
rect 588530 395325 588766 395561
rect 587570 388325 587806 388561
rect 587890 388325 588126 388561
rect 588210 388325 588446 388561
rect 588530 388325 588766 388561
rect 587570 381325 587806 381561
rect 587890 381325 588126 381561
rect 588210 381325 588446 381561
rect 588530 381325 588766 381561
rect 587570 374325 587806 374561
rect 587890 374325 588126 374561
rect 588210 374325 588446 374561
rect 588530 374325 588766 374561
rect 587570 367325 587806 367561
rect 587890 367325 588126 367561
rect 588210 367325 588446 367561
rect 588530 367325 588766 367561
rect 587570 360325 587806 360561
rect 587890 360325 588126 360561
rect 588210 360325 588446 360561
rect 588530 360325 588766 360561
rect 587570 353325 587806 353561
rect 587890 353325 588126 353561
rect 588210 353325 588446 353561
rect 588530 353325 588766 353561
rect 587570 346325 587806 346561
rect 587890 346325 588126 346561
rect 588210 346325 588446 346561
rect 588530 346325 588766 346561
rect 587570 339325 587806 339561
rect 587890 339325 588126 339561
rect 588210 339325 588446 339561
rect 588530 339325 588766 339561
rect 587570 332325 587806 332561
rect 587890 332325 588126 332561
rect 588210 332325 588446 332561
rect 588530 332325 588766 332561
rect 587570 325325 587806 325561
rect 587890 325325 588126 325561
rect 588210 325325 588446 325561
rect 588530 325325 588766 325561
rect 587570 318325 587806 318561
rect 587890 318325 588126 318561
rect 588210 318325 588446 318561
rect 588530 318325 588766 318561
rect 587570 311325 587806 311561
rect 587890 311325 588126 311561
rect 588210 311325 588446 311561
rect 588530 311325 588766 311561
rect 587570 304325 587806 304561
rect 587890 304325 588126 304561
rect 588210 304325 588446 304561
rect 588530 304325 588766 304561
rect 587570 297325 587806 297561
rect 587890 297325 588126 297561
rect 588210 297325 588446 297561
rect 588530 297325 588766 297561
rect 587570 290325 587806 290561
rect 587890 290325 588126 290561
rect 588210 290325 588446 290561
rect 588530 290325 588766 290561
rect 587570 283325 587806 283561
rect 587890 283325 588126 283561
rect 588210 283325 588446 283561
rect 588530 283325 588766 283561
rect 587570 276325 587806 276561
rect 587890 276325 588126 276561
rect 588210 276325 588446 276561
rect 588530 276325 588766 276561
rect 587570 269325 587806 269561
rect 587890 269325 588126 269561
rect 588210 269325 588446 269561
rect 588530 269325 588766 269561
rect 587570 262325 587806 262561
rect 587890 262325 588126 262561
rect 588210 262325 588446 262561
rect 588530 262325 588766 262561
rect 587570 255325 587806 255561
rect 587890 255325 588126 255561
rect 588210 255325 588446 255561
rect 588530 255325 588766 255561
rect 587570 248325 587806 248561
rect 587890 248325 588126 248561
rect 588210 248325 588446 248561
rect 588530 248325 588766 248561
rect 587570 241325 587806 241561
rect 587890 241325 588126 241561
rect 588210 241325 588446 241561
rect 588530 241325 588766 241561
rect 587570 234325 587806 234561
rect 587890 234325 588126 234561
rect 588210 234325 588446 234561
rect 588530 234325 588766 234561
rect 587570 227325 587806 227561
rect 587890 227325 588126 227561
rect 588210 227325 588446 227561
rect 588530 227325 588766 227561
rect 587570 220325 587806 220561
rect 587890 220325 588126 220561
rect 588210 220325 588446 220561
rect 588530 220325 588766 220561
rect 587570 213325 587806 213561
rect 587890 213325 588126 213561
rect 588210 213325 588446 213561
rect 588530 213325 588766 213561
rect 587570 206325 587806 206561
rect 587890 206325 588126 206561
rect 588210 206325 588446 206561
rect 588530 206325 588766 206561
rect 587570 199325 587806 199561
rect 587890 199325 588126 199561
rect 588210 199325 588446 199561
rect 588530 199325 588766 199561
rect 587570 192325 587806 192561
rect 587890 192325 588126 192561
rect 588210 192325 588446 192561
rect 588530 192325 588766 192561
rect 587570 185325 587806 185561
rect 587890 185325 588126 185561
rect 588210 185325 588446 185561
rect 588530 185325 588766 185561
rect 587570 178325 587806 178561
rect 587890 178325 588126 178561
rect 588210 178325 588446 178561
rect 588530 178325 588766 178561
rect 587570 171325 587806 171561
rect 587890 171325 588126 171561
rect 588210 171325 588446 171561
rect 588530 171325 588766 171561
rect 587570 164325 587806 164561
rect 587890 164325 588126 164561
rect 588210 164325 588446 164561
rect 588530 164325 588766 164561
rect 587570 157325 587806 157561
rect 587890 157325 588126 157561
rect 588210 157325 588446 157561
rect 588530 157325 588766 157561
rect 587570 150325 587806 150561
rect 587890 150325 588126 150561
rect 588210 150325 588446 150561
rect 588530 150325 588766 150561
rect 587570 143325 587806 143561
rect 587890 143325 588126 143561
rect 588210 143325 588446 143561
rect 588530 143325 588766 143561
rect 587570 136325 587806 136561
rect 587890 136325 588126 136561
rect 588210 136325 588446 136561
rect 588530 136325 588766 136561
rect 587570 129325 587806 129561
rect 587890 129325 588126 129561
rect 588210 129325 588446 129561
rect 588530 129325 588766 129561
rect 587570 122325 587806 122561
rect 587890 122325 588126 122561
rect 588210 122325 588446 122561
rect 588530 122325 588766 122561
rect 587570 115325 587806 115561
rect 587890 115325 588126 115561
rect 588210 115325 588446 115561
rect 588530 115325 588766 115561
rect 587570 108325 587806 108561
rect 587890 108325 588126 108561
rect 588210 108325 588446 108561
rect 588530 108325 588766 108561
rect 587570 101325 587806 101561
rect 587890 101325 588126 101561
rect 588210 101325 588446 101561
rect 588530 101325 588766 101561
rect 587570 94325 587806 94561
rect 587890 94325 588126 94561
rect 588210 94325 588446 94561
rect 588530 94325 588766 94561
rect 587570 87325 587806 87561
rect 587890 87325 588126 87561
rect 588210 87325 588446 87561
rect 588530 87325 588766 87561
rect 587570 80325 587806 80561
rect 587890 80325 588126 80561
rect 588210 80325 588446 80561
rect 588530 80325 588766 80561
rect 587570 73325 587806 73561
rect 587890 73325 588126 73561
rect 588210 73325 588446 73561
rect 588530 73325 588766 73561
rect 587570 66325 587806 66561
rect 587890 66325 588126 66561
rect 588210 66325 588446 66561
rect 588530 66325 588766 66561
rect 587570 59325 587806 59561
rect 587890 59325 588126 59561
rect 588210 59325 588446 59561
rect 588530 59325 588766 59561
rect 587570 52325 587806 52561
rect 587890 52325 588126 52561
rect 588210 52325 588446 52561
rect 588530 52325 588766 52561
rect 587570 45325 587806 45561
rect 587890 45325 588126 45561
rect 588210 45325 588446 45561
rect 588530 45325 588766 45561
rect 587570 38325 587806 38561
rect 587890 38325 588126 38561
rect 588210 38325 588446 38561
rect 588530 38325 588766 38561
rect 587570 31325 587806 31561
rect 587890 31325 588126 31561
rect 588210 31325 588446 31561
rect 588530 31325 588766 31561
rect 587570 24325 587806 24561
rect 587890 24325 588126 24561
rect 588210 24325 588446 24561
rect 588530 24325 588766 24561
rect 587570 17325 587806 17561
rect 587890 17325 588126 17561
rect 588210 17325 588446 17561
rect 588530 17325 588766 17561
rect 587570 10325 587806 10561
rect 587890 10325 588126 10561
rect 588210 10325 588446 10561
rect 588530 10325 588766 10561
rect 587570 3325 587806 3561
rect 587890 3325 588126 3561
rect 588210 3325 588446 3561
rect 588530 3325 588766 3561
<< metal5 >>
rect -3366 706198 587290 706230
rect -3366 705962 2918 706198
rect 3154 705962 9918 706198
rect 10154 705962 16918 706198
rect 17154 705962 23918 706198
rect 24154 705962 30918 706198
rect 31154 705962 37918 706198
rect 38154 705962 44918 706198
rect 45154 705962 51918 706198
rect 52154 705962 58918 706198
rect 59154 705962 65918 706198
rect 66154 705962 72918 706198
rect 73154 705962 79918 706198
rect 80154 705962 86918 706198
rect 87154 705962 93918 706198
rect 94154 705962 100918 706198
rect 101154 705962 107918 706198
rect 108154 705962 114918 706198
rect 115154 705962 121918 706198
rect 122154 705962 128918 706198
rect 129154 705962 135918 706198
rect 136154 705962 142918 706198
rect 143154 705962 149918 706198
rect 150154 705962 156918 706198
rect 157154 705962 163918 706198
rect 164154 705962 170918 706198
rect 171154 705962 177918 706198
rect 178154 705962 184918 706198
rect 185154 705962 191918 706198
rect 192154 705962 198918 706198
rect 199154 705962 205918 706198
rect 206154 705962 212918 706198
rect 213154 705962 219918 706198
rect 220154 705962 226918 706198
rect 227154 705962 233918 706198
rect 234154 705962 240918 706198
rect 241154 705962 247918 706198
rect 248154 705962 254918 706198
rect 255154 705962 261918 706198
rect 262154 705962 268918 706198
rect 269154 705962 275918 706198
rect 276154 705962 282918 706198
rect 283154 705962 289918 706198
rect 290154 705962 296918 706198
rect 297154 705962 303918 706198
rect 304154 705962 310918 706198
rect 311154 705962 317918 706198
rect 318154 705962 324918 706198
rect 325154 705962 331918 706198
rect 332154 705962 338918 706198
rect 339154 705962 345918 706198
rect 346154 705962 352918 706198
rect 353154 705962 359918 706198
rect 360154 705962 366918 706198
rect 367154 705962 373918 706198
rect 374154 705962 380918 706198
rect 381154 705962 387918 706198
rect 388154 705962 394918 706198
rect 395154 705962 401918 706198
rect 402154 705962 408918 706198
rect 409154 705962 415918 706198
rect 416154 705962 422918 706198
rect 423154 705962 429918 706198
rect 430154 705962 436918 706198
rect 437154 705962 443918 706198
rect 444154 705962 450918 706198
rect 451154 705962 457918 706198
rect 458154 705962 464918 706198
rect 465154 705962 471918 706198
rect 472154 705962 478918 706198
rect 479154 705962 485918 706198
rect 486154 705962 492918 706198
rect 493154 705962 499918 706198
rect 500154 705962 506918 706198
rect 507154 705962 513918 706198
rect 514154 705962 520918 706198
rect 521154 705962 527918 706198
rect 528154 705962 534918 706198
rect 535154 705962 541918 706198
rect 542154 705962 548918 706198
rect 549154 705962 555918 706198
rect 556154 705962 562918 706198
rect 563154 705962 569918 706198
rect 570154 705962 576918 706198
rect 577154 705962 587290 706198
rect -3366 705878 587290 705962
rect -3366 705642 2918 705878
rect 3154 705642 9918 705878
rect 10154 705642 16918 705878
rect 17154 705642 23918 705878
rect 24154 705642 30918 705878
rect 31154 705642 37918 705878
rect 38154 705642 44918 705878
rect 45154 705642 51918 705878
rect 52154 705642 58918 705878
rect 59154 705642 65918 705878
rect 66154 705642 72918 705878
rect 73154 705642 79918 705878
rect 80154 705642 86918 705878
rect 87154 705642 93918 705878
rect 94154 705642 100918 705878
rect 101154 705642 107918 705878
rect 108154 705642 114918 705878
rect 115154 705642 121918 705878
rect 122154 705642 128918 705878
rect 129154 705642 135918 705878
rect 136154 705642 142918 705878
rect 143154 705642 149918 705878
rect 150154 705642 156918 705878
rect 157154 705642 163918 705878
rect 164154 705642 170918 705878
rect 171154 705642 177918 705878
rect 178154 705642 184918 705878
rect 185154 705642 191918 705878
rect 192154 705642 198918 705878
rect 199154 705642 205918 705878
rect 206154 705642 212918 705878
rect 213154 705642 219918 705878
rect 220154 705642 226918 705878
rect 227154 705642 233918 705878
rect 234154 705642 240918 705878
rect 241154 705642 247918 705878
rect 248154 705642 254918 705878
rect 255154 705642 261918 705878
rect 262154 705642 268918 705878
rect 269154 705642 275918 705878
rect 276154 705642 282918 705878
rect 283154 705642 289918 705878
rect 290154 705642 296918 705878
rect 297154 705642 303918 705878
rect 304154 705642 310918 705878
rect 311154 705642 317918 705878
rect 318154 705642 324918 705878
rect 325154 705642 331918 705878
rect 332154 705642 338918 705878
rect 339154 705642 345918 705878
rect 346154 705642 352918 705878
rect 353154 705642 359918 705878
rect 360154 705642 366918 705878
rect 367154 705642 373918 705878
rect 374154 705642 380918 705878
rect 381154 705642 387918 705878
rect 388154 705642 394918 705878
rect 395154 705642 401918 705878
rect 402154 705642 408918 705878
rect 409154 705642 415918 705878
rect 416154 705642 422918 705878
rect 423154 705642 429918 705878
rect 430154 705642 436918 705878
rect 437154 705642 443918 705878
rect 444154 705642 450918 705878
rect 451154 705642 457918 705878
rect 458154 705642 464918 705878
rect 465154 705642 471918 705878
rect 472154 705642 478918 705878
rect 479154 705642 485918 705878
rect 486154 705642 492918 705878
rect 493154 705642 499918 705878
rect 500154 705642 506918 705878
rect 507154 705642 513918 705878
rect 514154 705642 520918 705878
rect 521154 705642 527918 705878
rect 528154 705642 534918 705878
rect 535154 705642 541918 705878
rect 542154 705642 548918 705878
rect 549154 705642 555918 705878
rect 556154 705642 562918 705878
rect 563154 705642 569918 705878
rect 570154 705642 576918 705878
rect 577154 705642 587290 705878
rect -3366 705610 587290 705642
rect -2406 705238 587122 705270
rect -2406 705002 -2374 705238
rect -2138 705002 -2054 705238
rect -1818 705002 1186 705238
rect 1422 705002 8186 705238
rect 8422 705002 15186 705238
rect 15422 705002 22186 705238
rect 22422 705002 29186 705238
rect 29422 705002 36186 705238
rect 36422 705002 43186 705238
rect 43422 705002 50186 705238
rect 50422 705002 57186 705238
rect 57422 705002 64186 705238
rect 64422 705002 71186 705238
rect 71422 705002 78186 705238
rect 78422 705002 85186 705238
rect 85422 705002 92186 705238
rect 92422 705002 99186 705238
rect 99422 705002 106186 705238
rect 106422 705002 113186 705238
rect 113422 705002 120186 705238
rect 120422 705002 127186 705238
rect 127422 705002 134186 705238
rect 134422 705002 141186 705238
rect 141422 705002 148186 705238
rect 148422 705002 155186 705238
rect 155422 705002 162186 705238
rect 162422 705002 169186 705238
rect 169422 705002 176186 705238
rect 176422 705002 183186 705238
rect 183422 705002 190186 705238
rect 190422 705002 197186 705238
rect 197422 705002 204186 705238
rect 204422 705002 211186 705238
rect 211422 705002 218186 705238
rect 218422 705002 225186 705238
rect 225422 705002 232186 705238
rect 232422 705002 239186 705238
rect 239422 705002 246186 705238
rect 246422 705002 253186 705238
rect 253422 705002 260186 705238
rect 260422 705002 267186 705238
rect 267422 705002 274186 705238
rect 274422 705002 281186 705238
rect 281422 705002 288186 705238
rect 288422 705002 295186 705238
rect 295422 705002 302186 705238
rect 302422 705002 309186 705238
rect 309422 705002 316186 705238
rect 316422 705002 323186 705238
rect 323422 705002 330186 705238
rect 330422 705002 337186 705238
rect 337422 705002 344186 705238
rect 344422 705002 351186 705238
rect 351422 705002 358186 705238
rect 358422 705002 365186 705238
rect 365422 705002 372186 705238
rect 372422 705002 379186 705238
rect 379422 705002 386186 705238
rect 386422 705002 393186 705238
rect 393422 705002 400186 705238
rect 400422 705002 407186 705238
rect 407422 705002 414186 705238
rect 414422 705002 421186 705238
rect 421422 705002 428186 705238
rect 428422 705002 435186 705238
rect 435422 705002 442186 705238
rect 442422 705002 449186 705238
rect 449422 705002 456186 705238
rect 456422 705002 463186 705238
rect 463422 705002 470186 705238
rect 470422 705002 477186 705238
rect 477422 705002 484186 705238
rect 484422 705002 491186 705238
rect 491422 705002 498186 705238
rect 498422 705002 505186 705238
rect 505422 705002 512186 705238
rect 512422 705002 519186 705238
rect 519422 705002 526186 705238
rect 526422 705002 533186 705238
rect 533422 705002 540186 705238
rect 540422 705002 547186 705238
rect 547422 705002 554186 705238
rect 554422 705002 561186 705238
rect 561422 705002 568186 705238
rect 568422 705002 575186 705238
rect 575422 705002 582186 705238
rect 582422 705002 585818 705238
rect 586054 705002 586138 705238
rect 586374 705002 586458 705238
rect 586694 705002 586778 705238
rect 587014 705002 587122 705238
rect -2406 704918 587122 705002
rect -2406 704682 -2374 704918
rect -2138 704682 -2054 704918
rect -1818 704682 1186 704918
rect 1422 704682 8186 704918
rect 8422 704682 15186 704918
rect 15422 704682 22186 704918
rect 22422 704682 29186 704918
rect 29422 704682 36186 704918
rect 36422 704682 43186 704918
rect 43422 704682 50186 704918
rect 50422 704682 57186 704918
rect 57422 704682 64186 704918
rect 64422 704682 71186 704918
rect 71422 704682 78186 704918
rect 78422 704682 85186 704918
rect 85422 704682 92186 704918
rect 92422 704682 99186 704918
rect 99422 704682 106186 704918
rect 106422 704682 113186 704918
rect 113422 704682 120186 704918
rect 120422 704682 127186 704918
rect 127422 704682 134186 704918
rect 134422 704682 141186 704918
rect 141422 704682 148186 704918
rect 148422 704682 155186 704918
rect 155422 704682 162186 704918
rect 162422 704682 169186 704918
rect 169422 704682 176186 704918
rect 176422 704682 183186 704918
rect 183422 704682 190186 704918
rect 190422 704682 197186 704918
rect 197422 704682 204186 704918
rect 204422 704682 211186 704918
rect 211422 704682 218186 704918
rect 218422 704682 225186 704918
rect 225422 704682 232186 704918
rect 232422 704682 239186 704918
rect 239422 704682 246186 704918
rect 246422 704682 253186 704918
rect 253422 704682 260186 704918
rect 260422 704682 267186 704918
rect 267422 704682 274186 704918
rect 274422 704682 281186 704918
rect 281422 704682 288186 704918
rect 288422 704682 295186 704918
rect 295422 704682 302186 704918
rect 302422 704682 309186 704918
rect 309422 704682 316186 704918
rect 316422 704682 323186 704918
rect 323422 704682 330186 704918
rect 330422 704682 337186 704918
rect 337422 704682 344186 704918
rect 344422 704682 351186 704918
rect 351422 704682 358186 704918
rect 358422 704682 365186 704918
rect 365422 704682 372186 704918
rect 372422 704682 379186 704918
rect 379422 704682 386186 704918
rect 386422 704682 393186 704918
rect 393422 704682 400186 704918
rect 400422 704682 407186 704918
rect 407422 704682 414186 704918
rect 414422 704682 421186 704918
rect 421422 704682 428186 704918
rect 428422 704682 435186 704918
rect 435422 704682 442186 704918
rect 442422 704682 449186 704918
rect 449422 704682 456186 704918
rect 456422 704682 463186 704918
rect 463422 704682 470186 704918
rect 470422 704682 477186 704918
rect 477422 704682 484186 704918
rect 484422 704682 491186 704918
rect 491422 704682 498186 704918
rect 498422 704682 505186 704918
rect 505422 704682 512186 704918
rect 512422 704682 519186 704918
rect 519422 704682 526186 704918
rect 526422 704682 533186 704918
rect 533422 704682 540186 704918
rect 540422 704682 547186 704918
rect 547422 704682 554186 704918
rect 554422 704682 561186 704918
rect 561422 704682 568186 704918
rect 568422 704682 575186 704918
rect 575422 704682 582186 704918
rect 582422 704682 585818 704918
rect 586054 704682 586138 704918
rect 586374 704682 586458 704918
rect 586694 704682 586778 704918
rect 587014 704682 587122 704918
rect -2406 704650 587122 704682
rect -4950 696561 588874 696603
rect -4950 696325 -4842 696561
rect -4606 696325 -4522 696561
rect -4286 696325 -4202 696561
rect -3966 696325 -3882 696561
rect -3646 696325 2918 696561
rect 3154 696325 9918 696561
rect 10154 696325 16918 696561
rect 17154 696325 23918 696561
rect 24154 696325 30918 696561
rect 31154 696325 37918 696561
rect 38154 696325 44918 696561
rect 45154 696325 51918 696561
rect 52154 696325 58918 696561
rect 59154 696325 65918 696561
rect 66154 696325 72918 696561
rect 73154 696325 79918 696561
rect 80154 696325 86918 696561
rect 87154 696325 93918 696561
rect 94154 696325 100918 696561
rect 101154 696325 107918 696561
rect 108154 696325 114918 696561
rect 115154 696325 121918 696561
rect 122154 696325 128918 696561
rect 129154 696325 135918 696561
rect 136154 696325 142918 696561
rect 143154 696325 149918 696561
rect 150154 696325 156918 696561
rect 157154 696325 163918 696561
rect 164154 696325 170918 696561
rect 171154 696325 177918 696561
rect 178154 696325 184918 696561
rect 185154 696325 191918 696561
rect 192154 696325 198918 696561
rect 199154 696325 205918 696561
rect 206154 696325 212918 696561
rect 213154 696325 219918 696561
rect 220154 696325 226918 696561
rect 227154 696325 233918 696561
rect 234154 696325 240918 696561
rect 241154 696325 247918 696561
rect 248154 696325 254918 696561
rect 255154 696325 261918 696561
rect 262154 696325 268918 696561
rect 269154 696325 275918 696561
rect 276154 696325 282918 696561
rect 283154 696325 289918 696561
rect 290154 696325 296918 696561
rect 297154 696325 303918 696561
rect 304154 696325 310918 696561
rect 311154 696325 317918 696561
rect 318154 696325 324918 696561
rect 325154 696325 331918 696561
rect 332154 696325 338918 696561
rect 339154 696325 345918 696561
rect 346154 696325 352918 696561
rect 353154 696325 359918 696561
rect 360154 696325 366918 696561
rect 367154 696325 373918 696561
rect 374154 696325 380918 696561
rect 381154 696325 387918 696561
rect 388154 696325 394918 696561
rect 395154 696325 401918 696561
rect 402154 696325 408918 696561
rect 409154 696325 415918 696561
rect 416154 696325 422918 696561
rect 423154 696325 429918 696561
rect 430154 696325 436918 696561
rect 437154 696325 443918 696561
rect 444154 696325 450918 696561
rect 451154 696325 457918 696561
rect 458154 696325 464918 696561
rect 465154 696325 471918 696561
rect 472154 696325 478918 696561
rect 479154 696325 485918 696561
rect 486154 696325 492918 696561
rect 493154 696325 499918 696561
rect 500154 696325 506918 696561
rect 507154 696325 513918 696561
rect 514154 696325 520918 696561
rect 521154 696325 527918 696561
rect 528154 696325 534918 696561
rect 535154 696325 541918 696561
rect 542154 696325 548918 696561
rect 549154 696325 555918 696561
rect 556154 696325 562918 696561
rect 563154 696325 569918 696561
rect 570154 696325 576918 696561
rect 577154 696325 587570 696561
rect 587806 696325 587890 696561
rect 588126 696325 588210 696561
rect 588446 696325 588530 696561
rect 588766 696325 588874 696561
rect -4950 696283 588874 696325
rect -4950 695494 588874 695536
rect -4950 695258 -3090 695494
rect -2854 695258 -2770 695494
rect -2534 695258 -2450 695494
rect -2214 695258 -2130 695494
rect -1894 695258 1186 695494
rect 1422 695258 8186 695494
rect 8422 695258 15186 695494
rect 15422 695258 22186 695494
rect 22422 695258 29186 695494
rect 29422 695258 36186 695494
rect 36422 695258 43186 695494
rect 43422 695258 50186 695494
rect 50422 695258 57186 695494
rect 57422 695258 64186 695494
rect 64422 695258 71186 695494
rect 71422 695258 78186 695494
rect 78422 695258 85186 695494
rect 85422 695258 92186 695494
rect 92422 695258 99186 695494
rect 99422 695258 106186 695494
rect 106422 695258 113186 695494
rect 113422 695258 120186 695494
rect 120422 695258 127186 695494
rect 127422 695258 134186 695494
rect 134422 695258 141186 695494
rect 141422 695258 148186 695494
rect 148422 695258 155186 695494
rect 155422 695258 162186 695494
rect 162422 695258 169186 695494
rect 169422 695258 176186 695494
rect 176422 695258 183186 695494
rect 183422 695258 190186 695494
rect 190422 695258 197186 695494
rect 197422 695258 204186 695494
rect 204422 695258 211186 695494
rect 211422 695258 218186 695494
rect 218422 695258 225186 695494
rect 225422 695258 232186 695494
rect 232422 695258 239186 695494
rect 239422 695258 246186 695494
rect 246422 695258 253186 695494
rect 253422 695258 260186 695494
rect 260422 695258 267186 695494
rect 267422 695258 274186 695494
rect 274422 695258 281186 695494
rect 281422 695258 288186 695494
rect 288422 695258 295186 695494
rect 295422 695258 302186 695494
rect 302422 695258 309186 695494
rect 309422 695258 316186 695494
rect 316422 695258 323186 695494
rect 323422 695258 330186 695494
rect 330422 695258 337186 695494
rect 337422 695258 344186 695494
rect 344422 695258 351186 695494
rect 351422 695258 358186 695494
rect 358422 695258 365186 695494
rect 365422 695258 372186 695494
rect 372422 695258 379186 695494
rect 379422 695258 386186 695494
rect 386422 695258 393186 695494
rect 393422 695258 400186 695494
rect 400422 695258 407186 695494
rect 407422 695258 414186 695494
rect 414422 695258 421186 695494
rect 421422 695258 428186 695494
rect 428422 695258 435186 695494
rect 435422 695258 442186 695494
rect 442422 695258 449186 695494
rect 449422 695258 456186 695494
rect 456422 695258 463186 695494
rect 463422 695258 470186 695494
rect 470422 695258 477186 695494
rect 477422 695258 484186 695494
rect 484422 695258 491186 695494
rect 491422 695258 498186 695494
rect 498422 695258 505186 695494
rect 505422 695258 512186 695494
rect 512422 695258 519186 695494
rect 519422 695258 526186 695494
rect 526422 695258 533186 695494
rect 533422 695258 540186 695494
rect 540422 695258 547186 695494
rect 547422 695258 554186 695494
rect 554422 695258 561186 695494
rect 561422 695258 568186 695494
rect 568422 695258 575186 695494
rect 575422 695258 582186 695494
rect 582422 695258 585818 695494
rect 586054 695258 586138 695494
rect 586374 695258 586458 695494
rect 586694 695258 586778 695494
rect 587014 695258 588874 695494
rect -4950 695216 588874 695258
rect -4950 689561 588874 689603
rect -4950 689325 -4842 689561
rect -4606 689325 -4522 689561
rect -4286 689325 -4202 689561
rect -3966 689325 -3882 689561
rect -3646 689325 2918 689561
rect 3154 689325 9918 689561
rect 10154 689325 16918 689561
rect 17154 689325 23918 689561
rect 24154 689325 30918 689561
rect 31154 689325 37918 689561
rect 38154 689325 44918 689561
rect 45154 689325 51918 689561
rect 52154 689325 58918 689561
rect 59154 689325 65918 689561
rect 66154 689325 72918 689561
rect 73154 689325 79918 689561
rect 80154 689325 86918 689561
rect 87154 689325 93918 689561
rect 94154 689325 100918 689561
rect 101154 689325 107918 689561
rect 108154 689325 114918 689561
rect 115154 689325 121918 689561
rect 122154 689325 128918 689561
rect 129154 689325 135918 689561
rect 136154 689325 142918 689561
rect 143154 689325 149918 689561
rect 150154 689325 156918 689561
rect 157154 689325 163918 689561
rect 164154 689325 170918 689561
rect 171154 689325 177918 689561
rect 178154 689325 184918 689561
rect 185154 689325 191918 689561
rect 192154 689325 198918 689561
rect 199154 689325 205918 689561
rect 206154 689325 212918 689561
rect 213154 689325 219918 689561
rect 220154 689325 226918 689561
rect 227154 689325 233918 689561
rect 234154 689325 240918 689561
rect 241154 689325 247918 689561
rect 248154 689325 254918 689561
rect 255154 689325 261918 689561
rect 262154 689325 268918 689561
rect 269154 689325 275918 689561
rect 276154 689325 282918 689561
rect 283154 689325 289918 689561
rect 290154 689325 296918 689561
rect 297154 689325 303918 689561
rect 304154 689325 310918 689561
rect 311154 689325 317918 689561
rect 318154 689325 324918 689561
rect 325154 689325 331918 689561
rect 332154 689325 338918 689561
rect 339154 689325 345918 689561
rect 346154 689325 352918 689561
rect 353154 689325 359918 689561
rect 360154 689325 366918 689561
rect 367154 689325 373918 689561
rect 374154 689325 380918 689561
rect 381154 689325 387918 689561
rect 388154 689325 394918 689561
rect 395154 689325 401918 689561
rect 402154 689325 408918 689561
rect 409154 689325 415918 689561
rect 416154 689325 422918 689561
rect 423154 689325 429918 689561
rect 430154 689325 436918 689561
rect 437154 689325 443918 689561
rect 444154 689325 450918 689561
rect 451154 689325 457918 689561
rect 458154 689325 464918 689561
rect 465154 689325 471918 689561
rect 472154 689325 478918 689561
rect 479154 689325 485918 689561
rect 486154 689325 492918 689561
rect 493154 689325 499918 689561
rect 500154 689325 506918 689561
rect 507154 689325 513918 689561
rect 514154 689325 520918 689561
rect 521154 689325 527918 689561
rect 528154 689325 534918 689561
rect 535154 689325 541918 689561
rect 542154 689325 548918 689561
rect 549154 689325 555918 689561
rect 556154 689325 562918 689561
rect 563154 689325 569918 689561
rect 570154 689325 576918 689561
rect 577154 689325 587570 689561
rect 587806 689325 587890 689561
rect 588126 689325 588210 689561
rect 588446 689325 588530 689561
rect 588766 689325 588874 689561
rect -4950 689283 588874 689325
rect -4950 688494 588874 688536
rect -4950 688258 -3090 688494
rect -2854 688258 -2770 688494
rect -2534 688258 -2450 688494
rect -2214 688258 -2130 688494
rect -1894 688258 1186 688494
rect 1422 688258 8186 688494
rect 8422 688258 15186 688494
rect 15422 688258 22186 688494
rect 22422 688258 29186 688494
rect 29422 688258 36186 688494
rect 36422 688258 43186 688494
rect 43422 688258 50186 688494
rect 50422 688258 57186 688494
rect 57422 688258 64186 688494
rect 64422 688258 71186 688494
rect 71422 688258 78186 688494
rect 78422 688258 85186 688494
rect 85422 688258 92186 688494
rect 92422 688258 99186 688494
rect 99422 688258 106186 688494
rect 106422 688258 113186 688494
rect 113422 688258 120186 688494
rect 120422 688258 127186 688494
rect 127422 688258 134186 688494
rect 134422 688258 141186 688494
rect 141422 688258 148186 688494
rect 148422 688258 155186 688494
rect 155422 688258 162186 688494
rect 162422 688258 169186 688494
rect 169422 688258 176186 688494
rect 176422 688258 183186 688494
rect 183422 688258 190186 688494
rect 190422 688258 197186 688494
rect 197422 688258 204186 688494
rect 204422 688258 211186 688494
rect 211422 688258 218186 688494
rect 218422 688258 225186 688494
rect 225422 688258 232186 688494
rect 232422 688258 239186 688494
rect 239422 688258 246186 688494
rect 246422 688258 253186 688494
rect 253422 688258 260186 688494
rect 260422 688258 267186 688494
rect 267422 688258 274186 688494
rect 274422 688258 281186 688494
rect 281422 688258 288186 688494
rect 288422 688258 295186 688494
rect 295422 688258 302186 688494
rect 302422 688258 309186 688494
rect 309422 688258 316186 688494
rect 316422 688258 323186 688494
rect 323422 688258 330186 688494
rect 330422 688258 337186 688494
rect 337422 688258 344186 688494
rect 344422 688258 351186 688494
rect 351422 688258 358186 688494
rect 358422 688258 365186 688494
rect 365422 688258 372186 688494
rect 372422 688258 379186 688494
rect 379422 688258 386186 688494
rect 386422 688258 393186 688494
rect 393422 688258 400186 688494
rect 400422 688258 407186 688494
rect 407422 688258 414186 688494
rect 414422 688258 421186 688494
rect 421422 688258 428186 688494
rect 428422 688258 435186 688494
rect 435422 688258 442186 688494
rect 442422 688258 449186 688494
rect 449422 688258 456186 688494
rect 456422 688258 463186 688494
rect 463422 688258 470186 688494
rect 470422 688258 477186 688494
rect 477422 688258 484186 688494
rect 484422 688258 491186 688494
rect 491422 688258 498186 688494
rect 498422 688258 505186 688494
rect 505422 688258 512186 688494
rect 512422 688258 519186 688494
rect 519422 688258 526186 688494
rect 526422 688258 533186 688494
rect 533422 688258 540186 688494
rect 540422 688258 547186 688494
rect 547422 688258 554186 688494
rect 554422 688258 561186 688494
rect 561422 688258 568186 688494
rect 568422 688258 575186 688494
rect 575422 688258 582186 688494
rect 582422 688258 585818 688494
rect 586054 688258 586138 688494
rect 586374 688258 586458 688494
rect 586694 688258 586778 688494
rect 587014 688258 588874 688494
rect -4950 688216 588874 688258
rect -4950 682561 588874 682603
rect -4950 682325 -4842 682561
rect -4606 682325 -4522 682561
rect -4286 682325 -4202 682561
rect -3966 682325 -3882 682561
rect -3646 682325 2918 682561
rect 3154 682325 9918 682561
rect 10154 682325 16918 682561
rect 17154 682325 23918 682561
rect 24154 682325 30918 682561
rect 31154 682325 37918 682561
rect 38154 682325 44918 682561
rect 45154 682325 51918 682561
rect 52154 682325 58918 682561
rect 59154 682325 65918 682561
rect 66154 682325 72918 682561
rect 73154 682325 79918 682561
rect 80154 682325 86918 682561
rect 87154 682325 93918 682561
rect 94154 682325 100918 682561
rect 101154 682325 107918 682561
rect 108154 682325 114918 682561
rect 115154 682325 121918 682561
rect 122154 682325 128918 682561
rect 129154 682325 135918 682561
rect 136154 682325 142918 682561
rect 143154 682325 149918 682561
rect 150154 682325 156918 682561
rect 157154 682325 163918 682561
rect 164154 682325 170918 682561
rect 171154 682325 177918 682561
rect 178154 682325 184918 682561
rect 185154 682325 191918 682561
rect 192154 682325 198918 682561
rect 199154 682325 205918 682561
rect 206154 682325 212918 682561
rect 213154 682325 219918 682561
rect 220154 682325 226918 682561
rect 227154 682325 233918 682561
rect 234154 682325 240918 682561
rect 241154 682325 247918 682561
rect 248154 682325 254918 682561
rect 255154 682325 261918 682561
rect 262154 682325 268918 682561
rect 269154 682325 275918 682561
rect 276154 682325 282918 682561
rect 283154 682325 289918 682561
rect 290154 682325 296918 682561
rect 297154 682325 303918 682561
rect 304154 682325 310918 682561
rect 311154 682325 317918 682561
rect 318154 682325 324918 682561
rect 325154 682325 331918 682561
rect 332154 682325 338918 682561
rect 339154 682325 345918 682561
rect 346154 682325 352918 682561
rect 353154 682325 359918 682561
rect 360154 682325 366918 682561
rect 367154 682325 373918 682561
rect 374154 682325 380918 682561
rect 381154 682325 387918 682561
rect 388154 682325 394918 682561
rect 395154 682325 401918 682561
rect 402154 682325 408918 682561
rect 409154 682325 415918 682561
rect 416154 682325 422918 682561
rect 423154 682325 429918 682561
rect 430154 682325 436918 682561
rect 437154 682325 443918 682561
rect 444154 682325 450918 682561
rect 451154 682325 457918 682561
rect 458154 682325 464918 682561
rect 465154 682325 471918 682561
rect 472154 682325 478918 682561
rect 479154 682325 485918 682561
rect 486154 682325 492918 682561
rect 493154 682325 499918 682561
rect 500154 682325 506918 682561
rect 507154 682325 513918 682561
rect 514154 682325 520918 682561
rect 521154 682325 527918 682561
rect 528154 682325 534918 682561
rect 535154 682325 541918 682561
rect 542154 682325 548918 682561
rect 549154 682325 555918 682561
rect 556154 682325 562918 682561
rect 563154 682325 569918 682561
rect 570154 682325 576918 682561
rect 577154 682325 587570 682561
rect 587806 682325 587890 682561
rect 588126 682325 588210 682561
rect 588446 682325 588530 682561
rect 588766 682325 588874 682561
rect -4950 682283 588874 682325
rect -4950 681494 588874 681536
rect -4950 681258 -3090 681494
rect -2854 681258 -2770 681494
rect -2534 681258 -2450 681494
rect -2214 681258 -2130 681494
rect -1894 681258 1186 681494
rect 1422 681258 8186 681494
rect 8422 681258 15186 681494
rect 15422 681258 22186 681494
rect 22422 681258 29186 681494
rect 29422 681258 36186 681494
rect 36422 681258 43186 681494
rect 43422 681258 50186 681494
rect 50422 681258 57186 681494
rect 57422 681258 64186 681494
rect 64422 681258 71186 681494
rect 71422 681258 78186 681494
rect 78422 681258 85186 681494
rect 85422 681258 92186 681494
rect 92422 681258 99186 681494
rect 99422 681258 106186 681494
rect 106422 681258 113186 681494
rect 113422 681258 120186 681494
rect 120422 681258 127186 681494
rect 127422 681258 134186 681494
rect 134422 681258 141186 681494
rect 141422 681258 148186 681494
rect 148422 681258 155186 681494
rect 155422 681258 162186 681494
rect 162422 681258 169186 681494
rect 169422 681258 176186 681494
rect 176422 681258 183186 681494
rect 183422 681258 190186 681494
rect 190422 681258 197186 681494
rect 197422 681258 204186 681494
rect 204422 681258 211186 681494
rect 211422 681258 218186 681494
rect 218422 681258 225186 681494
rect 225422 681258 232186 681494
rect 232422 681258 239186 681494
rect 239422 681258 246186 681494
rect 246422 681258 253186 681494
rect 253422 681258 260186 681494
rect 260422 681258 267186 681494
rect 267422 681258 274186 681494
rect 274422 681258 281186 681494
rect 281422 681258 288186 681494
rect 288422 681258 295186 681494
rect 295422 681258 302186 681494
rect 302422 681258 309186 681494
rect 309422 681258 316186 681494
rect 316422 681258 323186 681494
rect 323422 681258 330186 681494
rect 330422 681258 337186 681494
rect 337422 681258 344186 681494
rect 344422 681258 351186 681494
rect 351422 681258 358186 681494
rect 358422 681258 365186 681494
rect 365422 681258 372186 681494
rect 372422 681258 379186 681494
rect 379422 681258 386186 681494
rect 386422 681258 393186 681494
rect 393422 681258 400186 681494
rect 400422 681258 407186 681494
rect 407422 681258 414186 681494
rect 414422 681258 421186 681494
rect 421422 681258 428186 681494
rect 428422 681258 435186 681494
rect 435422 681258 442186 681494
rect 442422 681258 449186 681494
rect 449422 681258 456186 681494
rect 456422 681258 463186 681494
rect 463422 681258 470186 681494
rect 470422 681258 477186 681494
rect 477422 681258 484186 681494
rect 484422 681258 491186 681494
rect 491422 681258 498186 681494
rect 498422 681258 505186 681494
rect 505422 681258 512186 681494
rect 512422 681258 519186 681494
rect 519422 681258 526186 681494
rect 526422 681258 533186 681494
rect 533422 681258 540186 681494
rect 540422 681258 547186 681494
rect 547422 681258 554186 681494
rect 554422 681258 561186 681494
rect 561422 681258 568186 681494
rect 568422 681258 575186 681494
rect 575422 681258 582186 681494
rect 582422 681258 585818 681494
rect 586054 681258 586138 681494
rect 586374 681258 586458 681494
rect 586694 681258 586778 681494
rect 587014 681258 588874 681494
rect -4950 681216 588874 681258
rect -4950 675561 588874 675603
rect -4950 675325 -4842 675561
rect -4606 675325 -4522 675561
rect -4286 675325 -4202 675561
rect -3966 675325 -3882 675561
rect -3646 675325 2918 675561
rect 3154 675325 9918 675561
rect 10154 675325 16918 675561
rect 17154 675325 23918 675561
rect 24154 675325 30918 675561
rect 31154 675325 37918 675561
rect 38154 675325 44918 675561
rect 45154 675325 51918 675561
rect 52154 675325 58918 675561
rect 59154 675325 65918 675561
rect 66154 675325 72918 675561
rect 73154 675325 79918 675561
rect 80154 675325 86918 675561
rect 87154 675325 93918 675561
rect 94154 675325 100918 675561
rect 101154 675325 107918 675561
rect 108154 675325 114918 675561
rect 115154 675325 121918 675561
rect 122154 675325 128918 675561
rect 129154 675325 135918 675561
rect 136154 675325 142918 675561
rect 143154 675325 149918 675561
rect 150154 675325 156918 675561
rect 157154 675325 163918 675561
rect 164154 675325 170918 675561
rect 171154 675325 177918 675561
rect 178154 675325 184918 675561
rect 185154 675325 191918 675561
rect 192154 675325 198918 675561
rect 199154 675325 205918 675561
rect 206154 675325 212918 675561
rect 213154 675325 219918 675561
rect 220154 675325 226918 675561
rect 227154 675325 233918 675561
rect 234154 675325 240918 675561
rect 241154 675325 247918 675561
rect 248154 675325 254918 675561
rect 255154 675325 261918 675561
rect 262154 675325 268918 675561
rect 269154 675325 275918 675561
rect 276154 675325 282918 675561
rect 283154 675325 289918 675561
rect 290154 675325 296918 675561
rect 297154 675325 303918 675561
rect 304154 675325 310918 675561
rect 311154 675325 317918 675561
rect 318154 675325 324918 675561
rect 325154 675325 331918 675561
rect 332154 675325 338918 675561
rect 339154 675325 345918 675561
rect 346154 675325 352918 675561
rect 353154 675325 359918 675561
rect 360154 675325 366918 675561
rect 367154 675325 373918 675561
rect 374154 675325 380918 675561
rect 381154 675325 387918 675561
rect 388154 675325 394918 675561
rect 395154 675325 401918 675561
rect 402154 675325 408918 675561
rect 409154 675325 415918 675561
rect 416154 675325 422918 675561
rect 423154 675325 429918 675561
rect 430154 675325 436918 675561
rect 437154 675325 443918 675561
rect 444154 675325 450918 675561
rect 451154 675325 457918 675561
rect 458154 675325 464918 675561
rect 465154 675325 471918 675561
rect 472154 675325 478918 675561
rect 479154 675325 485918 675561
rect 486154 675325 492918 675561
rect 493154 675325 499918 675561
rect 500154 675325 506918 675561
rect 507154 675325 513918 675561
rect 514154 675325 520918 675561
rect 521154 675325 527918 675561
rect 528154 675325 534918 675561
rect 535154 675325 541918 675561
rect 542154 675325 548918 675561
rect 549154 675325 555918 675561
rect 556154 675325 562918 675561
rect 563154 675325 569918 675561
rect 570154 675325 576918 675561
rect 577154 675325 587570 675561
rect 587806 675325 587890 675561
rect 588126 675325 588210 675561
rect 588446 675325 588530 675561
rect 588766 675325 588874 675561
rect -4950 675283 588874 675325
rect -4950 674494 588874 674536
rect -4950 674258 -3090 674494
rect -2854 674258 -2770 674494
rect -2534 674258 -2450 674494
rect -2214 674258 -2130 674494
rect -1894 674258 1186 674494
rect 1422 674258 8186 674494
rect 8422 674258 15186 674494
rect 15422 674258 22186 674494
rect 22422 674258 29186 674494
rect 29422 674258 36186 674494
rect 36422 674258 43186 674494
rect 43422 674258 50186 674494
rect 50422 674258 57186 674494
rect 57422 674258 64186 674494
rect 64422 674258 71186 674494
rect 71422 674258 78186 674494
rect 78422 674258 85186 674494
rect 85422 674258 92186 674494
rect 92422 674258 99186 674494
rect 99422 674258 106186 674494
rect 106422 674258 113186 674494
rect 113422 674258 120186 674494
rect 120422 674258 127186 674494
rect 127422 674258 134186 674494
rect 134422 674258 141186 674494
rect 141422 674258 148186 674494
rect 148422 674258 155186 674494
rect 155422 674258 162186 674494
rect 162422 674258 169186 674494
rect 169422 674258 176186 674494
rect 176422 674258 183186 674494
rect 183422 674258 190186 674494
rect 190422 674258 197186 674494
rect 197422 674258 204186 674494
rect 204422 674258 211186 674494
rect 211422 674258 218186 674494
rect 218422 674258 225186 674494
rect 225422 674258 232186 674494
rect 232422 674258 239186 674494
rect 239422 674258 246186 674494
rect 246422 674258 253186 674494
rect 253422 674258 260186 674494
rect 260422 674258 267186 674494
rect 267422 674258 274186 674494
rect 274422 674258 281186 674494
rect 281422 674258 288186 674494
rect 288422 674258 295186 674494
rect 295422 674258 302186 674494
rect 302422 674258 309186 674494
rect 309422 674258 316186 674494
rect 316422 674258 323186 674494
rect 323422 674258 330186 674494
rect 330422 674258 337186 674494
rect 337422 674258 344186 674494
rect 344422 674258 351186 674494
rect 351422 674258 358186 674494
rect 358422 674258 365186 674494
rect 365422 674258 372186 674494
rect 372422 674258 379186 674494
rect 379422 674258 386186 674494
rect 386422 674258 393186 674494
rect 393422 674258 400186 674494
rect 400422 674258 407186 674494
rect 407422 674258 414186 674494
rect 414422 674258 421186 674494
rect 421422 674258 428186 674494
rect 428422 674258 435186 674494
rect 435422 674258 442186 674494
rect 442422 674258 449186 674494
rect 449422 674258 456186 674494
rect 456422 674258 463186 674494
rect 463422 674258 470186 674494
rect 470422 674258 477186 674494
rect 477422 674258 484186 674494
rect 484422 674258 491186 674494
rect 491422 674258 498186 674494
rect 498422 674258 505186 674494
rect 505422 674258 512186 674494
rect 512422 674258 519186 674494
rect 519422 674258 526186 674494
rect 526422 674258 533186 674494
rect 533422 674258 540186 674494
rect 540422 674258 547186 674494
rect 547422 674258 554186 674494
rect 554422 674258 561186 674494
rect 561422 674258 568186 674494
rect 568422 674258 575186 674494
rect 575422 674258 582186 674494
rect 582422 674258 585818 674494
rect 586054 674258 586138 674494
rect 586374 674258 586458 674494
rect 586694 674258 586778 674494
rect 587014 674258 588874 674494
rect -4950 674216 588874 674258
rect -4950 668561 588874 668603
rect -4950 668325 -4842 668561
rect -4606 668325 -4522 668561
rect -4286 668325 -4202 668561
rect -3966 668325 -3882 668561
rect -3646 668325 2918 668561
rect 3154 668325 9918 668561
rect 10154 668325 16918 668561
rect 17154 668325 23918 668561
rect 24154 668325 30918 668561
rect 31154 668325 37918 668561
rect 38154 668325 44918 668561
rect 45154 668325 51918 668561
rect 52154 668325 58918 668561
rect 59154 668325 65918 668561
rect 66154 668325 72918 668561
rect 73154 668325 79918 668561
rect 80154 668325 86918 668561
rect 87154 668325 93918 668561
rect 94154 668325 100918 668561
rect 101154 668325 107918 668561
rect 108154 668325 114918 668561
rect 115154 668325 121918 668561
rect 122154 668325 128918 668561
rect 129154 668325 135918 668561
rect 136154 668325 142918 668561
rect 143154 668325 149918 668561
rect 150154 668325 156918 668561
rect 157154 668325 163918 668561
rect 164154 668325 170918 668561
rect 171154 668325 177918 668561
rect 178154 668325 184918 668561
rect 185154 668325 191918 668561
rect 192154 668325 198918 668561
rect 199154 668325 205918 668561
rect 206154 668325 212918 668561
rect 213154 668325 219918 668561
rect 220154 668325 226918 668561
rect 227154 668325 233918 668561
rect 234154 668325 240918 668561
rect 241154 668325 247918 668561
rect 248154 668325 254918 668561
rect 255154 668325 261918 668561
rect 262154 668325 268918 668561
rect 269154 668325 275918 668561
rect 276154 668325 282918 668561
rect 283154 668325 289918 668561
rect 290154 668325 296918 668561
rect 297154 668325 303918 668561
rect 304154 668325 310918 668561
rect 311154 668325 317918 668561
rect 318154 668325 324918 668561
rect 325154 668325 331918 668561
rect 332154 668325 338918 668561
rect 339154 668325 345918 668561
rect 346154 668325 352918 668561
rect 353154 668325 359918 668561
rect 360154 668325 366918 668561
rect 367154 668325 373918 668561
rect 374154 668325 380918 668561
rect 381154 668325 387918 668561
rect 388154 668325 394918 668561
rect 395154 668325 401918 668561
rect 402154 668325 408918 668561
rect 409154 668325 415918 668561
rect 416154 668325 422918 668561
rect 423154 668325 429918 668561
rect 430154 668325 436918 668561
rect 437154 668325 443918 668561
rect 444154 668325 450918 668561
rect 451154 668325 457918 668561
rect 458154 668325 464918 668561
rect 465154 668325 471918 668561
rect 472154 668325 478918 668561
rect 479154 668325 485918 668561
rect 486154 668325 492918 668561
rect 493154 668325 499918 668561
rect 500154 668325 506918 668561
rect 507154 668325 513918 668561
rect 514154 668325 520918 668561
rect 521154 668325 527918 668561
rect 528154 668325 534918 668561
rect 535154 668325 541918 668561
rect 542154 668325 548918 668561
rect 549154 668325 555918 668561
rect 556154 668325 562918 668561
rect 563154 668325 569918 668561
rect 570154 668325 576918 668561
rect 577154 668325 587570 668561
rect 587806 668325 587890 668561
rect 588126 668325 588210 668561
rect 588446 668325 588530 668561
rect 588766 668325 588874 668561
rect -4950 668283 588874 668325
rect -4950 667494 588874 667536
rect -4950 667258 -3090 667494
rect -2854 667258 -2770 667494
rect -2534 667258 -2450 667494
rect -2214 667258 -2130 667494
rect -1894 667258 1186 667494
rect 1422 667258 8186 667494
rect 8422 667258 15186 667494
rect 15422 667258 22186 667494
rect 22422 667258 29186 667494
rect 29422 667258 36186 667494
rect 36422 667258 43186 667494
rect 43422 667258 50186 667494
rect 50422 667258 57186 667494
rect 57422 667258 64186 667494
rect 64422 667258 71186 667494
rect 71422 667258 78186 667494
rect 78422 667258 85186 667494
rect 85422 667258 92186 667494
rect 92422 667258 99186 667494
rect 99422 667258 106186 667494
rect 106422 667258 113186 667494
rect 113422 667258 120186 667494
rect 120422 667258 127186 667494
rect 127422 667258 134186 667494
rect 134422 667258 141186 667494
rect 141422 667258 148186 667494
rect 148422 667258 155186 667494
rect 155422 667258 162186 667494
rect 162422 667258 169186 667494
rect 169422 667258 176186 667494
rect 176422 667258 183186 667494
rect 183422 667258 190186 667494
rect 190422 667258 197186 667494
rect 197422 667258 204186 667494
rect 204422 667258 211186 667494
rect 211422 667258 218186 667494
rect 218422 667258 225186 667494
rect 225422 667258 232186 667494
rect 232422 667258 239186 667494
rect 239422 667258 246186 667494
rect 246422 667258 253186 667494
rect 253422 667258 260186 667494
rect 260422 667258 267186 667494
rect 267422 667258 274186 667494
rect 274422 667258 281186 667494
rect 281422 667258 288186 667494
rect 288422 667258 295186 667494
rect 295422 667258 302186 667494
rect 302422 667258 309186 667494
rect 309422 667258 316186 667494
rect 316422 667258 323186 667494
rect 323422 667258 330186 667494
rect 330422 667258 337186 667494
rect 337422 667258 344186 667494
rect 344422 667258 351186 667494
rect 351422 667258 358186 667494
rect 358422 667258 365186 667494
rect 365422 667258 372186 667494
rect 372422 667258 379186 667494
rect 379422 667258 386186 667494
rect 386422 667258 393186 667494
rect 393422 667258 400186 667494
rect 400422 667258 407186 667494
rect 407422 667258 414186 667494
rect 414422 667258 421186 667494
rect 421422 667258 428186 667494
rect 428422 667258 435186 667494
rect 435422 667258 442186 667494
rect 442422 667258 449186 667494
rect 449422 667258 456186 667494
rect 456422 667258 463186 667494
rect 463422 667258 470186 667494
rect 470422 667258 477186 667494
rect 477422 667258 484186 667494
rect 484422 667258 491186 667494
rect 491422 667258 498186 667494
rect 498422 667258 505186 667494
rect 505422 667258 512186 667494
rect 512422 667258 519186 667494
rect 519422 667258 526186 667494
rect 526422 667258 533186 667494
rect 533422 667258 540186 667494
rect 540422 667258 547186 667494
rect 547422 667258 554186 667494
rect 554422 667258 561186 667494
rect 561422 667258 568186 667494
rect 568422 667258 575186 667494
rect 575422 667258 582186 667494
rect 582422 667258 585818 667494
rect 586054 667258 586138 667494
rect 586374 667258 586458 667494
rect 586694 667258 586778 667494
rect 587014 667258 588874 667494
rect -4950 667216 588874 667258
rect -4950 661561 588874 661603
rect -4950 661325 -4842 661561
rect -4606 661325 -4522 661561
rect -4286 661325 -4202 661561
rect -3966 661325 -3882 661561
rect -3646 661325 2918 661561
rect 3154 661325 9918 661561
rect 10154 661325 16918 661561
rect 17154 661325 23918 661561
rect 24154 661325 30918 661561
rect 31154 661325 37918 661561
rect 38154 661325 44918 661561
rect 45154 661325 51918 661561
rect 52154 661325 58918 661561
rect 59154 661325 65918 661561
rect 66154 661325 72918 661561
rect 73154 661325 79918 661561
rect 80154 661325 86918 661561
rect 87154 661325 93918 661561
rect 94154 661325 100918 661561
rect 101154 661325 107918 661561
rect 108154 661325 114918 661561
rect 115154 661325 121918 661561
rect 122154 661325 128918 661561
rect 129154 661325 135918 661561
rect 136154 661325 142918 661561
rect 143154 661325 149918 661561
rect 150154 661325 156918 661561
rect 157154 661325 163918 661561
rect 164154 661325 170918 661561
rect 171154 661325 177918 661561
rect 178154 661325 184918 661561
rect 185154 661325 191918 661561
rect 192154 661325 198918 661561
rect 199154 661325 205918 661561
rect 206154 661325 212918 661561
rect 213154 661325 219918 661561
rect 220154 661325 226918 661561
rect 227154 661325 233918 661561
rect 234154 661325 240918 661561
rect 241154 661325 247918 661561
rect 248154 661325 254918 661561
rect 255154 661325 261918 661561
rect 262154 661325 268918 661561
rect 269154 661325 275918 661561
rect 276154 661325 282918 661561
rect 283154 661325 289918 661561
rect 290154 661325 296918 661561
rect 297154 661325 303918 661561
rect 304154 661325 310918 661561
rect 311154 661325 317918 661561
rect 318154 661325 324918 661561
rect 325154 661325 331918 661561
rect 332154 661325 338918 661561
rect 339154 661325 345918 661561
rect 346154 661325 352918 661561
rect 353154 661325 359918 661561
rect 360154 661325 366918 661561
rect 367154 661325 373918 661561
rect 374154 661325 380918 661561
rect 381154 661325 387918 661561
rect 388154 661325 394918 661561
rect 395154 661325 401918 661561
rect 402154 661325 408918 661561
rect 409154 661325 415918 661561
rect 416154 661325 422918 661561
rect 423154 661325 429918 661561
rect 430154 661325 436918 661561
rect 437154 661325 443918 661561
rect 444154 661325 450918 661561
rect 451154 661325 457918 661561
rect 458154 661325 464918 661561
rect 465154 661325 471918 661561
rect 472154 661325 478918 661561
rect 479154 661325 485918 661561
rect 486154 661325 492918 661561
rect 493154 661325 499918 661561
rect 500154 661325 506918 661561
rect 507154 661325 513918 661561
rect 514154 661325 520918 661561
rect 521154 661325 527918 661561
rect 528154 661325 534918 661561
rect 535154 661325 541918 661561
rect 542154 661325 548918 661561
rect 549154 661325 555918 661561
rect 556154 661325 562918 661561
rect 563154 661325 569918 661561
rect 570154 661325 576918 661561
rect 577154 661325 587570 661561
rect 587806 661325 587890 661561
rect 588126 661325 588210 661561
rect 588446 661325 588530 661561
rect 588766 661325 588874 661561
rect -4950 661283 588874 661325
rect -4950 660494 588874 660536
rect -4950 660258 -3090 660494
rect -2854 660258 -2770 660494
rect -2534 660258 -2450 660494
rect -2214 660258 -2130 660494
rect -1894 660258 1186 660494
rect 1422 660258 8186 660494
rect 8422 660258 15186 660494
rect 15422 660258 22186 660494
rect 22422 660258 29186 660494
rect 29422 660258 36186 660494
rect 36422 660258 43186 660494
rect 43422 660258 50186 660494
rect 50422 660258 57186 660494
rect 57422 660258 64186 660494
rect 64422 660258 71186 660494
rect 71422 660258 78186 660494
rect 78422 660258 85186 660494
rect 85422 660258 92186 660494
rect 92422 660258 99186 660494
rect 99422 660258 106186 660494
rect 106422 660258 113186 660494
rect 113422 660258 120186 660494
rect 120422 660258 127186 660494
rect 127422 660258 134186 660494
rect 134422 660258 141186 660494
rect 141422 660258 148186 660494
rect 148422 660258 155186 660494
rect 155422 660258 162186 660494
rect 162422 660258 169186 660494
rect 169422 660258 176186 660494
rect 176422 660258 183186 660494
rect 183422 660258 190186 660494
rect 190422 660258 197186 660494
rect 197422 660258 204186 660494
rect 204422 660258 211186 660494
rect 211422 660258 218186 660494
rect 218422 660258 225186 660494
rect 225422 660258 232186 660494
rect 232422 660258 239186 660494
rect 239422 660258 246186 660494
rect 246422 660258 253186 660494
rect 253422 660258 260186 660494
rect 260422 660258 267186 660494
rect 267422 660258 274186 660494
rect 274422 660258 281186 660494
rect 281422 660258 288186 660494
rect 288422 660258 295186 660494
rect 295422 660258 302186 660494
rect 302422 660258 309186 660494
rect 309422 660258 316186 660494
rect 316422 660258 323186 660494
rect 323422 660258 330186 660494
rect 330422 660258 337186 660494
rect 337422 660258 344186 660494
rect 344422 660258 351186 660494
rect 351422 660258 358186 660494
rect 358422 660258 365186 660494
rect 365422 660258 372186 660494
rect 372422 660258 379186 660494
rect 379422 660258 386186 660494
rect 386422 660258 393186 660494
rect 393422 660258 400186 660494
rect 400422 660258 407186 660494
rect 407422 660258 414186 660494
rect 414422 660258 421186 660494
rect 421422 660258 428186 660494
rect 428422 660258 435186 660494
rect 435422 660258 442186 660494
rect 442422 660258 449186 660494
rect 449422 660258 456186 660494
rect 456422 660258 463186 660494
rect 463422 660258 470186 660494
rect 470422 660258 477186 660494
rect 477422 660258 484186 660494
rect 484422 660258 491186 660494
rect 491422 660258 498186 660494
rect 498422 660258 505186 660494
rect 505422 660258 512186 660494
rect 512422 660258 519186 660494
rect 519422 660258 526186 660494
rect 526422 660258 533186 660494
rect 533422 660258 540186 660494
rect 540422 660258 547186 660494
rect 547422 660258 554186 660494
rect 554422 660258 561186 660494
rect 561422 660258 568186 660494
rect 568422 660258 575186 660494
rect 575422 660258 582186 660494
rect 582422 660258 585818 660494
rect 586054 660258 586138 660494
rect 586374 660258 586458 660494
rect 586694 660258 586778 660494
rect 587014 660258 588874 660494
rect -4950 660216 588874 660258
rect -4950 654561 588874 654603
rect -4950 654325 -4842 654561
rect -4606 654325 -4522 654561
rect -4286 654325 -4202 654561
rect -3966 654325 -3882 654561
rect -3646 654325 2918 654561
rect 3154 654325 9918 654561
rect 10154 654325 16918 654561
rect 17154 654325 23918 654561
rect 24154 654325 30918 654561
rect 31154 654325 37918 654561
rect 38154 654325 44918 654561
rect 45154 654325 51918 654561
rect 52154 654325 58918 654561
rect 59154 654325 65918 654561
rect 66154 654325 72918 654561
rect 73154 654325 79918 654561
rect 80154 654325 86918 654561
rect 87154 654325 93918 654561
rect 94154 654325 100918 654561
rect 101154 654325 107918 654561
rect 108154 654325 114918 654561
rect 115154 654325 121918 654561
rect 122154 654325 128918 654561
rect 129154 654325 135918 654561
rect 136154 654325 142918 654561
rect 143154 654325 149918 654561
rect 150154 654325 156918 654561
rect 157154 654325 163918 654561
rect 164154 654325 170918 654561
rect 171154 654325 177918 654561
rect 178154 654325 184918 654561
rect 185154 654325 191918 654561
rect 192154 654325 198918 654561
rect 199154 654325 205918 654561
rect 206154 654325 212918 654561
rect 213154 654325 219918 654561
rect 220154 654325 226918 654561
rect 227154 654325 233918 654561
rect 234154 654325 240918 654561
rect 241154 654325 247918 654561
rect 248154 654325 254918 654561
rect 255154 654325 261918 654561
rect 262154 654325 268918 654561
rect 269154 654325 275918 654561
rect 276154 654325 282918 654561
rect 283154 654325 289918 654561
rect 290154 654325 296918 654561
rect 297154 654325 303918 654561
rect 304154 654325 310918 654561
rect 311154 654325 317918 654561
rect 318154 654325 324918 654561
rect 325154 654325 331918 654561
rect 332154 654325 338918 654561
rect 339154 654325 345918 654561
rect 346154 654325 352918 654561
rect 353154 654325 359918 654561
rect 360154 654325 366918 654561
rect 367154 654325 373918 654561
rect 374154 654325 380918 654561
rect 381154 654325 387918 654561
rect 388154 654325 394918 654561
rect 395154 654325 401918 654561
rect 402154 654325 408918 654561
rect 409154 654325 415918 654561
rect 416154 654325 422918 654561
rect 423154 654325 429918 654561
rect 430154 654325 436918 654561
rect 437154 654325 443918 654561
rect 444154 654325 450918 654561
rect 451154 654325 457918 654561
rect 458154 654325 464918 654561
rect 465154 654325 471918 654561
rect 472154 654325 478918 654561
rect 479154 654325 485918 654561
rect 486154 654325 492918 654561
rect 493154 654325 499918 654561
rect 500154 654325 506918 654561
rect 507154 654325 513918 654561
rect 514154 654325 520918 654561
rect 521154 654325 527918 654561
rect 528154 654325 534918 654561
rect 535154 654325 541918 654561
rect 542154 654325 548918 654561
rect 549154 654325 555918 654561
rect 556154 654325 562918 654561
rect 563154 654325 569918 654561
rect 570154 654325 576918 654561
rect 577154 654325 587570 654561
rect 587806 654325 587890 654561
rect 588126 654325 588210 654561
rect 588446 654325 588530 654561
rect 588766 654325 588874 654561
rect -4950 654283 588874 654325
rect -4950 653494 588874 653536
rect -4950 653258 -3090 653494
rect -2854 653258 -2770 653494
rect -2534 653258 -2450 653494
rect -2214 653258 -2130 653494
rect -1894 653258 1186 653494
rect 1422 653258 8186 653494
rect 8422 653258 15186 653494
rect 15422 653258 22186 653494
rect 22422 653258 29186 653494
rect 29422 653258 36186 653494
rect 36422 653258 43186 653494
rect 43422 653258 50186 653494
rect 50422 653258 57186 653494
rect 57422 653258 64186 653494
rect 64422 653258 71186 653494
rect 71422 653258 78186 653494
rect 78422 653258 85186 653494
rect 85422 653258 92186 653494
rect 92422 653258 99186 653494
rect 99422 653258 106186 653494
rect 106422 653258 113186 653494
rect 113422 653258 120186 653494
rect 120422 653258 127186 653494
rect 127422 653258 134186 653494
rect 134422 653258 141186 653494
rect 141422 653258 148186 653494
rect 148422 653258 155186 653494
rect 155422 653258 162186 653494
rect 162422 653258 169186 653494
rect 169422 653258 176186 653494
rect 176422 653258 183186 653494
rect 183422 653258 190186 653494
rect 190422 653258 197186 653494
rect 197422 653258 204186 653494
rect 204422 653258 211186 653494
rect 211422 653258 218186 653494
rect 218422 653258 225186 653494
rect 225422 653258 232186 653494
rect 232422 653258 239186 653494
rect 239422 653258 246186 653494
rect 246422 653258 253186 653494
rect 253422 653258 260186 653494
rect 260422 653258 267186 653494
rect 267422 653258 274186 653494
rect 274422 653258 281186 653494
rect 281422 653258 288186 653494
rect 288422 653258 295186 653494
rect 295422 653258 302186 653494
rect 302422 653258 309186 653494
rect 309422 653258 316186 653494
rect 316422 653258 323186 653494
rect 323422 653258 330186 653494
rect 330422 653258 337186 653494
rect 337422 653258 344186 653494
rect 344422 653258 351186 653494
rect 351422 653258 358186 653494
rect 358422 653258 365186 653494
rect 365422 653258 372186 653494
rect 372422 653258 379186 653494
rect 379422 653258 386186 653494
rect 386422 653258 393186 653494
rect 393422 653258 400186 653494
rect 400422 653258 407186 653494
rect 407422 653258 414186 653494
rect 414422 653258 421186 653494
rect 421422 653258 428186 653494
rect 428422 653258 435186 653494
rect 435422 653258 442186 653494
rect 442422 653258 449186 653494
rect 449422 653258 456186 653494
rect 456422 653258 463186 653494
rect 463422 653258 470186 653494
rect 470422 653258 477186 653494
rect 477422 653258 484186 653494
rect 484422 653258 491186 653494
rect 491422 653258 498186 653494
rect 498422 653258 505186 653494
rect 505422 653258 512186 653494
rect 512422 653258 519186 653494
rect 519422 653258 526186 653494
rect 526422 653258 533186 653494
rect 533422 653258 540186 653494
rect 540422 653258 547186 653494
rect 547422 653258 554186 653494
rect 554422 653258 561186 653494
rect 561422 653258 568186 653494
rect 568422 653258 575186 653494
rect 575422 653258 582186 653494
rect 582422 653258 585818 653494
rect 586054 653258 586138 653494
rect 586374 653258 586458 653494
rect 586694 653258 586778 653494
rect 587014 653258 588874 653494
rect -4950 653216 588874 653258
rect -4950 647561 588874 647603
rect -4950 647325 -4842 647561
rect -4606 647325 -4522 647561
rect -4286 647325 -4202 647561
rect -3966 647325 -3882 647561
rect -3646 647325 2918 647561
rect 3154 647325 9918 647561
rect 10154 647325 16918 647561
rect 17154 647325 23918 647561
rect 24154 647325 30918 647561
rect 31154 647325 37918 647561
rect 38154 647325 44918 647561
rect 45154 647325 51918 647561
rect 52154 647325 58918 647561
rect 59154 647325 65918 647561
rect 66154 647325 72918 647561
rect 73154 647325 79918 647561
rect 80154 647325 86918 647561
rect 87154 647325 93918 647561
rect 94154 647325 100918 647561
rect 101154 647325 107918 647561
rect 108154 647325 114918 647561
rect 115154 647325 121918 647561
rect 122154 647325 128918 647561
rect 129154 647325 135918 647561
rect 136154 647325 142918 647561
rect 143154 647325 149918 647561
rect 150154 647325 156918 647561
rect 157154 647325 163918 647561
rect 164154 647325 170918 647561
rect 171154 647325 177918 647561
rect 178154 647325 184918 647561
rect 185154 647325 191918 647561
rect 192154 647325 198918 647561
rect 199154 647325 205918 647561
rect 206154 647325 212918 647561
rect 213154 647325 219918 647561
rect 220154 647325 226918 647561
rect 227154 647325 233918 647561
rect 234154 647325 240918 647561
rect 241154 647325 247918 647561
rect 248154 647325 254918 647561
rect 255154 647325 261918 647561
rect 262154 647325 268918 647561
rect 269154 647325 275918 647561
rect 276154 647325 282918 647561
rect 283154 647325 289918 647561
rect 290154 647325 296918 647561
rect 297154 647325 303918 647561
rect 304154 647325 310918 647561
rect 311154 647325 317918 647561
rect 318154 647325 324918 647561
rect 325154 647325 331918 647561
rect 332154 647325 338918 647561
rect 339154 647325 345918 647561
rect 346154 647325 352918 647561
rect 353154 647325 359918 647561
rect 360154 647325 366918 647561
rect 367154 647325 373918 647561
rect 374154 647325 380918 647561
rect 381154 647325 387918 647561
rect 388154 647325 394918 647561
rect 395154 647325 401918 647561
rect 402154 647325 408918 647561
rect 409154 647325 415918 647561
rect 416154 647325 422918 647561
rect 423154 647325 429918 647561
rect 430154 647325 436918 647561
rect 437154 647325 443918 647561
rect 444154 647325 450918 647561
rect 451154 647325 457918 647561
rect 458154 647325 464918 647561
rect 465154 647325 471918 647561
rect 472154 647325 478918 647561
rect 479154 647325 485918 647561
rect 486154 647325 492918 647561
rect 493154 647325 499918 647561
rect 500154 647325 506918 647561
rect 507154 647325 513918 647561
rect 514154 647325 520918 647561
rect 521154 647325 527918 647561
rect 528154 647325 534918 647561
rect 535154 647325 541918 647561
rect 542154 647325 548918 647561
rect 549154 647325 555918 647561
rect 556154 647325 562918 647561
rect 563154 647325 569918 647561
rect 570154 647325 576918 647561
rect 577154 647325 587570 647561
rect 587806 647325 587890 647561
rect 588126 647325 588210 647561
rect 588446 647325 588530 647561
rect 588766 647325 588874 647561
rect -4950 647283 588874 647325
rect -4950 646494 588874 646536
rect -4950 646258 -3090 646494
rect -2854 646258 -2770 646494
rect -2534 646258 -2450 646494
rect -2214 646258 -2130 646494
rect -1894 646258 1186 646494
rect 1422 646258 8186 646494
rect 8422 646258 15186 646494
rect 15422 646258 22186 646494
rect 22422 646258 29186 646494
rect 29422 646258 36186 646494
rect 36422 646258 43186 646494
rect 43422 646258 50186 646494
rect 50422 646258 57186 646494
rect 57422 646258 64186 646494
rect 64422 646258 71186 646494
rect 71422 646258 78186 646494
rect 78422 646258 85186 646494
rect 85422 646258 92186 646494
rect 92422 646258 99186 646494
rect 99422 646258 106186 646494
rect 106422 646258 113186 646494
rect 113422 646258 120186 646494
rect 120422 646258 127186 646494
rect 127422 646258 134186 646494
rect 134422 646258 141186 646494
rect 141422 646258 148186 646494
rect 148422 646258 155186 646494
rect 155422 646258 162186 646494
rect 162422 646258 169186 646494
rect 169422 646258 176186 646494
rect 176422 646258 183186 646494
rect 183422 646258 190186 646494
rect 190422 646258 197186 646494
rect 197422 646258 204186 646494
rect 204422 646258 211186 646494
rect 211422 646258 218186 646494
rect 218422 646258 225186 646494
rect 225422 646258 232186 646494
rect 232422 646258 239186 646494
rect 239422 646258 246186 646494
rect 246422 646258 253186 646494
rect 253422 646258 260186 646494
rect 260422 646258 267186 646494
rect 267422 646258 274186 646494
rect 274422 646258 281186 646494
rect 281422 646258 288186 646494
rect 288422 646258 295186 646494
rect 295422 646258 302186 646494
rect 302422 646258 309186 646494
rect 309422 646258 316186 646494
rect 316422 646258 323186 646494
rect 323422 646258 330186 646494
rect 330422 646258 337186 646494
rect 337422 646258 344186 646494
rect 344422 646258 351186 646494
rect 351422 646258 358186 646494
rect 358422 646258 365186 646494
rect 365422 646258 372186 646494
rect 372422 646258 379186 646494
rect 379422 646258 386186 646494
rect 386422 646258 393186 646494
rect 393422 646258 400186 646494
rect 400422 646258 407186 646494
rect 407422 646258 414186 646494
rect 414422 646258 421186 646494
rect 421422 646258 428186 646494
rect 428422 646258 435186 646494
rect 435422 646258 442186 646494
rect 442422 646258 449186 646494
rect 449422 646258 456186 646494
rect 456422 646258 463186 646494
rect 463422 646258 470186 646494
rect 470422 646258 477186 646494
rect 477422 646258 484186 646494
rect 484422 646258 491186 646494
rect 491422 646258 498186 646494
rect 498422 646258 505186 646494
rect 505422 646258 512186 646494
rect 512422 646258 519186 646494
rect 519422 646258 526186 646494
rect 526422 646258 533186 646494
rect 533422 646258 540186 646494
rect 540422 646258 547186 646494
rect 547422 646258 554186 646494
rect 554422 646258 561186 646494
rect 561422 646258 568186 646494
rect 568422 646258 575186 646494
rect 575422 646258 582186 646494
rect 582422 646258 585818 646494
rect 586054 646258 586138 646494
rect 586374 646258 586458 646494
rect 586694 646258 586778 646494
rect 587014 646258 588874 646494
rect -4950 646216 588874 646258
rect -4950 640561 588874 640603
rect -4950 640325 -4842 640561
rect -4606 640325 -4522 640561
rect -4286 640325 -4202 640561
rect -3966 640325 -3882 640561
rect -3646 640325 2918 640561
rect 3154 640325 9918 640561
rect 10154 640325 16918 640561
rect 17154 640325 23918 640561
rect 24154 640325 30918 640561
rect 31154 640325 37918 640561
rect 38154 640325 44918 640561
rect 45154 640325 51918 640561
rect 52154 640325 58918 640561
rect 59154 640325 65918 640561
rect 66154 640325 72918 640561
rect 73154 640325 79918 640561
rect 80154 640325 86918 640561
rect 87154 640325 93918 640561
rect 94154 640325 100918 640561
rect 101154 640325 107918 640561
rect 108154 640325 114918 640561
rect 115154 640325 121918 640561
rect 122154 640325 128918 640561
rect 129154 640325 135918 640561
rect 136154 640325 142918 640561
rect 143154 640325 149918 640561
rect 150154 640325 156918 640561
rect 157154 640325 163918 640561
rect 164154 640325 170918 640561
rect 171154 640325 177918 640561
rect 178154 640325 184918 640561
rect 185154 640325 191918 640561
rect 192154 640325 198918 640561
rect 199154 640325 205918 640561
rect 206154 640325 212918 640561
rect 213154 640325 219918 640561
rect 220154 640325 226918 640561
rect 227154 640325 233918 640561
rect 234154 640325 240918 640561
rect 241154 640325 247918 640561
rect 248154 640325 254918 640561
rect 255154 640325 261918 640561
rect 262154 640325 268918 640561
rect 269154 640325 275918 640561
rect 276154 640325 282918 640561
rect 283154 640325 289918 640561
rect 290154 640325 296918 640561
rect 297154 640325 303918 640561
rect 304154 640325 310918 640561
rect 311154 640325 317918 640561
rect 318154 640325 324918 640561
rect 325154 640325 331918 640561
rect 332154 640325 338918 640561
rect 339154 640325 345918 640561
rect 346154 640325 352918 640561
rect 353154 640325 359918 640561
rect 360154 640325 366918 640561
rect 367154 640325 373918 640561
rect 374154 640325 380918 640561
rect 381154 640325 387918 640561
rect 388154 640325 394918 640561
rect 395154 640325 401918 640561
rect 402154 640325 408918 640561
rect 409154 640325 415918 640561
rect 416154 640325 422918 640561
rect 423154 640325 429918 640561
rect 430154 640325 436918 640561
rect 437154 640325 443918 640561
rect 444154 640325 450918 640561
rect 451154 640325 457918 640561
rect 458154 640325 464918 640561
rect 465154 640325 471918 640561
rect 472154 640325 478918 640561
rect 479154 640325 485918 640561
rect 486154 640325 492918 640561
rect 493154 640325 499918 640561
rect 500154 640325 506918 640561
rect 507154 640325 513918 640561
rect 514154 640325 520918 640561
rect 521154 640325 527918 640561
rect 528154 640325 534918 640561
rect 535154 640325 541918 640561
rect 542154 640325 548918 640561
rect 549154 640325 555918 640561
rect 556154 640325 562918 640561
rect 563154 640325 569918 640561
rect 570154 640325 576918 640561
rect 577154 640325 587570 640561
rect 587806 640325 587890 640561
rect 588126 640325 588210 640561
rect 588446 640325 588530 640561
rect 588766 640325 588874 640561
rect -4950 640283 588874 640325
rect -4950 639494 588874 639536
rect -4950 639258 -3090 639494
rect -2854 639258 -2770 639494
rect -2534 639258 -2450 639494
rect -2214 639258 -2130 639494
rect -1894 639258 1186 639494
rect 1422 639258 8186 639494
rect 8422 639258 15186 639494
rect 15422 639258 22186 639494
rect 22422 639258 29186 639494
rect 29422 639258 36186 639494
rect 36422 639258 43186 639494
rect 43422 639258 50186 639494
rect 50422 639258 57186 639494
rect 57422 639258 64186 639494
rect 64422 639258 71186 639494
rect 71422 639258 78186 639494
rect 78422 639258 85186 639494
rect 85422 639258 92186 639494
rect 92422 639258 99186 639494
rect 99422 639258 106186 639494
rect 106422 639258 113186 639494
rect 113422 639258 120186 639494
rect 120422 639258 127186 639494
rect 127422 639258 134186 639494
rect 134422 639258 141186 639494
rect 141422 639258 148186 639494
rect 148422 639258 155186 639494
rect 155422 639258 162186 639494
rect 162422 639258 169186 639494
rect 169422 639258 176186 639494
rect 176422 639258 183186 639494
rect 183422 639258 190186 639494
rect 190422 639258 197186 639494
rect 197422 639258 204186 639494
rect 204422 639258 211186 639494
rect 211422 639258 218186 639494
rect 218422 639258 225186 639494
rect 225422 639258 232186 639494
rect 232422 639258 239186 639494
rect 239422 639258 246186 639494
rect 246422 639258 253186 639494
rect 253422 639258 260186 639494
rect 260422 639258 267186 639494
rect 267422 639258 274186 639494
rect 274422 639258 281186 639494
rect 281422 639258 288186 639494
rect 288422 639258 295186 639494
rect 295422 639258 302186 639494
rect 302422 639258 309186 639494
rect 309422 639258 316186 639494
rect 316422 639258 323186 639494
rect 323422 639258 330186 639494
rect 330422 639258 337186 639494
rect 337422 639258 344186 639494
rect 344422 639258 351186 639494
rect 351422 639258 358186 639494
rect 358422 639258 365186 639494
rect 365422 639258 372186 639494
rect 372422 639258 379186 639494
rect 379422 639258 386186 639494
rect 386422 639258 393186 639494
rect 393422 639258 400186 639494
rect 400422 639258 407186 639494
rect 407422 639258 414186 639494
rect 414422 639258 421186 639494
rect 421422 639258 428186 639494
rect 428422 639258 435186 639494
rect 435422 639258 442186 639494
rect 442422 639258 449186 639494
rect 449422 639258 456186 639494
rect 456422 639258 463186 639494
rect 463422 639258 470186 639494
rect 470422 639258 477186 639494
rect 477422 639258 484186 639494
rect 484422 639258 491186 639494
rect 491422 639258 498186 639494
rect 498422 639258 505186 639494
rect 505422 639258 512186 639494
rect 512422 639258 519186 639494
rect 519422 639258 526186 639494
rect 526422 639258 533186 639494
rect 533422 639258 540186 639494
rect 540422 639258 547186 639494
rect 547422 639258 554186 639494
rect 554422 639258 561186 639494
rect 561422 639258 568186 639494
rect 568422 639258 575186 639494
rect 575422 639258 582186 639494
rect 582422 639258 585818 639494
rect 586054 639258 586138 639494
rect 586374 639258 586458 639494
rect 586694 639258 586778 639494
rect 587014 639258 588874 639494
rect -4950 639216 588874 639258
rect -4950 633561 588874 633603
rect -4950 633325 -4842 633561
rect -4606 633325 -4522 633561
rect -4286 633325 -4202 633561
rect -3966 633325 -3882 633561
rect -3646 633325 2918 633561
rect 3154 633325 9918 633561
rect 10154 633325 16918 633561
rect 17154 633325 23918 633561
rect 24154 633325 30918 633561
rect 31154 633325 37918 633561
rect 38154 633325 44918 633561
rect 45154 633325 51918 633561
rect 52154 633325 58918 633561
rect 59154 633325 65918 633561
rect 66154 633325 72918 633561
rect 73154 633325 79918 633561
rect 80154 633325 86918 633561
rect 87154 633325 93918 633561
rect 94154 633325 100918 633561
rect 101154 633325 107918 633561
rect 108154 633325 114918 633561
rect 115154 633325 121918 633561
rect 122154 633325 128918 633561
rect 129154 633325 135918 633561
rect 136154 633325 142918 633561
rect 143154 633325 149918 633561
rect 150154 633325 156918 633561
rect 157154 633325 163918 633561
rect 164154 633325 170918 633561
rect 171154 633325 177918 633561
rect 178154 633325 184918 633561
rect 185154 633325 191918 633561
rect 192154 633325 198918 633561
rect 199154 633325 205918 633561
rect 206154 633325 212918 633561
rect 213154 633325 219918 633561
rect 220154 633325 226918 633561
rect 227154 633325 233918 633561
rect 234154 633325 240918 633561
rect 241154 633325 247918 633561
rect 248154 633325 254918 633561
rect 255154 633325 261918 633561
rect 262154 633325 268918 633561
rect 269154 633325 275918 633561
rect 276154 633325 282918 633561
rect 283154 633325 289918 633561
rect 290154 633325 296918 633561
rect 297154 633325 303918 633561
rect 304154 633325 310918 633561
rect 311154 633325 317918 633561
rect 318154 633325 324918 633561
rect 325154 633325 331918 633561
rect 332154 633325 338918 633561
rect 339154 633325 345918 633561
rect 346154 633325 352918 633561
rect 353154 633325 359918 633561
rect 360154 633325 366918 633561
rect 367154 633325 373918 633561
rect 374154 633325 380918 633561
rect 381154 633325 387918 633561
rect 388154 633325 394918 633561
rect 395154 633325 401918 633561
rect 402154 633325 408918 633561
rect 409154 633325 415918 633561
rect 416154 633325 422918 633561
rect 423154 633325 429918 633561
rect 430154 633325 436918 633561
rect 437154 633325 443918 633561
rect 444154 633325 450918 633561
rect 451154 633325 457918 633561
rect 458154 633325 464918 633561
rect 465154 633325 471918 633561
rect 472154 633325 478918 633561
rect 479154 633325 485918 633561
rect 486154 633325 492918 633561
rect 493154 633325 499918 633561
rect 500154 633325 506918 633561
rect 507154 633325 513918 633561
rect 514154 633325 520918 633561
rect 521154 633325 527918 633561
rect 528154 633325 534918 633561
rect 535154 633325 541918 633561
rect 542154 633325 548918 633561
rect 549154 633325 555918 633561
rect 556154 633325 562918 633561
rect 563154 633325 569918 633561
rect 570154 633325 576918 633561
rect 577154 633325 587570 633561
rect 587806 633325 587890 633561
rect 588126 633325 588210 633561
rect 588446 633325 588530 633561
rect 588766 633325 588874 633561
rect -4950 633283 588874 633325
rect -4950 632494 588874 632536
rect -4950 632258 -3090 632494
rect -2854 632258 -2770 632494
rect -2534 632258 -2450 632494
rect -2214 632258 -2130 632494
rect -1894 632258 1186 632494
rect 1422 632258 8186 632494
rect 8422 632258 15186 632494
rect 15422 632258 22186 632494
rect 22422 632258 29186 632494
rect 29422 632258 36186 632494
rect 36422 632258 43186 632494
rect 43422 632258 50186 632494
rect 50422 632258 57186 632494
rect 57422 632258 64186 632494
rect 64422 632258 71186 632494
rect 71422 632258 78186 632494
rect 78422 632258 85186 632494
rect 85422 632258 92186 632494
rect 92422 632258 99186 632494
rect 99422 632258 106186 632494
rect 106422 632258 113186 632494
rect 113422 632258 120186 632494
rect 120422 632258 127186 632494
rect 127422 632258 134186 632494
rect 134422 632258 141186 632494
rect 141422 632258 148186 632494
rect 148422 632258 155186 632494
rect 155422 632258 162186 632494
rect 162422 632258 169186 632494
rect 169422 632258 176186 632494
rect 176422 632258 183186 632494
rect 183422 632258 190186 632494
rect 190422 632258 197186 632494
rect 197422 632258 204186 632494
rect 204422 632258 211186 632494
rect 211422 632258 218186 632494
rect 218422 632258 225186 632494
rect 225422 632258 232186 632494
rect 232422 632258 239186 632494
rect 239422 632258 246186 632494
rect 246422 632258 253186 632494
rect 253422 632258 260186 632494
rect 260422 632258 267186 632494
rect 267422 632258 274186 632494
rect 274422 632258 281186 632494
rect 281422 632258 288186 632494
rect 288422 632258 295186 632494
rect 295422 632258 302186 632494
rect 302422 632258 309186 632494
rect 309422 632258 316186 632494
rect 316422 632258 323186 632494
rect 323422 632258 330186 632494
rect 330422 632258 337186 632494
rect 337422 632258 344186 632494
rect 344422 632258 351186 632494
rect 351422 632258 358186 632494
rect 358422 632258 365186 632494
rect 365422 632258 372186 632494
rect 372422 632258 379186 632494
rect 379422 632258 386186 632494
rect 386422 632258 393186 632494
rect 393422 632258 400186 632494
rect 400422 632258 407186 632494
rect 407422 632258 414186 632494
rect 414422 632258 421186 632494
rect 421422 632258 428186 632494
rect 428422 632258 435186 632494
rect 435422 632258 442186 632494
rect 442422 632258 449186 632494
rect 449422 632258 456186 632494
rect 456422 632258 463186 632494
rect 463422 632258 470186 632494
rect 470422 632258 477186 632494
rect 477422 632258 484186 632494
rect 484422 632258 491186 632494
rect 491422 632258 498186 632494
rect 498422 632258 505186 632494
rect 505422 632258 512186 632494
rect 512422 632258 519186 632494
rect 519422 632258 526186 632494
rect 526422 632258 533186 632494
rect 533422 632258 540186 632494
rect 540422 632258 547186 632494
rect 547422 632258 554186 632494
rect 554422 632258 561186 632494
rect 561422 632258 568186 632494
rect 568422 632258 575186 632494
rect 575422 632258 582186 632494
rect 582422 632258 585818 632494
rect 586054 632258 586138 632494
rect 586374 632258 586458 632494
rect 586694 632258 586778 632494
rect 587014 632258 588874 632494
rect -4950 632216 588874 632258
rect -4950 626561 588874 626603
rect -4950 626325 -4842 626561
rect -4606 626325 -4522 626561
rect -4286 626325 -4202 626561
rect -3966 626325 -3882 626561
rect -3646 626325 2918 626561
rect 3154 626325 9918 626561
rect 10154 626325 16918 626561
rect 17154 626325 23918 626561
rect 24154 626325 30918 626561
rect 31154 626325 37918 626561
rect 38154 626325 44918 626561
rect 45154 626325 51918 626561
rect 52154 626325 58918 626561
rect 59154 626325 65918 626561
rect 66154 626325 72918 626561
rect 73154 626325 79918 626561
rect 80154 626325 86918 626561
rect 87154 626325 93918 626561
rect 94154 626325 100918 626561
rect 101154 626325 107918 626561
rect 108154 626325 114918 626561
rect 115154 626325 121918 626561
rect 122154 626325 128918 626561
rect 129154 626325 135918 626561
rect 136154 626325 142918 626561
rect 143154 626325 149918 626561
rect 150154 626325 156918 626561
rect 157154 626325 163918 626561
rect 164154 626325 170918 626561
rect 171154 626325 177918 626561
rect 178154 626325 184918 626561
rect 185154 626325 191918 626561
rect 192154 626325 198918 626561
rect 199154 626325 205918 626561
rect 206154 626325 212918 626561
rect 213154 626325 219918 626561
rect 220154 626325 226918 626561
rect 227154 626325 233918 626561
rect 234154 626325 240918 626561
rect 241154 626325 247918 626561
rect 248154 626325 254918 626561
rect 255154 626325 261918 626561
rect 262154 626325 268918 626561
rect 269154 626325 275918 626561
rect 276154 626325 282918 626561
rect 283154 626325 289918 626561
rect 290154 626325 296918 626561
rect 297154 626325 303918 626561
rect 304154 626325 310918 626561
rect 311154 626325 317918 626561
rect 318154 626325 324918 626561
rect 325154 626325 331918 626561
rect 332154 626325 338918 626561
rect 339154 626325 345918 626561
rect 346154 626325 352918 626561
rect 353154 626325 359918 626561
rect 360154 626325 366918 626561
rect 367154 626325 373918 626561
rect 374154 626325 380918 626561
rect 381154 626325 387918 626561
rect 388154 626325 394918 626561
rect 395154 626325 401918 626561
rect 402154 626325 408918 626561
rect 409154 626325 415918 626561
rect 416154 626325 422918 626561
rect 423154 626325 429918 626561
rect 430154 626325 436918 626561
rect 437154 626325 443918 626561
rect 444154 626325 450918 626561
rect 451154 626325 457918 626561
rect 458154 626325 464918 626561
rect 465154 626325 471918 626561
rect 472154 626325 478918 626561
rect 479154 626325 485918 626561
rect 486154 626325 492918 626561
rect 493154 626325 499918 626561
rect 500154 626325 506918 626561
rect 507154 626325 513918 626561
rect 514154 626325 520918 626561
rect 521154 626325 527918 626561
rect 528154 626325 534918 626561
rect 535154 626325 541918 626561
rect 542154 626325 548918 626561
rect 549154 626325 555918 626561
rect 556154 626325 562918 626561
rect 563154 626325 569918 626561
rect 570154 626325 576918 626561
rect 577154 626325 587570 626561
rect 587806 626325 587890 626561
rect 588126 626325 588210 626561
rect 588446 626325 588530 626561
rect 588766 626325 588874 626561
rect -4950 626283 588874 626325
rect -4950 625494 588874 625536
rect -4950 625258 -3090 625494
rect -2854 625258 -2770 625494
rect -2534 625258 -2450 625494
rect -2214 625258 -2130 625494
rect -1894 625258 1186 625494
rect 1422 625258 8186 625494
rect 8422 625258 15186 625494
rect 15422 625258 22186 625494
rect 22422 625258 29186 625494
rect 29422 625258 36186 625494
rect 36422 625258 43186 625494
rect 43422 625258 50186 625494
rect 50422 625258 57186 625494
rect 57422 625258 64186 625494
rect 64422 625258 71186 625494
rect 71422 625258 78186 625494
rect 78422 625258 85186 625494
rect 85422 625258 92186 625494
rect 92422 625258 99186 625494
rect 99422 625258 106186 625494
rect 106422 625258 113186 625494
rect 113422 625258 120186 625494
rect 120422 625258 127186 625494
rect 127422 625258 134186 625494
rect 134422 625258 141186 625494
rect 141422 625258 148186 625494
rect 148422 625258 155186 625494
rect 155422 625258 162186 625494
rect 162422 625258 169186 625494
rect 169422 625258 176186 625494
rect 176422 625258 183186 625494
rect 183422 625258 190186 625494
rect 190422 625258 197186 625494
rect 197422 625258 204186 625494
rect 204422 625258 211186 625494
rect 211422 625258 218186 625494
rect 218422 625258 225186 625494
rect 225422 625258 232186 625494
rect 232422 625258 239186 625494
rect 239422 625258 246186 625494
rect 246422 625258 253186 625494
rect 253422 625258 260186 625494
rect 260422 625258 267186 625494
rect 267422 625258 274186 625494
rect 274422 625258 281186 625494
rect 281422 625258 288186 625494
rect 288422 625258 295186 625494
rect 295422 625258 302186 625494
rect 302422 625258 309186 625494
rect 309422 625258 316186 625494
rect 316422 625258 323186 625494
rect 323422 625258 330186 625494
rect 330422 625258 337186 625494
rect 337422 625258 344186 625494
rect 344422 625258 351186 625494
rect 351422 625258 358186 625494
rect 358422 625258 365186 625494
rect 365422 625258 372186 625494
rect 372422 625258 379186 625494
rect 379422 625258 386186 625494
rect 386422 625258 393186 625494
rect 393422 625258 400186 625494
rect 400422 625258 407186 625494
rect 407422 625258 414186 625494
rect 414422 625258 421186 625494
rect 421422 625258 428186 625494
rect 428422 625258 435186 625494
rect 435422 625258 442186 625494
rect 442422 625258 449186 625494
rect 449422 625258 456186 625494
rect 456422 625258 463186 625494
rect 463422 625258 470186 625494
rect 470422 625258 477186 625494
rect 477422 625258 484186 625494
rect 484422 625258 491186 625494
rect 491422 625258 498186 625494
rect 498422 625258 505186 625494
rect 505422 625258 512186 625494
rect 512422 625258 519186 625494
rect 519422 625258 526186 625494
rect 526422 625258 533186 625494
rect 533422 625258 540186 625494
rect 540422 625258 547186 625494
rect 547422 625258 554186 625494
rect 554422 625258 561186 625494
rect 561422 625258 568186 625494
rect 568422 625258 575186 625494
rect 575422 625258 582186 625494
rect 582422 625258 585818 625494
rect 586054 625258 586138 625494
rect 586374 625258 586458 625494
rect 586694 625258 586778 625494
rect 587014 625258 588874 625494
rect -4950 625216 588874 625258
rect -4950 619561 588874 619603
rect -4950 619325 -4842 619561
rect -4606 619325 -4522 619561
rect -4286 619325 -4202 619561
rect -3966 619325 -3882 619561
rect -3646 619325 2918 619561
rect 3154 619325 9918 619561
rect 10154 619325 16918 619561
rect 17154 619325 23918 619561
rect 24154 619325 30918 619561
rect 31154 619325 37918 619561
rect 38154 619325 44918 619561
rect 45154 619325 51918 619561
rect 52154 619325 58918 619561
rect 59154 619325 65918 619561
rect 66154 619325 72918 619561
rect 73154 619325 79918 619561
rect 80154 619325 86918 619561
rect 87154 619325 93918 619561
rect 94154 619325 100918 619561
rect 101154 619325 107918 619561
rect 108154 619325 114918 619561
rect 115154 619325 121918 619561
rect 122154 619325 128918 619561
rect 129154 619325 135918 619561
rect 136154 619325 142918 619561
rect 143154 619325 149918 619561
rect 150154 619325 156918 619561
rect 157154 619325 163918 619561
rect 164154 619325 170918 619561
rect 171154 619325 177918 619561
rect 178154 619325 184918 619561
rect 185154 619325 191918 619561
rect 192154 619325 198918 619561
rect 199154 619325 205918 619561
rect 206154 619325 212918 619561
rect 213154 619325 219918 619561
rect 220154 619325 226918 619561
rect 227154 619325 233918 619561
rect 234154 619325 240918 619561
rect 241154 619325 247918 619561
rect 248154 619325 254918 619561
rect 255154 619325 261918 619561
rect 262154 619325 268918 619561
rect 269154 619325 275918 619561
rect 276154 619325 282918 619561
rect 283154 619325 289918 619561
rect 290154 619325 296918 619561
rect 297154 619325 303918 619561
rect 304154 619325 310918 619561
rect 311154 619325 317918 619561
rect 318154 619325 324918 619561
rect 325154 619325 331918 619561
rect 332154 619325 338918 619561
rect 339154 619325 345918 619561
rect 346154 619325 352918 619561
rect 353154 619325 359918 619561
rect 360154 619325 366918 619561
rect 367154 619325 373918 619561
rect 374154 619325 380918 619561
rect 381154 619325 387918 619561
rect 388154 619325 394918 619561
rect 395154 619325 401918 619561
rect 402154 619325 408918 619561
rect 409154 619325 415918 619561
rect 416154 619325 422918 619561
rect 423154 619325 429918 619561
rect 430154 619325 436918 619561
rect 437154 619325 443918 619561
rect 444154 619325 450918 619561
rect 451154 619325 457918 619561
rect 458154 619325 464918 619561
rect 465154 619325 471918 619561
rect 472154 619325 478918 619561
rect 479154 619325 485918 619561
rect 486154 619325 492918 619561
rect 493154 619325 499918 619561
rect 500154 619325 506918 619561
rect 507154 619325 513918 619561
rect 514154 619325 520918 619561
rect 521154 619325 527918 619561
rect 528154 619325 534918 619561
rect 535154 619325 541918 619561
rect 542154 619325 548918 619561
rect 549154 619325 555918 619561
rect 556154 619325 562918 619561
rect 563154 619325 569918 619561
rect 570154 619325 576918 619561
rect 577154 619325 587570 619561
rect 587806 619325 587890 619561
rect 588126 619325 588210 619561
rect 588446 619325 588530 619561
rect 588766 619325 588874 619561
rect -4950 619283 588874 619325
rect -4950 618494 588874 618536
rect -4950 618258 -3090 618494
rect -2854 618258 -2770 618494
rect -2534 618258 -2450 618494
rect -2214 618258 -2130 618494
rect -1894 618258 1186 618494
rect 1422 618258 8186 618494
rect 8422 618258 15186 618494
rect 15422 618258 22186 618494
rect 22422 618258 29186 618494
rect 29422 618258 36186 618494
rect 36422 618258 43186 618494
rect 43422 618258 50186 618494
rect 50422 618258 57186 618494
rect 57422 618258 64186 618494
rect 64422 618258 71186 618494
rect 71422 618258 78186 618494
rect 78422 618258 85186 618494
rect 85422 618258 92186 618494
rect 92422 618258 99186 618494
rect 99422 618258 106186 618494
rect 106422 618258 113186 618494
rect 113422 618258 120186 618494
rect 120422 618258 127186 618494
rect 127422 618258 134186 618494
rect 134422 618258 141186 618494
rect 141422 618258 148186 618494
rect 148422 618258 155186 618494
rect 155422 618258 162186 618494
rect 162422 618258 169186 618494
rect 169422 618258 176186 618494
rect 176422 618258 183186 618494
rect 183422 618258 190186 618494
rect 190422 618258 197186 618494
rect 197422 618258 204186 618494
rect 204422 618258 211186 618494
rect 211422 618258 218186 618494
rect 218422 618258 225186 618494
rect 225422 618258 232186 618494
rect 232422 618258 239186 618494
rect 239422 618258 246186 618494
rect 246422 618258 253186 618494
rect 253422 618258 260186 618494
rect 260422 618258 267186 618494
rect 267422 618258 274186 618494
rect 274422 618258 281186 618494
rect 281422 618258 288186 618494
rect 288422 618258 295186 618494
rect 295422 618258 302186 618494
rect 302422 618258 309186 618494
rect 309422 618258 316186 618494
rect 316422 618258 323186 618494
rect 323422 618258 330186 618494
rect 330422 618258 337186 618494
rect 337422 618258 344186 618494
rect 344422 618258 351186 618494
rect 351422 618258 358186 618494
rect 358422 618258 365186 618494
rect 365422 618258 372186 618494
rect 372422 618258 379186 618494
rect 379422 618258 386186 618494
rect 386422 618258 393186 618494
rect 393422 618258 400186 618494
rect 400422 618258 407186 618494
rect 407422 618258 414186 618494
rect 414422 618258 421186 618494
rect 421422 618258 428186 618494
rect 428422 618258 435186 618494
rect 435422 618258 442186 618494
rect 442422 618258 449186 618494
rect 449422 618258 456186 618494
rect 456422 618258 463186 618494
rect 463422 618258 470186 618494
rect 470422 618258 477186 618494
rect 477422 618258 484186 618494
rect 484422 618258 491186 618494
rect 491422 618258 498186 618494
rect 498422 618258 505186 618494
rect 505422 618258 512186 618494
rect 512422 618258 519186 618494
rect 519422 618258 526186 618494
rect 526422 618258 533186 618494
rect 533422 618258 540186 618494
rect 540422 618258 547186 618494
rect 547422 618258 554186 618494
rect 554422 618258 561186 618494
rect 561422 618258 568186 618494
rect 568422 618258 575186 618494
rect 575422 618258 582186 618494
rect 582422 618258 585818 618494
rect 586054 618258 586138 618494
rect 586374 618258 586458 618494
rect 586694 618258 586778 618494
rect 587014 618258 588874 618494
rect -4950 618216 588874 618258
rect -4950 612561 588874 612603
rect -4950 612325 -4842 612561
rect -4606 612325 -4522 612561
rect -4286 612325 -4202 612561
rect -3966 612325 -3882 612561
rect -3646 612325 2918 612561
rect 3154 612325 9918 612561
rect 10154 612325 16918 612561
rect 17154 612325 23918 612561
rect 24154 612325 30918 612561
rect 31154 612325 37918 612561
rect 38154 612325 44918 612561
rect 45154 612325 51918 612561
rect 52154 612325 58918 612561
rect 59154 612325 65918 612561
rect 66154 612325 72918 612561
rect 73154 612325 79918 612561
rect 80154 612325 86918 612561
rect 87154 612325 93918 612561
rect 94154 612325 100918 612561
rect 101154 612325 107918 612561
rect 108154 612325 114918 612561
rect 115154 612325 121918 612561
rect 122154 612325 128918 612561
rect 129154 612325 135918 612561
rect 136154 612325 142918 612561
rect 143154 612325 149918 612561
rect 150154 612325 156918 612561
rect 157154 612325 163918 612561
rect 164154 612325 170918 612561
rect 171154 612325 177918 612561
rect 178154 612325 184918 612561
rect 185154 612325 191918 612561
rect 192154 612325 198918 612561
rect 199154 612325 205918 612561
rect 206154 612325 212918 612561
rect 213154 612325 219918 612561
rect 220154 612325 226918 612561
rect 227154 612325 233918 612561
rect 234154 612325 240918 612561
rect 241154 612325 247918 612561
rect 248154 612325 254918 612561
rect 255154 612325 261918 612561
rect 262154 612325 268918 612561
rect 269154 612325 275918 612561
rect 276154 612325 282918 612561
rect 283154 612325 289918 612561
rect 290154 612325 296918 612561
rect 297154 612325 303918 612561
rect 304154 612325 310918 612561
rect 311154 612325 317918 612561
rect 318154 612325 324918 612561
rect 325154 612325 331918 612561
rect 332154 612325 338918 612561
rect 339154 612325 345918 612561
rect 346154 612325 352918 612561
rect 353154 612325 359918 612561
rect 360154 612325 366918 612561
rect 367154 612325 373918 612561
rect 374154 612325 380918 612561
rect 381154 612325 387918 612561
rect 388154 612325 394918 612561
rect 395154 612325 401918 612561
rect 402154 612325 408918 612561
rect 409154 612325 415918 612561
rect 416154 612325 422918 612561
rect 423154 612325 429918 612561
rect 430154 612325 436918 612561
rect 437154 612325 443918 612561
rect 444154 612325 450918 612561
rect 451154 612325 457918 612561
rect 458154 612325 464918 612561
rect 465154 612325 471918 612561
rect 472154 612325 478918 612561
rect 479154 612325 485918 612561
rect 486154 612325 492918 612561
rect 493154 612325 499918 612561
rect 500154 612325 506918 612561
rect 507154 612325 513918 612561
rect 514154 612325 520918 612561
rect 521154 612325 527918 612561
rect 528154 612325 534918 612561
rect 535154 612325 541918 612561
rect 542154 612325 548918 612561
rect 549154 612325 555918 612561
rect 556154 612325 562918 612561
rect 563154 612325 569918 612561
rect 570154 612325 576918 612561
rect 577154 612325 587570 612561
rect 587806 612325 587890 612561
rect 588126 612325 588210 612561
rect 588446 612325 588530 612561
rect 588766 612325 588874 612561
rect -4950 612283 588874 612325
rect -4950 611494 588874 611536
rect -4950 611258 -3090 611494
rect -2854 611258 -2770 611494
rect -2534 611258 -2450 611494
rect -2214 611258 -2130 611494
rect -1894 611258 1186 611494
rect 1422 611258 8186 611494
rect 8422 611258 15186 611494
rect 15422 611258 22186 611494
rect 22422 611258 29186 611494
rect 29422 611258 36186 611494
rect 36422 611258 43186 611494
rect 43422 611258 50186 611494
rect 50422 611258 57186 611494
rect 57422 611258 64186 611494
rect 64422 611258 71186 611494
rect 71422 611258 78186 611494
rect 78422 611258 85186 611494
rect 85422 611258 92186 611494
rect 92422 611258 99186 611494
rect 99422 611258 106186 611494
rect 106422 611258 113186 611494
rect 113422 611258 120186 611494
rect 120422 611258 127186 611494
rect 127422 611258 134186 611494
rect 134422 611258 141186 611494
rect 141422 611258 148186 611494
rect 148422 611258 155186 611494
rect 155422 611258 162186 611494
rect 162422 611258 169186 611494
rect 169422 611258 176186 611494
rect 176422 611258 183186 611494
rect 183422 611258 190186 611494
rect 190422 611258 197186 611494
rect 197422 611258 204186 611494
rect 204422 611258 211186 611494
rect 211422 611258 218186 611494
rect 218422 611258 225186 611494
rect 225422 611258 232186 611494
rect 232422 611258 239186 611494
rect 239422 611258 246186 611494
rect 246422 611258 253186 611494
rect 253422 611258 260186 611494
rect 260422 611258 267186 611494
rect 267422 611258 274186 611494
rect 274422 611258 281186 611494
rect 281422 611258 288186 611494
rect 288422 611258 295186 611494
rect 295422 611258 302186 611494
rect 302422 611258 309186 611494
rect 309422 611258 316186 611494
rect 316422 611258 323186 611494
rect 323422 611258 330186 611494
rect 330422 611258 337186 611494
rect 337422 611258 344186 611494
rect 344422 611258 351186 611494
rect 351422 611258 358186 611494
rect 358422 611258 365186 611494
rect 365422 611258 372186 611494
rect 372422 611258 379186 611494
rect 379422 611258 386186 611494
rect 386422 611258 393186 611494
rect 393422 611258 400186 611494
rect 400422 611258 407186 611494
rect 407422 611258 414186 611494
rect 414422 611258 421186 611494
rect 421422 611258 428186 611494
rect 428422 611258 435186 611494
rect 435422 611258 442186 611494
rect 442422 611258 449186 611494
rect 449422 611258 456186 611494
rect 456422 611258 463186 611494
rect 463422 611258 470186 611494
rect 470422 611258 477186 611494
rect 477422 611258 484186 611494
rect 484422 611258 491186 611494
rect 491422 611258 498186 611494
rect 498422 611258 505186 611494
rect 505422 611258 512186 611494
rect 512422 611258 519186 611494
rect 519422 611258 526186 611494
rect 526422 611258 533186 611494
rect 533422 611258 540186 611494
rect 540422 611258 547186 611494
rect 547422 611258 554186 611494
rect 554422 611258 561186 611494
rect 561422 611258 568186 611494
rect 568422 611258 575186 611494
rect 575422 611258 582186 611494
rect 582422 611258 585818 611494
rect 586054 611258 586138 611494
rect 586374 611258 586458 611494
rect 586694 611258 586778 611494
rect 587014 611258 588874 611494
rect -4950 611216 588874 611258
rect -4950 605561 588874 605603
rect -4950 605325 -4842 605561
rect -4606 605325 -4522 605561
rect -4286 605325 -4202 605561
rect -3966 605325 -3882 605561
rect -3646 605325 2918 605561
rect 3154 605325 9918 605561
rect 10154 605325 16918 605561
rect 17154 605325 23918 605561
rect 24154 605325 30918 605561
rect 31154 605325 37918 605561
rect 38154 605325 44918 605561
rect 45154 605325 51918 605561
rect 52154 605325 58918 605561
rect 59154 605325 65918 605561
rect 66154 605325 72918 605561
rect 73154 605325 79918 605561
rect 80154 605325 86918 605561
rect 87154 605325 93918 605561
rect 94154 605325 100918 605561
rect 101154 605325 107918 605561
rect 108154 605325 114918 605561
rect 115154 605325 121918 605561
rect 122154 605325 128918 605561
rect 129154 605325 135918 605561
rect 136154 605325 142918 605561
rect 143154 605325 149918 605561
rect 150154 605325 156918 605561
rect 157154 605325 163918 605561
rect 164154 605325 170918 605561
rect 171154 605325 177918 605561
rect 178154 605325 184918 605561
rect 185154 605325 191918 605561
rect 192154 605325 198918 605561
rect 199154 605325 205918 605561
rect 206154 605325 212918 605561
rect 213154 605325 219918 605561
rect 220154 605325 226918 605561
rect 227154 605325 233918 605561
rect 234154 605325 240918 605561
rect 241154 605325 247918 605561
rect 248154 605325 254918 605561
rect 255154 605325 261918 605561
rect 262154 605325 268918 605561
rect 269154 605325 275918 605561
rect 276154 605325 282918 605561
rect 283154 605325 289918 605561
rect 290154 605325 296918 605561
rect 297154 605325 303918 605561
rect 304154 605325 310918 605561
rect 311154 605325 317918 605561
rect 318154 605325 324918 605561
rect 325154 605325 331918 605561
rect 332154 605325 338918 605561
rect 339154 605325 345918 605561
rect 346154 605325 352918 605561
rect 353154 605325 359918 605561
rect 360154 605325 366918 605561
rect 367154 605325 373918 605561
rect 374154 605325 380918 605561
rect 381154 605325 387918 605561
rect 388154 605325 394918 605561
rect 395154 605325 401918 605561
rect 402154 605325 408918 605561
rect 409154 605325 415918 605561
rect 416154 605325 422918 605561
rect 423154 605325 429918 605561
rect 430154 605325 436918 605561
rect 437154 605325 443918 605561
rect 444154 605325 450918 605561
rect 451154 605325 457918 605561
rect 458154 605325 464918 605561
rect 465154 605325 471918 605561
rect 472154 605325 478918 605561
rect 479154 605325 485918 605561
rect 486154 605325 492918 605561
rect 493154 605325 499918 605561
rect 500154 605325 506918 605561
rect 507154 605325 513918 605561
rect 514154 605325 520918 605561
rect 521154 605325 527918 605561
rect 528154 605325 534918 605561
rect 535154 605325 541918 605561
rect 542154 605325 548918 605561
rect 549154 605325 555918 605561
rect 556154 605325 562918 605561
rect 563154 605325 569918 605561
rect 570154 605325 576918 605561
rect 577154 605325 587570 605561
rect 587806 605325 587890 605561
rect 588126 605325 588210 605561
rect 588446 605325 588530 605561
rect 588766 605325 588874 605561
rect -4950 605283 588874 605325
rect -4950 604494 588874 604536
rect -4950 604258 -3090 604494
rect -2854 604258 -2770 604494
rect -2534 604258 -2450 604494
rect -2214 604258 -2130 604494
rect -1894 604258 1186 604494
rect 1422 604258 8186 604494
rect 8422 604258 15186 604494
rect 15422 604258 22186 604494
rect 22422 604258 29186 604494
rect 29422 604258 36186 604494
rect 36422 604258 43186 604494
rect 43422 604258 50186 604494
rect 50422 604258 57186 604494
rect 57422 604258 64186 604494
rect 64422 604258 71186 604494
rect 71422 604258 78186 604494
rect 78422 604258 85186 604494
rect 85422 604258 92186 604494
rect 92422 604258 99186 604494
rect 99422 604258 106186 604494
rect 106422 604258 113186 604494
rect 113422 604258 120186 604494
rect 120422 604258 127186 604494
rect 127422 604258 134186 604494
rect 134422 604258 141186 604494
rect 141422 604258 148186 604494
rect 148422 604258 155186 604494
rect 155422 604258 162186 604494
rect 162422 604258 169186 604494
rect 169422 604258 176186 604494
rect 176422 604258 183186 604494
rect 183422 604258 190186 604494
rect 190422 604258 197186 604494
rect 197422 604258 204186 604494
rect 204422 604258 211186 604494
rect 211422 604258 218186 604494
rect 218422 604258 225186 604494
rect 225422 604258 232186 604494
rect 232422 604258 239186 604494
rect 239422 604258 246186 604494
rect 246422 604258 253186 604494
rect 253422 604258 260186 604494
rect 260422 604258 267186 604494
rect 267422 604258 274186 604494
rect 274422 604258 281186 604494
rect 281422 604258 288186 604494
rect 288422 604258 295186 604494
rect 295422 604258 302186 604494
rect 302422 604258 309186 604494
rect 309422 604258 316186 604494
rect 316422 604258 323186 604494
rect 323422 604258 330186 604494
rect 330422 604258 337186 604494
rect 337422 604258 344186 604494
rect 344422 604258 351186 604494
rect 351422 604258 358186 604494
rect 358422 604258 365186 604494
rect 365422 604258 372186 604494
rect 372422 604258 379186 604494
rect 379422 604258 386186 604494
rect 386422 604258 393186 604494
rect 393422 604258 400186 604494
rect 400422 604258 407186 604494
rect 407422 604258 414186 604494
rect 414422 604258 421186 604494
rect 421422 604258 428186 604494
rect 428422 604258 435186 604494
rect 435422 604258 442186 604494
rect 442422 604258 449186 604494
rect 449422 604258 456186 604494
rect 456422 604258 463186 604494
rect 463422 604258 470186 604494
rect 470422 604258 477186 604494
rect 477422 604258 484186 604494
rect 484422 604258 491186 604494
rect 491422 604258 498186 604494
rect 498422 604258 505186 604494
rect 505422 604258 512186 604494
rect 512422 604258 519186 604494
rect 519422 604258 526186 604494
rect 526422 604258 533186 604494
rect 533422 604258 540186 604494
rect 540422 604258 547186 604494
rect 547422 604258 554186 604494
rect 554422 604258 561186 604494
rect 561422 604258 568186 604494
rect 568422 604258 575186 604494
rect 575422 604258 582186 604494
rect 582422 604258 585818 604494
rect 586054 604258 586138 604494
rect 586374 604258 586458 604494
rect 586694 604258 586778 604494
rect 587014 604258 588874 604494
rect -4950 604216 588874 604258
rect -4950 598561 588874 598603
rect -4950 598325 -4842 598561
rect -4606 598325 -4522 598561
rect -4286 598325 -4202 598561
rect -3966 598325 -3882 598561
rect -3646 598325 2918 598561
rect 3154 598325 9918 598561
rect 10154 598325 16918 598561
rect 17154 598325 23918 598561
rect 24154 598325 30918 598561
rect 31154 598325 37918 598561
rect 38154 598325 44918 598561
rect 45154 598325 51918 598561
rect 52154 598325 58918 598561
rect 59154 598325 65918 598561
rect 66154 598325 72918 598561
rect 73154 598325 79918 598561
rect 80154 598325 86918 598561
rect 87154 598325 93918 598561
rect 94154 598325 100918 598561
rect 101154 598325 107918 598561
rect 108154 598325 114918 598561
rect 115154 598325 121918 598561
rect 122154 598325 128918 598561
rect 129154 598325 135918 598561
rect 136154 598325 142918 598561
rect 143154 598325 149918 598561
rect 150154 598325 156918 598561
rect 157154 598325 163918 598561
rect 164154 598325 170918 598561
rect 171154 598325 177918 598561
rect 178154 598325 184918 598561
rect 185154 598325 191918 598561
rect 192154 598325 198918 598561
rect 199154 598325 205918 598561
rect 206154 598325 212918 598561
rect 213154 598325 219918 598561
rect 220154 598325 226918 598561
rect 227154 598325 233918 598561
rect 234154 598325 240918 598561
rect 241154 598325 247918 598561
rect 248154 598325 254918 598561
rect 255154 598325 261918 598561
rect 262154 598325 268918 598561
rect 269154 598325 275918 598561
rect 276154 598325 282918 598561
rect 283154 598325 289918 598561
rect 290154 598325 296918 598561
rect 297154 598325 303918 598561
rect 304154 598325 310918 598561
rect 311154 598325 317918 598561
rect 318154 598325 324918 598561
rect 325154 598325 331918 598561
rect 332154 598325 338918 598561
rect 339154 598325 345918 598561
rect 346154 598325 352918 598561
rect 353154 598325 359918 598561
rect 360154 598325 366918 598561
rect 367154 598325 373918 598561
rect 374154 598325 380918 598561
rect 381154 598325 387918 598561
rect 388154 598325 394918 598561
rect 395154 598325 401918 598561
rect 402154 598325 408918 598561
rect 409154 598325 415918 598561
rect 416154 598325 422918 598561
rect 423154 598325 429918 598561
rect 430154 598325 436918 598561
rect 437154 598325 443918 598561
rect 444154 598325 450918 598561
rect 451154 598325 457918 598561
rect 458154 598325 464918 598561
rect 465154 598325 471918 598561
rect 472154 598325 478918 598561
rect 479154 598325 485918 598561
rect 486154 598325 492918 598561
rect 493154 598325 499918 598561
rect 500154 598325 506918 598561
rect 507154 598325 513918 598561
rect 514154 598325 520918 598561
rect 521154 598325 527918 598561
rect 528154 598325 534918 598561
rect 535154 598325 541918 598561
rect 542154 598325 548918 598561
rect 549154 598325 555918 598561
rect 556154 598325 562918 598561
rect 563154 598325 569918 598561
rect 570154 598325 576918 598561
rect 577154 598325 587570 598561
rect 587806 598325 587890 598561
rect 588126 598325 588210 598561
rect 588446 598325 588530 598561
rect 588766 598325 588874 598561
rect -4950 598283 588874 598325
rect -4950 597494 588874 597536
rect -4950 597258 -3090 597494
rect -2854 597258 -2770 597494
rect -2534 597258 -2450 597494
rect -2214 597258 -2130 597494
rect -1894 597258 1186 597494
rect 1422 597258 8186 597494
rect 8422 597258 15186 597494
rect 15422 597258 22186 597494
rect 22422 597258 29186 597494
rect 29422 597258 36186 597494
rect 36422 597258 43186 597494
rect 43422 597258 50186 597494
rect 50422 597258 57186 597494
rect 57422 597258 64186 597494
rect 64422 597258 71186 597494
rect 71422 597258 78186 597494
rect 78422 597258 85186 597494
rect 85422 597258 92186 597494
rect 92422 597258 99186 597494
rect 99422 597258 106186 597494
rect 106422 597258 113186 597494
rect 113422 597258 120186 597494
rect 120422 597258 127186 597494
rect 127422 597258 134186 597494
rect 134422 597258 141186 597494
rect 141422 597258 148186 597494
rect 148422 597258 155186 597494
rect 155422 597258 162186 597494
rect 162422 597258 169186 597494
rect 169422 597258 176186 597494
rect 176422 597258 183186 597494
rect 183422 597258 190186 597494
rect 190422 597258 197186 597494
rect 197422 597258 204186 597494
rect 204422 597258 211186 597494
rect 211422 597258 218186 597494
rect 218422 597258 225186 597494
rect 225422 597258 232186 597494
rect 232422 597258 239186 597494
rect 239422 597258 246186 597494
rect 246422 597258 253186 597494
rect 253422 597258 260186 597494
rect 260422 597258 267186 597494
rect 267422 597258 274186 597494
rect 274422 597258 281186 597494
rect 281422 597258 288186 597494
rect 288422 597258 295186 597494
rect 295422 597258 302186 597494
rect 302422 597258 309186 597494
rect 309422 597258 316186 597494
rect 316422 597258 323186 597494
rect 323422 597258 330186 597494
rect 330422 597258 337186 597494
rect 337422 597258 344186 597494
rect 344422 597258 351186 597494
rect 351422 597258 358186 597494
rect 358422 597258 365186 597494
rect 365422 597258 372186 597494
rect 372422 597258 379186 597494
rect 379422 597258 386186 597494
rect 386422 597258 393186 597494
rect 393422 597258 400186 597494
rect 400422 597258 407186 597494
rect 407422 597258 414186 597494
rect 414422 597258 421186 597494
rect 421422 597258 428186 597494
rect 428422 597258 435186 597494
rect 435422 597258 442186 597494
rect 442422 597258 449186 597494
rect 449422 597258 456186 597494
rect 456422 597258 463186 597494
rect 463422 597258 470186 597494
rect 470422 597258 477186 597494
rect 477422 597258 484186 597494
rect 484422 597258 491186 597494
rect 491422 597258 498186 597494
rect 498422 597258 505186 597494
rect 505422 597258 512186 597494
rect 512422 597258 519186 597494
rect 519422 597258 526186 597494
rect 526422 597258 533186 597494
rect 533422 597258 540186 597494
rect 540422 597258 547186 597494
rect 547422 597258 554186 597494
rect 554422 597258 561186 597494
rect 561422 597258 568186 597494
rect 568422 597258 575186 597494
rect 575422 597258 582186 597494
rect 582422 597258 585818 597494
rect 586054 597258 586138 597494
rect 586374 597258 586458 597494
rect 586694 597258 586778 597494
rect 587014 597258 588874 597494
rect -4950 597216 588874 597258
rect -4950 591561 588874 591603
rect -4950 591325 -4842 591561
rect -4606 591325 -4522 591561
rect -4286 591325 -4202 591561
rect -3966 591325 -3882 591561
rect -3646 591325 2918 591561
rect 3154 591325 9918 591561
rect 10154 591325 16918 591561
rect 17154 591325 23918 591561
rect 24154 591325 30918 591561
rect 31154 591325 37918 591561
rect 38154 591325 44918 591561
rect 45154 591325 51918 591561
rect 52154 591325 58918 591561
rect 59154 591325 65918 591561
rect 66154 591325 72918 591561
rect 73154 591325 79918 591561
rect 80154 591325 86918 591561
rect 87154 591325 93918 591561
rect 94154 591325 100918 591561
rect 101154 591325 107918 591561
rect 108154 591325 114918 591561
rect 115154 591325 121918 591561
rect 122154 591325 128918 591561
rect 129154 591325 135918 591561
rect 136154 591325 142918 591561
rect 143154 591325 149918 591561
rect 150154 591325 156918 591561
rect 157154 591325 163918 591561
rect 164154 591325 170918 591561
rect 171154 591325 177918 591561
rect 178154 591325 184918 591561
rect 185154 591325 191918 591561
rect 192154 591325 198918 591561
rect 199154 591325 205918 591561
rect 206154 591325 212918 591561
rect 213154 591325 219918 591561
rect 220154 591325 226918 591561
rect 227154 591325 233918 591561
rect 234154 591325 240918 591561
rect 241154 591325 247918 591561
rect 248154 591325 254918 591561
rect 255154 591325 261918 591561
rect 262154 591325 268918 591561
rect 269154 591325 275918 591561
rect 276154 591325 282918 591561
rect 283154 591325 289918 591561
rect 290154 591325 296918 591561
rect 297154 591325 303918 591561
rect 304154 591325 310918 591561
rect 311154 591325 317918 591561
rect 318154 591325 324918 591561
rect 325154 591325 331918 591561
rect 332154 591325 338918 591561
rect 339154 591325 345918 591561
rect 346154 591325 352918 591561
rect 353154 591325 359918 591561
rect 360154 591325 366918 591561
rect 367154 591325 373918 591561
rect 374154 591325 380918 591561
rect 381154 591325 387918 591561
rect 388154 591325 394918 591561
rect 395154 591325 401918 591561
rect 402154 591325 408918 591561
rect 409154 591325 415918 591561
rect 416154 591325 422918 591561
rect 423154 591325 429918 591561
rect 430154 591325 436918 591561
rect 437154 591325 443918 591561
rect 444154 591325 450918 591561
rect 451154 591325 457918 591561
rect 458154 591325 464918 591561
rect 465154 591325 471918 591561
rect 472154 591325 478918 591561
rect 479154 591325 485918 591561
rect 486154 591325 492918 591561
rect 493154 591325 499918 591561
rect 500154 591325 506918 591561
rect 507154 591325 513918 591561
rect 514154 591325 520918 591561
rect 521154 591325 527918 591561
rect 528154 591325 534918 591561
rect 535154 591325 541918 591561
rect 542154 591325 548918 591561
rect 549154 591325 555918 591561
rect 556154 591325 562918 591561
rect 563154 591325 569918 591561
rect 570154 591325 576918 591561
rect 577154 591325 587570 591561
rect 587806 591325 587890 591561
rect 588126 591325 588210 591561
rect 588446 591325 588530 591561
rect 588766 591325 588874 591561
rect -4950 591283 588874 591325
rect -4950 590494 588874 590536
rect -4950 590258 -3090 590494
rect -2854 590258 -2770 590494
rect -2534 590258 -2450 590494
rect -2214 590258 -2130 590494
rect -1894 590258 1186 590494
rect 1422 590258 8186 590494
rect 8422 590258 15186 590494
rect 15422 590258 22186 590494
rect 22422 590258 29186 590494
rect 29422 590258 36186 590494
rect 36422 590258 43186 590494
rect 43422 590258 50186 590494
rect 50422 590258 57186 590494
rect 57422 590258 64186 590494
rect 64422 590258 71186 590494
rect 71422 590258 78186 590494
rect 78422 590258 85186 590494
rect 85422 590258 92186 590494
rect 92422 590258 99186 590494
rect 99422 590258 106186 590494
rect 106422 590258 113186 590494
rect 113422 590258 120186 590494
rect 120422 590258 127186 590494
rect 127422 590258 134186 590494
rect 134422 590258 141186 590494
rect 141422 590258 148186 590494
rect 148422 590258 155186 590494
rect 155422 590258 162186 590494
rect 162422 590258 169186 590494
rect 169422 590258 176186 590494
rect 176422 590258 183186 590494
rect 183422 590258 190186 590494
rect 190422 590258 197186 590494
rect 197422 590258 204186 590494
rect 204422 590258 211186 590494
rect 211422 590258 218186 590494
rect 218422 590258 225186 590494
rect 225422 590258 232186 590494
rect 232422 590258 239186 590494
rect 239422 590258 246186 590494
rect 246422 590258 253186 590494
rect 253422 590258 260186 590494
rect 260422 590258 267186 590494
rect 267422 590258 274186 590494
rect 274422 590258 281186 590494
rect 281422 590258 288186 590494
rect 288422 590258 295186 590494
rect 295422 590258 302186 590494
rect 302422 590258 309186 590494
rect 309422 590258 316186 590494
rect 316422 590258 323186 590494
rect 323422 590258 330186 590494
rect 330422 590258 337186 590494
rect 337422 590258 344186 590494
rect 344422 590258 351186 590494
rect 351422 590258 358186 590494
rect 358422 590258 365186 590494
rect 365422 590258 372186 590494
rect 372422 590258 379186 590494
rect 379422 590258 386186 590494
rect 386422 590258 393186 590494
rect 393422 590258 400186 590494
rect 400422 590258 407186 590494
rect 407422 590258 414186 590494
rect 414422 590258 421186 590494
rect 421422 590258 428186 590494
rect 428422 590258 435186 590494
rect 435422 590258 442186 590494
rect 442422 590258 449186 590494
rect 449422 590258 456186 590494
rect 456422 590258 463186 590494
rect 463422 590258 470186 590494
rect 470422 590258 477186 590494
rect 477422 590258 484186 590494
rect 484422 590258 491186 590494
rect 491422 590258 498186 590494
rect 498422 590258 505186 590494
rect 505422 590258 512186 590494
rect 512422 590258 519186 590494
rect 519422 590258 526186 590494
rect 526422 590258 533186 590494
rect 533422 590258 540186 590494
rect 540422 590258 547186 590494
rect 547422 590258 554186 590494
rect 554422 590258 561186 590494
rect 561422 590258 568186 590494
rect 568422 590258 575186 590494
rect 575422 590258 582186 590494
rect 582422 590258 585818 590494
rect 586054 590258 586138 590494
rect 586374 590258 586458 590494
rect 586694 590258 586778 590494
rect 587014 590258 588874 590494
rect -4950 590216 588874 590258
rect -4950 584561 588874 584603
rect -4950 584325 -4842 584561
rect -4606 584325 -4522 584561
rect -4286 584325 -4202 584561
rect -3966 584325 -3882 584561
rect -3646 584325 2918 584561
rect 3154 584325 9918 584561
rect 10154 584325 16918 584561
rect 17154 584325 23918 584561
rect 24154 584325 30918 584561
rect 31154 584325 37918 584561
rect 38154 584325 44918 584561
rect 45154 584325 51918 584561
rect 52154 584325 58918 584561
rect 59154 584325 65918 584561
rect 66154 584325 72918 584561
rect 73154 584325 79918 584561
rect 80154 584325 86918 584561
rect 87154 584325 93918 584561
rect 94154 584325 100918 584561
rect 101154 584325 107918 584561
rect 108154 584325 114918 584561
rect 115154 584325 121918 584561
rect 122154 584325 128918 584561
rect 129154 584325 135918 584561
rect 136154 584325 142918 584561
rect 143154 584325 149918 584561
rect 150154 584325 156918 584561
rect 157154 584325 163918 584561
rect 164154 584325 170918 584561
rect 171154 584325 177918 584561
rect 178154 584325 184918 584561
rect 185154 584325 191918 584561
rect 192154 584325 198918 584561
rect 199154 584325 205918 584561
rect 206154 584325 212918 584561
rect 213154 584325 219918 584561
rect 220154 584325 226918 584561
rect 227154 584325 233918 584561
rect 234154 584325 240918 584561
rect 241154 584325 247918 584561
rect 248154 584325 254918 584561
rect 255154 584325 261918 584561
rect 262154 584325 268918 584561
rect 269154 584325 275918 584561
rect 276154 584325 282918 584561
rect 283154 584325 289918 584561
rect 290154 584325 296918 584561
rect 297154 584325 303918 584561
rect 304154 584325 310918 584561
rect 311154 584325 317918 584561
rect 318154 584325 324918 584561
rect 325154 584325 331918 584561
rect 332154 584325 338918 584561
rect 339154 584325 345918 584561
rect 346154 584325 352918 584561
rect 353154 584325 359918 584561
rect 360154 584325 366918 584561
rect 367154 584325 373918 584561
rect 374154 584325 380918 584561
rect 381154 584325 387918 584561
rect 388154 584325 394918 584561
rect 395154 584325 401918 584561
rect 402154 584325 408918 584561
rect 409154 584325 415918 584561
rect 416154 584325 422918 584561
rect 423154 584325 429918 584561
rect 430154 584325 436918 584561
rect 437154 584325 443918 584561
rect 444154 584325 450918 584561
rect 451154 584325 457918 584561
rect 458154 584325 464918 584561
rect 465154 584325 471918 584561
rect 472154 584325 478918 584561
rect 479154 584325 485918 584561
rect 486154 584325 492918 584561
rect 493154 584325 499918 584561
rect 500154 584325 506918 584561
rect 507154 584325 513918 584561
rect 514154 584325 520918 584561
rect 521154 584325 527918 584561
rect 528154 584325 534918 584561
rect 535154 584325 541918 584561
rect 542154 584325 548918 584561
rect 549154 584325 555918 584561
rect 556154 584325 562918 584561
rect 563154 584325 569918 584561
rect 570154 584325 576918 584561
rect 577154 584325 587570 584561
rect 587806 584325 587890 584561
rect 588126 584325 588210 584561
rect 588446 584325 588530 584561
rect 588766 584325 588874 584561
rect -4950 584283 588874 584325
rect -4950 583494 588874 583536
rect -4950 583258 -3090 583494
rect -2854 583258 -2770 583494
rect -2534 583258 -2450 583494
rect -2214 583258 -2130 583494
rect -1894 583258 1186 583494
rect 1422 583258 8186 583494
rect 8422 583258 15186 583494
rect 15422 583258 22186 583494
rect 22422 583258 29186 583494
rect 29422 583258 36186 583494
rect 36422 583258 43186 583494
rect 43422 583258 50186 583494
rect 50422 583258 57186 583494
rect 57422 583258 64186 583494
rect 64422 583258 71186 583494
rect 71422 583258 78186 583494
rect 78422 583258 85186 583494
rect 85422 583258 92186 583494
rect 92422 583258 99186 583494
rect 99422 583258 106186 583494
rect 106422 583258 113186 583494
rect 113422 583258 120186 583494
rect 120422 583258 127186 583494
rect 127422 583258 134186 583494
rect 134422 583258 141186 583494
rect 141422 583258 148186 583494
rect 148422 583258 155186 583494
rect 155422 583258 162186 583494
rect 162422 583258 169186 583494
rect 169422 583258 176186 583494
rect 176422 583258 183186 583494
rect 183422 583258 190186 583494
rect 190422 583258 197186 583494
rect 197422 583258 204186 583494
rect 204422 583258 211186 583494
rect 211422 583258 218186 583494
rect 218422 583258 225186 583494
rect 225422 583258 232186 583494
rect 232422 583258 239186 583494
rect 239422 583258 246186 583494
rect 246422 583258 253186 583494
rect 253422 583258 260186 583494
rect 260422 583258 267186 583494
rect 267422 583258 274186 583494
rect 274422 583258 281186 583494
rect 281422 583258 288186 583494
rect 288422 583258 295186 583494
rect 295422 583258 302186 583494
rect 302422 583258 309186 583494
rect 309422 583258 316186 583494
rect 316422 583258 323186 583494
rect 323422 583258 330186 583494
rect 330422 583258 337186 583494
rect 337422 583258 344186 583494
rect 344422 583258 351186 583494
rect 351422 583258 358186 583494
rect 358422 583258 365186 583494
rect 365422 583258 372186 583494
rect 372422 583258 379186 583494
rect 379422 583258 386186 583494
rect 386422 583258 393186 583494
rect 393422 583258 400186 583494
rect 400422 583258 407186 583494
rect 407422 583258 414186 583494
rect 414422 583258 421186 583494
rect 421422 583258 428186 583494
rect 428422 583258 435186 583494
rect 435422 583258 442186 583494
rect 442422 583258 449186 583494
rect 449422 583258 456186 583494
rect 456422 583258 463186 583494
rect 463422 583258 470186 583494
rect 470422 583258 477186 583494
rect 477422 583258 484186 583494
rect 484422 583258 491186 583494
rect 491422 583258 498186 583494
rect 498422 583258 505186 583494
rect 505422 583258 512186 583494
rect 512422 583258 519186 583494
rect 519422 583258 526186 583494
rect 526422 583258 533186 583494
rect 533422 583258 540186 583494
rect 540422 583258 547186 583494
rect 547422 583258 554186 583494
rect 554422 583258 561186 583494
rect 561422 583258 568186 583494
rect 568422 583258 575186 583494
rect 575422 583258 582186 583494
rect 582422 583258 585818 583494
rect 586054 583258 586138 583494
rect 586374 583258 586458 583494
rect 586694 583258 586778 583494
rect 587014 583258 588874 583494
rect -4950 583216 588874 583258
rect -4950 577561 588874 577603
rect -4950 577325 -4842 577561
rect -4606 577325 -4522 577561
rect -4286 577325 -4202 577561
rect -3966 577325 -3882 577561
rect -3646 577325 2918 577561
rect 3154 577325 9918 577561
rect 10154 577325 16918 577561
rect 17154 577325 23918 577561
rect 24154 577325 30918 577561
rect 31154 577325 37918 577561
rect 38154 577325 44918 577561
rect 45154 577325 51918 577561
rect 52154 577325 58918 577561
rect 59154 577325 65918 577561
rect 66154 577325 72918 577561
rect 73154 577325 79918 577561
rect 80154 577325 86918 577561
rect 87154 577325 93918 577561
rect 94154 577325 100918 577561
rect 101154 577325 107918 577561
rect 108154 577325 114918 577561
rect 115154 577325 121918 577561
rect 122154 577325 128918 577561
rect 129154 577325 135918 577561
rect 136154 577325 142918 577561
rect 143154 577325 149918 577561
rect 150154 577325 156918 577561
rect 157154 577325 163918 577561
rect 164154 577325 170918 577561
rect 171154 577325 177918 577561
rect 178154 577325 184918 577561
rect 185154 577325 191918 577561
rect 192154 577325 198918 577561
rect 199154 577325 205918 577561
rect 206154 577325 212918 577561
rect 213154 577325 219918 577561
rect 220154 577325 226918 577561
rect 227154 577325 233918 577561
rect 234154 577325 240918 577561
rect 241154 577325 247918 577561
rect 248154 577325 254918 577561
rect 255154 577325 261918 577561
rect 262154 577325 268918 577561
rect 269154 577325 275918 577561
rect 276154 577325 282918 577561
rect 283154 577325 289918 577561
rect 290154 577325 296918 577561
rect 297154 577325 303918 577561
rect 304154 577325 310918 577561
rect 311154 577325 317918 577561
rect 318154 577325 324918 577561
rect 325154 577325 331918 577561
rect 332154 577325 338918 577561
rect 339154 577325 345918 577561
rect 346154 577325 352918 577561
rect 353154 577325 359918 577561
rect 360154 577325 366918 577561
rect 367154 577325 373918 577561
rect 374154 577325 380918 577561
rect 381154 577325 387918 577561
rect 388154 577325 394918 577561
rect 395154 577325 401918 577561
rect 402154 577325 408918 577561
rect 409154 577325 415918 577561
rect 416154 577325 422918 577561
rect 423154 577325 429918 577561
rect 430154 577325 436918 577561
rect 437154 577325 443918 577561
rect 444154 577325 450918 577561
rect 451154 577325 457918 577561
rect 458154 577325 464918 577561
rect 465154 577325 471918 577561
rect 472154 577325 478918 577561
rect 479154 577325 485918 577561
rect 486154 577325 492918 577561
rect 493154 577325 499918 577561
rect 500154 577325 506918 577561
rect 507154 577325 513918 577561
rect 514154 577325 520918 577561
rect 521154 577325 527918 577561
rect 528154 577325 534918 577561
rect 535154 577325 541918 577561
rect 542154 577325 548918 577561
rect 549154 577325 555918 577561
rect 556154 577325 562918 577561
rect 563154 577325 569918 577561
rect 570154 577325 576918 577561
rect 577154 577325 587570 577561
rect 587806 577325 587890 577561
rect 588126 577325 588210 577561
rect 588446 577325 588530 577561
rect 588766 577325 588874 577561
rect -4950 577283 588874 577325
rect -4950 576494 588874 576536
rect -4950 576258 -3090 576494
rect -2854 576258 -2770 576494
rect -2534 576258 -2450 576494
rect -2214 576258 -2130 576494
rect -1894 576258 1186 576494
rect 1422 576258 8186 576494
rect 8422 576258 15186 576494
rect 15422 576258 22186 576494
rect 22422 576258 29186 576494
rect 29422 576258 36186 576494
rect 36422 576258 43186 576494
rect 43422 576258 50186 576494
rect 50422 576258 57186 576494
rect 57422 576258 64186 576494
rect 64422 576258 71186 576494
rect 71422 576258 78186 576494
rect 78422 576258 85186 576494
rect 85422 576258 92186 576494
rect 92422 576258 99186 576494
rect 99422 576258 106186 576494
rect 106422 576258 113186 576494
rect 113422 576258 120186 576494
rect 120422 576258 127186 576494
rect 127422 576258 134186 576494
rect 134422 576258 141186 576494
rect 141422 576258 148186 576494
rect 148422 576258 155186 576494
rect 155422 576258 162186 576494
rect 162422 576258 169186 576494
rect 169422 576258 176186 576494
rect 176422 576258 183186 576494
rect 183422 576258 190186 576494
rect 190422 576258 197186 576494
rect 197422 576258 204186 576494
rect 204422 576258 211186 576494
rect 211422 576258 218186 576494
rect 218422 576258 225186 576494
rect 225422 576258 232186 576494
rect 232422 576258 239186 576494
rect 239422 576258 246186 576494
rect 246422 576258 253186 576494
rect 253422 576258 260186 576494
rect 260422 576258 267186 576494
rect 267422 576258 274186 576494
rect 274422 576258 281186 576494
rect 281422 576258 288186 576494
rect 288422 576258 295186 576494
rect 295422 576258 302186 576494
rect 302422 576258 309186 576494
rect 309422 576258 316186 576494
rect 316422 576258 323186 576494
rect 323422 576258 330186 576494
rect 330422 576258 337186 576494
rect 337422 576258 344186 576494
rect 344422 576258 351186 576494
rect 351422 576258 358186 576494
rect 358422 576258 365186 576494
rect 365422 576258 372186 576494
rect 372422 576258 379186 576494
rect 379422 576258 386186 576494
rect 386422 576258 393186 576494
rect 393422 576258 400186 576494
rect 400422 576258 407186 576494
rect 407422 576258 414186 576494
rect 414422 576258 421186 576494
rect 421422 576258 428186 576494
rect 428422 576258 435186 576494
rect 435422 576258 442186 576494
rect 442422 576258 449186 576494
rect 449422 576258 456186 576494
rect 456422 576258 463186 576494
rect 463422 576258 470186 576494
rect 470422 576258 477186 576494
rect 477422 576258 484186 576494
rect 484422 576258 491186 576494
rect 491422 576258 498186 576494
rect 498422 576258 505186 576494
rect 505422 576258 512186 576494
rect 512422 576258 519186 576494
rect 519422 576258 526186 576494
rect 526422 576258 533186 576494
rect 533422 576258 540186 576494
rect 540422 576258 547186 576494
rect 547422 576258 554186 576494
rect 554422 576258 561186 576494
rect 561422 576258 568186 576494
rect 568422 576258 575186 576494
rect 575422 576258 582186 576494
rect 582422 576258 585818 576494
rect 586054 576258 586138 576494
rect 586374 576258 586458 576494
rect 586694 576258 586778 576494
rect 587014 576258 588874 576494
rect -4950 576216 588874 576258
rect -4950 570561 588874 570603
rect -4950 570325 -4842 570561
rect -4606 570325 -4522 570561
rect -4286 570325 -4202 570561
rect -3966 570325 -3882 570561
rect -3646 570325 2918 570561
rect 3154 570325 9918 570561
rect 10154 570325 16918 570561
rect 17154 570325 23918 570561
rect 24154 570325 30918 570561
rect 31154 570325 37918 570561
rect 38154 570325 44918 570561
rect 45154 570325 51918 570561
rect 52154 570325 58918 570561
rect 59154 570325 65918 570561
rect 66154 570325 72918 570561
rect 73154 570325 79918 570561
rect 80154 570325 86918 570561
rect 87154 570325 93918 570561
rect 94154 570325 100918 570561
rect 101154 570325 107918 570561
rect 108154 570325 114918 570561
rect 115154 570325 121918 570561
rect 122154 570325 128918 570561
rect 129154 570325 135918 570561
rect 136154 570325 142918 570561
rect 143154 570325 149918 570561
rect 150154 570325 156918 570561
rect 157154 570325 163918 570561
rect 164154 570325 170918 570561
rect 171154 570325 177918 570561
rect 178154 570325 184918 570561
rect 185154 570325 191918 570561
rect 192154 570325 198918 570561
rect 199154 570325 205918 570561
rect 206154 570325 212918 570561
rect 213154 570325 219918 570561
rect 220154 570325 226918 570561
rect 227154 570325 233918 570561
rect 234154 570325 240918 570561
rect 241154 570325 247918 570561
rect 248154 570325 254918 570561
rect 255154 570325 261918 570561
rect 262154 570325 268918 570561
rect 269154 570325 275918 570561
rect 276154 570325 282918 570561
rect 283154 570325 289918 570561
rect 290154 570325 296918 570561
rect 297154 570325 303918 570561
rect 304154 570325 310918 570561
rect 311154 570325 317918 570561
rect 318154 570325 324918 570561
rect 325154 570325 331918 570561
rect 332154 570325 338918 570561
rect 339154 570325 345918 570561
rect 346154 570325 352918 570561
rect 353154 570325 359918 570561
rect 360154 570325 366918 570561
rect 367154 570325 373918 570561
rect 374154 570325 380918 570561
rect 381154 570325 387918 570561
rect 388154 570325 394918 570561
rect 395154 570325 401918 570561
rect 402154 570325 408918 570561
rect 409154 570325 415918 570561
rect 416154 570325 422918 570561
rect 423154 570325 429918 570561
rect 430154 570325 436918 570561
rect 437154 570325 443918 570561
rect 444154 570325 450918 570561
rect 451154 570325 457918 570561
rect 458154 570325 464918 570561
rect 465154 570325 471918 570561
rect 472154 570325 478918 570561
rect 479154 570325 485918 570561
rect 486154 570325 492918 570561
rect 493154 570325 499918 570561
rect 500154 570325 506918 570561
rect 507154 570325 513918 570561
rect 514154 570325 520918 570561
rect 521154 570325 527918 570561
rect 528154 570325 534918 570561
rect 535154 570325 541918 570561
rect 542154 570325 548918 570561
rect 549154 570325 555918 570561
rect 556154 570325 562918 570561
rect 563154 570325 569918 570561
rect 570154 570325 576918 570561
rect 577154 570325 587570 570561
rect 587806 570325 587890 570561
rect 588126 570325 588210 570561
rect 588446 570325 588530 570561
rect 588766 570325 588874 570561
rect -4950 570283 588874 570325
rect -4950 569494 588874 569536
rect -4950 569258 -3090 569494
rect -2854 569258 -2770 569494
rect -2534 569258 -2450 569494
rect -2214 569258 -2130 569494
rect -1894 569258 1186 569494
rect 1422 569258 8186 569494
rect 8422 569258 15186 569494
rect 15422 569258 22186 569494
rect 22422 569258 29186 569494
rect 29422 569258 36186 569494
rect 36422 569258 43186 569494
rect 43422 569258 50186 569494
rect 50422 569258 57186 569494
rect 57422 569258 64186 569494
rect 64422 569258 71186 569494
rect 71422 569258 78186 569494
rect 78422 569258 85186 569494
rect 85422 569258 92186 569494
rect 92422 569258 99186 569494
rect 99422 569258 106186 569494
rect 106422 569258 113186 569494
rect 113422 569258 120186 569494
rect 120422 569258 127186 569494
rect 127422 569258 134186 569494
rect 134422 569258 141186 569494
rect 141422 569258 148186 569494
rect 148422 569258 155186 569494
rect 155422 569258 162186 569494
rect 162422 569258 169186 569494
rect 169422 569258 176186 569494
rect 176422 569258 183186 569494
rect 183422 569258 190186 569494
rect 190422 569258 197186 569494
rect 197422 569258 204186 569494
rect 204422 569258 211186 569494
rect 211422 569258 218186 569494
rect 218422 569258 225186 569494
rect 225422 569258 232186 569494
rect 232422 569258 239186 569494
rect 239422 569258 246186 569494
rect 246422 569258 253186 569494
rect 253422 569258 260186 569494
rect 260422 569258 267186 569494
rect 267422 569258 274186 569494
rect 274422 569258 281186 569494
rect 281422 569258 288186 569494
rect 288422 569258 295186 569494
rect 295422 569258 302186 569494
rect 302422 569258 309186 569494
rect 309422 569258 316186 569494
rect 316422 569258 323186 569494
rect 323422 569258 330186 569494
rect 330422 569258 337186 569494
rect 337422 569258 344186 569494
rect 344422 569258 351186 569494
rect 351422 569258 358186 569494
rect 358422 569258 365186 569494
rect 365422 569258 372186 569494
rect 372422 569258 379186 569494
rect 379422 569258 386186 569494
rect 386422 569258 393186 569494
rect 393422 569258 400186 569494
rect 400422 569258 407186 569494
rect 407422 569258 414186 569494
rect 414422 569258 421186 569494
rect 421422 569258 428186 569494
rect 428422 569258 435186 569494
rect 435422 569258 442186 569494
rect 442422 569258 449186 569494
rect 449422 569258 456186 569494
rect 456422 569258 463186 569494
rect 463422 569258 470186 569494
rect 470422 569258 477186 569494
rect 477422 569258 484186 569494
rect 484422 569258 491186 569494
rect 491422 569258 498186 569494
rect 498422 569258 505186 569494
rect 505422 569258 512186 569494
rect 512422 569258 519186 569494
rect 519422 569258 526186 569494
rect 526422 569258 533186 569494
rect 533422 569258 540186 569494
rect 540422 569258 547186 569494
rect 547422 569258 554186 569494
rect 554422 569258 561186 569494
rect 561422 569258 568186 569494
rect 568422 569258 575186 569494
rect 575422 569258 582186 569494
rect 582422 569258 585818 569494
rect 586054 569258 586138 569494
rect 586374 569258 586458 569494
rect 586694 569258 586778 569494
rect 587014 569258 588874 569494
rect -4950 569216 588874 569258
rect -4950 563561 588874 563603
rect -4950 563325 -4842 563561
rect -4606 563325 -4522 563561
rect -4286 563325 -4202 563561
rect -3966 563325 -3882 563561
rect -3646 563325 2918 563561
rect 3154 563325 9918 563561
rect 10154 563325 16918 563561
rect 17154 563325 23918 563561
rect 24154 563325 30918 563561
rect 31154 563325 37918 563561
rect 38154 563325 44918 563561
rect 45154 563325 51918 563561
rect 52154 563325 58918 563561
rect 59154 563325 65918 563561
rect 66154 563325 72918 563561
rect 73154 563325 79918 563561
rect 80154 563325 86918 563561
rect 87154 563325 93918 563561
rect 94154 563325 100918 563561
rect 101154 563325 107918 563561
rect 108154 563325 114918 563561
rect 115154 563325 121918 563561
rect 122154 563325 128918 563561
rect 129154 563325 135918 563561
rect 136154 563325 142918 563561
rect 143154 563325 149918 563561
rect 150154 563325 156918 563561
rect 157154 563325 163918 563561
rect 164154 563325 170918 563561
rect 171154 563325 177918 563561
rect 178154 563325 184918 563561
rect 185154 563325 191918 563561
rect 192154 563325 198918 563561
rect 199154 563325 205918 563561
rect 206154 563325 212918 563561
rect 213154 563325 219918 563561
rect 220154 563325 226918 563561
rect 227154 563325 233918 563561
rect 234154 563325 240918 563561
rect 241154 563325 247918 563561
rect 248154 563325 254918 563561
rect 255154 563325 261918 563561
rect 262154 563325 268918 563561
rect 269154 563325 275918 563561
rect 276154 563325 282918 563561
rect 283154 563325 289918 563561
rect 290154 563325 296918 563561
rect 297154 563325 303918 563561
rect 304154 563325 310918 563561
rect 311154 563325 317918 563561
rect 318154 563325 324918 563561
rect 325154 563325 331918 563561
rect 332154 563325 338918 563561
rect 339154 563325 345918 563561
rect 346154 563325 352918 563561
rect 353154 563325 359918 563561
rect 360154 563325 366918 563561
rect 367154 563325 373918 563561
rect 374154 563325 380918 563561
rect 381154 563325 387918 563561
rect 388154 563325 394918 563561
rect 395154 563325 401918 563561
rect 402154 563325 408918 563561
rect 409154 563325 415918 563561
rect 416154 563325 422918 563561
rect 423154 563325 429918 563561
rect 430154 563325 436918 563561
rect 437154 563325 443918 563561
rect 444154 563325 450918 563561
rect 451154 563325 457918 563561
rect 458154 563325 464918 563561
rect 465154 563325 471918 563561
rect 472154 563325 478918 563561
rect 479154 563325 485918 563561
rect 486154 563325 492918 563561
rect 493154 563325 499918 563561
rect 500154 563325 506918 563561
rect 507154 563325 513918 563561
rect 514154 563325 520918 563561
rect 521154 563325 527918 563561
rect 528154 563325 534918 563561
rect 535154 563325 541918 563561
rect 542154 563325 548918 563561
rect 549154 563325 555918 563561
rect 556154 563325 562918 563561
rect 563154 563325 569918 563561
rect 570154 563325 576918 563561
rect 577154 563325 587570 563561
rect 587806 563325 587890 563561
rect 588126 563325 588210 563561
rect 588446 563325 588530 563561
rect 588766 563325 588874 563561
rect -4950 563283 588874 563325
rect -4950 562494 588874 562536
rect -4950 562258 -3090 562494
rect -2854 562258 -2770 562494
rect -2534 562258 -2450 562494
rect -2214 562258 -2130 562494
rect -1894 562258 1186 562494
rect 1422 562258 8186 562494
rect 8422 562258 15186 562494
rect 15422 562258 22186 562494
rect 22422 562258 29186 562494
rect 29422 562258 36186 562494
rect 36422 562258 43186 562494
rect 43422 562258 50186 562494
rect 50422 562258 57186 562494
rect 57422 562258 64186 562494
rect 64422 562258 71186 562494
rect 71422 562258 78186 562494
rect 78422 562258 85186 562494
rect 85422 562258 92186 562494
rect 92422 562258 99186 562494
rect 99422 562258 106186 562494
rect 106422 562258 113186 562494
rect 113422 562258 120186 562494
rect 120422 562258 127186 562494
rect 127422 562258 134186 562494
rect 134422 562258 141186 562494
rect 141422 562258 148186 562494
rect 148422 562258 155186 562494
rect 155422 562258 162186 562494
rect 162422 562258 169186 562494
rect 169422 562258 176186 562494
rect 176422 562258 183186 562494
rect 183422 562258 190186 562494
rect 190422 562258 197186 562494
rect 197422 562258 204186 562494
rect 204422 562258 211186 562494
rect 211422 562258 218186 562494
rect 218422 562258 225186 562494
rect 225422 562258 232186 562494
rect 232422 562258 239186 562494
rect 239422 562258 246186 562494
rect 246422 562258 253186 562494
rect 253422 562258 260186 562494
rect 260422 562258 267186 562494
rect 267422 562258 274186 562494
rect 274422 562258 281186 562494
rect 281422 562258 288186 562494
rect 288422 562258 295186 562494
rect 295422 562258 302186 562494
rect 302422 562258 309186 562494
rect 309422 562258 316186 562494
rect 316422 562258 323186 562494
rect 323422 562258 330186 562494
rect 330422 562258 337186 562494
rect 337422 562258 344186 562494
rect 344422 562258 351186 562494
rect 351422 562258 358186 562494
rect 358422 562258 365186 562494
rect 365422 562258 372186 562494
rect 372422 562258 379186 562494
rect 379422 562258 386186 562494
rect 386422 562258 393186 562494
rect 393422 562258 400186 562494
rect 400422 562258 407186 562494
rect 407422 562258 414186 562494
rect 414422 562258 421186 562494
rect 421422 562258 428186 562494
rect 428422 562258 435186 562494
rect 435422 562258 442186 562494
rect 442422 562258 449186 562494
rect 449422 562258 456186 562494
rect 456422 562258 463186 562494
rect 463422 562258 470186 562494
rect 470422 562258 477186 562494
rect 477422 562258 484186 562494
rect 484422 562258 491186 562494
rect 491422 562258 498186 562494
rect 498422 562258 505186 562494
rect 505422 562258 512186 562494
rect 512422 562258 519186 562494
rect 519422 562258 526186 562494
rect 526422 562258 533186 562494
rect 533422 562258 540186 562494
rect 540422 562258 547186 562494
rect 547422 562258 554186 562494
rect 554422 562258 561186 562494
rect 561422 562258 568186 562494
rect 568422 562258 575186 562494
rect 575422 562258 582186 562494
rect 582422 562258 585818 562494
rect 586054 562258 586138 562494
rect 586374 562258 586458 562494
rect 586694 562258 586778 562494
rect 587014 562258 588874 562494
rect -4950 562216 588874 562258
rect -4950 556561 588874 556603
rect -4950 556325 -4842 556561
rect -4606 556325 -4522 556561
rect -4286 556325 -4202 556561
rect -3966 556325 -3882 556561
rect -3646 556325 2918 556561
rect 3154 556325 9918 556561
rect 10154 556325 16918 556561
rect 17154 556325 23918 556561
rect 24154 556325 30918 556561
rect 31154 556325 37918 556561
rect 38154 556325 44918 556561
rect 45154 556325 51918 556561
rect 52154 556325 58918 556561
rect 59154 556325 65918 556561
rect 66154 556325 72918 556561
rect 73154 556325 79918 556561
rect 80154 556325 86918 556561
rect 87154 556325 93918 556561
rect 94154 556325 100918 556561
rect 101154 556325 107918 556561
rect 108154 556325 114918 556561
rect 115154 556325 121918 556561
rect 122154 556325 128918 556561
rect 129154 556325 135918 556561
rect 136154 556325 142918 556561
rect 143154 556325 149918 556561
rect 150154 556325 156918 556561
rect 157154 556325 163918 556561
rect 164154 556325 170918 556561
rect 171154 556325 177918 556561
rect 178154 556325 184918 556561
rect 185154 556325 191918 556561
rect 192154 556325 198918 556561
rect 199154 556325 205918 556561
rect 206154 556325 212918 556561
rect 213154 556325 219918 556561
rect 220154 556325 226918 556561
rect 227154 556325 233918 556561
rect 234154 556325 240918 556561
rect 241154 556325 247918 556561
rect 248154 556325 254918 556561
rect 255154 556325 261918 556561
rect 262154 556325 268918 556561
rect 269154 556325 275918 556561
rect 276154 556325 282918 556561
rect 283154 556325 289918 556561
rect 290154 556325 296918 556561
rect 297154 556325 303918 556561
rect 304154 556325 310918 556561
rect 311154 556325 317918 556561
rect 318154 556325 324918 556561
rect 325154 556325 331918 556561
rect 332154 556325 338918 556561
rect 339154 556325 345918 556561
rect 346154 556325 352918 556561
rect 353154 556325 359918 556561
rect 360154 556325 366918 556561
rect 367154 556325 373918 556561
rect 374154 556325 380918 556561
rect 381154 556325 387918 556561
rect 388154 556325 394918 556561
rect 395154 556325 401918 556561
rect 402154 556325 408918 556561
rect 409154 556325 415918 556561
rect 416154 556325 422918 556561
rect 423154 556325 429918 556561
rect 430154 556325 436918 556561
rect 437154 556325 443918 556561
rect 444154 556325 450918 556561
rect 451154 556325 457918 556561
rect 458154 556325 464918 556561
rect 465154 556325 471918 556561
rect 472154 556325 478918 556561
rect 479154 556325 485918 556561
rect 486154 556325 492918 556561
rect 493154 556325 499918 556561
rect 500154 556325 506918 556561
rect 507154 556325 513918 556561
rect 514154 556325 520918 556561
rect 521154 556325 527918 556561
rect 528154 556325 534918 556561
rect 535154 556325 541918 556561
rect 542154 556325 548918 556561
rect 549154 556325 555918 556561
rect 556154 556325 562918 556561
rect 563154 556325 569918 556561
rect 570154 556325 576918 556561
rect 577154 556325 587570 556561
rect 587806 556325 587890 556561
rect 588126 556325 588210 556561
rect 588446 556325 588530 556561
rect 588766 556325 588874 556561
rect -4950 556283 588874 556325
rect -4950 555494 588874 555536
rect -4950 555258 -3090 555494
rect -2854 555258 -2770 555494
rect -2534 555258 -2450 555494
rect -2214 555258 -2130 555494
rect -1894 555258 1186 555494
rect 1422 555258 8186 555494
rect 8422 555258 15186 555494
rect 15422 555258 22186 555494
rect 22422 555258 29186 555494
rect 29422 555258 36186 555494
rect 36422 555258 43186 555494
rect 43422 555258 50186 555494
rect 50422 555258 57186 555494
rect 57422 555258 64186 555494
rect 64422 555258 71186 555494
rect 71422 555258 78186 555494
rect 78422 555258 85186 555494
rect 85422 555258 92186 555494
rect 92422 555258 99186 555494
rect 99422 555258 106186 555494
rect 106422 555258 113186 555494
rect 113422 555258 120186 555494
rect 120422 555258 127186 555494
rect 127422 555258 134186 555494
rect 134422 555258 141186 555494
rect 141422 555258 148186 555494
rect 148422 555258 155186 555494
rect 155422 555258 162186 555494
rect 162422 555258 169186 555494
rect 169422 555258 176186 555494
rect 176422 555258 183186 555494
rect 183422 555258 190186 555494
rect 190422 555258 197186 555494
rect 197422 555258 204186 555494
rect 204422 555258 211186 555494
rect 211422 555258 218186 555494
rect 218422 555258 225186 555494
rect 225422 555258 232186 555494
rect 232422 555258 239186 555494
rect 239422 555258 246186 555494
rect 246422 555258 253186 555494
rect 253422 555258 260186 555494
rect 260422 555258 267186 555494
rect 267422 555258 274186 555494
rect 274422 555258 281186 555494
rect 281422 555258 288186 555494
rect 288422 555258 295186 555494
rect 295422 555258 302186 555494
rect 302422 555258 309186 555494
rect 309422 555258 316186 555494
rect 316422 555258 323186 555494
rect 323422 555258 330186 555494
rect 330422 555258 337186 555494
rect 337422 555258 344186 555494
rect 344422 555258 351186 555494
rect 351422 555258 358186 555494
rect 358422 555258 365186 555494
rect 365422 555258 372186 555494
rect 372422 555258 379186 555494
rect 379422 555258 386186 555494
rect 386422 555258 393186 555494
rect 393422 555258 400186 555494
rect 400422 555258 407186 555494
rect 407422 555258 414186 555494
rect 414422 555258 421186 555494
rect 421422 555258 428186 555494
rect 428422 555258 435186 555494
rect 435422 555258 442186 555494
rect 442422 555258 449186 555494
rect 449422 555258 456186 555494
rect 456422 555258 463186 555494
rect 463422 555258 470186 555494
rect 470422 555258 477186 555494
rect 477422 555258 484186 555494
rect 484422 555258 491186 555494
rect 491422 555258 498186 555494
rect 498422 555258 505186 555494
rect 505422 555258 512186 555494
rect 512422 555258 519186 555494
rect 519422 555258 526186 555494
rect 526422 555258 533186 555494
rect 533422 555258 540186 555494
rect 540422 555258 547186 555494
rect 547422 555258 554186 555494
rect 554422 555258 561186 555494
rect 561422 555258 568186 555494
rect 568422 555258 575186 555494
rect 575422 555258 582186 555494
rect 582422 555258 585818 555494
rect 586054 555258 586138 555494
rect 586374 555258 586458 555494
rect 586694 555258 586778 555494
rect 587014 555258 588874 555494
rect -4950 555216 588874 555258
rect -4950 549561 588874 549603
rect -4950 549325 -4842 549561
rect -4606 549325 -4522 549561
rect -4286 549325 -4202 549561
rect -3966 549325 -3882 549561
rect -3646 549325 2918 549561
rect 3154 549325 9918 549561
rect 10154 549325 16918 549561
rect 17154 549325 23918 549561
rect 24154 549325 30918 549561
rect 31154 549325 37918 549561
rect 38154 549325 44918 549561
rect 45154 549325 51918 549561
rect 52154 549325 58918 549561
rect 59154 549325 65918 549561
rect 66154 549325 72918 549561
rect 73154 549325 79918 549561
rect 80154 549325 86918 549561
rect 87154 549325 93918 549561
rect 94154 549325 100918 549561
rect 101154 549325 107918 549561
rect 108154 549325 114918 549561
rect 115154 549325 121918 549561
rect 122154 549325 128918 549561
rect 129154 549325 135918 549561
rect 136154 549325 142918 549561
rect 143154 549325 149918 549561
rect 150154 549325 156918 549561
rect 157154 549325 163918 549561
rect 164154 549325 170918 549561
rect 171154 549325 177918 549561
rect 178154 549325 184918 549561
rect 185154 549325 191918 549561
rect 192154 549325 198918 549561
rect 199154 549325 205918 549561
rect 206154 549325 212918 549561
rect 213154 549325 219918 549561
rect 220154 549325 226918 549561
rect 227154 549325 233918 549561
rect 234154 549325 240918 549561
rect 241154 549325 247918 549561
rect 248154 549325 254918 549561
rect 255154 549325 261918 549561
rect 262154 549325 268918 549561
rect 269154 549325 275918 549561
rect 276154 549325 282918 549561
rect 283154 549325 289918 549561
rect 290154 549325 296918 549561
rect 297154 549325 303918 549561
rect 304154 549325 310918 549561
rect 311154 549325 317918 549561
rect 318154 549325 324918 549561
rect 325154 549325 331918 549561
rect 332154 549325 338918 549561
rect 339154 549325 345918 549561
rect 346154 549325 352918 549561
rect 353154 549325 359918 549561
rect 360154 549325 366918 549561
rect 367154 549325 373918 549561
rect 374154 549325 380918 549561
rect 381154 549325 387918 549561
rect 388154 549325 394918 549561
rect 395154 549325 401918 549561
rect 402154 549325 408918 549561
rect 409154 549325 415918 549561
rect 416154 549325 422918 549561
rect 423154 549325 429918 549561
rect 430154 549325 436918 549561
rect 437154 549325 443918 549561
rect 444154 549325 450918 549561
rect 451154 549325 457918 549561
rect 458154 549325 464918 549561
rect 465154 549325 471918 549561
rect 472154 549325 478918 549561
rect 479154 549325 485918 549561
rect 486154 549325 492918 549561
rect 493154 549325 499918 549561
rect 500154 549325 506918 549561
rect 507154 549325 513918 549561
rect 514154 549325 520918 549561
rect 521154 549325 527918 549561
rect 528154 549325 534918 549561
rect 535154 549325 541918 549561
rect 542154 549325 548918 549561
rect 549154 549325 555918 549561
rect 556154 549325 562918 549561
rect 563154 549325 569918 549561
rect 570154 549325 576918 549561
rect 577154 549325 587570 549561
rect 587806 549325 587890 549561
rect 588126 549325 588210 549561
rect 588446 549325 588530 549561
rect 588766 549325 588874 549561
rect -4950 549283 588874 549325
rect -4950 548494 588874 548536
rect -4950 548258 -3090 548494
rect -2854 548258 -2770 548494
rect -2534 548258 -2450 548494
rect -2214 548258 -2130 548494
rect -1894 548258 1186 548494
rect 1422 548258 8186 548494
rect 8422 548258 15186 548494
rect 15422 548258 22186 548494
rect 22422 548258 29186 548494
rect 29422 548258 36186 548494
rect 36422 548258 43186 548494
rect 43422 548258 50186 548494
rect 50422 548258 57186 548494
rect 57422 548258 64186 548494
rect 64422 548258 71186 548494
rect 71422 548258 78186 548494
rect 78422 548258 85186 548494
rect 85422 548258 92186 548494
rect 92422 548258 99186 548494
rect 99422 548258 106186 548494
rect 106422 548258 113186 548494
rect 113422 548258 120186 548494
rect 120422 548258 127186 548494
rect 127422 548258 134186 548494
rect 134422 548258 141186 548494
rect 141422 548258 148186 548494
rect 148422 548258 155186 548494
rect 155422 548258 162186 548494
rect 162422 548258 169186 548494
rect 169422 548258 176186 548494
rect 176422 548258 183186 548494
rect 183422 548258 190186 548494
rect 190422 548258 197186 548494
rect 197422 548258 204186 548494
rect 204422 548258 211186 548494
rect 211422 548258 218186 548494
rect 218422 548258 225186 548494
rect 225422 548258 232186 548494
rect 232422 548258 239186 548494
rect 239422 548258 246186 548494
rect 246422 548258 253186 548494
rect 253422 548258 260186 548494
rect 260422 548258 267186 548494
rect 267422 548258 274186 548494
rect 274422 548258 281186 548494
rect 281422 548258 288186 548494
rect 288422 548258 295186 548494
rect 295422 548258 302186 548494
rect 302422 548258 309186 548494
rect 309422 548258 316186 548494
rect 316422 548258 323186 548494
rect 323422 548258 330186 548494
rect 330422 548258 337186 548494
rect 337422 548258 344186 548494
rect 344422 548258 351186 548494
rect 351422 548258 358186 548494
rect 358422 548258 365186 548494
rect 365422 548258 372186 548494
rect 372422 548258 379186 548494
rect 379422 548258 386186 548494
rect 386422 548258 393186 548494
rect 393422 548258 400186 548494
rect 400422 548258 407186 548494
rect 407422 548258 414186 548494
rect 414422 548258 421186 548494
rect 421422 548258 428186 548494
rect 428422 548258 435186 548494
rect 435422 548258 442186 548494
rect 442422 548258 449186 548494
rect 449422 548258 456186 548494
rect 456422 548258 463186 548494
rect 463422 548258 470186 548494
rect 470422 548258 477186 548494
rect 477422 548258 484186 548494
rect 484422 548258 491186 548494
rect 491422 548258 498186 548494
rect 498422 548258 505186 548494
rect 505422 548258 512186 548494
rect 512422 548258 519186 548494
rect 519422 548258 526186 548494
rect 526422 548258 533186 548494
rect 533422 548258 540186 548494
rect 540422 548258 547186 548494
rect 547422 548258 554186 548494
rect 554422 548258 561186 548494
rect 561422 548258 568186 548494
rect 568422 548258 575186 548494
rect 575422 548258 582186 548494
rect 582422 548258 585818 548494
rect 586054 548258 586138 548494
rect 586374 548258 586458 548494
rect 586694 548258 586778 548494
rect 587014 548258 588874 548494
rect -4950 548216 588874 548258
rect -4950 542561 588874 542603
rect -4950 542325 -4842 542561
rect -4606 542325 -4522 542561
rect -4286 542325 -4202 542561
rect -3966 542325 -3882 542561
rect -3646 542325 2918 542561
rect 3154 542325 9918 542561
rect 10154 542325 16918 542561
rect 17154 542325 23918 542561
rect 24154 542325 30918 542561
rect 31154 542325 37918 542561
rect 38154 542325 44918 542561
rect 45154 542325 51918 542561
rect 52154 542325 58918 542561
rect 59154 542325 65918 542561
rect 66154 542325 72918 542561
rect 73154 542325 79918 542561
rect 80154 542325 86918 542561
rect 87154 542325 93918 542561
rect 94154 542325 100918 542561
rect 101154 542325 107918 542561
rect 108154 542325 114918 542561
rect 115154 542325 121918 542561
rect 122154 542325 128918 542561
rect 129154 542325 135918 542561
rect 136154 542325 142918 542561
rect 143154 542325 149918 542561
rect 150154 542325 156918 542561
rect 157154 542325 163918 542561
rect 164154 542325 170918 542561
rect 171154 542325 177918 542561
rect 178154 542325 184918 542561
rect 185154 542325 191918 542561
rect 192154 542325 198918 542561
rect 199154 542325 205918 542561
rect 206154 542325 212918 542561
rect 213154 542325 219918 542561
rect 220154 542325 226918 542561
rect 227154 542325 233918 542561
rect 234154 542325 240918 542561
rect 241154 542325 247918 542561
rect 248154 542325 254918 542561
rect 255154 542325 261918 542561
rect 262154 542325 268918 542561
rect 269154 542325 275918 542561
rect 276154 542325 282918 542561
rect 283154 542325 289918 542561
rect 290154 542325 296918 542561
rect 297154 542325 303918 542561
rect 304154 542325 310918 542561
rect 311154 542325 317918 542561
rect 318154 542325 324918 542561
rect 325154 542325 331918 542561
rect 332154 542325 338918 542561
rect 339154 542325 345918 542561
rect 346154 542325 352918 542561
rect 353154 542325 359918 542561
rect 360154 542325 366918 542561
rect 367154 542325 373918 542561
rect 374154 542325 380918 542561
rect 381154 542325 387918 542561
rect 388154 542325 394918 542561
rect 395154 542325 401918 542561
rect 402154 542325 408918 542561
rect 409154 542325 415918 542561
rect 416154 542325 422918 542561
rect 423154 542325 429918 542561
rect 430154 542325 436918 542561
rect 437154 542325 443918 542561
rect 444154 542325 450918 542561
rect 451154 542325 457918 542561
rect 458154 542325 464918 542561
rect 465154 542325 471918 542561
rect 472154 542325 478918 542561
rect 479154 542325 485918 542561
rect 486154 542325 492918 542561
rect 493154 542325 499918 542561
rect 500154 542325 506918 542561
rect 507154 542325 513918 542561
rect 514154 542325 520918 542561
rect 521154 542325 527918 542561
rect 528154 542325 534918 542561
rect 535154 542325 541918 542561
rect 542154 542325 548918 542561
rect 549154 542325 555918 542561
rect 556154 542325 562918 542561
rect 563154 542325 569918 542561
rect 570154 542325 576918 542561
rect 577154 542325 587570 542561
rect 587806 542325 587890 542561
rect 588126 542325 588210 542561
rect 588446 542325 588530 542561
rect 588766 542325 588874 542561
rect -4950 542283 588874 542325
rect -4950 541494 588874 541536
rect -4950 541258 -3090 541494
rect -2854 541258 -2770 541494
rect -2534 541258 -2450 541494
rect -2214 541258 -2130 541494
rect -1894 541258 1186 541494
rect 1422 541258 8186 541494
rect 8422 541258 15186 541494
rect 15422 541258 22186 541494
rect 22422 541258 29186 541494
rect 29422 541258 36186 541494
rect 36422 541258 43186 541494
rect 43422 541258 50186 541494
rect 50422 541258 57186 541494
rect 57422 541258 64186 541494
rect 64422 541258 71186 541494
rect 71422 541258 78186 541494
rect 78422 541258 85186 541494
rect 85422 541258 92186 541494
rect 92422 541258 99186 541494
rect 99422 541258 106186 541494
rect 106422 541258 113186 541494
rect 113422 541258 120186 541494
rect 120422 541258 127186 541494
rect 127422 541258 134186 541494
rect 134422 541258 141186 541494
rect 141422 541258 148186 541494
rect 148422 541258 155186 541494
rect 155422 541258 162186 541494
rect 162422 541258 169186 541494
rect 169422 541258 176186 541494
rect 176422 541258 183186 541494
rect 183422 541258 190186 541494
rect 190422 541258 197186 541494
rect 197422 541258 204186 541494
rect 204422 541258 211186 541494
rect 211422 541258 218186 541494
rect 218422 541258 225186 541494
rect 225422 541258 232186 541494
rect 232422 541258 239186 541494
rect 239422 541258 246186 541494
rect 246422 541258 253186 541494
rect 253422 541258 260186 541494
rect 260422 541258 267186 541494
rect 267422 541258 274186 541494
rect 274422 541258 281186 541494
rect 281422 541258 288186 541494
rect 288422 541258 295186 541494
rect 295422 541258 302186 541494
rect 302422 541258 309186 541494
rect 309422 541258 316186 541494
rect 316422 541258 323186 541494
rect 323422 541258 330186 541494
rect 330422 541258 337186 541494
rect 337422 541258 344186 541494
rect 344422 541258 351186 541494
rect 351422 541258 358186 541494
rect 358422 541258 365186 541494
rect 365422 541258 372186 541494
rect 372422 541258 379186 541494
rect 379422 541258 386186 541494
rect 386422 541258 393186 541494
rect 393422 541258 400186 541494
rect 400422 541258 407186 541494
rect 407422 541258 414186 541494
rect 414422 541258 421186 541494
rect 421422 541258 428186 541494
rect 428422 541258 435186 541494
rect 435422 541258 442186 541494
rect 442422 541258 449186 541494
rect 449422 541258 456186 541494
rect 456422 541258 463186 541494
rect 463422 541258 470186 541494
rect 470422 541258 477186 541494
rect 477422 541258 484186 541494
rect 484422 541258 491186 541494
rect 491422 541258 498186 541494
rect 498422 541258 505186 541494
rect 505422 541258 512186 541494
rect 512422 541258 519186 541494
rect 519422 541258 526186 541494
rect 526422 541258 533186 541494
rect 533422 541258 540186 541494
rect 540422 541258 547186 541494
rect 547422 541258 554186 541494
rect 554422 541258 561186 541494
rect 561422 541258 568186 541494
rect 568422 541258 575186 541494
rect 575422 541258 582186 541494
rect 582422 541258 585818 541494
rect 586054 541258 586138 541494
rect 586374 541258 586458 541494
rect 586694 541258 586778 541494
rect 587014 541258 588874 541494
rect -4950 541216 588874 541258
rect -4950 535561 588874 535603
rect -4950 535325 -4842 535561
rect -4606 535325 -4522 535561
rect -4286 535325 -4202 535561
rect -3966 535325 -3882 535561
rect -3646 535325 2918 535561
rect 3154 535325 9918 535561
rect 10154 535325 16918 535561
rect 17154 535325 23918 535561
rect 24154 535325 30918 535561
rect 31154 535325 37918 535561
rect 38154 535325 44918 535561
rect 45154 535325 51918 535561
rect 52154 535325 58918 535561
rect 59154 535325 65918 535561
rect 66154 535325 72918 535561
rect 73154 535325 79918 535561
rect 80154 535325 86918 535561
rect 87154 535325 93918 535561
rect 94154 535325 100918 535561
rect 101154 535325 107918 535561
rect 108154 535325 114918 535561
rect 115154 535325 121918 535561
rect 122154 535325 128918 535561
rect 129154 535325 135918 535561
rect 136154 535325 142918 535561
rect 143154 535325 149918 535561
rect 150154 535325 156918 535561
rect 157154 535325 163918 535561
rect 164154 535325 170918 535561
rect 171154 535325 177918 535561
rect 178154 535325 184918 535561
rect 185154 535325 191918 535561
rect 192154 535325 198918 535561
rect 199154 535325 205918 535561
rect 206154 535325 212918 535561
rect 213154 535325 219918 535561
rect 220154 535325 226918 535561
rect 227154 535325 233918 535561
rect 234154 535325 240918 535561
rect 241154 535325 247918 535561
rect 248154 535325 254918 535561
rect 255154 535325 261918 535561
rect 262154 535325 268918 535561
rect 269154 535325 275918 535561
rect 276154 535325 282918 535561
rect 283154 535325 289918 535561
rect 290154 535325 296918 535561
rect 297154 535325 303918 535561
rect 304154 535325 310918 535561
rect 311154 535325 317918 535561
rect 318154 535325 324918 535561
rect 325154 535325 331918 535561
rect 332154 535325 338918 535561
rect 339154 535325 345918 535561
rect 346154 535325 352918 535561
rect 353154 535325 359918 535561
rect 360154 535325 366918 535561
rect 367154 535325 373918 535561
rect 374154 535325 380918 535561
rect 381154 535325 387918 535561
rect 388154 535325 394918 535561
rect 395154 535325 401918 535561
rect 402154 535325 408918 535561
rect 409154 535325 415918 535561
rect 416154 535325 422918 535561
rect 423154 535325 429918 535561
rect 430154 535325 436918 535561
rect 437154 535325 443918 535561
rect 444154 535325 450918 535561
rect 451154 535325 457918 535561
rect 458154 535325 464918 535561
rect 465154 535325 471918 535561
rect 472154 535325 478918 535561
rect 479154 535325 485918 535561
rect 486154 535325 492918 535561
rect 493154 535325 499918 535561
rect 500154 535325 506918 535561
rect 507154 535325 513918 535561
rect 514154 535325 520918 535561
rect 521154 535325 527918 535561
rect 528154 535325 534918 535561
rect 535154 535325 541918 535561
rect 542154 535325 548918 535561
rect 549154 535325 555918 535561
rect 556154 535325 562918 535561
rect 563154 535325 569918 535561
rect 570154 535325 576918 535561
rect 577154 535325 587570 535561
rect 587806 535325 587890 535561
rect 588126 535325 588210 535561
rect 588446 535325 588530 535561
rect 588766 535325 588874 535561
rect -4950 535283 588874 535325
rect -4950 534494 588874 534536
rect -4950 534258 -3090 534494
rect -2854 534258 -2770 534494
rect -2534 534258 -2450 534494
rect -2214 534258 -2130 534494
rect -1894 534258 1186 534494
rect 1422 534258 8186 534494
rect 8422 534258 15186 534494
rect 15422 534258 22186 534494
rect 22422 534258 29186 534494
rect 29422 534258 36186 534494
rect 36422 534258 43186 534494
rect 43422 534258 50186 534494
rect 50422 534258 57186 534494
rect 57422 534258 64186 534494
rect 64422 534258 71186 534494
rect 71422 534258 78186 534494
rect 78422 534258 85186 534494
rect 85422 534258 92186 534494
rect 92422 534258 99186 534494
rect 99422 534258 106186 534494
rect 106422 534258 113186 534494
rect 113422 534258 120186 534494
rect 120422 534258 127186 534494
rect 127422 534258 134186 534494
rect 134422 534258 141186 534494
rect 141422 534258 148186 534494
rect 148422 534258 155186 534494
rect 155422 534258 162186 534494
rect 162422 534258 169186 534494
rect 169422 534258 176186 534494
rect 176422 534258 183186 534494
rect 183422 534258 190186 534494
rect 190422 534258 197186 534494
rect 197422 534258 204186 534494
rect 204422 534258 211186 534494
rect 211422 534258 218186 534494
rect 218422 534258 225186 534494
rect 225422 534258 232186 534494
rect 232422 534258 239186 534494
rect 239422 534258 246186 534494
rect 246422 534258 253186 534494
rect 253422 534258 260186 534494
rect 260422 534258 267186 534494
rect 267422 534258 274186 534494
rect 274422 534258 281186 534494
rect 281422 534258 288186 534494
rect 288422 534258 295186 534494
rect 295422 534258 302186 534494
rect 302422 534258 309186 534494
rect 309422 534258 316186 534494
rect 316422 534258 323186 534494
rect 323422 534258 330186 534494
rect 330422 534258 337186 534494
rect 337422 534258 344186 534494
rect 344422 534258 351186 534494
rect 351422 534258 358186 534494
rect 358422 534258 365186 534494
rect 365422 534258 372186 534494
rect 372422 534258 379186 534494
rect 379422 534258 386186 534494
rect 386422 534258 393186 534494
rect 393422 534258 400186 534494
rect 400422 534258 407186 534494
rect 407422 534258 414186 534494
rect 414422 534258 421186 534494
rect 421422 534258 428186 534494
rect 428422 534258 435186 534494
rect 435422 534258 442186 534494
rect 442422 534258 449186 534494
rect 449422 534258 456186 534494
rect 456422 534258 463186 534494
rect 463422 534258 470186 534494
rect 470422 534258 477186 534494
rect 477422 534258 484186 534494
rect 484422 534258 491186 534494
rect 491422 534258 498186 534494
rect 498422 534258 505186 534494
rect 505422 534258 512186 534494
rect 512422 534258 519186 534494
rect 519422 534258 526186 534494
rect 526422 534258 533186 534494
rect 533422 534258 540186 534494
rect 540422 534258 547186 534494
rect 547422 534258 554186 534494
rect 554422 534258 561186 534494
rect 561422 534258 568186 534494
rect 568422 534258 575186 534494
rect 575422 534258 582186 534494
rect 582422 534258 585818 534494
rect 586054 534258 586138 534494
rect 586374 534258 586458 534494
rect 586694 534258 586778 534494
rect 587014 534258 588874 534494
rect -4950 534216 588874 534258
rect -4950 528561 588874 528603
rect -4950 528325 -4842 528561
rect -4606 528325 -4522 528561
rect -4286 528325 -4202 528561
rect -3966 528325 -3882 528561
rect -3646 528325 2918 528561
rect 3154 528325 9918 528561
rect 10154 528325 16918 528561
rect 17154 528325 23918 528561
rect 24154 528325 30918 528561
rect 31154 528325 37918 528561
rect 38154 528325 44918 528561
rect 45154 528325 51918 528561
rect 52154 528325 58918 528561
rect 59154 528325 65918 528561
rect 66154 528325 72918 528561
rect 73154 528325 79918 528561
rect 80154 528325 86918 528561
rect 87154 528325 93918 528561
rect 94154 528325 100918 528561
rect 101154 528325 107918 528561
rect 108154 528325 114918 528561
rect 115154 528325 121918 528561
rect 122154 528325 128918 528561
rect 129154 528325 135918 528561
rect 136154 528325 142918 528561
rect 143154 528325 149918 528561
rect 150154 528325 156918 528561
rect 157154 528325 163918 528561
rect 164154 528325 170918 528561
rect 171154 528325 177918 528561
rect 178154 528325 184918 528561
rect 185154 528325 191918 528561
rect 192154 528325 198918 528561
rect 199154 528325 205918 528561
rect 206154 528325 212918 528561
rect 213154 528325 219918 528561
rect 220154 528325 226918 528561
rect 227154 528325 233918 528561
rect 234154 528325 240918 528561
rect 241154 528325 247918 528561
rect 248154 528325 254918 528561
rect 255154 528325 261918 528561
rect 262154 528325 268918 528561
rect 269154 528325 275918 528561
rect 276154 528325 282918 528561
rect 283154 528325 289918 528561
rect 290154 528325 296918 528561
rect 297154 528325 303918 528561
rect 304154 528325 310918 528561
rect 311154 528325 317918 528561
rect 318154 528325 324918 528561
rect 325154 528325 331918 528561
rect 332154 528325 338918 528561
rect 339154 528325 345918 528561
rect 346154 528325 352918 528561
rect 353154 528325 359918 528561
rect 360154 528325 366918 528561
rect 367154 528325 373918 528561
rect 374154 528325 380918 528561
rect 381154 528325 387918 528561
rect 388154 528325 394918 528561
rect 395154 528325 401918 528561
rect 402154 528325 408918 528561
rect 409154 528325 415918 528561
rect 416154 528325 422918 528561
rect 423154 528325 429918 528561
rect 430154 528325 436918 528561
rect 437154 528325 443918 528561
rect 444154 528325 450918 528561
rect 451154 528325 457918 528561
rect 458154 528325 464918 528561
rect 465154 528325 471918 528561
rect 472154 528325 478918 528561
rect 479154 528325 485918 528561
rect 486154 528325 492918 528561
rect 493154 528325 499918 528561
rect 500154 528325 506918 528561
rect 507154 528325 513918 528561
rect 514154 528325 520918 528561
rect 521154 528325 527918 528561
rect 528154 528325 534918 528561
rect 535154 528325 541918 528561
rect 542154 528325 548918 528561
rect 549154 528325 555918 528561
rect 556154 528325 562918 528561
rect 563154 528325 569918 528561
rect 570154 528325 576918 528561
rect 577154 528325 587570 528561
rect 587806 528325 587890 528561
rect 588126 528325 588210 528561
rect 588446 528325 588530 528561
rect 588766 528325 588874 528561
rect -4950 528283 588874 528325
rect -4950 527494 588874 527536
rect -4950 527258 -3090 527494
rect -2854 527258 -2770 527494
rect -2534 527258 -2450 527494
rect -2214 527258 -2130 527494
rect -1894 527258 1186 527494
rect 1422 527258 8186 527494
rect 8422 527258 15186 527494
rect 15422 527258 22186 527494
rect 22422 527258 29186 527494
rect 29422 527258 36186 527494
rect 36422 527258 43186 527494
rect 43422 527258 50186 527494
rect 50422 527258 57186 527494
rect 57422 527258 64186 527494
rect 64422 527258 71186 527494
rect 71422 527258 78186 527494
rect 78422 527258 85186 527494
rect 85422 527258 92186 527494
rect 92422 527258 99186 527494
rect 99422 527258 106186 527494
rect 106422 527258 113186 527494
rect 113422 527258 120186 527494
rect 120422 527258 127186 527494
rect 127422 527258 134186 527494
rect 134422 527258 141186 527494
rect 141422 527258 148186 527494
rect 148422 527258 155186 527494
rect 155422 527258 162186 527494
rect 162422 527258 169186 527494
rect 169422 527258 176186 527494
rect 176422 527258 183186 527494
rect 183422 527258 190186 527494
rect 190422 527258 197186 527494
rect 197422 527258 204186 527494
rect 204422 527258 211186 527494
rect 211422 527258 218186 527494
rect 218422 527258 225186 527494
rect 225422 527258 232186 527494
rect 232422 527258 239186 527494
rect 239422 527258 246186 527494
rect 246422 527258 253186 527494
rect 253422 527258 260186 527494
rect 260422 527258 267186 527494
rect 267422 527258 274186 527494
rect 274422 527258 281186 527494
rect 281422 527258 288186 527494
rect 288422 527258 295186 527494
rect 295422 527258 302186 527494
rect 302422 527258 309186 527494
rect 309422 527258 316186 527494
rect 316422 527258 323186 527494
rect 323422 527258 330186 527494
rect 330422 527258 337186 527494
rect 337422 527258 344186 527494
rect 344422 527258 351186 527494
rect 351422 527258 358186 527494
rect 358422 527258 365186 527494
rect 365422 527258 372186 527494
rect 372422 527258 379186 527494
rect 379422 527258 386186 527494
rect 386422 527258 393186 527494
rect 393422 527258 400186 527494
rect 400422 527258 407186 527494
rect 407422 527258 414186 527494
rect 414422 527258 421186 527494
rect 421422 527258 428186 527494
rect 428422 527258 435186 527494
rect 435422 527258 442186 527494
rect 442422 527258 449186 527494
rect 449422 527258 456186 527494
rect 456422 527258 463186 527494
rect 463422 527258 470186 527494
rect 470422 527258 477186 527494
rect 477422 527258 484186 527494
rect 484422 527258 491186 527494
rect 491422 527258 498186 527494
rect 498422 527258 505186 527494
rect 505422 527258 512186 527494
rect 512422 527258 519186 527494
rect 519422 527258 526186 527494
rect 526422 527258 533186 527494
rect 533422 527258 540186 527494
rect 540422 527258 547186 527494
rect 547422 527258 554186 527494
rect 554422 527258 561186 527494
rect 561422 527258 568186 527494
rect 568422 527258 575186 527494
rect 575422 527258 582186 527494
rect 582422 527258 585818 527494
rect 586054 527258 586138 527494
rect 586374 527258 586458 527494
rect 586694 527258 586778 527494
rect 587014 527258 588874 527494
rect -4950 527216 588874 527258
rect -4950 521561 588874 521603
rect -4950 521325 -4842 521561
rect -4606 521325 -4522 521561
rect -4286 521325 -4202 521561
rect -3966 521325 -3882 521561
rect -3646 521325 2918 521561
rect 3154 521325 9918 521561
rect 10154 521325 16918 521561
rect 17154 521325 23918 521561
rect 24154 521325 30918 521561
rect 31154 521325 37918 521561
rect 38154 521325 44918 521561
rect 45154 521325 51918 521561
rect 52154 521325 58918 521561
rect 59154 521325 65918 521561
rect 66154 521325 72918 521561
rect 73154 521325 79918 521561
rect 80154 521325 86918 521561
rect 87154 521325 93918 521561
rect 94154 521325 100918 521561
rect 101154 521325 107918 521561
rect 108154 521325 114918 521561
rect 115154 521325 121918 521561
rect 122154 521325 128918 521561
rect 129154 521325 135918 521561
rect 136154 521325 142918 521561
rect 143154 521325 149918 521561
rect 150154 521325 156918 521561
rect 157154 521325 163918 521561
rect 164154 521325 170918 521561
rect 171154 521325 177918 521561
rect 178154 521325 184918 521561
rect 185154 521325 191918 521561
rect 192154 521325 198918 521561
rect 199154 521325 205918 521561
rect 206154 521325 212918 521561
rect 213154 521325 219918 521561
rect 220154 521325 226918 521561
rect 227154 521325 233918 521561
rect 234154 521325 240918 521561
rect 241154 521325 247918 521561
rect 248154 521325 254918 521561
rect 255154 521325 261918 521561
rect 262154 521325 268918 521561
rect 269154 521325 275918 521561
rect 276154 521325 282918 521561
rect 283154 521325 289918 521561
rect 290154 521325 296918 521561
rect 297154 521325 303918 521561
rect 304154 521325 310918 521561
rect 311154 521325 317918 521561
rect 318154 521325 324918 521561
rect 325154 521325 331918 521561
rect 332154 521325 338918 521561
rect 339154 521325 345918 521561
rect 346154 521325 352918 521561
rect 353154 521325 359918 521561
rect 360154 521325 366918 521561
rect 367154 521325 373918 521561
rect 374154 521325 380918 521561
rect 381154 521325 387918 521561
rect 388154 521325 394918 521561
rect 395154 521325 401918 521561
rect 402154 521325 408918 521561
rect 409154 521325 415918 521561
rect 416154 521325 422918 521561
rect 423154 521325 429918 521561
rect 430154 521325 436918 521561
rect 437154 521325 443918 521561
rect 444154 521325 450918 521561
rect 451154 521325 457918 521561
rect 458154 521325 464918 521561
rect 465154 521325 471918 521561
rect 472154 521325 478918 521561
rect 479154 521325 485918 521561
rect 486154 521325 492918 521561
rect 493154 521325 499918 521561
rect 500154 521325 506918 521561
rect 507154 521325 513918 521561
rect 514154 521325 520918 521561
rect 521154 521325 527918 521561
rect 528154 521325 534918 521561
rect 535154 521325 541918 521561
rect 542154 521325 548918 521561
rect 549154 521325 555918 521561
rect 556154 521325 562918 521561
rect 563154 521325 569918 521561
rect 570154 521325 576918 521561
rect 577154 521325 587570 521561
rect 587806 521325 587890 521561
rect 588126 521325 588210 521561
rect 588446 521325 588530 521561
rect 588766 521325 588874 521561
rect -4950 521283 588874 521325
rect -4950 520494 588874 520536
rect -4950 520258 -3090 520494
rect -2854 520258 -2770 520494
rect -2534 520258 -2450 520494
rect -2214 520258 -2130 520494
rect -1894 520258 1186 520494
rect 1422 520258 8186 520494
rect 8422 520258 15186 520494
rect 15422 520258 22186 520494
rect 22422 520258 29186 520494
rect 29422 520258 36186 520494
rect 36422 520258 43186 520494
rect 43422 520258 50186 520494
rect 50422 520258 57186 520494
rect 57422 520258 64186 520494
rect 64422 520258 71186 520494
rect 71422 520258 78186 520494
rect 78422 520258 85186 520494
rect 85422 520258 92186 520494
rect 92422 520258 99186 520494
rect 99422 520258 106186 520494
rect 106422 520258 113186 520494
rect 113422 520258 120186 520494
rect 120422 520258 127186 520494
rect 127422 520258 134186 520494
rect 134422 520258 141186 520494
rect 141422 520258 148186 520494
rect 148422 520258 155186 520494
rect 155422 520258 162186 520494
rect 162422 520258 169186 520494
rect 169422 520258 176186 520494
rect 176422 520258 183186 520494
rect 183422 520258 190186 520494
rect 190422 520258 197186 520494
rect 197422 520258 204186 520494
rect 204422 520258 211186 520494
rect 211422 520258 218186 520494
rect 218422 520258 225186 520494
rect 225422 520258 232186 520494
rect 232422 520258 239186 520494
rect 239422 520258 246186 520494
rect 246422 520258 253186 520494
rect 253422 520258 260186 520494
rect 260422 520258 267186 520494
rect 267422 520258 274186 520494
rect 274422 520258 281186 520494
rect 281422 520258 288186 520494
rect 288422 520258 295186 520494
rect 295422 520258 302186 520494
rect 302422 520258 309186 520494
rect 309422 520258 316186 520494
rect 316422 520258 323186 520494
rect 323422 520258 330186 520494
rect 330422 520258 337186 520494
rect 337422 520258 344186 520494
rect 344422 520258 351186 520494
rect 351422 520258 358186 520494
rect 358422 520258 365186 520494
rect 365422 520258 372186 520494
rect 372422 520258 379186 520494
rect 379422 520258 386186 520494
rect 386422 520258 393186 520494
rect 393422 520258 400186 520494
rect 400422 520258 407186 520494
rect 407422 520258 414186 520494
rect 414422 520258 421186 520494
rect 421422 520258 428186 520494
rect 428422 520258 435186 520494
rect 435422 520258 442186 520494
rect 442422 520258 449186 520494
rect 449422 520258 456186 520494
rect 456422 520258 463186 520494
rect 463422 520258 470186 520494
rect 470422 520258 477186 520494
rect 477422 520258 484186 520494
rect 484422 520258 491186 520494
rect 491422 520258 498186 520494
rect 498422 520258 505186 520494
rect 505422 520258 512186 520494
rect 512422 520258 519186 520494
rect 519422 520258 526186 520494
rect 526422 520258 533186 520494
rect 533422 520258 540186 520494
rect 540422 520258 547186 520494
rect 547422 520258 554186 520494
rect 554422 520258 561186 520494
rect 561422 520258 568186 520494
rect 568422 520258 575186 520494
rect 575422 520258 582186 520494
rect 582422 520258 585818 520494
rect 586054 520258 586138 520494
rect 586374 520258 586458 520494
rect 586694 520258 586778 520494
rect 587014 520258 588874 520494
rect -4950 520216 588874 520258
rect -4950 514561 588874 514603
rect -4950 514325 -4842 514561
rect -4606 514325 -4522 514561
rect -4286 514325 -4202 514561
rect -3966 514325 -3882 514561
rect -3646 514325 2918 514561
rect 3154 514325 9918 514561
rect 10154 514325 16918 514561
rect 17154 514325 23918 514561
rect 24154 514325 30918 514561
rect 31154 514325 37918 514561
rect 38154 514325 44918 514561
rect 45154 514325 51918 514561
rect 52154 514325 58918 514561
rect 59154 514325 65918 514561
rect 66154 514325 72918 514561
rect 73154 514325 79918 514561
rect 80154 514325 86918 514561
rect 87154 514325 93918 514561
rect 94154 514325 100918 514561
rect 101154 514325 107918 514561
rect 108154 514325 114918 514561
rect 115154 514325 121918 514561
rect 122154 514325 128918 514561
rect 129154 514325 135918 514561
rect 136154 514325 142918 514561
rect 143154 514325 149918 514561
rect 150154 514325 156918 514561
rect 157154 514325 163918 514561
rect 164154 514325 170918 514561
rect 171154 514325 177918 514561
rect 178154 514325 184918 514561
rect 185154 514325 191918 514561
rect 192154 514325 198918 514561
rect 199154 514325 205918 514561
rect 206154 514325 212918 514561
rect 213154 514325 219918 514561
rect 220154 514325 226918 514561
rect 227154 514325 233918 514561
rect 234154 514325 240918 514561
rect 241154 514325 247918 514561
rect 248154 514325 254918 514561
rect 255154 514325 261918 514561
rect 262154 514325 268918 514561
rect 269154 514325 275918 514561
rect 276154 514325 282918 514561
rect 283154 514325 289918 514561
rect 290154 514325 296918 514561
rect 297154 514325 303918 514561
rect 304154 514325 310918 514561
rect 311154 514325 317918 514561
rect 318154 514325 324918 514561
rect 325154 514325 331918 514561
rect 332154 514325 338918 514561
rect 339154 514325 345918 514561
rect 346154 514325 352918 514561
rect 353154 514325 359918 514561
rect 360154 514325 366918 514561
rect 367154 514325 373918 514561
rect 374154 514325 380918 514561
rect 381154 514325 387918 514561
rect 388154 514325 394918 514561
rect 395154 514325 401918 514561
rect 402154 514325 408918 514561
rect 409154 514325 415918 514561
rect 416154 514325 422918 514561
rect 423154 514325 429918 514561
rect 430154 514325 436918 514561
rect 437154 514325 443918 514561
rect 444154 514325 450918 514561
rect 451154 514325 457918 514561
rect 458154 514325 464918 514561
rect 465154 514325 471918 514561
rect 472154 514325 478918 514561
rect 479154 514325 485918 514561
rect 486154 514325 492918 514561
rect 493154 514325 499918 514561
rect 500154 514325 506918 514561
rect 507154 514325 513918 514561
rect 514154 514325 520918 514561
rect 521154 514325 527918 514561
rect 528154 514325 534918 514561
rect 535154 514325 541918 514561
rect 542154 514325 548918 514561
rect 549154 514325 555918 514561
rect 556154 514325 562918 514561
rect 563154 514325 569918 514561
rect 570154 514325 576918 514561
rect 577154 514325 587570 514561
rect 587806 514325 587890 514561
rect 588126 514325 588210 514561
rect 588446 514325 588530 514561
rect 588766 514325 588874 514561
rect -4950 514283 588874 514325
rect -4950 513494 588874 513536
rect -4950 513258 -3090 513494
rect -2854 513258 -2770 513494
rect -2534 513258 -2450 513494
rect -2214 513258 -2130 513494
rect -1894 513258 1186 513494
rect 1422 513258 8186 513494
rect 8422 513258 15186 513494
rect 15422 513258 22186 513494
rect 22422 513258 29186 513494
rect 29422 513258 36186 513494
rect 36422 513258 43186 513494
rect 43422 513258 50186 513494
rect 50422 513258 57186 513494
rect 57422 513258 64186 513494
rect 64422 513258 71186 513494
rect 71422 513258 78186 513494
rect 78422 513258 85186 513494
rect 85422 513258 92186 513494
rect 92422 513258 99186 513494
rect 99422 513258 106186 513494
rect 106422 513258 113186 513494
rect 113422 513258 120186 513494
rect 120422 513258 127186 513494
rect 127422 513258 134186 513494
rect 134422 513258 141186 513494
rect 141422 513258 148186 513494
rect 148422 513258 155186 513494
rect 155422 513258 162186 513494
rect 162422 513258 169186 513494
rect 169422 513258 176186 513494
rect 176422 513258 183186 513494
rect 183422 513258 190186 513494
rect 190422 513258 197186 513494
rect 197422 513258 204186 513494
rect 204422 513258 211186 513494
rect 211422 513258 218186 513494
rect 218422 513258 225186 513494
rect 225422 513258 232186 513494
rect 232422 513258 239186 513494
rect 239422 513258 246186 513494
rect 246422 513258 253186 513494
rect 253422 513258 260186 513494
rect 260422 513258 267186 513494
rect 267422 513258 274186 513494
rect 274422 513258 281186 513494
rect 281422 513258 288186 513494
rect 288422 513258 295186 513494
rect 295422 513258 302186 513494
rect 302422 513258 309186 513494
rect 309422 513258 316186 513494
rect 316422 513258 323186 513494
rect 323422 513258 330186 513494
rect 330422 513258 337186 513494
rect 337422 513258 344186 513494
rect 344422 513258 351186 513494
rect 351422 513258 358186 513494
rect 358422 513258 365186 513494
rect 365422 513258 372186 513494
rect 372422 513258 379186 513494
rect 379422 513258 386186 513494
rect 386422 513258 393186 513494
rect 393422 513258 400186 513494
rect 400422 513258 407186 513494
rect 407422 513258 414186 513494
rect 414422 513258 421186 513494
rect 421422 513258 428186 513494
rect 428422 513258 435186 513494
rect 435422 513258 442186 513494
rect 442422 513258 449186 513494
rect 449422 513258 456186 513494
rect 456422 513258 463186 513494
rect 463422 513258 470186 513494
rect 470422 513258 477186 513494
rect 477422 513258 484186 513494
rect 484422 513258 491186 513494
rect 491422 513258 498186 513494
rect 498422 513258 505186 513494
rect 505422 513258 512186 513494
rect 512422 513258 519186 513494
rect 519422 513258 526186 513494
rect 526422 513258 533186 513494
rect 533422 513258 540186 513494
rect 540422 513258 547186 513494
rect 547422 513258 554186 513494
rect 554422 513258 561186 513494
rect 561422 513258 568186 513494
rect 568422 513258 575186 513494
rect 575422 513258 582186 513494
rect 582422 513258 585818 513494
rect 586054 513258 586138 513494
rect 586374 513258 586458 513494
rect 586694 513258 586778 513494
rect 587014 513258 588874 513494
rect -4950 513216 588874 513258
rect -4950 507561 588874 507603
rect -4950 507325 -4842 507561
rect -4606 507325 -4522 507561
rect -4286 507325 -4202 507561
rect -3966 507325 -3882 507561
rect -3646 507325 2918 507561
rect 3154 507325 9918 507561
rect 10154 507325 16918 507561
rect 17154 507325 23918 507561
rect 24154 507325 30918 507561
rect 31154 507325 37918 507561
rect 38154 507325 44918 507561
rect 45154 507325 51918 507561
rect 52154 507325 58918 507561
rect 59154 507325 65918 507561
rect 66154 507325 72918 507561
rect 73154 507325 79918 507561
rect 80154 507325 86918 507561
rect 87154 507325 93918 507561
rect 94154 507325 100918 507561
rect 101154 507325 107918 507561
rect 108154 507325 114918 507561
rect 115154 507325 121918 507561
rect 122154 507325 128918 507561
rect 129154 507325 135918 507561
rect 136154 507325 142918 507561
rect 143154 507325 149918 507561
rect 150154 507325 156918 507561
rect 157154 507325 163918 507561
rect 164154 507325 170918 507561
rect 171154 507325 177918 507561
rect 178154 507325 184918 507561
rect 185154 507325 191918 507561
rect 192154 507325 198918 507561
rect 199154 507325 205918 507561
rect 206154 507325 212918 507561
rect 213154 507325 219918 507561
rect 220154 507325 226918 507561
rect 227154 507325 233918 507561
rect 234154 507325 240918 507561
rect 241154 507325 247918 507561
rect 248154 507325 254918 507561
rect 255154 507325 261918 507561
rect 262154 507325 268918 507561
rect 269154 507325 275918 507561
rect 276154 507325 282918 507561
rect 283154 507325 289918 507561
rect 290154 507325 296918 507561
rect 297154 507325 303918 507561
rect 304154 507325 310918 507561
rect 311154 507325 317918 507561
rect 318154 507325 324918 507561
rect 325154 507325 331918 507561
rect 332154 507325 338918 507561
rect 339154 507325 345918 507561
rect 346154 507325 352918 507561
rect 353154 507325 359918 507561
rect 360154 507325 366918 507561
rect 367154 507325 373918 507561
rect 374154 507325 380918 507561
rect 381154 507325 387918 507561
rect 388154 507325 394918 507561
rect 395154 507325 401918 507561
rect 402154 507325 408918 507561
rect 409154 507325 415918 507561
rect 416154 507325 422918 507561
rect 423154 507325 429918 507561
rect 430154 507325 436918 507561
rect 437154 507325 443918 507561
rect 444154 507325 450918 507561
rect 451154 507325 457918 507561
rect 458154 507325 464918 507561
rect 465154 507325 471918 507561
rect 472154 507325 478918 507561
rect 479154 507325 485918 507561
rect 486154 507325 492918 507561
rect 493154 507325 499918 507561
rect 500154 507325 506918 507561
rect 507154 507325 513918 507561
rect 514154 507325 520918 507561
rect 521154 507325 527918 507561
rect 528154 507325 534918 507561
rect 535154 507325 541918 507561
rect 542154 507325 548918 507561
rect 549154 507325 555918 507561
rect 556154 507325 562918 507561
rect 563154 507325 569918 507561
rect 570154 507325 576918 507561
rect 577154 507325 587570 507561
rect 587806 507325 587890 507561
rect 588126 507325 588210 507561
rect 588446 507325 588530 507561
rect 588766 507325 588874 507561
rect -4950 507283 588874 507325
rect -4950 506494 588874 506536
rect -4950 506258 -3090 506494
rect -2854 506258 -2770 506494
rect -2534 506258 -2450 506494
rect -2214 506258 -2130 506494
rect -1894 506258 1186 506494
rect 1422 506258 8186 506494
rect 8422 506258 15186 506494
rect 15422 506258 22186 506494
rect 22422 506258 29186 506494
rect 29422 506258 36186 506494
rect 36422 506258 43186 506494
rect 43422 506258 50186 506494
rect 50422 506258 57186 506494
rect 57422 506258 64186 506494
rect 64422 506258 71186 506494
rect 71422 506258 78186 506494
rect 78422 506258 85186 506494
rect 85422 506258 92186 506494
rect 92422 506258 99186 506494
rect 99422 506258 106186 506494
rect 106422 506258 113186 506494
rect 113422 506258 120186 506494
rect 120422 506258 127186 506494
rect 127422 506258 134186 506494
rect 134422 506258 141186 506494
rect 141422 506258 148186 506494
rect 148422 506258 155186 506494
rect 155422 506258 162186 506494
rect 162422 506258 169186 506494
rect 169422 506258 176186 506494
rect 176422 506258 183186 506494
rect 183422 506258 190186 506494
rect 190422 506258 197186 506494
rect 197422 506258 204186 506494
rect 204422 506258 211186 506494
rect 211422 506258 218186 506494
rect 218422 506258 225186 506494
rect 225422 506258 232186 506494
rect 232422 506258 239186 506494
rect 239422 506258 246186 506494
rect 246422 506258 253186 506494
rect 253422 506258 260186 506494
rect 260422 506258 267186 506494
rect 267422 506258 274186 506494
rect 274422 506258 281186 506494
rect 281422 506258 288186 506494
rect 288422 506258 295186 506494
rect 295422 506258 302186 506494
rect 302422 506258 309186 506494
rect 309422 506258 316186 506494
rect 316422 506258 323186 506494
rect 323422 506258 330186 506494
rect 330422 506258 337186 506494
rect 337422 506258 344186 506494
rect 344422 506258 351186 506494
rect 351422 506258 358186 506494
rect 358422 506258 365186 506494
rect 365422 506258 372186 506494
rect 372422 506258 379186 506494
rect 379422 506258 386186 506494
rect 386422 506258 393186 506494
rect 393422 506258 400186 506494
rect 400422 506258 407186 506494
rect 407422 506258 414186 506494
rect 414422 506258 421186 506494
rect 421422 506258 428186 506494
rect 428422 506258 435186 506494
rect 435422 506258 442186 506494
rect 442422 506258 449186 506494
rect 449422 506258 456186 506494
rect 456422 506258 463186 506494
rect 463422 506258 470186 506494
rect 470422 506258 477186 506494
rect 477422 506258 484186 506494
rect 484422 506258 491186 506494
rect 491422 506258 498186 506494
rect 498422 506258 505186 506494
rect 505422 506258 512186 506494
rect 512422 506258 519186 506494
rect 519422 506258 526186 506494
rect 526422 506258 533186 506494
rect 533422 506258 540186 506494
rect 540422 506258 547186 506494
rect 547422 506258 554186 506494
rect 554422 506258 561186 506494
rect 561422 506258 568186 506494
rect 568422 506258 575186 506494
rect 575422 506258 582186 506494
rect 582422 506258 585818 506494
rect 586054 506258 586138 506494
rect 586374 506258 586458 506494
rect 586694 506258 586778 506494
rect 587014 506258 588874 506494
rect -4950 506216 588874 506258
rect -4950 500561 588874 500603
rect -4950 500325 -4842 500561
rect -4606 500325 -4522 500561
rect -4286 500325 -4202 500561
rect -3966 500325 -3882 500561
rect -3646 500325 2918 500561
rect 3154 500325 9918 500561
rect 10154 500325 16918 500561
rect 17154 500325 23918 500561
rect 24154 500325 30918 500561
rect 31154 500325 37918 500561
rect 38154 500325 44918 500561
rect 45154 500325 51918 500561
rect 52154 500325 58918 500561
rect 59154 500325 65918 500561
rect 66154 500325 72918 500561
rect 73154 500325 79918 500561
rect 80154 500325 86918 500561
rect 87154 500325 93918 500561
rect 94154 500325 100918 500561
rect 101154 500325 107918 500561
rect 108154 500325 114918 500561
rect 115154 500325 121918 500561
rect 122154 500325 128918 500561
rect 129154 500325 135918 500561
rect 136154 500325 142918 500561
rect 143154 500325 149918 500561
rect 150154 500325 156918 500561
rect 157154 500325 163918 500561
rect 164154 500325 170918 500561
rect 171154 500325 177918 500561
rect 178154 500325 184918 500561
rect 185154 500325 191918 500561
rect 192154 500325 198918 500561
rect 199154 500325 205918 500561
rect 206154 500325 212918 500561
rect 213154 500325 219918 500561
rect 220154 500325 226918 500561
rect 227154 500325 233918 500561
rect 234154 500325 240918 500561
rect 241154 500325 247918 500561
rect 248154 500325 254918 500561
rect 255154 500325 261918 500561
rect 262154 500325 268918 500561
rect 269154 500325 275918 500561
rect 276154 500325 282918 500561
rect 283154 500325 289918 500561
rect 290154 500325 296918 500561
rect 297154 500325 303918 500561
rect 304154 500325 310918 500561
rect 311154 500325 317918 500561
rect 318154 500325 324918 500561
rect 325154 500325 331918 500561
rect 332154 500325 338918 500561
rect 339154 500325 345918 500561
rect 346154 500325 352918 500561
rect 353154 500325 359918 500561
rect 360154 500325 366918 500561
rect 367154 500325 373918 500561
rect 374154 500325 380918 500561
rect 381154 500325 387918 500561
rect 388154 500325 394918 500561
rect 395154 500325 401918 500561
rect 402154 500325 408918 500561
rect 409154 500325 415918 500561
rect 416154 500325 422918 500561
rect 423154 500325 429918 500561
rect 430154 500325 436918 500561
rect 437154 500325 443918 500561
rect 444154 500325 450918 500561
rect 451154 500325 457918 500561
rect 458154 500325 464918 500561
rect 465154 500325 471918 500561
rect 472154 500325 478918 500561
rect 479154 500325 485918 500561
rect 486154 500325 492918 500561
rect 493154 500325 499918 500561
rect 500154 500325 506918 500561
rect 507154 500325 513918 500561
rect 514154 500325 520918 500561
rect 521154 500325 527918 500561
rect 528154 500325 534918 500561
rect 535154 500325 541918 500561
rect 542154 500325 548918 500561
rect 549154 500325 555918 500561
rect 556154 500325 562918 500561
rect 563154 500325 569918 500561
rect 570154 500325 576918 500561
rect 577154 500325 587570 500561
rect 587806 500325 587890 500561
rect 588126 500325 588210 500561
rect 588446 500325 588530 500561
rect 588766 500325 588874 500561
rect -4950 500283 588874 500325
rect -4950 499494 588874 499536
rect -4950 499258 -3090 499494
rect -2854 499258 -2770 499494
rect -2534 499258 -2450 499494
rect -2214 499258 -2130 499494
rect -1894 499258 1186 499494
rect 1422 499258 8186 499494
rect 8422 499258 15186 499494
rect 15422 499258 22186 499494
rect 22422 499258 29186 499494
rect 29422 499258 36186 499494
rect 36422 499258 43186 499494
rect 43422 499258 50186 499494
rect 50422 499258 57186 499494
rect 57422 499258 64186 499494
rect 64422 499258 71186 499494
rect 71422 499258 78186 499494
rect 78422 499258 85186 499494
rect 85422 499258 92186 499494
rect 92422 499258 99186 499494
rect 99422 499258 106186 499494
rect 106422 499258 113186 499494
rect 113422 499258 120186 499494
rect 120422 499258 127186 499494
rect 127422 499258 134186 499494
rect 134422 499258 141186 499494
rect 141422 499258 148186 499494
rect 148422 499258 155186 499494
rect 155422 499258 162186 499494
rect 162422 499258 169186 499494
rect 169422 499258 176186 499494
rect 176422 499258 183186 499494
rect 183422 499258 190186 499494
rect 190422 499258 197186 499494
rect 197422 499258 204186 499494
rect 204422 499258 211186 499494
rect 211422 499258 218186 499494
rect 218422 499258 225186 499494
rect 225422 499258 232186 499494
rect 232422 499258 239186 499494
rect 239422 499258 246186 499494
rect 246422 499258 253186 499494
rect 253422 499258 260186 499494
rect 260422 499258 267186 499494
rect 267422 499258 274186 499494
rect 274422 499258 281186 499494
rect 281422 499258 288186 499494
rect 288422 499258 295186 499494
rect 295422 499258 302186 499494
rect 302422 499258 309186 499494
rect 309422 499258 316186 499494
rect 316422 499258 323186 499494
rect 323422 499258 330186 499494
rect 330422 499258 337186 499494
rect 337422 499258 344186 499494
rect 344422 499258 351186 499494
rect 351422 499258 358186 499494
rect 358422 499258 365186 499494
rect 365422 499258 372186 499494
rect 372422 499258 379186 499494
rect 379422 499258 386186 499494
rect 386422 499258 393186 499494
rect 393422 499258 400186 499494
rect 400422 499258 407186 499494
rect 407422 499258 414186 499494
rect 414422 499258 421186 499494
rect 421422 499258 428186 499494
rect 428422 499258 435186 499494
rect 435422 499258 442186 499494
rect 442422 499258 449186 499494
rect 449422 499258 456186 499494
rect 456422 499258 463186 499494
rect 463422 499258 470186 499494
rect 470422 499258 477186 499494
rect 477422 499258 484186 499494
rect 484422 499258 491186 499494
rect 491422 499258 498186 499494
rect 498422 499258 505186 499494
rect 505422 499258 512186 499494
rect 512422 499258 519186 499494
rect 519422 499258 526186 499494
rect 526422 499258 533186 499494
rect 533422 499258 540186 499494
rect 540422 499258 547186 499494
rect 547422 499258 554186 499494
rect 554422 499258 561186 499494
rect 561422 499258 568186 499494
rect 568422 499258 575186 499494
rect 575422 499258 582186 499494
rect 582422 499258 585818 499494
rect 586054 499258 586138 499494
rect 586374 499258 586458 499494
rect 586694 499258 586778 499494
rect 587014 499258 588874 499494
rect -4950 499216 588874 499258
rect -4950 493561 588874 493603
rect -4950 493325 -4842 493561
rect -4606 493325 -4522 493561
rect -4286 493325 -4202 493561
rect -3966 493325 -3882 493561
rect -3646 493325 2918 493561
rect 3154 493325 9918 493561
rect 10154 493325 16918 493561
rect 17154 493325 23918 493561
rect 24154 493325 30918 493561
rect 31154 493325 37918 493561
rect 38154 493325 44918 493561
rect 45154 493325 51918 493561
rect 52154 493325 58918 493561
rect 59154 493325 65918 493561
rect 66154 493325 72918 493561
rect 73154 493325 79918 493561
rect 80154 493325 86918 493561
rect 87154 493325 93918 493561
rect 94154 493325 100918 493561
rect 101154 493325 107918 493561
rect 108154 493325 114918 493561
rect 115154 493325 121918 493561
rect 122154 493325 128918 493561
rect 129154 493325 135918 493561
rect 136154 493325 142918 493561
rect 143154 493325 149918 493561
rect 150154 493325 156918 493561
rect 157154 493325 163918 493561
rect 164154 493325 170918 493561
rect 171154 493325 177918 493561
rect 178154 493325 184918 493561
rect 185154 493325 191918 493561
rect 192154 493325 198918 493561
rect 199154 493325 205918 493561
rect 206154 493325 212918 493561
rect 213154 493325 219918 493561
rect 220154 493325 226918 493561
rect 227154 493325 233918 493561
rect 234154 493325 240918 493561
rect 241154 493325 247918 493561
rect 248154 493325 254918 493561
rect 255154 493325 261918 493561
rect 262154 493325 268918 493561
rect 269154 493325 275918 493561
rect 276154 493325 282918 493561
rect 283154 493325 289918 493561
rect 290154 493325 296918 493561
rect 297154 493325 303918 493561
rect 304154 493325 310918 493561
rect 311154 493325 317918 493561
rect 318154 493325 324918 493561
rect 325154 493325 331918 493561
rect 332154 493325 338918 493561
rect 339154 493325 345918 493561
rect 346154 493325 352918 493561
rect 353154 493325 359918 493561
rect 360154 493325 366918 493561
rect 367154 493325 373918 493561
rect 374154 493325 380918 493561
rect 381154 493325 387918 493561
rect 388154 493325 394918 493561
rect 395154 493325 401918 493561
rect 402154 493325 408918 493561
rect 409154 493325 415918 493561
rect 416154 493325 422918 493561
rect 423154 493325 429918 493561
rect 430154 493325 436918 493561
rect 437154 493325 443918 493561
rect 444154 493325 450918 493561
rect 451154 493325 457918 493561
rect 458154 493325 464918 493561
rect 465154 493325 471918 493561
rect 472154 493325 478918 493561
rect 479154 493325 485918 493561
rect 486154 493325 492918 493561
rect 493154 493325 499918 493561
rect 500154 493325 506918 493561
rect 507154 493325 513918 493561
rect 514154 493325 520918 493561
rect 521154 493325 527918 493561
rect 528154 493325 534918 493561
rect 535154 493325 541918 493561
rect 542154 493325 548918 493561
rect 549154 493325 555918 493561
rect 556154 493325 562918 493561
rect 563154 493325 569918 493561
rect 570154 493325 576918 493561
rect 577154 493325 587570 493561
rect 587806 493325 587890 493561
rect 588126 493325 588210 493561
rect 588446 493325 588530 493561
rect 588766 493325 588874 493561
rect -4950 493283 588874 493325
rect -4950 492494 588874 492536
rect -4950 492258 -3090 492494
rect -2854 492258 -2770 492494
rect -2534 492258 -2450 492494
rect -2214 492258 -2130 492494
rect -1894 492258 1186 492494
rect 1422 492258 8186 492494
rect 8422 492258 15186 492494
rect 15422 492258 22186 492494
rect 22422 492258 29186 492494
rect 29422 492258 36186 492494
rect 36422 492258 43186 492494
rect 43422 492258 50186 492494
rect 50422 492258 57186 492494
rect 57422 492258 64186 492494
rect 64422 492258 71186 492494
rect 71422 492258 78186 492494
rect 78422 492258 85186 492494
rect 85422 492258 92186 492494
rect 92422 492258 99186 492494
rect 99422 492258 106186 492494
rect 106422 492258 113186 492494
rect 113422 492258 120186 492494
rect 120422 492258 127186 492494
rect 127422 492258 134186 492494
rect 134422 492258 141186 492494
rect 141422 492258 148186 492494
rect 148422 492258 155186 492494
rect 155422 492258 162186 492494
rect 162422 492258 169186 492494
rect 169422 492258 176186 492494
rect 176422 492258 183186 492494
rect 183422 492258 190186 492494
rect 190422 492258 197186 492494
rect 197422 492258 204186 492494
rect 204422 492258 211186 492494
rect 211422 492258 218186 492494
rect 218422 492258 225186 492494
rect 225422 492258 232186 492494
rect 232422 492258 239186 492494
rect 239422 492258 246186 492494
rect 246422 492258 253186 492494
rect 253422 492258 260186 492494
rect 260422 492258 267186 492494
rect 267422 492258 274186 492494
rect 274422 492258 281186 492494
rect 281422 492258 288186 492494
rect 288422 492258 295186 492494
rect 295422 492258 302186 492494
rect 302422 492258 309186 492494
rect 309422 492258 316186 492494
rect 316422 492258 323186 492494
rect 323422 492258 330186 492494
rect 330422 492258 337186 492494
rect 337422 492258 344186 492494
rect 344422 492258 351186 492494
rect 351422 492258 358186 492494
rect 358422 492258 365186 492494
rect 365422 492258 372186 492494
rect 372422 492258 379186 492494
rect 379422 492258 386186 492494
rect 386422 492258 393186 492494
rect 393422 492258 400186 492494
rect 400422 492258 407186 492494
rect 407422 492258 414186 492494
rect 414422 492258 421186 492494
rect 421422 492258 428186 492494
rect 428422 492258 435186 492494
rect 435422 492258 442186 492494
rect 442422 492258 449186 492494
rect 449422 492258 456186 492494
rect 456422 492258 463186 492494
rect 463422 492258 470186 492494
rect 470422 492258 477186 492494
rect 477422 492258 484186 492494
rect 484422 492258 491186 492494
rect 491422 492258 498186 492494
rect 498422 492258 505186 492494
rect 505422 492258 512186 492494
rect 512422 492258 519186 492494
rect 519422 492258 526186 492494
rect 526422 492258 533186 492494
rect 533422 492258 540186 492494
rect 540422 492258 547186 492494
rect 547422 492258 554186 492494
rect 554422 492258 561186 492494
rect 561422 492258 568186 492494
rect 568422 492258 575186 492494
rect 575422 492258 582186 492494
rect 582422 492258 585818 492494
rect 586054 492258 586138 492494
rect 586374 492258 586458 492494
rect 586694 492258 586778 492494
rect 587014 492258 588874 492494
rect -4950 492216 588874 492258
rect -4950 486561 588874 486603
rect -4950 486325 -4842 486561
rect -4606 486325 -4522 486561
rect -4286 486325 -4202 486561
rect -3966 486325 -3882 486561
rect -3646 486325 2918 486561
rect 3154 486325 9918 486561
rect 10154 486325 16918 486561
rect 17154 486325 23918 486561
rect 24154 486325 30918 486561
rect 31154 486325 37918 486561
rect 38154 486325 44918 486561
rect 45154 486325 51918 486561
rect 52154 486325 58918 486561
rect 59154 486325 65918 486561
rect 66154 486325 72918 486561
rect 73154 486325 79918 486561
rect 80154 486325 86918 486561
rect 87154 486325 93918 486561
rect 94154 486325 100918 486561
rect 101154 486325 107918 486561
rect 108154 486325 114918 486561
rect 115154 486325 121918 486561
rect 122154 486325 128918 486561
rect 129154 486325 135918 486561
rect 136154 486325 142918 486561
rect 143154 486325 149918 486561
rect 150154 486325 156918 486561
rect 157154 486325 163918 486561
rect 164154 486325 170918 486561
rect 171154 486325 177918 486561
rect 178154 486325 184918 486561
rect 185154 486325 191918 486561
rect 192154 486325 198918 486561
rect 199154 486325 205918 486561
rect 206154 486325 212918 486561
rect 213154 486325 219918 486561
rect 220154 486325 226918 486561
rect 227154 486325 233918 486561
rect 234154 486325 240918 486561
rect 241154 486325 247918 486561
rect 248154 486325 254918 486561
rect 255154 486325 261918 486561
rect 262154 486325 268918 486561
rect 269154 486325 275918 486561
rect 276154 486325 282918 486561
rect 283154 486325 289918 486561
rect 290154 486325 296918 486561
rect 297154 486325 303918 486561
rect 304154 486325 310918 486561
rect 311154 486325 317918 486561
rect 318154 486325 324918 486561
rect 325154 486325 331918 486561
rect 332154 486325 338918 486561
rect 339154 486325 345918 486561
rect 346154 486325 352918 486561
rect 353154 486325 359918 486561
rect 360154 486325 366918 486561
rect 367154 486325 373918 486561
rect 374154 486325 380918 486561
rect 381154 486325 387918 486561
rect 388154 486325 394918 486561
rect 395154 486325 401918 486561
rect 402154 486325 408918 486561
rect 409154 486325 415918 486561
rect 416154 486325 422918 486561
rect 423154 486325 429918 486561
rect 430154 486325 436918 486561
rect 437154 486325 443918 486561
rect 444154 486325 450918 486561
rect 451154 486325 457918 486561
rect 458154 486325 464918 486561
rect 465154 486325 471918 486561
rect 472154 486325 478918 486561
rect 479154 486325 485918 486561
rect 486154 486325 492918 486561
rect 493154 486325 499918 486561
rect 500154 486325 506918 486561
rect 507154 486325 513918 486561
rect 514154 486325 520918 486561
rect 521154 486325 527918 486561
rect 528154 486325 534918 486561
rect 535154 486325 541918 486561
rect 542154 486325 548918 486561
rect 549154 486325 555918 486561
rect 556154 486325 562918 486561
rect 563154 486325 569918 486561
rect 570154 486325 576918 486561
rect 577154 486325 587570 486561
rect 587806 486325 587890 486561
rect 588126 486325 588210 486561
rect 588446 486325 588530 486561
rect 588766 486325 588874 486561
rect -4950 486283 588874 486325
rect -4950 485494 588874 485536
rect -4950 485258 -3090 485494
rect -2854 485258 -2770 485494
rect -2534 485258 -2450 485494
rect -2214 485258 -2130 485494
rect -1894 485258 1186 485494
rect 1422 485258 8186 485494
rect 8422 485258 15186 485494
rect 15422 485258 22186 485494
rect 22422 485258 29186 485494
rect 29422 485258 36186 485494
rect 36422 485258 43186 485494
rect 43422 485258 50186 485494
rect 50422 485258 57186 485494
rect 57422 485258 64186 485494
rect 64422 485258 71186 485494
rect 71422 485258 78186 485494
rect 78422 485258 85186 485494
rect 85422 485258 92186 485494
rect 92422 485258 99186 485494
rect 99422 485258 106186 485494
rect 106422 485258 113186 485494
rect 113422 485258 120186 485494
rect 120422 485258 127186 485494
rect 127422 485258 134186 485494
rect 134422 485258 141186 485494
rect 141422 485258 148186 485494
rect 148422 485258 155186 485494
rect 155422 485258 162186 485494
rect 162422 485258 169186 485494
rect 169422 485258 176186 485494
rect 176422 485258 183186 485494
rect 183422 485258 190186 485494
rect 190422 485258 197186 485494
rect 197422 485258 204186 485494
rect 204422 485258 211186 485494
rect 211422 485258 218186 485494
rect 218422 485258 225186 485494
rect 225422 485258 232186 485494
rect 232422 485258 239186 485494
rect 239422 485258 246186 485494
rect 246422 485258 253186 485494
rect 253422 485258 260186 485494
rect 260422 485258 267186 485494
rect 267422 485258 274186 485494
rect 274422 485258 281186 485494
rect 281422 485258 288186 485494
rect 288422 485258 295186 485494
rect 295422 485258 302186 485494
rect 302422 485258 309186 485494
rect 309422 485258 316186 485494
rect 316422 485258 323186 485494
rect 323422 485258 330186 485494
rect 330422 485258 337186 485494
rect 337422 485258 344186 485494
rect 344422 485258 351186 485494
rect 351422 485258 358186 485494
rect 358422 485258 365186 485494
rect 365422 485258 372186 485494
rect 372422 485258 379186 485494
rect 379422 485258 386186 485494
rect 386422 485258 393186 485494
rect 393422 485258 400186 485494
rect 400422 485258 407186 485494
rect 407422 485258 414186 485494
rect 414422 485258 421186 485494
rect 421422 485258 428186 485494
rect 428422 485258 435186 485494
rect 435422 485258 442186 485494
rect 442422 485258 449186 485494
rect 449422 485258 456186 485494
rect 456422 485258 463186 485494
rect 463422 485258 470186 485494
rect 470422 485258 477186 485494
rect 477422 485258 484186 485494
rect 484422 485258 491186 485494
rect 491422 485258 498186 485494
rect 498422 485258 505186 485494
rect 505422 485258 512186 485494
rect 512422 485258 519186 485494
rect 519422 485258 526186 485494
rect 526422 485258 533186 485494
rect 533422 485258 540186 485494
rect 540422 485258 547186 485494
rect 547422 485258 554186 485494
rect 554422 485258 561186 485494
rect 561422 485258 568186 485494
rect 568422 485258 575186 485494
rect 575422 485258 582186 485494
rect 582422 485258 585818 485494
rect 586054 485258 586138 485494
rect 586374 485258 586458 485494
rect 586694 485258 586778 485494
rect 587014 485258 588874 485494
rect -4950 485216 588874 485258
rect -4950 479561 588874 479603
rect -4950 479325 -4842 479561
rect -4606 479325 -4522 479561
rect -4286 479325 -4202 479561
rect -3966 479325 -3882 479561
rect -3646 479325 2918 479561
rect 3154 479325 9918 479561
rect 10154 479325 16918 479561
rect 17154 479325 23918 479561
rect 24154 479325 30918 479561
rect 31154 479325 37918 479561
rect 38154 479325 44918 479561
rect 45154 479325 51918 479561
rect 52154 479325 58918 479561
rect 59154 479325 65918 479561
rect 66154 479325 72918 479561
rect 73154 479325 79918 479561
rect 80154 479325 86918 479561
rect 87154 479325 93918 479561
rect 94154 479325 100918 479561
rect 101154 479325 107918 479561
rect 108154 479325 114918 479561
rect 115154 479325 121918 479561
rect 122154 479325 128918 479561
rect 129154 479325 135918 479561
rect 136154 479325 142918 479561
rect 143154 479325 149918 479561
rect 150154 479325 156918 479561
rect 157154 479325 163918 479561
rect 164154 479325 170918 479561
rect 171154 479325 177918 479561
rect 178154 479325 184918 479561
rect 185154 479325 191918 479561
rect 192154 479325 198918 479561
rect 199154 479325 205918 479561
rect 206154 479325 212918 479561
rect 213154 479325 219918 479561
rect 220154 479325 226918 479561
rect 227154 479325 233918 479561
rect 234154 479325 240918 479561
rect 241154 479325 247918 479561
rect 248154 479325 254918 479561
rect 255154 479325 261918 479561
rect 262154 479325 268918 479561
rect 269154 479325 275918 479561
rect 276154 479325 282918 479561
rect 283154 479325 289918 479561
rect 290154 479325 296918 479561
rect 297154 479325 303918 479561
rect 304154 479325 310918 479561
rect 311154 479325 317918 479561
rect 318154 479325 324918 479561
rect 325154 479325 331918 479561
rect 332154 479325 338918 479561
rect 339154 479325 345918 479561
rect 346154 479325 352918 479561
rect 353154 479325 359918 479561
rect 360154 479325 366918 479561
rect 367154 479325 373918 479561
rect 374154 479325 380918 479561
rect 381154 479325 387918 479561
rect 388154 479325 394918 479561
rect 395154 479325 401918 479561
rect 402154 479325 408918 479561
rect 409154 479325 415918 479561
rect 416154 479325 422918 479561
rect 423154 479325 429918 479561
rect 430154 479325 436918 479561
rect 437154 479325 443918 479561
rect 444154 479325 450918 479561
rect 451154 479325 457918 479561
rect 458154 479325 464918 479561
rect 465154 479325 471918 479561
rect 472154 479325 478918 479561
rect 479154 479325 485918 479561
rect 486154 479325 492918 479561
rect 493154 479325 499918 479561
rect 500154 479325 506918 479561
rect 507154 479325 513918 479561
rect 514154 479325 520918 479561
rect 521154 479325 527918 479561
rect 528154 479325 534918 479561
rect 535154 479325 541918 479561
rect 542154 479325 548918 479561
rect 549154 479325 555918 479561
rect 556154 479325 562918 479561
rect 563154 479325 569918 479561
rect 570154 479325 576918 479561
rect 577154 479325 587570 479561
rect 587806 479325 587890 479561
rect 588126 479325 588210 479561
rect 588446 479325 588530 479561
rect 588766 479325 588874 479561
rect -4950 479283 588874 479325
rect -4950 478494 588874 478536
rect -4950 478258 -3090 478494
rect -2854 478258 -2770 478494
rect -2534 478258 -2450 478494
rect -2214 478258 -2130 478494
rect -1894 478258 1186 478494
rect 1422 478258 8186 478494
rect 8422 478258 15186 478494
rect 15422 478258 22186 478494
rect 22422 478258 29186 478494
rect 29422 478258 36186 478494
rect 36422 478258 43186 478494
rect 43422 478258 50186 478494
rect 50422 478258 57186 478494
rect 57422 478258 64186 478494
rect 64422 478258 71186 478494
rect 71422 478258 78186 478494
rect 78422 478258 85186 478494
rect 85422 478258 92186 478494
rect 92422 478258 99186 478494
rect 99422 478258 106186 478494
rect 106422 478258 113186 478494
rect 113422 478258 120186 478494
rect 120422 478258 127186 478494
rect 127422 478258 134186 478494
rect 134422 478258 141186 478494
rect 141422 478258 148186 478494
rect 148422 478258 155186 478494
rect 155422 478258 162186 478494
rect 162422 478258 169186 478494
rect 169422 478258 176186 478494
rect 176422 478258 183186 478494
rect 183422 478258 190186 478494
rect 190422 478258 197186 478494
rect 197422 478258 204186 478494
rect 204422 478258 211186 478494
rect 211422 478258 218186 478494
rect 218422 478258 225186 478494
rect 225422 478258 232186 478494
rect 232422 478258 239186 478494
rect 239422 478258 246186 478494
rect 246422 478258 253186 478494
rect 253422 478258 260186 478494
rect 260422 478258 267186 478494
rect 267422 478258 274186 478494
rect 274422 478258 281186 478494
rect 281422 478258 288186 478494
rect 288422 478258 295186 478494
rect 295422 478258 302186 478494
rect 302422 478258 309186 478494
rect 309422 478258 316186 478494
rect 316422 478258 323186 478494
rect 323422 478258 330186 478494
rect 330422 478258 337186 478494
rect 337422 478258 344186 478494
rect 344422 478258 351186 478494
rect 351422 478258 358186 478494
rect 358422 478258 365186 478494
rect 365422 478258 372186 478494
rect 372422 478258 379186 478494
rect 379422 478258 386186 478494
rect 386422 478258 393186 478494
rect 393422 478258 400186 478494
rect 400422 478258 407186 478494
rect 407422 478258 414186 478494
rect 414422 478258 421186 478494
rect 421422 478258 428186 478494
rect 428422 478258 435186 478494
rect 435422 478258 442186 478494
rect 442422 478258 449186 478494
rect 449422 478258 456186 478494
rect 456422 478258 463186 478494
rect 463422 478258 470186 478494
rect 470422 478258 477186 478494
rect 477422 478258 484186 478494
rect 484422 478258 491186 478494
rect 491422 478258 498186 478494
rect 498422 478258 505186 478494
rect 505422 478258 512186 478494
rect 512422 478258 519186 478494
rect 519422 478258 526186 478494
rect 526422 478258 533186 478494
rect 533422 478258 540186 478494
rect 540422 478258 547186 478494
rect 547422 478258 554186 478494
rect 554422 478258 561186 478494
rect 561422 478258 568186 478494
rect 568422 478258 575186 478494
rect 575422 478258 582186 478494
rect 582422 478258 585818 478494
rect 586054 478258 586138 478494
rect 586374 478258 586458 478494
rect 586694 478258 586778 478494
rect 587014 478258 588874 478494
rect -4950 478216 588874 478258
rect -4950 472561 588874 472603
rect -4950 472325 -4842 472561
rect -4606 472325 -4522 472561
rect -4286 472325 -4202 472561
rect -3966 472325 -3882 472561
rect -3646 472325 2918 472561
rect 3154 472325 9918 472561
rect 10154 472325 16918 472561
rect 17154 472325 23918 472561
rect 24154 472325 30918 472561
rect 31154 472325 37918 472561
rect 38154 472325 44918 472561
rect 45154 472325 51918 472561
rect 52154 472325 58918 472561
rect 59154 472325 65918 472561
rect 66154 472325 72918 472561
rect 73154 472325 79918 472561
rect 80154 472325 86918 472561
rect 87154 472325 93918 472561
rect 94154 472325 100918 472561
rect 101154 472325 107918 472561
rect 108154 472325 114918 472561
rect 115154 472325 121918 472561
rect 122154 472325 128918 472561
rect 129154 472325 135918 472561
rect 136154 472325 142918 472561
rect 143154 472325 149918 472561
rect 150154 472325 156918 472561
rect 157154 472325 163918 472561
rect 164154 472325 170918 472561
rect 171154 472325 177918 472561
rect 178154 472325 184918 472561
rect 185154 472325 191918 472561
rect 192154 472325 198918 472561
rect 199154 472325 205918 472561
rect 206154 472325 212918 472561
rect 213154 472325 219918 472561
rect 220154 472325 226918 472561
rect 227154 472325 233918 472561
rect 234154 472325 240918 472561
rect 241154 472325 247918 472561
rect 248154 472325 254918 472561
rect 255154 472325 261918 472561
rect 262154 472325 268918 472561
rect 269154 472325 275918 472561
rect 276154 472325 282918 472561
rect 283154 472325 289918 472561
rect 290154 472325 296918 472561
rect 297154 472325 303918 472561
rect 304154 472325 310918 472561
rect 311154 472325 317918 472561
rect 318154 472325 324918 472561
rect 325154 472325 331918 472561
rect 332154 472325 338918 472561
rect 339154 472325 345918 472561
rect 346154 472325 352918 472561
rect 353154 472325 359918 472561
rect 360154 472325 366918 472561
rect 367154 472325 373918 472561
rect 374154 472325 380918 472561
rect 381154 472325 387918 472561
rect 388154 472325 394918 472561
rect 395154 472325 401918 472561
rect 402154 472325 408918 472561
rect 409154 472325 415918 472561
rect 416154 472325 422918 472561
rect 423154 472325 429918 472561
rect 430154 472325 436918 472561
rect 437154 472325 443918 472561
rect 444154 472325 450918 472561
rect 451154 472325 457918 472561
rect 458154 472325 464918 472561
rect 465154 472325 471918 472561
rect 472154 472325 478918 472561
rect 479154 472325 485918 472561
rect 486154 472325 492918 472561
rect 493154 472325 499918 472561
rect 500154 472325 506918 472561
rect 507154 472325 513918 472561
rect 514154 472325 520918 472561
rect 521154 472325 527918 472561
rect 528154 472325 534918 472561
rect 535154 472325 541918 472561
rect 542154 472325 548918 472561
rect 549154 472325 555918 472561
rect 556154 472325 562918 472561
rect 563154 472325 569918 472561
rect 570154 472325 576918 472561
rect 577154 472325 587570 472561
rect 587806 472325 587890 472561
rect 588126 472325 588210 472561
rect 588446 472325 588530 472561
rect 588766 472325 588874 472561
rect -4950 472283 588874 472325
rect -4950 471494 588874 471536
rect -4950 471258 -3090 471494
rect -2854 471258 -2770 471494
rect -2534 471258 -2450 471494
rect -2214 471258 -2130 471494
rect -1894 471258 1186 471494
rect 1422 471258 8186 471494
rect 8422 471258 15186 471494
rect 15422 471258 22186 471494
rect 22422 471258 29186 471494
rect 29422 471258 36186 471494
rect 36422 471258 43186 471494
rect 43422 471258 50186 471494
rect 50422 471258 57186 471494
rect 57422 471258 64186 471494
rect 64422 471258 71186 471494
rect 71422 471258 78186 471494
rect 78422 471258 85186 471494
rect 85422 471258 92186 471494
rect 92422 471258 99186 471494
rect 99422 471258 106186 471494
rect 106422 471258 113186 471494
rect 113422 471258 120186 471494
rect 120422 471258 127186 471494
rect 127422 471258 134186 471494
rect 134422 471258 141186 471494
rect 141422 471258 148186 471494
rect 148422 471258 155186 471494
rect 155422 471258 162186 471494
rect 162422 471258 169186 471494
rect 169422 471258 176186 471494
rect 176422 471258 183186 471494
rect 183422 471258 190186 471494
rect 190422 471258 197186 471494
rect 197422 471258 204186 471494
rect 204422 471258 211186 471494
rect 211422 471258 218186 471494
rect 218422 471258 225186 471494
rect 225422 471258 232186 471494
rect 232422 471258 239186 471494
rect 239422 471258 246186 471494
rect 246422 471258 253186 471494
rect 253422 471258 260186 471494
rect 260422 471258 267186 471494
rect 267422 471258 274186 471494
rect 274422 471258 281186 471494
rect 281422 471258 288186 471494
rect 288422 471258 295186 471494
rect 295422 471258 302186 471494
rect 302422 471258 309186 471494
rect 309422 471258 316186 471494
rect 316422 471258 323186 471494
rect 323422 471258 330186 471494
rect 330422 471258 337186 471494
rect 337422 471258 344186 471494
rect 344422 471258 351186 471494
rect 351422 471258 358186 471494
rect 358422 471258 365186 471494
rect 365422 471258 372186 471494
rect 372422 471258 379186 471494
rect 379422 471258 386186 471494
rect 386422 471258 393186 471494
rect 393422 471258 400186 471494
rect 400422 471258 407186 471494
rect 407422 471258 414186 471494
rect 414422 471258 421186 471494
rect 421422 471258 428186 471494
rect 428422 471258 435186 471494
rect 435422 471258 442186 471494
rect 442422 471258 449186 471494
rect 449422 471258 456186 471494
rect 456422 471258 463186 471494
rect 463422 471258 470186 471494
rect 470422 471258 477186 471494
rect 477422 471258 484186 471494
rect 484422 471258 491186 471494
rect 491422 471258 498186 471494
rect 498422 471258 505186 471494
rect 505422 471258 512186 471494
rect 512422 471258 519186 471494
rect 519422 471258 526186 471494
rect 526422 471258 533186 471494
rect 533422 471258 540186 471494
rect 540422 471258 547186 471494
rect 547422 471258 554186 471494
rect 554422 471258 561186 471494
rect 561422 471258 568186 471494
rect 568422 471258 575186 471494
rect 575422 471258 582186 471494
rect 582422 471258 585818 471494
rect 586054 471258 586138 471494
rect 586374 471258 586458 471494
rect 586694 471258 586778 471494
rect 587014 471258 588874 471494
rect -4950 471216 588874 471258
rect -4950 465561 588874 465603
rect -4950 465325 -4842 465561
rect -4606 465325 -4522 465561
rect -4286 465325 -4202 465561
rect -3966 465325 -3882 465561
rect -3646 465325 2918 465561
rect 3154 465325 9918 465561
rect 10154 465325 16918 465561
rect 17154 465325 23918 465561
rect 24154 465325 30918 465561
rect 31154 465325 37918 465561
rect 38154 465325 44918 465561
rect 45154 465325 51918 465561
rect 52154 465325 58918 465561
rect 59154 465325 65918 465561
rect 66154 465325 72918 465561
rect 73154 465325 79918 465561
rect 80154 465325 86918 465561
rect 87154 465325 93918 465561
rect 94154 465325 100918 465561
rect 101154 465325 107918 465561
rect 108154 465325 114918 465561
rect 115154 465325 121918 465561
rect 122154 465325 128918 465561
rect 129154 465325 135918 465561
rect 136154 465325 142918 465561
rect 143154 465325 149918 465561
rect 150154 465325 156918 465561
rect 157154 465325 163918 465561
rect 164154 465325 170918 465561
rect 171154 465325 177918 465561
rect 178154 465325 184918 465561
rect 185154 465325 191918 465561
rect 192154 465325 198918 465561
rect 199154 465325 205918 465561
rect 206154 465325 212918 465561
rect 213154 465325 219918 465561
rect 220154 465325 226918 465561
rect 227154 465325 233918 465561
rect 234154 465325 240918 465561
rect 241154 465325 247918 465561
rect 248154 465325 254918 465561
rect 255154 465325 261918 465561
rect 262154 465325 268918 465561
rect 269154 465325 275918 465561
rect 276154 465325 282918 465561
rect 283154 465325 289918 465561
rect 290154 465325 296918 465561
rect 297154 465325 303918 465561
rect 304154 465325 310918 465561
rect 311154 465325 317918 465561
rect 318154 465325 324918 465561
rect 325154 465325 331918 465561
rect 332154 465325 338918 465561
rect 339154 465325 345918 465561
rect 346154 465325 352918 465561
rect 353154 465325 359918 465561
rect 360154 465325 366918 465561
rect 367154 465325 373918 465561
rect 374154 465325 380918 465561
rect 381154 465325 387918 465561
rect 388154 465325 394918 465561
rect 395154 465325 401918 465561
rect 402154 465325 408918 465561
rect 409154 465325 415918 465561
rect 416154 465325 422918 465561
rect 423154 465325 429918 465561
rect 430154 465325 436918 465561
rect 437154 465325 443918 465561
rect 444154 465325 450918 465561
rect 451154 465325 457918 465561
rect 458154 465325 464918 465561
rect 465154 465325 471918 465561
rect 472154 465325 478918 465561
rect 479154 465325 485918 465561
rect 486154 465325 492918 465561
rect 493154 465325 499918 465561
rect 500154 465325 506918 465561
rect 507154 465325 513918 465561
rect 514154 465325 520918 465561
rect 521154 465325 527918 465561
rect 528154 465325 534918 465561
rect 535154 465325 541918 465561
rect 542154 465325 548918 465561
rect 549154 465325 555918 465561
rect 556154 465325 562918 465561
rect 563154 465325 569918 465561
rect 570154 465325 576918 465561
rect 577154 465325 587570 465561
rect 587806 465325 587890 465561
rect 588126 465325 588210 465561
rect 588446 465325 588530 465561
rect 588766 465325 588874 465561
rect -4950 465283 588874 465325
rect -4950 464494 588874 464536
rect -4950 464258 -3090 464494
rect -2854 464258 -2770 464494
rect -2534 464258 -2450 464494
rect -2214 464258 -2130 464494
rect -1894 464258 1186 464494
rect 1422 464258 8186 464494
rect 8422 464258 15186 464494
rect 15422 464258 22186 464494
rect 22422 464258 29186 464494
rect 29422 464258 36186 464494
rect 36422 464258 43186 464494
rect 43422 464258 50186 464494
rect 50422 464258 57186 464494
rect 57422 464258 64186 464494
rect 64422 464258 71186 464494
rect 71422 464258 78186 464494
rect 78422 464258 85186 464494
rect 85422 464258 92186 464494
rect 92422 464258 99186 464494
rect 99422 464258 106186 464494
rect 106422 464258 113186 464494
rect 113422 464258 120186 464494
rect 120422 464258 127186 464494
rect 127422 464258 134186 464494
rect 134422 464258 141186 464494
rect 141422 464258 148186 464494
rect 148422 464258 155186 464494
rect 155422 464258 162186 464494
rect 162422 464258 169186 464494
rect 169422 464258 176186 464494
rect 176422 464258 183186 464494
rect 183422 464258 190186 464494
rect 190422 464258 197186 464494
rect 197422 464258 204186 464494
rect 204422 464258 211186 464494
rect 211422 464258 218186 464494
rect 218422 464258 225186 464494
rect 225422 464258 232186 464494
rect 232422 464258 239186 464494
rect 239422 464258 246186 464494
rect 246422 464258 253186 464494
rect 253422 464258 260186 464494
rect 260422 464258 267186 464494
rect 267422 464258 274186 464494
rect 274422 464258 281186 464494
rect 281422 464258 288186 464494
rect 288422 464258 295186 464494
rect 295422 464258 302186 464494
rect 302422 464258 309186 464494
rect 309422 464258 316186 464494
rect 316422 464258 323186 464494
rect 323422 464258 330186 464494
rect 330422 464258 337186 464494
rect 337422 464258 344186 464494
rect 344422 464258 351186 464494
rect 351422 464258 358186 464494
rect 358422 464258 365186 464494
rect 365422 464258 372186 464494
rect 372422 464258 379186 464494
rect 379422 464258 386186 464494
rect 386422 464258 393186 464494
rect 393422 464258 400186 464494
rect 400422 464258 407186 464494
rect 407422 464258 414186 464494
rect 414422 464258 421186 464494
rect 421422 464258 428186 464494
rect 428422 464258 435186 464494
rect 435422 464258 442186 464494
rect 442422 464258 449186 464494
rect 449422 464258 456186 464494
rect 456422 464258 463186 464494
rect 463422 464258 470186 464494
rect 470422 464258 477186 464494
rect 477422 464258 484186 464494
rect 484422 464258 491186 464494
rect 491422 464258 498186 464494
rect 498422 464258 505186 464494
rect 505422 464258 512186 464494
rect 512422 464258 519186 464494
rect 519422 464258 526186 464494
rect 526422 464258 533186 464494
rect 533422 464258 540186 464494
rect 540422 464258 547186 464494
rect 547422 464258 554186 464494
rect 554422 464258 561186 464494
rect 561422 464258 568186 464494
rect 568422 464258 575186 464494
rect 575422 464258 582186 464494
rect 582422 464258 585818 464494
rect 586054 464258 586138 464494
rect 586374 464258 586458 464494
rect 586694 464258 586778 464494
rect 587014 464258 588874 464494
rect -4950 464216 588874 464258
rect -4950 458561 588874 458603
rect -4950 458325 -4842 458561
rect -4606 458325 -4522 458561
rect -4286 458325 -4202 458561
rect -3966 458325 -3882 458561
rect -3646 458325 2918 458561
rect 3154 458325 9918 458561
rect 10154 458325 16918 458561
rect 17154 458325 23918 458561
rect 24154 458325 30918 458561
rect 31154 458325 37918 458561
rect 38154 458325 44918 458561
rect 45154 458325 51918 458561
rect 52154 458325 58918 458561
rect 59154 458325 65918 458561
rect 66154 458325 72918 458561
rect 73154 458325 79918 458561
rect 80154 458325 86918 458561
rect 87154 458325 93918 458561
rect 94154 458325 100918 458561
rect 101154 458325 107918 458561
rect 108154 458325 114918 458561
rect 115154 458325 121918 458561
rect 122154 458325 128918 458561
rect 129154 458325 135918 458561
rect 136154 458325 142918 458561
rect 143154 458325 149918 458561
rect 150154 458325 156918 458561
rect 157154 458325 163918 458561
rect 164154 458325 170918 458561
rect 171154 458325 177918 458561
rect 178154 458325 184918 458561
rect 185154 458325 191918 458561
rect 192154 458325 198918 458561
rect 199154 458325 205918 458561
rect 206154 458325 212918 458561
rect 213154 458325 219918 458561
rect 220154 458325 226918 458561
rect 227154 458325 233918 458561
rect 234154 458325 240918 458561
rect 241154 458325 247918 458561
rect 248154 458325 254918 458561
rect 255154 458325 261918 458561
rect 262154 458325 268918 458561
rect 269154 458325 275918 458561
rect 276154 458325 282918 458561
rect 283154 458325 289918 458561
rect 290154 458325 296918 458561
rect 297154 458325 303918 458561
rect 304154 458325 310918 458561
rect 311154 458325 317918 458561
rect 318154 458325 324918 458561
rect 325154 458325 331918 458561
rect 332154 458325 338918 458561
rect 339154 458325 345918 458561
rect 346154 458325 352918 458561
rect 353154 458325 359918 458561
rect 360154 458325 366918 458561
rect 367154 458325 373918 458561
rect 374154 458325 380918 458561
rect 381154 458325 387918 458561
rect 388154 458325 394918 458561
rect 395154 458325 401918 458561
rect 402154 458325 408918 458561
rect 409154 458325 415918 458561
rect 416154 458325 422918 458561
rect 423154 458325 429918 458561
rect 430154 458325 436918 458561
rect 437154 458325 443918 458561
rect 444154 458325 450918 458561
rect 451154 458325 457918 458561
rect 458154 458325 464918 458561
rect 465154 458325 471918 458561
rect 472154 458325 478918 458561
rect 479154 458325 485918 458561
rect 486154 458325 492918 458561
rect 493154 458325 499918 458561
rect 500154 458325 506918 458561
rect 507154 458325 513918 458561
rect 514154 458325 520918 458561
rect 521154 458325 527918 458561
rect 528154 458325 534918 458561
rect 535154 458325 541918 458561
rect 542154 458325 548918 458561
rect 549154 458325 555918 458561
rect 556154 458325 562918 458561
rect 563154 458325 569918 458561
rect 570154 458325 576918 458561
rect 577154 458325 587570 458561
rect 587806 458325 587890 458561
rect 588126 458325 588210 458561
rect 588446 458325 588530 458561
rect 588766 458325 588874 458561
rect -4950 458283 588874 458325
rect -4950 457494 588874 457536
rect -4950 457258 -3090 457494
rect -2854 457258 -2770 457494
rect -2534 457258 -2450 457494
rect -2214 457258 -2130 457494
rect -1894 457258 1186 457494
rect 1422 457258 8186 457494
rect 8422 457258 15186 457494
rect 15422 457258 22186 457494
rect 22422 457258 29186 457494
rect 29422 457258 36186 457494
rect 36422 457258 43186 457494
rect 43422 457258 50186 457494
rect 50422 457258 57186 457494
rect 57422 457258 64186 457494
rect 64422 457258 71186 457494
rect 71422 457258 78186 457494
rect 78422 457258 85186 457494
rect 85422 457258 92186 457494
rect 92422 457258 99186 457494
rect 99422 457258 106186 457494
rect 106422 457258 113186 457494
rect 113422 457258 120186 457494
rect 120422 457258 127186 457494
rect 127422 457258 134186 457494
rect 134422 457258 141186 457494
rect 141422 457258 148186 457494
rect 148422 457258 155186 457494
rect 155422 457258 162186 457494
rect 162422 457258 169186 457494
rect 169422 457258 176186 457494
rect 176422 457258 183186 457494
rect 183422 457258 190186 457494
rect 190422 457258 197186 457494
rect 197422 457258 204186 457494
rect 204422 457258 211186 457494
rect 211422 457258 218186 457494
rect 218422 457258 225186 457494
rect 225422 457258 232186 457494
rect 232422 457258 239186 457494
rect 239422 457258 246186 457494
rect 246422 457258 253186 457494
rect 253422 457258 260186 457494
rect 260422 457258 267186 457494
rect 267422 457258 274186 457494
rect 274422 457258 281186 457494
rect 281422 457258 288186 457494
rect 288422 457258 295186 457494
rect 295422 457258 302186 457494
rect 302422 457258 309186 457494
rect 309422 457258 316186 457494
rect 316422 457258 323186 457494
rect 323422 457258 330186 457494
rect 330422 457258 337186 457494
rect 337422 457258 344186 457494
rect 344422 457258 351186 457494
rect 351422 457258 358186 457494
rect 358422 457258 365186 457494
rect 365422 457258 372186 457494
rect 372422 457258 379186 457494
rect 379422 457258 386186 457494
rect 386422 457258 393186 457494
rect 393422 457258 400186 457494
rect 400422 457258 407186 457494
rect 407422 457258 414186 457494
rect 414422 457258 421186 457494
rect 421422 457258 428186 457494
rect 428422 457258 435186 457494
rect 435422 457258 442186 457494
rect 442422 457258 449186 457494
rect 449422 457258 456186 457494
rect 456422 457258 463186 457494
rect 463422 457258 470186 457494
rect 470422 457258 477186 457494
rect 477422 457258 484186 457494
rect 484422 457258 491186 457494
rect 491422 457258 498186 457494
rect 498422 457258 505186 457494
rect 505422 457258 512186 457494
rect 512422 457258 519186 457494
rect 519422 457258 526186 457494
rect 526422 457258 533186 457494
rect 533422 457258 540186 457494
rect 540422 457258 547186 457494
rect 547422 457258 554186 457494
rect 554422 457258 561186 457494
rect 561422 457258 568186 457494
rect 568422 457258 575186 457494
rect 575422 457258 582186 457494
rect 582422 457258 585818 457494
rect 586054 457258 586138 457494
rect 586374 457258 586458 457494
rect 586694 457258 586778 457494
rect 587014 457258 588874 457494
rect -4950 457216 588874 457258
rect -4950 451561 588874 451603
rect -4950 451325 -4842 451561
rect -4606 451325 -4522 451561
rect -4286 451325 -4202 451561
rect -3966 451325 -3882 451561
rect -3646 451325 2918 451561
rect 3154 451325 9918 451561
rect 10154 451325 16918 451561
rect 17154 451325 23918 451561
rect 24154 451325 30918 451561
rect 31154 451325 37918 451561
rect 38154 451325 44918 451561
rect 45154 451325 51918 451561
rect 52154 451325 58918 451561
rect 59154 451325 65918 451561
rect 66154 451325 72918 451561
rect 73154 451325 79918 451561
rect 80154 451325 86918 451561
rect 87154 451325 93918 451561
rect 94154 451325 100918 451561
rect 101154 451325 107918 451561
rect 108154 451325 114918 451561
rect 115154 451325 121918 451561
rect 122154 451325 128918 451561
rect 129154 451325 135918 451561
rect 136154 451325 142918 451561
rect 143154 451325 149918 451561
rect 150154 451325 156918 451561
rect 157154 451325 163918 451561
rect 164154 451325 170918 451561
rect 171154 451325 177918 451561
rect 178154 451325 184918 451561
rect 185154 451325 191918 451561
rect 192154 451325 198918 451561
rect 199154 451325 205918 451561
rect 206154 451325 212918 451561
rect 213154 451325 219918 451561
rect 220154 451325 226918 451561
rect 227154 451325 233918 451561
rect 234154 451325 240918 451561
rect 241154 451325 247918 451561
rect 248154 451325 254918 451561
rect 255154 451325 261918 451561
rect 262154 451325 268918 451561
rect 269154 451325 275918 451561
rect 276154 451325 282918 451561
rect 283154 451325 289918 451561
rect 290154 451325 296918 451561
rect 297154 451325 303918 451561
rect 304154 451325 310918 451561
rect 311154 451325 317918 451561
rect 318154 451325 324918 451561
rect 325154 451325 331918 451561
rect 332154 451325 338918 451561
rect 339154 451325 345918 451561
rect 346154 451325 352918 451561
rect 353154 451325 359918 451561
rect 360154 451325 366918 451561
rect 367154 451325 373918 451561
rect 374154 451325 380918 451561
rect 381154 451325 387918 451561
rect 388154 451325 394918 451561
rect 395154 451325 401918 451561
rect 402154 451325 408918 451561
rect 409154 451325 415918 451561
rect 416154 451325 422918 451561
rect 423154 451325 429918 451561
rect 430154 451325 436918 451561
rect 437154 451325 443918 451561
rect 444154 451325 450918 451561
rect 451154 451325 457918 451561
rect 458154 451325 464918 451561
rect 465154 451325 471918 451561
rect 472154 451325 478918 451561
rect 479154 451325 485918 451561
rect 486154 451325 492918 451561
rect 493154 451325 499918 451561
rect 500154 451325 506918 451561
rect 507154 451325 513918 451561
rect 514154 451325 520918 451561
rect 521154 451325 527918 451561
rect 528154 451325 534918 451561
rect 535154 451325 541918 451561
rect 542154 451325 548918 451561
rect 549154 451325 555918 451561
rect 556154 451325 562918 451561
rect 563154 451325 569918 451561
rect 570154 451325 576918 451561
rect 577154 451325 587570 451561
rect 587806 451325 587890 451561
rect 588126 451325 588210 451561
rect 588446 451325 588530 451561
rect 588766 451325 588874 451561
rect -4950 451283 588874 451325
rect -4950 450494 588874 450536
rect -4950 450258 -3090 450494
rect -2854 450258 -2770 450494
rect -2534 450258 -2450 450494
rect -2214 450258 -2130 450494
rect -1894 450258 1186 450494
rect 1422 450258 8186 450494
rect 8422 450258 15186 450494
rect 15422 450258 22186 450494
rect 22422 450258 29186 450494
rect 29422 450258 36186 450494
rect 36422 450258 43186 450494
rect 43422 450258 50186 450494
rect 50422 450258 57186 450494
rect 57422 450258 64186 450494
rect 64422 450258 71186 450494
rect 71422 450258 78186 450494
rect 78422 450258 85186 450494
rect 85422 450258 92186 450494
rect 92422 450258 99186 450494
rect 99422 450258 106186 450494
rect 106422 450258 113186 450494
rect 113422 450258 120186 450494
rect 120422 450258 127186 450494
rect 127422 450258 134186 450494
rect 134422 450258 141186 450494
rect 141422 450258 148186 450494
rect 148422 450258 155186 450494
rect 155422 450258 162186 450494
rect 162422 450258 169186 450494
rect 169422 450258 176186 450494
rect 176422 450258 183186 450494
rect 183422 450258 190186 450494
rect 190422 450258 197186 450494
rect 197422 450258 204186 450494
rect 204422 450258 211186 450494
rect 211422 450258 218186 450494
rect 218422 450258 225186 450494
rect 225422 450258 232186 450494
rect 232422 450258 239186 450494
rect 239422 450258 246186 450494
rect 246422 450258 253186 450494
rect 253422 450258 260186 450494
rect 260422 450258 267186 450494
rect 267422 450258 274186 450494
rect 274422 450258 281186 450494
rect 281422 450258 288186 450494
rect 288422 450258 295186 450494
rect 295422 450258 302186 450494
rect 302422 450258 309186 450494
rect 309422 450258 316186 450494
rect 316422 450258 323186 450494
rect 323422 450258 330186 450494
rect 330422 450258 337186 450494
rect 337422 450258 344186 450494
rect 344422 450258 351186 450494
rect 351422 450258 358186 450494
rect 358422 450258 365186 450494
rect 365422 450258 372186 450494
rect 372422 450258 379186 450494
rect 379422 450258 386186 450494
rect 386422 450258 393186 450494
rect 393422 450258 400186 450494
rect 400422 450258 407186 450494
rect 407422 450258 414186 450494
rect 414422 450258 421186 450494
rect 421422 450258 428186 450494
rect 428422 450258 435186 450494
rect 435422 450258 442186 450494
rect 442422 450258 449186 450494
rect 449422 450258 456186 450494
rect 456422 450258 463186 450494
rect 463422 450258 470186 450494
rect 470422 450258 477186 450494
rect 477422 450258 484186 450494
rect 484422 450258 491186 450494
rect 491422 450258 498186 450494
rect 498422 450258 505186 450494
rect 505422 450258 512186 450494
rect 512422 450258 519186 450494
rect 519422 450258 526186 450494
rect 526422 450258 533186 450494
rect 533422 450258 540186 450494
rect 540422 450258 547186 450494
rect 547422 450258 554186 450494
rect 554422 450258 561186 450494
rect 561422 450258 568186 450494
rect 568422 450258 575186 450494
rect 575422 450258 582186 450494
rect 582422 450258 585818 450494
rect 586054 450258 586138 450494
rect 586374 450258 586458 450494
rect 586694 450258 586778 450494
rect 587014 450258 588874 450494
rect -4950 450216 588874 450258
rect -4950 444561 588874 444603
rect -4950 444325 -4842 444561
rect -4606 444325 -4522 444561
rect -4286 444325 -4202 444561
rect -3966 444325 -3882 444561
rect -3646 444325 2918 444561
rect 3154 444325 9918 444561
rect 10154 444325 16918 444561
rect 17154 444325 23918 444561
rect 24154 444325 30918 444561
rect 31154 444325 37918 444561
rect 38154 444325 44918 444561
rect 45154 444325 51918 444561
rect 52154 444325 58918 444561
rect 59154 444325 65918 444561
rect 66154 444325 72918 444561
rect 73154 444325 79918 444561
rect 80154 444325 86918 444561
rect 87154 444325 93918 444561
rect 94154 444325 100918 444561
rect 101154 444325 107918 444561
rect 108154 444325 114918 444561
rect 115154 444325 121918 444561
rect 122154 444325 128918 444561
rect 129154 444325 135918 444561
rect 136154 444325 142918 444561
rect 143154 444325 149918 444561
rect 150154 444325 156918 444561
rect 157154 444325 163918 444561
rect 164154 444325 170918 444561
rect 171154 444325 177918 444561
rect 178154 444325 184918 444561
rect 185154 444325 191918 444561
rect 192154 444325 198918 444561
rect 199154 444325 205918 444561
rect 206154 444325 212918 444561
rect 213154 444325 219918 444561
rect 220154 444325 226918 444561
rect 227154 444325 233918 444561
rect 234154 444325 240918 444561
rect 241154 444325 247918 444561
rect 248154 444325 254918 444561
rect 255154 444325 261918 444561
rect 262154 444325 268918 444561
rect 269154 444325 275918 444561
rect 276154 444325 282918 444561
rect 283154 444325 289918 444561
rect 290154 444325 296918 444561
rect 297154 444325 303918 444561
rect 304154 444325 310918 444561
rect 311154 444325 317918 444561
rect 318154 444325 324918 444561
rect 325154 444325 331918 444561
rect 332154 444325 338918 444561
rect 339154 444325 345918 444561
rect 346154 444325 352918 444561
rect 353154 444325 359918 444561
rect 360154 444325 366918 444561
rect 367154 444325 373918 444561
rect 374154 444325 380918 444561
rect 381154 444325 387918 444561
rect 388154 444325 394918 444561
rect 395154 444325 401918 444561
rect 402154 444325 408918 444561
rect 409154 444325 415918 444561
rect 416154 444325 422918 444561
rect 423154 444325 429918 444561
rect 430154 444325 436918 444561
rect 437154 444325 443918 444561
rect 444154 444325 450918 444561
rect 451154 444325 457918 444561
rect 458154 444325 464918 444561
rect 465154 444325 471918 444561
rect 472154 444325 478918 444561
rect 479154 444325 485918 444561
rect 486154 444325 492918 444561
rect 493154 444325 499918 444561
rect 500154 444325 506918 444561
rect 507154 444325 513918 444561
rect 514154 444325 520918 444561
rect 521154 444325 527918 444561
rect 528154 444325 534918 444561
rect 535154 444325 541918 444561
rect 542154 444325 548918 444561
rect 549154 444325 555918 444561
rect 556154 444325 562918 444561
rect 563154 444325 569918 444561
rect 570154 444325 576918 444561
rect 577154 444325 587570 444561
rect 587806 444325 587890 444561
rect 588126 444325 588210 444561
rect 588446 444325 588530 444561
rect 588766 444325 588874 444561
rect -4950 444283 588874 444325
rect -4950 443494 588874 443536
rect -4950 443258 -3090 443494
rect -2854 443258 -2770 443494
rect -2534 443258 -2450 443494
rect -2214 443258 -2130 443494
rect -1894 443258 1186 443494
rect 1422 443258 8186 443494
rect 8422 443258 15186 443494
rect 15422 443258 22186 443494
rect 22422 443258 29186 443494
rect 29422 443258 36186 443494
rect 36422 443258 43186 443494
rect 43422 443258 50186 443494
rect 50422 443258 57186 443494
rect 57422 443258 64186 443494
rect 64422 443258 71186 443494
rect 71422 443258 78186 443494
rect 78422 443258 85186 443494
rect 85422 443258 92186 443494
rect 92422 443258 99186 443494
rect 99422 443258 106186 443494
rect 106422 443258 113186 443494
rect 113422 443258 120186 443494
rect 120422 443258 127186 443494
rect 127422 443258 134186 443494
rect 134422 443258 141186 443494
rect 141422 443258 148186 443494
rect 148422 443258 155186 443494
rect 155422 443258 162186 443494
rect 162422 443258 169186 443494
rect 169422 443258 176186 443494
rect 176422 443258 183186 443494
rect 183422 443258 190186 443494
rect 190422 443258 197186 443494
rect 197422 443258 204186 443494
rect 204422 443258 211186 443494
rect 211422 443258 218186 443494
rect 218422 443258 225186 443494
rect 225422 443258 232186 443494
rect 232422 443258 239186 443494
rect 239422 443258 246186 443494
rect 246422 443258 253186 443494
rect 253422 443258 260186 443494
rect 260422 443258 267186 443494
rect 267422 443258 274186 443494
rect 274422 443258 281186 443494
rect 281422 443258 288186 443494
rect 288422 443258 295186 443494
rect 295422 443258 302186 443494
rect 302422 443258 309186 443494
rect 309422 443258 316186 443494
rect 316422 443258 323186 443494
rect 323422 443258 330186 443494
rect 330422 443258 337186 443494
rect 337422 443258 344186 443494
rect 344422 443258 351186 443494
rect 351422 443258 358186 443494
rect 358422 443258 365186 443494
rect 365422 443258 372186 443494
rect 372422 443258 379186 443494
rect 379422 443258 386186 443494
rect 386422 443258 393186 443494
rect 393422 443258 400186 443494
rect 400422 443258 407186 443494
rect 407422 443258 414186 443494
rect 414422 443258 421186 443494
rect 421422 443258 428186 443494
rect 428422 443258 435186 443494
rect 435422 443258 442186 443494
rect 442422 443258 449186 443494
rect 449422 443258 456186 443494
rect 456422 443258 463186 443494
rect 463422 443258 470186 443494
rect 470422 443258 477186 443494
rect 477422 443258 484186 443494
rect 484422 443258 491186 443494
rect 491422 443258 498186 443494
rect 498422 443258 505186 443494
rect 505422 443258 512186 443494
rect 512422 443258 519186 443494
rect 519422 443258 526186 443494
rect 526422 443258 533186 443494
rect 533422 443258 540186 443494
rect 540422 443258 547186 443494
rect 547422 443258 554186 443494
rect 554422 443258 561186 443494
rect 561422 443258 568186 443494
rect 568422 443258 575186 443494
rect 575422 443258 582186 443494
rect 582422 443258 585818 443494
rect 586054 443258 586138 443494
rect 586374 443258 586458 443494
rect 586694 443258 586778 443494
rect 587014 443258 588874 443494
rect -4950 443216 588874 443258
rect -4950 437561 588874 437603
rect -4950 437325 -4842 437561
rect -4606 437325 -4522 437561
rect -4286 437325 -4202 437561
rect -3966 437325 -3882 437561
rect -3646 437325 2918 437561
rect 3154 437325 9918 437561
rect 10154 437325 16918 437561
rect 17154 437325 23918 437561
rect 24154 437325 30918 437561
rect 31154 437325 37918 437561
rect 38154 437325 44918 437561
rect 45154 437325 51918 437561
rect 52154 437325 58918 437561
rect 59154 437325 65918 437561
rect 66154 437325 72918 437561
rect 73154 437325 79918 437561
rect 80154 437325 86918 437561
rect 87154 437325 93918 437561
rect 94154 437325 100918 437561
rect 101154 437325 107918 437561
rect 108154 437325 114918 437561
rect 115154 437325 121918 437561
rect 122154 437325 128918 437561
rect 129154 437325 135918 437561
rect 136154 437325 142918 437561
rect 143154 437325 149918 437561
rect 150154 437325 156918 437561
rect 157154 437325 163918 437561
rect 164154 437325 170918 437561
rect 171154 437325 177918 437561
rect 178154 437325 184918 437561
rect 185154 437325 191918 437561
rect 192154 437325 198918 437561
rect 199154 437325 205918 437561
rect 206154 437325 212918 437561
rect 213154 437325 219918 437561
rect 220154 437325 226918 437561
rect 227154 437325 233918 437561
rect 234154 437325 240918 437561
rect 241154 437325 247918 437561
rect 248154 437325 254918 437561
rect 255154 437325 261918 437561
rect 262154 437325 268918 437561
rect 269154 437325 275918 437561
rect 276154 437325 282918 437561
rect 283154 437325 289918 437561
rect 290154 437325 296918 437561
rect 297154 437325 303918 437561
rect 304154 437325 310918 437561
rect 311154 437325 317918 437561
rect 318154 437325 324918 437561
rect 325154 437325 331918 437561
rect 332154 437325 338918 437561
rect 339154 437325 345918 437561
rect 346154 437325 352918 437561
rect 353154 437325 359918 437561
rect 360154 437325 366918 437561
rect 367154 437325 373918 437561
rect 374154 437325 380918 437561
rect 381154 437325 387918 437561
rect 388154 437325 394918 437561
rect 395154 437325 401918 437561
rect 402154 437325 408918 437561
rect 409154 437325 415918 437561
rect 416154 437325 422918 437561
rect 423154 437325 429918 437561
rect 430154 437325 436918 437561
rect 437154 437325 443918 437561
rect 444154 437325 450918 437561
rect 451154 437325 457918 437561
rect 458154 437325 464918 437561
rect 465154 437325 471918 437561
rect 472154 437325 478918 437561
rect 479154 437325 485918 437561
rect 486154 437325 492918 437561
rect 493154 437325 499918 437561
rect 500154 437325 506918 437561
rect 507154 437325 513918 437561
rect 514154 437325 520918 437561
rect 521154 437325 527918 437561
rect 528154 437325 534918 437561
rect 535154 437325 541918 437561
rect 542154 437325 548918 437561
rect 549154 437325 555918 437561
rect 556154 437325 562918 437561
rect 563154 437325 569918 437561
rect 570154 437325 576918 437561
rect 577154 437325 587570 437561
rect 587806 437325 587890 437561
rect 588126 437325 588210 437561
rect 588446 437325 588530 437561
rect 588766 437325 588874 437561
rect -4950 437283 588874 437325
rect -4950 436494 588874 436536
rect -4950 436258 -3090 436494
rect -2854 436258 -2770 436494
rect -2534 436258 -2450 436494
rect -2214 436258 -2130 436494
rect -1894 436258 1186 436494
rect 1422 436258 8186 436494
rect 8422 436258 15186 436494
rect 15422 436258 22186 436494
rect 22422 436258 29186 436494
rect 29422 436258 36186 436494
rect 36422 436258 43186 436494
rect 43422 436258 50186 436494
rect 50422 436258 57186 436494
rect 57422 436258 64186 436494
rect 64422 436258 71186 436494
rect 71422 436258 78186 436494
rect 78422 436258 85186 436494
rect 85422 436258 92186 436494
rect 92422 436258 99186 436494
rect 99422 436258 106186 436494
rect 106422 436258 113186 436494
rect 113422 436258 120186 436494
rect 120422 436258 127186 436494
rect 127422 436258 134186 436494
rect 134422 436258 141186 436494
rect 141422 436258 148186 436494
rect 148422 436258 155186 436494
rect 155422 436258 162186 436494
rect 162422 436258 169186 436494
rect 169422 436258 176186 436494
rect 176422 436258 183186 436494
rect 183422 436258 190186 436494
rect 190422 436258 197186 436494
rect 197422 436258 204186 436494
rect 204422 436258 211186 436494
rect 211422 436258 218186 436494
rect 218422 436258 225186 436494
rect 225422 436258 232186 436494
rect 232422 436258 239186 436494
rect 239422 436258 246186 436494
rect 246422 436258 253186 436494
rect 253422 436258 260186 436494
rect 260422 436258 267186 436494
rect 267422 436258 274186 436494
rect 274422 436258 281186 436494
rect 281422 436258 288186 436494
rect 288422 436258 295186 436494
rect 295422 436258 302186 436494
rect 302422 436258 309186 436494
rect 309422 436258 316186 436494
rect 316422 436258 323186 436494
rect 323422 436258 330186 436494
rect 330422 436258 337186 436494
rect 337422 436258 344186 436494
rect 344422 436258 351186 436494
rect 351422 436258 358186 436494
rect 358422 436258 365186 436494
rect 365422 436258 372186 436494
rect 372422 436258 379186 436494
rect 379422 436258 386186 436494
rect 386422 436258 393186 436494
rect 393422 436258 400186 436494
rect 400422 436258 407186 436494
rect 407422 436258 414186 436494
rect 414422 436258 421186 436494
rect 421422 436258 428186 436494
rect 428422 436258 435186 436494
rect 435422 436258 442186 436494
rect 442422 436258 449186 436494
rect 449422 436258 456186 436494
rect 456422 436258 463186 436494
rect 463422 436258 470186 436494
rect 470422 436258 477186 436494
rect 477422 436258 484186 436494
rect 484422 436258 491186 436494
rect 491422 436258 498186 436494
rect 498422 436258 505186 436494
rect 505422 436258 512186 436494
rect 512422 436258 519186 436494
rect 519422 436258 526186 436494
rect 526422 436258 533186 436494
rect 533422 436258 540186 436494
rect 540422 436258 547186 436494
rect 547422 436258 554186 436494
rect 554422 436258 561186 436494
rect 561422 436258 568186 436494
rect 568422 436258 575186 436494
rect 575422 436258 582186 436494
rect 582422 436258 585818 436494
rect 586054 436258 586138 436494
rect 586374 436258 586458 436494
rect 586694 436258 586778 436494
rect 587014 436258 588874 436494
rect -4950 436216 588874 436258
rect -4950 430561 588874 430603
rect -4950 430325 -4842 430561
rect -4606 430325 -4522 430561
rect -4286 430325 -4202 430561
rect -3966 430325 -3882 430561
rect -3646 430325 2918 430561
rect 3154 430325 9918 430561
rect 10154 430325 16918 430561
rect 17154 430325 23918 430561
rect 24154 430325 30918 430561
rect 31154 430325 37918 430561
rect 38154 430325 44918 430561
rect 45154 430325 51918 430561
rect 52154 430325 58918 430561
rect 59154 430325 65918 430561
rect 66154 430325 72918 430561
rect 73154 430325 79918 430561
rect 80154 430325 86918 430561
rect 87154 430325 93918 430561
rect 94154 430325 100918 430561
rect 101154 430325 107918 430561
rect 108154 430325 114918 430561
rect 115154 430325 121918 430561
rect 122154 430325 128918 430561
rect 129154 430325 135918 430561
rect 136154 430325 142918 430561
rect 143154 430325 149918 430561
rect 150154 430325 156918 430561
rect 157154 430325 163918 430561
rect 164154 430325 170918 430561
rect 171154 430325 177918 430561
rect 178154 430325 184918 430561
rect 185154 430325 191918 430561
rect 192154 430325 198918 430561
rect 199154 430325 205918 430561
rect 206154 430325 212918 430561
rect 213154 430325 219918 430561
rect 220154 430325 226918 430561
rect 227154 430325 233918 430561
rect 234154 430325 240918 430561
rect 241154 430325 247918 430561
rect 248154 430325 254918 430561
rect 255154 430325 261918 430561
rect 262154 430325 268918 430561
rect 269154 430325 275918 430561
rect 276154 430325 282918 430561
rect 283154 430325 289918 430561
rect 290154 430325 296918 430561
rect 297154 430325 303918 430561
rect 304154 430325 310918 430561
rect 311154 430325 317918 430561
rect 318154 430325 324918 430561
rect 325154 430325 331918 430561
rect 332154 430325 338918 430561
rect 339154 430325 345918 430561
rect 346154 430325 352918 430561
rect 353154 430325 359918 430561
rect 360154 430325 366918 430561
rect 367154 430325 373918 430561
rect 374154 430325 380918 430561
rect 381154 430325 387918 430561
rect 388154 430325 394918 430561
rect 395154 430325 401918 430561
rect 402154 430325 408918 430561
rect 409154 430325 415918 430561
rect 416154 430325 422918 430561
rect 423154 430325 429918 430561
rect 430154 430325 436918 430561
rect 437154 430325 443918 430561
rect 444154 430325 450918 430561
rect 451154 430325 457918 430561
rect 458154 430325 464918 430561
rect 465154 430325 471918 430561
rect 472154 430325 478918 430561
rect 479154 430325 485918 430561
rect 486154 430325 492918 430561
rect 493154 430325 499918 430561
rect 500154 430325 506918 430561
rect 507154 430325 513918 430561
rect 514154 430325 520918 430561
rect 521154 430325 527918 430561
rect 528154 430325 534918 430561
rect 535154 430325 541918 430561
rect 542154 430325 548918 430561
rect 549154 430325 555918 430561
rect 556154 430325 562918 430561
rect 563154 430325 569918 430561
rect 570154 430325 576918 430561
rect 577154 430325 587570 430561
rect 587806 430325 587890 430561
rect 588126 430325 588210 430561
rect 588446 430325 588530 430561
rect 588766 430325 588874 430561
rect -4950 430283 588874 430325
rect -4950 429494 588874 429536
rect -4950 429258 -3090 429494
rect -2854 429258 -2770 429494
rect -2534 429258 -2450 429494
rect -2214 429258 -2130 429494
rect -1894 429258 1186 429494
rect 1422 429258 8186 429494
rect 8422 429258 15186 429494
rect 15422 429258 22186 429494
rect 22422 429258 29186 429494
rect 29422 429258 36186 429494
rect 36422 429258 43186 429494
rect 43422 429258 50186 429494
rect 50422 429258 57186 429494
rect 57422 429258 64186 429494
rect 64422 429258 71186 429494
rect 71422 429258 78186 429494
rect 78422 429258 85186 429494
rect 85422 429258 92186 429494
rect 92422 429258 99186 429494
rect 99422 429258 106186 429494
rect 106422 429258 113186 429494
rect 113422 429258 120186 429494
rect 120422 429258 127186 429494
rect 127422 429258 134186 429494
rect 134422 429258 141186 429494
rect 141422 429258 148186 429494
rect 148422 429258 155186 429494
rect 155422 429258 162186 429494
rect 162422 429258 169186 429494
rect 169422 429258 176186 429494
rect 176422 429258 183186 429494
rect 183422 429258 190186 429494
rect 190422 429258 197186 429494
rect 197422 429258 204186 429494
rect 204422 429258 211186 429494
rect 211422 429258 218186 429494
rect 218422 429258 225186 429494
rect 225422 429258 232186 429494
rect 232422 429258 239186 429494
rect 239422 429258 246186 429494
rect 246422 429258 253186 429494
rect 253422 429258 260186 429494
rect 260422 429258 267186 429494
rect 267422 429258 274186 429494
rect 274422 429258 281186 429494
rect 281422 429258 288186 429494
rect 288422 429258 295186 429494
rect 295422 429258 302186 429494
rect 302422 429258 309186 429494
rect 309422 429258 316186 429494
rect 316422 429258 323186 429494
rect 323422 429258 330186 429494
rect 330422 429258 337186 429494
rect 337422 429258 344186 429494
rect 344422 429258 351186 429494
rect 351422 429258 358186 429494
rect 358422 429258 365186 429494
rect 365422 429258 372186 429494
rect 372422 429258 379186 429494
rect 379422 429258 386186 429494
rect 386422 429258 393186 429494
rect 393422 429258 400186 429494
rect 400422 429258 407186 429494
rect 407422 429258 414186 429494
rect 414422 429258 421186 429494
rect 421422 429258 428186 429494
rect 428422 429258 435186 429494
rect 435422 429258 442186 429494
rect 442422 429258 449186 429494
rect 449422 429258 456186 429494
rect 456422 429258 463186 429494
rect 463422 429258 470186 429494
rect 470422 429258 477186 429494
rect 477422 429258 484186 429494
rect 484422 429258 491186 429494
rect 491422 429258 498186 429494
rect 498422 429258 505186 429494
rect 505422 429258 512186 429494
rect 512422 429258 519186 429494
rect 519422 429258 526186 429494
rect 526422 429258 533186 429494
rect 533422 429258 540186 429494
rect 540422 429258 547186 429494
rect 547422 429258 554186 429494
rect 554422 429258 561186 429494
rect 561422 429258 568186 429494
rect 568422 429258 575186 429494
rect 575422 429258 582186 429494
rect 582422 429258 585818 429494
rect 586054 429258 586138 429494
rect 586374 429258 586458 429494
rect 586694 429258 586778 429494
rect 587014 429258 588874 429494
rect -4950 429216 588874 429258
rect -4950 423561 588874 423603
rect -4950 423325 -4842 423561
rect -4606 423325 -4522 423561
rect -4286 423325 -4202 423561
rect -3966 423325 -3882 423561
rect -3646 423325 2918 423561
rect 3154 423325 9918 423561
rect 10154 423325 16918 423561
rect 17154 423325 23918 423561
rect 24154 423325 30918 423561
rect 31154 423325 37918 423561
rect 38154 423325 44918 423561
rect 45154 423325 51918 423561
rect 52154 423325 58918 423561
rect 59154 423325 65918 423561
rect 66154 423325 72918 423561
rect 73154 423325 79918 423561
rect 80154 423325 86918 423561
rect 87154 423325 93918 423561
rect 94154 423325 100918 423561
rect 101154 423325 107918 423561
rect 108154 423325 114918 423561
rect 115154 423325 121918 423561
rect 122154 423325 128918 423561
rect 129154 423325 135918 423561
rect 136154 423325 142918 423561
rect 143154 423325 149918 423561
rect 150154 423325 156918 423561
rect 157154 423325 163918 423561
rect 164154 423325 170918 423561
rect 171154 423325 177918 423561
rect 178154 423325 184918 423561
rect 185154 423325 191918 423561
rect 192154 423325 198918 423561
rect 199154 423325 205918 423561
rect 206154 423325 212918 423561
rect 213154 423325 219918 423561
rect 220154 423325 226918 423561
rect 227154 423325 233918 423561
rect 234154 423325 240918 423561
rect 241154 423325 247918 423561
rect 248154 423325 254918 423561
rect 255154 423325 261918 423561
rect 262154 423325 268918 423561
rect 269154 423325 275918 423561
rect 276154 423325 282918 423561
rect 283154 423325 289918 423561
rect 290154 423325 296918 423561
rect 297154 423325 303918 423561
rect 304154 423325 310918 423561
rect 311154 423325 317918 423561
rect 318154 423325 324918 423561
rect 325154 423325 331918 423561
rect 332154 423325 338918 423561
rect 339154 423325 345918 423561
rect 346154 423325 352918 423561
rect 353154 423325 359918 423561
rect 360154 423325 366918 423561
rect 367154 423325 373918 423561
rect 374154 423325 380918 423561
rect 381154 423325 387918 423561
rect 388154 423325 394918 423561
rect 395154 423325 401918 423561
rect 402154 423325 408918 423561
rect 409154 423325 415918 423561
rect 416154 423325 422918 423561
rect 423154 423325 429918 423561
rect 430154 423325 436918 423561
rect 437154 423325 443918 423561
rect 444154 423325 450918 423561
rect 451154 423325 457918 423561
rect 458154 423325 464918 423561
rect 465154 423325 471918 423561
rect 472154 423325 478918 423561
rect 479154 423325 485918 423561
rect 486154 423325 492918 423561
rect 493154 423325 499918 423561
rect 500154 423325 506918 423561
rect 507154 423325 513918 423561
rect 514154 423325 520918 423561
rect 521154 423325 527918 423561
rect 528154 423325 534918 423561
rect 535154 423325 541918 423561
rect 542154 423325 548918 423561
rect 549154 423325 555918 423561
rect 556154 423325 562918 423561
rect 563154 423325 569918 423561
rect 570154 423325 576918 423561
rect 577154 423325 587570 423561
rect 587806 423325 587890 423561
rect 588126 423325 588210 423561
rect 588446 423325 588530 423561
rect 588766 423325 588874 423561
rect -4950 423283 588874 423325
rect -4950 422494 588874 422536
rect -4950 422258 -3090 422494
rect -2854 422258 -2770 422494
rect -2534 422258 -2450 422494
rect -2214 422258 -2130 422494
rect -1894 422258 1186 422494
rect 1422 422258 8186 422494
rect 8422 422258 15186 422494
rect 15422 422258 22186 422494
rect 22422 422258 29186 422494
rect 29422 422258 36186 422494
rect 36422 422258 43186 422494
rect 43422 422258 50186 422494
rect 50422 422258 57186 422494
rect 57422 422258 64186 422494
rect 64422 422258 71186 422494
rect 71422 422258 78186 422494
rect 78422 422258 85186 422494
rect 85422 422258 92186 422494
rect 92422 422258 99186 422494
rect 99422 422258 106186 422494
rect 106422 422258 113186 422494
rect 113422 422258 120186 422494
rect 120422 422258 127186 422494
rect 127422 422258 134186 422494
rect 134422 422258 141186 422494
rect 141422 422258 148186 422494
rect 148422 422258 155186 422494
rect 155422 422258 162186 422494
rect 162422 422258 169186 422494
rect 169422 422258 176186 422494
rect 176422 422258 183186 422494
rect 183422 422258 190186 422494
rect 190422 422258 197186 422494
rect 197422 422258 204186 422494
rect 204422 422258 211186 422494
rect 211422 422258 218186 422494
rect 218422 422258 225186 422494
rect 225422 422258 232186 422494
rect 232422 422258 239186 422494
rect 239422 422258 246186 422494
rect 246422 422258 253186 422494
rect 253422 422258 260186 422494
rect 260422 422258 267186 422494
rect 267422 422258 274186 422494
rect 274422 422258 281186 422494
rect 281422 422258 288186 422494
rect 288422 422258 295186 422494
rect 295422 422258 302186 422494
rect 302422 422258 309186 422494
rect 309422 422258 316186 422494
rect 316422 422258 323186 422494
rect 323422 422258 330186 422494
rect 330422 422258 337186 422494
rect 337422 422258 344186 422494
rect 344422 422258 351186 422494
rect 351422 422258 358186 422494
rect 358422 422258 365186 422494
rect 365422 422258 372186 422494
rect 372422 422258 379186 422494
rect 379422 422258 386186 422494
rect 386422 422258 393186 422494
rect 393422 422258 400186 422494
rect 400422 422258 407186 422494
rect 407422 422258 414186 422494
rect 414422 422258 421186 422494
rect 421422 422258 428186 422494
rect 428422 422258 435186 422494
rect 435422 422258 442186 422494
rect 442422 422258 449186 422494
rect 449422 422258 456186 422494
rect 456422 422258 463186 422494
rect 463422 422258 470186 422494
rect 470422 422258 477186 422494
rect 477422 422258 484186 422494
rect 484422 422258 491186 422494
rect 491422 422258 498186 422494
rect 498422 422258 505186 422494
rect 505422 422258 512186 422494
rect 512422 422258 519186 422494
rect 519422 422258 526186 422494
rect 526422 422258 533186 422494
rect 533422 422258 540186 422494
rect 540422 422258 547186 422494
rect 547422 422258 554186 422494
rect 554422 422258 561186 422494
rect 561422 422258 568186 422494
rect 568422 422258 575186 422494
rect 575422 422258 582186 422494
rect 582422 422258 585818 422494
rect 586054 422258 586138 422494
rect 586374 422258 586458 422494
rect 586694 422258 586778 422494
rect 587014 422258 588874 422494
rect -4950 422216 588874 422258
rect -4950 416561 588874 416603
rect -4950 416325 -4842 416561
rect -4606 416325 -4522 416561
rect -4286 416325 -4202 416561
rect -3966 416325 -3882 416561
rect -3646 416325 2918 416561
rect 3154 416325 9918 416561
rect 10154 416325 16918 416561
rect 17154 416325 23918 416561
rect 24154 416325 30918 416561
rect 31154 416325 37918 416561
rect 38154 416325 44918 416561
rect 45154 416325 51918 416561
rect 52154 416325 58918 416561
rect 59154 416325 65918 416561
rect 66154 416325 72918 416561
rect 73154 416325 79918 416561
rect 80154 416325 86918 416561
rect 87154 416325 93918 416561
rect 94154 416325 100918 416561
rect 101154 416325 107918 416561
rect 108154 416325 114918 416561
rect 115154 416325 121918 416561
rect 122154 416325 128918 416561
rect 129154 416325 135918 416561
rect 136154 416325 142918 416561
rect 143154 416325 149918 416561
rect 150154 416325 156918 416561
rect 157154 416325 163918 416561
rect 164154 416325 170918 416561
rect 171154 416325 177918 416561
rect 178154 416325 184918 416561
rect 185154 416325 191918 416561
rect 192154 416325 198918 416561
rect 199154 416325 205918 416561
rect 206154 416325 212918 416561
rect 213154 416325 219918 416561
rect 220154 416325 226918 416561
rect 227154 416325 233918 416561
rect 234154 416325 240918 416561
rect 241154 416325 247918 416561
rect 248154 416325 254918 416561
rect 255154 416325 261918 416561
rect 262154 416325 268918 416561
rect 269154 416325 275918 416561
rect 276154 416325 282918 416561
rect 283154 416325 289918 416561
rect 290154 416325 296918 416561
rect 297154 416325 303918 416561
rect 304154 416325 310918 416561
rect 311154 416325 317918 416561
rect 318154 416325 324918 416561
rect 325154 416325 331918 416561
rect 332154 416325 338918 416561
rect 339154 416325 345918 416561
rect 346154 416325 352918 416561
rect 353154 416325 359918 416561
rect 360154 416325 366918 416561
rect 367154 416325 373918 416561
rect 374154 416325 380918 416561
rect 381154 416325 387918 416561
rect 388154 416325 394918 416561
rect 395154 416325 401918 416561
rect 402154 416325 408918 416561
rect 409154 416325 415918 416561
rect 416154 416325 422918 416561
rect 423154 416325 429918 416561
rect 430154 416325 436918 416561
rect 437154 416325 443918 416561
rect 444154 416325 450918 416561
rect 451154 416325 457918 416561
rect 458154 416325 464918 416561
rect 465154 416325 471918 416561
rect 472154 416325 478918 416561
rect 479154 416325 485918 416561
rect 486154 416325 492918 416561
rect 493154 416325 499918 416561
rect 500154 416325 506918 416561
rect 507154 416325 513918 416561
rect 514154 416325 520918 416561
rect 521154 416325 522850 416561
rect 523086 416325 524782 416561
rect 525018 416325 526714 416561
rect 526950 416325 527918 416561
rect 528154 416325 534918 416561
rect 535154 416325 541918 416561
rect 542154 416325 548918 416561
rect 549154 416325 555918 416561
rect 556154 416325 562918 416561
rect 563154 416325 569918 416561
rect 570154 416325 576918 416561
rect 577154 416325 587570 416561
rect 587806 416325 587890 416561
rect 588126 416325 588210 416561
rect 588446 416325 588530 416561
rect 588766 416325 588874 416561
rect -4950 416283 588874 416325
rect -4950 415494 588874 415536
rect -4950 415258 -3090 415494
rect -2854 415258 -2770 415494
rect -2534 415258 -2450 415494
rect -2214 415258 -2130 415494
rect -1894 415258 1186 415494
rect 1422 415258 8186 415494
rect 8422 415258 15186 415494
rect 15422 415258 22186 415494
rect 22422 415258 29186 415494
rect 29422 415258 36186 415494
rect 36422 415258 43186 415494
rect 43422 415258 50186 415494
rect 50422 415258 57186 415494
rect 57422 415258 64186 415494
rect 64422 415258 71186 415494
rect 71422 415258 78186 415494
rect 78422 415258 85186 415494
rect 85422 415258 92186 415494
rect 92422 415258 99186 415494
rect 99422 415258 106186 415494
rect 106422 415258 113186 415494
rect 113422 415258 120186 415494
rect 120422 415258 127186 415494
rect 127422 415258 134186 415494
rect 134422 415258 141186 415494
rect 141422 415258 148186 415494
rect 148422 415258 155186 415494
rect 155422 415258 162186 415494
rect 162422 415258 169186 415494
rect 169422 415258 176186 415494
rect 176422 415258 183186 415494
rect 183422 415258 190186 415494
rect 190422 415258 197186 415494
rect 197422 415258 204186 415494
rect 204422 415258 211186 415494
rect 211422 415258 218186 415494
rect 218422 415258 225186 415494
rect 225422 415258 232186 415494
rect 232422 415258 239186 415494
rect 239422 415258 246186 415494
rect 246422 415258 253186 415494
rect 253422 415258 260186 415494
rect 260422 415258 267186 415494
rect 267422 415258 274186 415494
rect 274422 415258 281186 415494
rect 281422 415258 288186 415494
rect 288422 415258 295186 415494
rect 295422 415258 302186 415494
rect 302422 415258 309186 415494
rect 309422 415258 316186 415494
rect 316422 415258 323186 415494
rect 323422 415258 330186 415494
rect 330422 415258 337186 415494
rect 337422 415258 344186 415494
rect 344422 415258 351186 415494
rect 351422 415258 358186 415494
rect 358422 415258 365186 415494
rect 365422 415258 372186 415494
rect 372422 415258 379186 415494
rect 379422 415258 386186 415494
rect 386422 415258 393186 415494
rect 393422 415258 400186 415494
rect 400422 415258 407186 415494
rect 407422 415258 414186 415494
rect 414422 415258 421186 415494
rect 421422 415258 428186 415494
rect 428422 415258 435186 415494
rect 435422 415258 442186 415494
rect 442422 415258 449186 415494
rect 449422 415258 456186 415494
rect 456422 415258 463186 415494
rect 463422 415258 470186 415494
rect 470422 415258 477186 415494
rect 477422 415258 484186 415494
rect 484422 415258 491186 415494
rect 491422 415258 498186 415494
rect 498422 415258 505186 415494
rect 505422 415258 512186 415494
rect 512422 415258 519186 415494
rect 519422 415258 519952 415494
rect 520188 415258 521884 415494
rect 522120 415258 523816 415494
rect 524052 415258 525748 415494
rect 525984 415258 533186 415494
rect 533422 415258 540186 415494
rect 540422 415258 547186 415494
rect 547422 415258 554186 415494
rect 554422 415258 561186 415494
rect 561422 415258 568186 415494
rect 568422 415258 575186 415494
rect 575422 415258 582186 415494
rect 582422 415258 585818 415494
rect 586054 415258 586138 415494
rect 586374 415258 586458 415494
rect 586694 415258 586778 415494
rect 587014 415258 588874 415494
rect -4950 415216 588874 415258
rect -4950 409561 588874 409603
rect -4950 409325 -4842 409561
rect -4606 409325 -4522 409561
rect -4286 409325 -4202 409561
rect -3966 409325 -3882 409561
rect -3646 409325 2918 409561
rect 3154 409325 9918 409561
rect 10154 409325 16918 409561
rect 17154 409325 23918 409561
rect 24154 409325 30918 409561
rect 31154 409325 37918 409561
rect 38154 409325 44918 409561
rect 45154 409325 51918 409561
rect 52154 409325 58918 409561
rect 59154 409325 65918 409561
rect 66154 409325 72918 409561
rect 73154 409325 79918 409561
rect 80154 409325 86918 409561
rect 87154 409325 93918 409561
rect 94154 409325 100918 409561
rect 101154 409325 107918 409561
rect 108154 409325 114918 409561
rect 115154 409325 121918 409561
rect 122154 409325 128918 409561
rect 129154 409325 135918 409561
rect 136154 409325 142918 409561
rect 143154 409325 149918 409561
rect 150154 409325 156918 409561
rect 157154 409325 163918 409561
rect 164154 409325 170918 409561
rect 171154 409325 177918 409561
rect 178154 409325 184918 409561
rect 185154 409325 191918 409561
rect 192154 409325 198918 409561
rect 199154 409325 205918 409561
rect 206154 409325 212918 409561
rect 213154 409325 219918 409561
rect 220154 409325 226918 409561
rect 227154 409325 233918 409561
rect 234154 409325 240918 409561
rect 241154 409325 247918 409561
rect 248154 409325 254918 409561
rect 255154 409325 261918 409561
rect 262154 409325 268918 409561
rect 269154 409325 275918 409561
rect 276154 409325 282918 409561
rect 283154 409325 289918 409561
rect 290154 409325 296918 409561
rect 297154 409325 303918 409561
rect 304154 409325 310918 409561
rect 311154 409325 317918 409561
rect 318154 409325 324918 409561
rect 325154 409325 331918 409561
rect 332154 409325 338918 409561
rect 339154 409325 345918 409561
rect 346154 409325 352918 409561
rect 353154 409325 359918 409561
rect 360154 409325 366918 409561
rect 367154 409325 373918 409561
rect 374154 409325 380918 409561
rect 381154 409325 387918 409561
rect 388154 409325 394918 409561
rect 395154 409325 401918 409561
rect 402154 409325 408918 409561
rect 409154 409325 415918 409561
rect 416154 409325 422918 409561
rect 423154 409325 429918 409561
rect 430154 409325 436918 409561
rect 437154 409325 443918 409561
rect 444154 409325 450918 409561
rect 451154 409325 457918 409561
rect 458154 409325 464918 409561
rect 465154 409325 471918 409561
rect 472154 409325 478918 409561
rect 479154 409325 485918 409561
rect 486154 409325 492918 409561
rect 493154 409325 499918 409561
rect 500154 409325 506918 409561
rect 507154 409325 513918 409561
rect 514154 409325 520918 409561
rect 521154 409325 522850 409561
rect 523086 409325 524782 409561
rect 525018 409325 526714 409561
rect 526950 409325 527918 409561
rect 528154 409325 534918 409561
rect 535154 409325 541918 409561
rect 542154 409325 548918 409561
rect 549154 409325 555918 409561
rect 556154 409325 562918 409561
rect 563154 409325 569918 409561
rect 570154 409325 576918 409561
rect 577154 409325 587570 409561
rect 587806 409325 587890 409561
rect 588126 409325 588210 409561
rect 588446 409325 588530 409561
rect 588766 409325 588874 409561
rect -4950 409283 588874 409325
rect -4950 408494 588874 408536
rect -4950 408258 -3090 408494
rect -2854 408258 -2770 408494
rect -2534 408258 -2450 408494
rect -2214 408258 -2130 408494
rect -1894 408258 1186 408494
rect 1422 408258 8186 408494
rect 8422 408258 15186 408494
rect 15422 408258 22186 408494
rect 22422 408258 29186 408494
rect 29422 408258 36186 408494
rect 36422 408258 43186 408494
rect 43422 408258 50186 408494
rect 50422 408258 57186 408494
rect 57422 408258 64186 408494
rect 64422 408258 71186 408494
rect 71422 408258 78186 408494
rect 78422 408258 85186 408494
rect 85422 408258 92186 408494
rect 92422 408258 99186 408494
rect 99422 408258 106186 408494
rect 106422 408258 113186 408494
rect 113422 408258 120186 408494
rect 120422 408258 127186 408494
rect 127422 408258 134186 408494
rect 134422 408258 141186 408494
rect 141422 408258 148186 408494
rect 148422 408258 155186 408494
rect 155422 408258 162186 408494
rect 162422 408258 169186 408494
rect 169422 408258 176186 408494
rect 176422 408258 183186 408494
rect 183422 408258 190186 408494
rect 190422 408258 197186 408494
rect 197422 408258 204186 408494
rect 204422 408258 211186 408494
rect 211422 408258 218186 408494
rect 218422 408258 225186 408494
rect 225422 408258 232186 408494
rect 232422 408258 239186 408494
rect 239422 408258 246186 408494
rect 246422 408258 253186 408494
rect 253422 408258 260186 408494
rect 260422 408258 267186 408494
rect 267422 408258 274186 408494
rect 274422 408258 281186 408494
rect 281422 408258 288186 408494
rect 288422 408258 295186 408494
rect 295422 408258 302186 408494
rect 302422 408258 309186 408494
rect 309422 408258 316186 408494
rect 316422 408258 323186 408494
rect 323422 408258 330186 408494
rect 330422 408258 337186 408494
rect 337422 408258 344186 408494
rect 344422 408258 351186 408494
rect 351422 408258 358186 408494
rect 358422 408258 365186 408494
rect 365422 408258 372186 408494
rect 372422 408258 379186 408494
rect 379422 408258 386186 408494
rect 386422 408258 393186 408494
rect 393422 408258 400186 408494
rect 400422 408258 407186 408494
rect 407422 408258 414186 408494
rect 414422 408258 421186 408494
rect 421422 408258 428186 408494
rect 428422 408258 435186 408494
rect 435422 408258 442186 408494
rect 442422 408258 449186 408494
rect 449422 408258 456186 408494
rect 456422 408258 463186 408494
rect 463422 408258 470186 408494
rect 470422 408258 477186 408494
rect 477422 408258 484186 408494
rect 484422 408258 491186 408494
rect 491422 408258 498186 408494
rect 498422 408258 505186 408494
rect 505422 408258 512186 408494
rect 512422 408258 519186 408494
rect 519422 408258 519952 408494
rect 520188 408258 521884 408494
rect 522120 408258 523816 408494
rect 524052 408258 525748 408494
rect 525984 408258 533186 408494
rect 533422 408258 540186 408494
rect 540422 408258 547186 408494
rect 547422 408258 554186 408494
rect 554422 408258 561186 408494
rect 561422 408258 568186 408494
rect 568422 408258 575186 408494
rect 575422 408258 582186 408494
rect 582422 408258 585818 408494
rect 586054 408258 586138 408494
rect 586374 408258 586458 408494
rect 586694 408258 586778 408494
rect 587014 408258 588874 408494
rect -4950 408216 588874 408258
rect -4950 402561 588874 402603
rect -4950 402325 -4842 402561
rect -4606 402325 -4522 402561
rect -4286 402325 -4202 402561
rect -3966 402325 -3882 402561
rect -3646 402325 2918 402561
rect 3154 402325 9918 402561
rect 10154 402325 16918 402561
rect 17154 402325 23918 402561
rect 24154 402325 30918 402561
rect 31154 402325 37918 402561
rect 38154 402325 44918 402561
rect 45154 402325 51918 402561
rect 52154 402325 58918 402561
rect 59154 402325 65918 402561
rect 66154 402325 72918 402561
rect 73154 402325 79918 402561
rect 80154 402325 86918 402561
rect 87154 402325 93918 402561
rect 94154 402325 100918 402561
rect 101154 402325 107918 402561
rect 108154 402325 114918 402561
rect 115154 402325 121918 402561
rect 122154 402325 128918 402561
rect 129154 402325 135918 402561
rect 136154 402325 142918 402561
rect 143154 402325 149918 402561
rect 150154 402325 156918 402561
rect 157154 402325 163918 402561
rect 164154 402325 170918 402561
rect 171154 402325 177918 402561
rect 178154 402325 184918 402561
rect 185154 402325 191918 402561
rect 192154 402325 198918 402561
rect 199154 402325 205918 402561
rect 206154 402325 212918 402561
rect 213154 402325 219918 402561
rect 220154 402325 226918 402561
rect 227154 402325 233918 402561
rect 234154 402325 240918 402561
rect 241154 402325 247918 402561
rect 248154 402325 254918 402561
rect 255154 402325 261918 402561
rect 262154 402325 268918 402561
rect 269154 402325 275918 402561
rect 276154 402325 282918 402561
rect 283154 402325 289918 402561
rect 290154 402325 296918 402561
rect 297154 402325 303918 402561
rect 304154 402325 310918 402561
rect 311154 402325 317918 402561
rect 318154 402325 324918 402561
rect 325154 402325 331918 402561
rect 332154 402325 338918 402561
rect 339154 402325 345918 402561
rect 346154 402325 352918 402561
rect 353154 402325 359918 402561
rect 360154 402325 366918 402561
rect 367154 402325 373918 402561
rect 374154 402325 380918 402561
rect 381154 402325 387918 402561
rect 388154 402325 394918 402561
rect 395154 402325 401918 402561
rect 402154 402325 408918 402561
rect 409154 402325 415918 402561
rect 416154 402325 422918 402561
rect 423154 402325 429918 402561
rect 430154 402325 436918 402561
rect 437154 402325 443918 402561
rect 444154 402325 450918 402561
rect 451154 402325 457918 402561
rect 458154 402325 464918 402561
rect 465154 402325 471918 402561
rect 472154 402325 478918 402561
rect 479154 402325 485918 402561
rect 486154 402325 492918 402561
rect 493154 402325 499918 402561
rect 500154 402325 506918 402561
rect 507154 402325 513918 402561
rect 514154 402325 520918 402561
rect 521154 402325 522850 402561
rect 523086 402325 524782 402561
rect 525018 402325 526714 402561
rect 526950 402325 527918 402561
rect 528154 402325 534918 402561
rect 535154 402325 541918 402561
rect 542154 402325 548918 402561
rect 549154 402325 555918 402561
rect 556154 402325 562918 402561
rect 563154 402325 569918 402561
rect 570154 402325 576918 402561
rect 577154 402325 587570 402561
rect 587806 402325 587890 402561
rect 588126 402325 588210 402561
rect 588446 402325 588530 402561
rect 588766 402325 588874 402561
rect -4950 402283 588874 402325
rect -4950 401494 588874 401536
rect -4950 401258 -3090 401494
rect -2854 401258 -2770 401494
rect -2534 401258 -2450 401494
rect -2214 401258 -2130 401494
rect -1894 401258 1186 401494
rect 1422 401258 8186 401494
rect 8422 401258 15186 401494
rect 15422 401258 22186 401494
rect 22422 401258 29186 401494
rect 29422 401258 36186 401494
rect 36422 401258 43186 401494
rect 43422 401258 50186 401494
rect 50422 401258 57186 401494
rect 57422 401258 64186 401494
rect 64422 401258 71186 401494
rect 71422 401258 78186 401494
rect 78422 401258 85186 401494
rect 85422 401258 92186 401494
rect 92422 401258 99186 401494
rect 99422 401258 106186 401494
rect 106422 401258 113186 401494
rect 113422 401258 120186 401494
rect 120422 401258 127186 401494
rect 127422 401258 134186 401494
rect 134422 401258 141186 401494
rect 141422 401258 148186 401494
rect 148422 401258 155186 401494
rect 155422 401258 162186 401494
rect 162422 401258 169186 401494
rect 169422 401258 176186 401494
rect 176422 401258 183186 401494
rect 183422 401258 190186 401494
rect 190422 401258 197186 401494
rect 197422 401258 204186 401494
rect 204422 401258 211186 401494
rect 211422 401258 218186 401494
rect 218422 401258 225186 401494
rect 225422 401258 232186 401494
rect 232422 401258 239186 401494
rect 239422 401258 246186 401494
rect 246422 401258 253186 401494
rect 253422 401258 260186 401494
rect 260422 401258 267186 401494
rect 267422 401258 274186 401494
rect 274422 401258 281186 401494
rect 281422 401258 288186 401494
rect 288422 401258 295186 401494
rect 295422 401258 302186 401494
rect 302422 401258 309186 401494
rect 309422 401258 316186 401494
rect 316422 401258 323186 401494
rect 323422 401258 330186 401494
rect 330422 401258 337186 401494
rect 337422 401258 344186 401494
rect 344422 401258 351186 401494
rect 351422 401258 358186 401494
rect 358422 401258 365186 401494
rect 365422 401258 372186 401494
rect 372422 401258 379186 401494
rect 379422 401258 386186 401494
rect 386422 401258 393186 401494
rect 393422 401258 400186 401494
rect 400422 401258 407186 401494
rect 407422 401258 414186 401494
rect 414422 401258 421186 401494
rect 421422 401258 428186 401494
rect 428422 401258 435186 401494
rect 435422 401258 442186 401494
rect 442422 401258 449186 401494
rect 449422 401258 456186 401494
rect 456422 401258 463186 401494
rect 463422 401258 470186 401494
rect 470422 401258 477186 401494
rect 477422 401258 484186 401494
rect 484422 401258 491186 401494
rect 491422 401258 498186 401494
rect 498422 401258 505186 401494
rect 505422 401258 512186 401494
rect 512422 401258 519186 401494
rect 519422 401258 533186 401494
rect 533422 401258 540186 401494
rect 540422 401258 547186 401494
rect 547422 401258 554186 401494
rect 554422 401258 561186 401494
rect 561422 401258 568186 401494
rect 568422 401258 575186 401494
rect 575422 401258 582186 401494
rect 582422 401258 585818 401494
rect 586054 401258 586138 401494
rect 586374 401258 586458 401494
rect 586694 401258 586778 401494
rect 587014 401258 588874 401494
rect -4950 401216 588874 401258
rect -4950 395561 588874 395603
rect -4950 395325 -4842 395561
rect -4606 395325 -4522 395561
rect -4286 395325 -4202 395561
rect -3966 395325 -3882 395561
rect -3646 395325 2918 395561
rect 3154 395325 9918 395561
rect 10154 395325 16918 395561
rect 17154 395325 23918 395561
rect 24154 395325 30918 395561
rect 31154 395325 37918 395561
rect 38154 395325 44918 395561
rect 45154 395325 51918 395561
rect 52154 395325 58918 395561
rect 59154 395325 65918 395561
rect 66154 395325 72918 395561
rect 73154 395325 79918 395561
rect 80154 395325 86918 395561
rect 87154 395325 93918 395561
rect 94154 395325 100918 395561
rect 101154 395325 107918 395561
rect 108154 395325 114918 395561
rect 115154 395325 121918 395561
rect 122154 395325 128918 395561
rect 129154 395325 135918 395561
rect 136154 395325 142918 395561
rect 143154 395325 149918 395561
rect 150154 395325 156918 395561
rect 157154 395325 163918 395561
rect 164154 395325 170918 395561
rect 171154 395325 177918 395561
rect 178154 395325 184918 395561
rect 185154 395325 191918 395561
rect 192154 395325 198918 395561
rect 199154 395325 205918 395561
rect 206154 395325 212918 395561
rect 213154 395325 219918 395561
rect 220154 395325 226918 395561
rect 227154 395325 233918 395561
rect 234154 395325 240918 395561
rect 241154 395325 247918 395561
rect 248154 395325 254918 395561
rect 255154 395325 261918 395561
rect 262154 395325 268918 395561
rect 269154 395325 275918 395561
rect 276154 395325 282918 395561
rect 283154 395325 289918 395561
rect 290154 395325 296918 395561
rect 297154 395325 303918 395561
rect 304154 395325 310918 395561
rect 311154 395325 317918 395561
rect 318154 395325 324918 395561
rect 325154 395325 331918 395561
rect 332154 395325 338918 395561
rect 339154 395325 345918 395561
rect 346154 395325 352918 395561
rect 353154 395325 359918 395561
rect 360154 395325 366918 395561
rect 367154 395325 373918 395561
rect 374154 395325 380918 395561
rect 381154 395325 387918 395561
rect 388154 395325 394918 395561
rect 395154 395325 401918 395561
rect 402154 395325 408918 395561
rect 409154 395325 415918 395561
rect 416154 395325 422918 395561
rect 423154 395325 429918 395561
rect 430154 395325 436918 395561
rect 437154 395325 443918 395561
rect 444154 395325 450918 395561
rect 451154 395325 457918 395561
rect 458154 395325 464918 395561
rect 465154 395325 471918 395561
rect 472154 395325 478918 395561
rect 479154 395325 485918 395561
rect 486154 395325 492918 395561
rect 493154 395325 499918 395561
rect 500154 395325 506918 395561
rect 507154 395325 513918 395561
rect 514154 395325 520918 395561
rect 521154 395325 527918 395561
rect 528154 395325 534918 395561
rect 535154 395325 541918 395561
rect 542154 395325 548918 395561
rect 549154 395325 555918 395561
rect 556154 395325 562918 395561
rect 563154 395325 569918 395561
rect 570154 395325 576918 395561
rect 577154 395325 587570 395561
rect 587806 395325 587890 395561
rect 588126 395325 588210 395561
rect 588446 395325 588530 395561
rect 588766 395325 588874 395561
rect -4950 395283 588874 395325
rect -4950 394494 588874 394536
rect -4950 394258 -3090 394494
rect -2854 394258 -2770 394494
rect -2534 394258 -2450 394494
rect -2214 394258 -2130 394494
rect -1894 394258 1186 394494
rect 1422 394258 8186 394494
rect 8422 394258 15186 394494
rect 15422 394258 22186 394494
rect 22422 394258 29186 394494
rect 29422 394258 36186 394494
rect 36422 394258 43186 394494
rect 43422 394258 50186 394494
rect 50422 394258 57186 394494
rect 57422 394258 64186 394494
rect 64422 394258 71186 394494
rect 71422 394258 78186 394494
rect 78422 394258 85186 394494
rect 85422 394258 92186 394494
rect 92422 394258 99186 394494
rect 99422 394258 106186 394494
rect 106422 394258 113186 394494
rect 113422 394258 120186 394494
rect 120422 394258 127186 394494
rect 127422 394258 134186 394494
rect 134422 394258 141186 394494
rect 141422 394258 148186 394494
rect 148422 394258 155186 394494
rect 155422 394258 162186 394494
rect 162422 394258 169186 394494
rect 169422 394258 176186 394494
rect 176422 394258 183186 394494
rect 183422 394258 190186 394494
rect 190422 394258 197186 394494
rect 197422 394258 204186 394494
rect 204422 394258 211186 394494
rect 211422 394258 218186 394494
rect 218422 394258 225186 394494
rect 225422 394258 232186 394494
rect 232422 394258 239186 394494
rect 239422 394258 246186 394494
rect 246422 394258 253186 394494
rect 253422 394258 260186 394494
rect 260422 394258 267186 394494
rect 267422 394258 274186 394494
rect 274422 394258 281186 394494
rect 281422 394258 288186 394494
rect 288422 394258 295186 394494
rect 295422 394258 302186 394494
rect 302422 394258 309186 394494
rect 309422 394258 316186 394494
rect 316422 394258 323186 394494
rect 323422 394258 330186 394494
rect 330422 394258 337186 394494
rect 337422 394258 344186 394494
rect 344422 394258 351186 394494
rect 351422 394258 358186 394494
rect 358422 394258 365186 394494
rect 365422 394258 372186 394494
rect 372422 394258 379186 394494
rect 379422 394258 386186 394494
rect 386422 394258 393186 394494
rect 393422 394258 400186 394494
rect 400422 394258 407186 394494
rect 407422 394258 414186 394494
rect 414422 394258 421186 394494
rect 421422 394258 428186 394494
rect 428422 394258 435186 394494
rect 435422 394258 442186 394494
rect 442422 394258 449186 394494
rect 449422 394258 456186 394494
rect 456422 394258 463186 394494
rect 463422 394258 470186 394494
rect 470422 394258 477186 394494
rect 477422 394258 484186 394494
rect 484422 394258 491186 394494
rect 491422 394258 498186 394494
rect 498422 394258 505186 394494
rect 505422 394258 512186 394494
rect 512422 394258 519186 394494
rect 519422 394258 526186 394494
rect 526422 394258 533186 394494
rect 533422 394258 540186 394494
rect 540422 394258 547186 394494
rect 547422 394258 554186 394494
rect 554422 394258 561186 394494
rect 561422 394258 568186 394494
rect 568422 394258 575186 394494
rect 575422 394258 582186 394494
rect 582422 394258 585818 394494
rect 586054 394258 586138 394494
rect 586374 394258 586458 394494
rect 586694 394258 586778 394494
rect 587014 394258 588874 394494
rect -4950 394216 588874 394258
rect -4950 388561 588874 388603
rect -4950 388325 -4842 388561
rect -4606 388325 -4522 388561
rect -4286 388325 -4202 388561
rect -3966 388325 -3882 388561
rect -3646 388325 2918 388561
rect 3154 388325 9918 388561
rect 10154 388325 16918 388561
rect 17154 388325 23918 388561
rect 24154 388325 30918 388561
rect 31154 388325 37918 388561
rect 38154 388325 44918 388561
rect 45154 388325 51918 388561
rect 52154 388325 58918 388561
rect 59154 388325 65918 388561
rect 66154 388325 72918 388561
rect 73154 388325 79918 388561
rect 80154 388325 86918 388561
rect 87154 388325 93918 388561
rect 94154 388325 100918 388561
rect 101154 388325 107918 388561
rect 108154 388325 114918 388561
rect 115154 388325 121918 388561
rect 122154 388325 128918 388561
rect 129154 388325 135918 388561
rect 136154 388325 142918 388561
rect 143154 388325 149918 388561
rect 150154 388325 156918 388561
rect 157154 388325 163918 388561
rect 164154 388325 170918 388561
rect 171154 388325 177918 388561
rect 178154 388325 184918 388561
rect 185154 388325 191918 388561
rect 192154 388325 198918 388561
rect 199154 388325 205918 388561
rect 206154 388325 212918 388561
rect 213154 388325 219918 388561
rect 220154 388325 226918 388561
rect 227154 388325 233918 388561
rect 234154 388325 240918 388561
rect 241154 388325 247918 388561
rect 248154 388325 254918 388561
rect 255154 388325 261918 388561
rect 262154 388325 268918 388561
rect 269154 388325 275918 388561
rect 276154 388325 282918 388561
rect 283154 388325 289918 388561
rect 290154 388325 296918 388561
rect 297154 388325 303918 388561
rect 304154 388325 310918 388561
rect 311154 388325 317918 388561
rect 318154 388325 324918 388561
rect 325154 388325 331918 388561
rect 332154 388325 338918 388561
rect 339154 388325 345918 388561
rect 346154 388325 352918 388561
rect 353154 388325 359918 388561
rect 360154 388325 366918 388561
rect 367154 388325 373918 388561
rect 374154 388325 380918 388561
rect 381154 388325 387918 388561
rect 388154 388325 394918 388561
rect 395154 388325 401918 388561
rect 402154 388325 408918 388561
rect 409154 388325 415918 388561
rect 416154 388325 422918 388561
rect 423154 388325 429918 388561
rect 430154 388325 436918 388561
rect 437154 388325 443918 388561
rect 444154 388325 450918 388561
rect 451154 388325 457918 388561
rect 458154 388325 464918 388561
rect 465154 388325 471918 388561
rect 472154 388325 478918 388561
rect 479154 388325 485918 388561
rect 486154 388325 492918 388561
rect 493154 388325 499918 388561
rect 500154 388325 506918 388561
rect 507154 388325 513918 388561
rect 514154 388325 520918 388561
rect 521154 388325 527918 388561
rect 528154 388325 534918 388561
rect 535154 388325 541918 388561
rect 542154 388325 548918 388561
rect 549154 388325 555918 388561
rect 556154 388325 562918 388561
rect 563154 388325 569918 388561
rect 570154 388325 576918 388561
rect 577154 388325 587570 388561
rect 587806 388325 587890 388561
rect 588126 388325 588210 388561
rect 588446 388325 588530 388561
rect 588766 388325 588874 388561
rect -4950 388283 588874 388325
rect -4950 387494 588874 387536
rect -4950 387258 -3090 387494
rect -2854 387258 -2770 387494
rect -2534 387258 -2450 387494
rect -2214 387258 -2130 387494
rect -1894 387258 1186 387494
rect 1422 387258 8186 387494
rect 8422 387258 15186 387494
rect 15422 387258 22186 387494
rect 22422 387258 29186 387494
rect 29422 387258 36186 387494
rect 36422 387258 43186 387494
rect 43422 387258 50186 387494
rect 50422 387258 57186 387494
rect 57422 387258 64186 387494
rect 64422 387258 71186 387494
rect 71422 387258 78186 387494
rect 78422 387258 85186 387494
rect 85422 387258 92186 387494
rect 92422 387258 99186 387494
rect 99422 387258 106186 387494
rect 106422 387258 113186 387494
rect 113422 387258 120186 387494
rect 120422 387258 127186 387494
rect 127422 387258 134186 387494
rect 134422 387258 141186 387494
rect 141422 387258 148186 387494
rect 148422 387258 155186 387494
rect 155422 387258 162186 387494
rect 162422 387258 169186 387494
rect 169422 387258 176186 387494
rect 176422 387258 183186 387494
rect 183422 387258 190186 387494
rect 190422 387258 197186 387494
rect 197422 387258 204186 387494
rect 204422 387258 211186 387494
rect 211422 387258 218186 387494
rect 218422 387258 225186 387494
rect 225422 387258 232186 387494
rect 232422 387258 239186 387494
rect 239422 387258 246186 387494
rect 246422 387258 253186 387494
rect 253422 387258 260186 387494
rect 260422 387258 267186 387494
rect 267422 387258 274186 387494
rect 274422 387258 281186 387494
rect 281422 387258 288186 387494
rect 288422 387258 295186 387494
rect 295422 387258 302186 387494
rect 302422 387258 309186 387494
rect 309422 387258 316186 387494
rect 316422 387258 323186 387494
rect 323422 387258 330186 387494
rect 330422 387258 337186 387494
rect 337422 387258 344186 387494
rect 344422 387258 351186 387494
rect 351422 387258 358186 387494
rect 358422 387258 365186 387494
rect 365422 387258 372186 387494
rect 372422 387258 379186 387494
rect 379422 387258 386186 387494
rect 386422 387258 393186 387494
rect 393422 387258 400186 387494
rect 400422 387258 407186 387494
rect 407422 387258 414186 387494
rect 414422 387258 421186 387494
rect 421422 387258 428186 387494
rect 428422 387258 435186 387494
rect 435422 387258 442186 387494
rect 442422 387258 449186 387494
rect 449422 387258 456186 387494
rect 456422 387258 463186 387494
rect 463422 387258 470186 387494
rect 470422 387258 477186 387494
rect 477422 387258 484186 387494
rect 484422 387258 491186 387494
rect 491422 387258 498186 387494
rect 498422 387258 505186 387494
rect 505422 387258 512186 387494
rect 512422 387258 519186 387494
rect 519422 387258 526186 387494
rect 526422 387258 533186 387494
rect 533422 387258 540186 387494
rect 540422 387258 547186 387494
rect 547422 387258 554186 387494
rect 554422 387258 561186 387494
rect 561422 387258 568186 387494
rect 568422 387258 575186 387494
rect 575422 387258 582186 387494
rect 582422 387258 585818 387494
rect 586054 387258 586138 387494
rect 586374 387258 586458 387494
rect 586694 387258 586778 387494
rect 587014 387258 588874 387494
rect -4950 387216 588874 387258
rect -4950 381561 588874 381603
rect -4950 381325 -4842 381561
rect -4606 381325 -4522 381561
rect -4286 381325 -4202 381561
rect -3966 381325 -3882 381561
rect -3646 381325 2918 381561
rect 3154 381325 9918 381561
rect 10154 381325 16918 381561
rect 17154 381325 23918 381561
rect 24154 381325 30918 381561
rect 31154 381325 37918 381561
rect 38154 381325 44918 381561
rect 45154 381325 51918 381561
rect 52154 381325 58918 381561
rect 59154 381325 65918 381561
rect 66154 381325 72918 381561
rect 73154 381325 79918 381561
rect 80154 381325 86918 381561
rect 87154 381325 93918 381561
rect 94154 381325 100918 381561
rect 101154 381325 107918 381561
rect 108154 381325 114918 381561
rect 115154 381325 121918 381561
rect 122154 381325 128918 381561
rect 129154 381325 135918 381561
rect 136154 381325 142918 381561
rect 143154 381325 149918 381561
rect 150154 381325 156918 381561
rect 157154 381325 163918 381561
rect 164154 381325 170918 381561
rect 171154 381325 177918 381561
rect 178154 381325 184918 381561
rect 185154 381325 191918 381561
rect 192154 381325 198918 381561
rect 199154 381325 205918 381561
rect 206154 381325 212918 381561
rect 213154 381325 219918 381561
rect 220154 381325 226918 381561
rect 227154 381325 233918 381561
rect 234154 381325 240918 381561
rect 241154 381325 247918 381561
rect 248154 381325 254918 381561
rect 255154 381325 261918 381561
rect 262154 381325 268918 381561
rect 269154 381325 275918 381561
rect 276154 381325 282918 381561
rect 283154 381325 289918 381561
rect 290154 381325 296918 381561
rect 297154 381325 303918 381561
rect 304154 381325 310918 381561
rect 311154 381325 317918 381561
rect 318154 381325 324918 381561
rect 325154 381325 331918 381561
rect 332154 381325 338918 381561
rect 339154 381325 345918 381561
rect 346154 381325 352918 381561
rect 353154 381325 359918 381561
rect 360154 381325 366918 381561
rect 367154 381325 373918 381561
rect 374154 381325 380918 381561
rect 381154 381325 387918 381561
rect 388154 381325 394918 381561
rect 395154 381325 401918 381561
rect 402154 381325 408918 381561
rect 409154 381325 415918 381561
rect 416154 381325 422918 381561
rect 423154 381325 429918 381561
rect 430154 381325 436918 381561
rect 437154 381325 443918 381561
rect 444154 381325 450918 381561
rect 451154 381325 457918 381561
rect 458154 381325 464918 381561
rect 465154 381325 471918 381561
rect 472154 381325 478918 381561
rect 479154 381325 485918 381561
rect 486154 381325 492918 381561
rect 493154 381325 499918 381561
rect 500154 381325 506918 381561
rect 507154 381325 513918 381561
rect 514154 381325 527918 381561
rect 528154 381325 534918 381561
rect 535154 381325 541918 381561
rect 542154 381325 548918 381561
rect 549154 381325 555918 381561
rect 556154 381325 562918 381561
rect 563154 381325 569918 381561
rect 570154 381325 576918 381561
rect 577154 381325 587570 381561
rect 587806 381325 587890 381561
rect 588126 381325 588210 381561
rect 588446 381325 588530 381561
rect 588766 381325 588874 381561
rect -4950 381283 588874 381325
rect -4950 380494 588874 380536
rect -4950 380258 -3090 380494
rect -2854 380258 -2770 380494
rect -2534 380258 -2450 380494
rect -2214 380258 -2130 380494
rect -1894 380258 1186 380494
rect 1422 380258 8186 380494
rect 8422 380258 15186 380494
rect 15422 380258 22186 380494
rect 22422 380258 29186 380494
rect 29422 380258 36186 380494
rect 36422 380258 43186 380494
rect 43422 380258 50186 380494
rect 50422 380258 57186 380494
rect 57422 380258 64186 380494
rect 64422 380258 71186 380494
rect 71422 380258 78186 380494
rect 78422 380258 85186 380494
rect 85422 380258 92186 380494
rect 92422 380258 99186 380494
rect 99422 380258 106186 380494
rect 106422 380258 113186 380494
rect 113422 380258 120186 380494
rect 120422 380258 127186 380494
rect 127422 380258 134186 380494
rect 134422 380258 141186 380494
rect 141422 380258 148186 380494
rect 148422 380258 155186 380494
rect 155422 380258 162186 380494
rect 162422 380258 169186 380494
rect 169422 380258 176186 380494
rect 176422 380258 183186 380494
rect 183422 380258 190186 380494
rect 190422 380258 197186 380494
rect 197422 380258 204186 380494
rect 204422 380258 211186 380494
rect 211422 380258 218186 380494
rect 218422 380258 225186 380494
rect 225422 380258 232186 380494
rect 232422 380258 239186 380494
rect 239422 380258 246186 380494
rect 246422 380258 253186 380494
rect 253422 380258 260186 380494
rect 260422 380258 267186 380494
rect 267422 380258 274186 380494
rect 274422 380258 281186 380494
rect 281422 380258 288186 380494
rect 288422 380258 295186 380494
rect 295422 380258 302186 380494
rect 302422 380258 309186 380494
rect 309422 380258 316186 380494
rect 316422 380258 323186 380494
rect 323422 380258 330186 380494
rect 330422 380258 337186 380494
rect 337422 380258 344186 380494
rect 344422 380258 351186 380494
rect 351422 380258 358186 380494
rect 358422 380258 365186 380494
rect 365422 380258 372186 380494
rect 372422 380258 379186 380494
rect 379422 380258 386186 380494
rect 386422 380258 393186 380494
rect 393422 380258 400186 380494
rect 400422 380258 407186 380494
rect 407422 380258 414186 380494
rect 414422 380258 421186 380494
rect 421422 380258 428186 380494
rect 428422 380258 435186 380494
rect 435422 380258 442186 380494
rect 442422 380258 449186 380494
rect 449422 380258 456186 380494
rect 456422 380258 463186 380494
rect 463422 380258 470186 380494
rect 470422 380258 477186 380494
rect 477422 380258 484186 380494
rect 484422 380258 491186 380494
rect 491422 380258 498186 380494
rect 498422 380258 505186 380494
rect 505422 380258 512186 380494
rect 512422 380258 519186 380494
rect 519422 380258 533186 380494
rect 533422 380258 540186 380494
rect 540422 380258 547186 380494
rect 547422 380258 554186 380494
rect 554422 380258 561186 380494
rect 561422 380258 568186 380494
rect 568422 380258 575186 380494
rect 575422 380258 582186 380494
rect 582422 380258 585818 380494
rect 586054 380258 586138 380494
rect 586374 380258 586458 380494
rect 586694 380258 586778 380494
rect 587014 380258 588874 380494
rect -4950 380216 588874 380258
rect -4950 374561 588874 374603
rect -4950 374325 -4842 374561
rect -4606 374325 -4522 374561
rect -4286 374325 -4202 374561
rect -3966 374325 -3882 374561
rect -3646 374325 2918 374561
rect 3154 374325 9918 374561
rect 10154 374325 16918 374561
rect 17154 374325 23918 374561
rect 24154 374325 30918 374561
rect 31154 374325 37918 374561
rect 38154 374325 44918 374561
rect 45154 374325 51918 374561
rect 52154 374325 58918 374561
rect 59154 374325 65918 374561
rect 66154 374325 72918 374561
rect 73154 374325 79918 374561
rect 80154 374325 86918 374561
rect 87154 374325 93918 374561
rect 94154 374325 100918 374561
rect 101154 374325 107918 374561
rect 108154 374325 114918 374561
rect 115154 374325 121918 374561
rect 122154 374325 128918 374561
rect 129154 374325 135918 374561
rect 136154 374325 142918 374561
rect 143154 374325 149918 374561
rect 150154 374325 156918 374561
rect 157154 374325 163918 374561
rect 164154 374325 170918 374561
rect 171154 374325 177918 374561
rect 178154 374325 184918 374561
rect 185154 374325 191918 374561
rect 192154 374325 198918 374561
rect 199154 374325 205918 374561
rect 206154 374325 212918 374561
rect 213154 374325 219918 374561
rect 220154 374325 226918 374561
rect 227154 374325 233918 374561
rect 234154 374325 240918 374561
rect 241154 374325 247918 374561
rect 248154 374325 254918 374561
rect 255154 374325 261918 374561
rect 262154 374325 268918 374561
rect 269154 374325 275918 374561
rect 276154 374325 282918 374561
rect 283154 374325 289918 374561
rect 290154 374325 296918 374561
rect 297154 374325 303918 374561
rect 304154 374325 310918 374561
rect 311154 374325 317918 374561
rect 318154 374325 324918 374561
rect 325154 374325 331918 374561
rect 332154 374325 338918 374561
rect 339154 374325 345918 374561
rect 346154 374325 352918 374561
rect 353154 374325 359918 374561
rect 360154 374325 366918 374561
rect 367154 374325 373918 374561
rect 374154 374325 380918 374561
rect 381154 374325 387918 374561
rect 388154 374325 394918 374561
rect 395154 374325 401918 374561
rect 402154 374325 408918 374561
rect 409154 374325 415918 374561
rect 416154 374325 422918 374561
rect 423154 374325 429918 374561
rect 430154 374325 436918 374561
rect 437154 374325 443918 374561
rect 444154 374325 450918 374561
rect 451154 374325 457918 374561
rect 458154 374325 464918 374561
rect 465154 374325 471918 374561
rect 472154 374325 478918 374561
rect 479154 374325 485918 374561
rect 486154 374325 492918 374561
rect 493154 374325 499918 374561
rect 500154 374325 506918 374561
rect 507154 374325 513918 374561
rect 514154 374325 520918 374561
rect 521154 374325 522850 374561
rect 523086 374325 524782 374561
rect 525018 374325 526714 374561
rect 526950 374325 527918 374561
rect 528154 374325 534918 374561
rect 535154 374325 541918 374561
rect 542154 374325 548918 374561
rect 549154 374325 555918 374561
rect 556154 374325 562918 374561
rect 563154 374325 569918 374561
rect 570154 374325 576918 374561
rect 577154 374325 587570 374561
rect 587806 374325 587890 374561
rect 588126 374325 588210 374561
rect 588446 374325 588530 374561
rect 588766 374325 588874 374561
rect -4950 374283 588874 374325
rect -4950 373494 588874 373536
rect -4950 373258 -3090 373494
rect -2854 373258 -2770 373494
rect -2534 373258 -2450 373494
rect -2214 373258 -2130 373494
rect -1894 373258 1186 373494
rect 1422 373258 8186 373494
rect 8422 373258 15186 373494
rect 15422 373258 22186 373494
rect 22422 373258 29186 373494
rect 29422 373258 36186 373494
rect 36422 373258 43186 373494
rect 43422 373258 50186 373494
rect 50422 373258 57186 373494
rect 57422 373258 64186 373494
rect 64422 373258 71186 373494
rect 71422 373258 78186 373494
rect 78422 373258 85186 373494
rect 85422 373258 92186 373494
rect 92422 373258 99186 373494
rect 99422 373258 106186 373494
rect 106422 373258 113186 373494
rect 113422 373258 120186 373494
rect 120422 373258 127186 373494
rect 127422 373258 134186 373494
rect 134422 373258 141186 373494
rect 141422 373258 148186 373494
rect 148422 373258 155186 373494
rect 155422 373258 162186 373494
rect 162422 373258 169186 373494
rect 169422 373258 176186 373494
rect 176422 373258 183186 373494
rect 183422 373258 190186 373494
rect 190422 373258 197186 373494
rect 197422 373258 204186 373494
rect 204422 373258 211186 373494
rect 211422 373258 218186 373494
rect 218422 373258 225186 373494
rect 225422 373258 232186 373494
rect 232422 373258 239186 373494
rect 239422 373258 246186 373494
rect 246422 373258 253186 373494
rect 253422 373258 260186 373494
rect 260422 373258 267186 373494
rect 267422 373258 274186 373494
rect 274422 373258 281186 373494
rect 281422 373258 288186 373494
rect 288422 373258 295186 373494
rect 295422 373258 302186 373494
rect 302422 373258 309186 373494
rect 309422 373258 316186 373494
rect 316422 373258 323186 373494
rect 323422 373258 330186 373494
rect 330422 373258 337186 373494
rect 337422 373258 344186 373494
rect 344422 373258 351186 373494
rect 351422 373258 358186 373494
rect 358422 373258 365186 373494
rect 365422 373258 372186 373494
rect 372422 373258 379186 373494
rect 379422 373258 386186 373494
rect 386422 373258 393186 373494
rect 393422 373258 400186 373494
rect 400422 373258 407186 373494
rect 407422 373258 414186 373494
rect 414422 373258 421186 373494
rect 421422 373258 428186 373494
rect 428422 373258 435186 373494
rect 435422 373258 442186 373494
rect 442422 373258 449186 373494
rect 449422 373258 456186 373494
rect 456422 373258 463186 373494
rect 463422 373258 470186 373494
rect 470422 373258 477186 373494
rect 477422 373258 484186 373494
rect 484422 373258 491186 373494
rect 491422 373258 498186 373494
rect 498422 373258 505186 373494
rect 505422 373258 512186 373494
rect 512422 373258 519186 373494
rect 519422 373258 519952 373494
rect 520188 373258 521884 373494
rect 522120 373258 523816 373494
rect 524052 373258 525748 373494
rect 525984 373258 533186 373494
rect 533422 373258 540186 373494
rect 540422 373258 547186 373494
rect 547422 373258 554186 373494
rect 554422 373258 561186 373494
rect 561422 373258 568186 373494
rect 568422 373258 575186 373494
rect 575422 373258 582186 373494
rect 582422 373258 585818 373494
rect 586054 373258 586138 373494
rect 586374 373258 586458 373494
rect 586694 373258 586778 373494
rect 587014 373258 588874 373494
rect -4950 373216 588874 373258
rect -4950 367561 588874 367603
rect -4950 367325 -4842 367561
rect -4606 367325 -4522 367561
rect -4286 367325 -4202 367561
rect -3966 367325 -3882 367561
rect -3646 367325 2918 367561
rect 3154 367325 9918 367561
rect 10154 367325 16918 367561
rect 17154 367325 23918 367561
rect 24154 367325 30918 367561
rect 31154 367325 37918 367561
rect 38154 367325 44918 367561
rect 45154 367325 51918 367561
rect 52154 367325 58918 367561
rect 59154 367325 65918 367561
rect 66154 367325 72918 367561
rect 73154 367325 79918 367561
rect 80154 367325 86918 367561
rect 87154 367325 93918 367561
rect 94154 367325 100918 367561
rect 101154 367325 107918 367561
rect 108154 367325 114918 367561
rect 115154 367325 121918 367561
rect 122154 367325 128918 367561
rect 129154 367325 135918 367561
rect 136154 367325 142918 367561
rect 143154 367325 149918 367561
rect 150154 367325 156918 367561
rect 157154 367325 163918 367561
rect 164154 367325 170918 367561
rect 171154 367325 177918 367561
rect 178154 367325 184918 367561
rect 185154 367325 191918 367561
rect 192154 367325 198918 367561
rect 199154 367325 205918 367561
rect 206154 367325 212918 367561
rect 213154 367325 219918 367561
rect 220154 367325 226918 367561
rect 227154 367325 233918 367561
rect 234154 367325 240918 367561
rect 241154 367325 247918 367561
rect 248154 367325 254918 367561
rect 255154 367325 261918 367561
rect 262154 367325 268918 367561
rect 269154 367325 275918 367561
rect 276154 367325 282918 367561
rect 283154 367325 289918 367561
rect 290154 367325 317918 367561
rect 318154 367325 324918 367561
rect 325154 367325 331918 367561
rect 332154 367325 338918 367561
rect 339154 367325 345918 367561
rect 346154 367325 352918 367561
rect 353154 367325 359918 367561
rect 360154 367325 366918 367561
rect 367154 367325 373918 367561
rect 374154 367325 380918 367561
rect 381154 367325 387918 367561
rect 388154 367325 394918 367561
rect 395154 367325 401918 367561
rect 402154 367325 408918 367561
rect 409154 367325 415918 367561
rect 416154 367325 422918 367561
rect 423154 367325 429918 367561
rect 430154 367325 436918 367561
rect 437154 367325 443918 367561
rect 444154 367325 450918 367561
rect 451154 367325 457918 367561
rect 458154 367325 464918 367561
rect 465154 367325 471918 367561
rect 472154 367325 478918 367561
rect 479154 367325 485918 367561
rect 486154 367325 492918 367561
rect 493154 367325 499918 367561
rect 500154 367325 506918 367561
rect 507154 367325 513918 367561
rect 514154 367325 520918 367561
rect 521154 367325 522850 367561
rect 523086 367325 524782 367561
rect 525018 367325 526714 367561
rect 526950 367325 527918 367561
rect 528154 367325 534918 367561
rect 535154 367325 541918 367561
rect 542154 367325 548918 367561
rect 549154 367325 555918 367561
rect 556154 367325 562918 367561
rect 563154 367325 569918 367561
rect 570154 367325 576918 367561
rect 577154 367325 587570 367561
rect 587806 367325 587890 367561
rect 588126 367325 588210 367561
rect 588446 367325 588530 367561
rect 588766 367325 588874 367561
rect -4950 367283 588874 367325
rect -4950 366494 588874 366536
rect -4950 366258 -3090 366494
rect -2854 366258 -2770 366494
rect -2534 366258 -2450 366494
rect -2214 366258 -2130 366494
rect -1894 366258 1186 366494
rect 1422 366258 8186 366494
rect 8422 366258 15186 366494
rect 15422 366258 22186 366494
rect 22422 366258 29186 366494
rect 29422 366258 36186 366494
rect 36422 366258 43186 366494
rect 43422 366258 50186 366494
rect 50422 366258 57186 366494
rect 57422 366258 64186 366494
rect 64422 366258 71186 366494
rect 71422 366258 78186 366494
rect 78422 366258 85186 366494
rect 85422 366258 92186 366494
rect 92422 366258 99186 366494
rect 99422 366258 106186 366494
rect 106422 366258 113186 366494
rect 113422 366258 120186 366494
rect 120422 366258 127186 366494
rect 127422 366258 134186 366494
rect 134422 366258 141186 366494
rect 141422 366258 148186 366494
rect 148422 366258 155186 366494
rect 155422 366258 162186 366494
rect 162422 366258 169186 366494
rect 169422 366258 176186 366494
rect 176422 366258 183186 366494
rect 183422 366258 190186 366494
rect 190422 366258 197186 366494
rect 197422 366258 204186 366494
rect 204422 366258 211186 366494
rect 211422 366258 218186 366494
rect 218422 366258 225186 366494
rect 225422 366258 232186 366494
rect 232422 366258 239186 366494
rect 239422 366258 246186 366494
rect 246422 366258 253186 366494
rect 253422 366258 260186 366494
rect 260422 366258 267186 366494
rect 267422 366258 274186 366494
rect 274422 366258 281186 366494
rect 281422 366258 288186 366494
rect 288422 366258 316186 366494
rect 316422 366258 323186 366494
rect 323422 366258 330186 366494
rect 330422 366258 337186 366494
rect 337422 366258 344186 366494
rect 344422 366258 351186 366494
rect 351422 366258 358186 366494
rect 358422 366258 365186 366494
rect 365422 366258 372186 366494
rect 372422 366258 379186 366494
rect 379422 366258 386186 366494
rect 386422 366258 393186 366494
rect 393422 366258 400186 366494
rect 400422 366258 407186 366494
rect 407422 366258 414186 366494
rect 414422 366258 421186 366494
rect 421422 366258 428186 366494
rect 428422 366258 435186 366494
rect 435422 366258 442186 366494
rect 442422 366258 449186 366494
rect 449422 366258 456186 366494
rect 456422 366258 463186 366494
rect 463422 366258 470186 366494
rect 470422 366258 477186 366494
rect 477422 366258 484186 366494
rect 484422 366258 491186 366494
rect 491422 366258 498186 366494
rect 498422 366258 505186 366494
rect 505422 366258 512186 366494
rect 512422 366258 519186 366494
rect 519422 366258 519952 366494
rect 520188 366258 521884 366494
rect 522120 366258 523816 366494
rect 524052 366258 525748 366494
rect 525984 366258 533186 366494
rect 533422 366258 540186 366494
rect 540422 366258 547186 366494
rect 547422 366258 554186 366494
rect 554422 366258 561186 366494
rect 561422 366258 568186 366494
rect 568422 366258 575186 366494
rect 575422 366258 582186 366494
rect 582422 366258 585818 366494
rect 586054 366258 586138 366494
rect 586374 366258 586458 366494
rect 586694 366258 586778 366494
rect 587014 366258 588874 366494
rect -4950 366216 588874 366258
rect -4950 360561 588874 360603
rect -4950 360325 -4842 360561
rect -4606 360325 -4522 360561
rect -4286 360325 -4202 360561
rect -3966 360325 -3882 360561
rect -3646 360325 2918 360561
rect 3154 360325 9918 360561
rect 10154 360325 16918 360561
rect 17154 360325 23918 360561
rect 24154 360325 30918 360561
rect 31154 360325 37918 360561
rect 38154 360325 44918 360561
rect 45154 360325 51918 360561
rect 52154 360325 58918 360561
rect 59154 360325 65918 360561
rect 66154 360325 72918 360561
rect 73154 360325 79918 360561
rect 80154 360325 86918 360561
rect 87154 360325 93918 360561
rect 94154 360325 100918 360561
rect 101154 360325 107918 360561
rect 108154 360325 114918 360561
rect 115154 360325 121918 360561
rect 122154 360325 128918 360561
rect 129154 360325 135918 360561
rect 136154 360325 142918 360561
rect 143154 360325 149918 360561
rect 150154 360325 156918 360561
rect 157154 360325 163918 360561
rect 164154 360325 170918 360561
rect 171154 360325 177918 360561
rect 178154 360325 184918 360561
rect 185154 360325 191918 360561
rect 192154 360325 198918 360561
rect 199154 360325 205918 360561
rect 206154 360325 212918 360561
rect 213154 360325 219918 360561
rect 220154 360325 226918 360561
rect 227154 360325 233918 360561
rect 234154 360325 240918 360561
rect 241154 360325 247918 360561
rect 248154 360325 254918 360561
rect 255154 360325 261918 360561
rect 262154 360325 268918 360561
rect 269154 360325 275918 360561
rect 276154 360325 282918 360561
rect 283154 360325 289918 360561
rect 290154 360325 296918 360561
rect 297154 360325 303918 360561
rect 304154 360325 310918 360561
rect 311154 360325 317918 360561
rect 318154 360325 324918 360561
rect 325154 360325 331918 360561
rect 332154 360325 338918 360561
rect 339154 360325 345918 360561
rect 346154 360325 352918 360561
rect 353154 360325 359918 360561
rect 360154 360325 366918 360561
rect 367154 360325 373918 360561
rect 374154 360325 380918 360561
rect 381154 360325 387918 360561
rect 388154 360325 394918 360561
rect 395154 360325 401918 360561
rect 402154 360325 408918 360561
rect 409154 360325 415918 360561
rect 416154 360325 422918 360561
rect 423154 360325 429918 360561
rect 430154 360325 436918 360561
rect 437154 360325 443918 360561
rect 444154 360325 450918 360561
rect 451154 360325 457918 360561
rect 458154 360325 464918 360561
rect 465154 360325 471918 360561
rect 472154 360325 478918 360561
rect 479154 360325 485918 360561
rect 486154 360325 492918 360561
rect 493154 360325 499918 360561
rect 500154 360325 506918 360561
rect 507154 360325 513918 360561
rect 514154 360325 527918 360561
rect 528154 360325 534918 360561
rect 535154 360325 541918 360561
rect 542154 360325 548918 360561
rect 549154 360325 555918 360561
rect 556154 360325 562918 360561
rect 563154 360325 569918 360561
rect 570154 360325 576918 360561
rect 577154 360325 587570 360561
rect 587806 360325 587890 360561
rect 588126 360325 588210 360561
rect 588446 360325 588530 360561
rect 588766 360325 588874 360561
rect -4950 360283 588874 360325
rect -4950 359494 588874 359536
rect -4950 359258 -3090 359494
rect -2854 359258 -2770 359494
rect -2534 359258 -2450 359494
rect -2214 359258 -2130 359494
rect -1894 359258 1186 359494
rect 1422 359258 8186 359494
rect 8422 359258 15186 359494
rect 15422 359258 22186 359494
rect 22422 359258 29186 359494
rect 29422 359258 36186 359494
rect 36422 359258 43186 359494
rect 43422 359258 50186 359494
rect 50422 359258 57186 359494
rect 57422 359258 64186 359494
rect 64422 359258 71186 359494
rect 71422 359258 78186 359494
rect 78422 359258 85186 359494
rect 85422 359258 92186 359494
rect 92422 359258 99186 359494
rect 99422 359258 106186 359494
rect 106422 359258 113186 359494
rect 113422 359258 120186 359494
rect 120422 359258 127186 359494
rect 127422 359258 134186 359494
rect 134422 359258 141186 359494
rect 141422 359258 148186 359494
rect 148422 359258 155186 359494
rect 155422 359258 162186 359494
rect 162422 359258 169186 359494
rect 169422 359258 176186 359494
rect 176422 359258 183186 359494
rect 183422 359258 190186 359494
rect 190422 359258 197186 359494
rect 197422 359258 204186 359494
rect 204422 359258 211186 359494
rect 211422 359258 218186 359494
rect 218422 359258 225186 359494
rect 225422 359258 232186 359494
rect 232422 359258 239186 359494
rect 239422 359258 246186 359494
rect 246422 359258 253186 359494
rect 253422 359258 260186 359494
rect 260422 359258 267186 359494
rect 267422 359258 274186 359494
rect 274422 359258 281186 359494
rect 281422 359258 288186 359494
rect 288422 359258 295186 359494
rect 295422 359258 302186 359494
rect 302422 359258 309186 359494
rect 309422 359258 316186 359494
rect 316422 359258 323186 359494
rect 323422 359258 330186 359494
rect 330422 359258 337186 359494
rect 337422 359258 344186 359494
rect 344422 359258 351186 359494
rect 351422 359258 358186 359494
rect 358422 359258 365186 359494
rect 365422 359258 372186 359494
rect 372422 359258 379186 359494
rect 379422 359258 386186 359494
rect 386422 359258 393186 359494
rect 393422 359258 400186 359494
rect 400422 359258 407186 359494
rect 407422 359258 414186 359494
rect 414422 359258 421186 359494
rect 421422 359258 428186 359494
rect 428422 359258 435186 359494
rect 435422 359258 442186 359494
rect 442422 359258 449186 359494
rect 449422 359258 456186 359494
rect 456422 359258 463186 359494
rect 463422 359258 470186 359494
rect 470422 359258 477186 359494
rect 477422 359258 484186 359494
rect 484422 359258 491186 359494
rect 491422 359258 498186 359494
rect 498422 359258 505186 359494
rect 505422 359258 512186 359494
rect 512422 359258 519186 359494
rect 519422 359258 526186 359494
rect 526422 359258 533186 359494
rect 533422 359258 540186 359494
rect 540422 359258 547186 359494
rect 547422 359258 554186 359494
rect 554422 359258 561186 359494
rect 561422 359258 568186 359494
rect 568422 359258 575186 359494
rect 575422 359258 582186 359494
rect 582422 359258 585818 359494
rect 586054 359258 586138 359494
rect 586374 359258 586458 359494
rect 586694 359258 586778 359494
rect 587014 359258 588874 359494
rect -4950 359216 588874 359258
rect -4950 353561 588874 353603
rect -4950 353325 -4842 353561
rect -4606 353325 -4522 353561
rect -4286 353325 -4202 353561
rect -3966 353325 -3882 353561
rect -3646 353325 2918 353561
rect 3154 353325 9918 353561
rect 10154 353325 16918 353561
rect 17154 353325 23918 353561
rect 24154 353325 30918 353561
rect 31154 353325 37918 353561
rect 38154 353325 44918 353561
rect 45154 353325 51918 353561
rect 52154 353325 58918 353561
rect 59154 353325 65918 353561
rect 66154 353325 72918 353561
rect 73154 353325 79918 353561
rect 80154 353325 86918 353561
rect 87154 353325 93918 353561
rect 94154 353325 100918 353561
rect 101154 353325 107918 353561
rect 108154 353325 114918 353561
rect 115154 353325 121918 353561
rect 122154 353325 128918 353561
rect 129154 353325 135918 353561
rect 136154 353325 142918 353561
rect 143154 353325 149918 353561
rect 150154 353325 156918 353561
rect 157154 353325 163918 353561
rect 164154 353325 170918 353561
rect 171154 353325 177918 353561
rect 178154 353325 184918 353561
rect 185154 353325 191918 353561
rect 192154 353325 198918 353561
rect 199154 353325 205918 353561
rect 206154 353325 212918 353561
rect 213154 353325 219918 353561
rect 220154 353325 226918 353561
rect 227154 353325 233918 353561
rect 234154 353325 240918 353561
rect 241154 353325 247918 353561
rect 248154 353325 254918 353561
rect 255154 353325 261918 353561
rect 262154 353325 268918 353561
rect 269154 353325 275918 353561
rect 276154 353325 282918 353561
rect 283154 353325 289918 353561
rect 290154 353325 296918 353561
rect 297154 353325 303918 353561
rect 304154 353325 310918 353561
rect 311154 353325 317918 353561
rect 318154 353325 324918 353561
rect 325154 353325 331918 353561
rect 332154 353325 338918 353561
rect 339154 353325 345918 353561
rect 346154 353325 352918 353561
rect 353154 353325 359918 353561
rect 360154 353325 366918 353561
rect 367154 353325 373918 353561
rect 374154 353325 380918 353561
rect 381154 353325 387918 353561
rect 388154 353325 394918 353561
rect 395154 353325 401918 353561
rect 402154 353325 408918 353561
rect 409154 353325 415918 353561
rect 416154 353325 422918 353561
rect 423154 353325 429918 353561
rect 430154 353325 436918 353561
rect 437154 353325 443918 353561
rect 444154 353325 450918 353561
rect 451154 353325 457918 353561
rect 458154 353325 464918 353561
rect 465154 353325 471918 353561
rect 472154 353325 478918 353561
rect 479154 353325 485918 353561
rect 486154 353325 492918 353561
rect 493154 353325 499918 353561
rect 500154 353325 506918 353561
rect 507154 353325 513918 353561
rect 514154 353325 520918 353561
rect 521154 353325 527918 353561
rect 528154 353325 534918 353561
rect 535154 353325 541918 353561
rect 542154 353325 548918 353561
rect 549154 353325 555918 353561
rect 556154 353325 562918 353561
rect 563154 353325 569918 353561
rect 570154 353325 576918 353561
rect 577154 353325 587570 353561
rect 587806 353325 587890 353561
rect 588126 353325 588210 353561
rect 588446 353325 588530 353561
rect 588766 353325 588874 353561
rect -4950 353283 588874 353325
rect -4950 352494 588874 352536
rect -4950 352258 -3090 352494
rect -2854 352258 -2770 352494
rect -2534 352258 -2450 352494
rect -2214 352258 -2130 352494
rect -1894 352258 1186 352494
rect 1422 352258 8186 352494
rect 8422 352258 15186 352494
rect 15422 352258 22186 352494
rect 22422 352258 29186 352494
rect 29422 352258 36186 352494
rect 36422 352258 43186 352494
rect 43422 352258 50186 352494
rect 50422 352258 57186 352494
rect 57422 352258 64186 352494
rect 64422 352258 71186 352494
rect 71422 352258 78186 352494
rect 78422 352258 85186 352494
rect 85422 352258 92186 352494
rect 92422 352258 99186 352494
rect 99422 352258 106186 352494
rect 106422 352258 113186 352494
rect 113422 352258 120186 352494
rect 120422 352258 127186 352494
rect 127422 352258 134186 352494
rect 134422 352258 141186 352494
rect 141422 352258 148186 352494
rect 148422 352258 155186 352494
rect 155422 352258 162186 352494
rect 162422 352258 169186 352494
rect 169422 352258 176186 352494
rect 176422 352258 183186 352494
rect 183422 352258 190186 352494
rect 190422 352258 197186 352494
rect 197422 352258 204186 352494
rect 204422 352258 211186 352494
rect 211422 352258 218186 352494
rect 218422 352258 225186 352494
rect 225422 352258 232186 352494
rect 232422 352258 239186 352494
rect 239422 352258 246186 352494
rect 246422 352258 253186 352494
rect 253422 352258 260186 352494
rect 260422 352258 267186 352494
rect 267422 352258 274186 352494
rect 274422 352258 281186 352494
rect 281422 352258 288186 352494
rect 288422 352258 295186 352494
rect 295422 352258 302186 352494
rect 302422 352258 309186 352494
rect 309422 352258 316186 352494
rect 316422 352258 323186 352494
rect 323422 352258 330186 352494
rect 330422 352258 337186 352494
rect 337422 352258 344186 352494
rect 344422 352258 351186 352494
rect 351422 352258 358186 352494
rect 358422 352258 365186 352494
rect 365422 352258 372186 352494
rect 372422 352258 379186 352494
rect 379422 352258 386186 352494
rect 386422 352258 393186 352494
rect 393422 352258 400186 352494
rect 400422 352258 407186 352494
rect 407422 352258 414186 352494
rect 414422 352258 421186 352494
rect 421422 352258 428186 352494
rect 428422 352258 435186 352494
rect 435422 352258 442186 352494
rect 442422 352258 449186 352494
rect 449422 352258 456186 352494
rect 456422 352258 463186 352494
rect 463422 352258 470186 352494
rect 470422 352258 477186 352494
rect 477422 352258 484186 352494
rect 484422 352258 491186 352494
rect 491422 352258 498186 352494
rect 498422 352258 505186 352494
rect 505422 352258 512186 352494
rect 512422 352258 519186 352494
rect 519422 352258 526186 352494
rect 526422 352258 533186 352494
rect 533422 352258 540186 352494
rect 540422 352258 547186 352494
rect 547422 352258 554186 352494
rect 554422 352258 561186 352494
rect 561422 352258 568186 352494
rect 568422 352258 575186 352494
rect 575422 352258 582186 352494
rect 582422 352258 585818 352494
rect 586054 352258 586138 352494
rect 586374 352258 586458 352494
rect 586694 352258 586778 352494
rect 587014 352258 588874 352494
rect -4950 352216 588874 352258
rect -4950 346561 588874 346603
rect -4950 346325 -4842 346561
rect -4606 346325 -4522 346561
rect -4286 346325 -4202 346561
rect -3966 346325 -3882 346561
rect -3646 346325 2918 346561
rect 3154 346325 9918 346561
rect 10154 346325 16918 346561
rect 17154 346325 23918 346561
rect 24154 346325 30918 346561
rect 31154 346325 37918 346561
rect 38154 346325 44918 346561
rect 45154 346325 51918 346561
rect 52154 346325 58918 346561
rect 59154 346325 65918 346561
rect 66154 346325 72918 346561
rect 73154 346325 79918 346561
rect 80154 346325 86918 346561
rect 87154 346325 93918 346561
rect 94154 346325 100918 346561
rect 101154 346325 107918 346561
rect 108154 346325 114918 346561
rect 115154 346325 121918 346561
rect 122154 346325 128918 346561
rect 129154 346325 135918 346561
rect 136154 346325 142918 346561
rect 143154 346325 149918 346561
rect 150154 346325 156918 346561
rect 157154 346325 163918 346561
rect 164154 346325 170918 346561
rect 171154 346325 177918 346561
rect 178154 346325 184918 346561
rect 185154 346325 191918 346561
rect 192154 346325 198918 346561
rect 199154 346325 205918 346561
rect 206154 346325 212918 346561
rect 213154 346325 219918 346561
rect 220154 346325 226918 346561
rect 227154 346325 233918 346561
rect 234154 346325 240918 346561
rect 241154 346325 247918 346561
rect 248154 346325 254918 346561
rect 255154 346325 261918 346561
rect 262154 346325 268918 346561
rect 269154 346325 275918 346561
rect 276154 346325 282918 346561
rect 283154 346325 289918 346561
rect 290154 346325 296918 346561
rect 297154 346325 303918 346561
rect 304154 346325 310918 346561
rect 311154 346325 317918 346561
rect 318154 346325 324918 346561
rect 325154 346325 331918 346561
rect 332154 346325 338918 346561
rect 339154 346325 345918 346561
rect 346154 346325 352918 346561
rect 353154 346325 359918 346561
rect 360154 346325 366918 346561
rect 367154 346325 373918 346561
rect 374154 346325 380918 346561
rect 381154 346325 387918 346561
rect 388154 346325 394918 346561
rect 395154 346325 401918 346561
rect 402154 346325 408918 346561
rect 409154 346325 415918 346561
rect 416154 346325 422918 346561
rect 423154 346325 429918 346561
rect 430154 346325 436918 346561
rect 437154 346325 443918 346561
rect 444154 346325 450918 346561
rect 451154 346325 457918 346561
rect 458154 346325 464918 346561
rect 465154 346325 471918 346561
rect 472154 346325 478918 346561
rect 479154 346325 485918 346561
rect 486154 346325 492918 346561
rect 493154 346325 499918 346561
rect 500154 346325 506918 346561
rect 507154 346325 513918 346561
rect 514154 346325 520918 346561
rect 521154 346325 527918 346561
rect 528154 346325 534918 346561
rect 535154 346325 541918 346561
rect 542154 346325 548918 346561
rect 549154 346325 555918 346561
rect 556154 346325 562918 346561
rect 563154 346325 569918 346561
rect 570154 346325 576918 346561
rect 577154 346325 587570 346561
rect 587806 346325 587890 346561
rect 588126 346325 588210 346561
rect 588446 346325 588530 346561
rect 588766 346325 588874 346561
rect -4950 346283 588874 346325
rect -4950 345494 588874 345536
rect -4950 345258 -3090 345494
rect -2854 345258 -2770 345494
rect -2534 345258 -2450 345494
rect -2214 345258 -2130 345494
rect -1894 345258 1186 345494
rect 1422 345258 8186 345494
rect 8422 345258 15186 345494
rect 15422 345258 22186 345494
rect 22422 345258 29186 345494
rect 29422 345258 36186 345494
rect 36422 345258 43186 345494
rect 43422 345258 50186 345494
rect 50422 345258 57186 345494
rect 57422 345258 64186 345494
rect 64422 345258 71186 345494
rect 71422 345258 78186 345494
rect 78422 345258 85186 345494
rect 85422 345258 92186 345494
rect 92422 345258 99186 345494
rect 99422 345258 106186 345494
rect 106422 345258 113186 345494
rect 113422 345258 120186 345494
rect 120422 345258 127186 345494
rect 127422 345258 134186 345494
rect 134422 345258 141186 345494
rect 141422 345258 148186 345494
rect 148422 345258 155186 345494
rect 155422 345258 162186 345494
rect 162422 345258 169186 345494
rect 169422 345258 176186 345494
rect 176422 345258 183186 345494
rect 183422 345258 190186 345494
rect 190422 345258 197186 345494
rect 197422 345258 204186 345494
rect 204422 345258 211186 345494
rect 211422 345258 218186 345494
rect 218422 345258 225186 345494
rect 225422 345258 232186 345494
rect 232422 345258 239186 345494
rect 239422 345258 246186 345494
rect 246422 345258 253186 345494
rect 253422 345258 260186 345494
rect 260422 345258 267186 345494
rect 267422 345258 274186 345494
rect 274422 345258 281186 345494
rect 281422 345258 288186 345494
rect 288422 345258 295186 345494
rect 295422 345258 302186 345494
rect 302422 345258 309186 345494
rect 309422 345258 316186 345494
rect 316422 345258 323186 345494
rect 323422 345258 330186 345494
rect 330422 345258 337186 345494
rect 337422 345258 344186 345494
rect 344422 345258 351186 345494
rect 351422 345258 358186 345494
rect 358422 345258 365186 345494
rect 365422 345258 372186 345494
rect 372422 345258 379186 345494
rect 379422 345258 386186 345494
rect 386422 345258 393186 345494
rect 393422 345258 400186 345494
rect 400422 345258 407186 345494
rect 407422 345258 414186 345494
rect 414422 345258 421186 345494
rect 421422 345258 428186 345494
rect 428422 345258 435186 345494
rect 435422 345258 442186 345494
rect 442422 345258 449186 345494
rect 449422 345258 456186 345494
rect 456422 345258 463186 345494
rect 463422 345258 470186 345494
rect 470422 345258 477186 345494
rect 477422 345258 484186 345494
rect 484422 345258 491186 345494
rect 491422 345258 498186 345494
rect 498422 345258 505186 345494
rect 505422 345258 512186 345494
rect 512422 345258 519186 345494
rect 519422 345258 526186 345494
rect 526422 345258 533186 345494
rect 533422 345258 540186 345494
rect 540422 345258 547186 345494
rect 547422 345258 554186 345494
rect 554422 345258 561186 345494
rect 561422 345258 568186 345494
rect 568422 345258 575186 345494
rect 575422 345258 582186 345494
rect 582422 345258 585818 345494
rect 586054 345258 586138 345494
rect 586374 345258 586458 345494
rect 586694 345258 586778 345494
rect 587014 345258 588874 345494
rect -4950 345216 588874 345258
rect -4950 339561 588874 339603
rect -4950 339325 -4842 339561
rect -4606 339325 -4522 339561
rect -4286 339325 -4202 339561
rect -3966 339325 -3882 339561
rect -3646 339325 2918 339561
rect 3154 339325 9918 339561
rect 10154 339325 16918 339561
rect 17154 339325 23918 339561
rect 24154 339325 30918 339561
rect 31154 339325 37918 339561
rect 38154 339325 44918 339561
rect 45154 339325 51918 339561
rect 52154 339325 58918 339561
rect 59154 339325 65918 339561
rect 66154 339325 72918 339561
rect 73154 339325 79918 339561
rect 80154 339325 86918 339561
rect 87154 339325 93918 339561
rect 94154 339325 100918 339561
rect 101154 339325 107918 339561
rect 108154 339325 114918 339561
rect 115154 339325 121918 339561
rect 122154 339325 128918 339561
rect 129154 339325 135918 339561
rect 136154 339325 142918 339561
rect 143154 339325 149918 339561
rect 150154 339325 156918 339561
rect 157154 339325 163918 339561
rect 164154 339325 170918 339561
rect 171154 339325 177918 339561
rect 178154 339325 184918 339561
rect 185154 339325 191918 339561
rect 192154 339325 198918 339561
rect 199154 339325 205918 339561
rect 206154 339325 212918 339561
rect 213154 339325 219918 339561
rect 220154 339325 226918 339561
rect 227154 339325 233918 339561
rect 234154 339325 240918 339561
rect 241154 339325 247918 339561
rect 248154 339325 254918 339561
rect 255154 339325 261918 339561
rect 262154 339325 268918 339561
rect 269154 339325 275918 339561
rect 276154 339325 282918 339561
rect 283154 339325 289918 339561
rect 290154 339325 296918 339561
rect 297154 339325 303918 339561
rect 304154 339325 310918 339561
rect 311154 339325 317918 339561
rect 318154 339325 324918 339561
rect 325154 339325 331918 339561
rect 332154 339325 338918 339561
rect 339154 339325 345918 339561
rect 346154 339325 352918 339561
rect 353154 339325 359918 339561
rect 360154 339325 366918 339561
rect 367154 339325 373918 339561
rect 374154 339325 380918 339561
rect 381154 339325 387918 339561
rect 388154 339325 394918 339561
rect 395154 339325 401918 339561
rect 402154 339325 408918 339561
rect 409154 339325 415918 339561
rect 416154 339325 422918 339561
rect 423154 339325 429918 339561
rect 430154 339325 436918 339561
rect 437154 339325 443918 339561
rect 444154 339325 450918 339561
rect 451154 339325 457918 339561
rect 458154 339325 464918 339561
rect 465154 339325 471918 339561
rect 472154 339325 478918 339561
rect 479154 339325 485918 339561
rect 486154 339325 492918 339561
rect 493154 339325 499918 339561
rect 500154 339325 506918 339561
rect 507154 339325 513918 339561
rect 514154 339325 520918 339561
rect 521154 339325 522850 339561
rect 523086 339325 524782 339561
rect 525018 339325 526714 339561
rect 526950 339325 527918 339561
rect 528154 339325 534918 339561
rect 535154 339325 541918 339561
rect 542154 339325 548918 339561
rect 549154 339325 555918 339561
rect 556154 339325 562918 339561
rect 563154 339325 569918 339561
rect 570154 339325 576918 339561
rect 577154 339325 587570 339561
rect 587806 339325 587890 339561
rect 588126 339325 588210 339561
rect 588446 339325 588530 339561
rect 588766 339325 588874 339561
rect -4950 339283 588874 339325
rect -4950 338494 588874 338536
rect -4950 338258 -3090 338494
rect -2854 338258 -2770 338494
rect -2534 338258 -2450 338494
rect -2214 338258 -2130 338494
rect -1894 338258 1186 338494
rect 1422 338258 8186 338494
rect 8422 338258 15186 338494
rect 15422 338258 22186 338494
rect 22422 338258 29186 338494
rect 29422 338258 36186 338494
rect 36422 338258 43186 338494
rect 43422 338258 50186 338494
rect 50422 338258 57186 338494
rect 57422 338258 64186 338494
rect 64422 338258 71186 338494
rect 71422 338258 78186 338494
rect 78422 338258 85186 338494
rect 85422 338258 92186 338494
rect 92422 338258 99186 338494
rect 99422 338258 106186 338494
rect 106422 338258 113186 338494
rect 113422 338258 120186 338494
rect 120422 338258 127186 338494
rect 127422 338258 134186 338494
rect 134422 338258 141186 338494
rect 141422 338258 148186 338494
rect 148422 338258 155186 338494
rect 155422 338258 162186 338494
rect 162422 338258 169186 338494
rect 169422 338258 176186 338494
rect 176422 338258 183186 338494
rect 183422 338258 190186 338494
rect 190422 338258 197186 338494
rect 197422 338258 204186 338494
rect 204422 338258 211186 338494
rect 211422 338258 218186 338494
rect 218422 338258 225186 338494
rect 225422 338258 232186 338494
rect 232422 338258 239186 338494
rect 239422 338258 246186 338494
rect 246422 338258 253186 338494
rect 253422 338258 260186 338494
rect 260422 338258 267186 338494
rect 267422 338258 274186 338494
rect 274422 338258 281186 338494
rect 281422 338258 288186 338494
rect 288422 338258 295186 338494
rect 295422 338258 302186 338494
rect 302422 338258 309186 338494
rect 309422 338258 316186 338494
rect 316422 338258 323186 338494
rect 323422 338258 330186 338494
rect 330422 338258 337186 338494
rect 337422 338258 344186 338494
rect 344422 338258 351186 338494
rect 351422 338258 358186 338494
rect 358422 338258 365186 338494
rect 365422 338258 372186 338494
rect 372422 338258 379186 338494
rect 379422 338258 386186 338494
rect 386422 338258 393186 338494
rect 393422 338258 400186 338494
rect 400422 338258 407186 338494
rect 407422 338258 414186 338494
rect 414422 338258 421186 338494
rect 421422 338258 428186 338494
rect 428422 338258 435186 338494
rect 435422 338258 442186 338494
rect 442422 338258 449186 338494
rect 449422 338258 456186 338494
rect 456422 338258 463186 338494
rect 463422 338258 470186 338494
rect 470422 338258 477186 338494
rect 477422 338258 484186 338494
rect 484422 338258 491186 338494
rect 491422 338258 498186 338494
rect 498422 338258 505186 338494
rect 505422 338258 512186 338494
rect 512422 338258 519186 338494
rect 519422 338258 519952 338494
rect 520188 338258 521884 338494
rect 522120 338258 523816 338494
rect 524052 338258 525748 338494
rect 525984 338258 533186 338494
rect 533422 338258 540186 338494
rect 540422 338258 547186 338494
rect 547422 338258 554186 338494
rect 554422 338258 561186 338494
rect 561422 338258 568186 338494
rect 568422 338258 575186 338494
rect 575422 338258 582186 338494
rect 582422 338258 585818 338494
rect 586054 338258 586138 338494
rect 586374 338258 586458 338494
rect 586694 338258 586778 338494
rect 587014 338258 588874 338494
rect -4950 338216 588874 338258
rect -4950 332561 588874 332603
rect -4950 332325 -4842 332561
rect -4606 332325 -4522 332561
rect -4286 332325 -4202 332561
rect -3966 332325 -3882 332561
rect -3646 332325 2918 332561
rect 3154 332325 9918 332561
rect 10154 332325 16918 332561
rect 17154 332325 23918 332561
rect 24154 332325 30918 332561
rect 31154 332325 37918 332561
rect 38154 332325 44918 332561
rect 45154 332325 51918 332561
rect 52154 332325 58918 332561
rect 59154 332325 65918 332561
rect 66154 332325 72918 332561
rect 73154 332325 79918 332561
rect 80154 332325 86918 332561
rect 87154 332325 93918 332561
rect 94154 332325 100918 332561
rect 101154 332325 107918 332561
rect 108154 332325 114918 332561
rect 115154 332325 121918 332561
rect 122154 332325 128918 332561
rect 129154 332325 135918 332561
rect 136154 332325 142918 332561
rect 143154 332325 149918 332561
rect 150154 332325 156918 332561
rect 157154 332325 163918 332561
rect 164154 332325 170918 332561
rect 171154 332325 177918 332561
rect 178154 332325 184918 332561
rect 185154 332325 191918 332561
rect 192154 332325 198918 332561
rect 199154 332325 205918 332561
rect 206154 332325 212918 332561
rect 213154 332325 219918 332561
rect 220154 332325 226918 332561
rect 227154 332325 233918 332561
rect 234154 332325 240918 332561
rect 241154 332325 247918 332561
rect 248154 332325 254918 332561
rect 255154 332325 261918 332561
rect 262154 332325 268918 332561
rect 269154 332325 275918 332561
rect 276154 332325 282918 332561
rect 283154 332325 289918 332561
rect 290154 332325 296918 332561
rect 297154 332325 303918 332561
rect 304154 332325 310918 332561
rect 311154 332325 317918 332561
rect 318154 332325 324918 332561
rect 325154 332325 331918 332561
rect 332154 332325 338918 332561
rect 339154 332325 345918 332561
rect 346154 332325 352918 332561
rect 353154 332325 359918 332561
rect 360154 332325 366918 332561
rect 367154 332325 373918 332561
rect 374154 332325 380918 332561
rect 381154 332325 387918 332561
rect 388154 332325 394918 332561
rect 395154 332325 401918 332561
rect 402154 332325 408918 332561
rect 409154 332325 415918 332561
rect 416154 332325 422918 332561
rect 423154 332325 429918 332561
rect 430154 332325 436918 332561
rect 437154 332325 443918 332561
rect 444154 332325 450918 332561
rect 451154 332325 457918 332561
rect 458154 332325 464918 332561
rect 465154 332325 471918 332561
rect 472154 332325 478918 332561
rect 479154 332325 485918 332561
rect 486154 332325 492918 332561
rect 493154 332325 499918 332561
rect 500154 332325 506918 332561
rect 507154 332325 513918 332561
rect 514154 332325 520918 332561
rect 521154 332325 522850 332561
rect 523086 332325 524782 332561
rect 525018 332325 526714 332561
rect 526950 332325 527918 332561
rect 528154 332325 534918 332561
rect 535154 332325 541918 332561
rect 542154 332325 548918 332561
rect 549154 332325 555918 332561
rect 556154 332325 562918 332561
rect 563154 332325 569918 332561
rect 570154 332325 576918 332561
rect 577154 332325 587570 332561
rect 587806 332325 587890 332561
rect 588126 332325 588210 332561
rect 588446 332325 588530 332561
rect 588766 332325 588874 332561
rect -4950 332283 588874 332325
rect -4950 331494 588874 331536
rect -4950 331258 -3090 331494
rect -2854 331258 -2770 331494
rect -2534 331258 -2450 331494
rect -2214 331258 -2130 331494
rect -1894 331258 1186 331494
rect 1422 331258 8186 331494
rect 8422 331258 15186 331494
rect 15422 331258 22186 331494
rect 22422 331258 29186 331494
rect 29422 331258 36186 331494
rect 36422 331258 43186 331494
rect 43422 331258 50186 331494
rect 50422 331258 57186 331494
rect 57422 331258 64186 331494
rect 64422 331258 71186 331494
rect 71422 331258 78186 331494
rect 78422 331258 85186 331494
rect 85422 331258 92186 331494
rect 92422 331258 99186 331494
rect 99422 331258 106186 331494
rect 106422 331258 113186 331494
rect 113422 331258 120186 331494
rect 120422 331258 127186 331494
rect 127422 331258 134186 331494
rect 134422 331258 141186 331494
rect 141422 331258 148186 331494
rect 148422 331258 155186 331494
rect 155422 331258 162186 331494
rect 162422 331258 169186 331494
rect 169422 331258 176186 331494
rect 176422 331258 183186 331494
rect 183422 331258 190186 331494
rect 190422 331258 197186 331494
rect 197422 331258 204186 331494
rect 204422 331258 211186 331494
rect 211422 331258 218186 331494
rect 218422 331258 225186 331494
rect 225422 331258 232186 331494
rect 232422 331258 239186 331494
rect 239422 331258 246186 331494
rect 246422 331258 253186 331494
rect 253422 331258 260186 331494
rect 260422 331258 267186 331494
rect 267422 331258 274186 331494
rect 274422 331258 281186 331494
rect 281422 331258 288186 331494
rect 288422 331258 295186 331494
rect 295422 331258 302186 331494
rect 302422 331258 309186 331494
rect 309422 331258 316186 331494
rect 316422 331258 323186 331494
rect 323422 331258 330186 331494
rect 330422 331258 337186 331494
rect 337422 331258 344186 331494
rect 344422 331258 351186 331494
rect 351422 331258 358186 331494
rect 358422 331258 365186 331494
rect 365422 331258 372186 331494
rect 372422 331258 379186 331494
rect 379422 331258 386186 331494
rect 386422 331258 393186 331494
rect 393422 331258 400186 331494
rect 400422 331258 407186 331494
rect 407422 331258 414186 331494
rect 414422 331258 421186 331494
rect 421422 331258 428186 331494
rect 428422 331258 435186 331494
rect 435422 331258 442186 331494
rect 442422 331258 449186 331494
rect 449422 331258 456186 331494
rect 456422 331258 463186 331494
rect 463422 331258 470186 331494
rect 470422 331258 477186 331494
rect 477422 331258 484186 331494
rect 484422 331258 491186 331494
rect 491422 331258 498186 331494
rect 498422 331258 505186 331494
rect 505422 331258 512186 331494
rect 512422 331258 519186 331494
rect 519422 331258 519952 331494
rect 520188 331258 521884 331494
rect 522120 331258 523816 331494
rect 524052 331258 525748 331494
rect 525984 331258 533186 331494
rect 533422 331258 540186 331494
rect 540422 331258 547186 331494
rect 547422 331258 554186 331494
rect 554422 331258 561186 331494
rect 561422 331258 568186 331494
rect 568422 331258 575186 331494
rect 575422 331258 582186 331494
rect 582422 331258 585818 331494
rect 586054 331258 586138 331494
rect 586374 331258 586458 331494
rect 586694 331258 586778 331494
rect 587014 331258 588874 331494
rect -4950 331216 588874 331258
rect -4950 325561 588874 325603
rect -4950 325325 -4842 325561
rect -4606 325325 -4522 325561
rect -4286 325325 -4202 325561
rect -3966 325325 -3882 325561
rect -3646 325325 2918 325561
rect 3154 325325 9918 325561
rect 10154 325325 16918 325561
rect 17154 325325 23918 325561
rect 24154 325325 30918 325561
rect 31154 325325 37918 325561
rect 38154 325325 44918 325561
rect 45154 325325 51918 325561
rect 52154 325325 58918 325561
rect 59154 325325 65918 325561
rect 66154 325325 72918 325561
rect 73154 325325 79918 325561
rect 80154 325325 86918 325561
rect 87154 325325 93918 325561
rect 94154 325325 100918 325561
rect 101154 325325 107918 325561
rect 108154 325325 114918 325561
rect 115154 325325 121918 325561
rect 122154 325325 128918 325561
rect 129154 325325 135918 325561
rect 136154 325325 142918 325561
rect 143154 325325 149918 325561
rect 150154 325325 156918 325561
rect 157154 325325 163918 325561
rect 164154 325325 170918 325561
rect 171154 325325 177918 325561
rect 178154 325325 184918 325561
rect 185154 325325 191918 325561
rect 192154 325325 198918 325561
rect 199154 325325 205918 325561
rect 206154 325325 212918 325561
rect 213154 325325 219918 325561
rect 220154 325325 226918 325561
rect 227154 325325 233918 325561
rect 234154 325325 240918 325561
rect 241154 325325 247918 325561
rect 248154 325325 254918 325561
rect 255154 325325 261918 325561
rect 262154 325325 268918 325561
rect 269154 325325 275918 325561
rect 276154 325325 282918 325561
rect 283154 325325 289918 325561
rect 290154 325325 296918 325561
rect 297154 325325 303918 325561
rect 304154 325325 310918 325561
rect 311154 325325 317918 325561
rect 318154 325325 324918 325561
rect 325154 325325 331918 325561
rect 332154 325325 338918 325561
rect 339154 325325 345918 325561
rect 346154 325325 352918 325561
rect 353154 325325 359918 325561
rect 360154 325325 366918 325561
rect 367154 325325 373918 325561
rect 374154 325325 380918 325561
rect 381154 325325 387918 325561
rect 388154 325325 394918 325561
rect 395154 325325 401918 325561
rect 402154 325325 408918 325561
rect 409154 325325 415918 325561
rect 416154 325325 422918 325561
rect 423154 325325 429918 325561
rect 430154 325325 436918 325561
rect 437154 325325 443918 325561
rect 444154 325325 450918 325561
rect 451154 325325 457918 325561
rect 458154 325325 464918 325561
rect 465154 325325 471918 325561
rect 472154 325325 478918 325561
rect 479154 325325 485918 325561
rect 486154 325325 492918 325561
rect 493154 325325 499918 325561
rect 500154 325325 506918 325561
rect 507154 325325 513918 325561
rect 514154 325325 520918 325561
rect 521154 325325 522850 325561
rect 523086 325325 524782 325561
rect 525018 325325 526714 325561
rect 526950 325325 527918 325561
rect 528154 325325 534918 325561
rect 535154 325325 541918 325561
rect 542154 325325 548918 325561
rect 549154 325325 555918 325561
rect 556154 325325 562918 325561
rect 563154 325325 569918 325561
rect 570154 325325 576918 325561
rect 577154 325325 587570 325561
rect 587806 325325 587890 325561
rect 588126 325325 588210 325561
rect 588446 325325 588530 325561
rect 588766 325325 588874 325561
rect -4950 325283 588874 325325
rect -4950 324494 588874 324536
rect -4950 324258 -3090 324494
rect -2854 324258 -2770 324494
rect -2534 324258 -2450 324494
rect -2214 324258 -2130 324494
rect -1894 324258 1186 324494
rect 1422 324258 8186 324494
rect 8422 324258 15186 324494
rect 15422 324258 22186 324494
rect 22422 324258 29186 324494
rect 29422 324258 36186 324494
rect 36422 324258 43186 324494
rect 43422 324258 50186 324494
rect 50422 324258 57186 324494
rect 57422 324258 64186 324494
rect 64422 324258 71186 324494
rect 71422 324258 78186 324494
rect 78422 324258 85186 324494
rect 85422 324258 92186 324494
rect 92422 324258 99186 324494
rect 99422 324258 106186 324494
rect 106422 324258 113186 324494
rect 113422 324258 120186 324494
rect 120422 324258 127186 324494
rect 127422 324258 134186 324494
rect 134422 324258 141186 324494
rect 141422 324258 148186 324494
rect 148422 324258 155186 324494
rect 155422 324258 162186 324494
rect 162422 324258 169186 324494
rect 169422 324258 176186 324494
rect 176422 324258 183186 324494
rect 183422 324258 190186 324494
rect 190422 324258 197186 324494
rect 197422 324258 204186 324494
rect 204422 324258 211186 324494
rect 211422 324258 218186 324494
rect 218422 324258 225186 324494
rect 225422 324258 232186 324494
rect 232422 324258 239186 324494
rect 239422 324258 246186 324494
rect 246422 324258 253186 324494
rect 253422 324258 260186 324494
rect 260422 324258 267186 324494
rect 267422 324258 274186 324494
rect 274422 324258 281186 324494
rect 281422 324258 288186 324494
rect 288422 324258 295186 324494
rect 295422 324258 302186 324494
rect 302422 324258 309186 324494
rect 309422 324258 316186 324494
rect 316422 324258 323186 324494
rect 323422 324258 330186 324494
rect 330422 324258 337186 324494
rect 337422 324258 344186 324494
rect 344422 324258 351186 324494
rect 351422 324258 358186 324494
rect 358422 324258 365186 324494
rect 365422 324258 372186 324494
rect 372422 324258 379186 324494
rect 379422 324258 386186 324494
rect 386422 324258 393186 324494
rect 393422 324258 400186 324494
rect 400422 324258 407186 324494
rect 407422 324258 414186 324494
rect 414422 324258 421186 324494
rect 421422 324258 428186 324494
rect 428422 324258 435186 324494
rect 435422 324258 442186 324494
rect 442422 324258 449186 324494
rect 449422 324258 456186 324494
rect 456422 324258 463186 324494
rect 463422 324258 470186 324494
rect 470422 324258 477186 324494
rect 477422 324258 484186 324494
rect 484422 324258 491186 324494
rect 491422 324258 498186 324494
rect 498422 324258 505186 324494
rect 505422 324258 512186 324494
rect 512422 324258 519186 324494
rect 519422 324258 519952 324494
rect 520188 324258 521884 324494
rect 522120 324258 523816 324494
rect 524052 324258 525748 324494
rect 525984 324258 533186 324494
rect 533422 324258 540186 324494
rect 540422 324258 547186 324494
rect 547422 324258 554186 324494
rect 554422 324258 561186 324494
rect 561422 324258 568186 324494
rect 568422 324258 575186 324494
rect 575422 324258 582186 324494
rect 582422 324258 585818 324494
rect 586054 324258 586138 324494
rect 586374 324258 586458 324494
rect 586694 324258 586778 324494
rect 587014 324258 588874 324494
rect -4950 324216 588874 324258
rect -4950 318561 588874 318603
rect -4950 318325 -4842 318561
rect -4606 318325 -4522 318561
rect -4286 318325 -4202 318561
rect -3966 318325 -3882 318561
rect -3646 318325 2918 318561
rect 3154 318325 9918 318561
rect 10154 318325 16918 318561
rect 17154 318325 23918 318561
rect 24154 318325 30918 318561
rect 31154 318325 37918 318561
rect 38154 318325 44918 318561
rect 45154 318325 51918 318561
rect 52154 318325 58918 318561
rect 59154 318325 65918 318561
rect 66154 318325 72918 318561
rect 73154 318325 79918 318561
rect 80154 318325 86918 318561
rect 87154 318325 93918 318561
rect 94154 318325 100918 318561
rect 101154 318325 107918 318561
rect 108154 318325 114918 318561
rect 115154 318325 121918 318561
rect 122154 318325 128918 318561
rect 129154 318325 135918 318561
rect 136154 318325 142918 318561
rect 143154 318325 149918 318561
rect 150154 318325 156918 318561
rect 157154 318325 163918 318561
rect 164154 318325 170918 318561
rect 171154 318325 177918 318561
rect 178154 318325 184918 318561
rect 185154 318325 191918 318561
rect 192154 318325 198918 318561
rect 199154 318325 205918 318561
rect 206154 318325 212918 318561
rect 213154 318325 219918 318561
rect 220154 318325 226918 318561
rect 227154 318325 233918 318561
rect 234154 318325 240918 318561
rect 241154 318325 247918 318561
rect 248154 318325 254918 318561
rect 255154 318325 261918 318561
rect 262154 318325 268918 318561
rect 269154 318325 275918 318561
rect 276154 318325 282918 318561
rect 283154 318325 289918 318561
rect 290154 318325 296918 318561
rect 297154 318325 303918 318561
rect 304154 318325 310918 318561
rect 311154 318325 317918 318561
rect 318154 318325 324918 318561
rect 325154 318325 331918 318561
rect 332154 318325 338918 318561
rect 339154 318325 345918 318561
rect 346154 318325 352918 318561
rect 353154 318325 359918 318561
rect 360154 318325 366918 318561
rect 367154 318325 373918 318561
rect 374154 318325 380918 318561
rect 381154 318325 387918 318561
rect 388154 318325 394918 318561
rect 395154 318325 401918 318561
rect 402154 318325 408918 318561
rect 409154 318325 415918 318561
rect 416154 318325 422918 318561
rect 423154 318325 429918 318561
rect 430154 318325 436918 318561
rect 437154 318325 443918 318561
rect 444154 318325 450918 318561
rect 451154 318325 457918 318561
rect 458154 318325 464918 318561
rect 465154 318325 471918 318561
rect 472154 318325 478918 318561
rect 479154 318325 485918 318561
rect 486154 318325 492918 318561
rect 493154 318325 499918 318561
rect 500154 318325 506918 318561
rect 507154 318325 513918 318561
rect 514154 318325 520918 318561
rect 521154 318325 527918 318561
rect 528154 318325 534918 318561
rect 535154 318325 541918 318561
rect 542154 318325 548918 318561
rect 549154 318325 555918 318561
rect 556154 318325 562918 318561
rect 563154 318325 569918 318561
rect 570154 318325 576918 318561
rect 577154 318325 587570 318561
rect 587806 318325 587890 318561
rect 588126 318325 588210 318561
rect 588446 318325 588530 318561
rect 588766 318325 588874 318561
rect -4950 318283 588874 318325
rect -4950 317494 588874 317536
rect -4950 317258 -3090 317494
rect -2854 317258 -2770 317494
rect -2534 317258 -2450 317494
rect -2214 317258 -2130 317494
rect -1894 317258 1186 317494
rect 1422 317258 8186 317494
rect 8422 317258 15186 317494
rect 15422 317258 22186 317494
rect 22422 317258 29186 317494
rect 29422 317258 36186 317494
rect 36422 317258 43186 317494
rect 43422 317258 50186 317494
rect 50422 317258 57186 317494
rect 57422 317258 64186 317494
rect 64422 317258 71186 317494
rect 71422 317258 78186 317494
rect 78422 317258 85186 317494
rect 85422 317258 92186 317494
rect 92422 317258 99186 317494
rect 99422 317258 106186 317494
rect 106422 317258 113186 317494
rect 113422 317258 120186 317494
rect 120422 317258 127186 317494
rect 127422 317258 134186 317494
rect 134422 317258 141186 317494
rect 141422 317258 148186 317494
rect 148422 317258 155186 317494
rect 155422 317258 162186 317494
rect 162422 317258 169186 317494
rect 169422 317258 176186 317494
rect 176422 317258 183186 317494
rect 183422 317258 190186 317494
rect 190422 317258 197186 317494
rect 197422 317258 204186 317494
rect 204422 317258 211186 317494
rect 211422 317258 218186 317494
rect 218422 317258 225186 317494
rect 225422 317258 232186 317494
rect 232422 317258 239186 317494
rect 239422 317258 246186 317494
rect 246422 317258 253186 317494
rect 253422 317258 260186 317494
rect 260422 317258 267186 317494
rect 267422 317258 274186 317494
rect 274422 317258 281186 317494
rect 281422 317258 288186 317494
rect 288422 317258 295186 317494
rect 295422 317258 302186 317494
rect 302422 317258 309186 317494
rect 309422 317258 316186 317494
rect 316422 317258 323186 317494
rect 323422 317258 330186 317494
rect 330422 317258 337186 317494
rect 337422 317258 344186 317494
rect 344422 317258 351186 317494
rect 351422 317258 358186 317494
rect 358422 317258 365186 317494
rect 365422 317258 372186 317494
rect 372422 317258 379186 317494
rect 379422 317258 386186 317494
rect 386422 317258 393186 317494
rect 393422 317258 400186 317494
rect 400422 317258 407186 317494
rect 407422 317258 414186 317494
rect 414422 317258 421186 317494
rect 421422 317258 428186 317494
rect 428422 317258 435186 317494
rect 435422 317258 442186 317494
rect 442422 317258 449186 317494
rect 449422 317258 456186 317494
rect 456422 317258 463186 317494
rect 463422 317258 470186 317494
rect 470422 317258 477186 317494
rect 477422 317258 484186 317494
rect 484422 317258 491186 317494
rect 491422 317258 498186 317494
rect 498422 317258 505186 317494
rect 505422 317258 512186 317494
rect 512422 317258 519186 317494
rect 519422 317258 526186 317494
rect 526422 317258 533186 317494
rect 533422 317258 540186 317494
rect 540422 317258 547186 317494
rect 547422 317258 554186 317494
rect 554422 317258 561186 317494
rect 561422 317258 568186 317494
rect 568422 317258 575186 317494
rect 575422 317258 582186 317494
rect 582422 317258 585818 317494
rect 586054 317258 586138 317494
rect 586374 317258 586458 317494
rect 586694 317258 586778 317494
rect 587014 317258 588874 317494
rect -4950 317216 588874 317258
rect -4950 311561 588874 311603
rect -4950 311325 -4842 311561
rect -4606 311325 -4522 311561
rect -4286 311325 -4202 311561
rect -3966 311325 -3882 311561
rect -3646 311325 2918 311561
rect 3154 311325 9918 311561
rect 10154 311325 16918 311561
rect 17154 311325 23918 311561
rect 24154 311325 30918 311561
rect 31154 311325 37918 311561
rect 38154 311325 44918 311561
rect 45154 311325 51918 311561
rect 52154 311325 58918 311561
rect 59154 311325 65918 311561
rect 66154 311325 72918 311561
rect 73154 311325 79918 311561
rect 80154 311325 86918 311561
rect 87154 311325 93918 311561
rect 94154 311325 100918 311561
rect 101154 311325 107918 311561
rect 108154 311325 114918 311561
rect 115154 311325 121918 311561
rect 122154 311325 128918 311561
rect 129154 311325 135918 311561
rect 136154 311325 142918 311561
rect 143154 311325 149918 311561
rect 150154 311325 156918 311561
rect 157154 311325 163918 311561
rect 164154 311325 170918 311561
rect 171154 311325 177918 311561
rect 178154 311325 184918 311561
rect 185154 311325 191918 311561
rect 192154 311325 198918 311561
rect 199154 311325 205918 311561
rect 206154 311325 212918 311561
rect 213154 311325 219918 311561
rect 220154 311325 226918 311561
rect 227154 311325 233918 311561
rect 234154 311325 240918 311561
rect 241154 311325 247918 311561
rect 248154 311325 254918 311561
rect 255154 311325 261918 311561
rect 262154 311325 268918 311561
rect 269154 311325 275918 311561
rect 276154 311325 282918 311561
rect 283154 311325 289918 311561
rect 290154 311325 296918 311561
rect 297154 311325 303918 311561
rect 304154 311325 310918 311561
rect 311154 311325 317918 311561
rect 318154 311325 324918 311561
rect 325154 311325 331918 311561
rect 332154 311325 338918 311561
rect 339154 311325 345918 311561
rect 346154 311325 352918 311561
rect 353154 311325 359918 311561
rect 360154 311325 366918 311561
rect 367154 311325 373918 311561
rect 374154 311325 380918 311561
rect 381154 311325 387918 311561
rect 388154 311325 394918 311561
rect 395154 311325 401918 311561
rect 402154 311325 408918 311561
rect 409154 311325 415918 311561
rect 416154 311325 422918 311561
rect 423154 311325 429918 311561
rect 430154 311325 436918 311561
rect 437154 311325 443918 311561
rect 444154 311325 450918 311561
rect 451154 311325 457918 311561
rect 458154 311325 464918 311561
rect 465154 311325 471918 311561
rect 472154 311325 478918 311561
rect 479154 311325 485918 311561
rect 486154 311325 492918 311561
rect 493154 311325 499918 311561
rect 500154 311325 506918 311561
rect 507154 311325 513918 311561
rect 514154 311325 520918 311561
rect 521154 311325 527918 311561
rect 528154 311325 534918 311561
rect 535154 311325 541918 311561
rect 542154 311325 548918 311561
rect 549154 311325 555918 311561
rect 556154 311325 562918 311561
rect 563154 311325 569918 311561
rect 570154 311325 576918 311561
rect 577154 311325 587570 311561
rect 587806 311325 587890 311561
rect 588126 311325 588210 311561
rect 588446 311325 588530 311561
rect 588766 311325 588874 311561
rect -4950 311283 588874 311325
rect -4950 310494 588874 310536
rect -4950 310258 -3090 310494
rect -2854 310258 -2770 310494
rect -2534 310258 -2450 310494
rect -2214 310258 -2130 310494
rect -1894 310258 1186 310494
rect 1422 310258 8186 310494
rect 8422 310258 15186 310494
rect 15422 310258 22186 310494
rect 22422 310258 29186 310494
rect 29422 310258 36186 310494
rect 36422 310258 43186 310494
rect 43422 310258 50186 310494
rect 50422 310258 57186 310494
rect 57422 310258 64186 310494
rect 64422 310258 71186 310494
rect 71422 310258 78186 310494
rect 78422 310258 85186 310494
rect 85422 310258 92186 310494
rect 92422 310258 99186 310494
rect 99422 310258 106186 310494
rect 106422 310258 113186 310494
rect 113422 310258 120186 310494
rect 120422 310258 127186 310494
rect 127422 310258 134186 310494
rect 134422 310258 141186 310494
rect 141422 310258 148186 310494
rect 148422 310258 155186 310494
rect 155422 310258 162186 310494
rect 162422 310258 169186 310494
rect 169422 310258 176186 310494
rect 176422 310258 183186 310494
rect 183422 310258 190186 310494
rect 190422 310258 197186 310494
rect 197422 310258 204186 310494
rect 204422 310258 211186 310494
rect 211422 310258 218186 310494
rect 218422 310258 225186 310494
rect 225422 310258 232186 310494
rect 232422 310258 239186 310494
rect 239422 310258 246186 310494
rect 246422 310258 253186 310494
rect 253422 310258 260186 310494
rect 260422 310258 267186 310494
rect 267422 310258 274186 310494
rect 274422 310258 281186 310494
rect 281422 310258 288186 310494
rect 288422 310258 295186 310494
rect 295422 310258 302186 310494
rect 302422 310258 309186 310494
rect 309422 310258 316186 310494
rect 316422 310258 323186 310494
rect 323422 310258 330186 310494
rect 330422 310258 337186 310494
rect 337422 310258 344186 310494
rect 344422 310258 351186 310494
rect 351422 310258 358186 310494
rect 358422 310258 365186 310494
rect 365422 310258 372186 310494
rect 372422 310258 379186 310494
rect 379422 310258 386186 310494
rect 386422 310258 393186 310494
rect 393422 310258 400186 310494
rect 400422 310258 407186 310494
rect 407422 310258 414186 310494
rect 414422 310258 421186 310494
rect 421422 310258 428186 310494
rect 428422 310258 435186 310494
rect 435422 310258 442186 310494
rect 442422 310258 449186 310494
rect 449422 310258 456186 310494
rect 456422 310258 463186 310494
rect 463422 310258 470186 310494
rect 470422 310258 477186 310494
rect 477422 310258 484186 310494
rect 484422 310258 491186 310494
rect 491422 310258 498186 310494
rect 498422 310258 505186 310494
rect 505422 310258 512186 310494
rect 512422 310258 519186 310494
rect 519422 310258 526186 310494
rect 526422 310258 533186 310494
rect 533422 310258 540186 310494
rect 540422 310258 547186 310494
rect 547422 310258 554186 310494
rect 554422 310258 561186 310494
rect 561422 310258 568186 310494
rect 568422 310258 575186 310494
rect 575422 310258 582186 310494
rect 582422 310258 585818 310494
rect 586054 310258 586138 310494
rect 586374 310258 586458 310494
rect 586694 310258 586778 310494
rect 587014 310258 588874 310494
rect -4950 310216 588874 310258
rect -4950 304561 588874 304603
rect -4950 304325 -4842 304561
rect -4606 304325 -4522 304561
rect -4286 304325 -4202 304561
rect -3966 304325 -3882 304561
rect -3646 304325 2918 304561
rect 3154 304325 9918 304561
rect 10154 304325 16918 304561
rect 17154 304325 23918 304561
rect 24154 304325 30918 304561
rect 31154 304325 37918 304561
rect 38154 304325 44918 304561
rect 45154 304325 51918 304561
rect 52154 304325 58918 304561
rect 59154 304325 65918 304561
rect 66154 304325 72918 304561
rect 73154 304325 79918 304561
rect 80154 304325 86918 304561
rect 87154 304325 93918 304561
rect 94154 304325 100918 304561
rect 101154 304325 107918 304561
rect 108154 304325 114918 304561
rect 115154 304325 121918 304561
rect 122154 304325 128918 304561
rect 129154 304325 135918 304561
rect 136154 304325 142918 304561
rect 143154 304325 149918 304561
rect 150154 304325 156918 304561
rect 157154 304325 163918 304561
rect 164154 304325 170918 304561
rect 171154 304325 177918 304561
rect 178154 304325 184918 304561
rect 185154 304325 191918 304561
rect 192154 304325 198918 304561
rect 199154 304325 205918 304561
rect 206154 304325 212918 304561
rect 213154 304325 219918 304561
rect 220154 304325 226918 304561
rect 227154 304325 233918 304561
rect 234154 304325 240918 304561
rect 241154 304325 247918 304561
rect 248154 304325 254918 304561
rect 255154 304325 261918 304561
rect 262154 304325 268918 304561
rect 269154 304325 275918 304561
rect 276154 304325 282918 304561
rect 283154 304325 289918 304561
rect 290154 304325 296918 304561
rect 297154 304325 303918 304561
rect 304154 304325 310918 304561
rect 311154 304325 317918 304561
rect 318154 304325 324918 304561
rect 325154 304325 331918 304561
rect 332154 304325 338918 304561
rect 339154 304325 345918 304561
rect 346154 304325 352918 304561
rect 353154 304325 359918 304561
rect 360154 304325 366918 304561
rect 367154 304325 373918 304561
rect 374154 304325 380918 304561
rect 381154 304325 387918 304561
rect 388154 304325 394918 304561
rect 395154 304325 401918 304561
rect 402154 304325 408918 304561
rect 409154 304325 415918 304561
rect 416154 304325 422918 304561
rect 423154 304325 429918 304561
rect 430154 304325 436918 304561
rect 437154 304325 443918 304561
rect 444154 304325 450918 304561
rect 451154 304325 457918 304561
rect 458154 304325 464918 304561
rect 465154 304325 471918 304561
rect 472154 304325 478918 304561
rect 479154 304325 485918 304561
rect 486154 304325 492918 304561
rect 493154 304325 499918 304561
rect 500154 304325 506918 304561
rect 507154 304325 513918 304561
rect 514154 304325 520918 304561
rect 521154 304325 527918 304561
rect 528154 304325 534918 304561
rect 535154 304325 541918 304561
rect 542154 304325 548918 304561
rect 549154 304325 555918 304561
rect 556154 304325 562918 304561
rect 563154 304325 569918 304561
rect 570154 304325 576918 304561
rect 577154 304325 587570 304561
rect 587806 304325 587890 304561
rect 588126 304325 588210 304561
rect 588446 304325 588530 304561
rect 588766 304325 588874 304561
rect -4950 304283 588874 304325
rect -4950 303494 588874 303536
rect -4950 303258 -3090 303494
rect -2854 303258 -2770 303494
rect -2534 303258 -2450 303494
rect -2214 303258 -2130 303494
rect -1894 303258 1186 303494
rect 1422 303258 8186 303494
rect 8422 303258 15186 303494
rect 15422 303258 22186 303494
rect 22422 303258 29186 303494
rect 29422 303258 36186 303494
rect 36422 303258 43186 303494
rect 43422 303258 50186 303494
rect 50422 303258 57186 303494
rect 57422 303258 64186 303494
rect 64422 303258 71186 303494
rect 71422 303258 78186 303494
rect 78422 303258 85186 303494
rect 85422 303258 92186 303494
rect 92422 303258 99186 303494
rect 99422 303258 106186 303494
rect 106422 303258 113186 303494
rect 113422 303258 120186 303494
rect 120422 303258 127186 303494
rect 127422 303258 134186 303494
rect 134422 303258 141186 303494
rect 141422 303258 148186 303494
rect 148422 303258 155186 303494
rect 155422 303258 162186 303494
rect 162422 303258 169186 303494
rect 169422 303258 176186 303494
rect 176422 303258 183186 303494
rect 183422 303258 190186 303494
rect 190422 303258 197186 303494
rect 197422 303258 204186 303494
rect 204422 303258 211186 303494
rect 211422 303258 218186 303494
rect 218422 303258 225186 303494
rect 225422 303258 232186 303494
rect 232422 303258 239186 303494
rect 239422 303258 246186 303494
rect 246422 303258 253186 303494
rect 253422 303258 260186 303494
rect 260422 303258 267186 303494
rect 267422 303258 274186 303494
rect 274422 303258 281186 303494
rect 281422 303258 288186 303494
rect 288422 303258 295186 303494
rect 295422 303258 302186 303494
rect 302422 303258 309186 303494
rect 309422 303258 316186 303494
rect 316422 303258 323186 303494
rect 323422 303258 330186 303494
rect 330422 303258 337186 303494
rect 337422 303258 344186 303494
rect 344422 303258 351186 303494
rect 351422 303258 358186 303494
rect 358422 303258 365186 303494
rect 365422 303258 372186 303494
rect 372422 303258 379186 303494
rect 379422 303258 386186 303494
rect 386422 303258 393186 303494
rect 393422 303258 400186 303494
rect 400422 303258 407186 303494
rect 407422 303258 414186 303494
rect 414422 303258 421186 303494
rect 421422 303258 428186 303494
rect 428422 303258 435186 303494
rect 435422 303258 442186 303494
rect 442422 303258 449186 303494
rect 449422 303258 456186 303494
rect 456422 303258 463186 303494
rect 463422 303258 470186 303494
rect 470422 303258 477186 303494
rect 477422 303258 484186 303494
rect 484422 303258 491186 303494
rect 491422 303258 498186 303494
rect 498422 303258 505186 303494
rect 505422 303258 512186 303494
rect 512422 303258 519186 303494
rect 519422 303258 526186 303494
rect 526422 303258 533186 303494
rect 533422 303258 540186 303494
rect 540422 303258 547186 303494
rect 547422 303258 554186 303494
rect 554422 303258 561186 303494
rect 561422 303258 568186 303494
rect 568422 303258 575186 303494
rect 575422 303258 582186 303494
rect 582422 303258 585818 303494
rect 586054 303258 586138 303494
rect 586374 303258 586458 303494
rect 586694 303258 586778 303494
rect 587014 303258 588874 303494
rect -4950 303216 588874 303258
rect -4950 297561 588874 297603
rect -4950 297325 -4842 297561
rect -4606 297325 -4522 297561
rect -4286 297325 -4202 297561
rect -3966 297325 -3882 297561
rect -3646 297325 2918 297561
rect 3154 297325 9918 297561
rect 10154 297325 16918 297561
rect 17154 297325 23918 297561
rect 24154 297325 30918 297561
rect 31154 297325 37918 297561
rect 38154 297325 44918 297561
rect 45154 297325 51918 297561
rect 52154 297325 58918 297561
rect 59154 297325 65918 297561
rect 66154 297325 72918 297561
rect 73154 297325 79918 297561
rect 80154 297325 86918 297561
rect 87154 297325 93918 297561
rect 94154 297325 100918 297561
rect 101154 297325 107918 297561
rect 108154 297325 114918 297561
rect 115154 297325 121918 297561
rect 122154 297325 128918 297561
rect 129154 297325 135918 297561
rect 136154 297325 142918 297561
rect 143154 297325 149918 297561
rect 150154 297325 156918 297561
rect 157154 297325 163918 297561
rect 164154 297325 170918 297561
rect 171154 297325 177918 297561
rect 178154 297325 184918 297561
rect 185154 297325 191918 297561
rect 192154 297325 198918 297561
rect 199154 297325 205918 297561
rect 206154 297325 212918 297561
rect 213154 297325 219918 297561
rect 220154 297325 226918 297561
rect 227154 297325 233918 297561
rect 234154 297325 240918 297561
rect 241154 297325 247918 297561
rect 248154 297325 254918 297561
rect 255154 297325 261918 297561
rect 262154 297325 268918 297561
rect 269154 297325 275918 297561
rect 276154 297325 282918 297561
rect 283154 297325 289918 297561
rect 290154 297325 296918 297561
rect 297154 297325 303918 297561
rect 304154 297325 310918 297561
rect 311154 297325 317918 297561
rect 318154 297325 324918 297561
rect 325154 297325 331918 297561
rect 332154 297325 338918 297561
rect 339154 297325 345918 297561
rect 346154 297325 352918 297561
rect 353154 297325 359918 297561
rect 360154 297325 366918 297561
rect 367154 297325 373918 297561
rect 374154 297325 380918 297561
rect 381154 297325 387918 297561
rect 388154 297325 394918 297561
rect 395154 297325 401918 297561
rect 402154 297325 408918 297561
rect 409154 297325 415918 297561
rect 416154 297325 422918 297561
rect 423154 297325 429918 297561
rect 430154 297325 436918 297561
rect 437154 297325 443918 297561
rect 444154 297325 450918 297561
rect 451154 297325 457918 297561
rect 458154 297325 464918 297561
rect 465154 297325 471918 297561
rect 472154 297325 478918 297561
rect 479154 297325 485918 297561
rect 486154 297325 492918 297561
rect 493154 297325 499918 297561
rect 500154 297325 506918 297561
rect 507154 297325 513918 297561
rect 514154 297325 520918 297561
rect 521154 297325 522850 297561
rect 523086 297325 524782 297561
rect 525018 297325 526714 297561
rect 526950 297325 527918 297561
rect 528154 297325 534918 297561
rect 535154 297325 541918 297561
rect 542154 297325 548918 297561
rect 549154 297325 555918 297561
rect 556154 297325 562918 297561
rect 563154 297325 569918 297561
rect 570154 297325 576918 297561
rect 577154 297325 587570 297561
rect 587806 297325 587890 297561
rect 588126 297325 588210 297561
rect 588446 297325 588530 297561
rect 588766 297325 588874 297561
rect -4950 297283 588874 297325
rect -4950 296494 588874 296536
rect -4950 296258 -3090 296494
rect -2854 296258 -2770 296494
rect -2534 296258 -2450 296494
rect -2214 296258 -2130 296494
rect -1894 296258 1186 296494
rect 1422 296258 8186 296494
rect 8422 296258 15186 296494
rect 15422 296258 22186 296494
rect 22422 296258 29186 296494
rect 29422 296258 36186 296494
rect 36422 296258 43186 296494
rect 43422 296258 50186 296494
rect 50422 296258 57186 296494
rect 57422 296258 64186 296494
rect 64422 296258 71186 296494
rect 71422 296258 78186 296494
rect 78422 296258 85186 296494
rect 85422 296258 92186 296494
rect 92422 296258 99186 296494
rect 99422 296258 106186 296494
rect 106422 296258 113186 296494
rect 113422 296258 120186 296494
rect 120422 296258 127186 296494
rect 127422 296258 134186 296494
rect 134422 296258 141186 296494
rect 141422 296258 148186 296494
rect 148422 296258 155186 296494
rect 155422 296258 162186 296494
rect 162422 296258 169186 296494
rect 169422 296258 176186 296494
rect 176422 296258 183186 296494
rect 183422 296258 190186 296494
rect 190422 296258 197186 296494
rect 197422 296258 204186 296494
rect 204422 296258 211186 296494
rect 211422 296258 218186 296494
rect 218422 296258 225186 296494
rect 225422 296258 232186 296494
rect 232422 296258 239186 296494
rect 239422 296258 246186 296494
rect 246422 296258 253186 296494
rect 253422 296258 260186 296494
rect 260422 296258 267186 296494
rect 267422 296258 274186 296494
rect 274422 296258 281186 296494
rect 281422 296258 288186 296494
rect 288422 296258 295186 296494
rect 295422 296258 302186 296494
rect 302422 296258 309186 296494
rect 309422 296258 316186 296494
rect 316422 296258 323186 296494
rect 323422 296258 330186 296494
rect 330422 296258 337186 296494
rect 337422 296258 344186 296494
rect 344422 296258 351186 296494
rect 351422 296258 358186 296494
rect 358422 296258 365186 296494
rect 365422 296258 372186 296494
rect 372422 296258 379186 296494
rect 379422 296258 386186 296494
rect 386422 296258 393186 296494
rect 393422 296258 400186 296494
rect 400422 296258 407186 296494
rect 407422 296258 414186 296494
rect 414422 296258 421186 296494
rect 421422 296258 428186 296494
rect 428422 296258 435186 296494
rect 435422 296258 442186 296494
rect 442422 296258 449186 296494
rect 449422 296258 456186 296494
rect 456422 296258 463186 296494
rect 463422 296258 470186 296494
rect 470422 296258 477186 296494
rect 477422 296258 484186 296494
rect 484422 296258 491186 296494
rect 491422 296258 498186 296494
rect 498422 296258 505186 296494
rect 505422 296258 512186 296494
rect 512422 296258 519186 296494
rect 519422 296258 519952 296494
rect 520188 296258 521884 296494
rect 522120 296258 523816 296494
rect 524052 296258 525748 296494
rect 525984 296258 533186 296494
rect 533422 296258 540186 296494
rect 540422 296258 547186 296494
rect 547422 296258 554186 296494
rect 554422 296258 561186 296494
rect 561422 296258 568186 296494
rect 568422 296258 575186 296494
rect 575422 296258 582186 296494
rect 582422 296258 585818 296494
rect 586054 296258 586138 296494
rect 586374 296258 586458 296494
rect 586694 296258 586778 296494
rect 587014 296258 588874 296494
rect -4950 296216 588874 296258
rect -4950 290561 588874 290603
rect -4950 290325 -4842 290561
rect -4606 290325 -4522 290561
rect -4286 290325 -4202 290561
rect -3966 290325 -3882 290561
rect -3646 290325 2918 290561
rect 3154 290325 9918 290561
rect 10154 290325 16918 290561
rect 17154 290325 23918 290561
rect 24154 290325 30918 290561
rect 31154 290325 37918 290561
rect 38154 290325 44918 290561
rect 45154 290325 51918 290561
rect 52154 290325 58918 290561
rect 59154 290325 65918 290561
rect 66154 290325 72918 290561
rect 73154 290325 79918 290561
rect 80154 290325 86918 290561
rect 87154 290325 93918 290561
rect 94154 290325 100918 290561
rect 101154 290325 107918 290561
rect 108154 290325 114918 290561
rect 115154 290325 121918 290561
rect 122154 290325 128918 290561
rect 129154 290325 135918 290561
rect 136154 290325 142918 290561
rect 143154 290325 149918 290561
rect 150154 290325 156918 290561
rect 157154 290325 163918 290561
rect 164154 290325 170918 290561
rect 171154 290325 177918 290561
rect 178154 290325 184918 290561
rect 185154 290325 191918 290561
rect 192154 290325 198918 290561
rect 199154 290325 205918 290561
rect 206154 290325 212918 290561
rect 213154 290325 219918 290561
rect 220154 290325 226918 290561
rect 227154 290325 233918 290561
rect 234154 290325 240918 290561
rect 241154 290325 247918 290561
rect 248154 290325 254918 290561
rect 255154 290325 261918 290561
rect 262154 290325 268918 290561
rect 269154 290325 275918 290561
rect 276154 290325 282918 290561
rect 283154 290325 289918 290561
rect 290154 290325 296918 290561
rect 297154 290325 303918 290561
rect 304154 290325 310918 290561
rect 311154 290325 317918 290561
rect 318154 290325 324918 290561
rect 325154 290325 331918 290561
rect 332154 290325 338918 290561
rect 339154 290325 345918 290561
rect 346154 290325 352918 290561
rect 353154 290325 359918 290561
rect 360154 290325 366918 290561
rect 367154 290325 373918 290561
rect 374154 290325 380918 290561
rect 381154 290325 387918 290561
rect 388154 290325 394918 290561
rect 395154 290325 401918 290561
rect 402154 290325 408918 290561
rect 409154 290325 415918 290561
rect 416154 290325 422918 290561
rect 423154 290325 429918 290561
rect 430154 290325 436918 290561
rect 437154 290325 443918 290561
rect 444154 290325 450918 290561
rect 451154 290325 457918 290561
rect 458154 290325 464918 290561
rect 465154 290325 471918 290561
rect 472154 290325 478918 290561
rect 479154 290325 485918 290561
rect 486154 290325 492918 290561
rect 493154 290325 499918 290561
rect 500154 290325 506918 290561
rect 507154 290325 513918 290561
rect 514154 290325 520918 290561
rect 521154 290325 522850 290561
rect 523086 290325 524782 290561
rect 525018 290325 526714 290561
rect 526950 290325 527918 290561
rect 528154 290325 534918 290561
rect 535154 290325 541918 290561
rect 542154 290325 548918 290561
rect 549154 290325 555918 290561
rect 556154 290325 562918 290561
rect 563154 290325 569918 290561
rect 570154 290325 576918 290561
rect 577154 290325 587570 290561
rect 587806 290325 587890 290561
rect 588126 290325 588210 290561
rect 588446 290325 588530 290561
rect 588766 290325 588874 290561
rect -4950 290283 588874 290325
rect -4950 289494 588874 289536
rect -4950 289258 -3090 289494
rect -2854 289258 -2770 289494
rect -2534 289258 -2450 289494
rect -2214 289258 -2130 289494
rect -1894 289258 1186 289494
rect 1422 289258 8186 289494
rect 8422 289258 15186 289494
rect 15422 289258 22186 289494
rect 22422 289258 29186 289494
rect 29422 289258 36186 289494
rect 36422 289258 43186 289494
rect 43422 289258 50186 289494
rect 50422 289258 57186 289494
rect 57422 289258 64186 289494
rect 64422 289258 71186 289494
rect 71422 289258 78186 289494
rect 78422 289258 85186 289494
rect 85422 289258 92186 289494
rect 92422 289258 99186 289494
rect 99422 289258 106186 289494
rect 106422 289258 113186 289494
rect 113422 289258 120186 289494
rect 120422 289258 127186 289494
rect 127422 289258 134186 289494
rect 134422 289258 141186 289494
rect 141422 289258 148186 289494
rect 148422 289258 155186 289494
rect 155422 289258 162186 289494
rect 162422 289258 169186 289494
rect 169422 289258 176186 289494
rect 176422 289258 183186 289494
rect 183422 289258 190186 289494
rect 190422 289258 197186 289494
rect 197422 289258 204186 289494
rect 204422 289258 211186 289494
rect 211422 289258 218186 289494
rect 218422 289258 225186 289494
rect 225422 289258 232186 289494
rect 232422 289258 239186 289494
rect 239422 289258 246186 289494
rect 246422 289258 253186 289494
rect 253422 289258 260186 289494
rect 260422 289258 267186 289494
rect 267422 289258 274186 289494
rect 274422 289258 281186 289494
rect 281422 289258 288186 289494
rect 288422 289258 295186 289494
rect 295422 289258 302186 289494
rect 302422 289258 309186 289494
rect 309422 289258 316186 289494
rect 316422 289258 323186 289494
rect 323422 289258 330186 289494
rect 330422 289258 337186 289494
rect 337422 289258 344186 289494
rect 344422 289258 351186 289494
rect 351422 289258 358186 289494
rect 358422 289258 365186 289494
rect 365422 289258 372186 289494
rect 372422 289258 379186 289494
rect 379422 289258 386186 289494
rect 386422 289258 393186 289494
rect 393422 289258 400186 289494
rect 400422 289258 407186 289494
rect 407422 289258 414186 289494
rect 414422 289258 421186 289494
rect 421422 289258 428186 289494
rect 428422 289258 435186 289494
rect 435422 289258 442186 289494
rect 442422 289258 449186 289494
rect 449422 289258 456186 289494
rect 456422 289258 463186 289494
rect 463422 289258 470186 289494
rect 470422 289258 477186 289494
rect 477422 289258 484186 289494
rect 484422 289258 491186 289494
rect 491422 289258 498186 289494
rect 498422 289258 505186 289494
rect 505422 289258 512186 289494
rect 512422 289258 519186 289494
rect 519422 289258 519952 289494
rect 520188 289258 521884 289494
rect 522120 289258 523816 289494
rect 524052 289258 525748 289494
rect 525984 289258 533186 289494
rect 533422 289258 540186 289494
rect 540422 289258 547186 289494
rect 547422 289258 554186 289494
rect 554422 289258 561186 289494
rect 561422 289258 568186 289494
rect 568422 289258 575186 289494
rect 575422 289258 582186 289494
rect 582422 289258 585818 289494
rect 586054 289258 586138 289494
rect 586374 289258 586458 289494
rect 586694 289258 586778 289494
rect 587014 289258 588874 289494
rect -4950 289216 588874 289258
rect -4950 283561 588874 283603
rect -4950 283325 -4842 283561
rect -4606 283325 -4522 283561
rect -4286 283325 -4202 283561
rect -3966 283325 -3882 283561
rect -3646 283325 2918 283561
rect 3154 283325 9918 283561
rect 10154 283325 16918 283561
rect 17154 283325 23918 283561
rect 24154 283325 30918 283561
rect 31154 283325 37918 283561
rect 38154 283325 44918 283561
rect 45154 283325 51918 283561
rect 52154 283325 58918 283561
rect 59154 283325 65918 283561
rect 66154 283325 72918 283561
rect 73154 283325 79918 283561
rect 80154 283325 86918 283561
rect 87154 283325 93918 283561
rect 94154 283325 100918 283561
rect 101154 283325 107918 283561
rect 108154 283325 114918 283561
rect 115154 283325 121918 283561
rect 122154 283325 128918 283561
rect 129154 283325 135918 283561
rect 136154 283325 142918 283561
rect 143154 283325 149918 283561
rect 150154 283325 156918 283561
rect 157154 283325 163918 283561
rect 164154 283325 170918 283561
rect 171154 283325 177918 283561
rect 178154 283325 184918 283561
rect 185154 283325 191918 283561
rect 192154 283325 198918 283561
rect 199154 283325 205918 283561
rect 206154 283325 212918 283561
rect 213154 283325 219918 283561
rect 220154 283325 226918 283561
rect 227154 283325 233918 283561
rect 234154 283325 240918 283561
rect 241154 283325 247918 283561
rect 248154 283325 254918 283561
rect 255154 283325 261918 283561
rect 262154 283325 268918 283561
rect 269154 283325 275918 283561
rect 276154 283325 282918 283561
rect 283154 283325 289918 283561
rect 290154 283325 296918 283561
rect 297154 283325 303918 283561
rect 304154 283325 310918 283561
rect 311154 283325 317918 283561
rect 318154 283325 324918 283561
rect 325154 283325 331918 283561
rect 332154 283325 338918 283561
rect 339154 283325 345918 283561
rect 346154 283325 352918 283561
rect 353154 283325 359918 283561
rect 360154 283325 366918 283561
rect 367154 283325 373918 283561
rect 374154 283325 380918 283561
rect 381154 283325 387918 283561
rect 388154 283325 394918 283561
rect 395154 283325 401918 283561
rect 402154 283325 408918 283561
rect 409154 283325 415918 283561
rect 416154 283325 422918 283561
rect 423154 283325 429918 283561
rect 430154 283325 436918 283561
rect 437154 283325 443918 283561
rect 444154 283325 450918 283561
rect 451154 283325 457918 283561
rect 458154 283325 464918 283561
rect 465154 283325 471918 283561
rect 472154 283325 478918 283561
rect 479154 283325 485918 283561
rect 486154 283325 492918 283561
rect 493154 283325 499918 283561
rect 500154 283325 506918 283561
rect 507154 283325 513918 283561
rect 514154 283325 520918 283561
rect 521154 283325 522850 283561
rect 523086 283325 524782 283561
rect 525018 283325 526714 283561
rect 526950 283325 527918 283561
rect 528154 283325 534918 283561
rect 535154 283325 541918 283561
rect 542154 283325 548918 283561
rect 549154 283325 555918 283561
rect 556154 283325 562918 283561
rect 563154 283325 569918 283561
rect 570154 283325 576918 283561
rect 577154 283325 587570 283561
rect 587806 283325 587890 283561
rect 588126 283325 588210 283561
rect 588446 283325 588530 283561
rect 588766 283325 588874 283561
rect -4950 283283 588874 283325
rect -4950 282494 588874 282536
rect -4950 282258 -3090 282494
rect -2854 282258 -2770 282494
rect -2534 282258 -2450 282494
rect -2214 282258 -2130 282494
rect -1894 282258 1186 282494
rect 1422 282258 8186 282494
rect 8422 282258 15186 282494
rect 15422 282258 22186 282494
rect 22422 282258 29186 282494
rect 29422 282258 36186 282494
rect 36422 282258 43186 282494
rect 43422 282258 50186 282494
rect 50422 282258 57186 282494
rect 57422 282258 64186 282494
rect 64422 282258 71186 282494
rect 71422 282258 78186 282494
rect 78422 282258 85186 282494
rect 85422 282258 92186 282494
rect 92422 282258 99186 282494
rect 99422 282258 106186 282494
rect 106422 282258 113186 282494
rect 113422 282258 120186 282494
rect 120422 282258 127186 282494
rect 127422 282258 134186 282494
rect 134422 282258 141186 282494
rect 141422 282258 148186 282494
rect 148422 282258 155186 282494
rect 155422 282258 162186 282494
rect 162422 282258 169186 282494
rect 169422 282258 176186 282494
rect 176422 282258 183186 282494
rect 183422 282258 190186 282494
rect 190422 282258 197186 282494
rect 197422 282258 204186 282494
rect 204422 282258 211186 282494
rect 211422 282258 218186 282494
rect 218422 282258 225186 282494
rect 225422 282258 232186 282494
rect 232422 282258 239186 282494
rect 239422 282258 246186 282494
rect 246422 282258 253186 282494
rect 253422 282258 260186 282494
rect 260422 282258 267186 282494
rect 267422 282258 274186 282494
rect 274422 282258 281186 282494
rect 281422 282258 288186 282494
rect 288422 282258 295186 282494
rect 295422 282258 302186 282494
rect 302422 282258 309186 282494
rect 309422 282258 316186 282494
rect 316422 282258 323186 282494
rect 323422 282258 330186 282494
rect 330422 282258 337186 282494
rect 337422 282258 344186 282494
rect 344422 282258 351186 282494
rect 351422 282258 358186 282494
rect 358422 282258 365186 282494
rect 365422 282258 372186 282494
rect 372422 282258 379186 282494
rect 379422 282258 386186 282494
rect 386422 282258 393186 282494
rect 393422 282258 400186 282494
rect 400422 282258 407186 282494
rect 407422 282258 414186 282494
rect 414422 282258 421186 282494
rect 421422 282258 428186 282494
rect 428422 282258 435186 282494
rect 435422 282258 442186 282494
rect 442422 282258 449186 282494
rect 449422 282258 456186 282494
rect 456422 282258 463186 282494
rect 463422 282258 470186 282494
rect 470422 282258 477186 282494
rect 477422 282258 484186 282494
rect 484422 282258 491186 282494
rect 491422 282258 498186 282494
rect 498422 282258 505186 282494
rect 505422 282258 512186 282494
rect 512422 282258 519186 282494
rect 519422 282258 519952 282494
rect 520188 282258 521884 282494
rect 522120 282258 523816 282494
rect 524052 282258 525748 282494
rect 525984 282258 533186 282494
rect 533422 282258 540186 282494
rect 540422 282258 547186 282494
rect 547422 282258 554186 282494
rect 554422 282258 561186 282494
rect 561422 282258 568186 282494
rect 568422 282258 575186 282494
rect 575422 282258 582186 282494
rect 582422 282258 585818 282494
rect 586054 282258 586138 282494
rect 586374 282258 586458 282494
rect 586694 282258 586778 282494
rect 587014 282258 588874 282494
rect -4950 282216 588874 282258
rect -4950 276561 588874 276603
rect -4950 276325 -4842 276561
rect -4606 276325 -4522 276561
rect -4286 276325 -4202 276561
rect -3966 276325 -3882 276561
rect -3646 276325 2918 276561
rect 3154 276325 9918 276561
rect 10154 276325 16918 276561
rect 17154 276325 23918 276561
rect 24154 276325 30918 276561
rect 31154 276325 37918 276561
rect 38154 276325 44918 276561
rect 45154 276325 51918 276561
rect 52154 276325 58918 276561
rect 59154 276325 65918 276561
rect 66154 276325 72918 276561
rect 73154 276325 79918 276561
rect 80154 276325 86918 276561
rect 87154 276325 93918 276561
rect 94154 276325 100918 276561
rect 101154 276325 107918 276561
rect 108154 276325 114918 276561
rect 115154 276325 121918 276561
rect 122154 276325 128918 276561
rect 129154 276325 135918 276561
rect 136154 276325 142918 276561
rect 143154 276325 149918 276561
rect 150154 276325 156918 276561
rect 157154 276325 163918 276561
rect 164154 276325 170918 276561
rect 171154 276325 177918 276561
rect 178154 276325 184918 276561
rect 185154 276325 191918 276561
rect 192154 276325 198918 276561
rect 199154 276325 205918 276561
rect 206154 276325 212918 276561
rect 213154 276325 219918 276561
rect 220154 276325 226918 276561
rect 227154 276325 233918 276561
rect 234154 276325 240918 276561
rect 241154 276325 247918 276561
rect 248154 276325 254918 276561
rect 255154 276325 261918 276561
rect 262154 276325 268918 276561
rect 269154 276325 275918 276561
rect 276154 276325 282918 276561
rect 283154 276325 289918 276561
rect 290154 276325 296918 276561
rect 297154 276325 303918 276561
rect 304154 276325 310918 276561
rect 311154 276325 317918 276561
rect 318154 276325 324918 276561
rect 325154 276325 331918 276561
rect 332154 276325 338918 276561
rect 339154 276325 345918 276561
rect 346154 276325 352918 276561
rect 353154 276325 359918 276561
rect 360154 276325 366918 276561
rect 367154 276325 373918 276561
rect 374154 276325 380918 276561
rect 381154 276325 387918 276561
rect 388154 276325 394918 276561
rect 395154 276325 401918 276561
rect 402154 276325 408918 276561
rect 409154 276325 415918 276561
rect 416154 276325 422918 276561
rect 423154 276325 429918 276561
rect 430154 276325 436918 276561
rect 437154 276325 443918 276561
rect 444154 276325 450918 276561
rect 451154 276325 457918 276561
rect 458154 276325 464918 276561
rect 465154 276325 471918 276561
rect 472154 276325 478918 276561
rect 479154 276325 485918 276561
rect 486154 276325 492918 276561
rect 493154 276325 499918 276561
rect 500154 276325 506918 276561
rect 507154 276325 513918 276561
rect 514154 276325 520918 276561
rect 521154 276325 527918 276561
rect 528154 276325 534918 276561
rect 535154 276325 541918 276561
rect 542154 276325 548918 276561
rect 549154 276325 555918 276561
rect 556154 276325 562918 276561
rect 563154 276325 569918 276561
rect 570154 276325 576918 276561
rect 577154 276325 587570 276561
rect 587806 276325 587890 276561
rect 588126 276325 588210 276561
rect 588446 276325 588530 276561
rect 588766 276325 588874 276561
rect -4950 276283 588874 276325
rect -4950 275494 588874 275536
rect -4950 275258 -3090 275494
rect -2854 275258 -2770 275494
rect -2534 275258 -2450 275494
rect -2214 275258 -2130 275494
rect -1894 275258 1186 275494
rect 1422 275258 8186 275494
rect 8422 275258 15186 275494
rect 15422 275258 22186 275494
rect 22422 275258 29186 275494
rect 29422 275258 36186 275494
rect 36422 275258 43186 275494
rect 43422 275258 50186 275494
rect 50422 275258 57186 275494
rect 57422 275258 64186 275494
rect 64422 275258 71186 275494
rect 71422 275258 78186 275494
rect 78422 275258 85186 275494
rect 85422 275258 92186 275494
rect 92422 275258 99186 275494
rect 99422 275258 106186 275494
rect 106422 275258 113186 275494
rect 113422 275258 120186 275494
rect 120422 275258 127186 275494
rect 127422 275258 134186 275494
rect 134422 275258 141186 275494
rect 141422 275258 148186 275494
rect 148422 275258 155186 275494
rect 155422 275258 162186 275494
rect 162422 275258 169186 275494
rect 169422 275258 176186 275494
rect 176422 275258 183186 275494
rect 183422 275258 190186 275494
rect 190422 275258 197186 275494
rect 197422 275258 204186 275494
rect 204422 275258 211186 275494
rect 211422 275258 218186 275494
rect 218422 275258 225186 275494
rect 225422 275258 232186 275494
rect 232422 275258 239186 275494
rect 239422 275258 246186 275494
rect 246422 275258 253186 275494
rect 253422 275258 260186 275494
rect 260422 275258 267186 275494
rect 267422 275258 274186 275494
rect 274422 275258 281186 275494
rect 281422 275258 288186 275494
rect 288422 275258 295186 275494
rect 295422 275258 302186 275494
rect 302422 275258 309186 275494
rect 309422 275258 316186 275494
rect 316422 275258 323186 275494
rect 323422 275258 330186 275494
rect 330422 275258 337186 275494
rect 337422 275258 344186 275494
rect 344422 275258 351186 275494
rect 351422 275258 358186 275494
rect 358422 275258 365186 275494
rect 365422 275258 372186 275494
rect 372422 275258 379186 275494
rect 379422 275258 386186 275494
rect 386422 275258 393186 275494
rect 393422 275258 400186 275494
rect 400422 275258 407186 275494
rect 407422 275258 414186 275494
rect 414422 275258 421186 275494
rect 421422 275258 428186 275494
rect 428422 275258 435186 275494
rect 435422 275258 442186 275494
rect 442422 275258 449186 275494
rect 449422 275258 456186 275494
rect 456422 275258 463186 275494
rect 463422 275258 470186 275494
rect 470422 275258 477186 275494
rect 477422 275258 484186 275494
rect 484422 275258 491186 275494
rect 491422 275258 498186 275494
rect 498422 275258 505186 275494
rect 505422 275258 512186 275494
rect 512422 275258 519186 275494
rect 519422 275258 526186 275494
rect 526422 275258 533186 275494
rect 533422 275258 540186 275494
rect 540422 275258 547186 275494
rect 547422 275258 554186 275494
rect 554422 275258 561186 275494
rect 561422 275258 568186 275494
rect 568422 275258 575186 275494
rect 575422 275258 582186 275494
rect 582422 275258 585818 275494
rect 586054 275258 586138 275494
rect 586374 275258 586458 275494
rect 586694 275258 586778 275494
rect 587014 275258 588874 275494
rect -4950 275216 588874 275258
rect -4950 269561 588874 269603
rect -4950 269325 -4842 269561
rect -4606 269325 -4522 269561
rect -4286 269325 -4202 269561
rect -3966 269325 -3882 269561
rect -3646 269325 2918 269561
rect 3154 269325 9918 269561
rect 10154 269325 16918 269561
rect 17154 269325 23918 269561
rect 24154 269325 30918 269561
rect 31154 269325 37918 269561
rect 38154 269325 44918 269561
rect 45154 269325 51918 269561
rect 52154 269325 58918 269561
rect 59154 269325 65918 269561
rect 66154 269325 72918 269561
rect 73154 269325 79918 269561
rect 80154 269325 86918 269561
rect 87154 269325 93918 269561
rect 94154 269325 100918 269561
rect 101154 269325 107918 269561
rect 108154 269325 114918 269561
rect 115154 269325 121918 269561
rect 122154 269325 128918 269561
rect 129154 269325 135918 269561
rect 136154 269325 142918 269561
rect 143154 269325 149918 269561
rect 150154 269325 156918 269561
rect 157154 269325 163918 269561
rect 164154 269325 170918 269561
rect 171154 269325 177918 269561
rect 178154 269325 184918 269561
rect 185154 269325 191918 269561
rect 192154 269325 198918 269561
rect 199154 269325 205918 269561
rect 206154 269325 212918 269561
rect 213154 269325 219918 269561
rect 220154 269325 226918 269561
rect 227154 269325 233918 269561
rect 234154 269325 240918 269561
rect 241154 269325 247918 269561
rect 248154 269325 254918 269561
rect 255154 269325 261918 269561
rect 262154 269325 268918 269561
rect 269154 269325 275918 269561
rect 276154 269325 282918 269561
rect 283154 269325 289918 269561
rect 290154 269325 296918 269561
rect 297154 269325 303918 269561
rect 304154 269325 310918 269561
rect 311154 269325 317918 269561
rect 318154 269325 324918 269561
rect 325154 269325 331918 269561
rect 332154 269325 338918 269561
rect 339154 269325 345918 269561
rect 346154 269325 352918 269561
rect 353154 269325 359918 269561
rect 360154 269325 366918 269561
rect 367154 269325 373918 269561
rect 374154 269325 380918 269561
rect 381154 269325 387918 269561
rect 388154 269325 394918 269561
rect 395154 269325 401918 269561
rect 402154 269325 408918 269561
rect 409154 269325 415918 269561
rect 416154 269325 422918 269561
rect 423154 269325 429918 269561
rect 430154 269325 436918 269561
rect 437154 269325 443918 269561
rect 444154 269325 450918 269561
rect 451154 269325 457918 269561
rect 458154 269325 464918 269561
rect 465154 269325 471918 269561
rect 472154 269325 478918 269561
rect 479154 269325 485918 269561
rect 486154 269325 492918 269561
rect 493154 269325 499918 269561
rect 500154 269325 506918 269561
rect 507154 269325 513918 269561
rect 514154 269325 520918 269561
rect 521154 269325 527918 269561
rect 528154 269325 534918 269561
rect 535154 269325 541918 269561
rect 542154 269325 548918 269561
rect 549154 269325 555918 269561
rect 556154 269325 562918 269561
rect 563154 269325 569918 269561
rect 570154 269325 576918 269561
rect 577154 269325 587570 269561
rect 587806 269325 587890 269561
rect 588126 269325 588210 269561
rect 588446 269325 588530 269561
rect 588766 269325 588874 269561
rect -4950 269283 588874 269325
rect -4950 268494 588874 268536
rect -4950 268258 -3090 268494
rect -2854 268258 -2770 268494
rect -2534 268258 -2450 268494
rect -2214 268258 -2130 268494
rect -1894 268258 1186 268494
rect 1422 268258 8186 268494
rect 8422 268258 15186 268494
rect 15422 268258 22186 268494
rect 22422 268258 29186 268494
rect 29422 268258 36186 268494
rect 36422 268258 43186 268494
rect 43422 268258 50186 268494
rect 50422 268258 57186 268494
rect 57422 268258 64186 268494
rect 64422 268258 71186 268494
rect 71422 268258 78186 268494
rect 78422 268258 85186 268494
rect 85422 268258 92186 268494
rect 92422 268258 99186 268494
rect 99422 268258 106186 268494
rect 106422 268258 113186 268494
rect 113422 268258 120186 268494
rect 120422 268258 127186 268494
rect 127422 268258 134186 268494
rect 134422 268258 141186 268494
rect 141422 268258 148186 268494
rect 148422 268258 155186 268494
rect 155422 268258 162186 268494
rect 162422 268258 169186 268494
rect 169422 268258 176186 268494
rect 176422 268258 183186 268494
rect 183422 268258 190186 268494
rect 190422 268258 197186 268494
rect 197422 268258 204186 268494
rect 204422 268258 211186 268494
rect 211422 268258 218186 268494
rect 218422 268258 225186 268494
rect 225422 268258 232186 268494
rect 232422 268258 239186 268494
rect 239422 268258 246186 268494
rect 246422 268258 253186 268494
rect 253422 268258 260186 268494
rect 260422 268258 267186 268494
rect 267422 268258 274186 268494
rect 274422 268258 281186 268494
rect 281422 268258 288186 268494
rect 288422 268258 295186 268494
rect 295422 268258 302186 268494
rect 302422 268258 309186 268494
rect 309422 268258 316186 268494
rect 316422 268258 323186 268494
rect 323422 268258 330186 268494
rect 330422 268258 337186 268494
rect 337422 268258 344186 268494
rect 344422 268258 351186 268494
rect 351422 268258 358186 268494
rect 358422 268258 365186 268494
rect 365422 268258 372186 268494
rect 372422 268258 379186 268494
rect 379422 268258 386186 268494
rect 386422 268258 393186 268494
rect 393422 268258 400186 268494
rect 400422 268258 407186 268494
rect 407422 268258 414186 268494
rect 414422 268258 421186 268494
rect 421422 268258 428186 268494
rect 428422 268258 435186 268494
rect 435422 268258 442186 268494
rect 442422 268258 449186 268494
rect 449422 268258 456186 268494
rect 456422 268258 463186 268494
rect 463422 268258 470186 268494
rect 470422 268258 477186 268494
rect 477422 268258 484186 268494
rect 484422 268258 491186 268494
rect 491422 268258 498186 268494
rect 498422 268258 505186 268494
rect 505422 268258 512186 268494
rect 512422 268258 519186 268494
rect 519422 268258 526186 268494
rect 526422 268258 533186 268494
rect 533422 268258 540186 268494
rect 540422 268258 547186 268494
rect 547422 268258 554186 268494
rect 554422 268258 561186 268494
rect 561422 268258 568186 268494
rect 568422 268258 575186 268494
rect 575422 268258 582186 268494
rect 582422 268258 585818 268494
rect 586054 268258 586138 268494
rect 586374 268258 586458 268494
rect 586694 268258 586778 268494
rect 587014 268258 588874 268494
rect -4950 268216 588874 268258
rect -4950 262561 588874 262603
rect -4950 262325 -4842 262561
rect -4606 262325 -4522 262561
rect -4286 262325 -4202 262561
rect -3966 262325 -3882 262561
rect -3646 262325 2918 262561
rect 3154 262325 9918 262561
rect 10154 262325 16918 262561
rect 17154 262325 23918 262561
rect 24154 262325 30918 262561
rect 31154 262325 37918 262561
rect 38154 262325 44918 262561
rect 45154 262325 51918 262561
rect 52154 262325 58918 262561
rect 59154 262325 65918 262561
rect 66154 262325 72918 262561
rect 73154 262325 79918 262561
rect 80154 262325 86918 262561
rect 87154 262325 93918 262561
rect 94154 262325 100918 262561
rect 101154 262325 107918 262561
rect 108154 262325 114918 262561
rect 115154 262325 121918 262561
rect 122154 262325 128918 262561
rect 129154 262325 135918 262561
rect 136154 262325 142918 262561
rect 143154 262325 149918 262561
rect 150154 262325 156918 262561
rect 157154 262325 163918 262561
rect 164154 262325 170918 262561
rect 171154 262325 177918 262561
rect 178154 262325 184918 262561
rect 185154 262325 191918 262561
rect 192154 262325 198918 262561
rect 199154 262325 205918 262561
rect 206154 262325 212918 262561
rect 213154 262325 219918 262561
rect 220154 262325 226918 262561
rect 227154 262325 233918 262561
rect 234154 262325 240918 262561
rect 241154 262325 247918 262561
rect 248154 262325 254918 262561
rect 255154 262325 261918 262561
rect 262154 262325 268918 262561
rect 269154 262325 275918 262561
rect 276154 262325 282918 262561
rect 283154 262325 289918 262561
rect 290154 262325 296918 262561
rect 297154 262325 303918 262561
rect 304154 262325 310918 262561
rect 311154 262325 317918 262561
rect 318154 262325 324918 262561
rect 325154 262325 331918 262561
rect 332154 262325 338918 262561
rect 339154 262325 345918 262561
rect 346154 262325 352918 262561
rect 353154 262325 359918 262561
rect 360154 262325 366918 262561
rect 367154 262325 373918 262561
rect 374154 262325 380918 262561
rect 381154 262325 387918 262561
rect 388154 262325 394918 262561
rect 395154 262325 401918 262561
rect 402154 262325 408918 262561
rect 409154 262325 415918 262561
rect 416154 262325 422918 262561
rect 423154 262325 429918 262561
rect 430154 262325 436918 262561
rect 437154 262325 443918 262561
rect 444154 262325 450918 262561
rect 451154 262325 457918 262561
rect 458154 262325 464918 262561
rect 465154 262325 471918 262561
rect 472154 262325 478918 262561
rect 479154 262325 485918 262561
rect 486154 262325 492918 262561
rect 493154 262325 499918 262561
rect 500154 262325 506918 262561
rect 507154 262325 513918 262561
rect 514154 262325 520918 262561
rect 521154 262325 527918 262561
rect 528154 262325 534918 262561
rect 535154 262325 541918 262561
rect 542154 262325 548918 262561
rect 549154 262325 555918 262561
rect 556154 262325 562918 262561
rect 563154 262325 569918 262561
rect 570154 262325 576918 262561
rect 577154 262325 587570 262561
rect 587806 262325 587890 262561
rect 588126 262325 588210 262561
rect 588446 262325 588530 262561
rect 588766 262325 588874 262561
rect -4950 262283 588874 262325
rect -4950 261494 588874 261536
rect -4950 261258 -3090 261494
rect -2854 261258 -2770 261494
rect -2534 261258 -2450 261494
rect -2214 261258 -2130 261494
rect -1894 261258 1186 261494
rect 1422 261258 8186 261494
rect 8422 261258 15186 261494
rect 15422 261258 22186 261494
rect 22422 261258 29186 261494
rect 29422 261258 36186 261494
rect 36422 261258 43186 261494
rect 43422 261258 50186 261494
rect 50422 261258 57186 261494
rect 57422 261258 64186 261494
rect 64422 261258 71186 261494
rect 71422 261258 78186 261494
rect 78422 261258 85186 261494
rect 85422 261258 92186 261494
rect 92422 261258 99186 261494
rect 99422 261258 106186 261494
rect 106422 261258 113186 261494
rect 113422 261258 120186 261494
rect 120422 261258 127186 261494
rect 127422 261258 134186 261494
rect 134422 261258 141186 261494
rect 141422 261258 148186 261494
rect 148422 261258 155186 261494
rect 155422 261258 162186 261494
rect 162422 261258 169186 261494
rect 169422 261258 176186 261494
rect 176422 261258 183186 261494
rect 183422 261258 190186 261494
rect 190422 261258 197186 261494
rect 197422 261258 204186 261494
rect 204422 261258 211186 261494
rect 211422 261258 218186 261494
rect 218422 261258 225186 261494
rect 225422 261258 232186 261494
rect 232422 261258 239186 261494
rect 239422 261258 246186 261494
rect 246422 261258 253186 261494
rect 253422 261258 260186 261494
rect 260422 261258 267186 261494
rect 267422 261258 274186 261494
rect 274422 261258 281186 261494
rect 281422 261258 288186 261494
rect 288422 261258 295186 261494
rect 295422 261258 302186 261494
rect 302422 261258 309186 261494
rect 309422 261258 316186 261494
rect 316422 261258 323186 261494
rect 323422 261258 330186 261494
rect 330422 261258 337186 261494
rect 337422 261258 344186 261494
rect 344422 261258 351186 261494
rect 351422 261258 358186 261494
rect 358422 261258 365186 261494
rect 365422 261258 372186 261494
rect 372422 261258 379186 261494
rect 379422 261258 386186 261494
rect 386422 261258 393186 261494
rect 393422 261258 400186 261494
rect 400422 261258 407186 261494
rect 407422 261258 414186 261494
rect 414422 261258 421186 261494
rect 421422 261258 428186 261494
rect 428422 261258 435186 261494
rect 435422 261258 442186 261494
rect 442422 261258 449186 261494
rect 449422 261258 456186 261494
rect 456422 261258 463186 261494
rect 463422 261258 470186 261494
rect 470422 261258 477186 261494
rect 477422 261258 484186 261494
rect 484422 261258 491186 261494
rect 491422 261258 498186 261494
rect 498422 261258 505186 261494
rect 505422 261258 512186 261494
rect 512422 261258 519186 261494
rect 519422 261258 533186 261494
rect 533422 261258 540186 261494
rect 540422 261258 547186 261494
rect 547422 261258 554186 261494
rect 554422 261258 561186 261494
rect 561422 261258 568186 261494
rect 568422 261258 575186 261494
rect 575422 261258 582186 261494
rect 582422 261258 585818 261494
rect 586054 261258 586138 261494
rect 586374 261258 586458 261494
rect 586694 261258 586778 261494
rect 587014 261258 588874 261494
rect -4950 261216 588874 261258
rect -4950 255561 588874 255603
rect -4950 255325 -4842 255561
rect -4606 255325 -4522 255561
rect -4286 255325 -4202 255561
rect -3966 255325 -3882 255561
rect -3646 255325 2918 255561
rect 3154 255325 9918 255561
rect 10154 255325 16918 255561
rect 17154 255325 23918 255561
rect 24154 255325 30918 255561
rect 31154 255325 37918 255561
rect 38154 255325 44918 255561
rect 45154 255325 51918 255561
rect 52154 255325 58918 255561
rect 59154 255325 65918 255561
rect 66154 255325 72918 255561
rect 73154 255325 79918 255561
rect 80154 255325 86918 255561
rect 87154 255325 93918 255561
rect 94154 255325 100918 255561
rect 101154 255325 107918 255561
rect 108154 255325 114918 255561
rect 115154 255325 121918 255561
rect 122154 255325 128918 255561
rect 129154 255325 135918 255561
rect 136154 255325 142918 255561
rect 143154 255325 149918 255561
rect 150154 255325 156918 255561
rect 157154 255325 163918 255561
rect 164154 255325 170918 255561
rect 171154 255325 177918 255561
rect 178154 255325 184918 255561
rect 185154 255325 191918 255561
rect 192154 255325 198918 255561
rect 199154 255325 205918 255561
rect 206154 255325 212918 255561
rect 213154 255325 219918 255561
rect 220154 255325 226918 255561
rect 227154 255325 233918 255561
rect 234154 255325 240918 255561
rect 241154 255325 247918 255561
rect 248154 255325 254918 255561
rect 255154 255325 261918 255561
rect 262154 255325 268918 255561
rect 269154 255325 275918 255561
rect 276154 255325 282918 255561
rect 283154 255325 289918 255561
rect 290154 255325 296918 255561
rect 297154 255325 303918 255561
rect 304154 255325 310918 255561
rect 311154 255325 317918 255561
rect 318154 255325 324918 255561
rect 325154 255325 331918 255561
rect 332154 255325 338918 255561
rect 339154 255325 345918 255561
rect 346154 255325 352918 255561
rect 353154 255325 359918 255561
rect 360154 255325 366918 255561
rect 367154 255325 373918 255561
rect 374154 255325 380918 255561
rect 381154 255325 387918 255561
rect 388154 255325 394918 255561
rect 395154 255325 401918 255561
rect 402154 255325 408918 255561
rect 409154 255325 415918 255561
rect 416154 255325 422918 255561
rect 423154 255325 429918 255561
rect 430154 255325 436918 255561
rect 437154 255325 443918 255561
rect 444154 255325 450918 255561
rect 451154 255325 457918 255561
rect 458154 255325 464918 255561
rect 465154 255325 471918 255561
rect 472154 255325 478918 255561
rect 479154 255325 485918 255561
rect 486154 255325 492918 255561
rect 493154 255325 499918 255561
rect 500154 255325 506918 255561
rect 507154 255325 513918 255561
rect 514154 255325 520918 255561
rect 521154 255325 522850 255561
rect 523086 255325 524782 255561
rect 525018 255325 526714 255561
rect 526950 255325 527918 255561
rect 528154 255325 534918 255561
rect 535154 255325 541918 255561
rect 542154 255325 548918 255561
rect 549154 255325 555918 255561
rect 556154 255325 562918 255561
rect 563154 255325 569918 255561
rect 570154 255325 576918 255561
rect 577154 255325 587570 255561
rect 587806 255325 587890 255561
rect 588126 255325 588210 255561
rect 588446 255325 588530 255561
rect 588766 255325 588874 255561
rect -4950 255283 588874 255325
rect -4950 254494 588874 254536
rect -4950 254258 -3090 254494
rect -2854 254258 -2770 254494
rect -2534 254258 -2450 254494
rect -2214 254258 -2130 254494
rect -1894 254258 1186 254494
rect 1422 254258 8186 254494
rect 8422 254258 15186 254494
rect 15422 254258 22186 254494
rect 22422 254258 29186 254494
rect 29422 254258 36186 254494
rect 36422 254258 43186 254494
rect 43422 254258 50186 254494
rect 50422 254258 57186 254494
rect 57422 254258 64186 254494
rect 64422 254258 71186 254494
rect 71422 254258 78186 254494
rect 78422 254258 85186 254494
rect 85422 254258 92186 254494
rect 92422 254258 99186 254494
rect 99422 254258 106186 254494
rect 106422 254258 113186 254494
rect 113422 254258 120186 254494
rect 120422 254258 127186 254494
rect 127422 254258 134186 254494
rect 134422 254258 141186 254494
rect 141422 254258 148186 254494
rect 148422 254258 155186 254494
rect 155422 254258 162186 254494
rect 162422 254258 169186 254494
rect 169422 254258 176186 254494
rect 176422 254258 183186 254494
rect 183422 254258 190186 254494
rect 190422 254258 197186 254494
rect 197422 254258 204186 254494
rect 204422 254258 211186 254494
rect 211422 254258 218186 254494
rect 218422 254258 225186 254494
rect 225422 254258 232186 254494
rect 232422 254258 239186 254494
rect 239422 254258 246186 254494
rect 246422 254258 253186 254494
rect 253422 254258 260186 254494
rect 260422 254258 267186 254494
rect 267422 254258 274186 254494
rect 274422 254258 281186 254494
rect 281422 254258 288186 254494
rect 288422 254258 295186 254494
rect 295422 254258 302186 254494
rect 302422 254258 309186 254494
rect 309422 254258 316186 254494
rect 316422 254258 323186 254494
rect 323422 254258 330186 254494
rect 330422 254258 337186 254494
rect 337422 254258 344186 254494
rect 344422 254258 351186 254494
rect 351422 254258 358186 254494
rect 358422 254258 365186 254494
rect 365422 254258 372186 254494
rect 372422 254258 379186 254494
rect 379422 254258 386186 254494
rect 386422 254258 393186 254494
rect 393422 254258 400186 254494
rect 400422 254258 407186 254494
rect 407422 254258 414186 254494
rect 414422 254258 421186 254494
rect 421422 254258 428186 254494
rect 428422 254258 435186 254494
rect 435422 254258 442186 254494
rect 442422 254258 449186 254494
rect 449422 254258 456186 254494
rect 456422 254258 463186 254494
rect 463422 254258 470186 254494
rect 470422 254258 477186 254494
rect 477422 254258 484186 254494
rect 484422 254258 491186 254494
rect 491422 254258 498186 254494
rect 498422 254258 505186 254494
rect 505422 254258 512186 254494
rect 512422 254258 519186 254494
rect 519422 254258 519952 254494
rect 520188 254258 521884 254494
rect 522120 254258 523816 254494
rect 524052 254258 525748 254494
rect 525984 254258 533186 254494
rect 533422 254258 540186 254494
rect 540422 254258 547186 254494
rect 547422 254258 554186 254494
rect 554422 254258 561186 254494
rect 561422 254258 568186 254494
rect 568422 254258 575186 254494
rect 575422 254258 582186 254494
rect 582422 254258 585818 254494
rect 586054 254258 586138 254494
rect 586374 254258 586458 254494
rect 586694 254258 586778 254494
rect 587014 254258 588874 254494
rect -4950 254216 588874 254258
rect -4950 248561 588874 248603
rect -4950 248325 -4842 248561
rect -4606 248325 -4522 248561
rect -4286 248325 -4202 248561
rect -3966 248325 -3882 248561
rect -3646 248325 2918 248561
rect 3154 248325 9918 248561
rect 10154 248325 16918 248561
rect 17154 248325 23918 248561
rect 24154 248325 30918 248561
rect 31154 248325 37918 248561
rect 38154 248325 44918 248561
rect 45154 248325 51918 248561
rect 52154 248325 58918 248561
rect 59154 248325 65918 248561
rect 66154 248325 72918 248561
rect 73154 248325 79918 248561
rect 80154 248325 86918 248561
rect 87154 248325 93918 248561
rect 94154 248325 100918 248561
rect 101154 248325 107918 248561
rect 108154 248325 114918 248561
rect 115154 248325 121918 248561
rect 122154 248325 128918 248561
rect 129154 248325 135918 248561
rect 136154 248325 142918 248561
rect 143154 248325 149918 248561
rect 150154 248325 156918 248561
rect 157154 248325 163918 248561
rect 164154 248325 170918 248561
rect 171154 248325 177918 248561
rect 178154 248325 184918 248561
rect 185154 248325 191918 248561
rect 192154 248325 198918 248561
rect 199154 248325 205918 248561
rect 206154 248325 212918 248561
rect 213154 248325 219918 248561
rect 220154 248325 226918 248561
rect 227154 248325 233918 248561
rect 234154 248325 240918 248561
rect 241154 248325 247918 248561
rect 248154 248325 254918 248561
rect 255154 248325 261918 248561
rect 262154 248325 268918 248561
rect 269154 248325 275918 248561
rect 276154 248325 282918 248561
rect 283154 248325 289918 248561
rect 290154 248325 296918 248561
rect 297154 248325 303918 248561
rect 304154 248325 310918 248561
rect 311154 248325 317918 248561
rect 318154 248325 324918 248561
rect 325154 248325 331918 248561
rect 332154 248325 338918 248561
rect 339154 248325 345918 248561
rect 346154 248325 352918 248561
rect 353154 248325 359918 248561
rect 360154 248325 366918 248561
rect 367154 248325 373918 248561
rect 374154 248325 380918 248561
rect 381154 248325 387918 248561
rect 388154 248325 394918 248561
rect 395154 248325 401918 248561
rect 402154 248325 408918 248561
rect 409154 248325 415918 248561
rect 416154 248325 422918 248561
rect 423154 248325 429918 248561
rect 430154 248325 436918 248561
rect 437154 248325 443918 248561
rect 444154 248325 450918 248561
rect 451154 248325 457918 248561
rect 458154 248325 464918 248561
rect 465154 248325 471918 248561
rect 472154 248325 478918 248561
rect 479154 248325 485918 248561
rect 486154 248325 492918 248561
rect 493154 248325 499918 248561
rect 500154 248325 506918 248561
rect 507154 248325 513918 248561
rect 514154 248325 520918 248561
rect 521154 248325 522850 248561
rect 523086 248325 524782 248561
rect 525018 248325 526714 248561
rect 526950 248325 527918 248561
rect 528154 248325 534918 248561
rect 535154 248325 541918 248561
rect 542154 248325 548918 248561
rect 549154 248325 555918 248561
rect 556154 248325 562918 248561
rect 563154 248325 569918 248561
rect 570154 248325 576918 248561
rect 577154 248325 587570 248561
rect 587806 248325 587890 248561
rect 588126 248325 588210 248561
rect 588446 248325 588530 248561
rect 588766 248325 588874 248561
rect -4950 248283 588874 248325
rect -4950 247494 588874 247536
rect -4950 247258 -3090 247494
rect -2854 247258 -2770 247494
rect -2534 247258 -2450 247494
rect -2214 247258 -2130 247494
rect -1894 247258 1186 247494
rect 1422 247258 8186 247494
rect 8422 247258 15186 247494
rect 15422 247258 22186 247494
rect 22422 247258 29186 247494
rect 29422 247258 36186 247494
rect 36422 247258 43186 247494
rect 43422 247258 50186 247494
rect 50422 247258 57186 247494
rect 57422 247258 64186 247494
rect 64422 247258 71186 247494
rect 71422 247258 78186 247494
rect 78422 247258 85186 247494
rect 85422 247258 92186 247494
rect 92422 247258 99186 247494
rect 99422 247258 106186 247494
rect 106422 247258 113186 247494
rect 113422 247258 120186 247494
rect 120422 247258 127186 247494
rect 127422 247258 134186 247494
rect 134422 247258 141186 247494
rect 141422 247258 148186 247494
rect 148422 247258 155186 247494
rect 155422 247258 162186 247494
rect 162422 247258 169186 247494
rect 169422 247258 176186 247494
rect 176422 247258 183186 247494
rect 183422 247258 190186 247494
rect 190422 247258 197186 247494
rect 197422 247258 204186 247494
rect 204422 247258 211186 247494
rect 211422 247258 218186 247494
rect 218422 247258 225186 247494
rect 225422 247258 232186 247494
rect 232422 247258 239186 247494
rect 239422 247258 246186 247494
rect 246422 247258 253186 247494
rect 253422 247258 260186 247494
rect 260422 247258 267186 247494
rect 267422 247258 274186 247494
rect 274422 247258 281186 247494
rect 281422 247258 288186 247494
rect 288422 247258 295186 247494
rect 295422 247258 302186 247494
rect 302422 247258 309186 247494
rect 309422 247258 316186 247494
rect 316422 247258 323186 247494
rect 323422 247258 330186 247494
rect 330422 247258 337186 247494
rect 337422 247258 344186 247494
rect 344422 247258 351186 247494
rect 351422 247258 358186 247494
rect 358422 247258 365186 247494
rect 365422 247258 372186 247494
rect 372422 247258 379186 247494
rect 379422 247258 386186 247494
rect 386422 247258 393186 247494
rect 393422 247258 400186 247494
rect 400422 247258 407186 247494
rect 407422 247258 414186 247494
rect 414422 247258 421186 247494
rect 421422 247258 428186 247494
rect 428422 247258 435186 247494
rect 435422 247258 442186 247494
rect 442422 247258 449186 247494
rect 449422 247258 456186 247494
rect 456422 247258 463186 247494
rect 463422 247258 470186 247494
rect 470422 247258 477186 247494
rect 477422 247258 484186 247494
rect 484422 247258 491186 247494
rect 491422 247258 498186 247494
rect 498422 247258 505186 247494
rect 505422 247258 512186 247494
rect 512422 247258 519186 247494
rect 519422 247258 519952 247494
rect 520188 247258 521884 247494
rect 522120 247258 523816 247494
rect 524052 247258 525748 247494
rect 525984 247258 533186 247494
rect 533422 247258 540186 247494
rect 540422 247258 547186 247494
rect 547422 247258 554186 247494
rect 554422 247258 561186 247494
rect 561422 247258 568186 247494
rect 568422 247258 575186 247494
rect 575422 247258 582186 247494
rect 582422 247258 585818 247494
rect 586054 247258 586138 247494
rect 586374 247258 586458 247494
rect 586694 247258 586778 247494
rect 587014 247258 588874 247494
rect -4950 247216 588874 247258
rect -4950 241561 588874 241603
rect -4950 241325 -4842 241561
rect -4606 241325 -4522 241561
rect -4286 241325 -4202 241561
rect -3966 241325 -3882 241561
rect -3646 241325 2918 241561
rect 3154 241325 9918 241561
rect 10154 241325 16918 241561
rect 17154 241325 23918 241561
rect 24154 241325 30918 241561
rect 31154 241325 37918 241561
rect 38154 241325 44918 241561
rect 45154 241325 51918 241561
rect 52154 241325 58918 241561
rect 59154 241325 65918 241561
rect 66154 241325 72918 241561
rect 73154 241325 79918 241561
rect 80154 241325 86918 241561
rect 87154 241325 93918 241561
rect 94154 241325 100918 241561
rect 101154 241325 107918 241561
rect 108154 241325 114918 241561
rect 115154 241325 121918 241561
rect 122154 241325 128918 241561
rect 129154 241325 135918 241561
rect 136154 241325 142918 241561
rect 143154 241325 149918 241561
rect 150154 241325 156918 241561
rect 157154 241325 163918 241561
rect 164154 241325 170918 241561
rect 171154 241325 177918 241561
rect 178154 241325 184918 241561
rect 185154 241325 191918 241561
rect 192154 241325 198918 241561
rect 199154 241325 205918 241561
rect 206154 241325 212918 241561
rect 213154 241325 219918 241561
rect 220154 241325 226918 241561
rect 227154 241325 233918 241561
rect 234154 241325 240918 241561
rect 241154 241325 247918 241561
rect 248154 241325 254918 241561
rect 255154 241325 261918 241561
rect 262154 241325 268918 241561
rect 269154 241325 275918 241561
rect 276154 241325 282918 241561
rect 283154 241325 289918 241561
rect 290154 241325 296918 241561
rect 297154 241325 303918 241561
rect 304154 241325 310918 241561
rect 311154 241325 317918 241561
rect 318154 241325 324918 241561
rect 325154 241325 331918 241561
rect 332154 241325 338918 241561
rect 339154 241325 345918 241561
rect 346154 241325 352918 241561
rect 353154 241325 359918 241561
rect 360154 241325 366918 241561
rect 367154 241325 373918 241561
rect 374154 241325 380918 241561
rect 381154 241325 387918 241561
rect 388154 241325 394918 241561
rect 395154 241325 401918 241561
rect 402154 241325 408918 241561
rect 409154 241325 415918 241561
rect 416154 241325 422918 241561
rect 423154 241325 429918 241561
rect 430154 241325 436918 241561
rect 437154 241325 443918 241561
rect 444154 241325 450918 241561
rect 451154 241325 457918 241561
rect 458154 241325 464918 241561
rect 465154 241325 471918 241561
rect 472154 241325 478918 241561
rect 479154 241325 485918 241561
rect 486154 241325 492918 241561
rect 493154 241325 499918 241561
rect 500154 241325 506918 241561
rect 507154 241325 513918 241561
rect 514154 241325 527918 241561
rect 528154 241325 534918 241561
rect 535154 241325 541918 241561
rect 542154 241325 548918 241561
rect 549154 241325 555918 241561
rect 556154 241325 562918 241561
rect 563154 241325 569918 241561
rect 570154 241325 576918 241561
rect 577154 241325 587570 241561
rect 587806 241325 587890 241561
rect 588126 241325 588210 241561
rect 588446 241325 588530 241561
rect 588766 241325 588874 241561
rect -4950 241283 588874 241325
rect -4950 240494 588874 240536
rect -4950 240258 -3090 240494
rect -2854 240258 -2770 240494
rect -2534 240258 -2450 240494
rect -2214 240258 -2130 240494
rect -1894 240258 1186 240494
rect 1422 240258 8186 240494
rect 8422 240258 15186 240494
rect 15422 240258 22186 240494
rect 22422 240258 29186 240494
rect 29422 240258 36186 240494
rect 36422 240258 43186 240494
rect 43422 240258 50186 240494
rect 50422 240258 57186 240494
rect 57422 240258 64186 240494
rect 64422 240258 71186 240494
rect 71422 240258 78186 240494
rect 78422 240258 85186 240494
rect 85422 240258 92186 240494
rect 92422 240258 99186 240494
rect 99422 240258 106186 240494
rect 106422 240258 113186 240494
rect 113422 240258 120186 240494
rect 120422 240258 127186 240494
rect 127422 240258 134186 240494
rect 134422 240258 141186 240494
rect 141422 240258 148186 240494
rect 148422 240258 155186 240494
rect 155422 240258 162186 240494
rect 162422 240258 169186 240494
rect 169422 240258 176186 240494
rect 176422 240258 183186 240494
rect 183422 240258 190186 240494
rect 190422 240258 197186 240494
rect 197422 240258 204186 240494
rect 204422 240258 211186 240494
rect 211422 240258 218186 240494
rect 218422 240258 225186 240494
rect 225422 240258 232186 240494
rect 232422 240258 239186 240494
rect 239422 240258 246186 240494
rect 246422 240258 253186 240494
rect 253422 240258 260186 240494
rect 260422 240258 267186 240494
rect 267422 240258 274186 240494
rect 274422 240258 281186 240494
rect 281422 240258 288186 240494
rect 288422 240258 295186 240494
rect 295422 240258 302186 240494
rect 302422 240258 309186 240494
rect 309422 240258 316186 240494
rect 316422 240258 323186 240494
rect 323422 240258 330186 240494
rect 330422 240258 337186 240494
rect 337422 240258 344186 240494
rect 344422 240258 351186 240494
rect 351422 240258 358186 240494
rect 358422 240258 365186 240494
rect 365422 240258 372186 240494
rect 372422 240258 379186 240494
rect 379422 240258 386186 240494
rect 386422 240258 393186 240494
rect 393422 240258 400186 240494
rect 400422 240258 407186 240494
rect 407422 240258 414186 240494
rect 414422 240258 421186 240494
rect 421422 240258 428186 240494
rect 428422 240258 435186 240494
rect 435422 240258 442186 240494
rect 442422 240258 449186 240494
rect 449422 240258 456186 240494
rect 456422 240258 463186 240494
rect 463422 240258 470186 240494
rect 470422 240258 477186 240494
rect 477422 240258 484186 240494
rect 484422 240258 491186 240494
rect 491422 240258 498186 240494
rect 498422 240258 505186 240494
rect 505422 240258 512186 240494
rect 512422 240258 519186 240494
rect 519422 240258 533186 240494
rect 533422 240258 540186 240494
rect 540422 240258 547186 240494
rect 547422 240258 554186 240494
rect 554422 240258 561186 240494
rect 561422 240258 568186 240494
rect 568422 240258 575186 240494
rect 575422 240258 582186 240494
rect 582422 240258 585818 240494
rect 586054 240258 586138 240494
rect 586374 240258 586458 240494
rect 586694 240258 586778 240494
rect 587014 240258 588874 240494
rect -4950 240216 588874 240258
rect -4950 234561 588874 234603
rect -4950 234325 -4842 234561
rect -4606 234325 -4522 234561
rect -4286 234325 -4202 234561
rect -3966 234325 -3882 234561
rect -3646 234325 2918 234561
rect 3154 234325 9918 234561
rect 10154 234325 16918 234561
rect 17154 234325 23918 234561
rect 24154 234325 30918 234561
rect 31154 234325 37918 234561
rect 38154 234325 44918 234561
rect 45154 234325 51918 234561
rect 52154 234325 58918 234561
rect 59154 234325 65918 234561
rect 66154 234325 72918 234561
rect 73154 234325 79918 234561
rect 80154 234325 86918 234561
rect 87154 234325 93918 234561
rect 94154 234325 100918 234561
rect 101154 234325 107918 234561
rect 108154 234325 114918 234561
rect 115154 234325 121918 234561
rect 122154 234325 128918 234561
rect 129154 234325 135918 234561
rect 136154 234325 142918 234561
rect 143154 234325 149918 234561
rect 150154 234325 156918 234561
rect 157154 234325 163918 234561
rect 164154 234325 170918 234561
rect 171154 234325 177918 234561
rect 178154 234325 184918 234561
rect 185154 234325 191918 234561
rect 192154 234325 198918 234561
rect 199154 234325 205918 234561
rect 206154 234325 212918 234561
rect 213154 234325 219918 234561
rect 220154 234325 226918 234561
rect 227154 234325 233918 234561
rect 234154 234325 240918 234561
rect 241154 234325 247918 234561
rect 248154 234325 254918 234561
rect 255154 234325 261918 234561
rect 262154 234325 268918 234561
rect 269154 234325 275918 234561
rect 276154 234325 282918 234561
rect 283154 234325 289918 234561
rect 290154 234325 296918 234561
rect 297154 234325 303918 234561
rect 304154 234325 310918 234561
rect 311154 234325 317918 234561
rect 318154 234325 324918 234561
rect 325154 234325 331918 234561
rect 332154 234325 338918 234561
rect 339154 234325 345918 234561
rect 346154 234325 352918 234561
rect 353154 234325 359918 234561
rect 360154 234325 366918 234561
rect 367154 234325 373918 234561
rect 374154 234325 380918 234561
rect 381154 234325 387918 234561
rect 388154 234325 394918 234561
rect 395154 234325 401918 234561
rect 402154 234325 408918 234561
rect 409154 234325 415918 234561
rect 416154 234325 422918 234561
rect 423154 234325 429918 234561
rect 430154 234325 436918 234561
rect 437154 234325 443918 234561
rect 444154 234325 450918 234561
rect 451154 234325 457918 234561
rect 458154 234325 464918 234561
rect 465154 234325 471918 234561
rect 472154 234325 478918 234561
rect 479154 234325 485918 234561
rect 486154 234325 492918 234561
rect 493154 234325 499918 234561
rect 500154 234325 506918 234561
rect 507154 234325 513918 234561
rect 514154 234325 520918 234561
rect 521154 234325 527918 234561
rect 528154 234325 534918 234561
rect 535154 234325 541918 234561
rect 542154 234325 548918 234561
rect 549154 234325 555918 234561
rect 556154 234325 562918 234561
rect 563154 234325 569918 234561
rect 570154 234325 576918 234561
rect 577154 234325 587570 234561
rect 587806 234325 587890 234561
rect 588126 234325 588210 234561
rect 588446 234325 588530 234561
rect 588766 234325 588874 234561
rect -4950 234283 588874 234325
rect -4950 233494 588874 233536
rect -4950 233258 -3090 233494
rect -2854 233258 -2770 233494
rect -2534 233258 -2450 233494
rect -2214 233258 -2130 233494
rect -1894 233258 1186 233494
rect 1422 233258 8186 233494
rect 8422 233258 15186 233494
rect 15422 233258 22186 233494
rect 22422 233258 29186 233494
rect 29422 233258 36186 233494
rect 36422 233258 43186 233494
rect 43422 233258 50186 233494
rect 50422 233258 57186 233494
rect 57422 233258 64186 233494
rect 64422 233258 71186 233494
rect 71422 233258 78186 233494
rect 78422 233258 85186 233494
rect 85422 233258 92186 233494
rect 92422 233258 99186 233494
rect 99422 233258 106186 233494
rect 106422 233258 113186 233494
rect 113422 233258 120186 233494
rect 120422 233258 127186 233494
rect 127422 233258 134186 233494
rect 134422 233258 141186 233494
rect 141422 233258 148186 233494
rect 148422 233258 155186 233494
rect 155422 233258 162186 233494
rect 162422 233258 169186 233494
rect 169422 233258 176186 233494
rect 176422 233258 183186 233494
rect 183422 233258 190186 233494
rect 190422 233258 197186 233494
rect 197422 233258 204186 233494
rect 204422 233258 211186 233494
rect 211422 233258 218186 233494
rect 218422 233258 225186 233494
rect 225422 233258 232186 233494
rect 232422 233258 239186 233494
rect 239422 233258 246186 233494
rect 246422 233258 253186 233494
rect 253422 233258 260186 233494
rect 260422 233258 267186 233494
rect 267422 233258 274186 233494
rect 274422 233258 281186 233494
rect 281422 233258 288186 233494
rect 288422 233258 295186 233494
rect 295422 233258 302186 233494
rect 302422 233258 309186 233494
rect 309422 233258 316186 233494
rect 316422 233258 323186 233494
rect 323422 233258 330186 233494
rect 330422 233258 337186 233494
rect 337422 233258 344186 233494
rect 344422 233258 351186 233494
rect 351422 233258 358186 233494
rect 358422 233258 365186 233494
rect 365422 233258 372186 233494
rect 372422 233258 379186 233494
rect 379422 233258 386186 233494
rect 386422 233258 393186 233494
rect 393422 233258 400186 233494
rect 400422 233258 407186 233494
rect 407422 233258 414186 233494
rect 414422 233258 421186 233494
rect 421422 233258 428186 233494
rect 428422 233258 435186 233494
rect 435422 233258 442186 233494
rect 442422 233258 449186 233494
rect 449422 233258 456186 233494
rect 456422 233258 463186 233494
rect 463422 233258 470186 233494
rect 470422 233258 477186 233494
rect 477422 233258 484186 233494
rect 484422 233258 491186 233494
rect 491422 233258 498186 233494
rect 498422 233258 505186 233494
rect 505422 233258 512186 233494
rect 512422 233258 519186 233494
rect 519422 233258 526186 233494
rect 526422 233258 533186 233494
rect 533422 233258 540186 233494
rect 540422 233258 547186 233494
rect 547422 233258 554186 233494
rect 554422 233258 561186 233494
rect 561422 233258 568186 233494
rect 568422 233258 575186 233494
rect 575422 233258 582186 233494
rect 582422 233258 585818 233494
rect 586054 233258 586138 233494
rect 586374 233258 586458 233494
rect 586694 233258 586778 233494
rect 587014 233258 588874 233494
rect -4950 233216 588874 233258
rect -4950 227561 588874 227603
rect -4950 227325 -4842 227561
rect -4606 227325 -4522 227561
rect -4286 227325 -4202 227561
rect -3966 227325 -3882 227561
rect -3646 227325 2918 227561
rect 3154 227325 9918 227561
rect 10154 227325 16918 227561
rect 17154 227325 23918 227561
rect 24154 227325 30918 227561
rect 31154 227325 37918 227561
rect 38154 227325 44918 227561
rect 45154 227325 51918 227561
rect 52154 227325 58918 227561
rect 59154 227325 65918 227561
rect 66154 227325 72918 227561
rect 73154 227325 79918 227561
rect 80154 227325 86918 227561
rect 87154 227325 93918 227561
rect 94154 227325 100918 227561
rect 101154 227325 107918 227561
rect 108154 227325 114918 227561
rect 115154 227325 121918 227561
rect 122154 227325 128918 227561
rect 129154 227325 135918 227561
rect 136154 227325 142918 227561
rect 143154 227325 149918 227561
rect 150154 227325 156918 227561
rect 157154 227325 163918 227561
rect 164154 227325 170918 227561
rect 171154 227325 177918 227561
rect 178154 227325 184918 227561
rect 185154 227325 191918 227561
rect 192154 227325 198918 227561
rect 199154 227325 205918 227561
rect 206154 227325 212918 227561
rect 213154 227325 219918 227561
rect 220154 227325 226918 227561
rect 227154 227325 233918 227561
rect 234154 227325 240918 227561
rect 241154 227325 247918 227561
rect 248154 227325 254918 227561
rect 255154 227325 261918 227561
rect 262154 227325 268918 227561
rect 269154 227325 275918 227561
rect 276154 227325 282918 227561
rect 283154 227325 289918 227561
rect 290154 227325 296918 227561
rect 297154 227325 303918 227561
rect 304154 227325 310918 227561
rect 311154 227325 317918 227561
rect 318154 227325 324918 227561
rect 325154 227325 331918 227561
rect 332154 227325 338918 227561
rect 339154 227325 345918 227561
rect 346154 227325 352918 227561
rect 353154 227325 359918 227561
rect 360154 227325 366918 227561
rect 367154 227325 373918 227561
rect 374154 227325 380918 227561
rect 381154 227325 387918 227561
rect 388154 227325 394918 227561
rect 395154 227325 401918 227561
rect 402154 227325 408918 227561
rect 409154 227325 415918 227561
rect 416154 227325 422918 227561
rect 423154 227325 429918 227561
rect 430154 227325 436918 227561
rect 437154 227325 443918 227561
rect 444154 227325 450918 227561
rect 451154 227325 457918 227561
rect 458154 227325 464918 227561
rect 465154 227325 471918 227561
rect 472154 227325 478918 227561
rect 479154 227325 485918 227561
rect 486154 227325 492918 227561
rect 493154 227325 499918 227561
rect 500154 227325 506918 227561
rect 507154 227325 513918 227561
rect 514154 227325 520918 227561
rect 521154 227325 527918 227561
rect 528154 227325 534918 227561
rect 535154 227325 541918 227561
rect 542154 227325 548918 227561
rect 549154 227325 555918 227561
rect 556154 227325 562918 227561
rect 563154 227325 569918 227561
rect 570154 227325 576918 227561
rect 577154 227325 587570 227561
rect 587806 227325 587890 227561
rect 588126 227325 588210 227561
rect 588446 227325 588530 227561
rect 588766 227325 588874 227561
rect -4950 227283 588874 227325
rect -4950 226494 588874 226536
rect -4950 226258 -3090 226494
rect -2854 226258 -2770 226494
rect -2534 226258 -2450 226494
rect -2214 226258 -2130 226494
rect -1894 226258 1186 226494
rect 1422 226258 8186 226494
rect 8422 226258 15186 226494
rect 15422 226258 22186 226494
rect 22422 226258 29186 226494
rect 29422 226258 36186 226494
rect 36422 226258 43186 226494
rect 43422 226258 50186 226494
rect 50422 226258 57186 226494
rect 57422 226258 64186 226494
rect 64422 226258 71186 226494
rect 71422 226258 78186 226494
rect 78422 226258 85186 226494
rect 85422 226258 92186 226494
rect 92422 226258 99186 226494
rect 99422 226258 106186 226494
rect 106422 226258 113186 226494
rect 113422 226258 120186 226494
rect 120422 226258 127186 226494
rect 127422 226258 134186 226494
rect 134422 226258 141186 226494
rect 141422 226258 148186 226494
rect 148422 226258 155186 226494
rect 155422 226258 162186 226494
rect 162422 226258 169186 226494
rect 169422 226258 176186 226494
rect 176422 226258 183186 226494
rect 183422 226258 190186 226494
rect 190422 226258 197186 226494
rect 197422 226258 204186 226494
rect 204422 226258 211186 226494
rect 211422 226258 218186 226494
rect 218422 226258 225186 226494
rect 225422 226258 232186 226494
rect 232422 226258 239186 226494
rect 239422 226258 246186 226494
rect 246422 226258 253186 226494
rect 253422 226258 260186 226494
rect 260422 226258 267186 226494
rect 267422 226258 274186 226494
rect 274422 226258 281186 226494
rect 281422 226258 288186 226494
rect 288422 226258 295186 226494
rect 295422 226258 302186 226494
rect 302422 226258 309186 226494
rect 309422 226258 316186 226494
rect 316422 226258 323186 226494
rect 323422 226258 330186 226494
rect 330422 226258 337186 226494
rect 337422 226258 344186 226494
rect 344422 226258 351186 226494
rect 351422 226258 358186 226494
rect 358422 226258 365186 226494
rect 365422 226258 372186 226494
rect 372422 226258 379186 226494
rect 379422 226258 386186 226494
rect 386422 226258 393186 226494
rect 393422 226258 400186 226494
rect 400422 226258 407186 226494
rect 407422 226258 414186 226494
rect 414422 226258 421186 226494
rect 421422 226258 428186 226494
rect 428422 226258 435186 226494
rect 435422 226258 442186 226494
rect 442422 226258 449186 226494
rect 449422 226258 456186 226494
rect 456422 226258 463186 226494
rect 463422 226258 470186 226494
rect 470422 226258 477186 226494
rect 477422 226258 484186 226494
rect 484422 226258 491186 226494
rect 491422 226258 498186 226494
rect 498422 226258 505186 226494
rect 505422 226258 512186 226494
rect 512422 226258 519186 226494
rect 519422 226258 526186 226494
rect 526422 226258 533186 226494
rect 533422 226258 540186 226494
rect 540422 226258 547186 226494
rect 547422 226258 554186 226494
rect 554422 226258 561186 226494
rect 561422 226258 568186 226494
rect 568422 226258 575186 226494
rect 575422 226258 582186 226494
rect 582422 226258 585818 226494
rect 586054 226258 586138 226494
rect 586374 226258 586458 226494
rect 586694 226258 586778 226494
rect 587014 226258 588874 226494
rect -4950 226216 588874 226258
rect -4950 220561 588874 220603
rect -4950 220325 -4842 220561
rect -4606 220325 -4522 220561
rect -4286 220325 -4202 220561
rect -3966 220325 -3882 220561
rect -3646 220325 2918 220561
rect 3154 220325 9918 220561
rect 10154 220325 16918 220561
rect 17154 220325 23918 220561
rect 24154 220325 30918 220561
rect 31154 220325 37918 220561
rect 38154 220325 44918 220561
rect 45154 220325 51918 220561
rect 52154 220325 58918 220561
rect 59154 220325 65918 220561
rect 66154 220325 72918 220561
rect 73154 220325 79918 220561
rect 80154 220325 86918 220561
rect 87154 220325 93918 220561
rect 94154 220325 100918 220561
rect 101154 220325 107918 220561
rect 108154 220325 114918 220561
rect 115154 220325 121918 220561
rect 122154 220325 128918 220561
rect 129154 220325 135918 220561
rect 136154 220325 142918 220561
rect 143154 220325 149918 220561
rect 150154 220325 156918 220561
rect 157154 220325 163918 220561
rect 164154 220325 170918 220561
rect 171154 220325 177918 220561
rect 178154 220325 184918 220561
rect 185154 220325 191918 220561
rect 192154 220325 198918 220561
rect 199154 220325 205918 220561
rect 206154 220325 212918 220561
rect 213154 220325 219918 220561
rect 220154 220325 226918 220561
rect 227154 220325 233918 220561
rect 234154 220325 240918 220561
rect 241154 220325 247918 220561
rect 248154 220325 254918 220561
rect 255154 220325 261918 220561
rect 262154 220325 268918 220561
rect 269154 220325 275918 220561
rect 276154 220325 282918 220561
rect 283154 220325 289918 220561
rect 290154 220325 296918 220561
rect 297154 220325 303918 220561
rect 304154 220325 310918 220561
rect 311154 220325 317918 220561
rect 318154 220325 324918 220561
rect 325154 220325 331918 220561
rect 332154 220325 338918 220561
rect 339154 220325 345918 220561
rect 346154 220325 352918 220561
rect 353154 220325 359918 220561
rect 360154 220325 366918 220561
rect 367154 220325 373918 220561
rect 374154 220325 380918 220561
rect 381154 220325 387918 220561
rect 388154 220325 394918 220561
rect 395154 220325 401918 220561
rect 402154 220325 408918 220561
rect 409154 220325 415918 220561
rect 416154 220325 422918 220561
rect 423154 220325 429918 220561
rect 430154 220325 436918 220561
rect 437154 220325 443918 220561
rect 444154 220325 450918 220561
rect 451154 220325 457918 220561
rect 458154 220325 464918 220561
rect 465154 220325 471918 220561
rect 472154 220325 478918 220561
rect 479154 220325 485918 220561
rect 486154 220325 492918 220561
rect 493154 220325 499918 220561
rect 500154 220325 506918 220561
rect 507154 220325 513918 220561
rect 514154 220325 520918 220561
rect 521154 220325 527918 220561
rect 528154 220325 534918 220561
rect 535154 220325 541918 220561
rect 542154 220325 548918 220561
rect 549154 220325 555918 220561
rect 556154 220325 562918 220561
rect 563154 220325 569918 220561
rect 570154 220325 576918 220561
rect 577154 220325 587570 220561
rect 587806 220325 587890 220561
rect 588126 220325 588210 220561
rect 588446 220325 588530 220561
rect 588766 220325 588874 220561
rect -4950 220283 588874 220325
rect -4950 219494 588874 219536
rect -4950 219258 -3090 219494
rect -2854 219258 -2770 219494
rect -2534 219258 -2450 219494
rect -2214 219258 -2130 219494
rect -1894 219258 1186 219494
rect 1422 219258 8186 219494
rect 8422 219258 15186 219494
rect 15422 219258 22186 219494
rect 22422 219258 29186 219494
rect 29422 219258 36186 219494
rect 36422 219258 43186 219494
rect 43422 219258 50186 219494
rect 50422 219258 57186 219494
rect 57422 219258 64186 219494
rect 64422 219258 71186 219494
rect 71422 219258 78186 219494
rect 78422 219258 85186 219494
rect 85422 219258 92186 219494
rect 92422 219258 99186 219494
rect 99422 219258 106186 219494
rect 106422 219258 113186 219494
rect 113422 219258 120186 219494
rect 120422 219258 127186 219494
rect 127422 219258 134186 219494
rect 134422 219258 141186 219494
rect 141422 219258 148186 219494
rect 148422 219258 155186 219494
rect 155422 219258 162186 219494
rect 162422 219258 169186 219494
rect 169422 219258 176186 219494
rect 176422 219258 183186 219494
rect 183422 219258 190186 219494
rect 190422 219258 197186 219494
rect 197422 219258 204186 219494
rect 204422 219258 211186 219494
rect 211422 219258 218186 219494
rect 218422 219258 225186 219494
rect 225422 219258 232186 219494
rect 232422 219258 239186 219494
rect 239422 219258 246186 219494
rect 246422 219258 253186 219494
rect 253422 219258 260186 219494
rect 260422 219258 267186 219494
rect 267422 219258 274186 219494
rect 274422 219258 281186 219494
rect 281422 219258 288186 219494
rect 288422 219258 295186 219494
rect 295422 219258 302186 219494
rect 302422 219258 309186 219494
rect 309422 219258 316186 219494
rect 316422 219258 323186 219494
rect 323422 219258 330186 219494
rect 330422 219258 337186 219494
rect 337422 219258 344186 219494
rect 344422 219258 351186 219494
rect 351422 219258 358186 219494
rect 358422 219258 365186 219494
rect 365422 219258 372186 219494
rect 372422 219258 379186 219494
rect 379422 219258 386186 219494
rect 386422 219258 393186 219494
rect 393422 219258 400186 219494
rect 400422 219258 407186 219494
rect 407422 219258 414186 219494
rect 414422 219258 421186 219494
rect 421422 219258 428186 219494
rect 428422 219258 435186 219494
rect 435422 219258 442186 219494
rect 442422 219258 449186 219494
rect 449422 219258 456186 219494
rect 456422 219258 463186 219494
rect 463422 219258 470186 219494
rect 470422 219258 477186 219494
rect 477422 219258 484186 219494
rect 484422 219258 491186 219494
rect 491422 219258 498186 219494
rect 498422 219258 505186 219494
rect 505422 219258 512186 219494
rect 512422 219258 519186 219494
rect 519422 219258 526186 219494
rect 526422 219258 533186 219494
rect 533422 219258 540186 219494
rect 540422 219258 547186 219494
rect 547422 219258 554186 219494
rect 554422 219258 561186 219494
rect 561422 219258 568186 219494
rect 568422 219258 575186 219494
rect 575422 219258 582186 219494
rect 582422 219258 585818 219494
rect 586054 219258 586138 219494
rect 586374 219258 586458 219494
rect 586694 219258 586778 219494
rect 587014 219258 588874 219494
rect -4950 219216 588874 219258
rect -4950 213561 588874 213603
rect -4950 213325 -4842 213561
rect -4606 213325 -4522 213561
rect -4286 213325 -4202 213561
rect -3966 213325 -3882 213561
rect -3646 213325 2918 213561
rect 3154 213325 9918 213561
rect 10154 213325 16918 213561
rect 17154 213325 23918 213561
rect 24154 213325 30918 213561
rect 31154 213325 37918 213561
rect 38154 213325 44918 213561
rect 45154 213325 51918 213561
rect 52154 213325 58918 213561
rect 59154 213325 65918 213561
rect 66154 213325 72918 213561
rect 73154 213325 79918 213561
rect 80154 213325 86918 213561
rect 87154 213325 93918 213561
rect 94154 213325 100918 213561
rect 101154 213325 107918 213561
rect 108154 213325 114918 213561
rect 115154 213325 121918 213561
rect 122154 213325 128918 213561
rect 129154 213325 135918 213561
rect 136154 213325 142918 213561
rect 143154 213325 149918 213561
rect 150154 213325 156918 213561
rect 157154 213325 163918 213561
rect 164154 213325 170918 213561
rect 171154 213325 177918 213561
rect 178154 213325 184918 213561
rect 185154 213325 191918 213561
rect 192154 213325 198918 213561
rect 199154 213325 205918 213561
rect 206154 213325 212918 213561
rect 213154 213325 219918 213561
rect 220154 213325 226918 213561
rect 227154 213325 233918 213561
rect 234154 213325 240918 213561
rect 241154 213325 247918 213561
rect 248154 213325 254918 213561
rect 255154 213325 261918 213561
rect 262154 213325 268918 213561
rect 269154 213325 275918 213561
rect 276154 213325 282918 213561
rect 283154 213325 289918 213561
rect 290154 213325 296918 213561
rect 297154 213325 303918 213561
rect 304154 213325 310918 213561
rect 311154 213325 317918 213561
rect 318154 213325 324918 213561
rect 325154 213325 331918 213561
rect 332154 213325 338918 213561
rect 339154 213325 345918 213561
rect 346154 213325 352918 213561
rect 353154 213325 359918 213561
rect 360154 213325 366918 213561
rect 367154 213325 373918 213561
rect 374154 213325 380918 213561
rect 381154 213325 387918 213561
rect 388154 213325 394918 213561
rect 395154 213325 401918 213561
rect 402154 213325 408918 213561
rect 409154 213325 415918 213561
rect 416154 213325 422918 213561
rect 423154 213325 429918 213561
rect 430154 213325 436918 213561
rect 437154 213325 443918 213561
rect 444154 213325 450918 213561
rect 451154 213325 457918 213561
rect 458154 213325 464918 213561
rect 465154 213325 471918 213561
rect 472154 213325 478918 213561
rect 479154 213325 485918 213561
rect 486154 213325 492918 213561
rect 493154 213325 499918 213561
rect 500154 213325 506918 213561
rect 507154 213325 513918 213561
rect 514154 213325 520918 213561
rect 521154 213325 527918 213561
rect 528154 213325 534918 213561
rect 535154 213325 541918 213561
rect 542154 213325 548918 213561
rect 549154 213325 555918 213561
rect 556154 213325 562918 213561
rect 563154 213325 569918 213561
rect 570154 213325 576918 213561
rect 577154 213325 587570 213561
rect 587806 213325 587890 213561
rect 588126 213325 588210 213561
rect 588446 213325 588530 213561
rect 588766 213325 588874 213561
rect -4950 213283 588874 213325
rect -4950 212494 588874 212536
rect -4950 212258 -3090 212494
rect -2854 212258 -2770 212494
rect -2534 212258 -2450 212494
rect -2214 212258 -2130 212494
rect -1894 212258 1186 212494
rect 1422 212258 8186 212494
rect 8422 212258 15186 212494
rect 15422 212258 22186 212494
rect 22422 212258 29186 212494
rect 29422 212258 36186 212494
rect 36422 212258 43186 212494
rect 43422 212258 50186 212494
rect 50422 212258 57186 212494
rect 57422 212258 64186 212494
rect 64422 212258 71186 212494
rect 71422 212258 78186 212494
rect 78422 212258 85186 212494
rect 85422 212258 92186 212494
rect 92422 212258 99186 212494
rect 99422 212258 106186 212494
rect 106422 212258 113186 212494
rect 113422 212258 120186 212494
rect 120422 212258 127186 212494
rect 127422 212258 134186 212494
rect 134422 212258 141186 212494
rect 141422 212258 148186 212494
rect 148422 212258 155186 212494
rect 155422 212258 162186 212494
rect 162422 212258 169186 212494
rect 169422 212258 176186 212494
rect 176422 212258 183186 212494
rect 183422 212258 190186 212494
rect 190422 212258 197186 212494
rect 197422 212258 204186 212494
rect 204422 212258 211186 212494
rect 211422 212258 218186 212494
rect 218422 212258 225186 212494
rect 225422 212258 232186 212494
rect 232422 212258 239186 212494
rect 239422 212258 246186 212494
rect 246422 212258 253186 212494
rect 253422 212258 260186 212494
rect 260422 212258 267186 212494
rect 267422 212258 274186 212494
rect 274422 212258 281186 212494
rect 281422 212258 288186 212494
rect 288422 212258 295186 212494
rect 295422 212258 302186 212494
rect 302422 212258 309186 212494
rect 309422 212258 316186 212494
rect 316422 212258 323186 212494
rect 323422 212258 330186 212494
rect 330422 212258 337186 212494
rect 337422 212258 344186 212494
rect 344422 212258 351186 212494
rect 351422 212258 358186 212494
rect 358422 212258 365186 212494
rect 365422 212258 372186 212494
rect 372422 212258 379186 212494
rect 379422 212258 386186 212494
rect 386422 212258 393186 212494
rect 393422 212258 400186 212494
rect 400422 212258 407186 212494
rect 407422 212258 414186 212494
rect 414422 212258 421186 212494
rect 421422 212258 428186 212494
rect 428422 212258 435186 212494
rect 435422 212258 442186 212494
rect 442422 212258 449186 212494
rect 449422 212258 456186 212494
rect 456422 212258 463186 212494
rect 463422 212258 470186 212494
rect 470422 212258 477186 212494
rect 477422 212258 484186 212494
rect 484422 212258 491186 212494
rect 491422 212258 498186 212494
rect 498422 212258 505186 212494
rect 505422 212258 512186 212494
rect 512422 212258 519186 212494
rect 519422 212258 526186 212494
rect 526422 212258 533186 212494
rect 533422 212258 540186 212494
rect 540422 212258 547186 212494
rect 547422 212258 554186 212494
rect 554422 212258 561186 212494
rect 561422 212258 568186 212494
rect 568422 212258 575186 212494
rect 575422 212258 582186 212494
rect 582422 212258 585818 212494
rect 586054 212258 586138 212494
rect 586374 212258 586458 212494
rect 586694 212258 586778 212494
rect 587014 212258 588874 212494
rect -4950 212216 588874 212258
rect -4950 206561 588874 206603
rect -4950 206325 -4842 206561
rect -4606 206325 -4522 206561
rect -4286 206325 -4202 206561
rect -3966 206325 -3882 206561
rect -3646 206325 2918 206561
rect 3154 206325 9918 206561
rect 10154 206325 16918 206561
rect 17154 206325 23918 206561
rect 24154 206325 30918 206561
rect 31154 206325 37918 206561
rect 38154 206325 44918 206561
rect 45154 206325 51918 206561
rect 52154 206325 58918 206561
rect 59154 206325 65918 206561
rect 66154 206325 72918 206561
rect 73154 206325 79918 206561
rect 80154 206325 86918 206561
rect 87154 206325 93918 206561
rect 94154 206325 100918 206561
rect 101154 206325 107918 206561
rect 108154 206325 114918 206561
rect 115154 206325 121918 206561
rect 122154 206325 128918 206561
rect 129154 206325 135918 206561
rect 136154 206325 142918 206561
rect 143154 206325 149918 206561
rect 150154 206325 156918 206561
rect 157154 206325 163918 206561
rect 164154 206325 170918 206561
rect 171154 206325 177918 206561
rect 178154 206325 184918 206561
rect 185154 206325 191918 206561
rect 192154 206325 198918 206561
rect 199154 206325 205918 206561
rect 206154 206325 212918 206561
rect 213154 206325 219918 206561
rect 220154 206325 226918 206561
rect 227154 206325 233918 206561
rect 234154 206325 240918 206561
rect 241154 206325 247918 206561
rect 248154 206325 254918 206561
rect 255154 206325 261918 206561
rect 262154 206325 268918 206561
rect 269154 206325 275918 206561
rect 276154 206325 282918 206561
rect 283154 206325 289918 206561
rect 290154 206325 296918 206561
rect 297154 206325 303918 206561
rect 304154 206325 310918 206561
rect 311154 206325 317918 206561
rect 318154 206325 324918 206561
rect 325154 206325 331918 206561
rect 332154 206325 338918 206561
rect 339154 206325 345918 206561
rect 346154 206325 352918 206561
rect 353154 206325 359918 206561
rect 360154 206325 366918 206561
rect 367154 206325 373918 206561
rect 374154 206325 380918 206561
rect 381154 206325 387918 206561
rect 388154 206325 394918 206561
rect 395154 206325 401918 206561
rect 402154 206325 408918 206561
rect 409154 206325 415918 206561
rect 416154 206325 422918 206561
rect 423154 206325 429918 206561
rect 430154 206325 436918 206561
rect 437154 206325 443918 206561
rect 444154 206325 450918 206561
rect 451154 206325 457918 206561
rect 458154 206325 464918 206561
rect 465154 206325 471918 206561
rect 472154 206325 478918 206561
rect 479154 206325 485918 206561
rect 486154 206325 492918 206561
rect 493154 206325 499918 206561
rect 500154 206325 506918 206561
rect 507154 206325 513918 206561
rect 514154 206325 520918 206561
rect 521154 206325 527918 206561
rect 528154 206325 534918 206561
rect 535154 206325 541918 206561
rect 542154 206325 548918 206561
rect 549154 206325 555918 206561
rect 556154 206325 562918 206561
rect 563154 206325 569918 206561
rect 570154 206325 576918 206561
rect 577154 206325 587570 206561
rect 587806 206325 587890 206561
rect 588126 206325 588210 206561
rect 588446 206325 588530 206561
rect 588766 206325 588874 206561
rect -4950 206283 588874 206325
rect -4950 205494 588874 205536
rect -4950 205258 -3090 205494
rect -2854 205258 -2770 205494
rect -2534 205258 -2450 205494
rect -2214 205258 -2130 205494
rect -1894 205258 1186 205494
rect 1422 205258 8186 205494
rect 8422 205258 15186 205494
rect 15422 205258 22186 205494
rect 22422 205258 29186 205494
rect 29422 205258 36186 205494
rect 36422 205258 43186 205494
rect 43422 205258 50186 205494
rect 50422 205258 57186 205494
rect 57422 205258 64186 205494
rect 64422 205258 71186 205494
rect 71422 205258 78186 205494
rect 78422 205258 85186 205494
rect 85422 205258 92186 205494
rect 92422 205258 99186 205494
rect 99422 205258 106186 205494
rect 106422 205258 113186 205494
rect 113422 205258 120186 205494
rect 120422 205258 127186 205494
rect 127422 205258 134186 205494
rect 134422 205258 141186 205494
rect 141422 205258 148186 205494
rect 148422 205258 155186 205494
rect 155422 205258 162186 205494
rect 162422 205258 169186 205494
rect 169422 205258 176186 205494
rect 176422 205258 183186 205494
rect 183422 205258 190186 205494
rect 190422 205258 197186 205494
rect 197422 205258 204186 205494
rect 204422 205258 211186 205494
rect 211422 205258 218186 205494
rect 218422 205258 225186 205494
rect 225422 205258 232186 205494
rect 232422 205258 239186 205494
rect 239422 205258 246186 205494
rect 246422 205258 253186 205494
rect 253422 205258 260186 205494
rect 260422 205258 267186 205494
rect 267422 205258 274186 205494
rect 274422 205258 281186 205494
rect 281422 205258 288186 205494
rect 288422 205258 295186 205494
rect 295422 205258 302186 205494
rect 302422 205258 309186 205494
rect 309422 205258 316186 205494
rect 316422 205258 323186 205494
rect 323422 205258 330186 205494
rect 330422 205258 337186 205494
rect 337422 205258 344186 205494
rect 344422 205258 351186 205494
rect 351422 205258 358186 205494
rect 358422 205258 365186 205494
rect 365422 205258 372186 205494
rect 372422 205258 379186 205494
rect 379422 205258 386186 205494
rect 386422 205258 393186 205494
rect 393422 205258 400186 205494
rect 400422 205258 407186 205494
rect 407422 205258 414186 205494
rect 414422 205258 421186 205494
rect 421422 205258 428186 205494
rect 428422 205258 435186 205494
rect 435422 205258 442186 205494
rect 442422 205258 449186 205494
rect 449422 205258 456186 205494
rect 456422 205258 463186 205494
rect 463422 205258 470186 205494
rect 470422 205258 477186 205494
rect 477422 205258 484186 205494
rect 484422 205258 491186 205494
rect 491422 205258 498186 205494
rect 498422 205258 505186 205494
rect 505422 205258 512186 205494
rect 512422 205258 519186 205494
rect 519422 205258 526186 205494
rect 526422 205258 533186 205494
rect 533422 205258 540186 205494
rect 540422 205258 547186 205494
rect 547422 205258 554186 205494
rect 554422 205258 561186 205494
rect 561422 205258 568186 205494
rect 568422 205258 575186 205494
rect 575422 205258 582186 205494
rect 582422 205258 585818 205494
rect 586054 205258 586138 205494
rect 586374 205258 586458 205494
rect 586694 205258 586778 205494
rect 587014 205258 588874 205494
rect -4950 205216 588874 205258
rect -4950 199561 588874 199603
rect -4950 199325 -4842 199561
rect -4606 199325 -4522 199561
rect -4286 199325 -4202 199561
rect -3966 199325 -3882 199561
rect -3646 199325 2918 199561
rect 3154 199325 9918 199561
rect 10154 199325 16918 199561
rect 17154 199325 23918 199561
rect 24154 199325 30918 199561
rect 31154 199325 37918 199561
rect 38154 199325 44918 199561
rect 45154 199325 51918 199561
rect 52154 199325 58918 199561
rect 59154 199325 65918 199561
rect 66154 199325 72918 199561
rect 73154 199325 79918 199561
rect 80154 199325 86918 199561
rect 87154 199325 93918 199561
rect 94154 199325 100918 199561
rect 101154 199325 107918 199561
rect 108154 199325 114918 199561
rect 115154 199325 121918 199561
rect 122154 199325 128918 199561
rect 129154 199325 135918 199561
rect 136154 199325 142918 199561
rect 143154 199325 149918 199561
rect 150154 199325 156918 199561
rect 157154 199325 163918 199561
rect 164154 199325 170918 199561
rect 171154 199325 177918 199561
rect 178154 199325 184918 199561
rect 185154 199325 191918 199561
rect 192154 199325 198918 199561
rect 199154 199325 205918 199561
rect 206154 199325 212918 199561
rect 213154 199325 219918 199561
rect 220154 199325 226918 199561
rect 227154 199325 233918 199561
rect 234154 199325 240918 199561
rect 241154 199325 247918 199561
rect 248154 199325 254918 199561
rect 255154 199325 261918 199561
rect 262154 199325 268918 199561
rect 269154 199325 275918 199561
rect 276154 199325 282918 199561
rect 283154 199325 289918 199561
rect 290154 199325 317918 199561
rect 318154 199325 324918 199561
rect 325154 199325 331918 199561
rect 332154 199325 338918 199561
rect 339154 199325 345918 199561
rect 346154 199325 352918 199561
rect 353154 199325 359918 199561
rect 360154 199325 366918 199561
rect 367154 199325 373918 199561
rect 374154 199325 380918 199561
rect 381154 199325 387918 199561
rect 388154 199325 394918 199561
rect 395154 199325 401918 199561
rect 402154 199325 408918 199561
rect 409154 199325 415918 199561
rect 416154 199325 422918 199561
rect 423154 199325 429918 199561
rect 430154 199325 436918 199561
rect 437154 199325 443918 199561
rect 444154 199325 450918 199561
rect 451154 199325 457918 199561
rect 458154 199325 464918 199561
rect 465154 199325 471918 199561
rect 472154 199325 478918 199561
rect 479154 199325 485918 199561
rect 486154 199325 492918 199561
rect 493154 199325 499918 199561
rect 500154 199325 506918 199561
rect 507154 199325 513918 199561
rect 514154 199325 520918 199561
rect 521154 199325 527918 199561
rect 528154 199325 534918 199561
rect 535154 199325 541918 199561
rect 542154 199325 548918 199561
rect 549154 199325 555918 199561
rect 556154 199325 562918 199561
rect 563154 199325 569918 199561
rect 570154 199325 576918 199561
rect 577154 199325 587570 199561
rect 587806 199325 587890 199561
rect 588126 199325 588210 199561
rect 588446 199325 588530 199561
rect 588766 199325 588874 199561
rect -4950 199283 588874 199325
rect -4950 198494 588874 198536
rect -4950 198258 -3090 198494
rect -2854 198258 -2770 198494
rect -2534 198258 -2450 198494
rect -2214 198258 -2130 198494
rect -1894 198258 1186 198494
rect 1422 198258 8186 198494
rect 8422 198258 15186 198494
rect 15422 198258 22186 198494
rect 22422 198258 29186 198494
rect 29422 198258 36186 198494
rect 36422 198258 43186 198494
rect 43422 198258 50186 198494
rect 50422 198258 57186 198494
rect 57422 198258 64186 198494
rect 64422 198258 71186 198494
rect 71422 198258 78186 198494
rect 78422 198258 85186 198494
rect 85422 198258 92186 198494
rect 92422 198258 99186 198494
rect 99422 198258 106186 198494
rect 106422 198258 113186 198494
rect 113422 198258 120186 198494
rect 120422 198258 127186 198494
rect 127422 198258 134186 198494
rect 134422 198258 141186 198494
rect 141422 198258 148186 198494
rect 148422 198258 155186 198494
rect 155422 198258 162186 198494
rect 162422 198258 169186 198494
rect 169422 198258 176186 198494
rect 176422 198258 183186 198494
rect 183422 198258 190186 198494
rect 190422 198258 197186 198494
rect 197422 198258 204186 198494
rect 204422 198258 211186 198494
rect 211422 198258 218186 198494
rect 218422 198258 225186 198494
rect 225422 198258 232186 198494
rect 232422 198258 239186 198494
rect 239422 198258 246186 198494
rect 246422 198258 253186 198494
rect 253422 198258 260186 198494
rect 260422 198258 267186 198494
rect 267422 198258 274186 198494
rect 274422 198258 281186 198494
rect 281422 198258 288186 198494
rect 288422 198258 316186 198494
rect 316422 198258 323186 198494
rect 323422 198258 330186 198494
rect 330422 198258 337186 198494
rect 337422 198258 344186 198494
rect 344422 198258 351186 198494
rect 351422 198258 358186 198494
rect 358422 198258 365186 198494
rect 365422 198258 372186 198494
rect 372422 198258 379186 198494
rect 379422 198258 386186 198494
rect 386422 198258 393186 198494
rect 393422 198258 400186 198494
rect 400422 198258 407186 198494
rect 407422 198258 414186 198494
rect 414422 198258 421186 198494
rect 421422 198258 428186 198494
rect 428422 198258 435186 198494
rect 435422 198258 442186 198494
rect 442422 198258 449186 198494
rect 449422 198258 456186 198494
rect 456422 198258 463186 198494
rect 463422 198258 470186 198494
rect 470422 198258 477186 198494
rect 477422 198258 484186 198494
rect 484422 198258 491186 198494
rect 491422 198258 498186 198494
rect 498422 198258 505186 198494
rect 505422 198258 512186 198494
rect 512422 198258 519186 198494
rect 519422 198258 526186 198494
rect 526422 198258 533186 198494
rect 533422 198258 540186 198494
rect 540422 198258 547186 198494
rect 547422 198258 554186 198494
rect 554422 198258 561186 198494
rect 561422 198258 568186 198494
rect 568422 198258 575186 198494
rect 575422 198258 582186 198494
rect 582422 198258 585818 198494
rect 586054 198258 586138 198494
rect 586374 198258 586458 198494
rect 586694 198258 586778 198494
rect 587014 198258 588874 198494
rect -4950 198216 588874 198258
rect -4950 192561 588874 192603
rect -4950 192325 -4842 192561
rect -4606 192325 -4522 192561
rect -4286 192325 -4202 192561
rect -3966 192325 -3882 192561
rect -3646 192325 2918 192561
rect 3154 192325 9918 192561
rect 10154 192325 16918 192561
rect 17154 192325 23918 192561
rect 24154 192325 30918 192561
rect 31154 192325 37918 192561
rect 38154 192325 44918 192561
rect 45154 192325 51918 192561
rect 52154 192325 58918 192561
rect 59154 192325 65918 192561
rect 66154 192325 72918 192561
rect 73154 192325 79918 192561
rect 80154 192325 86918 192561
rect 87154 192325 93918 192561
rect 94154 192325 100918 192561
rect 101154 192325 107918 192561
rect 108154 192325 114918 192561
rect 115154 192325 121918 192561
rect 122154 192325 128918 192561
rect 129154 192325 135918 192561
rect 136154 192325 142918 192561
rect 143154 192325 149918 192561
rect 150154 192325 156918 192561
rect 157154 192325 163918 192561
rect 164154 192325 170918 192561
rect 171154 192325 177918 192561
rect 178154 192325 184918 192561
rect 185154 192325 191918 192561
rect 192154 192325 198918 192561
rect 199154 192325 205918 192561
rect 206154 192325 212918 192561
rect 213154 192325 219918 192561
rect 220154 192325 226918 192561
rect 227154 192325 233918 192561
rect 234154 192325 240918 192561
rect 241154 192325 247918 192561
rect 248154 192325 254918 192561
rect 255154 192325 261918 192561
rect 262154 192325 268918 192561
rect 269154 192325 275918 192561
rect 276154 192325 282918 192561
rect 283154 192325 289918 192561
rect 290154 192325 296918 192561
rect 297154 192325 303918 192561
rect 304154 192325 310918 192561
rect 311154 192325 317918 192561
rect 318154 192325 324918 192561
rect 325154 192325 331918 192561
rect 332154 192325 338918 192561
rect 339154 192325 345918 192561
rect 346154 192325 352918 192561
rect 353154 192325 359918 192561
rect 360154 192325 366918 192561
rect 367154 192325 373918 192561
rect 374154 192325 380918 192561
rect 381154 192325 387918 192561
rect 388154 192325 394918 192561
rect 395154 192325 401918 192561
rect 402154 192325 408918 192561
rect 409154 192325 415918 192561
rect 416154 192325 422918 192561
rect 423154 192325 429918 192561
rect 430154 192325 436918 192561
rect 437154 192325 443918 192561
rect 444154 192325 450918 192561
rect 451154 192325 457918 192561
rect 458154 192325 464918 192561
rect 465154 192325 471918 192561
rect 472154 192325 478918 192561
rect 479154 192325 485918 192561
rect 486154 192325 492918 192561
rect 493154 192325 499918 192561
rect 500154 192325 506918 192561
rect 507154 192325 513918 192561
rect 514154 192325 520918 192561
rect 521154 192325 527918 192561
rect 528154 192325 534918 192561
rect 535154 192325 541918 192561
rect 542154 192325 548918 192561
rect 549154 192325 555918 192561
rect 556154 192325 562918 192561
rect 563154 192325 569918 192561
rect 570154 192325 576918 192561
rect 577154 192325 587570 192561
rect 587806 192325 587890 192561
rect 588126 192325 588210 192561
rect 588446 192325 588530 192561
rect 588766 192325 588874 192561
rect -4950 192283 588874 192325
rect -4950 191494 588874 191536
rect -4950 191258 -3090 191494
rect -2854 191258 -2770 191494
rect -2534 191258 -2450 191494
rect -2214 191258 -2130 191494
rect -1894 191258 1186 191494
rect 1422 191258 8186 191494
rect 8422 191258 15186 191494
rect 15422 191258 22186 191494
rect 22422 191258 29186 191494
rect 29422 191258 36186 191494
rect 36422 191258 43186 191494
rect 43422 191258 50186 191494
rect 50422 191258 57186 191494
rect 57422 191258 64186 191494
rect 64422 191258 71186 191494
rect 71422 191258 78186 191494
rect 78422 191258 85186 191494
rect 85422 191258 92186 191494
rect 92422 191258 99186 191494
rect 99422 191258 106186 191494
rect 106422 191258 113186 191494
rect 113422 191258 120186 191494
rect 120422 191258 127186 191494
rect 127422 191258 134186 191494
rect 134422 191258 141186 191494
rect 141422 191258 148186 191494
rect 148422 191258 155186 191494
rect 155422 191258 162186 191494
rect 162422 191258 169186 191494
rect 169422 191258 176186 191494
rect 176422 191258 183186 191494
rect 183422 191258 190186 191494
rect 190422 191258 197186 191494
rect 197422 191258 204186 191494
rect 204422 191258 211186 191494
rect 211422 191258 218186 191494
rect 218422 191258 225186 191494
rect 225422 191258 232186 191494
rect 232422 191258 239186 191494
rect 239422 191258 246186 191494
rect 246422 191258 253186 191494
rect 253422 191258 260186 191494
rect 260422 191258 267186 191494
rect 267422 191258 274186 191494
rect 274422 191258 281186 191494
rect 281422 191258 288186 191494
rect 288422 191258 295186 191494
rect 295422 191258 302186 191494
rect 302422 191258 309186 191494
rect 309422 191258 316186 191494
rect 316422 191258 323186 191494
rect 323422 191258 330186 191494
rect 330422 191258 337186 191494
rect 337422 191258 344186 191494
rect 344422 191258 351186 191494
rect 351422 191258 358186 191494
rect 358422 191258 365186 191494
rect 365422 191258 372186 191494
rect 372422 191258 379186 191494
rect 379422 191258 386186 191494
rect 386422 191258 393186 191494
rect 393422 191258 400186 191494
rect 400422 191258 407186 191494
rect 407422 191258 414186 191494
rect 414422 191258 421186 191494
rect 421422 191258 428186 191494
rect 428422 191258 435186 191494
rect 435422 191258 442186 191494
rect 442422 191258 449186 191494
rect 449422 191258 456186 191494
rect 456422 191258 463186 191494
rect 463422 191258 470186 191494
rect 470422 191258 477186 191494
rect 477422 191258 484186 191494
rect 484422 191258 491186 191494
rect 491422 191258 498186 191494
rect 498422 191258 505186 191494
rect 505422 191258 512186 191494
rect 512422 191258 519186 191494
rect 519422 191258 526186 191494
rect 526422 191258 533186 191494
rect 533422 191258 540186 191494
rect 540422 191258 547186 191494
rect 547422 191258 554186 191494
rect 554422 191258 561186 191494
rect 561422 191258 568186 191494
rect 568422 191258 575186 191494
rect 575422 191258 582186 191494
rect 582422 191258 585818 191494
rect 586054 191258 586138 191494
rect 586374 191258 586458 191494
rect 586694 191258 586778 191494
rect 587014 191258 588874 191494
rect -4950 191216 588874 191258
rect -4950 185561 588874 185603
rect -4950 185325 -4842 185561
rect -4606 185325 -4522 185561
rect -4286 185325 -4202 185561
rect -3966 185325 -3882 185561
rect -3646 185325 2918 185561
rect 3154 185325 9918 185561
rect 10154 185325 16918 185561
rect 17154 185325 23918 185561
rect 24154 185325 30918 185561
rect 31154 185325 37918 185561
rect 38154 185325 44918 185561
rect 45154 185325 51918 185561
rect 52154 185325 58918 185561
rect 59154 185325 65918 185561
rect 66154 185325 72918 185561
rect 73154 185325 79918 185561
rect 80154 185325 86918 185561
rect 87154 185325 93918 185561
rect 94154 185325 100918 185561
rect 101154 185325 107918 185561
rect 108154 185325 114918 185561
rect 115154 185325 121918 185561
rect 122154 185325 128918 185561
rect 129154 185325 135918 185561
rect 136154 185325 142918 185561
rect 143154 185325 149918 185561
rect 150154 185325 156918 185561
rect 157154 185325 163918 185561
rect 164154 185325 170918 185561
rect 171154 185325 177918 185561
rect 178154 185325 184918 185561
rect 185154 185325 191918 185561
rect 192154 185325 198918 185561
rect 199154 185325 205918 185561
rect 206154 185325 212918 185561
rect 213154 185325 219918 185561
rect 220154 185325 226918 185561
rect 227154 185325 233918 185561
rect 234154 185325 240918 185561
rect 241154 185325 247918 185561
rect 248154 185325 254918 185561
rect 255154 185325 261918 185561
rect 262154 185325 268918 185561
rect 269154 185325 275918 185561
rect 276154 185325 282918 185561
rect 283154 185325 289918 185561
rect 290154 185325 296918 185561
rect 297154 185325 303918 185561
rect 304154 185325 310918 185561
rect 311154 185325 317918 185561
rect 318154 185325 324918 185561
rect 325154 185325 331918 185561
rect 332154 185325 338918 185561
rect 339154 185325 345918 185561
rect 346154 185325 352918 185561
rect 353154 185325 359918 185561
rect 360154 185325 366918 185561
rect 367154 185325 373918 185561
rect 374154 185325 380918 185561
rect 381154 185325 387918 185561
rect 388154 185325 394918 185561
rect 395154 185325 401918 185561
rect 402154 185325 408918 185561
rect 409154 185325 415918 185561
rect 416154 185325 422918 185561
rect 423154 185325 429918 185561
rect 430154 185325 436918 185561
rect 437154 185325 443918 185561
rect 444154 185325 450918 185561
rect 451154 185325 457918 185561
rect 458154 185325 464918 185561
rect 465154 185325 471918 185561
rect 472154 185325 478918 185561
rect 479154 185325 485918 185561
rect 486154 185325 492918 185561
rect 493154 185325 499918 185561
rect 500154 185325 506918 185561
rect 507154 185325 513918 185561
rect 514154 185325 520918 185561
rect 521154 185325 527918 185561
rect 528154 185325 534918 185561
rect 535154 185325 541918 185561
rect 542154 185325 548918 185561
rect 549154 185325 555918 185561
rect 556154 185325 562918 185561
rect 563154 185325 569918 185561
rect 570154 185325 576918 185561
rect 577154 185325 587570 185561
rect 587806 185325 587890 185561
rect 588126 185325 588210 185561
rect 588446 185325 588530 185561
rect 588766 185325 588874 185561
rect -4950 185283 588874 185325
rect -4950 184494 588874 184536
rect -4950 184258 -3090 184494
rect -2854 184258 -2770 184494
rect -2534 184258 -2450 184494
rect -2214 184258 -2130 184494
rect -1894 184258 1186 184494
rect 1422 184258 8186 184494
rect 8422 184258 15186 184494
rect 15422 184258 22186 184494
rect 22422 184258 29186 184494
rect 29422 184258 36186 184494
rect 36422 184258 43186 184494
rect 43422 184258 50186 184494
rect 50422 184258 57186 184494
rect 57422 184258 64186 184494
rect 64422 184258 71186 184494
rect 71422 184258 78186 184494
rect 78422 184258 85186 184494
rect 85422 184258 92186 184494
rect 92422 184258 99186 184494
rect 99422 184258 106186 184494
rect 106422 184258 113186 184494
rect 113422 184258 120186 184494
rect 120422 184258 127186 184494
rect 127422 184258 134186 184494
rect 134422 184258 141186 184494
rect 141422 184258 148186 184494
rect 148422 184258 155186 184494
rect 155422 184258 162186 184494
rect 162422 184258 169186 184494
rect 169422 184258 176186 184494
rect 176422 184258 183186 184494
rect 183422 184258 190186 184494
rect 190422 184258 197186 184494
rect 197422 184258 204186 184494
rect 204422 184258 211186 184494
rect 211422 184258 218186 184494
rect 218422 184258 225186 184494
rect 225422 184258 232186 184494
rect 232422 184258 239186 184494
rect 239422 184258 246186 184494
rect 246422 184258 253186 184494
rect 253422 184258 260186 184494
rect 260422 184258 267186 184494
rect 267422 184258 274186 184494
rect 274422 184258 281186 184494
rect 281422 184258 288186 184494
rect 288422 184258 295186 184494
rect 295422 184258 302186 184494
rect 302422 184258 309186 184494
rect 309422 184258 316186 184494
rect 316422 184258 323186 184494
rect 323422 184258 330186 184494
rect 330422 184258 337186 184494
rect 337422 184258 344186 184494
rect 344422 184258 351186 184494
rect 351422 184258 358186 184494
rect 358422 184258 365186 184494
rect 365422 184258 372186 184494
rect 372422 184258 379186 184494
rect 379422 184258 386186 184494
rect 386422 184258 393186 184494
rect 393422 184258 400186 184494
rect 400422 184258 407186 184494
rect 407422 184258 414186 184494
rect 414422 184258 421186 184494
rect 421422 184258 428186 184494
rect 428422 184258 435186 184494
rect 435422 184258 442186 184494
rect 442422 184258 449186 184494
rect 449422 184258 456186 184494
rect 456422 184258 463186 184494
rect 463422 184258 470186 184494
rect 470422 184258 477186 184494
rect 477422 184258 484186 184494
rect 484422 184258 491186 184494
rect 491422 184258 498186 184494
rect 498422 184258 505186 184494
rect 505422 184258 512186 184494
rect 512422 184258 519186 184494
rect 519422 184258 526186 184494
rect 526422 184258 533186 184494
rect 533422 184258 540186 184494
rect 540422 184258 547186 184494
rect 547422 184258 554186 184494
rect 554422 184258 561186 184494
rect 561422 184258 568186 184494
rect 568422 184258 575186 184494
rect 575422 184258 582186 184494
rect 582422 184258 585818 184494
rect 586054 184258 586138 184494
rect 586374 184258 586458 184494
rect 586694 184258 586778 184494
rect 587014 184258 588874 184494
rect -4950 184216 588874 184258
rect -4950 178561 588874 178603
rect -4950 178325 -4842 178561
rect -4606 178325 -4522 178561
rect -4286 178325 -4202 178561
rect -3966 178325 -3882 178561
rect -3646 178325 2918 178561
rect 3154 178325 9918 178561
rect 10154 178325 16918 178561
rect 17154 178325 23918 178561
rect 24154 178325 30918 178561
rect 31154 178325 37918 178561
rect 38154 178325 44918 178561
rect 45154 178325 51918 178561
rect 52154 178325 58918 178561
rect 59154 178325 65918 178561
rect 66154 178325 72918 178561
rect 73154 178325 79918 178561
rect 80154 178325 86918 178561
rect 87154 178325 93918 178561
rect 94154 178325 100918 178561
rect 101154 178325 107918 178561
rect 108154 178325 114918 178561
rect 115154 178325 121918 178561
rect 122154 178325 128918 178561
rect 129154 178325 135918 178561
rect 136154 178325 142918 178561
rect 143154 178325 149918 178561
rect 150154 178325 156918 178561
rect 157154 178325 163918 178561
rect 164154 178325 170918 178561
rect 171154 178325 177918 178561
rect 178154 178325 184918 178561
rect 185154 178325 191918 178561
rect 192154 178325 198918 178561
rect 199154 178325 205918 178561
rect 206154 178325 212918 178561
rect 213154 178325 219918 178561
rect 220154 178325 226918 178561
rect 227154 178325 233918 178561
rect 234154 178325 240918 178561
rect 241154 178325 247918 178561
rect 248154 178325 254918 178561
rect 255154 178325 261918 178561
rect 262154 178325 268918 178561
rect 269154 178325 275918 178561
rect 276154 178325 282918 178561
rect 283154 178325 289918 178561
rect 290154 178325 296918 178561
rect 297154 178325 303918 178561
rect 304154 178325 310918 178561
rect 311154 178325 317918 178561
rect 318154 178325 324918 178561
rect 325154 178325 331918 178561
rect 332154 178325 338918 178561
rect 339154 178325 345918 178561
rect 346154 178325 352918 178561
rect 353154 178325 359918 178561
rect 360154 178325 366918 178561
rect 367154 178325 373918 178561
rect 374154 178325 380918 178561
rect 381154 178325 387918 178561
rect 388154 178325 394918 178561
rect 395154 178325 401918 178561
rect 402154 178325 408918 178561
rect 409154 178325 415918 178561
rect 416154 178325 422918 178561
rect 423154 178325 429918 178561
rect 430154 178325 436918 178561
rect 437154 178325 443918 178561
rect 444154 178325 450918 178561
rect 451154 178325 457918 178561
rect 458154 178325 464918 178561
rect 465154 178325 471918 178561
rect 472154 178325 478918 178561
rect 479154 178325 485918 178561
rect 486154 178325 492918 178561
rect 493154 178325 499918 178561
rect 500154 178325 506918 178561
rect 507154 178325 513918 178561
rect 514154 178325 520918 178561
rect 521154 178325 527918 178561
rect 528154 178325 534918 178561
rect 535154 178325 541918 178561
rect 542154 178325 548918 178561
rect 549154 178325 555918 178561
rect 556154 178325 562918 178561
rect 563154 178325 569918 178561
rect 570154 178325 576918 178561
rect 577154 178325 587570 178561
rect 587806 178325 587890 178561
rect 588126 178325 588210 178561
rect 588446 178325 588530 178561
rect 588766 178325 588874 178561
rect -4950 178283 588874 178325
rect -4950 177494 588874 177536
rect -4950 177258 -3090 177494
rect -2854 177258 -2770 177494
rect -2534 177258 -2450 177494
rect -2214 177258 -2130 177494
rect -1894 177258 1186 177494
rect 1422 177258 8186 177494
rect 8422 177258 15186 177494
rect 15422 177258 22186 177494
rect 22422 177258 29186 177494
rect 29422 177258 36186 177494
rect 36422 177258 43186 177494
rect 43422 177258 50186 177494
rect 50422 177258 57186 177494
rect 57422 177258 64186 177494
rect 64422 177258 71186 177494
rect 71422 177258 78186 177494
rect 78422 177258 85186 177494
rect 85422 177258 92186 177494
rect 92422 177258 99186 177494
rect 99422 177258 106186 177494
rect 106422 177258 113186 177494
rect 113422 177258 120186 177494
rect 120422 177258 127186 177494
rect 127422 177258 134186 177494
rect 134422 177258 141186 177494
rect 141422 177258 148186 177494
rect 148422 177258 155186 177494
rect 155422 177258 162186 177494
rect 162422 177258 169186 177494
rect 169422 177258 176186 177494
rect 176422 177258 183186 177494
rect 183422 177258 190186 177494
rect 190422 177258 197186 177494
rect 197422 177258 204186 177494
rect 204422 177258 211186 177494
rect 211422 177258 218186 177494
rect 218422 177258 225186 177494
rect 225422 177258 232186 177494
rect 232422 177258 239186 177494
rect 239422 177258 246186 177494
rect 246422 177258 253186 177494
rect 253422 177258 260186 177494
rect 260422 177258 267186 177494
rect 267422 177258 274186 177494
rect 274422 177258 281186 177494
rect 281422 177258 288186 177494
rect 288422 177258 295186 177494
rect 295422 177258 302186 177494
rect 302422 177258 309186 177494
rect 309422 177258 316186 177494
rect 316422 177258 323186 177494
rect 323422 177258 330186 177494
rect 330422 177258 337186 177494
rect 337422 177258 344186 177494
rect 344422 177258 351186 177494
rect 351422 177258 358186 177494
rect 358422 177258 365186 177494
rect 365422 177258 372186 177494
rect 372422 177258 379186 177494
rect 379422 177258 386186 177494
rect 386422 177258 393186 177494
rect 393422 177258 400186 177494
rect 400422 177258 407186 177494
rect 407422 177258 414186 177494
rect 414422 177258 421186 177494
rect 421422 177258 428186 177494
rect 428422 177258 435186 177494
rect 435422 177258 442186 177494
rect 442422 177258 449186 177494
rect 449422 177258 456186 177494
rect 456422 177258 463186 177494
rect 463422 177258 470186 177494
rect 470422 177258 477186 177494
rect 477422 177258 484186 177494
rect 484422 177258 491186 177494
rect 491422 177258 498186 177494
rect 498422 177258 505186 177494
rect 505422 177258 512186 177494
rect 512422 177258 519186 177494
rect 519422 177258 526186 177494
rect 526422 177258 533186 177494
rect 533422 177258 540186 177494
rect 540422 177258 547186 177494
rect 547422 177258 554186 177494
rect 554422 177258 561186 177494
rect 561422 177258 568186 177494
rect 568422 177258 575186 177494
rect 575422 177258 582186 177494
rect 582422 177258 585818 177494
rect 586054 177258 586138 177494
rect 586374 177258 586458 177494
rect 586694 177258 586778 177494
rect 587014 177258 588874 177494
rect -4950 177216 588874 177258
rect -4950 171561 588874 171603
rect -4950 171325 -4842 171561
rect -4606 171325 -4522 171561
rect -4286 171325 -4202 171561
rect -3966 171325 -3882 171561
rect -3646 171325 2918 171561
rect 3154 171325 9918 171561
rect 10154 171325 16918 171561
rect 17154 171325 23918 171561
rect 24154 171325 30918 171561
rect 31154 171325 37918 171561
rect 38154 171325 44918 171561
rect 45154 171325 51918 171561
rect 52154 171325 58918 171561
rect 59154 171325 65918 171561
rect 66154 171325 72918 171561
rect 73154 171325 79918 171561
rect 80154 171325 86918 171561
rect 87154 171325 93918 171561
rect 94154 171325 100918 171561
rect 101154 171325 107918 171561
rect 108154 171325 114918 171561
rect 115154 171325 121918 171561
rect 122154 171325 128918 171561
rect 129154 171325 135918 171561
rect 136154 171325 142918 171561
rect 143154 171325 149918 171561
rect 150154 171325 156918 171561
rect 157154 171325 163918 171561
rect 164154 171325 170918 171561
rect 171154 171325 177918 171561
rect 178154 171325 184918 171561
rect 185154 171325 191918 171561
rect 192154 171325 198918 171561
rect 199154 171325 205918 171561
rect 206154 171325 212918 171561
rect 213154 171325 219918 171561
rect 220154 171325 226918 171561
rect 227154 171325 233918 171561
rect 234154 171325 240918 171561
rect 241154 171325 247918 171561
rect 248154 171325 254918 171561
rect 255154 171325 261918 171561
rect 262154 171325 268918 171561
rect 269154 171325 275918 171561
rect 276154 171325 282918 171561
rect 283154 171325 289918 171561
rect 290154 171325 296918 171561
rect 297154 171325 303918 171561
rect 304154 171325 310918 171561
rect 311154 171325 317918 171561
rect 318154 171325 324918 171561
rect 325154 171325 331918 171561
rect 332154 171325 338918 171561
rect 339154 171325 345918 171561
rect 346154 171325 352918 171561
rect 353154 171325 359918 171561
rect 360154 171325 366918 171561
rect 367154 171325 373918 171561
rect 374154 171325 380918 171561
rect 381154 171325 387918 171561
rect 388154 171325 394918 171561
rect 395154 171325 401918 171561
rect 402154 171325 408918 171561
rect 409154 171325 415918 171561
rect 416154 171325 422918 171561
rect 423154 171325 429918 171561
rect 430154 171325 436918 171561
rect 437154 171325 443918 171561
rect 444154 171325 450918 171561
rect 451154 171325 457918 171561
rect 458154 171325 464918 171561
rect 465154 171325 471918 171561
rect 472154 171325 478918 171561
rect 479154 171325 485918 171561
rect 486154 171325 492918 171561
rect 493154 171325 499918 171561
rect 500154 171325 506918 171561
rect 507154 171325 513918 171561
rect 514154 171325 520918 171561
rect 521154 171325 527918 171561
rect 528154 171325 534918 171561
rect 535154 171325 541918 171561
rect 542154 171325 548918 171561
rect 549154 171325 555918 171561
rect 556154 171325 562918 171561
rect 563154 171325 569918 171561
rect 570154 171325 576918 171561
rect 577154 171325 587570 171561
rect 587806 171325 587890 171561
rect 588126 171325 588210 171561
rect 588446 171325 588530 171561
rect 588766 171325 588874 171561
rect -4950 171283 588874 171325
rect -4950 170494 588874 170536
rect -4950 170258 -3090 170494
rect -2854 170258 -2770 170494
rect -2534 170258 -2450 170494
rect -2214 170258 -2130 170494
rect -1894 170258 1186 170494
rect 1422 170258 8186 170494
rect 8422 170258 15186 170494
rect 15422 170258 22186 170494
rect 22422 170258 29186 170494
rect 29422 170258 36186 170494
rect 36422 170258 43186 170494
rect 43422 170258 50186 170494
rect 50422 170258 57186 170494
rect 57422 170258 64186 170494
rect 64422 170258 71186 170494
rect 71422 170258 78186 170494
rect 78422 170258 85186 170494
rect 85422 170258 92186 170494
rect 92422 170258 99186 170494
rect 99422 170258 106186 170494
rect 106422 170258 113186 170494
rect 113422 170258 120186 170494
rect 120422 170258 127186 170494
rect 127422 170258 134186 170494
rect 134422 170258 141186 170494
rect 141422 170258 148186 170494
rect 148422 170258 155186 170494
rect 155422 170258 162186 170494
rect 162422 170258 169186 170494
rect 169422 170258 176186 170494
rect 176422 170258 183186 170494
rect 183422 170258 190186 170494
rect 190422 170258 197186 170494
rect 197422 170258 204186 170494
rect 204422 170258 211186 170494
rect 211422 170258 218186 170494
rect 218422 170258 225186 170494
rect 225422 170258 232186 170494
rect 232422 170258 239186 170494
rect 239422 170258 246186 170494
rect 246422 170258 253186 170494
rect 253422 170258 260186 170494
rect 260422 170258 267186 170494
rect 267422 170258 274186 170494
rect 274422 170258 281186 170494
rect 281422 170258 288186 170494
rect 288422 170258 295186 170494
rect 295422 170258 302186 170494
rect 302422 170258 309186 170494
rect 309422 170258 316186 170494
rect 316422 170258 323186 170494
rect 323422 170258 330186 170494
rect 330422 170258 337186 170494
rect 337422 170258 344186 170494
rect 344422 170258 351186 170494
rect 351422 170258 358186 170494
rect 358422 170258 365186 170494
rect 365422 170258 372186 170494
rect 372422 170258 379186 170494
rect 379422 170258 386186 170494
rect 386422 170258 393186 170494
rect 393422 170258 400186 170494
rect 400422 170258 407186 170494
rect 407422 170258 414186 170494
rect 414422 170258 421186 170494
rect 421422 170258 428186 170494
rect 428422 170258 435186 170494
rect 435422 170258 442186 170494
rect 442422 170258 449186 170494
rect 449422 170258 456186 170494
rect 456422 170258 463186 170494
rect 463422 170258 470186 170494
rect 470422 170258 477186 170494
rect 477422 170258 484186 170494
rect 484422 170258 491186 170494
rect 491422 170258 498186 170494
rect 498422 170258 505186 170494
rect 505422 170258 512186 170494
rect 512422 170258 519186 170494
rect 519422 170258 526186 170494
rect 526422 170258 533186 170494
rect 533422 170258 540186 170494
rect 540422 170258 547186 170494
rect 547422 170258 554186 170494
rect 554422 170258 561186 170494
rect 561422 170258 568186 170494
rect 568422 170258 575186 170494
rect 575422 170258 582186 170494
rect 582422 170258 585818 170494
rect 586054 170258 586138 170494
rect 586374 170258 586458 170494
rect 586694 170258 586778 170494
rect 587014 170258 588874 170494
rect -4950 170216 588874 170258
rect -4950 164561 588874 164603
rect -4950 164325 -4842 164561
rect -4606 164325 -4522 164561
rect -4286 164325 -4202 164561
rect -3966 164325 -3882 164561
rect -3646 164325 2918 164561
rect 3154 164325 9918 164561
rect 10154 164325 16918 164561
rect 17154 164325 23918 164561
rect 24154 164325 30918 164561
rect 31154 164325 37918 164561
rect 38154 164325 44918 164561
rect 45154 164325 51918 164561
rect 52154 164325 58918 164561
rect 59154 164325 65918 164561
rect 66154 164325 72918 164561
rect 73154 164325 79918 164561
rect 80154 164325 86918 164561
rect 87154 164325 93918 164561
rect 94154 164325 100918 164561
rect 101154 164325 107918 164561
rect 108154 164325 114918 164561
rect 115154 164325 121918 164561
rect 122154 164325 128918 164561
rect 129154 164325 135918 164561
rect 136154 164325 142918 164561
rect 143154 164325 149918 164561
rect 150154 164325 156918 164561
rect 157154 164325 163918 164561
rect 164154 164325 170918 164561
rect 171154 164325 177918 164561
rect 178154 164325 184918 164561
rect 185154 164325 191918 164561
rect 192154 164325 198918 164561
rect 199154 164325 205918 164561
rect 206154 164325 212918 164561
rect 213154 164325 219918 164561
rect 220154 164325 226918 164561
rect 227154 164325 233918 164561
rect 234154 164325 240918 164561
rect 241154 164325 247918 164561
rect 248154 164325 254918 164561
rect 255154 164325 261918 164561
rect 262154 164325 268918 164561
rect 269154 164325 275918 164561
rect 276154 164325 282918 164561
rect 283154 164325 289918 164561
rect 290154 164325 296918 164561
rect 297154 164325 303918 164561
rect 304154 164325 310918 164561
rect 311154 164325 317918 164561
rect 318154 164325 324918 164561
rect 325154 164325 331918 164561
rect 332154 164325 338918 164561
rect 339154 164325 345918 164561
rect 346154 164325 352918 164561
rect 353154 164325 359918 164561
rect 360154 164325 366918 164561
rect 367154 164325 373918 164561
rect 374154 164325 380918 164561
rect 381154 164325 387918 164561
rect 388154 164325 394918 164561
rect 395154 164325 401918 164561
rect 402154 164325 408918 164561
rect 409154 164325 415918 164561
rect 416154 164325 422918 164561
rect 423154 164325 429918 164561
rect 430154 164325 436918 164561
rect 437154 164325 443918 164561
rect 444154 164325 450918 164561
rect 451154 164325 457918 164561
rect 458154 164325 464918 164561
rect 465154 164325 471918 164561
rect 472154 164325 478918 164561
rect 479154 164325 485918 164561
rect 486154 164325 492918 164561
rect 493154 164325 499918 164561
rect 500154 164325 506918 164561
rect 507154 164325 513918 164561
rect 514154 164325 520918 164561
rect 521154 164325 527918 164561
rect 528154 164325 534918 164561
rect 535154 164325 541918 164561
rect 542154 164325 548918 164561
rect 549154 164325 555918 164561
rect 556154 164325 562918 164561
rect 563154 164325 569918 164561
rect 570154 164325 576918 164561
rect 577154 164325 587570 164561
rect 587806 164325 587890 164561
rect 588126 164325 588210 164561
rect 588446 164325 588530 164561
rect 588766 164325 588874 164561
rect -4950 164283 588874 164325
rect -4950 163494 588874 163536
rect -4950 163258 -3090 163494
rect -2854 163258 -2770 163494
rect -2534 163258 -2450 163494
rect -2214 163258 -2130 163494
rect -1894 163258 1186 163494
rect 1422 163258 8186 163494
rect 8422 163258 15186 163494
rect 15422 163258 22186 163494
rect 22422 163258 29186 163494
rect 29422 163258 36186 163494
rect 36422 163258 43186 163494
rect 43422 163258 50186 163494
rect 50422 163258 57186 163494
rect 57422 163258 64186 163494
rect 64422 163258 71186 163494
rect 71422 163258 78186 163494
rect 78422 163258 85186 163494
rect 85422 163258 92186 163494
rect 92422 163258 99186 163494
rect 99422 163258 106186 163494
rect 106422 163258 113186 163494
rect 113422 163258 120186 163494
rect 120422 163258 127186 163494
rect 127422 163258 134186 163494
rect 134422 163258 141186 163494
rect 141422 163258 148186 163494
rect 148422 163258 155186 163494
rect 155422 163258 162186 163494
rect 162422 163258 169186 163494
rect 169422 163258 176186 163494
rect 176422 163258 183186 163494
rect 183422 163258 190186 163494
rect 190422 163258 197186 163494
rect 197422 163258 204186 163494
rect 204422 163258 211186 163494
rect 211422 163258 218186 163494
rect 218422 163258 225186 163494
rect 225422 163258 232186 163494
rect 232422 163258 239186 163494
rect 239422 163258 246186 163494
rect 246422 163258 253186 163494
rect 253422 163258 260186 163494
rect 260422 163258 267186 163494
rect 267422 163258 274186 163494
rect 274422 163258 281186 163494
rect 281422 163258 288186 163494
rect 288422 163258 295186 163494
rect 295422 163258 302186 163494
rect 302422 163258 309186 163494
rect 309422 163258 316186 163494
rect 316422 163258 323186 163494
rect 323422 163258 330186 163494
rect 330422 163258 337186 163494
rect 337422 163258 344186 163494
rect 344422 163258 351186 163494
rect 351422 163258 358186 163494
rect 358422 163258 365186 163494
rect 365422 163258 372186 163494
rect 372422 163258 379186 163494
rect 379422 163258 386186 163494
rect 386422 163258 393186 163494
rect 393422 163258 400186 163494
rect 400422 163258 407186 163494
rect 407422 163258 414186 163494
rect 414422 163258 421186 163494
rect 421422 163258 428186 163494
rect 428422 163258 435186 163494
rect 435422 163258 442186 163494
rect 442422 163258 449186 163494
rect 449422 163258 456186 163494
rect 456422 163258 463186 163494
rect 463422 163258 470186 163494
rect 470422 163258 477186 163494
rect 477422 163258 484186 163494
rect 484422 163258 491186 163494
rect 491422 163258 498186 163494
rect 498422 163258 505186 163494
rect 505422 163258 512186 163494
rect 512422 163258 519186 163494
rect 519422 163258 526186 163494
rect 526422 163258 533186 163494
rect 533422 163258 540186 163494
rect 540422 163258 547186 163494
rect 547422 163258 554186 163494
rect 554422 163258 561186 163494
rect 561422 163258 568186 163494
rect 568422 163258 575186 163494
rect 575422 163258 582186 163494
rect 582422 163258 585818 163494
rect 586054 163258 586138 163494
rect 586374 163258 586458 163494
rect 586694 163258 586778 163494
rect 587014 163258 588874 163494
rect -4950 163216 588874 163258
rect -4950 157561 588874 157603
rect -4950 157325 -4842 157561
rect -4606 157325 -4522 157561
rect -4286 157325 -4202 157561
rect -3966 157325 -3882 157561
rect -3646 157325 2918 157561
rect 3154 157325 9918 157561
rect 10154 157325 16918 157561
rect 17154 157325 23918 157561
rect 24154 157325 30918 157561
rect 31154 157325 37918 157561
rect 38154 157325 44918 157561
rect 45154 157325 51918 157561
rect 52154 157325 58918 157561
rect 59154 157325 65918 157561
rect 66154 157325 72918 157561
rect 73154 157325 79918 157561
rect 80154 157325 86918 157561
rect 87154 157325 93918 157561
rect 94154 157325 100918 157561
rect 101154 157325 107918 157561
rect 108154 157325 114918 157561
rect 115154 157325 121918 157561
rect 122154 157325 128918 157561
rect 129154 157325 135918 157561
rect 136154 157325 142918 157561
rect 143154 157325 149918 157561
rect 150154 157325 156918 157561
rect 157154 157325 163918 157561
rect 164154 157325 170918 157561
rect 171154 157325 177918 157561
rect 178154 157325 184918 157561
rect 185154 157325 191918 157561
rect 192154 157325 198918 157561
rect 199154 157325 205918 157561
rect 206154 157325 212918 157561
rect 213154 157325 219918 157561
rect 220154 157325 226918 157561
rect 227154 157325 233918 157561
rect 234154 157325 240918 157561
rect 241154 157325 247918 157561
rect 248154 157325 254918 157561
rect 255154 157325 261918 157561
rect 262154 157325 268918 157561
rect 269154 157325 275918 157561
rect 276154 157325 282918 157561
rect 283154 157325 289918 157561
rect 290154 157325 296918 157561
rect 297154 157325 303918 157561
rect 304154 157325 310918 157561
rect 311154 157325 317918 157561
rect 318154 157325 324918 157561
rect 325154 157325 331918 157561
rect 332154 157325 338918 157561
rect 339154 157325 345918 157561
rect 346154 157325 352918 157561
rect 353154 157325 359918 157561
rect 360154 157325 366918 157561
rect 367154 157325 373918 157561
rect 374154 157325 380918 157561
rect 381154 157325 387918 157561
rect 388154 157325 394918 157561
rect 395154 157325 401918 157561
rect 402154 157325 408918 157561
rect 409154 157325 415918 157561
rect 416154 157325 422918 157561
rect 423154 157325 429918 157561
rect 430154 157325 436918 157561
rect 437154 157325 443918 157561
rect 444154 157325 450918 157561
rect 451154 157325 457918 157561
rect 458154 157325 464918 157561
rect 465154 157325 471918 157561
rect 472154 157325 478918 157561
rect 479154 157325 485918 157561
rect 486154 157325 492918 157561
rect 493154 157325 499918 157561
rect 500154 157325 506918 157561
rect 507154 157325 513918 157561
rect 514154 157325 520918 157561
rect 521154 157325 527918 157561
rect 528154 157325 534918 157561
rect 535154 157325 541918 157561
rect 542154 157325 548918 157561
rect 549154 157325 555918 157561
rect 556154 157325 562918 157561
rect 563154 157325 569918 157561
rect 570154 157325 576918 157561
rect 577154 157325 587570 157561
rect 587806 157325 587890 157561
rect 588126 157325 588210 157561
rect 588446 157325 588530 157561
rect 588766 157325 588874 157561
rect -4950 157283 588874 157325
rect -4950 156494 588874 156536
rect -4950 156258 -3090 156494
rect -2854 156258 -2770 156494
rect -2534 156258 -2450 156494
rect -2214 156258 -2130 156494
rect -1894 156258 1186 156494
rect 1422 156258 8186 156494
rect 8422 156258 15186 156494
rect 15422 156258 22186 156494
rect 22422 156258 29186 156494
rect 29422 156258 36186 156494
rect 36422 156258 43186 156494
rect 43422 156258 50186 156494
rect 50422 156258 57186 156494
rect 57422 156258 64186 156494
rect 64422 156258 71186 156494
rect 71422 156258 78186 156494
rect 78422 156258 85186 156494
rect 85422 156258 92186 156494
rect 92422 156258 99186 156494
rect 99422 156258 106186 156494
rect 106422 156258 113186 156494
rect 113422 156258 120186 156494
rect 120422 156258 127186 156494
rect 127422 156258 134186 156494
rect 134422 156258 141186 156494
rect 141422 156258 148186 156494
rect 148422 156258 155186 156494
rect 155422 156258 162186 156494
rect 162422 156258 169186 156494
rect 169422 156258 176186 156494
rect 176422 156258 183186 156494
rect 183422 156258 190186 156494
rect 190422 156258 197186 156494
rect 197422 156258 204186 156494
rect 204422 156258 211186 156494
rect 211422 156258 218186 156494
rect 218422 156258 225186 156494
rect 225422 156258 232186 156494
rect 232422 156258 239186 156494
rect 239422 156258 246186 156494
rect 246422 156258 253186 156494
rect 253422 156258 260186 156494
rect 260422 156258 267186 156494
rect 267422 156258 274186 156494
rect 274422 156258 281186 156494
rect 281422 156258 288186 156494
rect 288422 156258 295186 156494
rect 295422 156258 302186 156494
rect 302422 156258 309186 156494
rect 309422 156258 316186 156494
rect 316422 156258 323186 156494
rect 323422 156258 330186 156494
rect 330422 156258 337186 156494
rect 337422 156258 344186 156494
rect 344422 156258 351186 156494
rect 351422 156258 358186 156494
rect 358422 156258 365186 156494
rect 365422 156258 372186 156494
rect 372422 156258 379186 156494
rect 379422 156258 386186 156494
rect 386422 156258 393186 156494
rect 393422 156258 400186 156494
rect 400422 156258 407186 156494
rect 407422 156258 414186 156494
rect 414422 156258 421186 156494
rect 421422 156258 428186 156494
rect 428422 156258 435186 156494
rect 435422 156258 442186 156494
rect 442422 156258 449186 156494
rect 449422 156258 456186 156494
rect 456422 156258 463186 156494
rect 463422 156258 470186 156494
rect 470422 156258 477186 156494
rect 477422 156258 484186 156494
rect 484422 156258 491186 156494
rect 491422 156258 498186 156494
rect 498422 156258 505186 156494
rect 505422 156258 512186 156494
rect 512422 156258 519186 156494
rect 519422 156258 526186 156494
rect 526422 156258 533186 156494
rect 533422 156258 540186 156494
rect 540422 156258 547186 156494
rect 547422 156258 554186 156494
rect 554422 156258 561186 156494
rect 561422 156258 568186 156494
rect 568422 156258 575186 156494
rect 575422 156258 582186 156494
rect 582422 156258 585818 156494
rect 586054 156258 586138 156494
rect 586374 156258 586458 156494
rect 586694 156258 586778 156494
rect 587014 156258 588874 156494
rect -4950 156216 588874 156258
rect -4950 150561 588874 150603
rect -4950 150325 -4842 150561
rect -4606 150325 -4522 150561
rect -4286 150325 -4202 150561
rect -3966 150325 -3882 150561
rect -3646 150325 2918 150561
rect 3154 150325 9918 150561
rect 10154 150325 16918 150561
rect 17154 150325 23918 150561
rect 24154 150325 30918 150561
rect 31154 150325 37918 150561
rect 38154 150325 44918 150561
rect 45154 150325 51918 150561
rect 52154 150325 58918 150561
rect 59154 150325 65918 150561
rect 66154 150325 72918 150561
rect 73154 150325 79918 150561
rect 80154 150325 86918 150561
rect 87154 150325 93918 150561
rect 94154 150325 100918 150561
rect 101154 150325 107918 150561
rect 108154 150325 114918 150561
rect 115154 150325 121918 150561
rect 122154 150325 128918 150561
rect 129154 150325 135918 150561
rect 136154 150325 142918 150561
rect 143154 150325 149918 150561
rect 150154 150325 156918 150561
rect 157154 150325 163918 150561
rect 164154 150325 170918 150561
rect 171154 150325 177918 150561
rect 178154 150325 184918 150561
rect 185154 150325 191918 150561
rect 192154 150325 198918 150561
rect 199154 150325 205918 150561
rect 206154 150325 212918 150561
rect 213154 150325 219918 150561
rect 220154 150325 226918 150561
rect 227154 150325 233918 150561
rect 234154 150325 240918 150561
rect 241154 150325 247918 150561
rect 248154 150325 254918 150561
rect 255154 150325 261918 150561
rect 262154 150325 268918 150561
rect 269154 150325 275918 150561
rect 276154 150325 282918 150561
rect 283154 150325 289918 150561
rect 290154 150325 296918 150561
rect 297154 150325 303918 150561
rect 304154 150325 310918 150561
rect 311154 150325 317918 150561
rect 318154 150325 324918 150561
rect 325154 150325 331918 150561
rect 332154 150325 338918 150561
rect 339154 150325 345918 150561
rect 346154 150325 352918 150561
rect 353154 150325 359918 150561
rect 360154 150325 366918 150561
rect 367154 150325 373918 150561
rect 374154 150325 380918 150561
rect 381154 150325 387918 150561
rect 388154 150325 394918 150561
rect 395154 150325 401918 150561
rect 402154 150325 408918 150561
rect 409154 150325 415918 150561
rect 416154 150325 422918 150561
rect 423154 150325 429918 150561
rect 430154 150325 436918 150561
rect 437154 150325 443918 150561
rect 444154 150325 450918 150561
rect 451154 150325 457918 150561
rect 458154 150325 464918 150561
rect 465154 150325 471918 150561
rect 472154 150325 478918 150561
rect 479154 150325 485918 150561
rect 486154 150325 492918 150561
rect 493154 150325 499918 150561
rect 500154 150325 506918 150561
rect 507154 150325 513918 150561
rect 514154 150325 520918 150561
rect 521154 150325 527918 150561
rect 528154 150325 534918 150561
rect 535154 150325 541918 150561
rect 542154 150325 548918 150561
rect 549154 150325 555918 150561
rect 556154 150325 562918 150561
rect 563154 150325 569918 150561
rect 570154 150325 576918 150561
rect 577154 150325 587570 150561
rect 587806 150325 587890 150561
rect 588126 150325 588210 150561
rect 588446 150325 588530 150561
rect 588766 150325 588874 150561
rect -4950 150283 588874 150325
rect -4950 149494 588874 149536
rect -4950 149258 -3090 149494
rect -2854 149258 -2770 149494
rect -2534 149258 -2450 149494
rect -2214 149258 -2130 149494
rect -1894 149258 1186 149494
rect 1422 149258 8186 149494
rect 8422 149258 15186 149494
rect 15422 149258 22186 149494
rect 22422 149258 29186 149494
rect 29422 149258 36186 149494
rect 36422 149258 43186 149494
rect 43422 149258 50186 149494
rect 50422 149258 57186 149494
rect 57422 149258 64186 149494
rect 64422 149258 71186 149494
rect 71422 149258 78186 149494
rect 78422 149258 85186 149494
rect 85422 149258 92186 149494
rect 92422 149258 99186 149494
rect 99422 149258 106186 149494
rect 106422 149258 113186 149494
rect 113422 149258 120186 149494
rect 120422 149258 127186 149494
rect 127422 149258 134186 149494
rect 134422 149258 141186 149494
rect 141422 149258 148186 149494
rect 148422 149258 155186 149494
rect 155422 149258 162186 149494
rect 162422 149258 169186 149494
rect 169422 149258 176186 149494
rect 176422 149258 183186 149494
rect 183422 149258 190186 149494
rect 190422 149258 197186 149494
rect 197422 149258 204186 149494
rect 204422 149258 211186 149494
rect 211422 149258 218186 149494
rect 218422 149258 225186 149494
rect 225422 149258 232186 149494
rect 232422 149258 239186 149494
rect 239422 149258 246186 149494
rect 246422 149258 253186 149494
rect 253422 149258 260186 149494
rect 260422 149258 267186 149494
rect 267422 149258 274186 149494
rect 274422 149258 281186 149494
rect 281422 149258 288186 149494
rect 288422 149258 295186 149494
rect 295422 149258 302186 149494
rect 302422 149258 309186 149494
rect 309422 149258 316186 149494
rect 316422 149258 323186 149494
rect 323422 149258 330186 149494
rect 330422 149258 337186 149494
rect 337422 149258 344186 149494
rect 344422 149258 351186 149494
rect 351422 149258 358186 149494
rect 358422 149258 365186 149494
rect 365422 149258 372186 149494
rect 372422 149258 379186 149494
rect 379422 149258 386186 149494
rect 386422 149258 393186 149494
rect 393422 149258 400186 149494
rect 400422 149258 407186 149494
rect 407422 149258 414186 149494
rect 414422 149258 421186 149494
rect 421422 149258 428186 149494
rect 428422 149258 435186 149494
rect 435422 149258 442186 149494
rect 442422 149258 449186 149494
rect 449422 149258 456186 149494
rect 456422 149258 463186 149494
rect 463422 149258 470186 149494
rect 470422 149258 477186 149494
rect 477422 149258 484186 149494
rect 484422 149258 491186 149494
rect 491422 149258 498186 149494
rect 498422 149258 505186 149494
rect 505422 149258 512186 149494
rect 512422 149258 519186 149494
rect 519422 149258 526186 149494
rect 526422 149258 533186 149494
rect 533422 149258 540186 149494
rect 540422 149258 547186 149494
rect 547422 149258 554186 149494
rect 554422 149258 561186 149494
rect 561422 149258 568186 149494
rect 568422 149258 575186 149494
rect 575422 149258 582186 149494
rect 582422 149258 585818 149494
rect 586054 149258 586138 149494
rect 586374 149258 586458 149494
rect 586694 149258 586778 149494
rect 587014 149258 588874 149494
rect -4950 149216 588874 149258
rect -4950 143561 588874 143603
rect -4950 143325 -4842 143561
rect -4606 143325 -4522 143561
rect -4286 143325 -4202 143561
rect -3966 143325 -3882 143561
rect -3646 143325 2918 143561
rect 3154 143325 9918 143561
rect 10154 143325 16918 143561
rect 17154 143325 23918 143561
rect 24154 143325 30918 143561
rect 31154 143325 37918 143561
rect 38154 143325 44918 143561
rect 45154 143325 51918 143561
rect 52154 143325 58918 143561
rect 59154 143325 65918 143561
rect 66154 143325 72918 143561
rect 73154 143325 79918 143561
rect 80154 143325 86918 143561
rect 87154 143325 93918 143561
rect 94154 143325 100918 143561
rect 101154 143325 107918 143561
rect 108154 143325 114918 143561
rect 115154 143325 121918 143561
rect 122154 143325 128918 143561
rect 129154 143325 135918 143561
rect 136154 143325 142918 143561
rect 143154 143325 149918 143561
rect 150154 143325 156918 143561
rect 157154 143325 163918 143561
rect 164154 143325 170918 143561
rect 171154 143325 177918 143561
rect 178154 143325 184918 143561
rect 185154 143325 191918 143561
rect 192154 143325 198918 143561
rect 199154 143325 205918 143561
rect 206154 143325 212918 143561
rect 213154 143325 219918 143561
rect 220154 143325 226918 143561
rect 227154 143325 233918 143561
rect 234154 143325 240918 143561
rect 241154 143325 247918 143561
rect 248154 143325 254918 143561
rect 255154 143325 261918 143561
rect 262154 143325 268918 143561
rect 269154 143325 275918 143561
rect 276154 143325 282918 143561
rect 283154 143325 289918 143561
rect 290154 143325 296918 143561
rect 297154 143325 303918 143561
rect 304154 143325 310918 143561
rect 311154 143325 317918 143561
rect 318154 143325 324918 143561
rect 325154 143325 331918 143561
rect 332154 143325 338918 143561
rect 339154 143325 345918 143561
rect 346154 143325 352918 143561
rect 353154 143325 359918 143561
rect 360154 143325 366918 143561
rect 367154 143325 373918 143561
rect 374154 143325 380918 143561
rect 381154 143325 387918 143561
rect 388154 143325 394918 143561
rect 395154 143325 401918 143561
rect 402154 143325 408918 143561
rect 409154 143325 415918 143561
rect 416154 143325 422918 143561
rect 423154 143325 429918 143561
rect 430154 143325 436918 143561
rect 437154 143325 443918 143561
rect 444154 143325 450918 143561
rect 451154 143325 457918 143561
rect 458154 143325 464918 143561
rect 465154 143325 471918 143561
rect 472154 143325 478918 143561
rect 479154 143325 485918 143561
rect 486154 143325 492918 143561
rect 493154 143325 499918 143561
rect 500154 143325 506918 143561
rect 507154 143325 513918 143561
rect 514154 143325 520918 143561
rect 521154 143325 527918 143561
rect 528154 143325 534918 143561
rect 535154 143325 541918 143561
rect 542154 143325 548918 143561
rect 549154 143325 555918 143561
rect 556154 143325 562918 143561
rect 563154 143325 569918 143561
rect 570154 143325 576918 143561
rect 577154 143325 587570 143561
rect 587806 143325 587890 143561
rect 588126 143325 588210 143561
rect 588446 143325 588530 143561
rect 588766 143325 588874 143561
rect -4950 143283 588874 143325
rect -4950 142494 588874 142536
rect -4950 142258 -3090 142494
rect -2854 142258 -2770 142494
rect -2534 142258 -2450 142494
rect -2214 142258 -2130 142494
rect -1894 142258 1186 142494
rect 1422 142258 8186 142494
rect 8422 142258 15186 142494
rect 15422 142258 22186 142494
rect 22422 142258 29186 142494
rect 29422 142258 36186 142494
rect 36422 142258 43186 142494
rect 43422 142258 50186 142494
rect 50422 142258 57186 142494
rect 57422 142258 64186 142494
rect 64422 142258 71186 142494
rect 71422 142258 78186 142494
rect 78422 142258 85186 142494
rect 85422 142258 92186 142494
rect 92422 142258 99186 142494
rect 99422 142258 106186 142494
rect 106422 142258 113186 142494
rect 113422 142258 120186 142494
rect 120422 142258 127186 142494
rect 127422 142258 134186 142494
rect 134422 142258 141186 142494
rect 141422 142258 148186 142494
rect 148422 142258 155186 142494
rect 155422 142258 162186 142494
rect 162422 142258 169186 142494
rect 169422 142258 176186 142494
rect 176422 142258 183186 142494
rect 183422 142258 190186 142494
rect 190422 142258 197186 142494
rect 197422 142258 204186 142494
rect 204422 142258 211186 142494
rect 211422 142258 218186 142494
rect 218422 142258 225186 142494
rect 225422 142258 232186 142494
rect 232422 142258 239186 142494
rect 239422 142258 246186 142494
rect 246422 142258 253186 142494
rect 253422 142258 260186 142494
rect 260422 142258 267186 142494
rect 267422 142258 274186 142494
rect 274422 142258 281186 142494
rect 281422 142258 288186 142494
rect 288422 142258 295186 142494
rect 295422 142258 302186 142494
rect 302422 142258 309186 142494
rect 309422 142258 316186 142494
rect 316422 142258 323186 142494
rect 323422 142258 330186 142494
rect 330422 142258 337186 142494
rect 337422 142258 344186 142494
rect 344422 142258 351186 142494
rect 351422 142258 358186 142494
rect 358422 142258 365186 142494
rect 365422 142258 372186 142494
rect 372422 142258 379186 142494
rect 379422 142258 386186 142494
rect 386422 142258 393186 142494
rect 393422 142258 400186 142494
rect 400422 142258 407186 142494
rect 407422 142258 414186 142494
rect 414422 142258 421186 142494
rect 421422 142258 428186 142494
rect 428422 142258 435186 142494
rect 435422 142258 442186 142494
rect 442422 142258 449186 142494
rect 449422 142258 456186 142494
rect 456422 142258 463186 142494
rect 463422 142258 470186 142494
rect 470422 142258 477186 142494
rect 477422 142258 484186 142494
rect 484422 142258 491186 142494
rect 491422 142258 498186 142494
rect 498422 142258 505186 142494
rect 505422 142258 512186 142494
rect 512422 142258 519186 142494
rect 519422 142258 526186 142494
rect 526422 142258 533186 142494
rect 533422 142258 540186 142494
rect 540422 142258 547186 142494
rect 547422 142258 554186 142494
rect 554422 142258 561186 142494
rect 561422 142258 568186 142494
rect 568422 142258 575186 142494
rect 575422 142258 582186 142494
rect 582422 142258 585818 142494
rect 586054 142258 586138 142494
rect 586374 142258 586458 142494
rect 586694 142258 586778 142494
rect 587014 142258 588874 142494
rect -4950 142216 588874 142258
rect -4950 136561 588874 136603
rect -4950 136325 -4842 136561
rect -4606 136325 -4522 136561
rect -4286 136325 -4202 136561
rect -3966 136325 -3882 136561
rect -3646 136325 2918 136561
rect 3154 136325 9918 136561
rect 10154 136325 16918 136561
rect 17154 136325 23918 136561
rect 24154 136325 30918 136561
rect 31154 136325 37918 136561
rect 38154 136325 44918 136561
rect 45154 136325 51918 136561
rect 52154 136325 58918 136561
rect 59154 136325 65918 136561
rect 66154 136325 72918 136561
rect 73154 136325 79918 136561
rect 80154 136325 86918 136561
rect 87154 136325 93918 136561
rect 94154 136325 100918 136561
rect 101154 136325 107918 136561
rect 108154 136325 114918 136561
rect 115154 136325 121918 136561
rect 122154 136325 128918 136561
rect 129154 136325 135918 136561
rect 136154 136325 142918 136561
rect 143154 136325 149918 136561
rect 150154 136325 156918 136561
rect 157154 136325 163918 136561
rect 164154 136325 170918 136561
rect 171154 136325 177918 136561
rect 178154 136325 184918 136561
rect 185154 136325 191918 136561
rect 192154 136325 198918 136561
rect 199154 136325 205918 136561
rect 206154 136325 212918 136561
rect 213154 136325 219918 136561
rect 220154 136325 226918 136561
rect 227154 136325 233918 136561
rect 234154 136325 240918 136561
rect 241154 136325 247918 136561
rect 248154 136325 254918 136561
rect 255154 136325 261918 136561
rect 262154 136325 268918 136561
rect 269154 136325 275918 136561
rect 276154 136325 282918 136561
rect 283154 136325 289918 136561
rect 290154 136325 296918 136561
rect 297154 136325 303918 136561
rect 304154 136325 310918 136561
rect 311154 136325 317918 136561
rect 318154 136325 324918 136561
rect 325154 136325 331918 136561
rect 332154 136325 338918 136561
rect 339154 136325 345918 136561
rect 346154 136325 352918 136561
rect 353154 136325 359918 136561
rect 360154 136325 366918 136561
rect 367154 136325 373918 136561
rect 374154 136325 380918 136561
rect 381154 136325 387918 136561
rect 388154 136325 394918 136561
rect 395154 136325 401918 136561
rect 402154 136325 408918 136561
rect 409154 136325 415918 136561
rect 416154 136325 422918 136561
rect 423154 136325 429918 136561
rect 430154 136325 436918 136561
rect 437154 136325 443918 136561
rect 444154 136325 450918 136561
rect 451154 136325 457918 136561
rect 458154 136325 464918 136561
rect 465154 136325 471918 136561
rect 472154 136325 478918 136561
rect 479154 136325 485918 136561
rect 486154 136325 492918 136561
rect 493154 136325 499918 136561
rect 500154 136325 506918 136561
rect 507154 136325 513918 136561
rect 514154 136325 520918 136561
rect 521154 136325 527918 136561
rect 528154 136325 534918 136561
rect 535154 136325 541918 136561
rect 542154 136325 548918 136561
rect 549154 136325 555918 136561
rect 556154 136325 562918 136561
rect 563154 136325 569918 136561
rect 570154 136325 576918 136561
rect 577154 136325 587570 136561
rect 587806 136325 587890 136561
rect 588126 136325 588210 136561
rect 588446 136325 588530 136561
rect 588766 136325 588874 136561
rect -4950 136283 588874 136325
rect -4950 135494 588874 135536
rect -4950 135258 -3090 135494
rect -2854 135258 -2770 135494
rect -2534 135258 -2450 135494
rect -2214 135258 -2130 135494
rect -1894 135258 1186 135494
rect 1422 135258 8186 135494
rect 8422 135258 15186 135494
rect 15422 135258 22186 135494
rect 22422 135258 29186 135494
rect 29422 135258 36186 135494
rect 36422 135258 43186 135494
rect 43422 135258 50186 135494
rect 50422 135258 57186 135494
rect 57422 135258 64186 135494
rect 64422 135258 71186 135494
rect 71422 135258 78186 135494
rect 78422 135258 85186 135494
rect 85422 135258 92186 135494
rect 92422 135258 99186 135494
rect 99422 135258 106186 135494
rect 106422 135258 113186 135494
rect 113422 135258 120186 135494
rect 120422 135258 127186 135494
rect 127422 135258 134186 135494
rect 134422 135258 141186 135494
rect 141422 135258 148186 135494
rect 148422 135258 155186 135494
rect 155422 135258 162186 135494
rect 162422 135258 169186 135494
rect 169422 135258 176186 135494
rect 176422 135258 183186 135494
rect 183422 135258 190186 135494
rect 190422 135258 197186 135494
rect 197422 135258 204186 135494
rect 204422 135258 211186 135494
rect 211422 135258 218186 135494
rect 218422 135258 225186 135494
rect 225422 135258 232186 135494
rect 232422 135258 239186 135494
rect 239422 135258 246186 135494
rect 246422 135258 253186 135494
rect 253422 135258 260186 135494
rect 260422 135258 267186 135494
rect 267422 135258 274186 135494
rect 274422 135258 281186 135494
rect 281422 135258 288186 135494
rect 288422 135258 295186 135494
rect 295422 135258 302186 135494
rect 302422 135258 309186 135494
rect 309422 135258 316186 135494
rect 316422 135258 323186 135494
rect 323422 135258 330186 135494
rect 330422 135258 337186 135494
rect 337422 135258 344186 135494
rect 344422 135258 351186 135494
rect 351422 135258 358186 135494
rect 358422 135258 365186 135494
rect 365422 135258 372186 135494
rect 372422 135258 379186 135494
rect 379422 135258 386186 135494
rect 386422 135258 393186 135494
rect 393422 135258 400186 135494
rect 400422 135258 407186 135494
rect 407422 135258 414186 135494
rect 414422 135258 421186 135494
rect 421422 135258 428186 135494
rect 428422 135258 435186 135494
rect 435422 135258 442186 135494
rect 442422 135258 449186 135494
rect 449422 135258 456186 135494
rect 456422 135258 463186 135494
rect 463422 135258 470186 135494
rect 470422 135258 477186 135494
rect 477422 135258 484186 135494
rect 484422 135258 491186 135494
rect 491422 135258 498186 135494
rect 498422 135258 505186 135494
rect 505422 135258 512186 135494
rect 512422 135258 519186 135494
rect 519422 135258 526186 135494
rect 526422 135258 533186 135494
rect 533422 135258 540186 135494
rect 540422 135258 547186 135494
rect 547422 135258 554186 135494
rect 554422 135258 561186 135494
rect 561422 135258 568186 135494
rect 568422 135258 575186 135494
rect 575422 135258 582186 135494
rect 582422 135258 585818 135494
rect 586054 135258 586138 135494
rect 586374 135258 586458 135494
rect 586694 135258 586778 135494
rect 587014 135258 588874 135494
rect -4950 135216 588874 135258
rect -4950 129561 588874 129603
rect -4950 129325 -4842 129561
rect -4606 129325 -4522 129561
rect -4286 129325 -4202 129561
rect -3966 129325 -3882 129561
rect -3646 129325 2918 129561
rect 3154 129325 9918 129561
rect 10154 129325 16918 129561
rect 17154 129325 23918 129561
rect 24154 129325 30918 129561
rect 31154 129325 37918 129561
rect 38154 129325 44918 129561
rect 45154 129325 51918 129561
rect 52154 129325 58918 129561
rect 59154 129325 65918 129561
rect 66154 129325 72918 129561
rect 73154 129325 79918 129561
rect 80154 129325 86918 129561
rect 87154 129325 93918 129561
rect 94154 129325 100918 129561
rect 101154 129325 107918 129561
rect 108154 129325 114918 129561
rect 115154 129325 121918 129561
rect 122154 129325 128918 129561
rect 129154 129325 135918 129561
rect 136154 129325 142918 129561
rect 143154 129325 149918 129561
rect 150154 129325 156918 129561
rect 157154 129325 163918 129561
rect 164154 129325 170918 129561
rect 171154 129325 177918 129561
rect 178154 129325 184918 129561
rect 185154 129325 191918 129561
rect 192154 129325 198918 129561
rect 199154 129325 205918 129561
rect 206154 129325 212918 129561
rect 213154 129325 219918 129561
rect 220154 129325 226918 129561
rect 227154 129325 233918 129561
rect 234154 129325 240918 129561
rect 241154 129325 247918 129561
rect 248154 129325 254918 129561
rect 255154 129325 261918 129561
rect 262154 129325 268918 129561
rect 269154 129325 275918 129561
rect 276154 129325 282918 129561
rect 283154 129325 289918 129561
rect 290154 129325 296918 129561
rect 297154 129325 303918 129561
rect 304154 129325 310918 129561
rect 311154 129325 317918 129561
rect 318154 129325 324918 129561
rect 325154 129325 331918 129561
rect 332154 129325 338918 129561
rect 339154 129325 345918 129561
rect 346154 129325 352918 129561
rect 353154 129325 359918 129561
rect 360154 129325 366918 129561
rect 367154 129325 373918 129561
rect 374154 129325 380918 129561
rect 381154 129325 387918 129561
rect 388154 129325 394918 129561
rect 395154 129325 401918 129561
rect 402154 129325 408918 129561
rect 409154 129325 415918 129561
rect 416154 129325 422918 129561
rect 423154 129325 429918 129561
rect 430154 129325 436918 129561
rect 437154 129325 443918 129561
rect 444154 129325 450918 129561
rect 451154 129325 457918 129561
rect 458154 129325 464918 129561
rect 465154 129325 471918 129561
rect 472154 129325 478918 129561
rect 479154 129325 485918 129561
rect 486154 129325 492918 129561
rect 493154 129325 499918 129561
rect 500154 129325 506918 129561
rect 507154 129325 513918 129561
rect 514154 129325 520918 129561
rect 521154 129325 527918 129561
rect 528154 129325 534918 129561
rect 535154 129325 541918 129561
rect 542154 129325 548918 129561
rect 549154 129325 555918 129561
rect 556154 129325 562918 129561
rect 563154 129325 569918 129561
rect 570154 129325 576918 129561
rect 577154 129325 587570 129561
rect 587806 129325 587890 129561
rect 588126 129325 588210 129561
rect 588446 129325 588530 129561
rect 588766 129325 588874 129561
rect -4950 129283 588874 129325
rect -4950 128494 588874 128536
rect -4950 128258 -3090 128494
rect -2854 128258 -2770 128494
rect -2534 128258 -2450 128494
rect -2214 128258 -2130 128494
rect -1894 128258 1186 128494
rect 1422 128258 8186 128494
rect 8422 128258 15186 128494
rect 15422 128258 22186 128494
rect 22422 128258 29186 128494
rect 29422 128258 36186 128494
rect 36422 128258 43186 128494
rect 43422 128258 50186 128494
rect 50422 128258 57186 128494
rect 57422 128258 64186 128494
rect 64422 128258 71186 128494
rect 71422 128258 78186 128494
rect 78422 128258 85186 128494
rect 85422 128258 92186 128494
rect 92422 128258 99186 128494
rect 99422 128258 106186 128494
rect 106422 128258 113186 128494
rect 113422 128258 120186 128494
rect 120422 128258 127186 128494
rect 127422 128258 134186 128494
rect 134422 128258 141186 128494
rect 141422 128258 148186 128494
rect 148422 128258 155186 128494
rect 155422 128258 162186 128494
rect 162422 128258 169186 128494
rect 169422 128258 176186 128494
rect 176422 128258 183186 128494
rect 183422 128258 190186 128494
rect 190422 128258 197186 128494
rect 197422 128258 204186 128494
rect 204422 128258 211186 128494
rect 211422 128258 218186 128494
rect 218422 128258 225186 128494
rect 225422 128258 232186 128494
rect 232422 128258 239186 128494
rect 239422 128258 246186 128494
rect 246422 128258 253186 128494
rect 253422 128258 260186 128494
rect 260422 128258 267186 128494
rect 267422 128258 274186 128494
rect 274422 128258 281186 128494
rect 281422 128258 288186 128494
rect 288422 128258 295186 128494
rect 295422 128258 302186 128494
rect 302422 128258 309186 128494
rect 309422 128258 316186 128494
rect 316422 128258 323186 128494
rect 323422 128258 330186 128494
rect 330422 128258 337186 128494
rect 337422 128258 344186 128494
rect 344422 128258 351186 128494
rect 351422 128258 358186 128494
rect 358422 128258 365186 128494
rect 365422 128258 372186 128494
rect 372422 128258 379186 128494
rect 379422 128258 386186 128494
rect 386422 128258 393186 128494
rect 393422 128258 400186 128494
rect 400422 128258 407186 128494
rect 407422 128258 414186 128494
rect 414422 128258 421186 128494
rect 421422 128258 428186 128494
rect 428422 128258 435186 128494
rect 435422 128258 442186 128494
rect 442422 128258 449186 128494
rect 449422 128258 456186 128494
rect 456422 128258 463186 128494
rect 463422 128258 470186 128494
rect 470422 128258 477186 128494
rect 477422 128258 484186 128494
rect 484422 128258 491186 128494
rect 491422 128258 498186 128494
rect 498422 128258 505186 128494
rect 505422 128258 512186 128494
rect 512422 128258 519186 128494
rect 519422 128258 526186 128494
rect 526422 128258 533186 128494
rect 533422 128258 540186 128494
rect 540422 128258 547186 128494
rect 547422 128258 554186 128494
rect 554422 128258 561186 128494
rect 561422 128258 568186 128494
rect 568422 128258 575186 128494
rect 575422 128258 582186 128494
rect 582422 128258 585818 128494
rect 586054 128258 586138 128494
rect 586374 128258 586458 128494
rect 586694 128258 586778 128494
rect 587014 128258 588874 128494
rect -4950 128216 588874 128258
rect -4950 122561 588874 122603
rect -4950 122325 -4842 122561
rect -4606 122325 -4522 122561
rect -4286 122325 -4202 122561
rect -3966 122325 -3882 122561
rect -3646 122325 2918 122561
rect 3154 122325 9918 122561
rect 10154 122325 16918 122561
rect 17154 122325 23918 122561
rect 24154 122325 30918 122561
rect 31154 122325 37918 122561
rect 38154 122325 44918 122561
rect 45154 122325 51918 122561
rect 52154 122325 58918 122561
rect 59154 122325 65918 122561
rect 66154 122325 72918 122561
rect 73154 122325 79918 122561
rect 80154 122325 86918 122561
rect 87154 122325 93918 122561
rect 94154 122325 100918 122561
rect 101154 122325 107918 122561
rect 108154 122325 114918 122561
rect 115154 122325 121918 122561
rect 122154 122325 128918 122561
rect 129154 122325 135918 122561
rect 136154 122325 142918 122561
rect 143154 122325 149918 122561
rect 150154 122325 156918 122561
rect 157154 122325 163918 122561
rect 164154 122325 170918 122561
rect 171154 122325 177918 122561
rect 178154 122325 184918 122561
rect 185154 122325 191918 122561
rect 192154 122325 198918 122561
rect 199154 122325 205918 122561
rect 206154 122325 212918 122561
rect 213154 122325 219918 122561
rect 220154 122325 226918 122561
rect 227154 122325 233918 122561
rect 234154 122325 240918 122561
rect 241154 122325 247918 122561
rect 248154 122325 254918 122561
rect 255154 122325 261918 122561
rect 262154 122325 268918 122561
rect 269154 122325 275918 122561
rect 276154 122325 282918 122561
rect 283154 122325 289918 122561
rect 290154 122325 296918 122561
rect 297154 122325 303918 122561
rect 304154 122325 310918 122561
rect 311154 122325 317918 122561
rect 318154 122325 324918 122561
rect 325154 122325 331918 122561
rect 332154 122325 338918 122561
rect 339154 122325 345918 122561
rect 346154 122325 352918 122561
rect 353154 122325 359918 122561
rect 360154 122325 366918 122561
rect 367154 122325 373918 122561
rect 374154 122325 380918 122561
rect 381154 122325 387918 122561
rect 388154 122325 394918 122561
rect 395154 122325 401918 122561
rect 402154 122325 408918 122561
rect 409154 122325 415918 122561
rect 416154 122325 422918 122561
rect 423154 122325 429918 122561
rect 430154 122325 436918 122561
rect 437154 122325 443918 122561
rect 444154 122325 450918 122561
rect 451154 122325 457918 122561
rect 458154 122325 464918 122561
rect 465154 122325 471918 122561
rect 472154 122325 478918 122561
rect 479154 122325 485918 122561
rect 486154 122325 492918 122561
rect 493154 122325 499918 122561
rect 500154 122325 506918 122561
rect 507154 122325 513918 122561
rect 514154 122325 520918 122561
rect 521154 122325 527918 122561
rect 528154 122325 534918 122561
rect 535154 122325 541918 122561
rect 542154 122325 548918 122561
rect 549154 122325 555918 122561
rect 556154 122325 562918 122561
rect 563154 122325 569918 122561
rect 570154 122325 576918 122561
rect 577154 122325 587570 122561
rect 587806 122325 587890 122561
rect 588126 122325 588210 122561
rect 588446 122325 588530 122561
rect 588766 122325 588874 122561
rect -4950 122283 588874 122325
rect -4950 121494 588874 121536
rect -4950 121258 -3090 121494
rect -2854 121258 -2770 121494
rect -2534 121258 -2450 121494
rect -2214 121258 -2130 121494
rect -1894 121258 1186 121494
rect 1422 121258 8186 121494
rect 8422 121258 15186 121494
rect 15422 121258 22186 121494
rect 22422 121258 29186 121494
rect 29422 121258 36186 121494
rect 36422 121258 43186 121494
rect 43422 121258 50186 121494
rect 50422 121258 57186 121494
rect 57422 121258 64186 121494
rect 64422 121258 71186 121494
rect 71422 121258 78186 121494
rect 78422 121258 85186 121494
rect 85422 121258 92186 121494
rect 92422 121258 99186 121494
rect 99422 121258 106186 121494
rect 106422 121258 113186 121494
rect 113422 121258 120186 121494
rect 120422 121258 127186 121494
rect 127422 121258 134186 121494
rect 134422 121258 141186 121494
rect 141422 121258 148186 121494
rect 148422 121258 155186 121494
rect 155422 121258 162186 121494
rect 162422 121258 169186 121494
rect 169422 121258 176186 121494
rect 176422 121258 183186 121494
rect 183422 121258 190186 121494
rect 190422 121258 197186 121494
rect 197422 121258 204186 121494
rect 204422 121258 211186 121494
rect 211422 121258 218186 121494
rect 218422 121258 225186 121494
rect 225422 121258 232186 121494
rect 232422 121258 239186 121494
rect 239422 121258 246186 121494
rect 246422 121258 253186 121494
rect 253422 121258 260186 121494
rect 260422 121258 267186 121494
rect 267422 121258 274186 121494
rect 274422 121258 281186 121494
rect 281422 121258 288186 121494
rect 288422 121258 295186 121494
rect 295422 121258 302186 121494
rect 302422 121258 309186 121494
rect 309422 121258 316186 121494
rect 316422 121258 323186 121494
rect 323422 121258 330186 121494
rect 330422 121258 337186 121494
rect 337422 121258 344186 121494
rect 344422 121258 351186 121494
rect 351422 121258 358186 121494
rect 358422 121258 365186 121494
rect 365422 121258 372186 121494
rect 372422 121258 379186 121494
rect 379422 121258 386186 121494
rect 386422 121258 393186 121494
rect 393422 121258 400186 121494
rect 400422 121258 407186 121494
rect 407422 121258 414186 121494
rect 414422 121258 421186 121494
rect 421422 121258 428186 121494
rect 428422 121258 435186 121494
rect 435422 121258 442186 121494
rect 442422 121258 449186 121494
rect 449422 121258 456186 121494
rect 456422 121258 463186 121494
rect 463422 121258 470186 121494
rect 470422 121258 477186 121494
rect 477422 121258 484186 121494
rect 484422 121258 491186 121494
rect 491422 121258 498186 121494
rect 498422 121258 505186 121494
rect 505422 121258 512186 121494
rect 512422 121258 519186 121494
rect 519422 121258 526186 121494
rect 526422 121258 533186 121494
rect 533422 121258 540186 121494
rect 540422 121258 547186 121494
rect 547422 121258 554186 121494
rect 554422 121258 561186 121494
rect 561422 121258 568186 121494
rect 568422 121258 575186 121494
rect 575422 121258 582186 121494
rect 582422 121258 585818 121494
rect 586054 121258 586138 121494
rect 586374 121258 586458 121494
rect 586694 121258 586778 121494
rect 587014 121258 588874 121494
rect -4950 121216 588874 121258
rect -4950 115561 588874 115603
rect -4950 115325 -4842 115561
rect -4606 115325 -4522 115561
rect -4286 115325 -4202 115561
rect -3966 115325 -3882 115561
rect -3646 115325 2918 115561
rect 3154 115325 9918 115561
rect 10154 115325 16918 115561
rect 17154 115325 23918 115561
rect 24154 115325 30918 115561
rect 31154 115325 37918 115561
rect 38154 115325 44918 115561
rect 45154 115325 51918 115561
rect 52154 115325 58918 115561
rect 59154 115325 65918 115561
rect 66154 115325 72918 115561
rect 73154 115325 79918 115561
rect 80154 115325 86918 115561
rect 87154 115325 93918 115561
rect 94154 115325 100918 115561
rect 101154 115325 107918 115561
rect 108154 115325 114918 115561
rect 115154 115325 121918 115561
rect 122154 115325 128918 115561
rect 129154 115325 135918 115561
rect 136154 115325 142918 115561
rect 143154 115325 149918 115561
rect 150154 115325 156918 115561
rect 157154 115325 163918 115561
rect 164154 115325 170918 115561
rect 171154 115325 177918 115561
rect 178154 115325 184918 115561
rect 185154 115325 191918 115561
rect 192154 115325 198918 115561
rect 199154 115325 205918 115561
rect 206154 115325 212918 115561
rect 213154 115325 219918 115561
rect 220154 115325 226918 115561
rect 227154 115325 233918 115561
rect 234154 115325 240918 115561
rect 241154 115325 247918 115561
rect 248154 115325 254918 115561
rect 255154 115325 261918 115561
rect 262154 115325 268918 115561
rect 269154 115325 275918 115561
rect 276154 115325 282918 115561
rect 283154 115325 289918 115561
rect 290154 115325 296918 115561
rect 297154 115325 303918 115561
rect 304154 115325 310918 115561
rect 311154 115325 317918 115561
rect 318154 115325 324918 115561
rect 325154 115325 331918 115561
rect 332154 115325 338918 115561
rect 339154 115325 345918 115561
rect 346154 115325 352918 115561
rect 353154 115325 359918 115561
rect 360154 115325 366918 115561
rect 367154 115325 373918 115561
rect 374154 115325 380918 115561
rect 381154 115325 387918 115561
rect 388154 115325 394918 115561
rect 395154 115325 401918 115561
rect 402154 115325 408918 115561
rect 409154 115325 415918 115561
rect 416154 115325 422918 115561
rect 423154 115325 429918 115561
rect 430154 115325 436918 115561
rect 437154 115325 443918 115561
rect 444154 115325 450918 115561
rect 451154 115325 457918 115561
rect 458154 115325 464918 115561
rect 465154 115325 471918 115561
rect 472154 115325 478918 115561
rect 479154 115325 485918 115561
rect 486154 115325 492918 115561
rect 493154 115325 499918 115561
rect 500154 115325 506918 115561
rect 507154 115325 513918 115561
rect 514154 115325 520918 115561
rect 521154 115325 527918 115561
rect 528154 115325 534918 115561
rect 535154 115325 541918 115561
rect 542154 115325 548918 115561
rect 549154 115325 555918 115561
rect 556154 115325 562918 115561
rect 563154 115325 569918 115561
rect 570154 115325 576918 115561
rect 577154 115325 587570 115561
rect 587806 115325 587890 115561
rect 588126 115325 588210 115561
rect 588446 115325 588530 115561
rect 588766 115325 588874 115561
rect -4950 115283 588874 115325
rect -4950 114494 588874 114536
rect -4950 114258 -3090 114494
rect -2854 114258 -2770 114494
rect -2534 114258 -2450 114494
rect -2214 114258 -2130 114494
rect -1894 114258 1186 114494
rect 1422 114258 8186 114494
rect 8422 114258 15186 114494
rect 15422 114258 22186 114494
rect 22422 114258 29186 114494
rect 29422 114258 36186 114494
rect 36422 114258 43186 114494
rect 43422 114258 50186 114494
rect 50422 114258 57186 114494
rect 57422 114258 64186 114494
rect 64422 114258 71186 114494
rect 71422 114258 78186 114494
rect 78422 114258 85186 114494
rect 85422 114258 92186 114494
rect 92422 114258 99186 114494
rect 99422 114258 106186 114494
rect 106422 114258 113186 114494
rect 113422 114258 120186 114494
rect 120422 114258 127186 114494
rect 127422 114258 134186 114494
rect 134422 114258 141186 114494
rect 141422 114258 148186 114494
rect 148422 114258 155186 114494
rect 155422 114258 162186 114494
rect 162422 114258 169186 114494
rect 169422 114258 176186 114494
rect 176422 114258 183186 114494
rect 183422 114258 190186 114494
rect 190422 114258 197186 114494
rect 197422 114258 204186 114494
rect 204422 114258 211186 114494
rect 211422 114258 218186 114494
rect 218422 114258 225186 114494
rect 225422 114258 232186 114494
rect 232422 114258 239186 114494
rect 239422 114258 246186 114494
rect 246422 114258 253186 114494
rect 253422 114258 260186 114494
rect 260422 114258 267186 114494
rect 267422 114258 274186 114494
rect 274422 114258 281186 114494
rect 281422 114258 288186 114494
rect 288422 114258 295186 114494
rect 295422 114258 302186 114494
rect 302422 114258 309186 114494
rect 309422 114258 316186 114494
rect 316422 114258 323186 114494
rect 323422 114258 330186 114494
rect 330422 114258 337186 114494
rect 337422 114258 344186 114494
rect 344422 114258 351186 114494
rect 351422 114258 358186 114494
rect 358422 114258 365186 114494
rect 365422 114258 372186 114494
rect 372422 114258 379186 114494
rect 379422 114258 386186 114494
rect 386422 114258 393186 114494
rect 393422 114258 400186 114494
rect 400422 114258 407186 114494
rect 407422 114258 414186 114494
rect 414422 114258 421186 114494
rect 421422 114258 428186 114494
rect 428422 114258 435186 114494
rect 435422 114258 442186 114494
rect 442422 114258 449186 114494
rect 449422 114258 456186 114494
rect 456422 114258 463186 114494
rect 463422 114258 470186 114494
rect 470422 114258 477186 114494
rect 477422 114258 484186 114494
rect 484422 114258 491186 114494
rect 491422 114258 498186 114494
rect 498422 114258 505186 114494
rect 505422 114258 512186 114494
rect 512422 114258 519186 114494
rect 519422 114258 526186 114494
rect 526422 114258 533186 114494
rect 533422 114258 540186 114494
rect 540422 114258 547186 114494
rect 547422 114258 554186 114494
rect 554422 114258 561186 114494
rect 561422 114258 568186 114494
rect 568422 114258 575186 114494
rect 575422 114258 582186 114494
rect 582422 114258 585818 114494
rect 586054 114258 586138 114494
rect 586374 114258 586458 114494
rect 586694 114258 586778 114494
rect 587014 114258 588874 114494
rect -4950 114216 588874 114258
rect -4950 108561 588874 108603
rect -4950 108325 -4842 108561
rect -4606 108325 -4522 108561
rect -4286 108325 -4202 108561
rect -3966 108325 -3882 108561
rect -3646 108325 2918 108561
rect 3154 108325 9918 108561
rect 10154 108325 16918 108561
rect 17154 108325 23918 108561
rect 24154 108325 30918 108561
rect 31154 108325 37918 108561
rect 38154 108325 44918 108561
rect 45154 108325 51918 108561
rect 52154 108325 58918 108561
rect 59154 108325 65918 108561
rect 66154 108325 72918 108561
rect 73154 108325 79918 108561
rect 80154 108325 86918 108561
rect 87154 108325 93918 108561
rect 94154 108325 100918 108561
rect 101154 108325 107918 108561
rect 108154 108325 114918 108561
rect 115154 108325 121918 108561
rect 122154 108325 128918 108561
rect 129154 108325 135918 108561
rect 136154 108325 142918 108561
rect 143154 108325 149918 108561
rect 150154 108325 156918 108561
rect 157154 108325 163918 108561
rect 164154 108325 170918 108561
rect 171154 108325 177918 108561
rect 178154 108325 184918 108561
rect 185154 108325 191918 108561
rect 192154 108325 198918 108561
rect 199154 108325 205918 108561
rect 206154 108325 212918 108561
rect 213154 108325 219918 108561
rect 220154 108325 226918 108561
rect 227154 108325 233918 108561
rect 234154 108325 240918 108561
rect 241154 108325 247918 108561
rect 248154 108325 254918 108561
rect 255154 108325 261918 108561
rect 262154 108325 268918 108561
rect 269154 108325 275918 108561
rect 276154 108325 282918 108561
rect 283154 108325 289918 108561
rect 290154 108325 296918 108561
rect 297154 108325 303918 108561
rect 304154 108325 310918 108561
rect 311154 108325 317918 108561
rect 318154 108325 324918 108561
rect 325154 108325 331918 108561
rect 332154 108325 338918 108561
rect 339154 108325 345918 108561
rect 346154 108325 352918 108561
rect 353154 108325 359918 108561
rect 360154 108325 366918 108561
rect 367154 108325 373918 108561
rect 374154 108325 380918 108561
rect 381154 108325 387918 108561
rect 388154 108325 394918 108561
rect 395154 108325 401918 108561
rect 402154 108325 408918 108561
rect 409154 108325 415918 108561
rect 416154 108325 422918 108561
rect 423154 108325 429918 108561
rect 430154 108325 436918 108561
rect 437154 108325 443918 108561
rect 444154 108325 450918 108561
rect 451154 108325 457918 108561
rect 458154 108325 464918 108561
rect 465154 108325 471918 108561
rect 472154 108325 478918 108561
rect 479154 108325 485918 108561
rect 486154 108325 492918 108561
rect 493154 108325 499918 108561
rect 500154 108325 506918 108561
rect 507154 108325 513918 108561
rect 514154 108325 520918 108561
rect 521154 108325 527918 108561
rect 528154 108325 534918 108561
rect 535154 108325 541918 108561
rect 542154 108325 548918 108561
rect 549154 108325 555918 108561
rect 556154 108325 562918 108561
rect 563154 108325 569918 108561
rect 570154 108325 576918 108561
rect 577154 108325 587570 108561
rect 587806 108325 587890 108561
rect 588126 108325 588210 108561
rect 588446 108325 588530 108561
rect 588766 108325 588874 108561
rect -4950 108283 588874 108325
rect -4950 107494 588874 107536
rect -4950 107258 -3090 107494
rect -2854 107258 -2770 107494
rect -2534 107258 -2450 107494
rect -2214 107258 -2130 107494
rect -1894 107258 1186 107494
rect 1422 107258 8186 107494
rect 8422 107258 15186 107494
rect 15422 107258 22186 107494
rect 22422 107258 29186 107494
rect 29422 107258 36186 107494
rect 36422 107258 43186 107494
rect 43422 107258 50186 107494
rect 50422 107258 57186 107494
rect 57422 107258 64186 107494
rect 64422 107258 71186 107494
rect 71422 107258 78186 107494
rect 78422 107258 85186 107494
rect 85422 107258 92186 107494
rect 92422 107258 99186 107494
rect 99422 107258 106186 107494
rect 106422 107258 113186 107494
rect 113422 107258 120186 107494
rect 120422 107258 127186 107494
rect 127422 107258 134186 107494
rect 134422 107258 141186 107494
rect 141422 107258 148186 107494
rect 148422 107258 155186 107494
rect 155422 107258 162186 107494
rect 162422 107258 169186 107494
rect 169422 107258 176186 107494
rect 176422 107258 183186 107494
rect 183422 107258 190186 107494
rect 190422 107258 197186 107494
rect 197422 107258 204186 107494
rect 204422 107258 211186 107494
rect 211422 107258 218186 107494
rect 218422 107258 225186 107494
rect 225422 107258 232186 107494
rect 232422 107258 239186 107494
rect 239422 107258 246186 107494
rect 246422 107258 253186 107494
rect 253422 107258 260186 107494
rect 260422 107258 267186 107494
rect 267422 107258 274186 107494
rect 274422 107258 281186 107494
rect 281422 107258 288186 107494
rect 288422 107258 295186 107494
rect 295422 107258 302186 107494
rect 302422 107258 309186 107494
rect 309422 107258 316186 107494
rect 316422 107258 323186 107494
rect 323422 107258 330186 107494
rect 330422 107258 337186 107494
rect 337422 107258 344186 107494
rect 344422 107258 351186 107494
rect 351422 107258 358186 107494
rect 358422 107258 365186 107494
rect 365422 107258 372186 107494
rect 372422 107258 379186 107494
rect 379422 107258 386186 107494
rect 386422 107258 393186 107494
rect 393422 107258 400186 107494
rect 400422 107258 407186 107494
rect 407422 107258 414186 107494
rect 414422 107258 421186 107494
rect 421422 107258 428186 107494
rect 428422 107258 435186 107494
rect 435422 107258 442186 107494
rect 442422 107258 449186 107494
rect 449422 107258 456186 107494
rect 456422 107258 463186 107494
rect 463422 107258 470186 107494
rect 470422 107258 477186 107494
rect 477422 107258 484186 107494
rect 484422 107258 491186 107494
rect 491422 107258 498186 107494
rect 498422 107258 505186 107494
rect 505422 107258 512186 107494
rect 512422 107258 519186 107494
rect 519422 107258 526186 107494
rect 526422 107258 533186 107494
rect 533422 107258 540186 107494
rect 540422 107258 547186 107494
rect 547422 107258 554186 107494
rect 554422 107258 561186 107494
rect 561422 107258 568186 107494
rect 568422 107258 575186 107494
rect 575422 107258 582186 107494
rect 582422 107258 585818 107494
rect 586054 107258 586138 107494
rect 586374 107258 586458 107494
rect 586694 107258 586778 107494
rect 587014 107258 588874 107494
rect -4950 107216 588874 107258
rect -4950 101561 588874 101603
rect -4950 101325 -4842 101561
rect -4606 101325 -4522 101561
rect -4286 101325 -4202 101561
rect -3966 101325 -3882 101561
rect -3646 101325 2918 101561
rect 3154 101325 9918 101561
rect 10154 101325 16918 101561
rect 17154 101325 23918 101561
rect 24154 101325 30918 101561
rect 31154 101325 37918 101561
rect 38154 101325 44918 101561
rect 45154 101325 51918 101561
rect 52154 101325 58918 101561
rect 59154 101325 65918 101561
rect 66154 101325 72918 101561
rect 73154 101325 79918 101561
rect 80154 101325 86918 101561
rect 87154 101325 93918 101561
rect 94154 101325 100918 101561
rect 101154 101325 107918 101561
rect 108154 101325 114918 101561
rect 115154 101325 121918 101561
rect 122154 101325 128918 101561
rect 129154 101325 135918 101561
rect 136154 101325 142918 101561
rect 143154 101325 149918 101561
rect 150154 101325 156918 101561
rect 157154 101325 163918 101561
rect 164154 101325 170918 101561
rect 171154 101325 177918 101561
rect 178154 101325 184918 101561
rect 185154 101325 191918 101561
rect 192154 101325 198918 101561
rect 199154 101325 205918 101561
rect 206154 101325 212918 101561
rect 213154 101325 219918 101561
rect 220154 101325 226918 101561
rect 227154 101325 233918 101561
rect 234154 101325 240918 101561
rect 241154 101325 247918 101561
rect 248154 101325 254918 101561
rect 255154 101325 261918 101561
rect 262154 101325 268918 101561
rect 269154 101325 275918 101561
rect 276154 101325 282918 101561
rect 283154 101325 289918 101561
rect 290154 101325 296918 101561
rect 297154 101325 303918 101561
rect 304154 101325 310918 101561
rect 311154 101325 317918 101561
rect 318154 101325 324918 101561
rect 325154 101325 331918 101561
rect 332154 101325 338918 101561
rect 339154 101325 345918 101561
rect 346154 101325 352918 101561
rect 353154 101325 359918 101561
rect 360154 101325 366918 101561
rect 367154 101325 373918 101561
rect 374154 101325 380918 101561
rect 381154 101325 387918 101561
rect 388154 101325 394918 101561
rect 395154 101325 401918 101561
rect 402154 101325 408918 101561
rect 409154 101325 415918 101561
rect 416154 101325 422918 101561
rect 423154 101325 429918 101561
rect 430154 101325 436918 101561
rect 437154 101325 443918 101561
rect 444154 101325 450918 101561
rect 451154 101325 457918 101561
rect 458154 101325 464918 101561
rect 465154 101325 471918 101561
rect 472154 101325 478918 101561
rect 479154 101325 485918 101561
rect 486154 101325 492918 101561
rect 493154 101325 499918 101561
rect 500154 101325 506918 101561
rect 507154 101325 513918 101561
rect 514154 101325 520918 101561
rect 521154 101325 527918 101561
rect 528154 101325 534918 101561
rect 535154 101325 541918 101561
rect 542154 101325 548918 101561
rect 549154 101325 555918 101561
rect 556154 101325 562918 101561
rect 563154 101325 569918 101561
rect 570154 101325 576918 101561
rect 577154 101325 587570 101561
rect 587806 101325 587890 101561
rect 588126 101325 588210 101561
rect 588446 101325 588530 101561
rect 588766 101325 588874 101561
rect -4950 101283 588874 101325
rect -4950 100494 588874 100536
rect -4950 100258 -3090 100494
rect -2854 100258 -2770 100494
rect -2534 100258 -2450 100494
rect -2214 100258 -2130 100494
rect -1894 100258 1186 100494
rect 1422 100258 8186 100494
rect 8422 100258 15186 100494
rect 15422 100258 22186 100494
rect 22422 100258 29186 100494
rect 29422 100258 36186 100494
rect 36422 100258 43186 100494
rect 43422 100258 50186 100494
rect 50422 100258 57186 100494
rect 57422 100258 64186 100494
rect 64422 100258 71186 100494
rect 71422 100258 78186 100494
rect 78422 100258 85186 100494
rect 85422 100258 92186 100494
rect 92422 100258 99186 100494
rect 99422 100258 106186 100494
rect 106422 100258 113186 100494
rect 113422 100258 120186 100494
rect 120422 100258 127186 100494
rect 127422 100258 134186 100494
rect 134422 100258 141186 100494
rect 141422 100258 148186 100494
rect 148422 100258 155186 100494
rect 155422 100258 162186 100494
rect 162422 100258 169186 100494
rect 169422 100258 176186 100494
rect 176422 100258 183186 100494
rect 183422 100258 190186 100494
rect 190422 100258 197186 100494
rect 197422 100258 204186 100494
rect 204422 100258 211186 100494
rect 211422 100258 218186 100494
rect 218422 100258 225186 100494
rect 225422 100258 232186 100494
rect 232422 100258 239186 100494
rect 239422 100258 246186 100494
rect 246422 100258 253186 100494
rect 253422 100258 260186 100494
rect 260422 100258 267186 100494
rect 267422 100258 274186 100494
rect 274422 100258 281186 100494
rect 281422 100258 288186 100494
rect 288422 100258 295186 100494
rect 295422 100258 302186 100494
rect 302422 100258 309186 100494
rect 309422 100258 316186 100494
rect 316422 100258 323186 100494
rect 323422 100258 330186 100494
rect 330422 100258 337186 100494
rect 337422 100258 344186 100494
rect 344422 100258 351186 100494
rect 351422 100258 358186 100494
rect 358422 100258 365186 100494
rect 365422 100258 372186 100494
rect 372422 100258 379186 100494
rect 379422 100258 386186 100494
rect 386422 100258 393186 100494
rect 393422 100258 400186 100494
rect 400422 100258 407186 100494
rect 407422 100258 414186 100494
rect 414422 100258 421186 100494
rect 421422 100258 428186 100494
rect 428422 100258 435186 100494
rect 435422 100258 442186 100494
rect 442422 100258 449186 100494
rect 449422 100258 456186 100494
rect 456422 100258 463186 100494
rect 463422 100258 470186 100494
rect 470422 100258 477186 100494
rect 477422 100258 484186 100494
rect 484422 100258 491186 100494
rect 491422 100258 498186 100494
rect 498422 100258 505186 100494
rect 505422 100258 512186 100494
rect 512422 100258 519186 100494
rect 519422 100258 526186 100494
rect 526422 100258 533186 100494
rect 533422 100258 540186 100494
rect 540422 100258 547186 100494
rect 547422 100258 554186 100494
rect 554422 100258 561186 100494
rect 561422 100258 568186 100494
rect 568422 100258 575186 100494
rect 575422 100258 582186 100494
rect 582422 100258 585818 100494
rect 586054 100258 586138 100494
rect 586374 100258 586458 100494
rect 586694 100258 586778 100494
rect 587014 100258 588874 100494
rect -4950 100216 588874 100258
rect -4950 94561 588874 94603
rect -4950 94325 -4842 94561
rect -4606 94325 -4522 94561
rect -4286 94325 -4202 94561
rect -3966 94325 -3882 94561
rect -3646 94325 2918 94561
rect 3154 94325 9918 94561
rect 10154 94325 16918 94561
rect 17154 94325 23918 94561
rect 24154 94325 30918 94561
rect 31154 94325 37918 94561
rect 38154 94325 44918 94561
rect 45154 94325 51918 94561
rect 52154 94325 58918 94561
rect 59154 94325 65918 94561
rect 66154 94325 72918 94561
rect 73154 94325 79918 94561
rect 80154 94325 86918 94561
rect 87154 94325 93918 94561
rect 94154 94325 100918 94561
rect 101154 94325 107918 94561
rect 108154 94325 114918 94561
rect 115154 94325 121918 94561
rect 122154 94325 128918 94561
rect 129154 94325 135918 94561
rect 136154 94325 142918 94561
rect 143154 94325 149918 94561
rect 150154 94325 156918 94561
rect 157154 94325 163918 94561
rect 164154 94325 170918 94561
rect 171154 94325 177918 94561
rect 178154 94325 184918 94561
rect 185154 94325 191918 94561
rect 192154 94325 198918 94561
rect 199154 94325 205918 94561
rect 206154 94325 212918 94561
rect 213154 94325 219918 94561
rect 220154 94325 226918 94561
rect 227154 94325 233918 94561
rect 234154 94325 240918 94561
rect 241154 94325 247918 94561
rect 248154 94325 254918 94561
rect 255154 94325 261918 94561
rect 262154 94325 268918 94561
rect 269154 94325 275918 94561
rect 276154 94325 282918 94561
rect 283154 94325 289918 94561
rect 290154 94325 296918 94561
rect 297154 94325 303918 94561
rect 304154 94325 310918 94561
rect 311154 94325 317918 94561
rect 318154 94325 324918 94561
rect 325154 94325 331918 94561
rect 332154 94325 338918 94561
rect 339154 94325 345918 94561
rect 346154 94325 352918 94561
rect 353154 94325 359918 94561
rect 360154 94325 366918 94561
rect 367154 94325 373918 94561
rect 374154 94325 380918 94561
rect 381154 94325 387918 94561
rect 388154 94325 394918 94561
rect 395154 94325 401918 94561
rect 402154 94325 408918 94561
rect 409154 94325 415918 94561
rect 416154 94325 422918 94561
rect 423154 94325 429918 94561
rect 430154 94325 436918 94561
rect 437154 94325 443918 94561
rect 444154 94325 450918 94561
rect 451154 94325 457918 94561
rect 458154 94325 464918 94561
rect 465154 94325 471918 94561
rect 472154 94325 478918 94561
rect 479154 94325 485918 94561
rect 486154 94325 492918 94561
rect 493154 94325 499918 94561
rect 500154 94325 506918 94561
rect 507154 94325 513918 94561
rect 514154 94325 520918 94561
rect 521154 94325 527918 94561
rect 528154 94325 534918 94561
rect 535154 94325 541918 94561
rect 542154 94325 548918 94561
rect 549154 94325 555918 94561
rect 556154 94325 562918 94561
rect 563154 94325 569918 94561
rect 570154 94325 576918 94561
rect 577154 94325 587570 94561
rect 587806 94325 587890 94561
rect 588126 94325 588210 94561
rect 588446 94325 588530 94561
rect 588766 94325 588874 94561
rect -4950 94283 588874 94325
rect -4950 93494 588874 93536
rect -4950 93258 -3090 93494
rect -2854 93258 -2770 93494
rect -2534 93258 -2450 93494
rect -2214 93258 -2130 93494
rect -1894 93258 1186 93494
rect 1422 93258 8186 93494
rect 8422 93258 15186 93494
rect 15422 93258 22186 93494
rect 22422 93258 29186 93494
rect 29422 93258 36186 93494
rect 36422 93258 43186 93494
rect 43422 93258 50186 93494
rect 50422 93258 57186 93494
rect 57422 93258 64186 93494
rect 64422 93258 71186 93494
rect 71422 93258 78186 93494
rect 78422 93258 85186 93494
rect 85422 93258 92186 93494
rect 92422 93258 99186 93494
rect 99422 93258 106186 93494
rect 106422 93258 113186 93494
rect 113422 93258 120186 93494
rect 120422 93258 127186 93494
rect 127422 93258 134186 93494
rect 134422 93258 141186 93494
rect 141422 93258 148186 93494
rect 148422 93258 155186 93494
rect 155422 93258 162186 93494
rect 162422 93258 169186 93494
rect 169422 93258 176186 93494
rect 176422 93258 183186 93494
rect 183422 93258 190186 93494
rect 190422 93258 197186 93494
rect 197422 93258 204186 93494
rect 204422 93258 211186 93494
rect 211422 93258 218186 93494
rect 218422 93258 225186 93494
rect 225422 93258 232186 93494
rect 232422 93258 239186 93494
rect 239422 93258 246186 93494
rect 246422 93258 253186 93494
rect 253422 93258 260186 93494
rect 260422 93258 267186 93494
rect 267422 93258 274186 93494
rect 274422 93258 281186 93494
rect 281422 93258 288186 93494
rect 288422 93258 295186 93494
rect 295422 93258 302186 93494
rect 302422 93258 309186 93494
rect 309422 93258 316186 93494
rect 316422 93258 323186 93494
rect 323422 93258 330186 93494
rect 330422 93258 337186 93494
rect 337422 93258 344186 93494
rect 344422 93258 351186 93494
rect 351422 93258 358186 93494
rect 358422 93258 365186 93494
rect 365422 93258 372186 93494
rect 372422 93258 379186 93494
rect 379422 93258 386186 93494
rect 386422 93258 393186 93494
rect 393422 93258 400186 93494
rect 400422 93258 407186 93494
rect 407422 93258 414186 93494
rect 414422 93258 421186 93494
rect 421422 93258 428186 93494
rect 428422 93258 435186 93494
rect 435422 93258 442186 93494
rect 442422 93258 449186 93494
rect 449422 93258 456186 93494
rect 456422 93258 463186 93494
rect 463422 93258 470186 93494
rect 470422 93258 477186 93494
rect 477422 93258 484186 93494
rect 484422 93258 491186 93494
rect 491422 93258 498186 93494
rect 498422 93258 505186 93494
rect 505422 93258 512186 93494
rect 512422 93258 519186 93494
rect 519422 93258 526186 93494
rect 526422 93258 533186 93494
rect 533422 93258 540186 93494
rect 540422 93258 547186 93494
rect 547422 93258 554186 93494
rect 554422 93258 561186 93494
rect 561422 93258 568186 93494
rect 568422 93258 575186 93494
rect 575422 93258 582186 93494
rect 582422 93258 585818 93494
rect 586054 93258 586138 93494
rect 586374 93258 586458 93494
rect 586694 93258 586778 93494
rect 587014 93258 588874 93494
rect -4950 93216 588874 93258
rect -4950 87561 588874 87603
rect -4950 87325 -4842 87561
rect -4606 87325 -4522 87561
rect -4286 87325 -4202 87561
rect -3966 87325 -3882 87561
rect -3646 87325 2918 87561
rect 3154 87325 9918 87561
rect 10154 87325 16918 87561
rect 17154 87325 23918 87561
rect 24154 87325 30918 87561
rect 31154 87325 37918 87561
rect 38154 87325 44918 87561
rect 45154 87325 51918 87561
rect 52154 87325 58918 87561
rect 59154 87325 65918 87561
rect 66154 87325 72918 87561
rect 73154 87325 79918 87561
rect 80154 87325 86918 87561
rect 87154 87325 93918 87561
rect 94154 87325 100918 87561
rect 101154 87325 107918 87561
rect 108154 87325 114918 87561
rect 115154 87325 121918 87561
rect 122154 87325 128918 87561
rect 129154 87325 135918 87561
rect 136154 87325 142918 87561
rect 143154 87325 149918 87561
rect 150154 87325 156918 87561
rect 157154 87325 163918 87561
rect 164154 87325 170918 87561
rect 171154 87325 177918 87561
rect 178154 87325 184918 87561
rect 185154 87325 191918 87561
rect 192154 87325 198918 87561
rect 199154 87325 205918 87561
rect 206154 87325 212918 87561
rect 213154 87325 219918 87561
rect 220154 87325 226918 87561
rect 227154 87325 233918 87561
rect 234154 87325 240918 87561
rect 241154 87325 247918 87561
rect 248154 87325 254918 87561
rect 255154 87325 261918 87561
rect 262154 87325 268918 87561
rect 269154 87325 275918 87561
rect 276154 87325 282918 87561
rect 283154 87325 289918 87561
rect 290154 87325 296918 87561
rect 297154 87325 303918 87561
rect 304154 87325 310918 87561
rect 311154 87325 317918 87561
rect 318154 87325 324918 87561
rect 325154 87325 331918 87561
rect 332154 87325 338918 87561
rect 339154 87325 345918 87561
rect 346154 87325 352918 87561
rect 353154 87325 359918 87561
rect 360154 87325 366918 87561
rect 367154 87325 373918 87561
rect 374154 87325 380918 87561
rect 381154 87325 387918 87561
rect 388154 87325 394918 87561
rect 395154 87325 401918 87561
rect 402154 87325 408918 87561
rect 409154 87325 415918 87561
rect 416154 87325 422918 87561
rect 423154 87325 429918 87561
rect 430154 87325 436918 87561
rect 437154 87325 443918 87561
rect 444154 87325 450918 87561
rect 451154 87325 457918 87561
rect 458154 87325 464918 87561
rect 465154 87325 471918 87561
rect 472154 87325 478918 87561
rect 479154 87325 485918 87561
rect 486154 87325 492918 87561
rect 493154 87325 499918 87561
rect 500154 87325 506918 87561
rect 507154 87325 513918 87561
rect 514154 87325 520918 87561
rect 521154 87325 527918 87561
rect 528154 87325 534918 87561
rect 535154 87325 541918 87561
rect 542154 87325 548918 87561
rect 549154 87325 555918 87561
rect 556154 87325 562918 87561
rect 563154 87325 569918 87561
rect 570154 87325 576918 87561
rect 577154 87325 587570 87561
rect 587806 87325 587890 87561
rect 588126 87325 588210 87561
rect 588446 87325 588530 87561
rect 588766 87325 588874 87561
rect -4950 87283 588874 87325
rect -4950 86494 588874 86536
rect -4950 86258 -3090 86494
rect -2854 86258 -2770 86494
rect -2534 86258 -2450 86494
rect -2214 86258 -2130 86494
rect -1894 86258 1186 86494
rect 1422 86258 8186 86494
rect 8422 86258 15186 86494
rect 15422 86258 22186 86494
rect 22422 86258 29186 86494
rect 29422 86258 36186 86494
rect 36422 86258 43186 86494
rect 43422 86258 50186 86494
rect 50422 86258 57186 86494
rect 57422 86258 64186 86494
rect 64422 86258 71186 86494
rect 71422 86258 78186 86494
rect 78422 86258 85186 86494
rect 85422 86258 92186 86494
rect 92422 86258 99186 86494
rect 99422 86258 106186 86494
rect 106422 86258 113186 86494
rect 113422 86258 120186 86494
rect 120422 86258 127186 86494
rect 127422 86258 134186 86494
rect 134422 86258 141186 86494
rect 141422 86258 148186 86494
rect 148422 86258 155186 86494
rect 155422 86258 162186 86494
rect 162422 86258 169186 86494
rect 169422 86258 176186 86494
rect 176422 86258 183186 86494
rect 183422 86258 190186 86494
rect 190422 86258 197186 86494
rect 197422 86258 204186 86494
rect 204422 86258 211186 86494
rect 211422 86258 218186 86494
rect 218422 86258 225186 86494
rect 225422 86258 232186 86494
rect 232422 86258 239186 86494
rect 239422 86258 246186 86494
rect 246422 86258 253186 86494
rect 253422 86258 260186 86494
rect 260422 86258 267186 86494
rect 267422 86258 274186 86494
rect 274422 86258 281186 86494
rect 281422 86258 288186 86494
rect 288422 86258 295186 86494
rect 295422 86258 302186 86494
rect 302422 86258 309186 86494
rect 309422 86258 316186 86494
rect 316422 86258 323186 86494
rect 323422 86258 330186 86494
rect 330422 86258 337186 86494
rect 337422 86258 344186 86494
rect 344422 86258 351186 86494
rect 351422 86258 358186 86494
rect 358422 86258 365186 86494
rect 365422 86258 372186 86494
rect 372422 86258 379186 86494
rect 379422 86258 386186 86494
rect 386422 86258 393186 86494
rect 393422 86258 400186 86494
rect 400422 86258 407186 86494
rect 407422 86258 414186 86494
rect 414422 86258 421186 86494
rect 421422 86258 428186 86494
rect 428422 86258 435186 86494
rect 435422 86258 442186 86494
rect 442422 86258 449186 86494
rect 449422 86258 456186 86494
rect 456422 86258 463186 86494
rect 463422 86258 470186 86494
rect 470422 86258 477186 86494
rect 477422 86258 484186 86494
rect 484422 86258 491186 86494
rect 491422 86258 498186 86494
rect 498422 86258 505186 86494
rect 505422 86258 512186 86494
rect 512422 86258 519186 86494
rect 519422 86258 526186 86494
rect 526422 86258 533186 86494
rect 533422 86258 540186 86494
rect 540422 86258 547186 86494
rect 547422 86258 554186 86494
rect 554422 86258 561186 86494
rect 561422 86258 568186 86494
rect 568422 86258 575186 86494
rect 575422 86258 582186 86494
rect 582422 86258 585818 86494
rect 586054 86258 586138 86494
rect 586374 86258 586458 86494
rect 586694 86258 586778 86494
rect 587014 86258 588874 86494
rect -4950 86216 588874 86258
rect -4950 80561 588874 80603
rect -4950 80325 -4842 80561
rect -4606 80325 -4522 80561
rect -4286 80325 -4202 80561
rect -3966 80325 -3882 80561
rect -3646 80325 2918 80561
rect 3154 80325 9918 80561
rect 10154 80325 16918 80561
rect 17154 80325 23918 80561
rect 24154 80325 30918 80561
rect 31154 80325 37918 80561
rect 38154 80325 44918 80561
rect 45154 80325 51918 80561
rect 52154 80325 58918 80561
rect 59154 80325 65918 80561
rect 66154 80325 72918 80561
rect 73154 80325 79918 80561
rect 80154 80325 86918 80561
rect 87154 80325 93918 80561
rect 94154 80325 100918 80561
rect 101154 80325 107918 80561
rect 108154 80325 114918 80561
rect 115154 80325 121918 80561
rect 122154 80325 128918 80561
rect 129154 80325 135918 80561
rect 136154 80325 142918 80561
rect 143154 80325 149918 80561
rect 150154 80325 156918 80561
rect 157154 80325 163918 80561
rect 164154 80325 170918 80561
rect 171154 80325 177918 80561
rect 178154 80325 184918 80561
rect 185154 80325 191918 80561
rect 192154 80325 198918 80561
rect 199154 80325 205918 80561
rect 206154 80325 212918 80561
rect 213154 80325 219918 80561
rect 220154 80325 226918 80561
rect 227154 80325 233918 80561
rect 234154 80325 240918 80561
rect 241154 80325 247918 80561
rect 248154 80325 254918 80561
rect 255154 80325 261918 80561
rect 262154 80325 268918 80561
rect 269154 80325 275918 80561
rect 276154 80325 282918 80561
rect 283154 80325 289918 80561
rect 290154 80325 296918 80561
rect 297154 80325 303918 80561
rect 304154 80325 310918 80561
rect 311154 80325 317918 80561
rect 318154 80325 324918 80561
rect 325154 80325 331918 80561
rect 332154 80325 338918 80561
rect 339154 80325 345918 80561
rect 346154 80325 352918 80561
rect 353154 80325 359918 80561
rect 360154 80325 366918 80561
rect 367154 80325 373918 80561
rect 374154 80325 380918 80561
rect 381154 80325 387918 80561
rect 388154 80325 394918 80561
rect 395154 80325 401918 80561
rect 402154 80325 408918 80561
rect 409154 80325 415918 80561
rect 416154 80325 422918 80561
rect 423154 80325 429918 80561
rect 430154 80325 436918 80561
rect 437154 80325 443918 80561
rect 444154 80325 450918 80561
rect 451154 80325 457918 80561
rect 458154 80325 464918 80561
rect 465154 80325 471918 80561
rect 472154 80325 478918 80561
rect 479154 80325 485918 80561
rect 486154 80325 492918 80561
rect 493154 80325 499918 80561
rect 500154 80325 506918 80561
rect 507154 80325 513918 80561
rect 514154 80325 520918 80561
rect 521154 80325 527918 80561
rect 528154 80325 534918 80561
rect 535154 80325 541918 80561
rect 542154 80325 548918 80561
rect 549154 80325 555918 80561
rect 556154 80325 562918 80561
rect 563154 80325 569918 80561
rect 570154 80325 576918 80561
rect 577154 80325 587570 80561
rect 587806 80325 587890 80561
rect 588126 80325 588210 80561
rect 588446 80325 588530 80561
rect 588766 80325 588874 80561
rect -4950 80283 588874 80325
rect -4950 79494 588874 79536
rect -4950 79258 -3090 79494
rect -2854 79258 -2770 79494
rect -2534 79258 -2450 79494
rect -2214 79258 -2130 79494
rect -1894 79258 1186 79494
rect 1422 79258 8186 79494
rect 8422 79258 15186 79494
rect 15422 79258 22186 79494
rect 22422 79258 29186 79494
rect 29422 79258 36186 79494
rect 36422 79258 43186 79494
rect 43422 79258 50186 79494
rect 50422 79258 57186 79494
rect 57422 79258 64186 79494
rect 64422 79258 71186 79494
rect 71422 79258 78186 79494
rect 78422 79258 85186 79494
rect 85422 79258 92186 79494
rect 92422 79258 99186 79494
rect 99422 79258 106186 79494
rect 106422 79258 113186 79494
rect 113422 79258 120186 79494
rect 120422 79258 127186 79494
rect 127422 79258 134186 79494
rect 134422 79258 141186 79494
rect 141422 79258 148186 79494
rect 148422 79258 155186 79494
rect 155422 79258 162186 79494
rect 162422 79258 169186 79494
rect 169422 79258 176186 79494
rect 176422 79258 183186 79494
rect 183422 79258 190186 79494
rect 190422 79258 197186 79494
rect 197422 79258 204186 79494
rect 204422 79258 211186 79494
rect 211422 79258 218186 79494
rect 218422 79258 225186 79494
rect 225422 79258 232186 79494
rect 232422 79258 239186 79494
rect 239422 79258 246186 79494
rect 246422 79258 253186 79494
rect 253422 79258 260186 79494
rect 260422 79258 267186 79494
rect 267422 79258 274186 79494
rect 274422 79258 281186 79494
rect 281422 79258 288186 79494
rect 288422 79258 295186 79494
rect 295422 79258 302186 79494
rect 302422 79258 309186 79494
rect 309422 79258 316186 79494
rect 316422 79258 323186 79494
rect 323422 79258 330186 79494
rect 330422 79258 337186 79494
rect 337422 79258 344186 79494
rect 344422 79258 351186 79494
rect 351422 79258 358186 79494
rect 358422 79258 365186 79494
rect 365422 79258 372186 79494
rect 372422 79258 379186 79494
rect 379422 79258 386186 79494
rect 386422 79258 393186 79494
rect 393422 79258 400186 79494
rect 400422 79258 407186 79494
rect 407422 79258 414186 79494
rect 414422 79258 421186 79494
rect 421422 79258 428186 79494
rect 428422 79258 435186 79494
rect 435422 79258 442186 79494
rect 442422 79258 449186 79494
rect 449422 79258 456186 79494
rect 456422 79258 463186 79494
rect 463422 79258 470186 79494
rect 470422 79258 477186 79494
rect 477422 79258 484186 79494
rect 484422 79258 491186 79494
rect 491422 79258 498186 79494
rect 498422 79258 505186 79494
rect 505422 79258 512186 79494
rect 512422 79258 519186 79494
rect 519422 79258 526186 79494
rect 526422 79258 533186 79494
rect 533422 79258 540186 79494
rect 540422 79258 547186 79494
rect 547422 79258 554186 79494
rect 554422 79258 561186 79494
rect 561422 79258 568186 79494
rect 568422 79258 575186 79494
rect 575422 79258 582186 79494
rect 582422 79258 585818 79494
rect 586054 79258 586138 79494
rect 586374 79258 586458 79494
rect 586694 79258 586778 79494
rect 587014 79258 588874 79494
rect -4950 79216 588874 79258
rect -4950 73561 588874 73603
rect -4950 73325 -4842 73561
rect -4606 73325 -4522 73561
rect -4286 73325 -4202 73561
rect -3966 73325 -3882 73561
rect -3646 73325 2918 73561
rect 3154 73325 9918 73561
rect 10154 73325 16918 73561
rect 17154 73325 23918 73561
rect 24154 73325 30918 73561
rect 31154 73325 37918 73561
rect 38154 73325 44918 73561
rect 45154 73325 51918 73561
rect 52154 73325 58918 73561
rect 59154 73325 65918 73561
rect 66154 73325 72918 73561
rect 73154 73325 79918 73561
rect 80154 73325 86918 73561
rect 87154 73325 93918 73561
rect 94154 73325 100918 73561
rect 101154 73325 107918 73561
rect 108154 73325 114918 73561
rect 115154 73325 121918 73561
rect 122154 73325 128918 73561
rect 129154 73325 135918 73561
rect 136154 73325 142918 73561
rect 143154 73325 149918 73561
rect 150154 73325 156918 73561
rect 157154 73325 163918 73561
rect 164154 73325 170918 73561
rect 171154 73325 177918 73561
rect 178154 73325 184918 73561
rect 185154 73325 191918 73561
rect 192154 73325 198918 73561
rect 199154 73325 205918 73561
rect 206154 73325 212918 73561
rect 213154 73325 219918 73561
rect 220154 73325 226918 73561
rect 227154 73325 233918 73561
rect 234154 73325 240918 73561
rect 241154 73325 247918 73561
rect 248154 73325 254918 73561
rect 255154 73325 261918 73561
rect 262154 73325 268918 73561
rect 269154 73325 275918 73561
rect 276154 73325 282918 73561
rect 283154 73325 289918 73561
rect 290154 73325 296918 73561
rect 297154 73325 303918 73561
rect 304154 73325 310918 73561
rect 311154 73325 317918 73561
rect 318154 73325 324918 73561
rect 325154 73325 331918 73561
rect 332154 73325 338918 73561
rect 339154 73325 345918 73561
rect 346154 73325 352918 73561
rect 353154 73325 359918 73561
rect 360154 73325 366918 73561
rect 367154 73325 373918 73561
rect 374154 73325 380918 73561
rect 381154 73325 387918 73561
rect 388154 73325 394918 73561
rect 395154 73325 401918 73561
rect 402154 73325 408918 73561
rect 409154 73325 415918 73561
rect 416154 73325 422918 73561
rect 423154 73325 429918 73561
rect 430154 73325 436918 73561
rect 437154 73325 443918 73561
rect 444154 73325 450918 73561
rect 451154 73325 457918 73561
rect 458154 73325 464918 73561
rect 465154 73325 471918 73561
rect 472154 73325 478918 73561
rect 479154 73325 485918 73561
rect 486154 73325 492918 73561
rect 493154 73325 499918 73561
rect 500154 73325 506918 73561
rect 507154 73325 513918 73561
rect 514154 73325 520918 73561
rect 521154 73325 527918 73561
rect 528154 73325 534918 73561
rect 535154 73325 541918 73561
rect 542154 73325 548918 73561
rect 549154 73325 555918 73561
rect 556154 73325 562918 73561
rect 563154 73325 569918 73561
rect 570154 73325 576918 73561
rect 577154 73325 587570 73561
rect 587806 73325 587890 73561
rect 588126 73325 588210 73561
rect 588446 73325 588530 73561
rect 588766 73325 588874 73561
rect -4950 73283 588874 73325
rect -4950 72494 588874 72536
rect -4950 72258 -3090 72494
rect -2854 72258 -2770 72494
rect -2534 72258 -2450 72494
rect -2214 72258 -2130 72494
rect -1894 72258 1186 72494
rect 1422 72258 8186 72494
rect 8422 72258 15186 72494
rect 15422 72258 22186 72494
rect 22422 72258 29186 72494
rect 29422 72258 36186 72494
rect 36422 72258 43186 72494
rect 43422 72258 50186 72494
rect 50422 72258 57186 72494
rect 57422 72258 64186 72494
rect 64422 72258 71186 72494
rect 71422 72258 78186 72494
rect 78422 72258 85186 72494
rect 85422 72258 92186 72494
rect 92422 72258 99186 72494
rect 99422 72258 106186 72494
rect 106422 72258 113186 72494
rect 113422 72258 120186 72494
rect 120422 72258 127186 72494
rect 127422 72258 134186 72494
rect 134422 72258 141186 72494
rect 141422 72258 148186 72494
rect 148422 72258 155186 72494
rect 155422 72258 162186 72494
rect 162422 72258 169186 72494
rect 169422 72258 176186 72494
rect 176422 72258 183186 72494
rect 183422 72258 190186 72494
rect 190422 72258 197186 72494
rect 197422 72258 204186 72494
rect 204422 72258 211186 72494
rect 211422 72258 218186 72494
rect 218422 72258 225186 72494
rect 225422 72258 232186 72494
rect 232422 72258 239186 72494
rect 239422 72258 246186 72494
rect 246422 72258 253186 72494
rect 253422 72258 260186 72494
rect 260422 72258 267186 72494
rect 267422 72258 274186 72494
rect 274422 72258 281186 72494
rect 281422 72258 288186 72494
rect 288422 72258 295186 72494
rect 295422 72258 302186 72494
rect 302422 72258 309186 72494
rect 309422 72258 316186 72494
rect 316422 72258 323186 72494
rect 323422 72258 330186 72494
rect 330422 72258 337186 72494
rect 337422 72258 344186 72494
rect 344422 72258 351186 72494
rect 351422 72258 358186 72494
rect 358422 72258 365186 72494
rect 365422 72258 372186 72494
rect 372422 72258 379186 72494
rect 379422 72258 386186 72494
rect 386422 72258 393186 72494
rect 393422 72258 400186 72494
rect 400422 72258 407186 72494
rect 407422 72258 414186 72494
rect 414422 72258 421186 72494
rect 421422 72258 428186 72494
rect 428422 72258 435186 72494
rect 435422 72258 442186 72494
rect 442422 72258 449186 72494
rect 449422 72258 456186 72494
rect 456422 72258 463186 72494
rect 463422 72258 470186 72494
rect 470422 72258 477186 72494
rect 477422 72258 484186 72494
rect 484422 72258 491186 72494
rect 491422 72258 498186 72494
rect 498422 72258 505186 72494
rect 505422 72258 512186 72494
rect 512422 72258 519186 72494
rect 519422 72258 526186 72494
rect 526422 72258 533186 72494
rect 533422 72258 540186 72494
rect 540422 72258 547186 72494
rect 547422 72258 554186 72494
rect 554422 72258 561186 72494
rect 561422 72258 568186 72494
rect 568422 72258 575186 72494
rect 575422 72258 582186 72494
rect 582422 72258 585818 72494
rect 586054 72258 586138 72494
rect 586374 72258 586458 72494
rect 586694 72258 586778 72494
rect 587014 72258 588874 72494
rect -4950 72216 588874 72258
rect -4950 66561 588874 66603
rect -4950 66325 -4842 66561
rect -4606 66325 -4522 66561
rect -4286 66325 -4202 66561
rect -3966 66325 -3882 66561
rect -3646 66325 2918 66561
rect 3154 66325 9918 66561
rect 10154 66325 16918 66561
rect 17154 66325 23918 66561
rect 24154 66325 30918 66561
rect 31154 66325 37918 66561
rect 38154 66325 44918 66561
rect 45154 66325 51918 66561
rect 52154 66325 58918 66561
rect 59154 66325 65918 66561
rect 66154 66325 72918 66561
rect 73154 66325 79918 66561
rect 80154 66325 86918 66561
rect 87154 66325 93918 66561
rect 94154 66325 100918 66561
rect 101154 66325 107918 66561
rect 108154 66325 114918 66561
rect 115154 66325 121918 66561
rect 122154 66325 128918 66561
rect 129154 66325 135918 66561
rect 136154 66325 142918 66561
rect 143154 66325 149918 66561
rect 150154 66325 156918 66561
rect 157154 66325 163918 66561
rect 164154 66325 170918 66561
rect 171154 66325 177918 66561
rect 178154 66325 184918 66561
rect 185154 66325 191918 66561
rect 192154 66325 198918 66561
rect 199154 66325 205918 66561
rect 206154 66325 212918 66561
rect 213154 66325 219918 66561
rect 220154 66325 226918 66561
rect 227154 66325 233918 66561
rect 234154 66325 240918 66561
rect 241154 66325 247918 66561
rect 248154 66325 254918 66561
rect 255154 66325 261918 66561
rect 262154 66325 268918 66561
rect 269154 66325 275918 66561
rect 276154 66325 282918 66561
rect 283154 66325 289918 66561
rect 290154 66325 296918 66561
rect 297154 66325 303918 66561
rect 304154 66325 310918 66561
rect 311154 66325 317918 66561
rect 318154 66325 324918 66561
rect 325154 66325 331918 66561
rect 332154 66325 338918 66561
rect 339154 66325 345918 66561
rect 346154 66325 352918 66561
rect 353154 66325 359918 66561
rect 360154 66325 366918 66561
rect 367154 66325 373918 66561
rect 374154 66325 380918 66561
rect 381154 66325 387918 66561
rect 388154 66325 394918 66561
rect 395154 66325 401918 66561
rect 402154 66325 408918 66561
rect 409154 66325 415918 66561
rect 416154 66325 422918 66561
rect 423154 66325 429918 66561
rect 430154 66325 436918 66561
rect 437154 66325 443918 66561
rect 444154 66325 450918 66561
rect 451154 66325 457918 66561
rect 458154 66325 464918 66561
rect 465154 66325 471918 66561
rect 472154 66325 478918 66561
rect 479154 66325 485918 66561
rect 486154 66325 492918 66561
rect 493154 66325 499918 66561
rect 500154 66325 506918 66561
rect 507154 66325 513918 66561
rect 514154 66325 520918 66561
rect 521154 66325 527918 66561
rect 528154 66325 534918 66561
rect 535154 66325 541918 66561
rect 542154 66325 548918 66561
rect 549154 66325 555918 66561
rect 556154 66325 562918 66561
rect 563154 66325 569918 66561
rect 570154 66325 576918 66561
rect 577154 66325 587570 66561
rect 587806 66325 587890 66561
rect 588126 66325 588210 66561
rect 588446 66325 588530 66561
rect 588766 66325 588874 66561
rect -4950 66283 588874 66325
rect -4950 65494 588874 65536
rect -4950 65258 -3090 65494
rect -2854 65258 -2770 65494
rect -2534 65258 -2450 65494
rect -2214 65258 -2130 65494
rect -1894 65258 1186 65494
rect 1422 65258 8186 65494
rect 8422 65258 15186 65494
rect 15422 65258 22186 65494
rect 22422 65258 29186 65494
rect 29422 65258 36186 65494
rect 36422 65258 43186 65494
rect 43422 65258 50186 65494
rect 50422 65258 57186 65494
rect 57422 65258 64186 65494
rect 64422 65258 71186 65494
rect 71422 65258 78186 65494
rect 78422 65258 85186 65494
rect 85422 65258 92186 65494
rect 92422 65258 99186 65494
rect 99422 65258 106186 65494
rect 106422 65258 113186 65494
rect 113422 65258 120186 65494
rect 120422 65258 127186 65494
rect 127422 65258 134186 65494
rect 134422 65258 141186 65494
rect 141422 65258 148186 65494
rect 148422 65258 155186 65494
rect 155422 65258 162186 65494
rect 162422 65258 169186 65494
rect 169422 65258 176186 65494
rect 176422 65258 183186 65494
rect 183422 65258 190186 65494
rect 190422 65258 197186 65494
rect 197422 65258 204186 65494
rect 204422 65258 211186 65494
rect 211422 65258 218186 65494
rect 218422 65258 225186 65494
rect 225422 65258 232186 65494
rect 232422 65258 239186 65494
rect 239422 65258 246186 65494
rect 246422 65258 253186 65494
rect 253422 65258 260186 65494
rect 260422 65258 267186 65494
rect 267422 65258 274186 65494
rect 274422 65258 281186 65494
rect 281422 65258 288186 65494
rect 288422 65258 295186 65494
rect 295422 65258 302186 65494
rect 302422 65258 309186 65494
rect 309422 65258 316186 65494
rect 316422 65258 323186 65494
rect 323422 65258 330186 65494
rect 330422 65258 337186 65494
rect 337422 65258 344186 65494
rect 344422 65258 351186 65494
rect 351422 65258 358186 65494
rect 358422 65258 365186 65494
rect 365422 65258 372186 65494
rect 372422 65258 379186 65494
rect 379422 65258 386186 65494
rect 386422 65258 393186 65494
rect 393422 65258 400186 65494
rect 400422 65258 407186 65494
rect 407422 65258 414186 65494
rect 414422 65258 421186 65494
rect 421422 65258 428186 65494
rect 428422 65258 435186 65494
rect 435422 65258 442186 65494
rect 442422 65258 449186 65494
rect 449422 65258 456186 65494
rect 456422 65258 463186 65494
rect 463422 65258 470186 65494
rect 470422 65258 477186 65494
rect 477422 65258 484186 65494
rect 484422 65258 491186 65494
rect 491422 65258 498186 65494
rect 498422 65258 505186 65494
rect 505422 65258 512186 65494
rect 512422 65258 519186 65494
rect 519422 65258 526186 65494
rect 526422 65258 533186 65494
rect 533422 65258 540186 65494
rect 540422 65258 547186 65494
rect 547422 65258 554186 65494
rect 554422 65258 561186 65494
rect 561422 65258 568186 65494
rect 568422 65258 575186 65494
rect 575422 65258 582186 65494
rect 582422 65258 585818 65494
rect 586054 65258 586138 65494
rect 586374 65258 586458 65494
rect 586694 65258 586778 65494
rect 587014 65258 588874 65494
rect -4950 65216 588874 65258
rect -4950 59561 588874 59603
rect -4950 59325 -4842 59561
rect -4606 59325 -4522 59561
rect -4286 59325 -4202 59561
rect -3966 59325 -3882 59561
rect -3646 59325 2918 59561
rect 3154 59325 9918 59561
rect 10154 59325 16918 59561
rect 17154 59325 23918 59561
rect 24154 59325 30918 59561
rect 31154 59325 37918 59561
rect 38154 59325 44918 59561
rect 45154 59325 51918 59561
rect 52154 59325 58918 59561
rect 59154 59325 65918 59561
rect 66154 59325 72918 59561
rect 73154 59325 79918 59561
rect 80154 59325 86918 59561
rect 87154 59325 93918 59561
rect 94154 59325 100918 59561
rect 101154 59325 107918 59561
rect 108154 59325 114918 59561
rect 115154 59325 121918 59561
rect 122154 59325 128918 59561
rect 129154 59325 135918 59561
rect 136154 59325 142918 59561
rect 143154 59325 149918 59561
rect 150154 59325 156918 59561
rect 157154 59325 163918 59561
rect 164154 59325 170918 59561
rect 171154 59325 177918 59561
rect 178154 59325 184918 59561
rect 185154 59325 191918 59561
rect 192154 59325 198918 59561
rect 199154 59325 205918 59561
rect 206154 59325 212918 59561
rect 213154 59325 219918 59561
rect 220154 59325 226918 59561
rect 227154 59325 233918 59561
rect 234154 59325 240918 59561
rect 241154 59325 247918 59561
rect 248154 59325 254918 59561
rect 255154 59325 261918 59561
rect 262154 59325 268918 59561
rect 269154 59325 275918 59561
rect 276154 59325 282918 59561
rect 283154 59325 289918 59561
rect 290154 59325 296918 59561
rect 297154 59325 303918 59561
rect 304154 59325 310918 59561
rect 311154 59325 317918 59561
rect 318154 59325 324918 59561
rect 325154 59325 331918 59561
rect 332154 59325 338918 59561
rect 339154 59325 345918 59561
rect 346154 59325 352918 59561
rect 353154 59325 359918 59561
rect 360154 59325 366918 59561
rect 367154 59325 373918 59561
rect 374154 59325 380918 59561
rect 381154 59325 387918 59561
rect 388154 59325 394918 59561
rect 395154 59325 401918 59561
rect 402154 59325 408918 59561
rect 409154 59325 415918 59561
rect 416154 59325 422918 59561
rect 423154 59325 429918 59561
rect 430154 59325 436918 59561
rect 437154 59325 443918 59561
rect 444154 59325 450918 59561
rect 451154 59325 457918 59561
rect 458154 59325 464918 59561
rect 465154 59325 471918 59561
rect 472154 59325 478918 59561
rect 479154 59325 485918 59561
rect 486154 59325 492918 59561
rect 493154 59325 499918 59561
rect 500154 59325 506918 59561
rect 507154 59325 513918 59561
rect 514154 59325 520918 59561
rect 521154 59325 527918 59561
rect 528154 59325 534918 59561
rect 535154 59325 541918 59561
rect 542154 59325 548918 59561
rect 549154 59325 555918 59561
rect 556154 59325 562918 59561
rect 563154 59325 569918 59561
rect 570154 59325 576918 59561
rect 577154 59325 587570 59561
rect 587806 59325 587890 59561
rect 588126 59325 588210 59561
rect 588446 59325 588530 59561
rect 588766 59325 588874 59561
rect -4950 59283 588874 59325
rect -4950 58494 588874 58536
rect -4950 58258 -3090 58494
rect -2854 58258 -2770 58494
rect -2534 58258 -2450 58494
rect -2214 58258 -2130 58494
rect -1894 58258 1186 58494
rect 1422 58258 8186 58494
rect 8422 58258 15186 58494
rect 15422 58258 22186 58494
rect 22422 58258 29186 58494
rect 29422 58258 36186 58494
rect 36422 58258 43186 58494
rect 43422 58258 50186 58494
rect 50422 58258 57186 58494
rect 57422 58258 64186 58494
rect 64422 58258 71186 58494
rect 71422 58258 78186 58494
rect 78422 58258 85186 58494
rect 85422 58258 92186 58494
rect 92422 58258 99186 58494
rect 99422 58258 106186 58494
rect 106422 58258 113186 58494
rect 113422 58258 120186 58494
rect 120422 58258 127186 58494
rect 127422 58258 134186 58494
rect 134422 58258 141186 58494
rect 141422 58258 148186 58494
rect 148422 58258 155186 58494
rect 155422 58258 162186 58494
rect 162422 58258 169186 58494
rect 169422 58258 176186 58494
rect 176422 58258 183186 58494
rect 183422 58258 190186 58494
rect 190422 58258 197186 58494
rect 197422 58258 204186 58494
rect 204422 58258 211186 58494
rect 211422 58258 218186 58494
rect 218422 58258 225186 58494
rect 225422 58258 232186 58494
rect 232422 58258 239186 58494
rect 239422 58258 246186 58494
rect 246422 58258 253186 58494
rect 253422 58258 260186 58494
rect 260422 58258 267186 58494
rect 267422 58258 274186 58494
rect 274422 58258 281186 58494
rect 281422 58258 288186 58494
rect 288422 58258 295186 58494
rect 295422 58258 302186 58494
rect 302422 58258 309186 58494
rect 309422 58258 316186 58494
rect 316422 58258 323186 58494
rect 323422 58258 330186 58494
rect 330422 58258 337186 58494
rect 337422 58258 344186 58494
rect 344422 58258 351186 58494
rect 351422 58258 358186 58494
rect 358422 58258 365186 58494
rect 365422 58258 372186 58494
rect 372422 58258 379186 58494
rect 379422 58258 386186 58494
rect 386422 58258 393186 58494
rect 393422 58258 400186 58494
rect 400422 58258 407186 58494
rect 407422 58258 414186 58494
rect 414422 58258 421186 58494
rect 421422 58258 428186 58494
rect 428422 58258 435186 58494
rect 435422 58258 442186 58494
rect 442422 58258 449186 58494
rect 449422 58258 456186 58494
rect 456422 58258 463186 58494
rect 463422 58258 470186 58494
rect 470422 58258 477186 58494
rect 477422 58258 484186 58494
rect 484422 58258 491186 58494
rect 491422 58258 498186 58494
rect 498422 58258 505186 58494
rect 505422 58258 512186 58494
rect 512422 58258 519186 58494
rect 519422 58258 526186 58494
rect 526422 58258 533186 58494
rect 533422 58258 540186 58494
rect 540422 58258 547186 58494
rect 547422 58258 554186 58494
rect 554422 58258 561186 58494
rect 561422 58258 568186 58494
rect 568422 58258 575186 58494
rect 575422 58258 582186 58494
rect 582422 58258 585818 58494
rect 586054 58258 586138 58494
rect 586374 58258 586458 58494
rect 586694 58258 586778 58494
rect 587014 58258 588874 58494
rect -4950 58216 588874 58258
rect -4950 52561 588874 52603
rect -4950 52325 -4842 52561
rect -4606 52325 -4522 52561
rect -4286 52325 -4202 52561
rect -3966 52325 -3882 52561
rect -3646 52325 2918 52561
rect 3154 52325 9918 52561
rect 10154 52325 16918 52561
rect 17154 52325 23918 52561
rect 24154 52325 30918 52561
rect 31154 52325 37918 52561
rect 38154 52325 44918 52561
rect 45154 52325 51918 52561
rect 52154 52325 58918 52561
rect 59154 52325 65918 52561
rect 66154 52325 72918 52561
rect 73154 52325 79918 52561
rect 80154 52325 86918 52561
rect 87154 52325 93918 52561
rect 94154 52325 100918 52561
rect 101154 52325 107918 52561
rect 108154 52325 114918 52561
rect 115154 52325 121918 52561
rect 122154 52325 128918 52561
rect 129154 52325 135918 52561
rect 136154 52325 142918 52561
rect 143154 52325 149918 52561
rect 150154 52325 156918 52561
rect 157154 52325 163918 52561
rect 164154 52325 170918 52561
rect 171154 52325 177918 52561
rect 178154 52325 184918 52561
rect 185154 52325 191918 52561
rect 192154 52325 198918 52561
rect 199154 52325 205918 52561
rect 206154 52325 212918 52561
rect 213154 52325 219918 52561
rect 220154 52325 226918 52561
rect 227154 52325 233918 52561
rect 234154 52325 240918 52561
rect 241154 52325 247918 52561
rect 248154 52325 254918 52561
rect 255154 52325 261918 52561
rect 262154 52325 268918 52561
rect 269154 52325 275918 52561
rect 276154 52325 282918 52561
rect 283154 52325 289918 52561
rect 290154 52325 296918 52561
rect 297154 52325 303918 52561
rect 304154 52325 310918 52561
rect 311154 52325 317918 52561
rect 318154 52325 324918 52561
rect 325154 52325 331918 52561
rect 332154 52325 338918 52561
rect 339154 52325 345918 52561
rect 346154 52325 352918 52561
rect 353154 52325 359918 52561
rect 360154 52325 366918 52561
rect 367154 52325 373918 52561
rect 374154 52325 380918 52561
rect 381154 52325 387918 52561
rect 388154 52325 394918 52561
rect 395154 52325 401918 52561
rect 402154 52325 408918 52561
rect 409154 52325 415918 52561
rect 416154 52325 422918 52561
rect 423154 52325 429918 52561
rect 430154 52325 436918 52561
rect 437154 52325 443918 52561
rect 444154 52325 450918 52561
rect 451154 52325 457918 52561
rect 458154 52325 464918 52561
rect 465154 52325 471918 52561
rect 472154 52325 478918 52561
rect 479154 52325 485918 52561
rect 486154 52325 492918 52561
rect 493154 52325 499918 52561
rect 500154 52325 506918 52561
rect 507154 52325 513918 52561
rect 514154 52325 520918 52561
rect 521154 52325 527918 52561
rect 528154 52325 534918 52561
rect 535154 52325 541918 52561
rect 542154 52325 548918 52561
rect 549154 52325 555918 52561
rect 556154 52325 562918 52561
rect 563154 52325 569918 52561
rect 570154 52325 576918 52561
rect 577154 52325 587570 52561
rect 587806 52325 587890 52561
rect 588126 52325 588210 52561
rect 588446 52325 588530 52561
rect 588766 52325 588874 52561
rect -4950 52283 588874 52325
rect -4950 51494 588874 51536
rect -4950 51258 -3090 51494
rect -2854 51258 -2770 51494
rect -2534 51258 -2450 51494
rect -2214 51258 -2130 51494
rect -1894 51258 1186 51494
rect 1422 51258 8186 51494
rect 8422 51258 15186 51494
rect 15422 51258 22186 51494
rect 22422 51258 29186 51494
rect 29422 51258 36186 51494
rect 36422 51258 43186 51494
rect 43422 51258 50186 51494
rect 50422 51258 57186 51494
rect 57422 51258 64186 51494
rect 64422 51258 71186 51494
rect 71422 51258 78186 51494
rect 78422 51258 85186 51494
rect 85422 51258 92186 51494
rect 92422 51258 99186 51494
rect 99422 51258 106186 51494
rect 106422 51258 113186 51494
rect 113422 51258 120186 51494
rect 120422 51258 127186 51494
rect 127422 51258 134186 51494
rect 134422 51258 141186 51494
rect 141422 51258 148186 51494
rect 148422 51258 155186 51494
rect 155422 51258 162186 51494
rect 162422 51258 169186 51494
rect 169422 51258 176186 51494
rect 176422 51258 183186 51494
rect 183422 51258 190186 51494
rect 190422 51258 197186 51494
rect 197422 51258 204186 51494
rect 204422 51258 211186 51494
rect 211422 51258 218186 51494
rect 218422 51258 225186 51494
rect 225422 51258 232186 51494
rect 232422 51258 239186 51494
rect 239422 51258 246186 51494
rect 246422 51258 253186 51494
rect 253422 51258 260186 51494
rect 260422 51258 267186 51494
rect 267422 51258 274186 51494
rect 274422 51258 281186 51494
rect 281422 51258 288186 51494
rect 288422 51258 295186 51494
rect 295422 51258 302186 51494
rect 302422 51258 309186 51494
rect 309422 51258 316186 51494
rect 316422 51258 323186 51494
rect 323422 51258 330186 51494
rect 330422 51258 337186 51494
rect 337422 51258 344186 51494
rect 344422 51258 351186 51494
rect 351422 51258 358186 51494
rect 358422 51258 365186 51494
rect 365422 51258 372186 51494
rect 372422 51258 379186 51494
rect 379422 51258 386186 51494
rect 386422 51258 393186 51494
rect 393422 51258 400186 51494
rect 400422 51258 407186 51494
rect 407422 51258 414186 51494
rect 414422 51258 421186 51494
rect 421422 51258 428186 51494
rect 428422 51258 435186 51494
rect 435422 51258 442186 51494
rect 442422 51258 449186 51494
rect 449422 51258 456186 51494
rect 456422 51258 463186 51494
rect 463422 51258 470186 51494
rect 470422 51258 477186 51494
rect 477422 51258 484186 51494
rect 484422 51258 491186 51494
rect 491422 51258 498186 51494
rect 498422 51258 505186 51494
rect 505422 51258 512186 51494
rect 512422 51258 519186 51494
rect 519422 51258 526186 51494
rect 526422 51258 533186 51494
rect 533422 51258 540186 51494
rect 540422 51258 547186 51494
rect 547422 51258 554186 51494
rect 554422 51258 561186 51494
rect 561422 51258 568186 51494
rect 568422 51258 575186 51494
rect 575422 51258 582186 51494
rect 582422 51258 585818 51494
rect 586054 51258 586138 51494
rect 586374 51258 586458 51494
rect 586694 51258 586778 51494
rect 587014 51258 588874 51494
rect -4950 51216 588874 51258
rect -4950 45561 588874 45603
rect -4950 45325 -4842 45561
rect -4606 45325 -4522 45561
rect -4286 45325 -4202 45561
rect -3966 45325 -3882 45561
rect -3646 45325 2918 45561
rect 3154 45325 9918 45561
rect 10154 45325 16918 45561
rect 17154 45325 23918 45561
rect 24154 45325 30918 45561
rect 31154 45325 37918 45561
rect 38154 45325 44918 45561
rect 45154 45325 51918 45561
rect 52154 45325 58918 45561
rect 59154 45325 65918 45561
rect 66154 45325 72918 45561
rect 73154 45325 79918 45561
rect 80154 45325 86918 45561
rect 87154 45325 93918 45561
rect 94154 45325 100918 45561
rect 101154 45325 107918 45561
rect 108154 45325 114918 45561
rect 115154 45325 121918 45561
rect 122154 45325 128918 45561
rect 129154 45325 135918 45561
rect 136154 45325 142918 45561
rect 143154 45325 149918 45561
rect 150154 45325 156918 45561
rect 157154 45325 163918 45561
rect 164154 45325 170918 45561
rect 171154 45325 177918 45561
rect 178154 45325 184918 45561
rect 185154 45325 191918 45561
rect 192154 45325 198918 45561
rect 199154 45325 205918 45561
rect 206154 45325 212918 45561
rect 213154 45325 219918 45561
rect 220154 45325 226918 45561
rect 227154 45325 233918 45561
rect 234154 45325 240918 45561
rect 241154 45325 247918 45561
rect 248154 45325 254918 45561
rect 255154 45325 261918 45561
rect 262154 45325 268918 45561
rect 269154 45325 275918 45561
rect 276154 45325 282918 45561
rect 283154 45325 289918 45561
rect 290154 45325 296918 45561
rect 297154 45325 303918 45561
rect 304154 45325 310918 45561
rect 311154 45325 317918 45561
rect 318154 45325 324918 45561
rect 325154 45325 331918 45561
rect 332154 45325 338918 45561
rect 339154 45325 345918 45561
rect 346154 45325 352918 45561
rect 353154 45325 359918 45561
rect 360154 45325 366918 45561
rect 367154 45325 373918 45561
rect 374154 45325 380918 45561
rect 381154 45325 387918 45561
rect 388154 45325 394918 45561
rect 395154 45325 401918 45561
rect 402154 45325 408918 45561
rect 409154 45325 415918 45561
rect 416154 45325 422918 45561
rect 423154 45325 429918 45561
rect 430154 45325 436918 45561
rect 437154 45325 443918 45561
rect 444154 45325 450918 45561
rect 451154 45325 457918 45561
rect 458154 45325 464918 45561
rect 465154 45325 471918 45561
rect 472154 45325 478918 45561
rect 479154 45325 485918 45561
rect 486154 45325 492918 45561
rect 493154 45325 499918 45561
rect 500154 45325 506918 45561
rect 507154 45325 513918 45561
rect 514154 45325 520918 45561
rect 521154 45325 527918 45561
rect 528154 45325 534918 45561
rect 535154 45325 541918 45561
rect 542154 45325 548918 45561
rect 549154 45325 555918 45561
rect 556154 45325 562918 45561
rect 563154 45325 569918 45561
rect 570154 45325 576918 45561
rect 577154 45325 587570 45561
rect 587806 45325 587890 45561
rect 588126 45325 588210 45561
rect 588446 45325 588530 45561
rect 588766 45325 588874 45561
rect -4950 45283 588874 45325
rect -4950 44494 588874 44536
rect -4950 44258 -3090 44494
rect -2854 44258 -2770 44494
rect -2534 44258 -2450 44494
rect -2214 44258 -2130 44494
rect -1894 44258 1186 44494
rect 1422 44258 8186 44494
rect 8422 44258 15186 44494
rect 15422 44258 22186 44494
rect 22422 44258 29186 44494
rect 29422 44258 36186 44494
rect 36422 44258 43186 44494
rect 43422 44258 50186 44494
rect 50422 44258 57186 44494
rect 57422 44258 64186 44494
rect 64422 44258 71186 44494
rect 71422 44258 78186 44494
rect 78422 44258 85186 44494
rect 85422 44258 92186 44494
rect 92422 44258 99186 44494
rect 99422 44258 106186 44494
rect 106422 44258 113186 44494
rect 113422 44258 120186 44494
rect 120422 44258 127186 44494
rect 127422 44258 134186 44494
rect 134422 44258 141186 44494
rect 141422 44258 148186 44494
rect 148422 44258 155186 44494
rect 155422 44258 162186 44494
rect 162422 44258 169186 44494
rect 169422 44258 176186 44494
rect 176422 44258 183186 44494
rect 183422 44258 190186 44494
rect 190422 44258 197186 44494
rect 197422 44258 204186 44494
rect 204422 44258 211186 44494
rect 211422 44258 218186 44494
rect 218422 44258 225186 44494
rect 225422 44258 232186 44494
rect 232422 44258 239186 44494
rect 239422 44258 246186 44494
rect 246422 44258 253186 44494
rect 253422 44258 260186 44494
rect 260422 44258 267186 44494
rect 267422 44258 274186 44494
rect 274422 44258 281186 44494
rect 281422 44258 288186 44494
rect 288422 44258 295186 44494
rect 295422 44258 302186 44494
rect 302422 44258 309186 44494
rect 309422 44258 316186 44494
rect 316422 44258 323186 44494
rect 323422 44258 330186 44494
rect 330422 44258 337186 44494
rect 337422 44258 344186 44494
rect 344422 44258 351186 44494
rect 351422 44258 358186 44494
rect 358422 44258 365186 44494
rect 365422 44258 372186 44494
rect 372422 44258 379186 44494
rect 379422 44258 386186 44494
rect 386422 44258 393186 44494
rect 393422 44258 400186 44494
rect 400422 44258 407186 44494
rect 407422 44258 414186 44494
rect 414422 44258 421186 44494
rect 421422 44258 428186 44494
rect 428422 44258 435186 44494
rect 435422 44258 442186 44494
rect 442422 44258 449186 44494
rect 449422 44258 456186 44494
rect 456422 44258 463186 44494
rect 463422 44258 470186 44494
rect 470422 44258 477186 44494
rect 477422 44258 484186 44494
rect 484422 44258 491186 44494
rect 491422 44258 498186 44494
rect 498422 44258 505186 44494
rect 505422 44258 512186 44494
rect 512422 44258 519186 44494
rect 519422 44258 526186 44494
rect 526422 44258 533186 44494
rect 533422 44258 540186 44494
rect 540422 44258 547186 44494
rect 547422 44258 554186 44494
rect 554422 44258 561186 44494
rect 561422 44258 568186 44494
rect 568422 44258 575186 44494
rect 575422 44258 582186 44494
rect 582422 44258 585818 44494
rect 586054 44258 586138 44494
rect 586374 44258 586458 44494
rect 586694 44258 586778 44494
rect 587014 44258 588874 44494
rect -4950 44216 588874 44258
rect -4950 38561 588874 38603
rect -4950 38325 -4842 38561
rect -4606 38325 -4522 38561
rect -4286 38325 -4202 38561
rect -3966 38325 -3882 38561
rect -3646 38325 2918 38561
rect 3154 38325 9918 38561
rect 10154 38325 16918 38561
rect 17154 38325 23918 38561
rect 24154 38325 30918 38561
rect 31154 38325 37918 38561
rect 38154 38325 44918 38561
rect 45154 38325 51918 38561
rect 52154 38325 58918 38561
rect 59154 38325 65918 38561
rect 66154 38325 72918 38561
rect 73154 38325 79918 38561
rect 80154 38325 86918 38561
rect 87154 38325 93918 38561
rect 94154 38325 100918 38561
rect 101154 38325 107918 38561
rect 108154 38325 114918 38561
rect 115154 38325 121918 38561
rect 122154 38325 128918 38561
rect 129154 38325 135918 38561
rect 136154 38325 142918 38561
rect 143154 38325 149918 38561
rect 150154 38325 156918 38561
rect 157154 38325 163918 38561
rect 164154 38325 170918 38561
rect 171154 38325 177918 38561
rect 178154 38325 184918 38561
rect 185154 38325 191918 38561
rect 192154 38325 198918 38561
rect 199154 38325 205918 38561
rect 206154 38325 212918 38561
rect 213154 38325 219918 38561
rect 220154 38325 226918 38561
rect 227154 38325 233918 38561
rect 234154 38325 240918 38561
rect 241154 38325 247918 38561
rect 248154 38325 254918 38561
rect 255154 38325 261918 38561
rect 262154 38325 268918 38561
rect 269154 38325 275918 38561
rect 276154 38325 282918 38561
rect 283154 38325 289918 38561
rect 290154 38325 296918 38561
rect 297154 38325 303918 38561
rect 304154 38325 310918 38561
rect 311154 38325 317918 38561
rect 318154 38325 324918 38561
rect 325154 38325 331918 38561
rect 332154 38325 338918 38561
rect 339154 38325 345918 38561
rect 346154 38325 352918 38561
rect 353154 38325 359918 38561
rect 360154 38325 366918 38561
rect 367154 38325 373918 38561
rect 374154 38325 380918 38561
rect 381154 38325 387918 38561
rect 388154 38325 394918 38561
rect 395154 38325 401918 38561
rect 402154 38325 408918 38561
rect 409154 38325 415918 38561
rect 416154 38325 422918 38561
rect 423154 38325 429918 38561
rect 430154 38325 436918 38561
rect 437154 38325 443918 38561
rect 444154 38325 450918 38561
rect 451154 38325 457918 38561
rect 458154 38325 464918 38561
rect 465154 38325 471918 38561
rect 472154 38325 478918 38561
rect 479154 38325 485918 38561
rect 486154 38325 492918 38561
rect 493154 38325 499918 38561
rect 500154 38325 506918 38561
rect 507154 38325 513918 38561
rect 514154 38325 520918 38561
rect 521154 38325 527918 38561
rect 528154 38325 534918 38561
rect 535154 38325 541918 38561
rect 542154 38325 548918 38561
rect 549154 38325 555918 38561
rect 556154 38325 562918 38561
rect 563154 38325 569918 38561
rect 570154 38325 576918 38561
rect 577154 38325 587570 38561
rect 587806 38325 587890 38561
rect 588126 38325 588210 38561
rect 588446 38325 588530 38561
rect 588766 38325 588874 38561
rect -4950 38283 588874 38325
rect -4950 37494 588874 37536
rect -4950 37258 -3090 37494
rect -2854 37258 -2770 37494
rect -2534 37258 -2450 37494
rect -2214 37258 -2130 37494
rect -1894 37258 1186 37494
rect 1422 37258 8186 37494
rect 8422 37258 15186 37494
rect 15422 37258 22186 37494
rect 22422 37258 29186 37494
rect 29422 37258 36186 37494
rect 36422 37258 43186 37494
rect 43422 37258 50186 37494
rect 50422 37258 57186 37494
rect 57422 37258 64186 37494
rect 64422 37258 71186 37494
rect 71422 37258 78186 37494
rect 78422 37258 85186 37494
rect 85422 37258 92186 37494
rect 92422 37258 99186 37494
rect 99422 37258 106186 37494
rect 106422 37258 113186 37494
rect 113422 37258 120186 37494
rect 120422 37258 127186 37494
rect 127422 37258 134186 37494
rect 134422 37258 141186 37494
rect 141422 37258 148186 37494
rect 148422 37258 155186 37494
rect 155422 37258 162186 37494
rect 162422 37258 169186 37494
rect 169422 37258 176186 37494
rect 176422 37258 183186 37494
rect 183422 37258 190186 37494
rect 190422 37258 197186 37494
rect 197422 37258 204186 37494
rect 204422 37258 211186 37494
rect 211422 37258 218186 37494
rect 218422 37258 225186 37494
rect 225422 37258 232186 37494
rect 232422 37258 239186 37494
rect 239422 37258 246186 37494
rect 246422 37258 253186 37494
rect 253422 37258 260186 37494
rect 260422 37258 267186 37494
rect 267422 37258 274186 37494
rect 274422 37258 281186 37494
rect 281422 37258 288186 37494
rect 288422 37258 295186 37494
rect 295422 37258 302186 37494
rect 302422 37258 309186 37494
rect 309422 37258 316186 37494
rect 316422 37258 323186 37494
rect 323422 37258 330186 37494
rect 330422 37258 337186 37494
rect 337422 37258 344186 37494
rect 344422 37258 351186 37494
rect 351422 37258 358186 37494
rect 358422 37258 365186 37494
rect 365422 37258 372186 37494
rect 372422 37258 379186 37494
rect 379422 37258 386186 37494
rect 386422 37258 393186 37494
rect 393422 37258 400186 37494
rect 400422 37258 407186 37494
rect 407422 37258 414186 37494
rect 414422 37258 421186 37494
rect 421422 37258 428186 37494
rect 428422 37258 435186 37494
rect 435422 37258 442186 37494
rect 442422 37258 449186 37494
rect 449422 37258 456186 37494
rect 456422 37258 463186 37494
rect 463422 37258 470186 37494
rect 470422 37258 477186 37494
rect 477422 37258 484186 37494
rect 484422 37258 491186 37494
rect 491422 37258 498186 37494
rect 498422 37258 505186 37494
rect 505422 37258 512186 37494
rect 512422 37258 519186 37494
rect 519422 37258 526186 37494
rect 526422 37258 533186 37494
rect 533422 37258 540186 37494
rect 540422 37258 547186 37494
rect 547422 37258 554186 37494
rect 554422 37258 561186 37494
rect 561422 37258 568186 37494
rect 568422 37258 575186 37494
rect 575422 37258 582186 37494
rect 582422 37258 585818 37494
rect 586054 37258 586138 37494
rect 586374 37258 586458 37494
rect 586694 37258 586778 37494
rect 587014 37258 588874 37494
rect -4950 37216 588874 37258
rect -4950 31561 588874 31603
rect -4950 31325 -4842 31561
rect -4606 31325 -4522 31561
rect -4286 31325 -4202 31561
rect -3966 31325 -3882 31561
rect -3646 31325 2918 31561
rect 3154 31325 9918 31561
rect 10154 31325 16918 31561
rect 17154 31325 23918 31561
rect 24154 31325 30918 31561
rect 31154 31325 37918 31561
rect 38154 31325 44918 31561
rect 45154 31325 51918 31561
rect 52154 31325 58918 31561
rect 59154 31325 65918 31561
rect 66154 31325 72918 31561
rect 73154 31325 79918 31561
rect 80154 31325 86918 31561
rect 87154 31325 93918 31561
rect 94154 31325 100918 31561
rect 101154 31325 107918 31561
rect 108154 31325 114918 31561
rect 115154 31325 121918 31561
rect 122154 31325 128918 31561
rect 129154 31325 135918 31561
rect 136154 31325 142918 31561
rect 143154 31325 149918 31561
rect 150154 31325 156918 31561
rect 157154 31325 163918 31561
rect 164154 31325 170918 31561
rect 171154 31325 177918 31561
rect 178154 31325 184918 31561
rect 185154 31325 191918 31561
rect 192154 31325 198918 31561
rect 199154 31325 205918 31561
rect 206154 31325 212918 31561
rect 213154 31325 219918 31561
rect 220154 31325 226918 31561
rect 227154 31325 233918 31561
rect 234154 31325 240918 31561
rect 241154 31325 247918 31561
rect 248154 31325 254918 31561
rect 255154 31325 261918 31561
rect 262154 31325 268918 31561
rect 269154 31325 275918 31561
rect 276154 31325 282918 31561
rect 283154 31325 289918 31561
rect 290154 31325 296918 31561
rect 297154 31325 303918 31561
rect 304154 31325 310918 31561
rect 311154 31325 317918 31561
rect 318154 31325 324918 31561
rect 325154 31325 331918 31561
rect 332154 31325 338918 31561
rect 339154 31325 345918 31561
rect 346154 31325 352918 31561
rect 353154 31325 359918 31561
rect 360154 31325 366918 31561
rect 367154 31325 373918 31561
rect 374154 31325 380918 31561
rect 381154 31325 387918 31561
rect 388154 31325 394918 31561
rect 395154 31325 401918 31561
rect 402154 31325 408918 31561
rect 409154 31325 415918 31561
rect 416154 31325 422918 31561
rect 423154 31325 429918 31561
rect 430154 31325 436918 31561
rect 437154 31325 443918 31561
rect 444154 31325 450918 31561
rect 451154 31325 457918 31561
rect 458154 31325 464918 31561
rect 465154 31325 471918 31561
rect 472154 31325 478918 31561
rect 479154 31325 485918 31561
rect 486154 31325 492918 31561
rect 493154 31325 499918 31561
rect 500154 31325 506918 31561
rect 507154 31325 513918 31561
rect 514154 31325 520918 31561
rect 521154 31325 527918 31561
rect 528154 31325 534918 31561
rect 535154 31325 541918 31561
rect 542154 31325 548918 31561
rect 549154 31325 555918 31561
rect 556154 31325 562918 31561
rect 563154 31325 569918 31561
rect 570154 31325 576918 31561
rect 577154 31325 587570 31561
rect 587806 31325 587890 31561
rect 588126 31325 588210 31561
rect 588446 31325 588530 31561
rect 588766 31325 588874 31561
rect -4950 31283 588874 31325
rect -4950 30494 588874 30536
rect -4950 30258 -3090 30494
rect -2854 30258 -2770 30494
rect -2534 30258 -2450 30494
rect -2214 30258 -2130 30494
rect -1894 30258 1186 30494
rect 1422 30258 8186 30494
rect 8422 30258 15186 30494
rect 15422 30258 22186 30494
rect 22422 30258 29186 30494
rect 29422 30258 36186 30494
rect 36422 30258 43186 30494
rect 43422 30258 50186 30494
rect 50422 30258 57186 30494
rect 57422 30258 64186 30494
rect 64422 30258 71186 30494
rect 71422 30258 78186 30494
rect 78422 30258 85186 30494
rect 85422 30258 92186 30494
rect 92422 30258 99186 30494
rect 99422 30258 106186 30494
rect 106422 30258 113186 30494
rect 113422 30258 120186 30494
rect 120422 30258 127186 30494
rect 127422 30258 134186 30494
rect 134422 30258 141186 30494
rect 141422 30258 148186 30494
rect 148422 30258 155186 30494
rect 155422 30258 162186 30494
rect 162422 30258 169186 30494
rect 169422 30258 176186 30494
rect 176422 30258 183186 30494
rect 183422 30258 190186 30494
rect 190422 30258 197186 30494
rect 197422 30258 204186 30494
rect 204422 30258 211186 30494
rect 211422 30258 218186 30494
rect 218422 30258 225186 30494
rect 225422 30258 232186 30494
rect 232422 30258 239186 30494
rect 239422 30258 246186 30494
rect 246422 30258 253186 30494
rect 253422 30258 260186 30494
rect 260422 30258 267186 30494
rect 267422 30258 274186 30494
rect 274422 30258 281186 30494
rect 281422 30258 288186 30494
rect 288422 30258 295186 30494
rect 295422 30258 302186 30494
rect 302422 30258 309186 30494
rect 309422 30258 316186 30494
rect 316422 30258 323186 30494
rect 323422 30258 330186 30494
rect 330422 30258 337186 30494
rect 337422 30258 344186 30494
rect 344422 30258 351186 30494
rect 351422 30258 358186 30494
rect 358422 30258 365186 30494
rect 365422 30258 372186 30494
rect 372422 30258 379186 30494
rect 379422 30258 386186 30494
rect 386422 30258 393186 30494
rect 393422 30258 400186 30494
rect 400422 30258 407186 30494
rect 407422 30258 414186 30494
rect 414422 30258 421186 30494
rect 421422 30258 428186 30494
rect 428422 30258 435186 30494
rect 435422 30258 442186 30494
rect 442422 30258 449186 30494
rect 449422 30258 456186 30494
rect 456422 30258 463186 30494
rect 463422 30258 470186 30494
rect 470422 30258 477186 30494
rect 477422 30258 484186 30494
rect 484422 30258 491186 30494
rect 491422 30258 498186 30494
rect 498422 30258 505186 30494
rect 505422 30258 512186 30494
rect 512422 30258 519186 30494
rect 519422 30258 526186 30494
rect 526422 30258 533186 30494
rect 533422 30258 540186 30494
rect 540422 30258 547186 30494
rect 547422 30258 554186 30494
rect 554422 30258 561186 30494
rect 561422 30258 568186 30494
rect 568422 30258 575186 30494
rect 575422 30258 582186 30494
rect 582422 30258 585818 30494
rect 586054 30258 586138 30494
rect 586374 30258 586458 30494
rect 586694 30258 586778 30494
rect 587014 30258 588874 30494
rect -4950 30216 588874 30258
rect -4950 24561 588874 24603
rect -4950 24325 -4842 24561
rect -4606 24325 -4522 24561
rect -4286 24325 -4202 24561
rect -3966 24325 -3882 24561
rect -3646 24325 2918 24561
rect 3154 24325 9918 24561
rect 10154 24325 16918 24561
rect 17154 24325 23918 24561
rect 24154 24325 30918 24561
rect 31154 24325 37918 24561
rect 38154 24325 44918 24561
rect 45154 24325 51918 24561
rect 52154 24325 58918 24561
rect 59154 24325 65918 24561
rect 66154 24325 72918 24561
rect 73154 24325 79918 24561
rect 80154 24325 86918 24561
rect 87154 24325 93918 24561
rect 94154 24325 100918 24561
rect 101154 24325 107918 24561
rect 108154 24325 114918 24561
rect 115154 24325 121918 24561
rect 122154 24325 128918 24561
rect 129154 24325 135918 24561
rect 136154 24325 142918 24561
rect 143154 24325 149918 24561
rect 150154 24325 156918 24561
rect 157154 24325 163918 24561
rect 164154 24325 170918 24561
rect 171154 24325 177918 24561
rect 178154 24325 184918 24561
rect 185154 24325 191918 24561
rect 192154 24325 198918 24561
rect 199154 24325 205918 24561
rect 206154 24325 212918 24561
rect 213154 24325 219918 24561
rect 220154 24325 226918 24561
rect 227154 24325 233918 24561
rect 234154 24325 240918 24561
rect 241154 24325 247918 24561
rect 248154 24325 254918 24561
rect 255154 24325 261918 24561
rect 262154 24325 268918 24561
rect 269154 24325 275918 24561
rect 276154 24325 282918 24561
rect 283154 24325 289918 24561
rect 290154 24325 296918 24561
rect 297154 24325 303918 24561
rect 304154 24325 310918 24561
rect 311154 24325 317918 24561
rect 318154 24325 324918 24561
rect 325154 24325 331918 24561
rect 332154 24325 338918 24561
rect 339154 24325 345918 24561
rect 346154 24325 352918 24561
rect 353154 24325 359918 24561
rect 360154 24325 366918 24561
rect 367154 24325 373918 24561
rect 374154 24325 380918 24561
rect 381154 24325 387918 24561
rect 388154 24325 394918 24561
rect 395154 24325 401918 24561
rect 402154 24325 408918 24561
rect 409154 24325 415918 24561
rect 416154 24325 422918 24561
rect 423154 24325 429918 24561
rect 430154 24325 436918 24561
rect 437154 24325 443918 24561
rect 444154 24325 450918 24561
rect 451154 24325 457918 24561
rect 458154 24325 464918 24561
rect 465154 24325 471918 24561
rect 472154 24325 478918 24561
rect 479154 24325 485918 24561
rect 486154 24325 492918 24561
rect 493154 24325 499918 24561
rect 500154 24325 506918 24561
rect 507154 24325 513918 24561
rect 514154 24325 520918 24561
rect 521154 24325 527918 24561
rect 528154 24325 534918 24561
rect 535154 24325 541918 24561
rect 542154 24325 548918 24561
rect 549154 24325 555918 24561
rect 556154 24325 562918 24561
rect 563154 24325 569918 24561
rect 570154 24325 576918 24561
rect 577154 24325 587570 24561
rect 587806 24325 587890 24561
rect 588126 24325 588210 24561
rect 588446 24325 588530 24561
rect 588766 24325 588874 24561
rect -4950 24283 588874 24325
rect -4950 23494 588874 23536
rect -4950 23258 -3090 23494
rect -2854 23258 -2770 23494
rect -2534 23258 -2450 23494
rect -2214 23258 -2130 23494
rect -1894 23258 1186 23494
rect 1422 23258 8186 23494
rect 8422 23258 15186 23494
rect 15422 23258 22186 23494
rect 22422 23258 29186 23494
rect 29422 23258 36186 23494
rect 36422 23258 43186 23494
rect 43422 23258 50186 23494
rect 50422 23258 57186 23494
rect 57422 23258 64186 23494
rect 64422 23258 71186 23494
rect 71422 23258 78186 23494
rect 78422 23258 85186 23494
rect 85422 23258 92186 23494
rect 92422 23258 99186 23494
rect 99422 23258 106186 23494
rect 106422 23258 113186 23494
rect 113422 23258 120186 23494
rect 120422 23258 127186 23494
rect 127422 23258 134186 23494
rect 134422 23258 141186 23494
rect 141422 23258 148186 23494
rect 148422 23258 155186 23494
rect 155422 23258 162186 23494
rect 162422 23258 169186 23494
rect 169422 23258 176186 23494
rect 176422 23258 183186 23494
rect 183422 23258 190186 23494
rect 190422 23258 197186 23494
rect 197422 23258 204186 23494
rect 204422 23258 211186 23494
rect 211422 23258 218186 23494
rect 218422 23258 225186 23494
rect 225422 23258 232186 23494
rect 232422 23258 239186 23494
rect 239422 23258 246186 23494
rect 246422 23258 253186 23494
rect 253422 23258 260186 23494
rect 260422 23258 267186 23494
rect 267422 23258 274186 23494
rect 274422 23258 281186 23494
rect 281422 23258 288186 23494
rect 288422 23258 295186 23494
rect 295422 23258 302186 23494
rect 302422 23258 309186 23494
rect 309422 23258 316186 23494
rect 316422 23258 323186 23494
rect 323422 23258 330186 23494
rect 330422 23258 337186 23494
rect 337422 23258 344186 23494
rect 344422 23258 351186 23494
rect 351422 23258 358186 23494
rect 358422 23258 365186 23494
rect 365422 23258 372186 23494
rect 372422 23258 379186 23494
rect 379422 23258 386186 23494
rect 386422 23258 393186 23494
rect 393422 23258 400186 23494
rect 400422 23258 407186 23494
rect 407422 23258 414186 23494
rect 414422 23258 421186 23494
rect 421422 23258 428186 23494
rect 428422 23258 435186 23494
rect 435422 23258 442186 23494
rect 442422 23258 449186 23494
rect 449422 23258 456186 23494
rect 456422 23258 463186 23494
rect 463422 23258 470186 23494
rect 470422 23258 477186 23494
rect 477422 23258 484186 23494
rect 484422 23258 491186 23494
rect 491422 23258 498186 23494
rect 498422 23258 505186 23494
rect 505422 23258 512186 23494
rect 512422 23258 519186 23494
rect 519422 23258 526186 23494
rect 526422 23258 533186 23494
rect 533422 23258 540186 23494
rect 540422 23258 547186 23494
rect 547422 23258 554186 23494
rect 554422 23258 561186 23494
rect 561422 23258 568186 23494
rect 568422 23258 575186 23494
rect 575422 23258 582186 23494
rect 582422 23258 585818 23494
rect 586054 23258 586138 23494
rect 586374 23258 586458 23494
rect 586694 23258 586778 23494
rect 587014 23258 588874 23494
rect -4950 23216 588874 23258
rect -4950 17561 588874 17603
rect -4950 17325 -4842 17561
rect -4606 17325 -4522 17561
rect -4286 17325 -4202 17561
rect -3966 17325 -3882 17561
rect -3646 17325 2918 17561
rect 3154 17325 9918 17561
rect 10154 17325 16918 17561
rect 17154 17325 23918 17561
rect 24154 17325 30918 17561
rect 31154 17325 37918 17561
rect 38154 17325 44918 17561
rect 45154 17325 51918 17561
rect 52154 17325 58918 17561
rect 59154 17325 65918 17561
rect 66154 17325 72918 17561
rect 73154 17325 79918 17561
rect 80154 17325 86918 17561
rect 87154 17325 93918 17561
rect 94154 17325 100918 17561
rect 101154 17325 107918 17561
rect 108154 17325 114918 17561
rect 115154 17325 121918 17561
rect 122154 17325 128918 17561
rect 129154 17325 135918 17561
rect 136154 17325 142918 17561
rect 143154 17325 149918 17561
rect 150154 17325 156918 17561
rect 157154 17325 163918 17561
rect 164154 17325 170918 17561
rect 171154 17325 177918 17561
rect 178154 17325 184918 17561
rect 185154 17325 191918 17561
rect 192154 17325 198918 17561
rect 199154 17325 205918 17561
rect 206154 17325 212918 17561
rect 213154 17325 219918 17561
rect 220154 17325 226918 17561
rect 227154 17325 233918 17561
rect 234154 17325 240918 17561
rect 241154 17325 247918 17561
rect 248154 17325 254918 17561
rect 255154 17325 261918 17561
rect 262154 17325 268918 17561
rect 269154 17325 275918 17561
rect 276154 17325 282918 17561
rect 283154 17325 289918 17561
rect 290154 17325 296918 17561
rect 297154 17325 303918 17561
rect 304154 17325 310918 17561
rect 311154 17325 317918 17561
rect 318154 17325 324918 17561
rect 325154 17325 331918 17561
rect 332154 17325 338918 17561
rect 339154 17325 345918 17561
rect 346154 17325 352918 17561
rect 353154 17325 359918 17561
rect 360154 17325 366918 17561
rect 367154 17325 373918 17561
rect 374154 17325 380918 17561
rect 381154 17325 387918 17561
rect 388154 17325 394918 17561
rect 395154 17325 401918 17561
rect 402154 17325 408918 17561
rect 409154 17325 415918 17561
rect 416154 17325 422918 17561
rect 423154 17325 429918 17561
rect 430154 17325 436918 17561
rect 437154 17325 443918 17561
rect 444154 17325 450918 17561
rect 451154 17325 457918 17561
rect 458154 17325 464918 17561
rect 465154 17325 471918 17561
rect 472154 17325 478918 17561
rect 479154 17325 485918 17561
rect 486154 17325 492918 17561
rect 493154 17325 499918 17561
rect 500154 17325 506918 17561
rect 507154 17325 513918 17561
rect 514154 17325 520918 17561
rect 521154 17325 527918 17561
rect 528154 17325 534918 17561
rect 535154 17325 541918 17561
rect 542154 17325 548918 17561
rect 549154 17325 555918 17561
rect 556154 17325 562918 17561
rect 563154 17325 569918 17561
rect 570154 17325 576918 17561
rect 577154 17325 587570 17561
rect 587806 17325 587890 17561
rect 588126 17325 588210 17561
rect 588446 17325 588530 17561
rect 588766 17325 588874 17561
rect -4950 17283 588874 17325
rect -4950 16494 588874 16536
rect -4950 16258 -3090 16494
rect -2854 16258 -2770 16494
rect -2534 16258 -2450 16494
rect -2214 16258 -2130 16494
rect -1894 16258 1186 16494
rect 1422 16258 8186 16494
rect 8422 16258 15186 16494
rect 15422 16258 22186 16494
rect 22422 16258 29186 16494
rect 29422 16258 36186 16494
rect 36422 16258 43186 16494
rect 43422 16258 50186 16494
rect 50422 16258 57186 16494
rect 57422 16258 64186 16494
rect 64422 16258 71186 16494
rect 71422 16258 78186 16494
rect 78422 16258 85186 16494
rect 85422 16258 92186 16494
rect 92422 16258 99186 16494
rect 99422 16258 106186 16494
rect 106422 16258 113186 16494
rect 113422 16258 120186 16494
rect 120422 16258 127186 16494
rect 127422 16258 134186 16494
rect 134422 16258 141186 16494
rect 141422 16258 148186 16494
rect 148422 16258 155186 16494
rect 155422 16258 162186 16494
rect 162422 16258 169186 16494
rect 169422 16258 176186 16494
rect 176422 16258 183186 16494
rect 183422 16258 190186 16494
rect 190422 16258 197186 16494
rect 197422 16258 204186 16494
rect 204422 16258 211186 16494
rect 211422 16258 218186 16494
rect 218422 16258 225186 16494
rect 225422 16258 232186 16494
rect 232422 16258 239186 16494
rect 239422 16258 246186 16494
rect 246422 16258 253186 16494
rect 253422 16258 260186 16494
rect 260422 16258 267186 16494
rect 267422 16258 274186 16494
rect 274422 16258 281186 16494
rect 281422 16258 288186 16494
rect 288422 16258 295186 16494
rect 295422 16258 302186 16494
rect 302422 16258 309186 16494
rect 309422 16258 316186 16494
rect 316422 16258 323186 16494
rect 323422 16258 330186 16494
rect 330422 16258 337186 16494
rect 337422 16258 344186 16494
rect 344422 16258 351186 16494
rect 351422 16258 358186 16494
rect 358422 16258 365186 16494
rect 365422 16258 372186 16494
rect 372422 16258 379186 16494
rect 379422 16258 386186 16494
rect 386422 16258 393186 16494
rect 393422 16258 400186 16494
rect 400422 16258 407186 16494
rect 407422 16258 414186 16494
rect 414422 16258 421186 16494
rect 421422 16258 428186 16494
rect 428422 16258 435186 16494
rect 435422 16258 442186 16494
rect 442422 16258 449186 16494
rect 449422 16258 456186 16494
rect 456422 16258 463186 16494
rect 463422 16258 470186 16494
rect 470422 16258 477186 16494
rect 477422 16258 484186 16494
rect 484422 16258 491186 16494
rect 491422 16258 498186 16494
rect 498422 16258 505186 16494
rect 505422 16258 512186 16494
rect 512422 16258 519186 16494
rect 519422 16258 526186 16494
rect 526422 16258 533186 16494
rect 533422 16258 540186 16494
rect 540422 16258 547186 16494
rect 547422 16258 554186 16494
rect 554422 16258 561186 16494
rect 561422 16258 568186 16494
rect 568422 16258 575186 16494
rect 575422 16258 582186 16494
rect 582422 16258 585818 16494
rect 586054 16258 586138 16494
rect 586374 16258 586458 16494
rect 586694 16258 586778 16494
rect 587014 16258 588874 16494
rect -4950 16216 588874 16258
rect -4950 10561 588874 10603
rect -4950 10325 -4842 10561
rect -4606 10325 -4522 10561
rect -4286 10325 -4202 10561
rect -3966 10325 -3882 10561
rect -3646 10325 2918 10561
rect 3154 10325 9918 10561
rect 10154 10325 16918 10561
rect 17154 10325 23918 10561
rect 24154 10325 30918 10561
rect 31154 10325 37918 10561
rect 38154 10325 44918 10561
rect 45154 10325 51918 10561
rect 52154 10325 58918 10561
rect 59154 10325 65918 10561
rect 66154 10325 72918 10561
rect 73154 10325 79918 10561
rect 80154 10325 86918 10561
rect 87154 10325 93918 10561
rect 94154 10325 100918 10561
rect 101154 10325 107918 10561
rect 108154 10325 114918 10561
rect 115154 10325 121918 10561
rect 122154 10325 128918 10561
rect 129154 10325 135918 10561
rect 136154 10325 142918 10561
rect 143154 10325 149918 10561
rect 150154 10325 156918 10561
rect 157154 10325 163918 10561
rect 164154 10325 170918 10561
rect 171154 10325 177918 10561
rect 178154 10325 184918 10561
rect 185154 10325 191918 10561
rect 192154 10325 198918 10561
rect 199154 10325 205918 10561
rect 206154 10325 212918 10561
rect 213154 10325 219918 10561
rect 220154 10325 226918 10561
rect 227154 10325 233918 10561
rect 234154 10325 240918 10561
rect 241154 10325 247918 10561
rect 248154 10325 254918 10561
rect 255154 10325 261918 10561
rect 262154 10325 268918 10561
rect 269154 10325 275918 10561
rect 276154 10325 282918 10561
rect 283154 10325 289918 10561
rect 290154 10325 296918 10561
rect 297154 10325 303918 10561
rect 304154 10325 310918 10561
rect 311154 10325 317918 10561
rect 318154 10325 324918 10561
rect 325154 10325 331918 10561
rect 332154 10325 338918 10561
rect 339154 10325 345918 10561
rect 346154 10325 352918 10561
rect 353154 10325 359918 10561
rect 360154 10325 366918 10561
rect 367154 10325 373918 10561
rect 374154 10325 380918 10561
rect 381154 10325 387918 10561
rect 388154 10325 394918 10561
rect 395154 10325 401918 10561
rect 402154 10325 408918 10561
rect 409154 10325 415918 10561
rect 416154 10325 422918 10561
rect 423154 10325 429918 10561
rect 430154 10325 436918 10561
rect 437154 10325 443918 10561
rect 444154 10325 450918 10561
rect 451154 10325 457918 10561
rect 458154 10325 464918 10561
rect 465154 10325 471918 10561
rect 472154 10325 478918 10561
rect 479154 10325 485918 10561
rect 486154 10325 492918 10561
rect 493154 10325 499918 10561
rect 500154 10325 506918 10561
rect 507154 10325 513918 10561
rect 514154 10325 520918 10561
rect 521154 10325 527918 10561
rect 528154 10325 534918 10561
rect 535154 10325 541918 10561
rect 542154 10325 548918 10561
rect 549154 10325 555918 10561
rect 556154 10325 562918 10561
rect 563154 10325 569918 10561
rect 570154 10325 576918 10561
rect 577154 10325 587570 10561
rect 587806 10325 587890 10561
rect 588126 10325 588210 10561
rect 588446 10325 588530 10561
rect 588766 10325 588874 10561
rect -4950 10283 588874 10325
rect -4950 9494 588874 9536
rect -4950 9258 -3090 9494
rect -2854 9258 -2770 9494
rect -2534 9258 -2450 9494
rect -2214 9258 -2130 9494
rect -1894 9258 1186 9494
rect 1422 9258 8186 9494
rect 8422 9258 15186 9494
rect 15422 9258 22186 9494
rect 22422 9258 29186 9494
rect 29422 9258 36186 9494
rect 36422 9258 43186 9494
rect 43422 9258 50186 9494
rect 50422 9258 57186 9494
rect 57422 9258 64186 9494
rect 64422 9258 71186 9494
rect 71422 9258 78186 9494
rect 78422 9258 85186 9494
rect 85422 9258 92186 9494
rect 92422 9258 99186 9494
rect 99422 9258 106186 9494
rect 106422 9258 113186 9494
rect 113422 9258 120186 9494
rect 120422 9258 127186 9494
rect 127422 9258 134186 9494
rect 134422 9258 141186 9494
rect 141422 9258 148186 9494
rect 148422 9258 155186 9494
rect 155422 9258 162186 9494
rect 162422 9258 169186 9494
rect 169422 9258 176186 9494
rect 176422 9258 183186 9494
rect 183422 9258 190186 9494
rect 190422 9258 197186 9494
rect 197422 9258 204186 9494
rect 204422 9258 211186 9494
rect 211422 9258 218186 9494
rect 218422 9258 225186 9494
rect 225422 9258 232186 9494
rect 232422 9258 239186 9494
rect 239422 9258 246186 9494
rect 246422 9258 253186 9494
rect 253422 9258 260186 9494
rect 260422 9258 267186 9494
rect 267422 9258 274186 9494
rect 274422 9258 281186 9494
rect 281422 9258 288186 9494
rect 288422 9258 295186 9494
rect 295422 9258 302186 9494
rect 302422 9258 309186 9494
rect 309422 9258 316186 9494
rect 316422 9258 323186 9494
rect 323422 9258 330186 9494
rect 330422 9258 337186 9494
rect 337422 9258 344186 9494
rect 344422 9258 351186 9494
rect 351422 9258 358186 9494
rect 358422 9258 365186 9494
rect 365422 9258 372186 9494
rect 372422 9258 379186 9494
rect 379422 9258 386186 9494
rect 386422 9258 393186 9494
rect 393422 9258 400186 9494
rect 400422 9258 407186 9494
rect 407422 9258 414186 9494
rect 414422 9258 421186 9494
rect 421422 9258 428186 9494
rect 428422 9258 435186 9494
rect 435422 9258 442186 9494
rect 442422 9258 449186 9494
rect 449422 9258 456186 9494
rect 456422 9258 463186 9494
rect 463422 9258 470186 9494
rect 470422 9258 477186 9494
rect 477422 9258 484186 9494
rect 484422 9258 491186 9494
rect 491422 9258 498186 9494
rect 498422 9258 505186 9494
rect 505422 9258 512186 9494
rect 512422 9258 519186 9494
rect 519422 9258 526186 9494
rect 526422 9258 533186 9494
rect 533422 9258 540186 9494
rect 540422 9258 547186 9494
rect 547422 9258 554186 9494
rect 554422 9258 561186 9494
rect 561422 9258 568186 9494
rect 568422 9258 575186 9494
rect 575422 9258 582186 9494
rect 582422 9258 585818 9494
rect 586054 9258 586138 9494
rect 586374 9258 586458 9494
rect 586694 9258 586778 9494
rect 587014 9258 588874 9494
rect -4950 9216 588874 9258
rect -4950 3561 588874 3603
rect -4950 3325 -4842 3561
rect -4606 3325 -4522 3561
rect -4286 3325 -4202 3561
rect -3966 3325 -3882 3561
rect -3646 3325 2918 3561
rect 3154 3325 9918 3561
rect 10154 3325 16918 3561
rect 17154 3325 23918 3561
rect 24154 3325 30918 3561
rect 31154 3325 37918 3561
rect 38154 3325 44918 3561
rect 45154 3325 51918 3561
rect 52154 3325 58918 3561
rect 59154 3325 65918 3561
rect 66154 3325 72918 3561
rect 73154 3325 79918 3561
rect 80154 3325 86918 3561
rect 87154 3325 93918 3561
rect 94154 3325 100918 3561
rect 101154 3325 107918 3561
rect 108154 3325 114918 3561
rect 115154 3325 121918 3561
rect 122154 3325 128918 3561
rect 129154 3325 135918 3561
rect 136154 3325 142918 3561
rect 143154 3325 149918 3561
rect 150154 3325 156918 3561
rect 157154 3325 163918 3561
rect 164154 3325 170918 3561
rect 171154 3325 177918 3561
rect 178154 3325 184918 3561
rect 185154 3325 191918 3561
rect 192154 3325 198918 3561
rect 199154 3325 205918 3561
rect 206154 3325 212918 3561
rect 213154 3325 219918 3561
rect 220154 3325 226918 3561
rect 227154 3325 233918 3561
rect 234154 3325 240918 3561
rect 241154 3325 247918 3561
rect 248154 3325 254918 3561
rect 255154 3325 261918 3561
rect 262154 3325 268918 3561
rect 269154 3325 275918 3561
rect 276154 3325 282918 3561
rect 283154 3325 289918 3561
rect 290154 3325 296918 3561
rect 297154 3325 303918 3561
rect 304154 3325 310918 3561
rect 311154 3325 317918 3561
rect 318154 3325 324918 3561
rect 325154 3325 331918 3561
rect 332154 3325 338918 3561
rect 339154 3325 345918 3561
rect 346154 3325 352918 3561
rect 353154 3325 359918 3561
rect 360154 3325 366918 3561
rect 367154 3325 373918 3561
rect 374154 3325 380918 3561
rect 381154 3325 387918 3561
rect 388154 3325 394918 3561
rect 395154 3325 401918 3561
rect 402154 3325 408918 3561
rect 409154 3325 415918 3561
rect 416154 3325 422918 3561
rect 423154 3325 429918 3561
rect 430154 3325 436918 3561
rect 437154 3325 443918 3561
rect 444154 3325 450918 3561
rect 451154 3325 457918 3561
rect 458154 3325 464918 3561
rect 465154 3325 471918 3561
rect 472154 3325 478918 3561
rect 479154 3325 485918 3561
rect 486154 3325 492918 3561
rect 493154 3325 499918 3561
rect 500154 3325 506918 3561
rect 507154 3325 513918 3561
rect 514154 3325 520918 3561
rect 521154 3325 527918 3561
rect 528154 3325 534918 3561
rect 535154 3325 541918 3561
rect 542154 3325 548918 3561
rect 549154 3325 555918 3561
rect 556154 3325 562918 3561
rect 563154 3325 569918 3561
rect 570154 3325 576918 3561
rect 577154 3325 587570 3561
rect 587806 3325 587890 3561
rect 588126 3325 588210 3561
rect 588446 3325 588530 3561
rect 588766 3325 588874 3561
rect -4950 3283 588874 3325
rect -4950 2494 588874 2536
rect -4950 2258 -3090 2494
rect -2854 2258 -2770 2494
rect -2534 2258 -2450 2494
rect -2214 2258 -2130 2494
rect -1894 2258 1186 2494
rect 1422 2258 8186 2494
rect 8422 2258 15186 2494
rect 15422 2258 22186 2494
rect 22422 2258 29186 2494
rect 29422 2258 36186 2494
rect 36422 2258 43186 2494
rect 43422 2258 50186 2494
rect 50422 2258 57186 2494
rect 57422 2258 64186 2494
rect 64422 2258 71186 2494
rect 71422 2258 78186 2494
rect 78422 2258 85186 2494
rect 85422 2258 92186 2494
rect 92422 2258 99186 2494
rect 99422 2258 106186 2494
rect 106422 2258 113186 2494
rect 113422 2258 120186 2494
rect 120422 2258 127186 2494
rect 127422 2258 134186 2494
rect 134422 2258 141186 2494
rect 141422 2258 148186 2494
rect 148422 2258 155186 2494
rect 155422 2258 162186 2494
rect 162422 2258 169186 2494
rect 169422 2258 176186 2494
rect 176422 2258 183186 2494
rect 183422 2258 190186 2494
rect 190422 2258 197186 2494
rect 197422 2258 204186 2494
rect 204422 2258 211186 2494
rect 211422 2258 218186 2494
rect 218422 2258 225186 2494
rect 225422 2258 232186 2494
rect 232422 2258 239186 2494
rect 239422 2258 246186 2494
rect 246422 2258 253186 2494
rect 253422 2258 260186 2494
rect 260422 2258 267186 2494
rect 267422 2258 274186 2494
rect 274422 2258 281186 2494
rect 281422 2258 288186 2494
rect 288422 2258 295186 2494
rect 295422 2258 302186 2494
rect 302422 2258 309186 2494
rect 309422 2258 316186 2494
rect 316422 2258 323186 2494
rect 323422 2258 330186 2494
rect 330422 2258 337186 2494
rect 337422 2258 344186 2494
rect 344422 2258 351186 2494
rect 351422 2258 358186 2494
rect 358422 2258 365186 2494
rect 365422 2258 372186 2494
rect 372422 2258 379186 2494
rect 379422 2258 386186 2494
rect 386422 2258 393186 2494
rect 393422 2258 400186 2494
rect 400422 2258 407186 2494
rect 407422 2258 414186 2494
rect 414422 2258 421186 2494
rect 421422 2258 428186 2494
rect 428422 2258 435186 2494
rect 435422 2258 442186 2494
rect 442422 2258 449186 2494
rect 449422 2258 456186 2494
rect 456422 2258 463186 2494
rect 463422 2258 470186 2494
rect 470422 2258 477186 2494
rect 477422 2258 484186 2494
rect 484422 2258 491186 2494
rect 491422 2258 498186 2494
rect 498422 2258 505186 2494
rect 505422 2258 512186 2494
rect 512422 2258 519186 2494
rect 519422 2258 526186 2494
rect 526422 2258 533186 2494
rect 533422 2258 540186 2494
rect 540422 2258 547186 2494
rect 547422 2258 554186 2494
rect 554422 2258 561186 2494
rect 561422 2258 568186 2494
rect 568422 2258 575186 2494
rect 575422 2258 582186 2494
rect 582422 2258 585818 2494
rect 586054 2258 586138 2494
rect 586374 2258 586458 2494
rect 586694 2258 586778 2494
rect 587014 2258 588874 2494
rect -4950 2216 588874 2258
rect -2406 -746 587122 -714
rect -2406 -982 -2374 -746
rect -2138 -982 -2054 -746
rect -1818 -982 1186 -746
rect 1422 -982 8186 -746
rect 8422 -982 15186 -746
rect 15422 -982 22186 -746
rect 22422 -982 29186 -746
rect 29422 -982 36186 -746
rect 36422 -982 43186 -746
rect 43422 -982 50186 -746
rect 50422 -982 57186 -746
rect 57422 -982 64186 -746
rect 64422 -982 71186 -746
rect 71422 -982 78186 -746
rect 78422 -982 85186 -746
rect 85422 -982 92186 -746
rect 92422 -982 99186 -746
rect 99422 -982 106186 -746
rect 106422 -982 113186 -746
rect 113422 -982 120186 -746
rect 120422 -982 127186 -746
rect 127422 -982 134186 -746
rect 134422 -982 141186 -746
rect 141422 -982 148186 -746
rect 148422 -982 155186 -746
rect 155422 -982 162186 -746
rect 162422 -982 169186 -746
rect 169422 -982 176186 -746
rect 176422 -982 183186 -746
rect 183422 -982 190186 -746
rect 190422 -982 197186 -746
rect 197422 -982 204186 -746
rect 204422 -982 211186 -746
rect 211422 -982 218186 -746
rect 218422 -982 225186 -746
rect 225422 -982 232186 -746
rect 232422 -982 239186 -746
rect 239422 -982 246186 -746
rect 246422 -982 253186 -746
rect 253422 -982 260186 -746
rect 260422 -982 267186 -746
rect 267422 -982 274186 -746
rect 274422 -982 281186 -746
rect 281422 -982 288186 -746
rect 288422 -982 295186 -746
rect 295422 -982 302186 -746
rect 302422 -982 309186 -746
rect 309422 -982 316186 -746
rect 316422 -982 323186 -746
rect 323422 -982 330186 -746
rect 330422 -982 337186 -746
rect 337422 -982 344186 -746
rect 344422 -982 351186 -746
rect 351422 -982 358186 -746
rect 358422 -982 365186 -746
rect 365422 -982 372186 -746
rect 372422 -982 379186 -746
rect 379422 -982 386186 -746
rect 386422 -982 393186 -746
rect 393422 -982 400186 -746
rect 400422 -982 407186 -746
rect 407422 -982 414186 -746
rect 414422 -982 421186 -746
rect 421422 -982 428186 -746
rect 428422 -982 435186 -746
rect 435422 -982 442186 -746
rect 442422 -982 449186 -746
rect 449422 -982 456186 -746
rect 456422 -982 463186 -746
rect 463422 -982 470186 -746
rect 470422 -982 477186 -746
rect 477422 -982 484186 -746
rect 484422 -982 491186 -746
rect 491422 -982 498186 -746
rect 498422 -982 505186 -746
rect 505422 -982 512186 -746
rect 512422 -982 519186 -746
rect 519422 -982 526186 -746
rect 526422 -982 533186 -746
rect 533422 -982 540186 -746
rect 540422 -982 547186 -746
rect 547422 -982 554186 -746
rect 554422 -982 561186 -746
rect 561422 -982 568186 -746
rect 568422 -982 575186 -746
rect 575422 -982 582186 -746
rect 582422 -982 585818 -746
rect 586054 -982 586138 -746
rect 586374 -982 586458 -746
rect 586694 -982 586778 -746
rect 587014 -982 587122 -746
rect -2406 -1066 587122 -982
rect -2406 -1302 -2374 -1066
rect -2138 -1302 -2054 -1066
rect -1818 -1302 1186 -1066
rect 1422 -1302 8186 -1066
rect 8422 -1302 15186 -1066
rect 15422 -1302 22186 -1066
rect 22422 -1302 29186 -1066
rect 29422 -1302 36186 -1066
rect 36422 -1302 43186 -1066
rect 43422 -1302 50186 -1066
rect 50422 -1302 57186 -1066
rect 57422 -1302 64186 -1066
rect 64422 -1302 71186 -1066
rect 71422 -1302 78186 -1066
rect 78422 -1302 85186 -1066
rect 85422 -1302 92186 -1066
rect 92422 -1302 99186 -1066
rect 99422 -1302 106186 -1066
rect 106422 -1302 113186 -1066
rect 113422 -1302 120186 -1066
rect 120422 -1302 127186 -1066
rect 127422 -1302 134186 -1066
rect 134422 -1302 141186 -1066
rect 141422 -1302 148186 -1066
rect 148422 -1302 155186 -1066
rect 155422 -1302 162186 -1066
rect 162422 -1302 169186 -1066
rect 169422 -1302 176186 -1066
rect 176422 -1302 183186 -1066
rect 183422 -1302 190186 -1066
rect 190422 -1302 197186 -1066
rect 197422 -1302 204186 -1066
rect 204422 -1302 211186 -1066
rect 211422 -1302 218186 -1066
rect 218422 -1302 225186 -1066
rect 225422 -1302 232186 -1066
rect 232422 -1302 239186 -1066
rect 239422 -1302 246186 -1066
rect 246422 -1302 253186 -1066
rect 253422 -1302 260186 -1066
rect 260422 -1302 267186 -1066
rect 267422 -1302 274186 -1066
rect 274422 -1302 281186 -1066
rect 281422 -1302 288186 -1066
rect 288422 -1302 295186 -1066
rect 295422 -1302 302186 -1066
rect 302422 -1302 309186 -1066
rect 309422 -1302 316186 -1066
rect 316422 -1302 323186 -1066
rect 323422 -1302 330186 -1066
rect 330422 -1302 337186 -1066
rect 337422 -1302 344186 -1066
rect 344422 -1302 351186 -1066
rect 351422 -1302 358186 -1066
rect 358422 -1302 365186 -1066
rect 365422 -1302 372186 -1066
rect 372422 -1302 379186 -1066
rect 379422 -1302 386186 -1066
rect 386422 -1302 393186 -1066
rect 393422 -1302 400186 -1066
rect 400422 -1302 407186 -1066
rect 407422 -1302 414186 -1066
rect 414422 -1302 421186 -1066
rect 421422 -1302 428186 -1066
rect 428422 -1302 435186 -1066
rect 435422 -1302 442186 -1066
rect 442422 -1302 449186 -1066
rect 449422 -1302 456186 -1066
rect 456422 -1302 463186 -1066
rect 463422 -1302 470186 -1066
rect 470422 -1302 477186 -1066
rect 477422 -1302 484186 -1066
rect 484422 -1302 491186 -1066
rect 491422 -1302 498186 -1066
rect 498422 -1302 505186 -1066
rect 505422 -1302 512186 -1066
rect 512422 -1302 519186 -1066
rect 519422 -1302 526186 -1066
rect 526422 -1302 533186 -1066
rect 533422 -1302 540186 -1066
rect 540422 -1302 547186 -1066
rect 547422 -1302 554186 -1066
rect 554422 -1302 561186 -1066
rect 561422 -1302 568186 -1066
rect 568422 -1302 575186 -1066
rect 575422 -1302 582186 -1066
rect 582422 -1302 585818 -1066
rect 586054 -1302 586138 -1066
rect 586374 -1302 586458 -1066
rect 586694 -1302 586778 -1066
rect 587014 -1302 587122 -1066
rect -2406 -1334 587122 -1302
rect -3366 -1706 587290 -1674
rect -3366 -1942 2918 -1706
rect 3154 -1942 9918 -1706
rect 10154 -1942 16918 -1706
rect 17154 -1942 23918 -1706
rect 24154 -1942 30918 -1706
rect 31154 -1942 37918 -1706
rect 38154 -1942 44918 -1706
rect 45154 -1942 51918 -1706
rect 52154 -1942 58918 -1706
rect 59154 -1942 65918 -1706
rect 66154 -1942 72918 -1706
rect 73154 -1942 79918 -1706
rect 80154 -1942 86918 -1706
rect 87154 -1942 93918 -1706
rect 94154 -1942 100918 -1706
rect 101154 -1942 107918 -1706
rect 108154 -1942 114918 -1706
rect 115154 -1942 121918 -1706
rect 122154 -1942 128918 -1706
rect 129154 -1942 135918 -1706
rect 136154 -1942 142918 -1706
rect 143154 -1942 149918 -1706
rect 150154 -1942 156918 -1706
rect 157154 -1942 163918 -1706
rect 164154 -1942 170918 -1706
rect 171154 -1942 177918 -1706
rect 178154 -1942 184918 -1706
rect 185154 -1942 191918 -1706
rect 192154 -1942 198918 -1706
rect 199154 -1942 205918 -1706
rect 206154 -1942 212918 -1706
rect 213154 -1942 219918 -1706
rect 220154 -1942 226918 -1706
rect 227154 -1942 233918 -1706
rect 234154 -1942 240918 -1706
rect 241154 -1942 247918 -1706
rect 248154 -1942 254918 -1706
rect 255154 -1942 261918 -1706
rect 262154 -1942 268918 -1706
rect 269154 -1942 275918 -1706
rect 276154 -1942 282918 -1706
rect 283154 -1942 289918 -1706
rect 290154 -1942 296918 -1706
rect 297154 -1942 303918 -1706
rect 304154 -1942 310918 -1706
rect 311154 -1942 317918 -1706
rect 318154 -1942 324918 -1706
rect 325154 -1942 331918 -1706
rect 332154 -1942 338918 -1706
rect 339154 -1942 345918 -1706
rect 346154 -1942 352918 -1706
rect 353154 -1942 359918 -1706
rect 360154 -1942 366918 -1706
rect 367154 -1942 373918 -1706
rect 374154 -1942 380918 -1706
rect 381154 -1942 387918 -1706
rect 388154 -1942 394918 -1706
rect 395154 -1942 401918 -1706
rect 402154 -1942 408918 -1706
rect 409154 -1942 415918 -1706
rect 416154 -1942 422918 -1706
rect 423154 -1942 429918 -1706
rect 430154 -1942 436918 -1706
rect 437154 -1942 443918 -1706
rect 444154 -1942 450918 -1706
rect 451154 -1942 457918 -1706
rect 458154 -1942 464918 -1706
rect 465154 -1942 471918 -1706
rect 472154 -1942 478918 -1706
rect 479154 -1942 485918 -1706
rect 486154 -1942 492918 -1706
rect 493154 -1942 499918 -1706
rect 500154 -1942 506918 -1706
rect 507154 -1942 513918 -1706
rect 514154 -1942 520918 -1706
rect 521154 -1942 527918 -1706
rect 528154 -1942 534918 -1706
rect 535154 -1942 541918 -1706
rect 542154 -1942 548918 -1706
rect 549154 -1942 555918 -1706
rect 556154 -1942 562918 -1706
rect 563154 -1942 569918 -1706
rect 570154 -1942 576918 -1706
rect 577154 -1942 587290 -1706
rect -3366 -2026 587290 -1942
rect -3366 -2262 2918 -2026
rect 3154 -2262 9918 -2026
rect 10154 -2262 16918 -2026
rect 17154 -2262 23918 -2026
rect 24154 -2262 30918 -2026
rect 31154 -2262 37918 -2026
rect 38154 -2262 44918 -2026
rect 45154 -2262 51918 -2026
rect 52154 -2262 58918 -2026
rect 59154 -2262 65918 -2026
rect 66154 -2262 72918 -2026
rect 73154 -2262 79918 -2026
rect 80154 -2262 86918 -2026
rect 87154 -2262 93918 -2026
rect 94154 -2262 100918 -2026
rect 101154 -2262 107918 -2026
rect 108154 -2262 114918 -2026
rect 115154 -2262 121918 -2026
rect 122154 -2262 128918 -2026
rect 129154 -2262 135918 -2026
rect 136154 -2262 142918 -2026
rect 143154 -2262 149918 -2026
rect 150154 -2262 156918 -2026
rect 157154 -2262 163918 -2026
rect 164154 -2262 170918 -2026
rect 171154 -2262 177918 -2026
rect 178154 -2262 184918 -2026
rect 185154 -2262 191918 -2026
rect 192154 -2262 198918 -2026
rect 199154 -2262 205918 -2026
rect 206154 -2262 212918 -2026
rect 213154 -2262 219918 -2026
rect 220154 -2262 226918 -2026
rect 227154 -2262 233918 -2026
rect 234154 -2262 240918 -2026
rect 241154 -2262 247918 -2026
rect 248154 -2262 254918 -2026
rect 255154 -2262 261918 -2026
rect 262154 -2262 268918 -2026
rect 269154 -2262 275918 -2026
rect 276154 -2262 282918 -2026
rect 283154 -2262 289918 -2026
rect 290154 -2262 296918 -2026
rect 297154 -2262 303918 -2026
rect 304154 -2262 310918 -2026
rect 311154 -2262 317918 -2026
rect 318154 -2262 324918 -2026
rect 325154 -2262 331918 -2026
rect 332154 -2262 338918 -2026
rect 339154 -2262 345918 -2026
rect 346154 -2262 352918 -2026
rect 353154 -2262 359918 -2026
rect 360154 -2262 366918 -2026
rect 367154 -2262 373918 -2026
rect 374154 -2262 380918 -2026
rect 381154 -2262 387918 -2026
rect 388154 -2262 394918 -2026
rect 395154 -2262 401918 -2026
rect 402154 -2262 408918 -2026
rect 409154 -2262 415918 -2026
rect 416154 -2262 422918 -2026
rect 423154 -2262 429918 -2026
rect 430154 -2262 436918 -2026
rect 437154 -2262 443918 -2026
rect 444154 -2262 450918 -2026
rect 451154 -2262 457918 -2026
rect 458154 -2262 464918 -2026
rect 465154 -2262 471918 -2026
rect 472154 -2262 478918 -2026
rect 479154 -2262 485918 -2026
rect 486154 -2262 492918 -2026
rect 493154 -2262 499918 -2026
rect 500154 -2262 506918 -2026
rect 507154 -2262 513918 -2026
rect 514154 -2262 520918 -2026
rect 521154 -2262 527918 -2026
rect 528154 -2262 534918 -2026
rect 535154 -2262 541918 -2026
rect 542154 -2262 548918 -2026
rect 549154 -2262 555918 -2026
rect 556154 -2262 562918 -2026
rect 563154 -2262 569918 -2026
rect 570154 -2262 576918 -2026
rect 577154 -2262 587290 -2026
rect -3366 -2294 587290 -2262
use mux16x1_project  mprj1
timestamp 0
transform 1 0 518000 0 1 400000
box 0 552 10000 22000
use mux16x1_project  mprj2
timestamp 0
transform 1 0 518000 0 1 360000
box 0 552 10000 22000
use mux16x1_project  mprj3
timestamp 0
transform 1 0 518000 0 1 320000
box 0 552 10000 22000
use mux16x1_project  mprj4
timestamp 0
transform 1 0 518000 0 1 280000
box 0 552 10000 22000
use mux16x1_project  mprj5
timestamp 0
transform 1 0 518000 0 1 240000
box 0 552 10000 22000
use sky130_osu_ring_oscillator_mpr2aa_8_b0r1  ro1
timestamp 0
transform 1 0 295144 0 1 489170
box 0 0 16345 2492
use sky130_osu_ring_oscillator_mpr2at_8_b0r1  ro2
timestamp 0
transform 1 0 292553 0 1 470600
box 2591 0 21079 2522
use sky130_osu_ring_oscillator_mpr2ca_8_b0r1  ro3
timestamp 0
transform 1 0 295144 0 1 449600
box 3 0 17148 2491
use sky130_osu_ring_oscillator_mpr2ct_8_b0r1  ro4
timestamp 0
transform 1 0 295147 0 1 428859
box -3 -259 17782 2233
use sky130_osu_ring_oscillator_mpr2ea_8_b0r1  ro5
timestamp 0
transform 1 0 293164 0 1 407600
box 1980 0 18866 2492
use sky130_osu_ring_oscillator_mpr2et_8_b0r1  ro6
timestamp 0
transform 1 0 292719 0 1 386600
box 2425 0 21548 2493
use sky130_osu_ring_oscillator_mpr2xa_8_b0r1  ro7
timestamp 0
transform 1 0 293378 0 1 365600
box 1766 0 17585 2493
use sky130_osu_ring_oscillator_mpr2ya_8_b0r1  ro8
timestamp 0
transform 1 0 295144 0 1 344600
box 5 0 15825 2493
use sky130_osu_ring_oscillator_mpr2aa_8_b0r2  ro9
timestamp 0
transform 1 0 293262 0 1 323600
box 1882 0 18237 2492
use sky130_osu_ring_oscillator_mpr2at_8_b0r2  ro10
timestamp 0
transform 1 0 295144 0 1 302600
box 4 0 18521 2522
use sky130_osu_ring_oscillator_mpr2ca_8_b0r2  ro11
timestamp 0
transform 1 0 293154 0 1 281600
box 1990 0 19207 2494
use sky130_osu_ring_oscillator_mpr2ct_8_b0r2  ro12
timestamp 0
transform 1 0 295144 0 1 260600
box 1 0 17784 2493
use sky130_osu_ring_oscillator_mpr2ea_8_b0r2  ro13
timestamp 0
transform 1 0 293164 0 1 239600
box 1980 0 18865 2492
use sky130_osu_ring_oscillator_mpr2et_8_b0r2  ro14
timestamp 0
transform 1 0 292718 0 1 218600
box 2426 0 21546 2495
use sky130_osu_ring_oscillator_mpr2xa_8_b0r2  ro15
timestamp 0
transform 1 0 295143 0 1 197599
box 1 1 15820 2494
use sky130_osu_ring_oscillator_mpr2ya_8_b0r2  ro16
timestamp 0
transform 1 0 295144 0 1 176800
box 0 0 15821 2493
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal4 s -3198 -2126 -1786 706062 0 FreeSans 7680 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -2406 -1334 587122 -714 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -2406 704650 587122 705270 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 585710 -2126 587122 706062 0 FreeSans 7680 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 1144 -2294 1464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 8144 -2294 8464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 15144 -2294 15464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 22144 -2294 22464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 29144 -2294 29464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 36144 -2294 36464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 43144 -2294 43464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 50144 -2294 50464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 57144 -2294 57464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 64144 -2294 64464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 71144 -2294 71464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 78144 -2294 78464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 85144 -2294 85464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 92144 -2294 92464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 99144 -2294 99464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 106144 -2294 106464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 113144 -2294 113464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 120144 -2294 120464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 127144 -2294 127464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 134144 -2294 134464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 141144 -2294 141464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 148144 -2294 148464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 155144 -2294 155464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 162144 -2294 162464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 169144 -2294 169464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 176144 -2294 176464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 183144 -2294 183464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 190144 -2294 190464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 197144 -2294 197464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 204144 -2294 204464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 211144 -2294 211464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 218144 -2294 218464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 225144 -2294 225464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 232144 -2294 232464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 239144 -2294 239464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 246144 -2294 246464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 253144 -2294 253464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 260144 -2294 260464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 267144 -2294 267464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 274144 -2294 274464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 281144 -2294 281464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 288144 -2294 288464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 295144 -2294 295464 196236 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 295144 200640 295464 364236 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 295144 368640 295464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 302144 -2294 302464 196236 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 302144 200640 302464 364236 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 302144 368640 302464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 309144 -2294 309464 196236 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 309144 200640 309464 364236 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 309144 368640 309464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 316144 -2294 316464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 323144 -2294 323464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 330144 -2294 330464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 337144 -2294 337464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 344144 -2294 344464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 351144 -2294 351464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 358144 -2294 358464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 365144 -2294 365464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 372144 -2294 372464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 379144 -2294 379464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 386144 -2294 386464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 393144 -2294 393464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 400144 -2294 400464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 407144 -2294 407464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 414144 -2294 414464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 421144 -2294 421464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 428144 -2294 428464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 435144 -2294 435464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 442144 -2294 442464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 449144 -2294 449464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 456144 -2294 456464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 463144 -2294 463464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 470144 -2294 470464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 477144 -2294 477464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 484144 -2294 484464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 491144 -2294 491464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 498144 -2294 498464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 505144 -2294 505464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 512144 -2294 512464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 519144 -2294 519464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 -2294 526464 240008 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 261752 526464 280008 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 301752 526464 320008 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 341752 526464 360008 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 381752 526464 400008 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 526144 421752 526464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 533144 -2294 533464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 540144 -2294 540464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 547144 -2294 547464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 554144 -2294 554464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 561144 -2294 561464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 568144 -2294 568464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 575144 -2294 575464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 582144 -2294 582464 706230 0 FreeSans 1920 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 2216 588874 2536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 9216 588874 9536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 16216 588874 16536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 23216 588874 23536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 30216 588874 30536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 37216 588874 37536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 44216 588874 44536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 51216 588874 51536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 58216 588874 58536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 65216 588874 65536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 72216 588874 72536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 79216 588874 79536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 86216 588874 86536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 93216 588874 93536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 100216 588874 100536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 107216 588874 107536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 114216 588874 114536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 121216 588874 121536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 128216 588874 128536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 135216 588874 135536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 142216 588874 142536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 149216 588874 149536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 156216 588874 156536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 163216 588874 163536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 170216 588874 170536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 177216 588874 177536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 184216 588874 184536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 191216 588874 191536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 198216 588874 198536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 205216 588874 205536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 212216 588874 212536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 219216 588874 219536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 226216 588874 226536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 233216 588874 233536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 240216 588874 240536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 247216 588874 247536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 254216 588874 254536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 261216 588874 261536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 268216 588874 268536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 275216 588874 275536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 282216 588874 282536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 289216 588874 289536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 296216 588874 296536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 303216 588874 303536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 310216 588874 310536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 317216 588874 317536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 324216 588874 324536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 331216 588874 331536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 338216 588874 338536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 345216 588874 345536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 352216 588874 352536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 359216 588874 359536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 366216 588874 366536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 373216 588874 373536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 380216 588874 380536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 387216 588874 387536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 394216 588874 394536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 401216 588874 401536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 408216 588874 408536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 415216 588874 415536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 422216 588874 422536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 429216 588874 429536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 436216 588874 436536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 443216 588874 443536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 450216 588874 450536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 457216 588874 457536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 464216 588874 464536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 471216 588874 471536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 478216 588874 478536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 485216 588874 485536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 492216 588874 492536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 499216 588874 499536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 506216 588874 506536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 513216 588874 513536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 520216 588874 520536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 527216 588874 527536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 534216 588874 534536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 541216 588874 541536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 548216 588874 548536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 555216 588874 555536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 562216 588874 562536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 569216 588874 569536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 576216 588874 576536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 583216 588874 583536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 590216 588874 590536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 597216 588874 597536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 604216 588874 604536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 611216 588874 611536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 618216 588874 618536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 625216 588874 625536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 632216 588874 632536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 639216 588874 639536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 646216 588874 646536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 653216 588874 653536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 660216 588874 660536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 667216 588874 667536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 674216 588874 674536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 681216 588874 681536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 688216 588874 688536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -4950 695216 588874 695536 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s -4950 -3878 -3538 707814 0 FreeSans 7680 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3366 -2294 587290 -1674 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3366 705610 587290 706230 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 587462 -3878 588874 707814 0 FreeSans 7680 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 2876 -2294 3196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 9876 -2294 10196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 16876 -2294 17196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 23876 -2294 24196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 30876 -2294 31196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 37876 -2294 38196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 44876 -2294 45196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 51876 -2294 52196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 58876 -2294 59196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 65876 -2294 66196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 72876 -2294 73196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 79876 -2294 80196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 86876 -2294 87196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 93876 -2294 94196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 100876 -2294 101196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 107876 -2294 108196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 114876 -2294 115196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 121876 -2294 122196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 128876 -2294 129196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 135876 -2294 136196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 142876 -2294 143196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 149876 -2294 150196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 156876 -2294 157196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 163876 -2294 164196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 170876 -2294 171196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 177876 -2294 178196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 184876 -2294 185196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 191876 -2294 192196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 198876 -2294 199196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 205876 -2294 206196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 212876 -2294 213196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 219876 -2294 220196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 226876 -2294 227196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 233876 -2294 234196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 240876 -2294 241196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 247876 -2294 248196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 254876 -2294 255196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 261876 -2294 262196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 268876 -2294 269196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 275876 -2294 276196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 282876 -2294 283196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 289876 -2294 290196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 296876 -2294 297196 196236 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 296876 200640 297196 364236 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 296876 368640 297196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 303876 -2294 304196 196236 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 303876 200640 304196 364236 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 303876 368640 304196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 310876 -2294 311196 196236 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 310876 200547 311196 364236 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 310876 368547 311196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 317876 -2294 318196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 324876 -2294 325196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 331876 -2294 332196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 338876 -2294 339196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 345876 -2294 346196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 352876 -2294 353196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 359876 -2294 360196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 366876 -2294 367196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 373876 -2294 374196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 380876 -2294 381196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 387876 -2294 388196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 394876 -2294 395196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 401876 -2294 402196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 408876 -2294 409196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 415876 -2294 416196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 422876 -2294 423196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 429876 -2294 430196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 436876 -2294 437196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 443876 -2294 444196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 450876 -2294 451196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 457876 -2294 458196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 464876 -2294 465196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 471876 -2294 472196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 478876 -2294 479196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 485876 -2294 486196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 492876 -2294 493196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 499876 -2294 500196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 506876 -2294 507196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 513876 -2294 514196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 -2294 521196 240008 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 261752 521196 280008 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 301752 521196 320008 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 341752 521196 360008 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 381752 521196 400008 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 520876 421752 521196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 527876 -2294 528196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 534876 -2294 535196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 541876 -2294 542196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 548876 -2294 549196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 555876 -2294 556196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 562876 -2294 563196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 569876 -2294 570196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 576876 -2294 577196 706230 0 FreeSans 1920 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 3283 588874 3603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 10283 588874 10603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 17283 588874 17603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 24283 588874 24603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 31283 588874 31603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 38283 588874 38603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 45283 588874 45603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 52283 588874 52603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 59283 588874 59603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 66283 588874 66603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 73283 588874 73603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 80283 588874 80603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 87283 588874 87603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 94283 588874 94603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 101283 588874 101603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 108283 588874 108603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 115283 588874 115603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 122283 588874 122603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 129283 588874 129603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 136283 588874 136603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 143283 588874 143603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 150283 588874 150603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 157283 588874 157603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 164283 588874 164603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 171283 588874 171603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 178283 588874 178603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 185283 588874 185603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 192283 588874 192603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 199283 588874 199603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 206283 588874 206603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 213283 588874 213603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 220283 588874 220603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 227283 588874 227603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 234283 588874 234603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 241283 588874 241603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 248283 588874 248603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 255283 588874 255603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 262283 588874 262603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 269283 588874 269603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 276283 588874 276603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 283283 588874 283603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 290283 588874 290603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 297283 588874 297603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 304283 588874 304603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 311283 588874 311603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 318283 588874 318603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 325283 588874 325603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 332283 588874 332603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 339283 588874 339603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 346283 588874 346603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 353283 588874 353603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 360283 588874 360603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 367283 588874 367603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 374283 588874 374603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 381283 588874 381603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 388283 588874 388603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 395283 588874 395603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 402283 588874 402603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 409283 588874 409603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 416283 588874 416603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 423283 588874 423603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 430283 588874 430603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 437283 588874 437603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 444283 588874 444603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 451283 588874 451603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 458283 588874 458603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 465283 588874 465603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 472283 588874 472603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 479283 588874 479603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 486283 588874 486603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 493283 588874 493603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 500283 588874 500603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 507283 588874 507603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 514283 588874 514603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 521283 588874 521603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 528283 588874 528603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 535283 588874 535603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 542283 588874 542603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 549283 588874 549603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 556283 588874 556603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 563283 588874 563603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 570283 588874 570603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 577283 588874 577603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 584283 588874 584603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 591283 588874 591603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 598283 588874 598603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 605283 588874 605603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 612283 588874 612603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 619283 588874 619603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 626283 588874 626603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 633283 588874 633603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 640283 588874 640603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 647283 588874 647603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 654283 588874 654603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 661283 588874 661603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 668283 588874 668603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 675283 588874 675603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 682283 588874 682603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 689283 588874 689603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -4950 696283 588874 696603 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 145 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 146 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 147 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 148 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 149 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 150 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 151 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 152 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 153 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 154 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 155 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 156 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 157 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 158 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 159 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 160 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 161 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 162 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 163 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 164 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 165 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 166 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 167 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 168 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 169 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 170 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 171 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 172 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 173 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 174 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 175 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 176 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 177 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 178 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 179 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 180 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 181 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 182 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 183 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 184 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 185 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 186 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 187 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 188 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 189 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 190 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 191 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 192 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 193 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 194 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 195 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 196 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 197 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 198 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 199 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 200 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 201 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 202 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 203 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 204 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 205 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 206 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 207 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 208 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 209 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 210 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 211 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 212 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 213 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 214 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 215 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 216 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 217 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 218 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 219 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 220 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 221 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 222 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 223 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 224 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 225 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 226 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 227 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 228 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 229 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 230 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 231 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 232 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 233 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 234 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 235 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 236 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 237 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 238 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 239 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 240 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 241 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 242 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 243 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 244 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 245 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 246 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 247 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 248 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 249 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 250 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
