magic
tech sky130A
magscale 1 2
timestamp 1699645154
<< viali >>
rect 301934 490569 301968 490603
rect 295770 450109 295804 450143
rect 299087 450109 299121 450143
rect 299342 430593 299376 430627
rect 298982 410601 299016 410635
rect 305512 410601 305546 410635
rect 303587 390609 303621 390643
rect 307712 370617 307746 370651
rect 299340 270589 299374 270623
rect 298981 250597 299015 250631
rect 305511 250597 305545 250631
rect 303587 230605 303621 230639
rect 295503 210613 295537 210647
rect 307711 210613 307745 210647
<< metal1 >>
rect 289722 490900 289728 490952
rect 289780 490940 289786 490952
rect 292040 490940 292068 491208
rect 289780 490912 292068 490940
rect 289780 490900 289786 490912
rect 301958 490609 301964 490612
rect 301922 490603 301964 490609
rect 301922 490569 301934 490603
rect 301922 490563 301964 490569
rect 301958 490560 301964 490563
rect 302016 490560 302022 490612
rect 295616 490228 295668 490234
rect 295616 490170 295668 490176
rect 298744 490228 298796 490234
rect 298744 490170 298796 490176
rect 305092 490228 305144 490234
rect 305092 490170 305144 490176
rect 308232 490056 308260 490202
rect 311158 490056 311164 490068
rect 308232 490028 311164 490056
rect 311158 490016 311164 490028
rect 311216 490016 311222 490068
rect 298738 487228 298744 487280
rect 298796 487268 298802 487280
rect 322198 487268 322204 487280
rect 298796 487240 322204 487268
rect 298796 487228 298802 487240
rect 322198 487228 322204 487240
rect 322256 487228 322262 487280
rect 301958 487160 301964 487212
rect 302016 487200 302022 487212
rect 327718 487200 327724 487212
rect 302016 487172 327724 487200
rect 302016 487160 302022 487172
rect 327718 487160 327724 487172
rect 327776 487160 327782 487212
rect 289722 451188 289728 451240
rect 289780 451228 289786 451240
rect 289780 451200 292068 451228
rect 289780 451188 289786 451200
rect 302424 450226 302476 450232
rect 302424 450168 302476 450174
rect 305736 450226 305788 450232
rect 305736 450168 305788 450174
rect 295758 450143 295816 450149
rect 295758 450109 295770 450143
rect 295804 450140 295816 450143
rect 295886 450140 295892 450152
rect 295804 450112 295892 450140
rect 295804 450109 295816 450112
rect 295758 450103 295816 450109
rect 295886 450100 295892 450112
rect 295944 450100 295950 450152
rect 299075 450143 299133 450149
rect 299075 450109 299087 450143
rect 299121 450140 299133 450143
rect 299198 450140 299204 450152
rect 299121 450112 299204 450140
rect 299121 450109 299133 450112
rect 299075 450103 299133 450109
rect 299198 450100 299204 450112
rect 299256 450100 299262 450152
rect 309060 450140 309088 450200
rect 311250 450140 311256 450152
rect 309060 450112 311256 450140
rect 311250 450100 311256 450112
rect 311308 450100 311314 450152
rect 299198 447244 299204 447296
rect 299256 447284 299262 447296
rect 323578 447284 323584 447296
rect 299256 447256 323584 447284
rect 299256 447244 299262 447256
rect 323578 447244 323584 447256
rect 323636 447244 323642 447296
rect 302418 447176 302424 447228
rect 302476 447216 302482 447228
rect 329098 447216 329104 447228
rect 302476 447188 329104 447216
rect 302476 447176 302482 447188
rect 329098 447176 329104 447188
rect 329156 447176 329162 447228
rect 305730 447108 305736 447160
rect 305788 447148 305794 447160
rect 333238 447148 333244 447160
rect 305788 447120 333244 447148
rect 305788 447108 305794 447120
rect 333238 447108 333244 447120
rect 333296 447108 333302 447160
rect 289722 431196 289728 431248
rect 289780 431236 289786 431248
rect 289780 431208 292068 431236
rect 289780 431196 289786 431208
rect 292040 431206 292068 431208
rect 299290 430584 299296 430636
rect 299348 430633 299354 430636
rect 299348 430627 299388 430633
rect 299376 430593 299388 430627
rect 299348 430587 299388 430593
rect 299348 430584 299354 430587
rect 296622 430216 296628 430228
rect 295918 430188 296628 430216
rect 296622 430176 296628 430188
rect 296680 430176 296686 430228
rect 302792 430226 302844 430232
rect 302792 430168 302844 430174
rect 306196 430226 306248 430232
rect 306196 430168 306248 430174
rect 309704 430148 309732 430200
rect 312538 430148 312544 430160
rect 309704 430120 312544 430148
rect 312538 430108 312544 430120
rect 312596 430108 312602 430160
rect 299290 426504 299296 426556
rect 299348 426544 299354 426556
rect 324958 426544 324964 426556
rect 299348 426516 324964 426544
rect 299348 426504 299354 426516
rect 324958 426504 324964 426516
rect 325016 426504 325022 426556
rect 302786 426436 302792 426488
rect 302844 426476 302850 426488
rect 330478 426476 330484 426488
rect 302844 426448 330484 426476
rect 302844 426436 302850 426448
rect 330478 426436 330484 426448
rect 330536 426436 330542 426488
rect 296622 418072 296628 418124
rect 296680 418112 296686 418124
rect 517514 418112 517520 418124
rect 296680 418084 517520 418112
rect 296680 418072 296686 418084
rect 517514 418072 517520 418084
rect 517572 418072 517578 418124
rect 319438 413992 319444 414044
rect 319496 414032 319502 414044
rect 517514 414032 517520 414044
rect 319496 414004 517520 414032
rect 319496 413992 319502 414004
rect 517514 413992 517520 414004
rect 517572 413992 517578 414044
rect 320818 412632 320824 412684
rect 320876 412672 320882 412684
rect 517514 412672 517520 412684
rect 320876 412644 517520 412672
rect 320876 412632 320882 412644
rect 517514 412632 517520 412644
rect 517572 412632 517578 412684
rect 289722 411204 289728 411256
rect 289780 411244 289786 411256
rect 289780 411216 292068 411244
rect 289780 411204 289786 411216
rect 292040 411206 292068 411216
rect 298922 410592 298928 410644
rect 298980 410641 298986 410644
rect 298980 410635 299028 410641
rect 298980 410601 298982 410635
rect 299016 410601 299028 410635
rect 298980 410595 299028 410601
rect 298980 410592 298986 410595
rect 305454 410592 305460 410644
rect 305512 410641 305518 410644
rect 305512 410635 305558 410641
rect 305546 410601 305558 410635
rect 305512 410595 305558 410601
rect 305512 410592 305518 410595
rect 295708 410226 295760 410232
rect 295708 410168 295760 410174
rect 302240 410226 302292 410232
rect 311342 410224 311348 410236
rect 308784 410196 311348 410224
rect 311342 410184 311348 410196
rect 311400 410184 311406 410236
rect 302240 410168 302292 410174
rect 295702 408416 295708 408468
rect 295760 408456 295766 408468
rect 518158 408456 518164 408468
rect 295760 408428 518164 408456
rect 295760 408416 295766 408428
rect 518158 408416 518164 408428
rect 518216 408416 518222 408468
rect 298922 407532 298928 407584
rect 298980 407572 298986 407584
rect 298980 407544 306374 407572
rect 298980 407532 298986 407544
rect 302234 407464 302240 407516
rect 302292 407504 302298 407516
rect 302292 407476 305408 407504
rect 302292 407464 302298 407476
rect 305380 407300 305408 407476
rect 306346 407368 306374 407544
rect 326338 407368 326344 407380
rect 306346 407340 326344 407368
rect 326338 407328 326344 407340
rect 326396 407328 326402 407380
rect 331858 407300 331864 407312
rect 305380 407272 331864 407300
rect 331858 407260 331864 407272
rect 331916 407260 331922 407312
rect 305454 407192 305460 407244
rect 305512 407232 305518 407244
rect 334618 407232 334624 407244
rect 305512 407204 334624 407232
rect 305512 407192 305518 407204
rect 334618 407192 334624 407204
rect 334676 407192 334682 407244
rect 315298 407124 315304 407176
rect 315356 407164 315362 407176
rect 517514 407164 517520 407176
rect 315356 407136 517520 407164
rect 315356 407124 315362 407136
rect 517514 407124 517520 407136
rect 517572 407124 517578 407176
rect 316678 405696 316684 405748
rect 316736 405736 316742 405748
rect 517514 405736 517520 405748
rect 316736 405708 517520 405736
rect 316736 405696 316742 405708
rect 517514 405696 517520 405708
rect 517572 405696 517578 405748
rect 318058 401616 318064 401668
rect 318116 401656 318122 401668
rect 517514 401656 517520 401668
rect 318116 401628 517520 401656
rect 318116 401616 318122 401628
rect 517514 401616 517520 401628
rect 517572 401616 517578 401668
rect 289722 391212 289728 391264
rect 289780 391252 289786 391264
rect 289780 391224 292068 391252
rect 289780 391212 289786 391224
rect 292040 391206 292068 391224
rect 301596 391232 301648 391238
rect 301596 391174 301648 391180
rect 305368 391232 305420 391238
rect 309134 391180 309140 391232
rect 309192 391180 309198 391232
rect 305368 391174 305420 391180
rect 303614 390649 303620 390652
rect 303575 390643 303620 390649
rect 303575 390609 303587 390643
rect 303575 390603 303620 390609
rect 303614 390600 303620 390603
rect 303672 390600 303678 390652
rect 313918 390232 313924 390244
rect 296168 390226 296220 390232
rect 296168 390168 296220 390174
rect 299848 390226 299900 390232
rect 299848 390168 299900 390174
rect 307300 390226 307352 390232
rect 310992 390204 313924 390232
rect 310992 390200 311020 390204
rect 313918 390192 313924 390204
rect 313976 390192 313982 390244
rect 307300 390168 307352 390174
rect 296162 387744 296168 387796
rect 296220 387784 296226 387796
rect 319438 387784 319444 387796
rect 296220 387756 319444 387784
rect 296220 387744 296226 387756
rect 319438 387744 319444 387756
rect 319496 387744 319502 387796
rect 299842 386860 299848 386912
rect 299900 386900 299906 386912
rect 300762 386900 300768 386912
rect 299900 386872 300768 386900
rect 299900 386860 299906 386872
rect 300762 386860 300768 386872
rect 300820 386860 300826 386912
rect 322198 382168 322204 382220
rect 322256 382208 322262 382220
rect 517514 382208 517520 382220
rect 322256 382180 517520 382208
rect 322256 382168 322262 382180
rect 517514 382168 517520 382180
rect 517572 382168 517578 382220
rect 323578 379448 323584 379500
rect 323636 379488 323642 379500
rect 517514 379488 517520 379500
rect 323636 379460 517520 379488
rect 323636 379448 323642 379460
rect 517514 379448 517520 379460
rect 517572 379448 517578 379500
rect 324958 378088 324964 378140
rect 325016 378128 325022 378140
rect 517514 378128 517520 378140
rect 325016 378100 517520 378128
rect 325016 378088 325022 378100
rect 517514 378088 517520 378100
rect 517572 378088 517578 378140
rect 326338 376660 326344 376712
rect 326396 376700 326402 376712
rect 517514 376700 517520 376712
rect 326396 376672 517520 376700
rect 326396 376660 326402 376672
rect 517514 376660 517520 376672
rect 517572 376660 517578 376712
rect 300762 375300 300768 375352
rect 300820 375340 300826 375352
rect 517514 375340 517520 375352
rect 300820 375312 517520 375340
rect 300820 375300 300826 375312
rect 517514 375300 517520 375312
rect 517572 375300 517578 375352
rect 292040 371056 292068 371206
rect 289740 371028 292068 371056
rect 289740 370932 289768 371028
rect 289722 370880 289728 370932
rect 289780 370880 289786 370932
rect 307700 370651 307758 370657
rect 307700 370617 307712 370651
rect 307746 370648 307758 370651
rect 309778 370648 309784 370660
rect 307746 370620 309784 370648
rect 307746 370617 307758 370620
rect 307700 370611 307758 370617
rect 309778 370608 309784 370620
rect 309836 370608 309842 370660
rect 306852 370444 306880 370570
rect 306926 370444 306932 370456
rect 306852 370416 306932 370444
rect 306926 370404 306932 370416
rect 306984 370404 306990 370456
rect 295524 370226 295576 370232
rect 295524 370168 295576 370174
rect 298560 370226 298612 370232
rect 301774 370214 301780 370226
rect 301622 370186 301780 370214
rect 301774 370174 301780 370186
rect 301832 370174 301838 370226
rect 304810 370214 304816 370226
rect 304658 370186 304816 370214
rect 304810 370174 304816 370186
rect 304868 370174 304874 370226
rect 298560 370168 298612 370174
rect 295518 368432 295524 368484
rect 295576 368472 295582 368484
rect 295576 368444 296714 368472
rect 295576 368432 295582 368444
rect 296686 368404 296714 368444
rect 298554 368432 298560 368484
rect 298612 368472 298618 368484
rect 517514 368472 517520 368484
rect 298612 368444 517520 368472
rect 298612 368432 298618 368444
rect 517514 368432 517520 368444
rect 517572 368432 517578 368484
rect 320818 368404 320824 368416
rect 296686 368376 320824 368404
rect 320818 368364 320824 368376
rect 320876 368364 320882 368416
rect 319438 365712 319444 365764
rect 319496 365752 319502 365764
rect 517514 365752 517520 365764
rect 319496 365724 517520 365752
rect 319496 365712 319502 365724
rect 517514 365712 517520 365724
rect 517572 365712 517578 365764
rect 320818 364352 320824 364404
rect 320876 364392 320882 364404
rect 517514 364392 517520 364404
rect 320876 364364 517520 364392
rect 320876 364352 320882 364364
rect 517514 364352 517520 364364
rect 517572 364352 517578 364404
rect 322198 361564 322204 361616
rect 322256 361604 322262 361616
rect 517514 361604 517520 361616
rect 322256 361576 517520 361604
rect 322256 361564 322262 361576
rect 517514 361564 517520 361576
rect 517572 361564 517578 361616
rect 327718 342184 327724 342236
rect 327776 342224 327782 342236
rect 517514 342224 517520 342236
rect 327776 342196 517520 342224
rect 327776 342184 327782 342196
rect 517514 342184 517520 342196
rect 517572 342184 517578 342236
rect 329098 339396 329104 339448
rect 329156 339436 329162 339448
rect 517514 339436 517520 339448
rect 329156 339408 517520 339436
rect 329156 339396 329162 339408
rect 517514 339396 517520 339408
rect 517572 339396 517578 339448
rect 330478 338036 330484 338088
rect 330536 338076 330542 338088
rect 517514 338076 517520 338088
rect 330536 338048 517520 338076
rect 330536 338036 330542 338048
rect 517514 338036 517520 338048
rect 517572 338036 517578 338088
rect 331858 336676 331864 336728
rect 331916 336716 331922 336728
rect 517514 336716 517520 336728
rect 331916 336688 517520 336716
rect 331916 336676 331922 336688
rect 517514 336676 517520 336688
rect 517572 336676 517578 336728
rect 302142 333888 302148 333940
rect 302200 333928 302206 333940
rect 517514 333928 517520 333940
rect 302200 333900 517520 333928
rect 302200 333888 302206 333900
rect 517514 333888 517520 333900
rect 517572 333888 517578 333940
rect 323578 327088 323584 327140
rect 323636 327128 323642 327140
rect 517514 327128 517520 327140
rect 323636 327100 517520 327128
rect 323636 327088 323642 327100
rect 517514 327088 517520 327100
rect 517572 327088 517578 327140
rect 324958 325660 324964 325712
rect 325016 325700 325022 325712
rect 517514 325700 517520 325712
rect 325016 325672 517520 325700
rect 325016 325660 325022 325672
rect 517514 325660 517520 325672
rect 517572 325660 517578 325712
rect 326338 324300 326344 324352
rect 326396 324340 326402 324352
rect 517514 324340 517520 324352
rect 326396 324312 517520 324340
rect 326396 324300 326402 324312
rect 517514 324300 517520 324312
rect 517572 324300 517578 324352
rect 327718 321580 327724 321632
rect 327776 321620 327782 321632
rect 517514 321620 517520 321632
rect 327776 321592 517520 321620
rect 327776 321580 327782 321592
rect 517514 321580 517520 321592
rect 517572 321580 517578 321632
rect 333238 299412 333244 299464
rect 333296 299452 333302 299464
rect 517514 299452 517520 299464
rect 333296 299424 517520 299452
rect 333296 299412 333302 299424
rect 517514 299412 517520 299424
rect 517572 299412 517578 299464
rect 334618 296624 334624 296676
rect 334676 296664 334682 296676
rect 517514 296664 517520 296676
rect 334676 296636 517520 296664
rect 334676 296624 334682 296636
rect 517514 296624 517520 296636
rect 517572 296624 517578 296676
rect 304902 293904 304908 293956
rect 304960 293944 304966 293956
rect 517514 293944 517520 293956
rect 304960 293916 517520 293944
rect 304960 293904 304966 293916
rect 517514 293904 517520 293916
rect 517572 293904 517578 293956
rect 289722 291388 289728 291440
rect 289780 291428 289786 291440
rect 289780 291400 292160 291428
rect 289780 291388 289786 291400
rect 292132 291292 292160 291400
rect 292040 291264 292160 291292
rect 292040 291220 292068 291264
rect 292040 291192 292146 291220
rect 295800 290226 295852 290232
rect 305736 290226 305788 290232
rect 295800 290168 295852 290174
rect 299106 290164 299112 290216
rect 299164 290164 299170 290216
rect 302418 290164 302424 290216
rect 302476 290164 302482 290216
rect 305736 290168 305788 290174
rect 309060 290136 309088 290200
rect 311434 290136 311440 290148
rect 309060 290108 311440 290136
rect 311434 290096 311440 290108
rect 311492 290096 311498 290148
rect 302344 288408 302556 288436
rect 295794 288328 295800 288380
rect 295852 288368 295858 288380
rect 295852 288340 296714 288368
rect 295852 288328 295858 288340
rect 296686 288232 296714 288340
rect 299106 288328 299112 288380
rect 299164 288368 299170 288380
rect 302344 288368 302372 288408
rect 299164 288340 302372 288368
rect 299164 288328 299170 288340
rect 302418 288328 302424 288380
rect 302476 288328 302482 288380
rect 302528 288368 302556 288408
rect 518526 288368 518532 288380
rect 302528 288340 518532 288368
rect 518526 288328 518532 288340
rect 518584 288328 518590 288380
rect 302436 288300 302464 288328
rect 323578 288300 323584 288312
rect 302436 288272 323584 288300
rect 323578 288260 323584 288272
rect 323636 288260 323642 288312
rect 315298 288232 315304 288244
rect 296686 288204 315304 288232
rect 315298 288192 315304 288204
rect 315356 288192 315362 288244
rect 305730 287716 305736 287768
rect 305788 287756 305794 287768
rect 305788 287728 306374 287756
rect 305788 287716 305794 287728
rect 306346 287688 306374 287728
rect 517514 287688 517520 287700
rect 306346 287660 517520 287688
rect 517514 287648 517520 287660
rect 517572 287648 517578 287700
rect 329098 284316 329104 284368
rect 329156 284356 329162 284368
rect 517514 284356 517520 284368
rect 329156 284328 517520 284356
rect 329156 284316 329162 284328
rect 517514 284316 517520 284328
rect 517572 284316 517578 284368
rect 289722 271396 289728 271448
rect 289780 271436 289786 271448
rect 289780 271408 292068 271436
rect 289780 271396 289786 271408
rect 292040 271206 292068 271408
rect 299290 270580 299296 270632
rect 299348 270629 299354 270632
rect 299348 270623 299386 270629
rect 299374 270589 299386 270623
rect 299348 270583 299386 270589
rect 299348 270580 299354 270583
rect 295892 270226 295944 270232
rect 295892 270168 295944 270174
rect 302792 270226 302844 270232
rect 302792 270168 302844 270174
rect 306196 270226 306248 270232
rect 309718 270212 310008 270214
rect 312630 270212 312636 270224
rect 309718 270186 312636 270212
rect 309980 270184 312636 270186
rect 306196 270168 306248 270174
rect 312630 270172 312636 270184
rect 312688 270172 312694 270224
rect 306190 267656 306196 267708
rect 306248 267696 306254 267708
rect 518710 267696 518716 267708
rect 306248 267668 518716 267696
rect 306248 267656 306254 267668
rect 518710 267656 518716 267668
rect 518768 267656 518774 267708
rect 302786 267588 302792 267640
rect 302844 267628 302850 267640
rect 324958 267628 324964 267640
rect 302844 267600 324964 267628
rect 302844 267588 302850 267600
rect 324958 267588 324964 267600
rect 325016 267588 325022 267640
rect 299290 267520 299296 267572
rect 299348 267560 299354 267572
rect 319438 267560 319444 267572
rect 299348 267532 319444 267560
rect 299348 267520 299354 267532
rect 319438 267520 319444 267532
rect 319496 267520 319502 267572
rect 295886 267452 295892 267504
rect 295944 267492 295950 267504
rect 316678 267492 316684 267504
rect 295944 267464 316684 267492
rect 295944 267452 295950 267464
rect 316678 267452 316684 267464
rect 316736 267452 316742 267504
rect 311158 262148 311164 262200
rect 311216 262188 311222 262200
rect 517514 262188 517520 262200
rect 311216 262160 517520 262188
rect 311216 262148 311222 262160
rect 517514 262148 517520 262160
rect 517572 262148 517578 262200
rect 311250 259360 311256 259412
rect 311308 259400 311314 259412
rect 517514 259400 517520 259412
rect 311308 259372 517520 259400
rect 311308 259360 311314 259372
rect 517514 259360 517520 259372
rect 517572 259360 517578 259412
rect 312538 258000 312544 258052
rect 312596 258040 312602 258052
rect 517514 258040 517520 258052
rect 312596 258012 517520 258040
rect 312596 258000 312602 258012
rect 517514 258000 517520 258012
rect 517572 258000 517578 258052
rect 311342 256640 311348 256692
rect 311400 256680 311406 256692
rect 517514 256680 517520 256692
rect 311400 256652 517520 256680
rect 311400 256640 311406 256652
rect 517514 256640 517520 256652
rect 517572 256640 517578 256692
rect 313918 255212 313924 255264
rect 313976 255252 313982 255264
rect 517514 255252 517520 255264
rect 313976 255224 517520 255252
rect 313976 255212 313982 255224
rect 517514 255212 517520 255224
rect 517572 255212 517578 255264
rect 309778 253852 309784 253904
rect 309836 253892 309842 253904
rect 517514 253892 517520 253904
rect 309836 253864 517520 253892
rect 309836 253852 309842 253864
rect 517514 253852 517520 253864
rect 517572 253852 517578 253904
rect 289722 251404 289728 251456
rect 289780 251444 289786 251456
rect 289780 251416 292068 251444
rect 289780 251404 289786 251416
rect 292040 251206 292068 251416
rect 298646 251240 298652 251252
rect 298296 251220 298652 251240
rect 298218 251212 298652 251220
rect 298218 251192 298324 251212
rect 298646 251200 298652 251212
rect 298704 251200 298710 251252
rect 298922 250588 298928 250640
rect 298980 250637 298986 250640
rect 298980 250631 299027 250637
rect 298980 250597 298981 250631
rect 299015 250597 299027 250631
rect 298980 250591 299027 250597
rect 298980 250588 298986 250591
rect 305454 250588 305460 250640
rect 305512 250637 305518 250640
rect 305512 250631 305557 250637
rect 305545 250597 305557 250631
rect 305512 250591 305557 250597
rect 305512 250588 305518 250591
rect 295708 250226 295760 250232
rect 295708 250168 295760 250174
rect 302240 250226 302292 250232
rect 311802 250220 311808 250232
rect 308784 250192 311808 250220
rect 311802 250180 311808 250192
rect 311860 250180 311866 250232
rect 302240 250168 302292 250174
rect 298940 248424 299474 248452
rect 295702 248344 295708 248396
rect 295760 248384 295766 248396
rect 298940 248384 298968 248424
rect 295760 248356 298968 248384
rect 299446 248384 299474 248424
rect 518250 248384 518256 248396
rect 299446 248356 518256 248384
rect 295760 248344 295766 248356
rect 518250 248344 518256 248356
rect 518308 248344 518314 248396
rect 311434 248276 311440 248328
rect 311492 248316 311498 248328
rect 517514 248316 517520 248328
rect 311492 248288 517520 248316
rect 311492 248276 311498 248288
rect 517514 248276 517520 248288
rect 517572 248276 517578 248328
rect 302234 248208 302240 248260
rect 302292 248248 302298 248260
rect 326338 248248 326344 248260
rect 302292 248220 326344 248248
rect 302292 248208 302298 248220
rect 326338 248208 326344 248220
rect 326396 248208 326402 248260
rect 305454 248140 305460 248192
rect 305512 248180 305518 248192
rect 329098 248180 329104 248192
rect 305512 248152 329104 248180
rect 305512 248140 305518 248152
rect 329098 248140 329104 248152
rect 329156 248140 329162 248192
rect 298922 248072 298928 248124
rect 298980 248112 298986 248124
rect 320818 248112 320824 248124
rect 298980 248084 320824 248112
rect 298980 248072 298986 248084
rect 320818 248072 320824 248084
rect 320876 248072 320882 248124
rect 312630 246984 312636 247036
rect 312688 247024 312694 247036
rect 517514 247024 517520 247036
rect 312688 246996 517520 247024
rect 312688 246984 312694 246996
rect 517514 246984 517520 246996
rect 517572 246984 517578 247036
rect 311802 245556 311808 245608
rect 311860 245596 311866 245608
rect 517514 245596 517520 245608
rect 311860 245568 517520 245596
rect 311860 245556 311866 245568
rect 517514 245556 517520 245568
rect 517572 245556 517578 245608
rect 313918 242904 313924 242956
rect 313976 242944 313982 242956
rect 517514 242944 517520 242956
rect 313976 242916 517520 242944
rect 313976 242904 313982 242916
rect 517514 242904 517520 242916
rect 517572 242904 517578 242956
rect 289722 231412 289728 231464
rect 289780 231452 289786 231464
rect 289780 231424 292068 231452
rect 289780 231412 289786 231424
rect 292040 231207 292068 231424
rect 303614 230645 303620 230648
rect 303575 230639 303620 230645
rect 303575 230605 303587 230639
rect 303575 230599 303620 230605
rect 303614 230596 303620 230599
rect 303672 230596 303678 230648
rect 310992 230432 311020 230496
rect 313918 230432 313924 230444
rect 310992 230404 313924 230432
rect 313918 230392 313924 230404
rect 313976 230392 313982 230444
rect 296168 230226 296220 230232
rect 296168 230168 296220 230174
rect 299848 230226 299900 230232
rect 299848 230168 299900 230174
rect 307300 230226 307352 230232
rect 307300 230168 307352 230174
rect 296162 227672 296168 227724
rect 296220 227712 296226 227724
rect 518158 227712 518164 227724
rect 296220 227684 518164 227712
rect 296220 227672 296226 227684
rect 518158 227672 518164 227684
rect 518216 227672 518222 227724
rect 299842 227604 299848 227656
rect 299900 227644 299906 227656
rect 518342 227644 518348 227656
rect 299900 227616 518348 227644
rect 299900 227604 299906 227616
rect 518342 227604 518348 227616
rect 518400 227604 518406 227656
rect 303614 227536 303620 227588
rect 303672 227576 303678 227588
rect 518434 227576 518440 227588
rect 303672 227548 518440 227576
rect 303672 227536 303678 227548
rect 518434 227536 518440 227548
rect 518492 227536 518498 227588
rect 307294 227468 307300 227520
rect 307352 227508 307358 227520
rect 518618 227508 518624 227520
rect 307352 227480 518624 227508
rect 307352 227468 307358 227480
rect 518618 227468 518624 227480
rect 518676 227468 518682 227520
rect 580902 211868 580908 211880
rect 291948 211840 580908 211868
rect 291948 211664 291976 211840
rect 580902 211828 580908 211840
rect 580960 211828 580966 211880
rect 291948 211636 292068 211664
rect 289722 211352 289728 211404
rect 289780 211392 289786 211404
rect 292040 211392 292068 211636
rect 289780 211364 292068 211392
rect 289780 211352 289786 211364
rect 292040 211206 292068 211364
rect 295518 210653 295524 210656
rect 295491 210647 295524 210653
rect 295491 210613 295503 210647
rect 295491 210607 295524 210613
rect 295518 210604 295524 210607
rect 295576 210604 295582 210656
rect 307699 210647 307757 210653
rect 307699 210613 307711 210647
rect 307745 210644 307757 210647
rect 307745 210616 316034 210644
rect 307745 210613 307757 210616
rect 307699 210607 307757 210613
rect 298560 210226 298612 210232
rect 298560 210168 298612 210174
rect 301596 210226 301648 210232
rect 301596 210168 301648 210174
rect 304632 210226 304684 210232
rect 304632 210168 304684 210174
rect 316006 210168 316034 210616
rect 518250 210168 518256 210180
rect 316006 210140 518256 210168
rect 518250 210128 518256 210140
rect 518308 210128 518314 210180
rect 304626 208292 304632 208344
rect 304684 208332 304690 208344
rect 518526 208332 518532 208344
rect 304684 208304 518532 208332
rect 304684 208292 304690 208304
rect 518526 208292 518532 208304
rect 518584 208292 518590 208344
rect 301590 208224 301596 208276
rect 301648 208264 301654 208276
rect 327718 208264 327724 208276
rect 301648 208236 327724 208264
rect 301648 208224 301654 208236
rect 327718 208224 327724 208236
rect 327776 208224 327782 208276
rect 298554 208156 298560 208208
rect 298612 208196 298618 208208
rect 322198 208196 322204 208208
rect 298612 208168 322204 208196
rect 298612 208156 298618 208168
rect 322198 208156 322204 208168
rect 322256 208156 322262 208208
rect 295518 208088 295524 208140
rect 295576 208128 295582 208140
rect 318058 208128 318064 208140
rect 295576 208100 318064 208128
rect 295576 208088 295582 208100
rect 318058 208088 318064 208100
rect 318116 208088 318122 208140
<< via1 >>
rect 289728 490900 289780 490952
rect 301964 490603 302016 490612
rect 301964 490569 301968 490603
rect 301968 490569 302016 490603
rect 301964 490560 302016 490569
rect 295616 490176 295668 490228
rect 298744 490176 298796 490228
rect 305092 490176 305144 490228
rect 311164 490016 311216 490068
rect 298744 487228 298796 487280
rect 322204 487228 322256 487280
rect 301964 487160 302016 487212
rect 327724 487160 327776 487212
rect 289728 451188 289780 451240
rect 302424 450174 302476 450226
rect 305736 450174 305788 450226
rect 295892 450100 295944 450152
rect 299204 450100 299256 450152
rect 311256 450100 311308 450152
rect 299204 447244 299256 447296
rect 323584 447244 323636 447296
rect 302424 447176 302476 447228
rect 329104 447176 329156 447228
rect 305736 447108 305788 447160
rect 333244 447108 333296 447160
rect 289728 431196 289780 431248
rect 299296 430627 299348 430636
rect 299296 430593 299342 430627
rect 299342 430593 299348 430627
rect 299296 430584 299348 430593
rect 296628 430176 296680 430228
rect 302792 430174 302844 430226
rect 306196 430174 306248 430226
rect 312544 430108 312596 430160
rect 299296 426504 299348 426556
rect 324964 426504 325016 426556
rect 302792 426436 302844 426488
rect 330484 426436 330536 426488
rect 296628 418072 296680 418124
rect 517520 418072 517572 418124
rect 319444 413992 319496 414044
rect 517520 413992 517572 414044
rect 320824 412632 320876 412684
rect 517520 412632 517572 412684
rect 289728 411204 289780 411256
rect 298928 410592 298980 410644
rect 305460 410592 305512 410644
rect 295708 410174 295760 410226
rect 302240 410174 302292 410226
rect 311348 410184 311400 410236
rect 295708 408416 295760 408468
rect 518164 408416 518216 408468
rect 298928 407532 298980 407584
rect 302240 407464 302292 407516
rect 326344 407328 326396 407380
rect 331864 407260 331916 407312
rect 305460 407192 305512 407244
rect 334624 407192 334676 407244
rect 315304 407124 315356 407176
rect 517520 407124 517572 407176
rect 316684 405696 316736 405748
rect 517520 405696 517572 405748
rect 318064 401616 318116 401668
rect 517520 401616 517572 401668
rect 289728 391212 289780 391264
rect 301596 391180 301648 391232
rect 305368 391180 305420 391232
rect 309140 391180 309192 391232
rect 303620 390643 303672 390652
rect 303620 390609 303621 390643
rect 303621 390609 303672 390643
rect 303620 390600 303672 390609
rect 296168 390174 296220 390226
rect 299848 390174 299900 390226
rect 307300 390174 307352 390226
rect 313924 390192 313976 390244
rect 296168 387744 296220 387796
rect 319444 387744 319496 387796
rect 299848 386860 299900 386912
rect 300768 386860 300820 386912
rect 322204 382168 322256 382220
rect 517520 382168 517572 382220
rect 323584 379448 323636 379500
rect 517520 379448 517572 379500
rect 324964 378088 325016 378140
rect 517520 378088 517572 378140
rect 326344 376660 326396 376712
rect 517520 376660 517572 376712
rect 300768 375300 300820 375352
rect 517520 375300 517572 375352
rect 289728 370880 289780 370932
rect 309784 370608 309836 370660
rect 306932 370404 306984 370456
rect 295524 370174 295576 370226
rect 298560 370174 298612 370226
rect 301780 370174 301832 370226
rect 304816 370174 304868 370226
rect 295524 368432 295576 368484
rect 298560 368432 298612 368484
rect 517520 368432 517572 368484
rect 320824 368364 320876 368416
rect 319444 365712 319496 365764
rect 517520 365712 517572 365764
rect 320824 364352 320876 364404
rect 517520 364352 517572 364404
rect 322204 361564 322256 361616
rect 517520 361564 517572 361616
rect 327724 342184 327776 342236
rect 517520 342184 517572 342236
rect 329104 339396 329156 339448
rect 517520 339396 517572 339448
rect 330484 338036 330536 338088
rect 517520 338036 517572 338088
rect 331864 336676 331916 336728
rect 517520 336676 517572 336728
rect 302148 333888 302200 333940
rect 517520 333888 517572 333940
rect 323584 327088 323636 327140
rect 517520 327088 517572 327140
rect 324964 325660 325016 325712
rect 517520 325660 517572 325712
rect 326344 324300 326396 324352
rect 517520 324300 517572 324352
rect 327724 321580 327776 321632
rect 517520 321580 517572 321632
rect 333244 299412 333296 299464
rect 517520 299412 517572 299464
rect 334624 296624 334676 296676
rect 517520 296624 517572 296676
rect 304908 293904 304960 293956
rect 517520 293904 517572 293956
rect 289728 291388 289780 291440
rect 295800 290174 295852 290226
rect 299112 290164 299164 290216
rect 302424 290164 302476 290216
rect 305736 290174 305788 290226
rect 311440 290096 311492 290148
rect 295800 288328 295852 288380
rect 299112 288328 299164 288380
rect 302424 288328 302476 288380
rect 518532 288328 518584 288380
rect 323584 288260 323636 288312
rect 315304 288192 315356 288244
rect 305736 287716 305788 287768
rect 517520 287648 517572 287700
rect 329104 284316 329156 284368
rect 517520 284316 517572 284368
rect 289728 271396 289780 271448
rect 299296 270623 299348 270632
rect 299296 270589 299340 270623
rect 299340 270589 299348 270623
rect 299296 270580 299348 270589
rect 295892 270174 295944 270226
rect 302792 270174 302844 270226
rect 306196 270174 306248 270226
rect 312636 270172 312688 270224
rect 306196 267656 306248 267708
rect 518716 267656 518768 267708
rect 302792 267588 302844 267640
rect 324964 267588 325016 267640
rect 299296 267520 299348 267572
rect 319444 267520 319496 267572
rect 295892 267452 295944 267504
rect 316684 267452 316736 267504
rect 311164 262148 311216 262200
rect 517520 262148 517572 262200
rect 311256 259360 311308 259412
rect 517520 259360 517572 259412
rect 312544 258000 312596 258052
rect 517520 258000 517572 258052
rect 311348 256640 311400 256692
rect 517520 256640 517572 256692
rect 313924 255212 313976 255264
rect 517520 255212 517572 255264
rect 309784 253852 309836 253904
rect 517520 253852 517572 253904
rect 289728 251404 289780 251456
rect 298652 251200 298704 251252
rect 298928 250588 298980 250640
rect 305460 250631 305512 250640
rect 305460 250597 305511 250631
rect 305511 250597 305512 250631
rect 305460 250588 305512 250597
rect 295708 250174 295760 250226
rect 302240 250174 302292 250226
rect 311808 250180 311860 250232
rect 295708 248344 295760 248396
rect 518256 248344 518308 248396
rect 311440 248276 311492 248328
rect 517520 248276 517572 248328
rect 302240 248208 302292 248260
rect 326344 248208 326396 248260
rect 305460 248140 305512 248192
rect 329104 248140 329156 248192
rect 298928 248072 298980 248124
rect 320824 248072 320876 248124
rect 312636 246984 312688 247036
rect 517520 246984 517572 247036
rect 311808 245556 311860 245608
rect 517520 245556 517572 245608
rect 313924 242904 313976 242956
rect 517520 242904 517572 242956
rect 289728 231412 289780 231464
rect 303620 230639 303672 230648
rect 303620 230605 303621 230639
rect 303621 230605 303672 230639
rect 303620 230596 303672 230605
rect 313924 230392 313976 230444
rect 296168 230174 296220 230226
rect 299848 230174 299900 230226
rect 307300 230174 307352 230226
rect 296168 227672 296220 227724
rect 518164 227672 518216 227724
rect 299848 227604 299900 227656
rect 518348 227604 518400 227656
rect 303620 227536 303672 227588
rect 518440 227536 518492 227588
rect 307300 227468 307352 227520
rect 518624 227468 518676 227520
rect 580908 211828 580960 211880
rect 289728 211352 289780 211404
rect 295524 210647 295576 210656
rect 295524 210613 295537 210647
rect 295537 210613 295576 210647
rect 295524 210604 295576 210613
rect 298560 210174 298612 210226
rect 301596 210174 301648 210226
rect 304632 210174 304684 210226
rect 518256 210128 518308 210180
rect 304632 208292 304684 208344
rect 518532 208292 518584 208344
rect 301596 208224 301648 208276
rect 327724 208224 327776 208276
rect 298560 208156 298612 208208
rect 322204 208156 322256 208208
rect 295524 208088 295576 208140
rect 318064 208088 318116 208140
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 289728 490952 289780 490958
rect 289728 490894 289780 490900
rect 289740 451246 289768 490894
rect 294769 490592 294778 490648
rect 294834 490592 294843 490648
rect 297925 490592 297934 490648
rect 297990 490592 297999 490648
rect 301080 490592 301089 490648
rect 301145 490592 301154 490648
rect 301964 490612 302016 490618
rect 304237 490592 304246 490648
rect 304302 490592 304311 490648
rect 301964 490554 302016 490560
rect 295616 490228 295668 490234
rect 295616 490170 295668 490176
rect 298744 490228 298796 490234
rect 298744 490170 298796 490176
rect 295628 487257 295656 490170
rect 298756 487286 298784 490170
rect 298744 487280 298796 487286
rect 295614 487248 295670 487257
rect 298744 487222 298796 487228
rect 301976 487218 302004 490554
rect 307417 490385 307445 490620
rect 307403 490376 307459 490385
rect 307403 490311 307459 490320
rect 305092 490228 305144 490234
rect 305092 490170 305144 490176
rect 305104 487257 305132 490170
rect 311164 490068 311216 490074
rect 311164 490010 311216 490016
rect 305090 487248 305146 487257
rect 295614 487183 295670 487192
rect 301964 487212 302016 487218
rect 305090 487183 305146 487192
rect 301964 487154 302016 487160
rect 289728 451240 289780 451246
rect 289728 451182 289780 451188
rect 289740 431254 289768 451182
rect 294524 451166 294954 451194
rect 294524 450945 294552 451166
rect 301551 451152 301560 451208
rect 301616 451152 301625 451208
rect 304868 451152 304877 451208
rect 304933 451152 304942 451208
rect 307772 451166 308221 451194
rect 307772 450945 307800 451166
rect 294510 450936 294566 450945
rect 294510 450871 294566 450880
rect 307758 450936 307814 450945
rect 307758 450871 307814 450880
rect 298257 450537 298285 450772
rect 298257 450528 298338 450537
rect 298257 450486 298282 450528
rect 298282 450463 298338 450472
rect 302424 450226 302476 450232
rect 302424 450168 302476 450174
rect 305736 450226 305788 450232
rect 305736 450168 305788 450174
rect 295892 450152 295944 450158
rect 295892 450094 295944 450100
rect 299204 450152 299256 450158
rect 299204 450094 299256 450100
rect 295904 447273 295932 450094
rect 299216 447302 299244 450094
rect 299204 447296 299256 447302
rect 295890 447264 295946 447273
rect 299204 447238 299256 447244
rect 302436 447234 302464 450168
rect 295890 447199 295946 447208
rect 302424 447228 302476 447234
rect 302424 447170 302476 447176
rect 305748 447166 305776 450168
rect 305736 447160 305788 447166
rect 305736 447102 305788 447108
rect 289728 431248 289780 431254
rect 289728 431190 289780 431196
rect 298190 431216 298246 431225
rect 289740 411262 289768 431190
rect 298246 431174 298526 431202
rect 298190 431151 298246 431160
rect 294694 431080 294750 431089
rect 301594 431080 301650 431089
rect 294750 431038 295082 431066
rect 294694 431015 294750 431024
rect 301650 431038 301970 431066
rect 301594 431015 301650 431024
rect 308402 430944 308458 430953
rect 305288 430902 305414 430930
rect 305288 430794 305316 430902
rect 308458 430902 308858 430930
rect 308402 430879 308458 430888
rect 305104 430766 305316 430794
rect 304998 430672 305054 430681
rect 299296 430636 299348 430642
rect 305104 430658 305132 430766
rect 305054 430630 305132 430658
rect 304998 430607 305054 430616
rect 299296 430578 299348 430584
rect 296628 430228 296680 430234
rect 296628 430170 296680 430176
rect 296640 418130 296668 430170
rect 299308 426562 299336 430578
rect 302792 430226 302844 430232
rect 302792 430168 302844 430174
rect 306196 430226 306248 430232
rect 306196 430168 306248 430174
rect 299296 426556 299348 426562
rect 299296 426498 299348 426504
rect 302804 426494 302832 430168
rect 302792 426488 302844 426494
rect 306208 426465 306236 430168
rect 302792 426430 302844 426436
rect 306194 426456 306250 426465
rect 306194 426391 306250 426400
rect 296628 418124 296680 418130
rect 296628 418066 296680 418072
rect 298190 411360 298246 411369
rect 298112 411318 298190 411346
rect 289728 411256 289780 411262
rect 289728 411198 289780 411204
rect 298112 411210 298140 411318
rect 298190 411295 298246 411304
rect 289740 391270 289768 411198
rect 298112 411182 298168 411210
rect 294889 410394 294917 410652
rect 298928 410644 298980 410650
rect 298928 410586 298980 410592
rect 294889 410366 294920 410394
rect 294892 410122 294920 410366
rect 295708 410226 295760 410232
rect 295708 410168 295760 410174
rect 295154 410136 295210 410145
rect 294892 410094 295154 410122
rect 295154 410071 295210 410080
rect 295720 408474 295748 410168
rect 295708 408468 295760 408474
rect 295708 408410 295760 408416
rect 298940 407590 298968 410586
rect 301419 410394 301447 410652
rect 304684 410394 304712 410652
rect 305460 410644 305512 410650
rect 305460 410586 305512 410592
rect 301419 410366 301452 410394
rect 304684 410366 304764 410394
rect 301424 410122 301452 410366
rect 302240 410226 302292 410232
rect 302240 410168 302292 410174
rect 301594 410136 301650 410145
rect 301424 410094 301594 410122
rect 301594 410071 301650 410080
rect 298928 407584 298980 407590
rect 298928 407526 298980 407532
rect 302252 407522 302280 410168
rect 304736 410145 304764 410366
rect 304722 410136 304778 410145
rect 304722 410071 304778 410080
rect 302240 407516 302292 407522
rect 302240 407458 302292 407464
rect 305472 407250 305500 410586
rect 307949 410394 307977 410652
rect 307949 410366 307984 410394
rect 307956 410122 307984 410366
rect 308218 410136 308274 410145
rect 307956 410094 308218 410122
rect 308218 410071 308274 410080
rect 305460 407244 305512 407250
rect 305460 407186 305512 407192
rect 295338 391504 295394 391513
rect 299202 391504 299258 391513
rect 295338 391439 295394 391448
rect 299047 391462 299202 391490
rect 289728 391264 289780 391270
rect 289728 391206 289780 391212
rect 289740 370938 289768 391206
rect 295352 391204 295380 391439
rect 298190 391232 298246 391241
rect 299047 391218 299075 391462
rect 299202 391439 299258 391448
rect 298246 391204 299075 391218
rect 301594 391232 301650 391241
rect 298246 391190 299061 391204
rect 298190 391167 298246 391176
rect 301594 391167 301650 391176
rect 305368 391232 305420 391238
rect 305368 391174 305420 391180
rect 309140 391232 309192 391238
rect 309140 391174 309192 391180
rect 305380 391105 305408 391174
rect 309152 391105 309180 391174
rect 305366 391096 305422 391105
rect 305366 391031 305422 391040
rect 309138 391096 309194 391105
rect 309138 391031 309194 391040
rect 303620 390652 303672 390658
rect 303620 390594 303672 390600
rect 296168 390226 296220 390232
rect 296168 390168 296220 390174
rect 299848 390226 299900 390232
rect 299848 390168 299900 390174
rect 296180 387802 296208 390168
rect 296168 387796 296220 387802
rect 296168 387738 296220 387744
rect 299860 386918 299888 390168
rect 299848 386912 299900 386918
rect 299848 386854 299900 386860
rect 300768 386912 300820 386918
rect 303632 386889 303660 390594
rect 307300 390226 307352 390232
rect 307300 390168 307352 390174
rect 307312 386889 307340 390168
rect 300768 386854 300820 386860
rect 303618 386880 303674 386889
rect 300780 375358 300808 386854
rect 303618 386815 303674 386824
rect 307298 386880 307354 386889
rect 307298 386815 307354 386824
rect 300768 375352 300820 375358
rect 300768 375294 300820 375300
rect 289728 370932 289780 370938
rect 289728 370874 289780 370880
rect 289740 291446 289768 370874
rect 294676 370410 294704 370668
rect 297728 370546 297756 370668
rect 297728 370518 297772 370546
rect 294616 370382 294704 370410
rect 294510 370016 294566 370025
rect 294616 370002 294644 370382
rect 295524 370226 295576 370232
rect 295524 370168 295576 370174
rect 294566 369974 294644 370002
rect 294510 369951 294566 369960
rect 295536 368490 295564 370168
rect 297744 370002 297772 370518
rect 298560 370226 298612 370232
rect 298560 370168 298612 370174
rect 298006 370016 298062 370025
rect 297744 369974 298006 370002
rect 298006 369951 298062 369960
rect 298572 368490 298600 370168
rect 300780 370025 300808 370668
rect 303832 370410 303860 370668
rect 309784 370660 309836 370666
rect 309784 370602 309836 370608
rect 306932 370456 306984 370462
rect 303832 370382 303936 370410
rect 306932 370398 306984 370404
rect 301780 370226 301832 370232
rect 301780 370168 301832 370174
rect 300766 370016 300822 370025
rect 300766 369951 300822 369960
rect 295524 368484 295576 368490
rect 295524 368426 295576 368432
rect 298560 368484 298612 368490
rect 298560 368426 298612 368432
rect 301792 364334 301820 370168
rect 303908 370002 303936 370382
rect 304816 370226 304868 370232
rect 304816 370168 304868 370174
rect 304170 370016 304226 370025
rect 303908 369974 304170 370002
rect 304170 369951 304226 369960
rect 304828 364334 304856 370168
rect 306944 370025 306972 370398
rect 306930 370016 306986 370025
rect 306930 369951 306986 369960
rect 301792 364306 302188 364334
rect 304828 364306 304948 364334
rect 302160 333946 302188 364306
rect 302148 333940 302200 333946
rect 302148 333882 302200 333888
rect 304920 293962 304948 364306
rect 304908 293956 304960 293962
rect 304908 293898 304960 293904
rect 304899 291488 304908 291544
rect 304964 291488 304973 291544
rect 289728 291440 289780 291446
rect 300122 291408 300178 291417
rect 289728 291382 289780 291388
rect 289740 271454 289768 291382
rect 299837 291366 300122 291394
rect 306746 291408 306802 291417
rect 306470 291366 306746 291394
rect 300122 291343 300178 291352
rect 306746 291343 306802 291352
rect 294602 291272 294658 291281
rect 298098 291272 298154 291281
rect 294658 291230 294985 291258
rect 294602 291207 294658 291216
rect 298154 291230 298302 291258
rect 298098 291207 298154 291216
rect 295800 290226 295852 290232
rect 305736 290226 305788 290232
rect 295800 290168 295852 290174
rect 299112 290216 299164 290222
rect 295812 288386 295840 290168
rect 299112 290158 299164 290164
rect 302424 290216 302476 290222
rect 305736 290168 305788 290174
rect 302424 290158 302476 290164
rect 299124 288386 299152 290158
rect 302436 288386 302464 290158
rect 295800 288380 295852 288386
rect 295800 288322 295852 288328
rect 299112 288380 299164 288386
rect 299112 288322 299164 288328
rect 302424 288380 302476 288386
rect 302424 288322 302476 288328
rect 305748 287774 305776 290168
rect 305736 287768 305788 287774
rect 305736 287710 305788 287716
rect 294685 271496 294694 271552
rect 294750 271496 294759 271552
rect 298489 271496 298498 271552
rect 298554 271496 298563 271552
rect 301401 271496 301410 271552
rect 301466 271496 301475 271552
rect 304989 271496 304998 271552
rect 305054 271496 305063 271552
rect 308301 271496 308310 271552
rect 308366 271496 308375 271552
rect 289728 271448 289780 271454
rect 289728 271390 289780 271396
rect 289740 251462 289768 271390
rect 299296 270632 299348 270638
rect 299296 270574 299348 270580
rect 295892 270226 295944 270232
rect 295892 270168 295944 270174
rect 295904 267510 295932 270168
rect 299308 267578 299336 270574
rect 302792 270226 302844 270232
rect 302792 270168 302844 270174
rect 306196 270226 306248 270232
rect 306196 270168 306248 270174
rect 302804 267646 302832 270168
rect 306208 267714 306236 270168
rect 306196 267708 306248 267714
rect 306196 267650 306248 267656
rect 302792 267640 302844 267646
rect 302792 267582 302844 267588
rect 299296 267572 299348 267578
rect 299296 267514 299348 267520
rect 295892 267504 295944 267510
rect 295892 267446 295944 267452
rect 309796 253910 309824 370602
rect 311176 262206 311204 490010
rect 322204 487280 322256 487286
rect 322204 487222 322256 487228
rect 311256 450152 311308 450158
rect 311256 450094 311308 450100
rect 311164 262200 311216 262206
rect 311164 262142 311216 262148
rect 311268 259418 311296 450094
rect 312544 430160 312596 430166
rect 312544 430102 312596 430108
rect 311348 410236 311400 410242
rect 311348 410178 311400 410184
rect 311256 259412 311308 259418
rect 311256 259354 311308 259360
rect 311360 256698 311388 410178
rect 311440 290148 311492 290154
rect 311440 290090 311492 290096
rect 311348 256692 311400 256698
rect 311348 256634 311400 256640
rect 309784 253904 309836 253910
rect 309784 253846 309836 253852
rect 298650 251560 298706 251569
rect 301410 251560 301466 251569
rect 298650 251495 298706 251504
rect 301332 251518 301410 251546
rect 289728 251456 289780 251462
rect 289728 251398 289780 251404
rect 294878 251424 294934 251433
rect 289740 231470 289768 251398
rect 294878 251359 294934 251368
rect 294888 251124 294916 251359
rect 298664 251258 298692 251495
rect 298652 251252 298704 251258
rect 298652 251194 298704 251200
rect 301332 251138 301360 251518
rect 308218 251560 308274 251569
rect 301410 251495 301466 251504
rect 307864 251518 308218 251546
rect 307864 251138 307892 251518
rect 308218 251495 308274 251504
rect 308954 251560 309010 251569
rect 309010 251518 309180 251546
rect 308954 251495 309010 251504
rect 301332 251110 301432 251138
rect 307864 251110 307962 251138
rect 304669 251016 304725 251025
rect 304669 250951 304725 250960
rect 298928 250640 298980 250646
rect 298928 250582 298980 250588
rect 305460 250640 305512 250646
rect 305460 250582 305512 250588
rect 295708 250226 295760 250232
rect 295708 250168 295760 250174
rect 295720 248402 295748 250168
rect 295708 248396 295760 248402
rect 295708 248338 295760 248344
rect 298940 248130 298968 250582
rect 302240 250226 302292 250232
rect 302240 250168 302292 250174
rect 302252 248266 302280 250168
rect 302240 248260 302292 248266
rect 302240 248202 302292 248208
rect 305472 248198 305500 250582
rect 305460 248192 305512 248198
rect 305460 248134 305512 248140
rect 298928 248124 298980 248130
rect 298928 248066 298980 248072
rect 309152 233345 309180 251518
rect 311452 248334 311480 290090
rect 312556 258058 312584 430102
rect 319444 414044 319496 414050
rect 319444 413986 319496 413992
rect 315304 407176 315356 407182
rect 315304 407118 315356 407124
rect 313924 390244 313976 390250
rect 313924 390186 313976 390192
rect 312636 270224 312688 270230
rect 312636 270166 312688 270172
rect 312544 258052 312596 258058
rect 312544 257994 312596 258000
rect 311808 250232 311860 250238
rect 311808 250174 311860 250180
rect 311440 248328 311492 248334
rect 311440 248270 311492 248276
rect 311820 245614 311848 250174
rect 312648 247042 312676 270166
rect 313936 255270 313964 390186
rect 315316 288250 315344 407118
rect 316684 405748 316736 405754
rect 316684 405690 316736 405696
rect 315304 288244 315356 288250
rect 315304 288186 315356 288192
rect 316696 267510 316724 405690
rect 318064 401668 318116 401674
rect 318064 401610 318116 401616
rect 316684 267504 316736 267510
rect 316684 267446 316736 267452
rect 313924 255264 313976 255270
rect 313924 255206 313976 255212
rect 312636 247036 312688 247042
rect 312636 246978 312688 246984
rect 311808 245608 311860 245614
rect 311808 245550 311860 245556
rect 313924 242956 313976 242962
rect 313924 242898 313976 242904
rect 309138 233336 309194 233345
rect 309138 233271 309194 233280
rect 289728 231464 289780 231470
rect 295338 231432 295394 231441
rect 289728 231406 289780 231412
rect 289740 211410 289768 231406
rect 295335 231376 295338 231418
rect 295335 231367 295394 231376
rect 299033 231432 299089 231441
rect 299033 231367 299089 231376
rect 295335 231132 295363 231367
rect 299047 231010 299075 231367
rect 299032 230996 299075 231010
rect 299032 230982 299061 230996
rect 296168 230226 296220 230232
rect 299032 230217 299060 230982
rect 303620 230648 303672 230654
rect 302745 230616 302801 230625
rect 303620 230590 303672 230596
rect 306457 230616 306513 230625
rect 302745 230551 302801 230560
rect 299848 230226 299900 230232
rect 296168 230168 296220 230174
rect 299018 230208 299074 230217
rect 296180 227730 296208 230168
rect 299848 230168 299900 230174
rect 299018 230143 299074 230152
rect 296168 227724 296220 227730
rect 296168 227666 296220 227672
rect 299860 227662 299888 230168
rect 299848 227656 299900 227662
rect 299848 227598 299900 227604
rect 303632 227594 303660 230590
rect 306457 230551 306513 230560
rect 310150 230616 310206 230625
rect 310150 230551 310206 230560
rect 313936 230450 313964 242898
rect 313924 230444 313976 230450
rect 313924 230386 313976 230392
rect 307300 230226 307352 230232
rect 307300 230168 307352 230174
rect 303620 227588 303672 227594
rect 303620 227530 303672 227536
rect 307312 227526 307340 230168
rect 307300 227520 307352 227526
rect 307300 227462 307352 227468
rect 307022 213344 307078 213353
rect 307022 213279 307078 213288
rect 303894 213208 303950 213217
rect 303894 213143 303950 213152
rect 303908 211857 303936 213143
rect 307036 211857 307064 213279
rect 303894 211848 303950 211857
rect 303894 211783 303950 211792
rect 307022 211848 307078 211857
rect 307022 211783 307078 211792
rect 306930 211576 306986 211585
rect 306930 211511 306986 211520
rect 303817 211440 303873 211449
rect 289728 211404 289780 211410
rect 306944 211426 306972 211511
rect 303817 211375 303873 211384
rect 306883 211398 306972 211426
rect 289728 211346 289780 211352
rect 300765 211168 300821 211177
rect 303831 211140 303859 211375
rect 306883 211140 306911 211398
rect 300765 211103 300821 211112
rect 295524 210656 295576 210662
rect 295524 210598 295576 210604
rect 294708 210497 294736 210596
rect 294694 210488 294750 210497
rect 294694 210423 294750 210432
rect 295536 208146 295564 210598
rect 297744 210497 297772 210596
rect 297730 210488 297786 210497
rect 297730 210423 297786 210432
rect 298560 210226 298612 210232
rect 298560 210168 298612 210174
rect 301596 210226 301648 210232
rect 301596 210168 301648 210174
rect 304632 210226 304684 210232
rect 304632 210168 304684 210174
rect 298572 208214 298600 210168
rect 301608 208282 301636 210168
rect 304644 208350 304672 210168
rect 304632 208344 304684 208350
rect 304632 208286 304684 208292
rect 301596 208276 301648 208282
rect 301596 208218 301648 208224
rect 298560 208208 298612 208214
rect 298560 208150 298612 208156
rect 318076 208146 318104 401610
rect 319456 387802 319484 413986
rect 320824 412684 320876 412690
rect 320824 412626 320876 412632
rect 319444 387796 319496 387802
rect 319444 387738 319496 387744
rect 320836 368422 320864 412626
rect 322216 382226 322244 487222
rect 327724 487212 327776 487218
rect 327724 487154 327776 487160
rect 323584 447296 323636 447302
rect 323584 447238 323636 447244
rect 322204 382220 322256 382226
rect 322204 382162 322256 382168
rect 323596 379506 323624 447238
rect 324964 426556 325016 426562
rect 324964 426498 325016 426504
rect 323584 379500 323636 379506
rect 323584 379442 323636 379448
rect 324976 378146 325004 426498
rect 326344 407380 326396 407386
rect 326344 407322 326396 407328
rect 324964 378140 325016 378146
rect 324964 378082 325016 378088
rect 326356 376718 326384 407322
rect 326344 376712 326396 376718
rect 326344 376654 326396 376660
rect 320824 368416 320876 368422
rect 320824 368358 320876 368364
rect 319444 365764 319496 365770
rect 319444 365706 319496 365712
rect 319456 267578 319484 365706
rect 320824 364404 320876 364410
rect 320824 364346 320876 364352
rect 319444 267572 319496 267578
rect 319444 267514 319496 267520
rect 320836 248130 320864 364346
rect 322204 361616 322256 361622
rect 322204 361558 322256 361564
rect 320824 248124 320876 248130
rect 320824 248066 320876 248072
rect 322216 208214 322244 361558
rect 327736 342242 327764 487154
rect 329104 447228 329156 447234
rect 329104 447170 329156 447176
rect 327724 342236 327776 342242
rect 327724 342178 327776 342184
rect 329116 339454 329144 447170
rect 333244 447160 333296 447166
rect 333244 447102 333296 447108
rect 330484 426488 330536 426494
rect 330484 426430 330536 426436
rect 329104 339448 329156 339454
rect 329104 339390 329156 339396
rect 330496 338094 330524 426430
rect 331864 407312 331916 407318
rect 331864 407254 331916 407260
rect 330484 338088 330536 338094
rect 330484 338030 330536 338036
rect 331876 336734 331904 407254
rect 331864 336728 331916 336734
rect 331864 336670 331916 336676
rect 323584 327140 323636 327146
rect 323584 327082 323636 327088
rect 323596 288318 323624 327082
rect 324964 325712 325016 325718
rect 324964 325654 325016 325660
rect 323584 288312 323636 288318
rect 323584 288254 323636 288260
rect 324976 267646 325004 325654
rect 326344 324352 326396 324358
rect 326344 324294 326396 324300
rect 324964 267640 325016 267646
rect 324964 267582 325016 267588
rect 326356 248266 326384 324294
rect 327724 321632 327776 321638
rect 327724 321574 327776 321580
rect 326344 248260 326396 248266
rect 326344 248202 326396 248208
rect 327736 208282 327764 321574
rect 333256 299470 333284 447102
rect 520660 421382 521226 421410
rect 528678 421382 529336 421410
rect 517520 418124 517572 418130
rect 517520 418066 517572 418072
rect 517532 416945 517560 418066
rect 517518 416936 517574 416945
rect 517518 416871 517574 416880
rect 518162 415576 518218 415585
rect 518162 415511 518218 415520
rect 517518 414216 517574 414225
rect 517518 414151 517574 414160
rect 517532 414050 517560 414151
rect 517520 414044 517572 414050
rect 517520 413986 517572 413992
rect 517518 412856 517574 412865
rect 517518 412791 517574 412800
rect 517532 412690 517560 412791
rect 517520 412684 517572 412690
rect 517520 412626 517572 412632
rect 518176 408474 518204 415511
rect 518164 408468 518216 408474
rect 518164 408410 518216 408416
rect 517518 407416 517574 407425
rect 517518 407351 517574 407360
rect 334624 407244 334676 407250
rect 334624 407186 334676 407192
rect 333244 299464 333296 299470
rect 333244 299406 333296 299412
rect 334636 296682 334664 407186
rect 517532 407182 517560 407351
rect 517520 407176 517572 407182
rect 517520 407118 517572 407124
rect 517518 406056 517574 406065
rect 517518 405991 517574 406000
rect 517532 405754 517560 405991
rect 517520 405748 517572 405754
rect 517520 405690 517572 405696
rect 518254 404696 518310 404705
rect 518254 404631 518310 404640
rect 518162 403336 518218 403345
rect 518162 403271 518218 403280
rect 517518 401976 517574 401985
rect 517518 401911 517574 401920
rect 517532 401674 517560 401911
rect 517520 401668 517572 401674
rect 517520 401610 517572 401616
rect 517520 382220 517572 382226
rect 517520 382162 517572 382168
rect 517532 381041 517560 382162
rect 517518 381032 517574 381041
rect 517518 380967 517574 380976
rect 517520 379500 517572 379506
rect 517520 379442 517572 379448
rect 517532 378321 517560 379442
rect 517518 378312 517574 378321
rect 517518 378247 517574 378256
rect 517520 378140 517572 378146
rect 517520 378082 517572 378088
rect 517532 376961 517560 378082
rect 517518 376952 517574 376961
rect 517518 376887 517574 376896
rect 517520 376712 517572 376718
rect 517520 376654 517572 376660
rect 517532 375601 517560 376654
rect 517518 375592 517574 375601
rect 517518 375527 517574 375536
rect 517520 375352 517572 375358
rect 517520 375294 517572 375300
rect 517532 374241 517560 375294
rect 517518 374232 517574 374241
rect 517518 374167 517574 374176
rect 517518 372872 517574 372881
rect 517518 372807 517574 372816
rect 517532 368490 517560 372807
rect 517520 368484 517572 368490
rect 517520 368426 517572 368432
rect 517518 366072 517574 366081
rect 517518 366007 517574 366016
rect 517532 365770 517560 366007
rect 517520 365764 517572 365770
rect 517520 365706 517572 365712
rect 517518 364712 517574 364721
rect 517518 364647 517574 364656
rect 517532 364410 517560 364647
rect 517520 364404 517572 364410
rect 517520 364346 517572 364352
rect 517518 361992 517574 362001
rect 517518 361927 517574 361936
rect 517532 361622 517560 361927
rect 517520 361616 517572 361622
rect 517520 361558 517572 361564
rect 517520 342236 517572 342242
rect 517520 342178 517572 342184
rect 517532 341057 517560 342178
rect 517518 341048 517574 341057
rect 517518 340983 517574 340992
rect 517520 339448 517572 339454
rect 517520 339390 517572 339396
rect 517532 338337 517560 339390
rect 517518 338328 517574 338337
rect 517518 338263 517574 338272
rect 517520 338088 517572 338094
rect 517520 338030 517572 338036
rect 517532 336977 517560 338030
rect 517518 336968 517574 336977
rect 517518 336903 517574 336912
rect 517520 336728 517572 336734
rect 517520 336670 517572 336676
rect 517532 335617 517560 336670
rect 517518 335608 517574 335617
rect 517518 335543 517574 335552
rect 517520 333940 517572 333946
rect 517520 333882 517572 333888
rect 517532 332897 517560 333882
rect 517518 332888 517574 332897
rect 517518 332823 517574 332832
rect 517518 327448 517574 327457
rect 517518 327383 517574 327392
rect 517532 327146 517560 327383
rect 517520 327140 517572 327146
rect 517520 327082 517572 327088
rect 517518 326088 517574 326097
rect 517518 326023 517574 326032
rect 517532 325718 517560 326023
rect 517520 325712 517572 325718
rect 517520 325654 517572 325660
rect 517518 324728 517574 324737
rect 517518 324663 517574 324672
rect 517532 324358 517560 324663
rect 517520 324352 517572 324358
rect 517520 324294 517572 324300
rect 517518 322008 517574 322017
rect 517518 321943 517574 321952
rect 517532 321638 517560 321943
rect 517520 321632 517572 321638
rect 517520 321574 517572 321580
rect 517520 299464 517572 299470
rect 517520 299406 517572 299412
rect 517532 298353 517560 299406
rect 517518 298344 517574 298353
rect 517518 298279 517574 298288
rect 334624 296676 334676 296682
rect 334624 296618 334676 296624
rect 517520 296676 517572 296682
rect 517520 296618 517572 296624
rect 517532 295633 517560 296618
rect 517518 295624 517574 295633
rect 517518 295559 517574 295568
rect 517520 293956 517572 293962
rect 517520 293898 517572 293904
rect 517532 292913 517560 293898
rect 517518 292904 517574 292913
rect 517518 292839 517574 292848
rect 517520 287700 517572 287706
rect 517520 287642 517572 287648
rect 517532 287473 517560 287642
rect 517518 287464 517574 287473
rect 517518 287399 517574 287408
rect 517518 284744 517574 284753
rect 517518 284679 517574 284688
rect 517532 284374 517560 284679
rect 329104 284368 329156 284374
rect 329104 284310 329156 284316
rect 517520 284368 517572 284374
rect 517520 284310 517572 284316
rect 329116 248198 329144 284310
rect 517520 262200 517572 262206
rect 517520 262142 517572 262148
rect 517532 261089 517560 262142
rect 517518 261080 517574 261089
rect 517518 261015 517574 261024
rect 517520 259412 517572 259418
rect 517520 259354 517572 259360
rect 517532 258369 517560 259354
rect 517518 258360 517574 258369
rect 517518 258295 517574 258304
rect 517520 258052 517572 258058
rect 517520 257994 517572 258000
rect 517532 257009 517560 257994
rect 517518 257000 517574 257009
rect 517518 256935 517574 256944
rect 517520 256692 517572 256698
rect 517520 256634 517572 256640
rect 517532 255649 517560 256634
rect 517518 255640 517574 255649
rect 517518 255575 517574 255584
rect 517520 255264 517572 255270
rect 517520 255206 517572 255212
rect 517532 254289 517560 255206
rect 517518 254280 517574 254289
rect 517518 254215 517574 254224
rect 517520 253904 517572 253910
rect 517520 253846 517572 253852
rect 517532 252929 517560 253846
rect 517518 252920 517574 252929
rect 517518 252855 517574 252864
rect 517520 248328 517572 248334
rect 517520 248270 517572 248276
rect 329104 248192 329156 248198
rect 329104 248134 329156 248140
rect 517532 247489 517560 248270
rect 517518 247480 517574 247489
rect 517518 247415 517574 247424
rect 517520 247036 517572 247042
rect 517520 246978 517572 246984
rect 517532 246129 517560 246978
rect 517518 246120 517574 246129
rect 517518 246055 517574 246064
rect 517520 245608 517572 245614
rect 517520 245550 517572 245556
rect 517532 244769 517560 245550
rect 517518 244760 517574 244769
rect 517518 244695 517574 244704
rect 517518 243400 517574 243409
rect 517518 243335 517574 243344
rect 517532 242962 517560 243335
rect 517520 242956 517572 242962
rect 517520 242898 517572 242904
rect 518176 227730 518204 403271
rect 518268 248402 518296 404631
rect 520660 402974 520688 421382
rect 523682 421288 523738 421297
rect 523682 421223 523738 421232
rect 526166 421288 526222 421297
rect 526166 421223 526222 421232
rect 529308 404977 529336 421382
rect 529294 404968 529350 404977
rect 529294 404903 529350 404912
rect 520660 402946 520872 402974
rect 520844 381426 520872 402946
rect 523682 383752 523738 383761
rect 523682 383687 523738 383696
rect 526166 383752 526222 383761
rect 526166 383687 526222 383696
rect 523696 381956 523724 383687
rect 526180 381956 526208 383687
rect 529308 381426 529336 404903
rect 520844 381398 521226 381426
rect 528678 381398 529336 381426
rect 520844 373994 520872 381398
rect 520660 373966 520872 373994
rect 529124 373994 529152 381398
rect 529124 373966 529336 373994
rect 518530 367432 518586 367441
rect 518530 367367 518586 367376
rect 518346 363352 518402 363361
rect 518346 363287 518402 363296
rect 518256 248396 518308 248402
rect 518256 248338 518308 248344
rect 518254 242040 518310 242049
rect 518254 241975 518310 241984
rect 518164 227724 518216 227730
rect 518164 227666 518216 227672
rect 518268 210186 518296 241975
rect 518360 227662 518388 363287
rect 518438 323368 518494 323377
rect 518438 323303 518494 323312
rect 518348 227656 518400 227662
rect 518348 227598 518400 227604
rect 518452 227594 518480 323303
rect 518544 288386 518572 367367
rect 520660 364334 520688 373966
rect 520660 364306 520872 364334
rect 520844 341442 520872 364306
rect 529308 345014 529336 373966
rect 529124 344986 529336 345014
rect 529124 341442 529152 344986
rect 520844 341414 521226 341442
rect 528678 341414 529152 341442
rect 520844 335354 520872 341414
rect 523682 341320 523738 341329
rect 523682 341255 523738 341264
rect 526166 341320 526222 341329
rect 526166 341255 526222 341264
rect 520660 335326 520872 335354
rect 529124 335354 529152 341414
rect 529124 335326 529336 335354
rect 520660 325694 520688 335326
rect 520660 325666 520872 325694
rect 520844 301458 520872 325666
rect 529308 306374 529336 335326
rect 529032 306346 529336 306374
rect 526166 303648 526222 303657
rect 526166 303583 526222 303592
rect 523682 302288 523738 302297
rect 523682 302223 523738 302232
rect 523696 301852 523724 302223
rect 526180 301852 526208 303583
rect 529032 301866 529060 306346
rect 580170 302288 580226 302297
rect 580170 302223 580226 302232
rect 528678 301838 529336 301866
rect 520844 301430 521226 301458
rect 520844 296714 520872 301430
rect 520660 296686 520872 296714
rect 518532 288380 518584 288386
rect 518532 288322 518584 288328
rect 518714 286104 518770 286113
rect 518714 286039 518770 286048
rect 518622 283384 518678 283393
rect 518622 283319 518678 283328
rect 518530 282024 518586 282033
rect 518530 281959 518586 281968
rect 518440 227588 518492 227594
rect 518440 227530 518492 227536
rect 518256 210180 518308 210186
rect 518256 210122 518308 210128
rect 518544 208350 518572 281959
rect 518636 227526 518664 283319
rect 518728 267714 518756 286039
rect 520660 267734 520688 296686
rect 529308 267734 529336 301838
rect 580184 298761 580212 302223
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 518716 267708 518768 267714
rect 520660 267706 520872 267734
rect 518716 267650 518768 267656
rect 520844 263673 520872 267706
rect 529032 267706 529336 267734
rect 523682 264616 523738 264625
rect 523682 264551 523738 264560
rect 526166 264616 526222 264625
rect 526166 264551 526222 264560
rect 520830 263664 520886 263673
rect 520830 263599 520886 263608
rect 520844 261882 520872 263599
rect 520844 261854 521226 261882
rect 523696 261868 523724 264551
rect 526180 261868 526208 264551
rect 529032 261882 529060 267706
rect 580262 263664 580318 263673
rect 580262 263599 580318 263608
rect 528678 261854 529060 261882
rect 580276 245585 580304 263599
rect 580262 245576 580318 245585
rect 580262 245511 580318 245520
rect 518624 227520 518676 227526
rect 518624 227462 518676 227468
rect 580446 213344 580502 213353
rect 580446 213279 580502 213288
rect 580262 213208 580318 213217
rect 580262 213143 580318 213152
rect 518532 208344 518584 208350
rect 518532 208286 518584 208292
rect 327724 208276 327776 208282
rect 327724 208218 327776 208224
rect 322204 208208 322256 208214
rect 322204 208150 322256 208156
rect 295524 208140 295576 208146
rect 295524 208082 295576 208088
rect 318064 208140 318116 208146
rect 318064 208082 318116 208088
rect 580276 126041 580304 213143
rect 580460 165889 580488 213279
rect 580908 211880 580960 211886
rect 580908 211822 580960 211828
rect 580920 205737 580948 211822
rect 580906 205728 580962 205737
rect 580906 205663 580962 205672
rect 580446 165880 580502 165889
rect 580446 165815 580502 165824
rect 580262 126032 580318 126041
rect 580262 125967 580318 125976
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
<< via2 >>
rect 294778 490592 294834 490648
rect 297934 490592 297990 490648
rect 301089 490592 301145 490648
rect 304246 490592 304302 490648
rect 295614 487192 295670 487248
rect 307403 490320 307459 490376
rect 305090 487192 305146 487248
rect 301560 451152 301616 451208
rect 304877 451152 304933 451208
rect 294510 450880 294566 450936
rect 307758 450880 307814 450936
rect 298282 450472 298338 450528
rect 295890 447208 295946 447264
rect 298190 431160 298246 431216
rect 294694 431024 294750 431080
rect 301594 431024 301650 431080
rect 308402 430888 308458 430944
rect 304998 430616 305054 430672
rect 306194 426400 306250 426456
rect 298190 411304 298246 411360
rect 295154 410080 295210 410136
rect 301594 410080 301650 410136
rect 304722 410080 304778 410136
rect 308218 410080 308274 410136
rect 295338 391448 295394 391504
rect 298190 391176 298246 391232
rect 299202 391448 299258 391504
rect 301594 391180 301596 391232
rect 301596 391180 301648 391232
rect 301648 391180 301650 391232
rect 301594 391176 301650 391180
rect 305366 391040 305422 391096
rect 309138 391040 309194 391096
rect 303618 386824 303674 386880
rect 307298 386824 307354 386880
rect 294510 369960 294566 370016
rect 298006 369960 298062 370016
rect 300766 369960 300822 370016
rect 304170 369960 304226 370016
rect 306930 369960 306986 370016
rect 304908 291488 304964 291544
rect 300122 291352 300178 291408
rect 306746 291352 306802 291408
rect 294602 291216 294658 291272
rect 298098 291216 298154 291272
rect 294694 271496 294750 271552
rect 298498 271496 298554 271552
rect 301410 271496 301466 271552
rect 304998 271496 305054 271552
rect 308310 271496 308366 271552
rect 298650 251504 298706 251560
rect 294878 251368 294934 251424
rect 301410 251504 301466 251560
rect 308218 251504 308274 251560
rect 308954 251504 309010 251560
rect 304669 250960 304725 251016
rect 309138 233280 309194 233336
rect 295338 231376 295394 231432
rect 299033 231376 299089 231432
rect 302745 230560 302801 230616
rect 299018 230152 299074 230208
rect 306457 230560 306513 230616
rect 310150 230560 310206 230616
rect 307022 213288 307078 213344
rect 303894 213152 303950 213208
rect 303894 211792 303950 211848
rect 307022 211792 307078 211848
rect 306930 211520 306986 211576
rect 303817 211384 303873 211440
rect 300765 211112 300821 211168
rect 294694 210432 294750 210488
rect 297730 210432 297786 210488
rect 517518 416880 517574 416936
rect 518162 415520 518218 415576
rect 517518 414160 517574 414216
rect 517518 412800 517574 412856
rect 517518 407360 517574 407416
rect 517518 406000 517574 406056
rect 518254 404640 518310 404696
rect 518162 403280 518218 403336
rect 517518 401920 517574 401976
rect 517518 380976 517574 381032
rect 517518 378256 517574 378312
rect 517518 376896 517574 376952
rect 517518 375536 517574 375592
rect 517518 374176 517574 374232
rect 517518 372816 517574 372872
rect 517518 366016 517574 366072
rect 517518 364656 517574 364712
rect 517518 361936 517574 361992
rect 517518 340992 517574 341048
rect 517518 338272 517574 338328
rect 517518 336912 517574 336968
rect 517518 335552 517574 335608
rect 517518 332832 517574 332888
rect 517518 327392 517574 327448
rect 517518 326032 517574 326088
rect 517518 324672 517574 324728
rect 517518 321952 517574 322008
rect 517518 298288 517574 298344
rect 517518 295568 517574 295624
rect 517518 292848 517574 292904
rect 517518 287408 517574 287464
rect 517518 284688 517574 284744
rect 517518 261024 517574 261080
rect 517518 258304 517574 258360
rect 517518 256944 517574 257000
rect 517518 255584 517574 255640
rect 517518 254224 517574 254280
rect 517518 252864 517574 252920
rect 517518 247424 517574 247480
rect 517518 246064 517574 246120
rect 517518 244704 517574 244760
rect 517518 243344 517574 243400
rect 523682 421232 523738 421288
rect 526166 421232 526222 421288
rect 529294 404912 529350 404968
rect 523682 383696 523738 383752
rect 526166 383696 526222 383752
rect 518530 367376 518586 367432
rect 518346 363296 518402 363352
rect 518254 241984 518310 242040
rect 518438 323312 518494 323368
rect 523682 341264 523738 341320
rect 526166 341264 526222 341320
rect 526166 303592 526222 303648
rect 523682 302232 523738 302288
rect 580170 302232 580226 302288
rect 518714 286048 518770 286104
rect 518622 283328 518678 283384
rect 518530 281968 518586 282024
rect 580170 298696 580226 298752
rect 523682 264560 523738 264616
rect 526166 264560 526222 264616
rect 520830 263608 520886 263664
rect 580262 263608 580318 263664
rect 580262 245520 580318 245576
rect 580446 213288 580502 213344
rect 580262 213152 580318 213208
rect 580906 205672 580962 205728
rect 580446 165824 580502 165880
rect 580262 125976 580318 126032
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect 294773 490652 294839 490653
rect 297929 490652 297995 490653
rect 301084 490652 301150 490653
rect 304241 490652 304307 490653
rect 294773 490648 294828 490652
rect 294892 490650 294898 490652
rect 294773 490592 294778 490648
rect 294773 490588 294828 490592
rect 294892 490590 294930 490650
rect 297929 490648 297956 490652
rect 298020 490650 298026 490652
rect 297929 490592 297934 490648
rect 294892 490588 294898 490590
rect 297929 490588 297956 490592
rect 298020 490590 298086 490650
rect 298020 490588 298026 490590
rect 301078 490588 301084 490652
rect 301148 490650 301154 490652
rect 301148 490590 301240 490650
rect 301148 490588 301154 490590
rect 304206 490588 304212 490652
rect 304276 490650 304307 490652
rect 304276 490648 304368 490650
rect 304302 490592 304368 490648
rect 304276 490590 304368 490592
rect 304276 490588 304307 490590
rect 294773 490587 294839 490588
rect 297929 490587 297995 490588
rect 301084 490587 301150 490588
rect 304241 490587 304307 490588
rect 307398 490380 307464 490381
rect 307334 490378 307340 490380
rect 307307 490318 307340 490378
rect 307404 490376 307464 490380
rect 307459 490320 307464 490376
rect 307334 490316 307340 490318
rect 307404 490316 307464 490320
rect 307398 490315 307464 490316
rect -960 488596 480 488836
rect 295609 487250 295675 487253
rect 296478 487250 296484 487252
rect 295609 487248 296484 487250
rect 295609 487192 295614 487248
rect 295670 487192 296484 487248
rect 295609 487190 296484 487192
rect 295609 487187 295675 487190
rect 296478 487188 296484 487190
rect 296548 487188 296554 487252
rect 305085 487250 305151 487253
rect 306230 487250 306236 487252
rect 305085 487248 306236 487250
rect 305085 487192 305090 487248
rect 305146 487192 306236 487248
rect 305085 487190 306236 487192
rect 305085 487187 305151 487190
rect 306230 487188 306236 487190
rect 306300 487188 306306 487252
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect 301262 451148 301268 451212
rect 301332 451210 301338 451212
rect 301555 451210 301621 451213
rect 301332 451208 301621 451210
rect 301332 451152 301560 451208
rect 301616 451152 301621 451208
rect 301332 451150 301621 451152
rect 301332 451148 301338 451150
rect 301555 451147 301621 451150
rect 304574 451148 304580 451212
rect 304644 451210 304650 451212
rect 304872 451210 304938 451213
rect 304644 451208 304938 451210
rect 304644 451152 304877 451208
rect 304933 451152 304938 451208
rect 304644 451150 304938 451152
rect 304644 451148 304650 451150
rect 304872 451147 304938 451150
rect 294505 450940 294571 450941
rect 307753 450940 307819 450941
rect 294454 450876 294460 450940
rect 294524 450938 294571 450940
rect 294524 450936 294616 450938
rect 294566 450880 294616 450936
rect 294524 450878 294616 450880
rect 294524 450876 294571 450878
rect 307702 450876 307708 450940
rect 307772 450938 307819 450940
rect 307772 450936 307864 450938
rect 307814 450880 307864 450936
rect 307772 450878 307864 450880
rect 307772 450876 307819 450878
rect 294505 450875 294571 450876
rect 307753 450875 307819 450876
rect 298134 450468 298140 450532
rect 298204 450530 298210 450532
rect 298277 450530 298343 450533
rect 298204 450528 298343 450530
rect 298204 450472 298282 450528
rect 298338 450472 298343 450528
rect 298204 450470 298343 450472
rect 298204 450468 298210 450470
rect 298277 450467 298343 450470
rect -960 449428 480 449668
rect 295885 447266 295951 447269
rect 296294 447266 296300 447268
rect 295885 447264 296300 447266
rect 295885 447208 295890 447264
rect 295946 447208 296300 447264
rect 295885 447206 296300 447208
rect 295885 447203 295951 447206
rect 296294 447204 296300 447206
rect 296364 447204 296370 447268
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect 298185 431220 298251 431221
rect 298134 431156 298140 431220
rect 298204 431218 298251 431220
rect 299238 431218 299244 431220
rect 298204 431216 299244 431218
rect 298246 431160 299244 431216
rect 298204 431158 299244 431160
rect 298204 431156 298251 431158
rect 299238 431156 299244 431158
rect 299308 431156 299314 431220
rect 298185 431155 298251 431156
rect 294454 431020 294460 431084
rect 294524 431082 294530 431084
rect 294689 431082 294755 431085
rect 294524 431080 294755 431082
rect 294524 431024 294694 431080
rect 294750 431024 294755 431080
rect 294524 431022 294755 431024
rect 294524 431020 294530 431022
rect 294689 431019 294755 431022
rect 301446 431020 301452 431084
rect 301516 431082 301522 431084
rect 301589 431082 301655 431085
rect 301516 431080 301655 431082
rect 301516 431024 301594 431080
rect 301650 431024 301655 431080
rect 301516 431022 301655 431024
rect 301516 431020 301522 431022
rect 301589 431019 301655 431022
rect 308254 430884 308260 430948
rect 308324 430946 308330 430948
rect 308397 430946 308463 430949
rect 308324 430944 308463 430946
rect 308324 430888 308402 430944
rect 308458 430888 308463 430944
rect 308324 430886 308463 430888
rect 308324 430884 308330 430886
rect 308397 430883 308463 430886
rect 304758 430612 304764 430676
rect 304828 430674 304834 430676
rect 304993 430674 305059 430677
rect 304828 430672 305059 430674
rect 304828 430616 304998 430672
rect 305054 430616 305059 430672
rect 304828 430614 305059 430616
rect 304828 430612 304834 430614
rect 304993 430611 305059 430614
rect 306046 426396 306052 426460
rect 306116 426458 306122 426460
rect 306189 426458 306255 426461
rect 306116 426456 306255 426458
rect 306116 426400 306194 426456
rect 306250 426400 306255 426456
rect 306116 426398 306255 426400
rect 306116 426396 306122 426398
rect 306189 426395 306255 426398
rect -960 423452 480 423692
rect 523534 421228 523540 421292
rect 523604 421290 523610 421292
rect 523677 421290 523743 421293
rect 523604 421288 523743 421290
rect 523604 421232 523682 421288
rect 523738 421232 523743 421288
rect 523604 421230 523743 421232
rect 523604 421228 523610 421230
rect 523677 421227 523743 421230
rect 526161 421290 526227 421293
rect 526294 421290 526300 421292
rect 526161 421288 526300 421290
rect 526161 421232 526166 421288
rect 526222 421232 526300 421288
rect 526161 421230 526300 421232
rect 526161 421227 526227 421230
rect 526294 421228 526300 421230
rect 526364 421228 526370 421292
rect 296478 421092 296484 421156
rect 296548 421154 296554 421156
rect 296548 421094 509250 421154
rect 296548 421092 296554 421094
rect 509190 421018 509250 421094
rect 509190 420958 520076 421018
rect 296294 418372 296300 418436
rect 296364 418434 296370 418436
rect 296364 418374 509250 418434
rect 296364 418372 296370 418374
rect 509190 418298 509250 418374
rect 509190 418238 520076 418298
rect 583520 418148 584960 418388
rect 517513 416938 517579 416941
rect 517513 416936 520076 416938
rect 517513 416880 517518 416936
rect 517574 416880 520076 416936
rect 517513 416878 520076 416880
rect 517513 416875 517579 416878
rect 518157 415578 518223 415581
rect 518157 415576 520076 415578
rect 518157 415520 518162 415576
rect 518218 415520 520076 415576
rect 518157 415518 520076 415520
rect 518157 415515 518223 415518
rect 517513 414218 517579 414221
rect 517513 414216 520076 414218
rect 517513 414160 517518 414216
rect 517574 414160 520076 414216
rect 517513 414158 520076 414160
rect 517513 414155 517579 414158
rect 517513 412858 517579 412861
rect 517513 412856 520076 412858
rect 517513 412800 517518 412856
rect 517574 412800 520076 412856
rect 517513 412798 520076 412800
rect 517513 412795 517579 412798
rect 298185 411362 298251 411365
rect 299238 411362 299244 411364
rect 298185 411360 299244 411362
rect 298185 411304 298190 411360
rect 298246 411304 299244 411360
rect 298185 411302 299244 411304
rect 298185 411299 298251 411302
rect 299238 411300 299244 411302
rect 299308 411300 299314 411364
rect 531446 410954 531452 410956
rect 529828 410894 531452 410954
rect 531446 410892 531452 410894
rect 531516 410892 531522 410956
rect -960 410396 480 410636
rect 295149 410140 295215 410141
rect 301589 410140 301655 410141
rect 304717 410140 304783 410141
rect 308213 410140 308279 410141
rect 295149 410138 295196 410140
rect 295104 410136 295196 410138
rect 295104 410080 295154 410136
rect 295104 410078 295196 410080
rect 295149 410076 295196 410078
rect 295260 410076 295266 410140
rect 301589 410138 301636 410140
rect 301544 410136 301636 410138
rect 301544 410080 301594 410136
rect 301544 410078 301636 410080
rect 301589 410076 301636 410078
rect 301700 410076 301706 410140
rect 304717 410138 304764 410140
rect 304672 410136 304764 410138
rect 304672 410080 304722 410136
rect 304672 410078 304764 410080
rect 304717 410076 304764 410078
rect 304828 410076 304834 410140
rect 308213 410138 308260 410140
rect 308168 410136 308260 410138
rect 308168 410080 308218 410136
rect 308168 410078 308260 410080
rect 308213 410076 308260 410078
rect 308324 410076 308330 410140
rect 295149 410075 295215 410076
rect 301589 410075 301655 410076
rect 304717 410075 304783 410076
rect 308213 410075 308279 410076
rect 517513 407418 517579 407421
rect 517513 407416 520076 407418
rect 517513 407360 517518 407416
rect 517574 407360 520076 407416
rect 517513 407358 520076 407360
rect 517513 407355 517579 407358
rect 517513 406058 517579 406061
rect 517513 406056 520076 406058
rect 517513 406000 517518 406056
rect 517574 406000 520076 406056
rect 517513 405998 520076 406000
rect 517513 405995 517579 405998
rect 529289 404970 529355 404973
rect 583520 404970 584960 405060
rect 529289 404968 584960 404970
rect 529289 404912 529294 404968
rect 529350 404912 584960 404968
rect 529289 404910 584960 404912
rect 529289 404907 529355 404910
rect 583520 404820 584960 404910
rect 518249 404698 518315 404701
rect 518249 404696 520076 404698
rect 518249 404640 518254 404696
rect 518310 404640 520076 404696
rect 518249 404638 520076 404640
rect 518249 404635 518315 404638
rect 518157 403338 518223 403341
rect 518157 403336 520076 403338
rect 518157 403280 518162 403336
rect 518218 403280 520076 403336
rect 518157 403278 520076 403280
rect 518157 403275 518223 403278
rect 517513 401978 517579 401981
rect 517513 401976 520076 401978
rect 517513 401920 517518 401976
rect 517574 401920 520076 401976
rect 517513 401918 520076 401920
rect 517513 401915 517579 401918
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect 295190 391444 295196 391508
rect 295260 391506 295266 391508
rect 295333 391506 295399 391509
rect 299197 391508 299263 391509
rect 299197 391506 299244 391508
rect 295260 391504 295399 391506
rect 295260 391448 295338 391504
rect 295394 391448 295399 391504
rect 295260 391446 295399 391448
rect 299152 391504 299244 391506
rect 299152 391448 299202 391504
rect 299152 391446 299244 391448
rect 295260 391444 295266 391446
rect 295333 391443 295399 391446
rect 299197 391444 299244 391446
rect 299308 391444 299314 391508
rect 299197 391443 299263 391444
rect 298185 391236 298251 391237
rect 298134 391234 298140 391236
rect 298094 391174 298140 391234
rect 298204 391232 298251 391236
rect 301589 391236 301655 391237
rect 301589 391234 301636 391236
rect 298246 391176 298251 391232
rect 298134 391172 298140 391174
rect 298204 391172 298251 391176
rect 301544 391232 301636 391234
rect 301544 391176 301594 391232
rect 301544 391174 301636 391176
rect 298185 391171 298251 391172
rect 301589 391172 301636 391174
rect 301700 391172 301706 391236
rect 301589 391171 301655 391172
rect 304758 391036 304764 391100
rect 304828 391098 304834 391100
rect 305361 391098 305427 391101
rect 304828 391096 305427 391098
rect 304828 391040 305366 391096
rect 305422 391040 305427 391096
rect 304828 391038 305427 391040
rect 304828 391036 304834 391038
rect 305361 391035 305427 391038
rect 307702 391036 307708 391100
rect 307772 391098 307778 391100
rect 309133 391098 309199 391101
rect 307772 391096 309199 391098
rect 307772 391040 309138 391096
rect 309194 391040 309199 391096
rect 307772 391038 309199 391040
rect 307772 391036 307778 391038
rect 309133 391035 309199 391038
rect 303613 386882 303679 386885
rect 304758 386882 304764 386884
rect 303613 386880 304764 386882
rect 303613 386824 303618 386880
rect 303674 386824 304764 386880
rect 303613 386822 304764 386824
rect 303613 386819 303679 386822
rect 304758 386820 304764 386822
rect 304828 386820 304834 386884
rect 307293 386882 307359 386885
rect 307518 386882 307524 386884
rect 307293 386880 307524 386882
rect 307293 386824 307298 386880
rect 307354 386824 307524 386880
rect 307293 386822 307524 386824
rect 307293 386819 307359 386822
rect 307518 386820 307524 386822
rect 307588 386820 307594 386884
rect -960 384284 480 384524
rect 523534 383692 523540 383756
rect 523604 383754 523610 383756
rect 523677 383754 523743 383757
rect 523604 383752 523743 383754
rect 523604 383696 523682 383752
rect 523738 383696 523743 383752
rect 523604 383694 523743 383696
rect 523604 383692 523610 383694
rect 523677 383691 523743 383694
rect 526161 383754 526227 383757
rect 526294 383754 526300 383756
rect 526161 383752 526300 383754
rect 526161 383696 526166 383752
rect 526222 383696 526300 383752
rect 526161 383694 526300 383696
rect 526161 383691 526227 383694
rect 526294 383692 526300 383694
rect 526364 383692 526370 383756
rect 517513 381034 517579 381037
rect 517513 381032 520076 381034
rect 517513 380976 517518 381032
rect 517574 380976 520076 381032
rect 517513 380974 520076 380976
rect 517513 380971 517579 380974
rect 517513 378314 517579 378317
rect 517513 378312 520076 378314
rect 517513 378256 517518 378312
rect 517574 378256 520076 378312
rect 583520 378300 584960 378540
rect 517513 378254 520076 378256
rect 517513 378251 517579 378254
rect 517513 376954 517579 376957
rect 517513 376952 520076 376954
rect 517513 376896 517518 376952
rect 517574 376896 520076 376952
rect 517513 376894 520076 376896
rect 517513 376891 517579 376894
rect 517513 375594 517579 375597
rect 517513 375592 520076 375594
rect 517513 375536 517518 375592
rect 517574 375536 520076 375592
rect 517513 375534 520076 375536
rect 517513 375531 517579 375534
rect 517513 374234 517579 374237
rect 517513 374232 520076 374234
rect 517513 374176 517518 374232
rect 517574 374176 520076 374232
rect 517513 374174 520076 374176
rect 517513 374171 517579 374174
rect 517513 372874 517579 372877
rect 517513 372872 520076 372874
rect 517513 372816 517518 372872
rect 517574 372816 520076 372872
rect 517513 372814 520076 372816
rect 517513 372811 517579 372814
rect -960 371228 480 371468
rect 531446 370970 531452 370972
rect 529828 370910 531452 370970
rect 531446 370908 531452 370910
rect 531516 370908 531522 370972
rect 294505 370020 294571 370021
rect 294454 369956 294460 370020
rect 294524 370018 294571 370020
rect 298001 370018 298067 370021
rect 300761 370020 300827 370021
rect 298134 370018 298140 370020
rect 294524 370016 294616 370018
rect 294566 369960 294616 370016
rect 294524 369958 294616 369960
rect 298001 370016 298140 370018
rect 298001 369960 298006 370016
rect 298062 369960 298140 370016
rect 298001 369958 298140 369960
rect 294524 369956 294571 369958
rect 294505 369955 294571 369956
rect 298001 369955 298067 369958
rect 298134 369956 298140 369958
rect 298204 369956 298210 370020
rect 300710 369956 300716 370020
rect 300780 370018 300827 370020
rect 304165 370020 304231 370021
rect 306925 370020 306991 370021
rect 304165 370018 304212 370020
rect 300780 370016 300872 370018
rect 300822 369960 300872 370016
rect 300780 369958 300872 369960
rect 304120 370016 304212 370018
rect 304120 369960 304170 370016
rect 304120 369958 304212 369960
rect 300780 369956 300827 369958
rect 300761 369955 300827 369956
rect 304165 369956 304212 369958
rect 304276 369956 304282 370020
rect 306925 370018 306972 370020
rect 306880 370016 306972 370018
rect 306880 369960 306930 370016
rect 306880 369958 306972 369960
rect 306925 369956 306972 369958
rect 307036 369956 307042 370020
rect 304165 369955 304231 369956
rect 306925 369955 306991 369956
rect 518525 367434 518591 367437
rect 518525 367432 520076 367434
rect 518525 367376 518530 367432
rect 518586 367376 520076 367432
rect 518525 367374 520076 367376
rect 518525 367371 518591 367374
rect 517513 366074 517579 366077
rect 517513 366072 520076 366074
rect 517513 366016 517518 366072
rect 517574 366016 520076 366072
rect 517513 366014 520076 366016
rect 517513 366011 517579 366014
rect 583520 364972 584960 365212
rect 517513 364714 517579 364717
rect 517513 364712 520076 364714
rect 517513 364656 517518 364712
rect 517574 364656 520076 364712
rect 517513 364654 520076 364656
rect 517513 364651 517579 364654
rect 518341 363354 518407 363357
rect 518341 363352 520076 363354
rect 518341 363296 518346 363352
rect 518402 363296 520076 363352
rect 518341 363294 520076 363296
rect 518341 363291 518407 363294
rect 517513 361994 517579 361997
rect 517513 361992 520076 361994
rect 517513 361936 517518 361992
rect 517574 361936 520076 361992
rect 517513 361934 520076 361936
rect 517513 361931 517579 361934
rect -960 358308 480 358548
rect 527030 351868 527036 351932
rect 527100 351930 527106 351932
rect 583520 351930 584960 352020
rect 527100 351870 584960 351930
rect 527100 351868 527106 351870
rect 583520 351780 584960 351870
rect -960 345252 480 345492
rect 523534 341260 523540 341324
rect 523604 341322 523610 341324
rect 523677 341322 523743 341325
rect 523604 341320 523743 341322
rect 523604 341264 523682 341320
rect 523738 341264 523743 341320
rect 523604 341262 523743 341264
rect 523604 341260 523610 341262
rect 523677 341259 523743 341262
rect 526161 341322 526227 341325
rect 526294 341322 526300 341324
rect 526161 341320 526300 341322
rect 526161 341264 526166 341320
rect 526222 341264 526300 341320
rect 526161 341262 526300 341264
rect 526161 341259 526227 341262
rect 526294 341260 526300 341262
rect 526364 341260 526370 341324
rect 517513 341050 517579 341053
rect 517513 341048 520076 341050
rect 517513 340992 517518 341048
rect 517574 340992 520076 341048
rect 517513 340990 520076 340992
rect 517513 340987 517579 340990
rect 583520 338452 584960 338692
rect 517513 338330 517579 338333
rect 517513 338328 520076 338330
rect 517513 338272 517518 338328
rect 517574 338272 520076 338328
rect 517513 338270 520076 338272
rect 517513 338267 517579 338270
rect 517513 336970 517579 336973
rect 517513 336968 520076 336970
rect 517513 336912 517518 336968
rect 517574 336912 520076 336968
rect 517513 336910 520076 336912
rect 517513 336907 517579 336910
rect 517513 335610 517579 335613
rect 517513 335608 520076 335610
rect 517513 335552 517518 335608
rect 517574 335552 520076 335608
rect 517513 335550 520076 335552
rect 517513 335547 517579 335550
rect 304758 334188 304764 334252
rect 304828 334250 304834 334252
rect 304828 334190 520076 334250
rect 304828 334188 304834 334190
rect 517513 332890 517579 332893
rect 517513 332888 520076 332890
rect 517513 332832 517518 332888
rect 517574 332832 520076 332888
rect 517513 332830 520076 332832
rect 517513 332827 517579 332830
rect -960 332196 480 332436
rect 531446 330986 531452 330988
rect 529828 330926 531452 330986
rect 531446 330924 531452 330926
rect 531516 330924 531522 330988
rect 517513 327450 517579 327453
rect 517513 327448 520076 327450
rect 517513 327392 517518 327448
rect 517574 327392 520076 327448
rect 517513 327390 520076 327392
rect 517513 327387 517579 327390
rect 517513 326090 517579 326093
rect 517513 326088 520076 326090
rect 517513 326032 517518 326088
rect 517574 326032 520076 326088
rect 517513 326030 520076 326032
rect 517513 326027 517579 326030
rect 583520 325124 584960 325364
rect 517513 324730 517579 324733
rect 517513 324728 520076 324730
rect 517513 324672 517518 324728
rect 517574 324672 520076 324728
rect 517513 324670 520076 324672
rect 517513 324667 517579 324670
rect 518433 323370 518499 323373
rect 518433 323368 520076 323370
rect 518433 323312 518438 323368
rect 518494 323312 520076 323368
rect 518433 323310 520076 323312
rect 518433 323307 518499 323310
rect 517513 322010 517579 322013
rect 517513 322008 520076 322010
rect 517513 321952 517518 322008
rect 517574 321952 520076 322008
rect 517513 321950 520076 321952
rect 517513 321947 517579 321950
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 526161 303650 526227 303653
rect 526294 303650 526300 303652
rect 526161 303648 526300 303650
rect 526161 303592 526166 303648
rect 526222 303592 526300 303648
rect 526161 303590 526300 303592
rect 526161 303587 526227 303590
rect 526294 303588 526300 303590
rect 526364 303588 526370 303652
rect 523534 302228 523540 302292
rect 523604 302290 523610 302292
rect 523677 302290 523743 302293
rect 524270 302290 524276 302292
rect 523604 302288 524276 302290
rect 523604 302232 523682 302288
rect 523738 302232 524276 302288
rect 523604 302230 524276 302232
rect 523604 302228 523610 302230
rect 523677 302227 523743 302230
rect 524270 302228 524276 302230
rect 524340 302290 524346 302292
rect 580165 302290 580231 302293
rect 524340 302288 580231 302290
rect 524340 302232 580170 302288
rect 580226 302232 580231 302288
rect 524340 302230 580231 302232
rect 524340 302228 524346 302230
rect 580165 302227 580231 302230
rect 306230 301004 306236 301068
rect 306300 301066 306306 301068
rect 306300 301006 520076 301066
rect 306300 301004 306306 301006
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 517513 298346 517579 298349
rect 517513 298344 520076 298346
rect 517513 298288 517518 298344
rect 517574 298288 520076 298344
rect 517513 298286 520076 298288
rect 517513 298283 517579 298286
rect 306046 296924 306052 296988
rect 306116 296986 306122 296988
rect 306116 296926 520076 296986
rect 306116 296924 306122 296926
rect 517513 295626 517579 295629
rect 517513 295624 520076 295626
rect 517513 295568 517518 295624
rect 517574 295568 520076 295624
rect 517513 295566 520076 295568
rect 517513 295563 517579 295566
rect 307518 294204 307524 294268
rect 307588 294266 307594 294268
rect 307588 294206 520076 294266
rect 307588 294204 307594 294206
rect -960 293028 480 293268
rect 517513 292906 517579 292909
rect 517513 292904 520076 292906
rect 517513 292848 517518 292904
rect 517574 292848 520076 292904
rect 517513 292846 520076 292848
rect 517513 292843 517579 292846
rect 304206 291484 304212 291548
rect 304276 291546 304282 291548
rect 304758 291546 304764 291548
rect 304276 291486 304764 291546
rect 304276 291484 304282 291486
rect 304758 291484 304764 291486
rect 304828 291546 304834 291548
rect 304903 291546 304969 291549
rect 304828 291544 304969 291546
rect 304828 291488 304908 291544
rect 304964 291488 304969 291544
rect 304828 291486 304969 291488
rect 304828 291484 304834 291486
rect 304903 291483 304969 291486
rect 300117 291412 300183 291413
rect 306741 291412 306807 291413
rect 300117 291410 300164 291412
rect 300072 291408 300164 291410
rect 300072 291352 300122 291408
rect 300072 291350 300164 291352
rect 300117 291348 300164 291350
rect 300228 291348 300234 291412
rect 306741 291410 306788 291412
rect 306696 291408 306788 291410
rect 306696 291352 306746 291408
rect 306696 291350 306788 291352
rect 306741 291348 306788 291350
rect 306852 291348 306858 291412
rect 300117 291347 300183 291348
rect 306741 291347 306807 291348
rect 294454 291212 294460 291276
rect 294524 291274 294530 291276
rect 294597 291274 294663 291277
rect 298093 291276 298159 291277
rect 298093 291274 298140 291276
rect 294524 291272 294663 291274
rect 294524 291216 294602 291272
rect 294658 291216 294663 291272
rect 294524 291214 294663 291216
rect 298048 291272 298140 291274
rect 298204 291274 298210 291276
rect 299238 291274 299244 291276
rect 298048 291216 298098 291272
rect 298048 291214 298140 291216
rect 294524 291212 294530 291214
rect 294597 291211 294663 291214
rect 298093 291212 298140 291214
rect 298204 291214 299244 291274
rect 298204 291212 298210 291214
rect 299238 291212 299244 291214
rect 299308 291212 299314 291276
rect 298093 291211 298159 291212
rect 531446 291002 531452 291004
rect 529828 290942 531452 291002
rect 531446 290940 531452 290942
rect 531516 290940 531522 291004
rect 517513 287466 517579 287469
rect 517513 287464 520076 287466
rect 517513 287408 517518 287464
rect 517574 287408 520076 287464
rect 517513 287406 520076 287408
rect 517513 287403 517579 287406
rect 518709 286106 518775 286109
rect 518709 286104 520076 286106
rect 518709 286048 518714 286104
rect 518770 286048 520076 286104
rect 518709 286046 520076 286048
rect 518709 286043 518775 286046
rect 583520 285276 584960 285516
rect 517513 284746 517579 284749
rect 517513 284744 520076 284746
rect 517513 284688 517518 284744
rect 517574 284688 520076 284744
rect 517513 284686 520076 284688
rect 517513 284683 517579 284686
rect 518617 283386 518683 283389
rect 518617 283384 520076 283386
rect 518617 283328 518622 283384
rect 518678 283328 520076 283384
rect 518617 283326 520076 283328
rect 518617 283323 518683 283326
rect 518525 282026 518591 282029
rect 518525 282024 520076 282026
rect 518525 281968 518530 282024
rect 518586 281968 520076 282024
rect 518525 281966 520076 281968
rect 518525 281963 518591 281966
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect 300894 271764 300900 271828
rect 300964 271764 300970 271828
rect 300902 271690 300962 271764
rect 300902 271630 301514 271690
rect 301454 271557 301514 271630
rect 307702 271628 307708 271692
rect 307772 271690 307778 271692
rect 307772 271630 308322 271690
rect 307772 271628 307778 271630
rect 308262 271557 308322 271630
rect 294689 271556 294755 271557
rect 294638 271492 294644 271556
rect 294708 271554 294755 271556
rect 298493 271554 298559 271557
rect 301405 271556 301514 271557
rect 304993 271556 305059 271557
rect 308262 271556 308371 271557
rect 299238 271554 299244 271556
rect 294708 271552 294800 271554
rect 294750 271496 294800 271552
rect 294708 271494 294800 271496
rect 298493 271552 299244 271554
rect 298493 271496 298498 271552
rect 298554 271496 299244 271552
rect 298493 271494 299244 271496
rect 294708 271492 294755 271494
rect 294689 271491 294755 271492
rect 298493 271491 298559 271494
rect 299238 271492 299244 271494
rect 299308 271492 299314 271556
rect 301405 271552 301452 271556
rect 301516 271554 301522 271556
rect 301405 271496 301410 271552
rect 301405 271492 301452 271496
rect 301516 271494 301604 271554
rect 301516 271492 301522 271494
rect 304942 271492 304948 271556
rect 305012 271554 305059 271556
rect 305012 271552 305104 271554
rect 305054 271496 305104 271552
rect 305012 271494 305104 271496
rect 305012 271492 305059 271494
rect 308254 271492 308260 271556
rect 308324 271554 308371 271556
rect 308324 271552 308412 271554
rect 308366 271496 308412 271552
rect 308324 271494 308412 271496
rect 308324 271492 308371 271494
rect 301405 271491 301471 271492
rect 304993 271491 305059 271492
rect 308305 271491 308371 271492
rect -960 267052 480 267292
rect 523677 264618 523743 264621
rect 524270 264618 524276 264620
rect 523677 264616 524276 264618
rect 523677 264560 523682 264616
rect 523738 264560 524276 264616
rect 523677 264558 524276 264560
rect 523677 264555 523743 264558
rect 524270 264556 524276 264558
rect 524340 264556 524346 264620
rect 526161 264618 526227 264621
rect 526294 264618 526300 264620
rect 526161 264616 526300 264618
rect 526161 264560 526166 264616
rect 526222 264560 526300 264616
rect 526161 264558 526300 264560
rect 526161 264555 526227 264558
rect 526294 264556 526300 264558
rect 526364 264556 526370 264620
rect 520825 263666 520891 263669
rect 580257 263666 580323 263669
rect 520825 263664 580323 263666
rect 520825 263608 520830 263664
rect 520886 263608 580262 263664
rect 580318 263608 580323 263664
rect 520825 263606 580323 263608
rect 520825 263603 520891 263606
rect 580257 263603 580323 263606
rect 517513 261082 517579 261085
rect 517513 261080 520076 261082
rect 517513 261024 517518 261080
rect 517574 261024 520076 261080
rect 517513 261022 520076 261024
rect 517513 261019 517579 261022
rect 583520 258756 584960 258996
rect 517513 258362 517579 258365
rect 517513 258360 520076 258362
rect 517513 258304 517518 258360
rect 517574 258304 520076 258360
rect 517513 258302 520076 258304
rect 517513 258299 517579 258302
rect 517513 257002 517579 257005
rect 517513 257000 520076 257002
rect 517513 256944 517518 257000
rect 517574 256944 520076 257000
rect 517513 256942 520076 256944
rect 517513 256939 517579 256942
rect 517513 255642 517579 255645
rect 517513 255640 520076 255642
rect 517513 255584 517518 255640
rect 517574 255584 520076 255640
rect 517513 255582 520076 255584
rect 517513 255579 517579 255582
rect 517513 254282 517579 254285
rect 517513 254280 520076 254282
rect -960 253996 480 254236
rect 517513 254224 517518 254280
rect 517574 254224 520076 254280
rect 517513 254222 520076 254224
rect 517513 254219 517579 254222
rect 517513 252922 517579 252925
rect 517513 252920 520076 252922
rect 517513 252864 517518 252920
rect 517574 252864 520076 252920
rect 517513 252862 520076 252864
rect 517513 252859 517579 252862
rect 298645 251562 298711 251565
rect 301405 251564 301471 251565
rect 308213 251564 308279 251565
rect 299238 251562 299244 251564
rect 298645 251560 299244 251562
rect 298645 251504 298650 251560
rect 298706 251504 299244 251560
rect 298645 251502 299244 251504
rect 298645 251499 298711 251502
rect 299238 251500 299244 251502
rect 299308 251500 299314 251564
rect 301405 251562 301452 251564
rect 301360 251560 301452 251562
rect 301516 251562 301522 251564
rect 302734 251562 302740 251564
rect 301360 251504 301410 251560
rect 301360 251502 301452 251504
rect 301405 251500 301452 251502
rect 301516 251502 302740 251562
rect 301516 251500 301522 251502
rect 302734 251500 302740 251502
rect 302804 251500 302810 251564
rect 308213 251562 308260 251564
rect 308168 251560 308260 251562
rect 308324 251562 308330 251564
rect 308949 251562 309015 251565
rect 308324 251560 309015 251562
rect 308168 251504 308218 251560
rect 308324 251504 308954 251560
rect 309010 251504 309015 251560
rect 308168 251502 308260 251504
rect 308213 251500 308260 251502
rect 308324 251502 309015 251504
rect 308324 251500 308330 251502
rect 301405 251499 301471 251500
rect 308213 251499 308279 251500
rect 308949 251499 309015 251502
rect 294873 251426 294939 251429
rect 295374 251426 295380 251428
rect 294873 251424 295380 251426
rect 294873 251368 294878 251424
rect 294934 251368 295380 251424
rect 294873 251366 295380 251368
rect 294873 251363 294939 251366
rect 295374 251364 295380 251366
rect 295444 251364 295450 251428
rect 304664 251018 304730 251021
rect 304942 251018 304948 251020
rect 304664 251016 304948 251018
rect 304664 250960 304669 251016
rect 304725 250960 304948 251016
rect 304664 250958 304948 250960
rect 304664 250955 304730 250958
rect 304942 250956 304948 250958
rect 305012 250956 305018 251020
rect 531446 251018 531452 251020
rect 529828 250958 531452 251018
rect 531446 250956 531452 250958
rect 531516 250956 531522 251020
rect 517513 247482 517579 247485
rect 517513 247480 520076 247482
rect 517513 247424 517518 247480
rect 517574 247424 520076 247480
rect 517513 247422 520076 247424
rect 517513 247419 517579 247422
rect 517513 246122 517579 246125
rect 517513 246120 520076 246122
rect 517513 246064 517518 246120
rect 517574 246064 520076 246120
rect 517513 246062 520076 246064
rect 517513 246059 517579 246062
rect 580257 245578 580323 245581
rect 583520 245578 584960 245668
rect 580257 245576 584960 245578
rect 580257 245520 580262 245576
rect 580318 245520 584960 245576
rect 580257 245518 584960 245520
rect 580257 245515 580323 245518
rect 583520 245428 584960 245518
rect 517513 244762 517579 244765
rect 517513 244760 520076 244762
rect 517513 244704 517518 244760
rect 517574 244704 520076 244760
rect 517513 244702 520076 244704
rect 517513 244699 517579 244702
rect 517513 243402 517579 243405
rect 517513 243400 520076 243402
rect 517513 243344 517518 243400
rect 517574 243344 520076 243400
rect 517513 243342 520076 243344
rect 517513 243339 517579 243342
rect 518249 242042 518315 242045
rect 518249 242040 520076 242042
rect 518249 241984 518254 242040
rect 518310 241984 520076 242040
rect 518249 241982 520076 241984
rect 518249 241979 518315 241982
rect -960 240940 480 241180
rect 309133 233338 309199 233341
rect 309726 233338 309732 233340
rect 309133 233336 309732 233338
rect 309133 233280 309138 233336
rect 309194 233280 309732 233336
rect 309133 233278 309732 233280
rect 309133 233275 309199 233278
rect 309726 233276 309732 233278
rect 309796 233276 309802 233340
rect 583520 232236 584960 232476
rect 295333 231436 295399 231437
rect 295333 231434 295380 231436
rect 295288 231432 295380 231434
rect 295288 231376 295338 231432
rect 295288 231374 295380 231376
rect 295333 231372 295380 231374
rect 295444 231372 295450 231436
rect 299028 231434 299094 231437
rect 299238 231434 299244 231436
rect 299028 231432 299244 231434
rect 299028 231376 299033 231432
rect 299089 231376 299244 231432
rect 299028 231374 299244 231376
rect 295333 231371 295399 231372
rect 299028 231371 299094 231374
rect 299238 231372 299244 231374
rect 299308 231372 299314 231436
rect 302740 230618 302806 230621
rect 306452 230620 306518 230621
rect 302918 230618 302924 230620
rect 302740 230616 302924 230618
rect 302740 230560 302745 230616
rect 302801 230560 302924 230616
rect 302740 230558 302924 230560
rect 302740 230555 302806 230558
rect 302918 230556 302924 230558
rect 302988 230556 302994 230620
rect 306414 230556 306420 230620
rect 306484 230618 306518 230620
rect 306484 230616 306576 230618
rect 306513 230560 306576 230616
rect 306484 230558 306576 230560
rect 306484 230556 306518 230558
rect 309726 230556 309732 230620
rect 309796 230618 309802 230620
rect 310145 230618 310211 230621
rect 309796 230616 310211 230618
rect 309796 230560 310150 230616
rect 310206 230560 310211 230616
rect 309796 230558 310211 230560
rect 309796 230556 309802 230558
rect 306452 230555 306518 230556
rect 310145 230555 310211 230558
rect 298134 230148 298140 230212
rect 298204 230210 298210 230212
rect 299013 230210 299079 230213
rect 298204 230208 299079 230210
rect 298204 230152 299018 230208
rect 299074 230152 299079 230208
rect 298204 230150 299079 230152
rect 298204 230148 298210 230150
rect 299013 230147 299079 230150
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 307017 213346 307083 213349
rect 309726 213346 309732 213348
rect 307017 213344 309732 213346
rect 307017 213288 307022 213344
rect 307078 213288 309732 213344
rect 307017 213286 309732 213288
rect 307017 213283 307083 213286
rect 309726 213284 309732 213286
rect 309796 213346 309802 213348
rect 580441 213346 580507 213349
rect 309796 213344 580507 213346
rect 309796 213288 580446 213344
rect 580502 213288 580507 213344
rect 309796 213286 580507 213288
rect 309796 213284 309802 213286
rect 580441 213283 580507 213286
rect 303889 213210 303955 213213
rect 306414 213210 306420 213212
rect 303889 213208 306420 213210
rect 303889 213152 303894 213208
rect 303950 213152 306420 213208
rect 303889 213150 306420 213152
rect 303889 213147 303955 213150
rect 306414 213148 306420 213150
rect 306484 213210 306490 213212
rect 580257 213210 580323 213213
rect 306484 213208 580323 213210
rect 306484 213152 580262 213208
rect 580318 213152 580323 213208
rect 306484 213150 580323 213152
rect 306484 213148 306490 213150
rect 580257 213147 580323 213150
rect 303889 211850 303955 211853
rect 307017 211850 307083 211853
rect 303846 211848 303955 211850
rect 303846 211792 303894 211848
rect 303950 211792 303955 211848
rect 303846 211787 303955 211792
rect 306974 211848 307083 211850
rect 306974 211792 307022 211848
rect 307078 211792 307083 211848
rect 306974 211787 307083 211792
rect 303846 211445 303906 211787
rect 306974 211581 307034 211787
rect 306925 211576 307034 211581
rect 306925 211520 306930 211576
rect 306986 211520 307034 211576
rect 306925 211518 307034 211520
rect 306925 211515 306991 211518
rect 303812 211440 303906 211445
rect 303812 211384 303817 211440
rect 303873 211384 303906 211440
rect 303812 211382 303906 211384
rect 303812 211379 303878 211382
rect 300760 211170 300826 211173
rect 302734 211170 302740 211172
rect 300760 211168 302740 211170
rect 300760 211112 300765 211168
rect 300821 211112 302740 211168
rect 300760 211110 302740 211112
rect 300760 211107 300826 211110
rect 302734 211108 302740 211110
rect 302804 211108 302810 211172
rect 294689 210490 294755 210493
rect 295374 210490 295380 210492
rect 294689 210488 295380 210490
rect 294689 210432 294694 210488
rect 294750 210432 295380 210488
rect 294689 210430 295380 210432
rect 294689 210427 294755 210430
rect 295374 210428 295380 210430
rect 295444 210428 295450 210492
rect 297725 210490 297791 210493
rect 298134 210490 298140 210492
rect 297725 210488 298140 210490
rect 297725 210432 297730 210488
rect 297786 210432 298140 210488
rect 297725 210430 298140 210432
rect 297725 210427 297791 210430
rect 298134 210428 298140 210430
rect 298204 210428 298210 210492
rect 580901 205730 580967 205733
rect 583520 205730 584960 205820
rect 580901 205728 584960 205730
rect 580901 205672 580906 205728
rect 580962 205672 584960 205728
rect 580901 205670 584960 205672
rect 580901 205667 580967 205670
rect 583520 205580 584960 205670
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 580441 165882 580507 165885
rect 583520 165882 584960 165972
rect 580441 165880 584960 165882
rect 580441 165824 580446 165880
rect 580502 165824 584960 165880
rect 580441 165822 584960 165824
rect 580441 165819 580507 165822
rect 583520 165732 584960 165822
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 580257 126034 580323 126037
rect 583520 126034 584960 126124
rect 580257 126032 584960 126034
rect 580257 125976 580262 126032
rect 580318 125976 584960 126032
rect 580257 125974 584960 125976
rect 580257 125971 580323 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 302918 86124 302924 86188
rect 302988 86186 302994 86188
rect 583520 86186 584960 86276
rect 302988 86126 584960 86186
rect 302988 86124 302994 86126
rect 583520 86036 584960 86126
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 298134 46276 298140 46340
rect 298204 46338 298210 46340
rect 583520 46338 584960 46428
rect 298204 46278 584960 46338
rect 298204 46276 298210 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 531814 19756 531820 19820
rect 531884 19818 531890 19820
rect 583520 19818 584960 19908
rect 531884 19758 584960 19818
rect 531884 19756 531890 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 295926 6564 295932 6628
rect 295996 6626 296002 6628
rect 583520 6626 584960 6716
rect 295996 6566 584960 6626
rect 295996 6564 296002 6566
rect 583520 6476 584960 6566
<< via3 >>
rect 294828 490648 294892 490652
rect 294828 490592 294834 490648
rect 294834 490592 294892 490648
rect 294828 490588 294892 490592
rect 297956 490648 298020 490652
rect 297956 490592 297990 490648
rect 297990 490592 298020 490648
rect 297956 490588 298020 490592
rect 301084 490648 301148 490652
rect 301084 490592 301089 490648
rect 301089 490592 301145 490648
rect 301145 490592 301148 490648
rect 301084 490588 301148 490592
rect 304212 490648 304276 490652
rect 304212 490592 304246 490648
rect 304246 490592 304276 490648
rect 304212 490588 304276 490592
rect 307340 490376 307404 490380
rect 307340 490320 307403 490376
rect 307403 490320 307404 490376
rect 307340 490316 307404 490320
rect 296484 487188 296548 487252
rect 306236 487188 306300 487252
rect 301268 451148 301332 451212
rect 304580 451148 304644 451212
rect 294460 450936 294524 450940
rect 294460 450880 294510 450936
rect 294510 450880 294524 450936
rect 294460 450876 294524 450880
rect 307708 450936 307772 450940
rect 307708 450880 307758 450936
rect 307758 450880 307772 450936
rect 307708 450876 307772 450880
rect 298140 450468 298204 450532
rect 296300 447204 296364 447268
rect 298140 431216 298204 431220
rect 298140 431160 298190 431216
rect 298190 431160 298204 431216
rect 298140 431156 298204 431160
rect 299244 431156 299308 431220
rect 294460 431020 294524 431084
rect 301452 431020 301516 431084
rect 308260 430884 308324 430948
rect 304764 430612 304828 430676
rect 306052 426396 306116 426460
rect 523540 421228 523604 421292
rect 526300 421228 526364 421292
rect 296484 421092 296548 421156
rect 296300 418372 296364 418436
rect 299244 411300 299308 411364
rect 531452 410892 531516 410956
rect 295196 410136 295260 410140
rect 295196 410080 295210 410136
rect 295210 410080 295260 410136
rect 295196 410076 295260 410080
rect 301636 410136 301700 410140
rect 301636 410080 301650 410136
rect 301650 410080 301700 410136
rect 301636 410076 301700 410080
rect 304764 410136 304828 410140
rect 304764 410080 304778 410136
rect 304778 410080 304828 410136
rect 304764 410076 304828 410080
rect 308260 410136 308324 410140
rect 308260 410080 308274 410136
rect 308274 410080 308324 410136
rect 308260 410076 308324 410080
rect 295196 391444 295260 391508
rect 299244 391504 299308 391508
rect 299244 391448 299258 391504
rect 299258 391448 299308 391504
rect 299244 391444 299308 391448
rect 298140 391232 298204 391236
rect 298140 391176 298190 391232
rect 298190 391176 298204 391232
rect 298140 391172 298204 391176
rect 301636 391232 301700 391236
rect 301636 391176 301650 391232
rect 301650 391176 301700 391232
rect 301636 391172 301700 391176
rect 304764 391036 304828 391100
rect 307708 391036 307772 391100
rect 304764 386820 304828 386884
rect 307524 386820 307588 386884
rect 523540 383692 523604 383756
rect 526300 383692 526364 383756
rect 531452 370908 531516 370972
rect 294460 370016 294524 370020
rect 294460 369960 294510 370016
rect 294510 369960 294524 370016
rect 294460 369956 294524 369960
rect 298140 369956 298204 370020
rect 300716 370016 300780 370020
rect 300716 369960 300766 370016
rect 300766 369960 300780 370016
rect 300716 369956 300780 369960
rect 304212 370016 304276 370020
rect 304212 369960 304226 370016
rect 304226 369960 304276 370016
rect 304212 369956 304276 369960
rect 306972 370016 307036 370020
rect 306972 369960 306986 370016
rect 306986 369960 307036 370016
rect 306972 369956 307036 369960
rect 527036 351868 527100 351932
rect 523540 341260 523604 341324
rect 526300 341260 526364 341324
rect 304764 334188 304828 334252
rect 531452 330924 531516 330988
rect 526300 303588 526364 303652
rect 523540 302228 523604 302292
rect 524276 302228 524340 302292
rect 306236 301004 306300 301068
rect 306052 296924 306116 296988
rect 307524 294204 307588 294268
rect 304212 291484 304276 291548
rect 304764 291484 304828 291548
rect 300164 291408 300228 291412
rect 300164 291352 300178 291408
rect 300178 291352 300228 291408
rect 300164 291348 300228 291352
rect 306788 291408 306852 291412
rect 306788 291352 306802 291408
rect 306802 291352 306852 291408
rect 306788 291348 306852 291352
rect 294460 291212 294524 291276
rect 298140 291272 298204 291276
rect 298140 291216 298154 291272
rect 298154 291216 298204 291272
rect 298140 291212 298204 291216
rect 299244 291212 299308 291276
rect 531452 290940 531516 291004
rect 300900 271764 300964 271828
rect 307708 271628 307772 271692
rect 294644 271552 294708 271556
rect 294644 271496 294694 271552
rect 294694 271496 294708 271552
rect 294644 271492 294708 271496
rect 299244 271492 299308 271556
rect 301452 271552 301516 271556
rect 301452 271496 301466 271552
rect 301466 271496 301516 271552
rect 301452 271492 301516 271496
rect 304948 271552 305012 271556
rect 304948 271496 304998 271552
rect 304998 271496 305012 271552
rect 304948 271492 305012 271496
rect 308260 271552 308324 271556
rect 308260 271496 308310 271552
rect 308310 271496 308324 271552
rect 308260 271492 308324 271496
rect 524276 264556 524340 264620
rect 526300 264556 526364 264620
rect 299244 251500 299308 251564
rect 301452 251560 301516 251564
rect 301452 251504 301466 251560
rect 301466 251504 301516 251560
rect 301452 251500 301516 251504
rect 302740 251500 302804 251564
rect 308260 251560 308324 251564
rect 308260 251504 308274 251560
rect 308274 251504 308324 251560
rect 308260 251500 308324 251504
rect 295380 251364 295444 251428
rect 304948 250956 305012 251020
rect 531452 250956 531516 251020
rect 309732 233276 309796 233340
rect 295380 231432 295444 231436
rect 295380 231376 295394 231432
rect 295394 231376 295444 231432
rect 295380 231372 295444 231376
rect 299244 231372 299308 231436
rect 302924 230556 302988 230620
rect 306420 230616 306484 230620
rect 306420 230560 306457 230616
rect 306457 230560 306484 230616
rect 306420 230556 306484 230560
rect 309732 230556 309796 230620
rect 298140 230148 298204 230212
rect 309732 213284 309796 213348
rect 306420 213148 306484 213212
rect 302740 211108 302804 211172
rect 295380 210428 295444 210492
rect 298140 210428 298204 210492
rect 302924 86124 302988 86188
rect 298140 46276 298204 46340
rect 531820 19756 531884 19820
rect 295932 6564 295996 6628
<< metal4 >>
rect -3236 705918 -2636 706100
rect -3236 705682 -3054 705918
rect -2818 705682 -2636 705918
rect -3236 675494 -2636 705682
rect -3236 675258 -3054 675494
rect -2818 675258 -2636 675494
rect -3236 638294 -2636 675258
rect -3236 638058 -3054 638294
rect -2818 638058 -2636 638294
rect -3236 601094 -2636 638058
rect -3236 600858 -3054 601094
rect -2818 600858 -2636 601094
rect -3236 563894 -2636 600858
rect -3236 563658 -3054 563894
rect -2818 563658 -2636 563894
rect -3236 526694 -2636 563658
rect -3236 526458 -3054 526694
rect -2818 526458 -2636 526694
rect -3236 489494 -2636 526458
rect -3236 489258 -3054 489494
rect -2818 489258 -2636 489494
rect -3236 452294 -2636 489258
rect -3236 452058 -3054 452294
rect -2818 452058 -2636 452294
rect -3236 415094 -2636 452058
rect -3236 414858 -3054 415094
rect -2818 414858 -2636 415094
rect -3236 377894 -2636 414858
rect -3236 377658 -3054 377894
rect -2818 377658 -2636 377894
rect -3236 340694 -2636 377658
rect -3236 340458 -3054 340694
rect -2818 340458 -2636 340694
rect -3236 303494 -2636 340458
rect -3236 303258 -3054 303494
rect -2818 303258 -2636 303494
rect -3236 266294 -2636 303258
rect -3236 266058 -3054 266294
rect -2818 266058 -2636 266294
rect -3236 229094 -2636 266058
rect -3236 228858 -3054 229094
rect -2818 228858 -2636 229094
rect -3236 191894 -2636 228858
rect -3236 191658 -3054 191894
rect -2818 191658 -2636 191894
rect -3236 154694 -2636 191658
rect -3236 154458 -3054 154694
rect -2818 154458 -2636 154694
rect -3236 117494 -2636 154458
rect -3236 117258 -3054 117494
rect -2818 117258 -2636 117494
rect -3236 80294 -2636 117258
rect -3236 80058 -3054 80294
rect -2818 80058 -2636 80294
rect -3236 43094 -2636 80058
rect -3236 42858 -3054 43094
rect -2818 42858 -2636 43094
rect -3236 5894 -2636 42858
rect -3236 5658 -3054 5894
rect -2818 5658 -2636 5894
rect -3236 -1746 -2636 5658
rect -2296 704978 -1696 705160
rect -2296 704742 -2114 704978
rect -1878 704742 -1696 704978
rect -2296 671894 -1696 704742
rect -2296 671658 -2114 671894
rect -1878 671658 -1696 671894
rect -2296 634694 -1696 671658
rect -2296 634458 -2114 634694
rect -1878 634458 -1696 634694
rect -2296 597494 -1696 634458
rect -2296 597258 -2114 597494
rect -1878 597258 -1696 597494
rect -2296 560294 -1696 597258
rect -2296 560058 -2114 560294
rect -1878 560058 -1696 560294
rect -2296 523094 -1696 560058
rect -2296 522858 -2114 523094
rect -1878 522858 -1696 523094
rect -2296 485894 -1696 522858
rect -2296 485658 -2114 485894
rect -1878 485658 -1696 485894
rect -2296 448694 -1696 485658
rect -2296 448458 -2114 448694
rect -1878 448458 -1696 448694
rect -2296 411494 -1696 448458
rect -2296 411258 -2114 411494
rect -1878 411258 -1696 411494
rect -2296 374294 -1696 411258
rect -2296 374058 -2114 374294
rect -1878 374058 -1696 374294
rect -2296 337094 -1696 374058
rect -2296 336858 -2114 337094
rect -1878 336858 -1696 337094
rect -2296 299894 -1696 336858
rect -2296 299658 -2114 299894
rect -1878 299658 -1696 299894
rect -2296 262694 -1696 299658
rect -2296 262458 -2114 262694
rect -1878 262458 -1696 262694
rect -2296 225494 -1696 262458
rect -2296 225258 -2114 225494
rect -1878 225258 -1696 225494
rect -2296 188294 -1696 225258
rect -2296 188058 -2114 188294
rect -1878 188058 -1696 188294
rect -2296 151094 -1696 188058
rect -2296 150858 -2114 151094
rect -1878 150858 -1696 151094
rect -2296 113894 -1696 150858
rect -2296 113658 -2114 113894
rect -1878 113658 -1696 113894
rect -2296 76694 -1696 113658
rect -2296 76458 -2114 76694
rect -1878 76458 -1696 76694
rect -2296 39494 -1696 76458
rect -2296 39258 -2114 39494
rect -1878 39258 -1696 39494
rect -2296 2294 -1696 39258
rect -2296 2058 -2114 2294
rect -1878 2058 -1696 2294
rect -2296 -806 -1696 2058
rect -2296 -1042 -2114 -806
rect -1878 -1042 -1696 -806
rect -2296 -1224 -1696 -1042
rect 804 704978 1404 706100
rect 804 704742 986 704978
rect 1222 704742 1404 704978
rect 804 671894 1404 704742
rect 804 671658 986 671894
rect 1222 671658 1404 671894
rect 804 634694 1404 671658
rect 804 634458 986 634694
rect 1222 634458 1404 634694
rect 804 597494 1404 634458
rect 804 597258 986 597494
rect 1222 597258 1404 597494
rect 804 560294 1404 597258
rect 804 560058 986 560294
rect 1222 560058 1404 560294
rect 804 523094 1404 560058
rect 804 522858 986 523094
rect 1222 522858 1404 523094
rect 804 485894 1404 522858
rect 804 485658 986 485894
rect 1222 485658 1404 485894
rect 804 448694 1404 485658
rect 804 448458 986 448694
rect 1222 448458 1404 448694
rect 804 411494 1404 448458
rect 804 411258 986 411494
rect 1222 411258 1404 411494
rect 804 374294 1404 411258
rect 804 374058 986 374294
rect 1222 374058 1404 374294
rect 804 337094 1404 374058
rect 804 336858 986 337094
rect 1222 336858 1404 337094
rect 804 299894 1404 336858
rect 804 299658 986 299894
rect 1222 299658 1404 299894
rect 804 262694 1404 299658
rect 804 262458 986 262694
rect 1222 262458 1404 262694
rect 804 225494 1404 262458
rect 804 225258 986 225494
rect 1222 225258 1404 225494
rect 804 188294 1404 225258
rect 804 188058 986 188294
rect 1222 188058 1404 188294
rect 804 151094 1404 188058
rect 804 150858 986 151094
rect 1222 150858 1404 151094
rect 804 113894 1404 150858
rect 804 113658 986 113894
rect 1222 113658 1404 113894
rect 804 76694 1404 113658
rect 804 76458 986 76694
rect 1222 76458 1404 76694
rect 804 39494 1404 76458
rect 804 39258 986 39494
rect 1222 39258 1404 39494
rect 804 2294 1404 39258
rect 804 2058 986 2294
rect 1222 2058 1404 2294
rect 804 -806 1404 2058
rect 804 -1042 986 -806
rect 1222 -1042 1404 -806
rect -3236 -1982 -3054 -1746
rect -2818 -1982 -2636 -1746
rect -3236 -2164 -2636 -1982
rect 804 -2164 1404 -1042
rect 4404 705918 5004 706100
rect 4404 705682 4586 705918
rect 4822 705682 5004 705918
rect 4404 675494 5004 705682
rect 4404 675258 4586 675494
rect 4822 675258 5004 675494
rect 4404 638294 5004 675258
rect 4404 638058 4586 638294
rect 4822 638058 5004 638294
rect 4404 601094 5004 638058
rect 4404 600858 4586 601094
rect 4822 600858 5004 601094
rect 4404 563894 5004 600858
rect 4404 563658 4586 563894
rect 4822 563658 5004 563894
rect 4404 526694 5004 563658
rect 4404 526458 4586 526694
rect 4822 526458 5004 526694
rect 4404 489494 5004 526458
rect 4404 489258 4586 489494
rect 4822 489258 5004 489494
rect 4404 452294 5004 489258
rect 4404 452058 4586 452294
rect 4822 452058 5004 452294
rect 4404 415094 5004 452058
rect 4404 414858 4586 415094
rect 4822 414858 5004 415094
rect 4404 377894 5004 414858
rect 4404 377658 4586 377894
rect 4822 377658 5004 377894
rect 4404 340694 5004 377658
rect 4404 340458 4586 340694
rect 4822 340458 5004 340694
rect 4404 303494 5004 340458
rect 4404 303258 4586 303494
rect 4822 303258 5004 303494
rect 4404 266294 5004 303258
rect 4404 266058 4586 266294
rect 4822 266058 5004 266294
rect 4404 229094 5004 266058
rect 4404 228858 4586 229094
rect 4822 228858 5004 229094
rect 4404 191894 5004 228858
rect 4404 191658 4586 191894
rect 4822 191658 5004 191894
rect 4404 154694 5004 191658
rect 4404 154458 4586 154694
rect 4822 154458 5004 154694
rect 4404 117494 5004 154458
rect 4404 117258 4586 117494
rect 4822 117258 5004 117494
rect 4404 80294 5004 117258
rect 4404 80058 4586 80294
rect 4822 80058 5004 80294
rect 4404 43094 5004 80058
rect 4404 42858 4586 43094
rect 4822 42858 5004 43094
rect 4404 5894 5004 42858
rect 4404 5658 4586 5894
rect 4822 5658 5004 5894
rect 4404 -1746 5004 5658
rect 4404 -1982 4586 -1746
rect 4822 -1982 5004 -1746
rect 4404 -2164 5004 -1982
rect 38004 704978 38604 706100
rect 38004 704742 38186 704978
rect 38422 704742 38604 704978
rect 38004 671894 38604 704742
rect 38004 671658 38186 671894
rect 38422 671658 38604 671894
rect 38004 634694 38604 671658
rect 38004 634458 38186 634694
rect 38422 634458 38604 634694
rect 38004 597494 38604 634458
rect 38004 597258 38186 597494
rect 38422 597258 38604 597494
rect 38004 560294 38604 597258
rect 38004 560058 38186 560294
rect 38422 560058 38604 560294
rect 38004 523094 38604 560058
rect 38004 522858 38186 523094
rect 38422 522858 38604 523094
rect 38004 485894 38604 522858
rect 38004 485658 38186 485894
rect 38422 485658 38604 485894
rect 38004 448694 38604 485658
rect 38004 448458 38186 448694
rect 38422 448458 38604 448694
rect 38004 411494 38604 448458
rect 38004 411258 38186 411494
rect 38422 411258 38604 411494
rect 38004 374294 38604 411258
rect 38004 374058 38186 374294
rect 38422 374058 38604 374294
rect 38004 337094 38604 374058
rect 38004 336858 38186 337094
rect 38422 336858 38604 337094
rect 38004 299894 38604 336858
rect 38004 299658 38186 299894
rect 38422 299658 38604 299894
rect 38004 262694 38604 299658
rect 38004 262458 38186 262694
rect 38422 262458 38604 262694
rect 38004 225494 38604 262458
rect 38004 225258 38186 225494
rect 38422 225258 38604 225494
rect 38004 188294 38604 225258
rect 38004 188058 38186 188294
rect 38422 188058 38604 188294
rect 38004 151094 38604 188058
rect 38004 150858 38186 151094
rect 38422 150858 38604 151094
rect 38004 113894 38604 150858
rect 38004 113658 38186 113894
rect 38422 113658 38604 113894
rect 38004 76694 38604 113658
rect 38004 76458 38186 76694
rect 38422 76458 38604 76694
rect 38004 39494 38604 76458
rect 38004 39258 38186 39494
rect 38422 39258 38604 39494
rect 38004 2294 38604 39258
rect 38004 2058 38186 2294
rect 38422 2058 38604 2294
rect 38004 -806 38604 2058
rect 38004 -1042 38186 -806
rect 38422 -1042 38604 -806
rect 38004 -2164 38604 -1042
rect 41604 705918 42204 706100
rect 41604 705682 41786 705918
rect 42022 705682 42204 705918
rect 41604 675494 42204 705682
rect 41604 675258 41786 675494
rect 42022 675258 42204 675494
rect 41604 638294 42204 675258
rect 41604 638058 41786 638294
rect 42022 638058 42204 638294
rect 41604 601094 42204 638058
rect 41604 600858 41786 601094
rect 42022 600858 42204 601094
rect 41604 563894 42204 600858
rect 41604 563658 41786 563894
rect 42022 563658 42204 563894
rect 41604 526694 42204 563658
rect 41604 526458 41786 526694
rect 42022 526458 42204 526694
rect 41604 489494 42204 526458
rect 41604 489258 41786 489494
rect 42022 489258 42204 489494
rect 41604 452294 42204 489258
rect 41604 452058 41786 452294
rect 42022 452058 42204 452294
rect 41604 415094 42204 452058
rect 41604 414858 41786 415094
rect 42022 414858 42204 415094
rect 41604 377894 42204 414858
rect 41604 377658 41786 377894
rect 42022 377658 42204 377894
rect 41604 340694 42204 377658
rect 41604 340458 41786 340694
rect 42022 340458 42204 340694
rect 41604 303494 42204 340458
rect 41604 303258 41786 303494
rect 42022 303258 42204 303494
rect 41604 266294 42204 303258
rect 41604 266058 41786 266294
rect 42022 266058 42204 266294
rect 41604 229094 42204 266058
rect 41604 228858 41786 229094
rect 42022 228858 42204 229094
rect 41604 191894 42204 228858
rect 41604 191658 41786 191894
rect 42022 191658 42204 191894
rect 41604 154694 42204 191658
rect 41604 154458 41786 154694
rect 42022 154458 42204 154694
rect 41604 117494 42204 154458
rect 41604 117258 41786 117494
rect 42022 117258 42204 117494
rect 41604 80294 42204 117258
rect 41604 80058 41786 80294
rect 42022 80058 42204 80294
rect 41604 43094 42204 80058
rect 41604 42858 41786 43094
rect 42022 42858 42204 43094
rect 41604 5894 42204 42858
rect 41604 5658 41786 5894
rect 42022 5658 42204 5894
rect 41604 -1746 42204 5658
rect 41604 -1982 41786 -1746
rect 42022 -1982 42204 -1746
rect 41604 -2164 42204 -1982
rect 75204 704978 75804 706100
rect 75204 704742 75386 704978
rect 75622 704742 75804 704978
rect 75204 671894 75804 704742
rect 75204 671658 75386 671894
rect 75622 671658 75804 671894
rect 75204 634694 75804 671658
rect 75204 634458 75386 634694
rect 75622 634458 75804 634694
rect 75204 597494 75804 634458
rect 75204 597258 75386 597494
rect 75622 597258 75804 597494
rect 75204 560294 75804 597258
rect 75204 560058 75386 560294
rect 75622 560058 75804 560294
rect 75204 523094 75804 560058
rect 75204 522858 75386 523094
rect 75622 522858 75804 523094
rect 75204 485894 75804 522858
rect 75204 485658 75386 485894
rect 75622 485658 75804 485894
rect 75204 448694 75804 485658
rect 75204 448458 75386 448694
rect 75622 448458 75804 448694
rect 75204 411494 75804 448458
rect 75204 411258 75386 411494
rect 75622 411258 75804 411494
rect 75204 374294 75804 411258
rect 75204 374058 75386 374294
rect 75622 374058 75804 374294
rect 75204 337094 75804 374058
rect 75204 336858 75386 337094
rect 75622 336858 75804 337094
rect 75204 299894 75804 336858
rect 75204 299658 75386 299894
rect 75622 299658 75804 299894
rect 75204 262694 75804 299658
rect 75204 262458 75386 262694
rect 75622 262458 75804 262694
rect 75204 225494 75804 262458
rect 75204 225258 75386 225494
rect 75622 225258 75804 225494
rect 75204 188294 75804 225258
rect 75204 188058 75386 188294
rect 75622 188058 75804 188294
rect 75204 151094 75804 188058
rect 75204 150858 75386 151094
rect 75622 150858 75804 151094
rect 75204 113894 75804 150858
rect 75204 113658 75386 113894
rect 75622 113658 75804 113894
rect 75204 76694 75804 113658
rect 75204 76458 75386 76694
rect 75622 76458 75804 76694
rect 75204 39494 75804 76458
rect 75204 39258 75386 39494
rect 75622 39258 75804 39494
rect 75204 2294 75804 39258
rect 75204 2058 75386 2294
rect 75622 2058 75804 2294
rect 75204 -806 75804 2058
rect 75204 -1042 75386 -806
rect 75622 -1042 75804 -806
rect 75204 -2164 75804 -1042
rect 78804 705918 79404 706100
rect 78804 705682 78986 705918
rect 79222 705682 79404 705918
rect 78804 675494 79404 705682
rect 78804 675258 78986 675494
rect 79222 675258 79404 675494
rect 78804 638294 79404 675258
rect 78804 638058 78986 638294
rect 79222 638058 79404 638294
rect 78804 601094 79404 638058
rect 78804 600858 78986 601094
rect 79222 600858 79404 601094
rect 78804 563894 79404 600858
rect 78804 563658 78986 563894
rect 79222 563658 79404 563894
rect 78804 526694 79404 563658
rect 78804 526458 78986 526694
rect 79222 526458 79404 526694
rect 78804 489494 79404 526458
rect 78804 489258 78986 489494
rect 79222 489258 79404 489494
rect 78804 452294 79404 489258
rect 78804 452058 78986 452294
rect 79222 452058 79404 452294
rect 78804 415094 79404 452058
rect 78804 414858 78986 415094
rect 79222 414858 79404 415094
rect 78804 377894 79404 414858
rect 78804 377658 78986 377894
rect 79222 377658 79404 377894
rect 78804 340694 79404 377658
rect 78804 340458 78986 340694
rect 79222 340458 79404 340694
rect 78804 303494 79404 340458
rect 78804 303258 78986 303494
rect 79222 303258 79404 303494
rect 78804 266294 79404 303258
rect 78804 266058 78986 266294
rect 79222 266058 79404 266294
rect 78804 229094 79404 266058
rect 78804 228858 78986 229094
rect 79222 228858 79404 229094
rect 78804 191894 79404 228858
rect 78804 191658 78986 191894
rect 79222 191658 79404 191894
rect 78804 154694 79404 191658
rect 78804 154458 78986 154694
rect 79222 154458 79404 154694
rect 78804 117494 79404 154458
rect 78804 117258 78986 117494
rect 79222 117258 79404 117494
rect 78804 80294 79404 117258
rect 78804 80058 78986 80294
rect 79222 80058 79404 80294
rect 78804 43094 79404 80058
rect 78804 42858 78986 43094
rect 79222 42858 79404 43094
rect 78804 5894 79404 42858
rect 78804 5658 78986 5894
rect 79222 5658 79404 5894
rect 78804 -1746 79404 5658
rect 78804 -1982 78986 -1746
rect 79222 -1982 79404 -1746
rect 78804 -2164 79404 -1982
rect 112404 704978 113004 706100
rect 112404 704742 112586 704978
rect 112822 704742 113004 704978
rect 112404 671894 113004 704742
rect 112404 671658 112586 671894
rect 112822 671658 113004 671894
rect 112404 634694 113004 671658
rect 112404 634458 112586 634694
rect 112822 634458 113004 634694
rect 112404 597494 113004 634458
rect 112404 597258 112586 597494
rect 112822 597258 113004 597494
rect 112404 560294 113004 597258
rect 112404 560058 112586 560294
rect 112822 560058 113004 560294
rect 112404 523094 113004 560058
rect 112404 522858 112586 523094
rect 112822 522858 113004 523094
rect 112404 485894 113004 522858
rect 112404 485658 112586 485894
rect 112822 485658 113004 485894
rect 112404 448694 113004 485658
rect 112404 448458 112586 448694
rect 112822 448458 113004 448694
rect 112404 411494 113004 448458
rect 112404 411258 112586 411494
rect 112822 411258 113004 411494
rect 112404 374294 113004 411258
rect 112404 374058 112586 374294
rect 112822 374058 113004 374294
rect 112404 337094 113004 374058
rect 112404 336858 112586 337094
rect 112822 336858 113004 337094
rect 112404 299894 113004 336858
rect 112404 299658 112586 299894
rect 112822 299658 113004 299894
rect 112404 262694 113004 299658
rect 112404 262458 112586 262694
rect 112822 262458 113004 262694
rect 112404 225494 113004 262458
rect 112404 225258 112586 225494
rect 112822 225258 113004 225494
rect 112404 188294 113004 225258
rect 112404 188058 112586 188294
rect 112822 188058 113004 188294
rect 112404 151094 113004 188058
rect 112404 150858 112586 151094
rect 112822 150858 113004 151094
rect 112404 113894 113004 150858
rect 112404 113658 112586 113894
rect 112822 113658 113004 113894
rect 112404 76694 113004 113658
rect 112404 76458 112586 76694
rect 112822 76458 113004 76694
rect 112404 39494 113004 76458
rect 112404 39258 112586 39494
rect 112822 39258 113004 39494
rect 112404 2294 113004 39258
rect 112404 2058 112586 2294
rect 112822 2058 113004 2294
rect 112404 -806 113004 2058
rect 112404 -1042 112586 -806
rect 112822 -1042 113004 -806
rect 112404 -2164 113004 -1042
rect 116004 705918 116604 706100
rect 116004 705682 116186 705918
rect 116422 705682 116604 705918
rect 116004 675494 116604 705682
rect 116004 675258 116186 675494
rect 116422 675258 116604 675494
rect 116004 638294 116604 675258
rect 116004 638058 116186 638294
rect 116422 638058 116604 638294
rect 116004 601094 116604 638058
rect 116004 600858 116186 601094
rect 116422 600858 116604 601094
rect 116004 563894 116604 600858
rect 116004 563658 116186 563894
rect 116422 563658 116604 563894
rect 116004 526694 116604 563658
rect 116004 526458 116186 526694
rect 116422 526458 116604 526694
rect 116004 489494 116604 526458
rect 116004 489258 116186 489494
rect 116422 489258 116604 489494
rect 116004 452294 116604 489258
rect 116004 452058 116186 452294
rect 116422 452058 116604 452294
rect 116004 415094 116604 452058
rect 116004 414858 116186 415094
rect 116422 414858 116604 415094
rect 116004 377894 116604 414858
rect 116004 377658 116186 377894
rect 116422 377658 116604 377894
rect 116004 340694 116604 377658
rect 116004 340458 116186 340694
rect 116422 340458 116604 340694
rect 116004 303494 116604 340458
rect 116004 303258 116186 303494
rect 116422 303258 116604 303494
rect 116004 266294 116604 303258
rect 116004 266058 116186 266294
rect 116422 266058 116604 266294
rect 116004 229094 116604 266058
rect 116004 228858 116186 229094
rect 116422 228858 116604 229094
rect 116004 191894 116604 228858
rect 116004 191658 116186 191894
rect 116422 191658 116604 191894
rect 116004 154694 116604 191658
rect 116004 154458 116186 154694
rect 116422 154458 116604 154694
rect 116004 117494 116604 154458
rect 116004 117258 116186 117494
rect 116422 117258 116604 117494
rect 116004 80294 116604 117258
rect 116004 80058 116186 80294
rect 116422 80058 116604 80294
rect 116004 43094 116604 80058
rect 116004 42858 116186 43094
rect 116422 42858 116604 43094
rect 116004 5894 116604 42858
rect 116004 5658 116186 5894
rect 116422 5658 116604 5894
rect 116004 -1746 116604 5658
rect 116004 -1982 116186 -1746
rect 116422 -1982 116604 -1746
rect 116004 -2164 116604 -1982
rect 149604 704978 150204 706100
rect 149604 704742 149786 704978
rect 150022 704742 150204 704978
rect 149604 671894 150204 704742
rect 149604 671658 149786 671894
rect 150022 671658 150204 671894
rect 149604 634694 150204 671658
rect 149604 634458 149786 634694
rect 150022 634458 150204 634694
rect 149604 597494 150204 634458
rect 149604 597258 149786 597494
rect 150022 597258 150204 597494
rect 149604 560294 150204 597258
rect 149604 560058 149786 560294
rect 150022 560058 150204 560294
rect 149604 523094 150204 560058
rect 149604 522858 149786 523094
rect 150022 522858 150204 523094
rect 149604 485894 150204 522858
rect 149604 485658 149786 485894
rect 150022 485658 150204 485894
rect 149604 448694 150204 485658
rect 149604 448458 149786 448694
rect 150022 448458 150204 448694
rect 149604 411494 150204 448458
rect 149604 411258 149786 411494
rect 150022 411258 150204 411494
rect 149604 374294 150204 411258
rect 149604 374058 149786 374294
rect 150022 374058 150204 374294
rect 149604 337094 150204 374058
rect 149604 336858 149786 337094
rect 150022 336858 150204 337094
rect 149604 299894 150204 336858
rect 149604 299658 149786 299894
rect 150022 299658 150204 299894
rect 149604 262694 150204 299658
rect 149604 262458 149786 262694
rect 150022 262458 150204 262694
rect 149604 225494 150204 262458
rect 149604 225258 149786 225494
rect 150022 225258 150204 225494
rect 149604 188294 150204 225258
rect 149604 188058 149786 188294
rect 150022 188058 150204 188294
rect 149604 151094 150204 188058
rect 149604 150858 149786 151094
rect 150022 150858 150204 151094
rect 149604 113894 150204 150858
rect 149604 113658 149786 113894
rect 150022 113658 150204 113894
rect 149604 76694 150204 113658
rect 149604 76458 149786 76694
rect 150022 76458 150204 76694
rect 149604 39494 150204 76458
rect 149604 39258 149786 39494
rect 150022 39258 150204 39494
rect 149604 2294 150204 39258
rect 149604 2058 149786 2294
rect 150022 2058 150204 2294
rect 149604 -806 150204 2058
rect 149604 -1042 149786 -806
rect 150022 -1042 150204 -806
rect 149604 -2164 150204 -1042
rect 153204 705918 153804 706100
rect 153204 705682 153386 705918
rect 153622 705682 153804 705918
rect 153204 675494 153804 705682
rect 153204 675258 153386 675494
rect 153622 675258 153804 675494
rect 153204 638294 153804 675258
rect 153204 638058 153386 638294
rect 153622 638058 153804 638294
rect 153204 601094 153804 638058
rect 153204 600858 153386 601094
rect 153622 600858 153804 601094
rect 153204 563894 153804 600858
rect 153204 563658 153386 563894
rect 153622 563658 153804 563894
rect 153204 526694 153804 563658
rect 153204 526458 153386 526694
rect 153622 526458 153804 526694
rect 153204 489494 153804 526458
rect 153204 489258 153386 489494
rect 153622 489258 153804 489494
rect 153204 452294 153804 489258
rect 153204 452058 153386 452294
rect 153622 452058 153804 452294
rect 153204 415094 153804 452058
rect 153204 414858 153386 415094
rect 153622 414858 153804 415094
rect 153204 377894 153804 414858
rect 153204 377658 153386 377894
rect 153622 377658 153804 377894
rect 153204 340694 153804 377658
rect 153204 340458 153386 340694
rect 153622 340458 153804 340694
rect 153204 303494 153804 340458
rect 153204 303258 153386 303494
rect 153622 303258 153804 303494
rect 153204 266294 153804 303258
rect 153204 266058 153386 266294
rect 153622 266058 153804 266294
rect 153204 229094 153804 266058
rect 153204 228858 153386 229094
rect 153622 228858 153804 229094
rect 153204 191894 153804 228858
rect 153204 191658 153386 191894
rect 153622 191658 153804 191894
rect 153204 154694 153804 191658
rect 153204 154458 153386 154694
rect 153622 154458 153804 154694
rect 153204 117494 153804 154458
rect 153204 117258 153386 117494
rect 153622 117258 153804 117494
rect 153204 80294 153804 117258
rect 153204 80058 153386 80294
rect 153622 80058 153804 80294
rect 153204 43094 153804 80058
rect 153204 42858 153386 43094
rect 153622 42858 153804 43094
rect 153204 5894 153804 42858
rect 153204 5658 153386 5894
rect 153622 5658 153804 5894
rect 153204 -1746 153804 5658
rect 153204 -1982 153386 -1746
rect 153622 -1982 153804 -1746
rect 153204 -2164 153804 -1982
rect 186804 704978 187404 706100
rect 186804 704742 186986 704978
rect 187222 704742 187404 704978
rect 186804 671894 187404 704742
rect 186804 671658 186986 671894
rect 187222 671658 187404 671894
rect 186804 634694 187404 671658
rect 186804 634458 186986 634694
rect 187222 634458 187404 634694
rect 186804 597494 187404 634458
rect 186804 597258 186986 597494
rect 187222 597258 187404 597494
rect 186804 560294 187404 597258
rect 186804 560058 186986 560294
rect 187222 560058 187404 560294
rect 186804 523094 187404 560058
rect 186804 522858 186986 523094
rect 187222 522858 187404 523094
rect 186804 485894 187404 522858
rect 186804 485658 186986 485894
rect 187222 485658 187404 485894
rect 186804 448694 187404 485658
rect 186804 448458 186986 448694
rect 187222 448458 187404 448694
rect 186804 411494 187404 448458
rect 186804 411258 186986 411494
rect 187222 411258 187404 411494
rect 186804 374294 187404 411258
rect 186804 374058 186986 374294
rect 187222 374058 187404 374294
rect 186804 337094 187404 374058
rect 186804 336858 186986 337094
rect 187222 336858 187404 337094
rect 186804 299894 187404 336858
rect 186804 299658 186986 299894
rect 187222 299658 187404 299894
rect 186804 262694 187404 299658
rect 186804 262458 186986 262694
rect 187222 262458 187404 262694
rect 186804 225494 187404 262458
rect 186804 225258 186986 225494
rect 187222 225258 187404 225494
rect 186804 188294 187404 225258
rect 186804 188058 186986 188294
rect 187222 188058 187404 188294
rect 186804 151094 187404 188058
rect 186804 150858 186986 151094
rect 187222 150858 187404 151094
rect 186804 113894 187404 150858
rect 186804 113658 186986 113894
rect 187222 113658 187404 113894
rect 186804 76694 187404 113658
rect 186804 76458 186986 76694
rect 187222 76458 187404 76694
rect 186804 39494 187404 76458
rect 186804 39258 186986 39494
rect 187222 39258 187404 39494
rect 186804 2294 187404 39258
rect 186804 2058 186986 2294
rect 187222 2058 187404 2294
rect 186804 -806 187404 2058
rect 186804 -1042 186986 -806
rect 187222 -1042 187404 -806
rect 186804 -2164 187404 -1042
rect 190404 705918 191004 706100
rect 190404 705682 190586 705918
rect 190822 705682 191004 705918
rect 190404 675494 191004 705682
rect 190404 675258 190586 675494
rect 190822 675258 191004 675494
rect 190404 638294 191004 675258
rect 190404 638058 190586 638294
rect 190822 638058 191004 638294
rect 190404 601094 191004 638058
rect 190404 600858 190586 601094
rect 190822 600858 191004 601094
rect 190404 563894 191004 600858
rect 190404 563658 190586 563894
rect 190822 563658 191004 563894
rect 190404 526694 191004 563658
rect 190404 526458 190586 526694
rect 190822 526458 191004 526694
rect 190404 489494 191004 526458
rect 190404 489258 190586 489494
rect 190822 489258 191004 489494
rect 190404 452294 191004 489258
rect 190404 452058 190586 452294
rect 190822 452058 191004 452294
rect 190404 415094 191004 452058
rect 190404 414858 190586 415094
rect 190822 414858 191004 415094
rect 190404 377894 191004 414858
rect 190404 377658 190586 377894
rect 190822 377658 191004 377894
rect 190404 340694 191004 377658
rect 190404 340458 190586 340694
rect 190822 340458 191004 340694
rect 190404 303494 191004 340458
rect 190404 303258 190586 303494
rect 190822 303258 191004 303494
rect 190404 266294 191004 303258
rect 190404 266058 190586 266294
rect 190822 266058 191004 266294
rect 190404 229094 191004 266058
rect 190404 228858 190586 229094
rect 190822 228858 191004 229094
rect 190404 191894 191004 228858
rect 190404 191658 190586 191894
rect 190822 191658 191004 191894
rect 190404 154694 191004 191658
rect 190404 154458 190586 154694
rect 190822 154458 191004 154694
rect 190404 117494 191004 154458
rect 190404 117258 190586 117494
rect 190822 117258 191004 117494
rect 190404 80294 191004 117258
rect 190404 80058 190586 80294
rect 190822 80058 191004 80294
rect 190404 43094 191004 80058
rect 190404 42858 190586 43094
rect 190822 42858 191004 43094
rect 190404 5894 191004 42858
rect 190404 5658 190586 5894
rect 190822 5658 191004 5894
rect 190404 -1746 191004 5658
rect 190404 -1982 190586 -1746
rect 190822 -1982 191004 -1746
rect 190404 -2164 191004 -1982
rect 224004 704978 224604 706100
rect 224004 704742 224186 704978
rect 224422 704742 224604 704978
rect 224004 671894 224604 704742
rect 224004 671658 224186 671894
rect 224422 671658 224604 671894
rect 224004 634694 224604 671658
rect 224004 634458 224186 634694
rect 224422 634458 224604 634694
rect 224004 597494 224604 634458
rect 224004 597258 224186 597494
rect 224422 597258 224604 597494
rect 224004 560294 224604 597258
rect 224004 560058 224186 560294
rect 224422 560058 224604 560294
rect 224004 523094 224604 560058
rect 224004 522858 224186 523094
rect 224422 522858 224604 523094
rect 224004 485894 224604 522858
rect 224004 485658 224186 485894
rect 224422 485658 224604 485894
rect 224004 448694 224604 485658
rect 224004 448458 224186 448694
rect 224422 448458 224604 448694
rect 224004 411494 224604 448458
rect 224004 411258 224186 411494
rect 224422 411258 224604 411494
rect 224004 374294 224604 411258
rect 224004 374058 224186 374294
rect 224422 374058 224604 374294
rect 224004 337094 224604 374058
rect 224004 336858 224186 337094
rect 224422 336858 224604 337094
rect 224004 299894 224604 336858
rect 224004 299658 224186 299894
rect 224422 299658 224604 299894
rect 224004 262694 224604 299658
rect 224004 262458 224186 262694
rect 224422 262458 224604 262694
rect 224004 225494 224604 262458
rect 224004 225258 224186 225494
rect 224422 225258 224604 225494
rect 224004 188294 224604 225258
rect 224004 188058 224186 188294
rect 224422 188058 224604 188294
rect 224004 151094 224604 188058
rect 224004 150858 224186 151094
rect 224422 150858 224604 151094
rect 224004 113894 224604 150858
rect 224004 113658 224186 113894
rect 224422 113658 224604 113894
rect 224004 76694 224604 113658
rect 224004 76458 224186 76694
rect 224422 76458 224604 76694
rect 224004 39494 224604 76458
rect 224004 39258 224186 39494
rect 224422 39258 224604 39494
rect 224004 2294 224604 39258
rect 224004 2058 224186 2294
rect 224422 2058 224604 2294
rect 224004 -806 224604 2058
rect 224004 -1042 224186 -806
rect 224422 -1042 224604 -806
rect 224004 -2164 224604 -1042
rect 227604 705918 228204 706100
rect 227604 705682 227786 705918
rect 228022 705682 228204 705918
rect 227604 675494 228204 705682
rect 227604 675258 227786 675494
rect 228022 675258 228204 675494
rect 227604 638294 228204 675258
rect 227604 638058 227786 638294
rect 228022 638058 228204 638294
rect 227604 601094 228204 638058
rect 227604 600858 227786 601094
rect 228022 600858 228204 601094
rect 227604 563894 228204 600858
rect 227604 563658 227786 563894
rect 228022 563658 228204 563894
rect 227604 526694 228204 563658
rect 227604 526458 227786 526694
rect 228022 526458 228204 526694
rect 227604 489494 228204 526458
rect 227604 489258 227786 489494
rect 228022 489258 228204 489494
rect 227604 452294 228204 489258
rect 227604 452058 227786 452294
rect 228022 452058 228204 452294
rect 227604 415094 228204 452058
rect 227604 414858 227786 415094
rect 228022 414858 228204 415094
rect 227604 377894 228204 414858
rect 227604 377658 227786 377894
rect 228022 377658 228204 377894
rect 227604 340694 228204 377658
rect 227604 340458 227786 340694
rect 228022 340458 228204 340694
rect 227604 303494 228204 340458
rect 227604 303258 227786 303494
rect 228022 303258 228204 303494
rect 227604 266294 228204 303258
rect 227604 266058 227786 266294
rect 228022 266058 228204 266294
rect 227604 229094 228204 266058
rect 227604 228858 227786 229094
rect 228022 228858 228204 229094
rect 227604 191894 228204 228858
rect 227604 191658 227786 191894
rect 228022 191658 228204 191894
rect 227604 154694 228204 191658
rect 227604 154458 227786 154694
rect 228022 154458 228204 154694
rect 227604 117494 228204 154458
rect 227604 117258 227786 117494
rect 228022 117258 228204 117494
rect 227604 80294 228204 117258
rect 227604 80058 227786 80294
rect 228022 80058 228204 80294
rect 227604 43094 228204 80058
rect 227604 42858 227786 43094
rect 228022 42858 228204 43094
rect 227604 5894 228204 42858
rect 227604 5658 227786 5894
rect 228022 5658 228204 5894
rect 227604 -1746 228204 5658
rect 227604 -1982 227786 -1746
rect 228022 -1982 228204 -1746
rect 227604 -2164 228204 -1982
rect 261204 704978 261804 706100
rect 261204 704742 261386 704978
rect 261622 704742 261804 704978
rect 261204 671894 261804 704742
rect 261204 671658 261386 671894
rect 261622 671658 261804 671894
rect 261204 634694 261804 671658
rect 261204 634458 261386 634694
rect 261622 634458 261804 634694
rect 261204 597494 261804 634458
rect 261204 597258 261386 597494
rect 261622 597258 261804 597494
rect 261204 560294 261804 597258
rect 261204 560058 261386 560294
rect 261622 560058 261804 560294
rect 261204 523094 261804 560058
rect 261204 522858 261386 523094
rect 261622 522858 261804 523094
rect 261204 485894 261804 522858
rect 261204 485658 261386 485894
rect 261622 485658 261804 485894
rect 261204 448694 261804 485658
rect 261204 448458 261386 448694
rect 261622 448458 261804 448694
rect 261204 411494 261804 448458
rect 261204 411258 261386 411494
rect 261622 411258 261804 411494
rect 261204 374294 261804 411258
rect 261204 374058 261386 374294
rect 261622 374058 261804 374294
rect 261204 337094 261804 374058
rect 261204 336858 261386 337094
rect 261622 336858 261804 337094
rect 261204 299894 261804 336858
rect 261204 299658 261386 299894
rect 261622 299658 261804 299894
rect 261204 262694 261804 299658
rect 261204 262458 261386 262694
rect 261622 262458 261804 262694
rect 261204 225494 261804 262458
rect 261204 225258 261386 225494
rect 261622 225258 261804 225494
rect 261204 188294 261804 225258
rect 261204 188058 261386 188294
rect 261622 188058 261804 188294
rect 261204 151094 261804 188058
rect 261204 150858 261386 151094
rect 261622 150858 261804 151094
rect 261204 113894 261804 150858
rect 261204 113658 261386 113894
rect 261622 113658 261804 113894
rect 261204 76694 261804 113658
rect 261204 76458 261386 76694
rect 261622 76458 261804 76694
rect 261204 39494 261804 76458
rect 261204 39258 261386 39494
rect 261622 39258 261804 39494
rect 261204 2294 261804 39258
rect 261204 2058 261386 2294
rect 261622 2058 261804 2294
rect 261204 -806 261804 2058
rect 261204 -1042 261386 -806
rect 261622 -1042 261804 -806
rect 261204 -2164 261804 -1042
rect 264804 705918 265404 706100
rect 264804 705682 264986 705918
rect 265222 705682 265404 705918
rect 264804 675494 265404 705682
rect 264804 675258 264986 675494
rect 265222 675258 265404 675494
rect 264804 638294 265404 675258
rect 264804 638058 264986 638294
rect 265222 638058 265404 638294
rect 264804 601094 265404 638058
rect 264804 600858 264986 601094
rect 265222 600858 265404 601094
rect 264804 563894 265404 600858
rect 264804 563658 264986 563894
rect 265222 563658 265404 563894
rect 264804 526694 265404 563658
rect 264804 526458 264986 526694
rect 265222 526458 265404 526694
rect 264804 489494 265404 526458
rect 298404 704978 299004 706100
rect 298404 704742 298586 704978
rect 298822 704742 299004 704978
rect 298404 671894 299004 704742
rect 298404 671658 298586 671894
rect 298822 671658 299004 671894
rect 298404 634694 299004 671658
rect 298404 634458 298586 634694
rect 298822 634458 299004 634694
rect 298404 597494 299004 634458
rect 298404 597258 298586 597494
rect 298822 597258 299004 597494
rect 298404 560294 299004 597258
rect 298404 560058 298586 560294
rect 298822 560058 299004 560294
rect 298404 523094 299004 560058
rect 298404 522858 298586 523094
rect 298822 522858 299004 523094
rect 294827 490652 294893 490653
rect 294827 490588 294828 490652
rect 294892 490588 294893 490652
rect 294827 490587 294893 490588
rect 297955 490652 298021 490653
rect 297955 490588 297956 490652
rect 298020 490588 298021 490652
rect 297955 490587 298021 490588
rect 294830 489930 294890 490587
rect 264804 489258 264986 489494
rect 265222 489258 265404 489494
rect 264804 452294 265404 489258
rect 264804 452058 264986 452294
rect 265222 452058 265404 452294
rect 264804 415094 265404 452058
rect 294462 489870 294890 489930
rect 294462 450941 294522 489870
rect 296483 487252 296549 487253
rect 296483 487188 296484 487252
rect 296548 487188 296549 487252
rect 296483 487187 296549 487188
rect 294459 450940 294525 450941
rect 294459 450876 294460 450940
rect 294524 450876 294525 450940
rect 294459 450875 294525 450876
rect 294462 431085 294522 450875
rect 296299 447268 296365 447269
rect 296299 447204 296300 447268
rect 296364 447204 296365 447268
rect 296299 447203 296365 447204
rect 294459 431084 294525 431085
rect 294459 431020 294460 431084
rect 294524 431020 294525 431084
rect 294459 431019 294525 431020
rect 294462 422310 294522 431019
rect 294462 422250 295258 422310
rect 264804 414858 264986 415094
rect 265222 414858 265404 415094
rect 264804 377894 265404 414858
rect 295198 410141 295258 422250
rect 296302 418437 296362 447203
rect 296486 421157 296546 487187
rect 297958 453930 298018 490587
rect 298404 485894 299004 522858
rect 302004 705918 302604 706100
rect 302004 705682 302186 705918
rect 302422 705682 302604 705918
rect 302004 675494 302604 705682
rect 302004 675258 302186 675494
rect 302422 675258 302604 675494
rect 302004 638294 302604 675258
rect 302004 638058 302186 638294
rect 302422 638058 302604 638294
rect 302004 601094 302604 638058
rect 302004 600858 302186 601094
rect 302422 600858 302604 601094
rect 302004 563894 302604 600858
rect 302004 563658 302186 563894
rect 302422 563658 302604 563894
rect 302004 526694 302604 563658
rect 302004 526458 302186 526694
rect 302422 526458 302604 526694
rect 301083 490652 301149 490653
rect 301083 490588 301084 490652
rect 301148 490588 301149 490652
rect 301083 490587 301149 490588
rect 301086 489930 301146 490587
rect 301086 489870 301514 489930
rect 298404 485658 298586 485894
rect 298822 485658 299004 485894
rect 297958 453870 298202 453930
rect 298142 450533 298202 453870
rect 298139 450532 298205 450533
rect 298139 450468 298140 450532
rect 298204 450468 298205 450532
rect 298139 450467 298205 450468
rect 298142 431221 298202 450467
rect 298404 448694 299004 485658
rect 301267 451212 301333 451213
rect 301267 451148 301268 451212
rect 301332 451210 301333 451212
rect 301454 451210 301514 489870
rect 301332 451150 301514 451210
rect 301332 451148 301333 451150
rect 301267 451147 301333 451148
rect 298404 448458 298586 448694
rect 298822 448458 299004 448694
rect 298139 431220 298205 431221
rect 298139 431156 298140 431220
rect 298204 431156 298205 431220
rect 298139 431155 298205 431156
rect 296483 421156 296549 421157
rect 296483 421092 296484 421156
rect 296548 421092 296549 421156
rect 296483 421091 296549 421092
rect 296299 418436 296365 418437
rect 296299 418372 296300 418436
rect 296364 418372 296365 418436
rect 296299 418371 296365 418372
rect 298404 411494 299004 448458
rect 299243 431220 299309 431221
rect 299243 431156 299244 431220
rect 299308 431156 299309 431220
rect 299243 431155 299309 431156
rect 298404 411258 298586 411494
rect 298822 411258 299004 411494
rect 299246 411365 299306 431155
rect 301454 431085 301514 451150
rect 302004 489494 302604 526458
rect 335604 704978 336204 706100
rect 335604 704742 335786 704978
rect 336022 704742 336204 704978
rect 335604 671894 336204 704742
rect 335604 671658 335786 671894
rect 336022 671658 336204 671894
rect 335604 634694 336204 671658
rect 335604 634458 335786 634694
rect 336022 634458 336204 634694
rect 335604 597494 336204 634458
rect 335604 597258 335786 597494
rect 336022 597258 336204 597494
rect 335604 560294 336204 597258
rect 335604 560058 335786 560294
rect 336022 560058 336204 560294
rect 335604 523094 336204 560058
rect 335604 522858 335786 523094
rect 336022 522858 336204 523094
rect 304211 490652 304277 490653
rect 304211 490588 304212 490652
rect 304276 490588 304277 490652
rect 304211 490587 304277 490588
rect 302004 489258 302186 489494
rect 302422 489258 302604 489494
rect 302004 452294 302604 489258
rect 304214 460950 304274 490587
rect 307339 490380 307405 490381
rect 307339 490316 307340 490380
rect 307404 490316 307405 490380
rect 307339 490315 307405 490316
rect 307342 489930 307402 490315
rect 307342 489870 307586 489930
rect 306235 487252 306301 487253
rect 306235 487188 306236 487252
rect 306300 487188 306301 487252
rect 306235 487187 306301 487188
rect 304214 460890 304826 460950
rect 302004 452058 302186 452294
rect 302422 452058 302604 452294
rect 301451 431084 301517 431085
rect 301451 431020 301452 431084
rect 301516 431020 301517 431084
rect 301451 431019 301517 431020
rect 301454 422310 301514 431019
rect 301454 422250 301698 422310
rect 299243 411364 299309 411365
rect 299243 411300 299244 411364
rect 299308 411300 299309 411364
rect 299243 411299 299309 411300
rect 295195 410140 295261 410141
rect 295195 410076 295196 410140
rect 295260 410076 295261 410140
rect 295195 410075 295261 410076
rect 295198 391509 295258 410075
rect 295195 391508 295261 391509
rect 295195 391444 295196 391508
rect 295260 391444 295261 391508
rect 295195 391443 295261 391444
rect 264804 377658 264986 377894
rect 265222 377658 265404 377894
rect 264804 340694 265404 377658
rect 295198 374010 295258 391443
rect 298139 391236 298205 391237
rect 298139 391172 298140 391236
rect 298204 391172 298205 391236
rect 298139 391171 298205 391172
rect 294462 373950 295258 374010
rect 294462 370021 294522 373950
rect 298142 370021 298202 391171
rect 298404 374294 299004 411258
rect 299246 391509 299306 411299
rect 301638 410141 301698 422250
rect 302004 415094 302604 452058
rect 304579 451212 304645 451213
rect 304579 451148 304580 451212
rect 304644 451210 304645 451212
rect 304766 451210 304826 460890
rect 304644 451150 304826 451210
rect 304644 451148 304645 451150
rect 304579 451147 304645 451148
rect 304766 430677 304826 451150
rect 304763 430676 304829 430677
rect 304763 430612 304764 430676
rect 304828 430612 304829 430676
rect 304763 430611 304829 430612
rect 302004 414858 302186 415094
rect 302422 414858 302604 415094
rect 301635 410140 301701 410141
rect 301635 410076 301636 410140
rect 301700 410076 301701 410140
rect 301635 410075 301701 410076
rect 299243 391508 299309 391509
rect 299243 391444 299244 391508
rect 299308 391444 299309 391508
rect 299243 391443 299309 391444
rect 301638 391237 301698 410075
rect 301635 391236 301701 391237
rect 301635 391172 301636 391236
rect 301700 391172 301701 391236
rect 301635 391171 301701 391172
rect 301638 389190 301698 391171
rect 298404 374058 298586 374294
rect 298822 374058 299004 374294
rect 298404 372781 299004 374058
rect 301454 389130 301698 389190
rect 301454 374010 301514 389130
rect 300718 373950 301514 374010
rect 302004 377894 302604 414858
rect 304766 410141 304826 430611
rect 306051 426460 306117 426461
rect 306051 426396 306052 426460
rect 306116 426396 306117 426460
rect 306051 426395 306117 426396
rect 304763 410140 304829 410141
rect 304763 410076 304764 410140
rect 304828 410076 304829 410140
rect 304763 410075 304829 410076
rect 304766 391101 304826 410075
rect 304763 391100 304829 391101
rect 304763 391036 304764 391100
rect 304828 391036 304829 391100
rect 304763 391035 304829 391036
rect 304766 389190 304826 391035
rect 302004 377658 302186 377894
rect 302422 377658 302604 377894
rect 300718 370021 300778 373950
rect 302004 372781 302604 377658
rect 304582 389130 304826 389190
rect 304582 374010 304642 389130
rect 304763 386884 304829 386885
rect 304763 386820 304764 386884
rect 304828 386820 304829 386884
rect 304763 386819 304829 386820
rect 304214 373950 304642 374010
rect 304214 370021 304274 373950
rect 294459 370020 294525 370021
rect 294459 369956 294460 370020
rect 294524 369956 294525 370020
rect 294459 369955 294525 369956
rect 298139 370020 298205 370021
rect 298139 369956 298140 370020
rect 298204 369956 298205 370020
rect 298139 369955 298205 369956
rect 300715 370020 300781 370021
rect 300715 369956 300716 370020
rect 300780 369956 300781 370020
rect 300715 369955 300781 369956
rect 304211 370020 304277 370021
rect 304211 369956 304212 370020
rect 304276 369956 304277 370020
rect 304211 369955 304277 369956
rect 264804 340458 264986 340694
rect 265222 340458 265404 340694
rect 264804 303494 265404 340458
rect 264804 303258 264986 303494
rect 265222 303258 265404 303494
rect 264804 266294 265404 303258
rect 294462 291277 294522 369955
rect 298142 291277 298202 369955
rect 298404 337094 299004 368377
rect 298404 336858 298586 337094
rect 298822 336858 299004 337094
rect 298404 299894 299004 336858
rect 298404 299658 298586 299894
rect 298822 299658 299004 299894
rect 294459 291276 294525 291277
rect 294459 291212 294460 291276
rect 294524 291212 294525 291276
rect 294459 291211 294525 291212
rect 298139 291276 298205 291277
rect 298139 291212 298140 291276
rect 298204 291212 298205 291276
rect 298139 291211 298205 291212
rect 294462 287070 294522 291211
rect 294462 287010 294706 287070
rect 294646 271557 294706 287010
rect 294643 271556 294709 271557
rect 294643 271492 294644 271556
rect 294708 271492 294709 271556
rect 294643 271491 294709 271492
rect 294646 267750 294706 271491
rect 294646 267690 295258 267750
rect 264804 266058 264986 266294
rect 265222 266058 265404 266294
rect 264804 229094 265404 266058
rect 295198 252650 295258 267690
rect 298404 262694 299004 299658
rect 300718 296730 300778 369955
rect 300166 296670 300778 296730
rect 302004 340694 302604 368377
rect 302004 340458 302186 340694
rect 302422 340458 302604 340694
rect 302004 303494 302604 340458
rect 302004 303258 302186 303494
rect 302422 303258 302604 303494
rect 300166 291413 300226 296670
rect 300163 291412 300229 291413
rect 300163 291348 300164 291412
rect 300228 291348 300229 291412
rect 300163 291347 300229 291348
rect 299243 291276 299309 291277
rect 299243 291212 299244 291276
rect 299308 291212 299309 291276
rect 299243 291211 299309 291212
rect 299246 271557 299306 291211
rect 300166 287070 300226 291347
rect 300166 287010 300778 287070
rect 300718 273730 300778 287010
rect 300718 273670 300962 273730
rect 300902 271829 300962 273670
rect 300899 271828 300965 271829
rect 300899 271764 300900 271828
rect 300964 271764 300965 271828
rect 300899 271763 300965 271764
rect 299243 271556 299309 271557
rect 299243 271492 299244 271556
rect 299308 271492 299309 271556
rect 299243 271491 299309 271492
rect 301451 271556 301517 271557
rect 301451 271492 301452 271556
rect 301516 271492 301517 271556
rect 301451 271491 301517 271492
rect 298404 262458 298586 262694
rect 298822 262458 299004 262694
rect 295198 252590 295442 252650
rect 295382 251429 295442 252590
rect 295379 251428 295445 251429
rect 295379 251364 295380 251428
rect 295444 251364 295445 251428
rect 295379 251363 295445 251364
rect 295382 231437 295442 251363
rect 295379 231436 295445 231437
rect 295379 231372 295380 231436
rect 295444 231372 295445 231436
rect 295379 231371 295445 231372
rect 264804 228858 264986 229094
rect 265222 228858 265404 229094
rect 264804 191894 265404 228858
rect 295382 210493 295442 231371
rect 298139 230212 298205 230213
rect 298139 230148 298140 230212
rect 298204 230148 298205 230212
rect 298139 230147 298205 230148
rect 298142 210493 298202 230147
rect 298404 225494 299004 262458
rect 299246 251565 299306 271491
rect 301454 251565 301514 271491
rect 302004 266294 302604 303258
rect 304214 291549 304274 369955
rect 304766 334253 304826 386819
rect 304763 334252 304829 334253
rect 304763 334188 304764 334252
rect 304828 334188 304829 334252
rect 304763 334187 304829 334188
rect 306054 296989 306114 426395
rect 306238 301069 306298 487187
rect 307526 460950 307586 489870
rect 335604 485894 336204 522858
rect 335604 485658 335786 485894
rect 336022 485658 336204 485894
rect 307526 460890 307770 460950
rect 307710 450941 307770 460890
rect 307707 450940 307773 450941
rect 307707 450876 307708 450940
rect 307772 450876 307773 450940
rect 307707 450875 307773 450876
rect 307710 441630 307770 450875
rect 335604 448694 336204 485658
rect 335604 448458 335786 448694
rect 336022 448458 336204 448694
rect 307710 441570 308322 441630
rect 308262 430949 308322 441570
rect 308259 430948 308325 430949
rect 308259 430884 308260 430948
rect 308324 430884 308325 430948
rect 308259 430883 308325 430884
rect 308262 410141 308322 430883
rect 335604 411494 336204 448458
rect 335604 411258 335786 411494
rect 336022 411258 336204 411494
rect 308259 410140 308325 410141
rect 308259 410076 308260 410140
rect 308324 410076 308325 410140
rect 308259 410075 308325 410076
rect 308262 402990 308322 410075
rect 307894 402930 308322 402990
rect 307894 398850 307954 402930
rect 307710 398790 307954 398850
rect 307710 391101 307770 398790
rect 307707 391100 307773 391101
rect 307707 391036 307708 391100
rect 307772 391036 307773 391100
rect 307707 391035 307773 391036
rect 307710 389190 307770 391035
rect 307342 389130 307770 389190
rect 307342 374010 307402 389130
rect 307523 386884 307589 386885
rect 307523 386820 307524 386884
rect 307588 386820 307589 386884
rect 307523 386819 307589 386820
rect 306974 373950 307402 374010
rect 306974 370021 307034 373950
rect 306971 370020 307037 370021
rect 306971 369956 306972 370020
rect 307036 369956 307037 370020
rect 306971 369955 307037 369956
rect 306235 301068 306301 301069
rect 306235 301004 306236 301068
rect 306300 301004 306301 301068
rect 306235 301003 306301 301004
rect 306051 296988 306117 296989
rect 306051 296924 306052 296988
rect 306116 296924 306117 296988
rect 306051 296923 306117 296924
rect 306974 296730 307034 369955
rect 306790 296670 307034 296730
rect 304211 291548 304277 291549
rect 304211 291484 304212 291548
rect 304276 291484 304277 291548
rect 304211 291483 304277 291484
rect 304763 291548 304829 291549
rect 304763 291484 304764 291548
rect 304828 291484 304829 291548
rect 304763 291483 304829 291484
rect 304766 287070 304826 291483
rect 306790 291413 306850 296670
rect 307526 294269 307586 386819
rect 335604 374294 336204 411258
rect 335604 374058 335786 374294
rect 336022 374058 336204 374294
rect 335604 337094 336204 374058
rect 335604 336858 335786 337094
rect 336022 336858 336204 337094
rect 335604 299894 336204 336858
rect 335604 299658 335786 299894
rect 336022 299658 336204 299894
rect 307523 294268 307589 294269
rect 307523 294204 307524 294268
rect 307588 294204 307589 294268
rect 307523 294203 307589 294204
rect 306787 291412 306853 291413
rect 306787 291348 306788 291412
rect 306852 291348 306853 291412
rect 306787 291347 306853 291348
rect 306790 287070 306850 291347
rect 304766 287010 305010 287070
rect 306790 287010 307770 287070
rect 304950 271557 305010 287010
rect 307710 271693 307770 287010
rect 307707 271692 307773 271693
rect 307707 271628 307708 271692
rect 307772 271628 307773 271692
rect 307707 271627 307773 271628
rect 304947 271556 305013 271557
rect 304947 271492 304948 271556
rect 305012 271492 305013 271556
rect 304947 271491 305013 271492
rect 308259 271556 308325 271557
rect 308259 271492 308260 271556
rect 308324 271492 308325 271556
rect 308259 271491 308325 271492
rect 302004 266058 302186 266294
rect 302422 266058 302604 266294
rect 299243 251564 299309 251565
rect 299243 251500 299244 251564
rect 299308 251500 299309 251564
rect 299243 251499 299309 251500
rect 301451 251564 301517 251565
rect 301451 251500 301452 251564
rect 301516 251500 301517 251564
rect 301451 251499 301517 251500
rect 299246 231437 299306 251499
rect 299243 231436 299309 231437
rect 299243 231372 299244 231436
rect 299308 231372 299309 231436
rect 299243 231371 299309 231372
rect 298404 225258 298586 225494
rect 298822 225258 299004 225494
rect 298404 212781 299004 225258
rect 302004 229094 302604 266058
rect 302739 251564 302805 251565
rect 302739 251500 302740 251564
rect 302804 251500 302805 251564
rect 302739 251499 302805 251500
rect 302742 248430 302802 251499
rect 304950 251021 305010 271491
rect 308262 251565 308322 271491
rect 335604 262694 336204 299658
rect 335604 262458 335786 262694
rect 336022 262458 336204 262694
rect 308259 251564 308325 251565
rect 308259 251500 308260 251564
rect 308324 251500 308325 251564
rect 308259 251499 308325 251500
rect 304947 251020 305013 251021
rect 304947 250956 304948 251020
rect 305012 250956 305013 251020
rect 304947 250955 305013 250956
rect 304950 248430 305010 250955
rect 302742 248370 302986 248430
rect 304950 248370 306298 248430
rect 302926 230621 302986 248370
rect 306238 234630 306298 248370
rect 306238 234570 306482 234630
rect 306422 230621 306482 234570
rect 309731 233340 309797 233341
rect 309731 233276 309732 233340
rect 309796 233276 309797 233340
rect 309731 233275 309797 233276
rect 309734 230621 309794 233275
rect 302923 230620 302989 230621
rect 302923 230556 302924 230620
rect 302988 230556 302989 230620
rect 302923 230555 302989 230556
rect 306419 230620 306485 230621
rect 306419 230556 306420 230620
rect 306484 230556 306485 230620
rect 306419 230555 306485 230556
rect 309731 230620 309797 230621
rect 309731 230556 309732 230620
rect 309796 230556 309797 230620
rect 309731 230555 309797 230556
rect 302004 228858 302186 229094
rect 302422 228858 302604 229094
rect 302004 212781 302604 228858
rect 302739 211172 302805 211173
rect 302739 211108 302740 211172
rect 302804 211170 302805 211172
rect 302926 211170 302986 230555
rect 306422 213213 306482 230555
rect 309734 213349 309794 230555
rect 335604 225494 336204 262458
rect 335604 225258 335786 225494
rect 336022 225258 336204 225494
rect 309731 213348 309797 213349
rect 309731 213284 309732 213348
rect 309796 213284 309797 213348
rect 309731 213283 309797 213284
rect 306419 213212 306485 213213
rect 306419 213148 306420 213212
rect 306484 213148 306485 213212
rect 306419 213147 306485 213148
rect 302804 211110 302986 211170
rect 302804 211108 302805 211110
rect 302739 211107 302805 211108
rect 295379 210492 295445 210493
rect 295379 210428 295380 210492
rect 295444 210428 295445 210492
rect 295379 210427 295445 210428
rect 298139 210492 298205 210493
rect 298139 210428 298140 210492
rect 298204 210428 298205 210492
rect 298139 210427 298205 210428
rect 295382 209790 295442 210427
rect 295382 209730 295994 209790
rect 264804 191658 264986 191894
rect 265222 191658 265404 191894
rect 264804 154694 265404 191658
rect 264804 154458 264986 154694
rect 265222 154458 265404 154694
rect 264804 117494 265404 154458
rect 264804 117258 264986 117494
rect 265222 117258 265404 117494
rect 264804 80294 265404 117258
rect 264804 80058 264986 80294
rect 265222 80058 265404 80294
rect 264804 43094 265404 80058
rect 264804 42858 264986 43094
rect 265222 42858 265404 43094
rect 264804 5894 265404 42858
rect 295934 6629 295994 209730
rect 298142 46341 298202 210427
rect 298404 188294 299004 208377
rect 298404 188058 298586 188294
rect 298822 188058 299004 188294
rect 298404 151094 299004 188058
rect 298404 150858 298586 151094
rect 298822 150858 299004 151094
rect 298404 113894 299004 150858
rect 298404 113658 298586 113894
rect 298822 113658 299004 113894
rect 298404 76694 299004 113658
rect 298404 76458 298586 76694
rect 298822 76458 299004 76694
rect 298139 46340 298205 46341
rect 298139 46276 298140 46340
rect 298204 46276 298205 46340
rect 298139 46275 298205 46276
rect 298404 39494 299004 76458
rect 298404 39258 298586 39494
rect 298822 39258 299004 39494
rect 295931 6628 295997 6629
rect 295931 6564 295932 6628
rect 295996 6564 295997 6628
rect 295931 6563 295997 6564
rect 264804 5658 264986 5894
rect 265222 5658 265404 5894
rect 264804 -1746 265404 5658
rect 264804 -1982 264986 -1746
rect 265222 -1982 265404 -1746
rect 264804 -2164 265404 -1982
rect 298404 2294 299004 39258
rect 298404 2058 298586 2294
rect 298822 2058 299004 2294
rect 298404 -806 299004 2058
rect 298404 -1042 298586 -806
rect 298822 -1042 299004 -806
rect 298404 -2164 299004 -1042
rect 302004 191894 302604 208377
rect 302004 191658 302186 191894
rect 302422 191658 302604 191894
rect 302004 154694 302604 191658
rect 302004 154458 302186 154694
rect 302422 154458 302604 154694
rect 302004 117494 302604 154458
rect 302004 117258 302186 117494
rect 302422 117258 302604 117494
rect 302004 80294 302604 117258
rect 302926 86189 302986 211110
rect 335604 188294 336204 225258
rect 335604 188058 335786 188294
rect 336022 188058 336204 188294
rect 335604 151094 336204 188058
rect 335604 150858 335786 151094
rect 336022 150858 336204 151094
rect 335604 113894 336204 150858
rect 335604 113658 335786 113894
rect 336022 113658 336204 113894
rect 302923 86188 302989 86189
rect 302923 86124 302924 86188
rect 302988 86124 302989 86188
rect 302923 86123 302989 86124
rect 302004 80058 302186 80294
rect 302422 80058 302604 80294
rect 302004 43094 302604 80058
rect 302004 42858 302186 43094
rect 302422 42858 302604 43094
rect 302004 5894 302604 42858
rect 302004 5658 302186 5894
rect 302422 5658 302604 5894
rect 302004 -1746 302604 5658
rect 302004 -1982 302186 -1746
rect 302422 -1982 302604 -1746
rect 302004 -2164 302604 -1982
rect 335604 76694 336204 113658
rect 335604 76458 335786 76694
rect 336022 76458 336204 76694
rect 335604 39494 336204 76458
rect 335604 39258 335786 39494
rect 336022 39258 336204 39494
rect 335604 2294 336204 39258
rect 335604 2058 335786 2294
rect 336022 2058 336204 2294
rect 335604 -806 336204 2058
rect 335604 -1042 335786 -806
rect 336022 -1042 336204 -806
rect 335604 -2164 336204 -1042
rect 339204 705918 339804 706100
rect 339204 705682 339386 705918
rect 339622 705682 339804 705918
rect 339204 675494 339804 705682
rect 339204 675258 339386 675494
rect 339622 675258 339804 675494
rect 339204 638294 339804 675258
rect 339204 638058 339386 638294
rect 339622 638058 339804 638294
rect 339204 601094 339804 638058
rect 339204 600858 339386 601094
rect 339622 600858 339804 601094
rect 339204 563894 339804 600858
rect 339204 563658 339386 563894
rect 339622 563658 339804 563894
rect 339204 526694 339804 563658
rect 339204 526458 339386 526694
rect 339622 526458 339804 526694
rect 339204 489494 339804 526458
rect 339204 489258 339386 489494
rect 339622 489258 339804 489494
rect 339204 452294 339804 489258
rect 339204 452058 339386 452294
rect 339622 452058 339804 452294
rect 339204 415094 339804 452058
rect 339204 414858 339386 415094
rect 339622 414858 339804 415094
rect 339204 377894 339804 414858
rect 339204 377658 339386 377894
rect 339622 377658 339804 377894
rect 339204 340694 339804 377658
rect 339204 340458 339386 340694
rect 339622 340458 339804 340694
rect 339204 303494 339804 340458
rect 339204 303258 339386 303494
rect 339622 303258 339804 303494
rect 339204 266294 339804 303258
rect 339204 266058 339386 266294
rect 339622 266058 339804 266294
rect 339204 229094 339804 266058
rect 339204 228858 339386 229094
rect 339622 228858 339804 229094
rect 339204 191894 339804 228858
rect 339204 191658 339386 191894
rect 339622 191658 339804 191894
rect 339204 154694 339804 191658
rect 339204 154458 339386 154694
rect 339622 154458 339804 154694
rect 339204 117494 339804 154458
rect 339204 117258 339386 117494
rect 339622 117258 339804 117494
rect 339204 80294 339804 117258
rect 339204 80058 339386 80294
rect 339622 80058 339804 80294
rect 339204 43094 339804 80058
rect 339204 42858 339386 43094
rect 339622 42858 339804 43094
rect 339204 5894 339804 42858
rect 339204 5658 339386 5894
rect 339622 5658 339804 5894
rect 339204 -1746 339804 5658
rect 339204 -1982 339386 -1746
rect 339622 -1982 339804 -1746
rect 339204 -2164 339804 -1982
rect 372804 704978 373404 706100
rect 372804 704742 372986 704978
rect 373222 704742 373404 704978
rect 372804 671894 373404 704742
rect 372804 671658 372986 671894
rect 373222 671658 373404 671894
rect 372804 634694 373404 671658
rect 372804 634458 372986 634694
rect 373222 634458 373404 634694
rect 372804 597494 373404 634458
rect 372804 597258 372986 597494
rect 373222 597258 373404 597494
rect 372804 560294 373404 597258
rect 372804 560058 372986 560294
rect 373222 560058 373404 560294
rect 372804 523094 373404 560058
rect 372804 522858 372986 523094
rect 373222 522858 373404 523094
rect 372804 485894 373404 522858
rect 372804 485658 372986 485894
rect 373222 485658 373404 485894
rect 372804 448694 373404 485658
rect 372804 448458 372986 448694
rect 373222 448458 373404 448694
rect 372804 411494 373404 448458
rect 372804 411258 372986 411494
rect 373222 411258 373404 411494
rect 372804 374294 373404 411258
rect 372804 374058 372986 374294
rect 373222 374058 373404 374294
rect 372804 337094 373404 374058
rect 372804 336858 372986 337094
rect 373222 336858 373404 337094
rect 372804 299894 373404 336858
rect 372804 299658 372986 299894
rect 373222 299658 373404 299894
rect 372804 262694 373404 299658
rect 372804 262458 372986 262694
rect 373222 262458 373404 262694
rect 372804 225494 373404 262458
rect 372804 225258 372986 225494
rect 373222 225258 373404 225494
rect 372804 188294 373404 225258
rect 372804 188058 372986 188294
rect 373222 188058 373404 188294
rect 372804 151094 373404 188058
rect 372804 150858 372986 151094
rect 373222 150858 373404 151094
rect 372804 113894 373404 150858
rect 372804 113658 372986 113894
rect 373222 113658 373404 113894
rect 372804 76694 373404 113658
rect 372804 76458 372986 76694
rect 373222 76458 373404 76694
rect 372804 39494 373404 76458
rect 372804 39258 372986 39494
rect 373222 39258 373404 39494
rect 372804 2294 373404 39258
rect 372804 2058 372986 2294
rect 373222 2058 373404 2294
rect 372804 -806 373404 2058
rect 372804 -1042 372986 -806
rect 373222 -1042 373404 -806
rect 372804 -2164 373404 -1042
rect 376404 705918 377004 706100
rect 376404 705682 376586 705918
rect 376822 705682 377004 705918
rect 376404 675494 377004 705682
rect 376404 675258 376586 675494
rect 376822 675258 377004 675494
rect 376404 638294 377004 675258
rect 376404 638058 376586 638294
rect 376822 638058 377004 638294
rect 376404 601094 377004 638058
rect 376404 600858 376586 601094
rect 376822 600858 377004 601094
rect 376404 563894 377004 600858
rect 376404 563658 376586 563894
rect 376822 563658 377004 563894
rect 376404 526694 377004 563658
rect 376404 526458 376586 526694
rect 376822 526458 377004 526694
rect 376404 489494 377004 526458
rect 376404 489258 376586 489494
rect 376822 489258 377004 489494
rect 376404 452294 377004 489258
rect 376404 452058 376586 452294
rect 376822 452058 377004 452294
rect 376404 415094 377004 452058
rect 376404 414858 376586 415094
rect 376822 414858 377004 415094
rect 376404 377894 377004 414858
rect 376404 377658 376586 377894
rect 376822 377658 377004 377894
rect 376404 340694 377004 377658
rect 376404 340458 376586 340694
rect 376822 340458 377004 340694
rect 376404 303494 377004 340458
rect 376404 303258 376586 303494
rect 376822 303258 377004 303494
rect 376404 266294 377004 303258
rect 376404 266058 376586 266294
rect 376822 266058 377004 266294
rect 376404 229094 377004 266058
rect 376404 228858 376586 229094
rect 376822 228858 377004 229094
rect 376404 191894 377004 228858
rect 376404 191658 376586 191894
rect 376822 191658 377004 191894
rect 376404 154694 377004 191658
rect 376404 154458 376586 154694
rect 376822 154458 377004 154694
rect 376404 117494 377004 154458
rect 376404 117258 376586 117494
rect 376822 117258 377004 117494
rect 376404 80294 377004 117258
rect 376404 80058 376586 80294
rect 376822 80058 377004 80294
rect 376404 43094 377004 80058
rect 376404 42858 376586 43094
rect 376822 42858 377004 43094
rect 376404 5894 377004 42858
rect 376404 5658 376586 5894
rect 376822 5658 377004 5894
rect 376404 -1746 377004 5658
rect 376404 -1982 376586 -1746
rect 376822 -1982 377004 -1746
rect 376404 -2164 377004 -1982
rect 410004 704978 410604 706100
rect 410004 704742 410186 704978
rect 410422 704742 410604 704978
rect 410004 671894 410604 704742
rect 410004 671658 410186 671894
rect 410422 671658 410604 671894
rect 410004 634694 410604 671658
rect 410004 634458 410186 634694
rect 410422 634458 410604 634694
rect 410004 597494 410604 634458
rect 410004 597258 410186 597494
rect 410422 597258 410604 597494
rect 410004 560294 410604 597258
rect 410004 560058 410186 560294
rect 410422 560058 410604 560294
rect 410004 523094 410604 560058
rect 410004 522858 410186 523094
rect 410422 522858 410604 523094
rect 410004 485894 410604 522858
rect 410004 485658 410186 485894
rect 410422 485658 410604 485894
rect 410004 448694 410604 485658
rect 410004 448458 410186 448694
rect 410422 448458 410604 448694
rect 410004 411494 410604 448458
rect 410004 411258 410186 411494
rect 410422 411258 410604 411494
rect 410004 374294 410604 411258
rect 410004 374058 410186 374294
rect 410422 374058 410604 374294
rect 410004 337094 410604 374058
rect 410004 336858 410186 337094
rect 410422 336858 410604 337094
rect 410004 299894 410604 336858
rect 410004 299658 410186 299894
rect 410422 299658 410604 299894
rect 410004 262694 410604 299658
rect 410004 262458 410186 262694
rect 410422 262458 410604 262694
rect 410004 225494 410604 262458
rect 410004 225258 410186 225494
rect 410422 225258 410604 225494
rect 410004 188294 410604 225258
rect 410004 188058 410186 188294
rect 410422 188058 410604 188294
rect 410004 151094 410604 188058
rect 410004 150858 410186 151094
rect 410422 150858 410604 151094
rect 410004 113894 410604 150858
rect 410004 113658 410186 113894
rect 410422 113658 410604 113894
rect 410004 76694 410604 113658
rect 410004 76458 410186 76694
rect 410422 76458 410604 76694
rect 410004 39494 410604 76458
rect 410004 39258 410186 39494
rect 410422 39258 410604 39494
rect 410004 2294 410604 39258
rect 410004 2058 410186 2294
rect 410422 2058 410604 2294
rect 410004 -806 410604 2058
rect 410004 -1042 410186 -806
rect 410422 -1042 410604 -806
rect 410004 -2164 410604 -1042
rect 413604 705918 414204 706100
rect 413604 705682 413786 705918
rect 414022 705682 414204 705918
rect 413604 675494 414204 705682
rect 413604 675258 413786 675494
rect 414022 675258 414204 675494
rect 413604 638294 414204 675258
rect 413604 638058 413786 638294
rect 414022 638058 414204 638294
rect 413604 601094 414204 638058
rect 413604 600858 413786 601094
rect 414022 600858 414204 601094
rect 413604 563894 414204 600858
rect 413604 563658 413786 563894
rect 414022 563658 414204 563894
rect 413604 526694 414204 563658
rect 413604 526458 413786 526694
rect 414022 526458 414204 526694
rect 413604 489494 414204 526458
rect 413604 489258 413786 489494
rect 414022 489258 414204 489494
rect 413604 452294 414204 489258
rect 413604 452058 413786 452294
rect 414022 452058 414204 452294
rect 413604 415094 414204 452058
rect 413604 414858 413786 415094
rect 414022 414858 414204 415094
rect 413604 377894 414204 414858
rect 413604 377658 413786 377894
rect 414022 377658 414204 377894
rect 413604 340694 414204 377658
rect 413604 340458 413786 340694
rect 414022 340458 414204 340694
rect 413604 303494 414204 340458
rect 413604 303258 413786 303494
rect 414022 303258 414204 303494
rect 413604 266294 414204 303258
rect 413604 266058 413786 266294
rect 414022 266058 414204 266294
rect 413604 229094 414204 266058
rect 413604 228858 413786 229094
rect 414022 228858 414204 229094
rect 413604 191894 414204 228858
rect 413604 191658 413786 191894
rect 414022 191658 414204 191894
rect 413604 154694 414204 191658
rect 413604 154458 413786 154694
rect 414022 154458 414204 154694
rect 413604 117494 414204 154458
rect 413604 117258 413786 117494
rect 414022 117258 414204 117494
rect 413604 80294 414204 117258
rect 413604 80058 413786 80294
rect 414022 80058 414204 80294
rect 413604 43094 414204 80058
rect 413604 42858 413786 43094
rect 414022 42858 414204 43094
rect 413604 5894 414204 42858
rect 413604 5658 413786 5894
rect 414022 5658 414204 5894
rect 413604 -1746 414204 5658
rect 413604 -1982 413786 -1746
rect 414022 -1982 414204 -1746
rect 413604 -2164 414204 -1982
rect 447204 704978 447804 706100
rect 447204 704742 447386 704978
rect 447622 704742 447804 704978
rect 447204 671894 447804 704742
rect 447204 671658 447386 671894
rect 447622 671658 447804 671894
rect 447204 634694 447804 671658
rect 447204 634458 447386 634694
rect 447622 634458 447804 634694
rect 447204 597494 447804 634458
rect 447204 597258 447386 597494
rect 447622 597258 447804 597494
rect 447204 560294 447804 597258
rect 447204 560058 447386 560294
rect 447622 560058 447804 560294
rect 447204 523094 447804 560058
rect 447204 522858 447386 523094
rect 447622 522858 447804 523094
rect 447204 485894 447804 522858
rect 447204 485658 447386 485894
rect 447622 485658 447804 485894
rect 447204 448694 447804 485658
rect 447204 448458 447386 448694
rect 447622 448458 447804 448694
rect 447204 411494 447804 448458
rect 447204 411258 447386 411494
rect 447622 411258 447804 411494
rect 447204 374294 447804 411258
rect 447204 374058 447386 374294
rect 447622 374058 447804 374294
rect 447204 337094 447804 374058
rect 447204 336858 447386 337094
rect 447622 336858 447804 337094
rect 447204 299894 447804 336858
rect 447204 299658 447386 299894
rect 447622 299658 447804 299894
rect 447204 262694 447804 299658
rect 447204 262458 447386 262694
rect 447622 262458 447804 262694
rect 447204 225494 447804 262458
rect 447204 225258 447386 225494
rect 447622 225258 447804 225494
rect 447204 188294 447804 225258
rect 447204 188058 447386 188294
rect 447622 188058 447804 188294
rect 447204 151094 447804 188058
rect 447204 150858 447386 151094
rect 447622 150858 447804 151094
rect 447204 113894 447804 150858
rect 447204 113658 447386 113894
rect 447622 113658 447804 113894
rect 447204 76694 447804 113658
rect 447204 76458 447386 76694
rect 447622 76458 447804 76694
rect 447204 39494 447804 76458
rect 447204 39258 447386 39494
rect 447622 39258 447804 39494
rect 447204 2294 447804 39258
rect 447204 2058 447386 2294
rect 447622 2058 447804 2294
rect 447204 -806 447804 2058
rect 447204 -1042 447386 -806
rect 447622 -1042 447804 -806
rect 447204 -2164 447804 -1042
rect 450804 705918 451404 706100
rect 450804 705682 450986 705918
rect 451222 705682 451404 705918
rect 450804 675494 451404 705682
rect 450804 675258 450986 675494
rect 451222 675258 451404 675494
rect 450804 638294 451404 675258
rect 450804 638058 450986 638294
rect 451222 638058 451404 638294
rect 450804 601094 451404 638058
rect 450804 600858 450986 601094
rect 451222 600858 451404 601094
rect 450804 563894 451404 600858
rect 450804 563658 450986 563894
rect 451222 563658 451404 563894
rect 450804 526694 451404 563658
rect 450804 526458 450986 526694
rect 451222 526458 451404 526694
rect 450804 489494 451404 526458
rect 450804 489258 450986 489494
rect 451222 489258 451404 489494
rect 450804 452294 451404 489258
rect 450804 452058 450986 452294
rect 451222 452058 451404 452294
rect 450804 415094 451404 452058
rect 450804 414858 450986 415094
rect 451222 414858 451404 415094
rect 450804 377894 451404 414858
rect 450804 377658 450986 377894
rect 451222 377658 451404 377894
rect 450804 340694 451404 377658
rect 450804 340458 450986 340694
rect 451222 340458 451404 340694
rect 450804 303494 451404 340458
rect 450804 303258 450986 303494
rect 451222 303258 451404 303494
rect 450804 266294 451404 303258
rect 450804 266058 450986 266294
rect 451222 266058 451404 266294
rect 450804 229094 451404 266058
rect 450804 228858 450986 229094
rect 451222 228858 451404 229094
rect 450804 191894 451404 228858
rect 450804 191658 450986 191894
rect 451222 191658 451404 191894
rect 450804 154694 451404 191658
rect 450804 154458 450986 154694
rect 451222 154458 451404 154694
rect 450804 117494 451404 154458
rect 450804 117258 450986 117494
rect 451222 117258 451404 117494
rect 450804 80294 451404 117258
rect 450804 80058 450986 80294
rect 451222 80058 451404 80294
rect 450804 43094 451404 80058
rect 450804 42858 450986 43094
rect 451222 42858 451404 43094
rect 450804 5894 451404 42858
rect 450804 5658 450986 5894
rect 451222 5658 451404 5894
rect 450804 -1746 451404 5658
rect 450804 -1982 450986 -1746
rect 451222 -1982 451404 -1746
rect 450804 -2164 451404 -1982
rect 484404 704978 485004 706100
rect 484404 704742 484586 704978
rect 484822 704742 485004 704978
rect 484404 671894 485004 704742
rect 484404 671658 484586 671894
rect 484822 671658 485004 671894
rect 484404 634694 485004 671658
rect 484404 634458 484586 634694
rect 484822 634458 485004 634694
rect 484404 597494 485004 634458
rect 484404 597258 484586 597494
rect 484822 597258 485004 597494
rect 484404 560294 485004 597258
rect 484404 560058 484586 560294
rect 484822 560058 485004 560294
rect 484404 523094 485004 560058
rect 484404 522858 484586 523094
rect 484822 522858 485004 523094
rect 484404 485894 485004 522858
rect 484404 485658 484586 485894
rect 484822 485658 485004 485894
rect 484404 448694 485004 485658
rect 484404 448458 484586 448694
rect 484822 448458 485004 448694
rect 484404 411494 485004 448458
rect 484404 411258 484586 411494
rect 484822 411258 485004 411494
rect 484404 374294 485004 411258
rect 484404 374058 484586 374294
rect 484822 374058 485004 374294
rect 484404 337094 485004 374058
rect 484404 336858 484586 337094
rect 484822 336858 485004 337094
rect 484404 299894 485004 336858
rect 484404 299658 484586 299894
rect 484822 299658 485004 299894
rect 484404 262694 485004 299658
rect 484404 262458 484586 262694
rect 484822 262458 485004 262694
rect 484404 225494 485004 262458
rect 484404 225258 484586 225494
rect 484822 225258 485004 225494
rect 484404 188294 485004 225258
rect 484404 188058 484586 188294
rect 484822 188058 485004 188294
rect 484404 151094 485004 188058
rect 484404 150858 484586 151094
rect 484822 150858 485004 151094
rect 484404 113894 485004 150858
rect 484404 113658 484586 113894
rect 484822 113658 485004 113894
rect 484404 76694 485004 113658
rect 484404 76458 484586 76694
rect 484822 76458 485004 76694
rect 484404 39494 485004 76458
rect 484404 39258 484586 39494
rect 484822 39258 485004 39494
rect 484404 2294 485004 39258
rect 484404 2058 484586 2294
rect 484822 2058 485004 2294
rect 484404 -806 485004 2058
rect 484404 -1042 484586 -806
rect 484822 -1042 485004 -806
rect 484404 -2164 485004 -1042
rect 488004 705918 488604 706100
rect 488004 705682 488186 705918
rect 488422 705682 488604 705918
rect 488004 675494 488604 705682
rect 488004 675258 488186 675494
rect 488422 675258 488604 675494
rect 488004 638294 488604 675258
rect 488004 638058 488186 638294
rect 488422 638058 488604 638294
rect 488004 601094 488604 638058
rect 488004 600858 488186 601094
rect 488422 600858 488604 601094
rect 488004 563894 488604 600858
rect 488004 563658 488186 563894
rect 488422 563658 488604 563894
rect 488004 526694 488604 563658
rect 488004 526458 488186 526694
rect 488422 526458 488604 526694
rect 488004 489494 488604 526458
rect 488004 489258 488186 489494
rect 488422 489258 488604 489494
rect 488004 452294 488604 489258
rect 488004 452058 488186 452294
rect 488422 452058 488604 452294
rect 488004 415094 488604 452058
rect 521604 704978 522204 706100
rect 521604 704742 521786 704978
rect 522022 704742 522204 704978
rect 521604 671894 522204 704742
rect 521604 671658 521786 671894
rect 522022 671658 522204 671894
rect 521604 634694 522204 671658
rect 521604 634458 521786 634694
rect 522022 634458 522204 634694
rect 521604 597494 522204 634458
rect 521604 597258 521786 597494
rect 522022 597258 522204 597494
rect 521604 560294 522204 597258
rect 521604 560058 521786 560294
rect 522022 560058 522204 560294
rect 521604 523094 522204 560058
rect 521604 522858 521786 523094
rect 522022 522858 522204 523094
rect 521604 485894 522204 522858
rect 521604 485658 521786 485894
rect 522022 485658 522204 485894
rect 521604 448694 522204 485658
rect 521604 448458 521786 448694
rect 522022 448458 522204 448694
rect 521604 421752 522204 448458
rect 525204 705918 525804 706100
rect 525204 705682 525386 705918
rect 525622 705682 525804 705918
rect 525204 675494 525804 705682
rect 525204 675258 525386 675494
rect 525622 675258 525804 675494
rect 525204 638294 525804 675258
rect 525204 638058 525386 638294
rect 525622 638058 525804 638294
rect 525204 601094 525804 638058
rect 525204 600858 525386 601094
rect 525622 600858 525804 601094
rect 525204 563894 525804 600858
rect 525204 563658 525386 563894
rect 525622 563658 525804 563894
rect 525204 526694 525804 563658
rect 525204 526458 525386 526694
rect 525622 526458 525804 526694
rect 525204 489494 525804 526458
rect 525204 489258 525386 489494
rect 525622 489258 525804 489494
rect 525204 452294 525804 489258
rect 525204 452058 525386 452294
rect 525622 452058 525804 452294
rect 525204 421752 525804 452058
rect 558804 704978 559404 706100
rect 558804 704742 558986 704978
rect 559222 704742 559404 704978
rect 558804 671894 559404 704742
rect 558804 671658 558986 671894
rect 559222 671658 559404 671894
rect 558804 634694 559404 671658
rect 558804 634458 558986 634694
rect 559222 634458 559404 634694
rect 558804 597494 559404 634458
rect 558804 597258 558986 597494
rect 559222 597258 559404 597494
rect 558804 560294 559404 597258
rect 558804 560058 558986 560294
rect 559222 560058 559404 560294
rect 558804 523094 559404 560058
rect 558804 522858 558986 523094
rect 559222 522858 559404 523094
rect 558804 485894 559404 522858
rect 558804 485658 558986 485894
rect 559222 485658 559404 485894
rect 558804 448694 559404 485658
rect 558804 448458 558986 448694
rect 559222 448458 559404 448694
rect 523539 421292 523605 421293
rect 523539 421228 523540 421292
rect 523604 421228 523605 421292
rect 523539 421227 523605 421228
rect 526299 421292 526365 421293
rect 526299 421228 526300 421292
rect 526364 421228 526365 421292
rect 526299 421227 526365 421228
rect 488004 414858 488186 415094
rect 488422 414858 488604 415094
rect 488004 377894 488604 414858
rect 523542 383757 523602 421227
rect 526302 383757 526362 421227
rect 558804 411494 559404 448458
rect 558804 411258 558986 411494
rect 559222 411258 559404 411494
rect 531451 410956 531517 410957
rect 531451 410892 531452 410956
rect 531516 410892 531517 410956
rect 531451 410891 531517 410892
rect 523539 383756 523605 383757
rect 523539 383692 523540 383756
rect 523604 383692 523605 383756
rect 523539 383691 523605 383692
rect 526299 383756 526365 383757
rect 526299 383692 526300 383756
rect 526364 383692 526365 383756
rect 526299 383691 526365 383692
rect 488004 377658 488186 377894
rect 488422 377658 488604 377894
rect 488004 340694 488604 377658
rect 523542 341325 523602 383691
rect 526302 374010 526362 383691
rect 526302 373950 526546 374010
rect 526486 354690 526546 373950
rect 531454 370973 531514 410891
rect 558804 374294 559404 411258
rect 558804 374058 558986 374294
rect 559222 374058 559404 374294
rect 531451 370972 531517 370973
rect 531451 370908 531452 370972
rect 531516 370908 531517 370972
rect 531451 370907 531517 370908
rect 526486 354630 527098 354690
rect 527038 351933 527098 354630
rect 527035 351932 527101 351933
rect 527035 351868 527036 351932
rect 527100 351868 527101 351932
rect 527035 351867 527101 351868
rect 527038 345030 527098 351867
rect 526302 344970 527098 345030
rect 526302 341325 526362 344970
rect 523539 341324 523605 341325
rect 523539 341260 523540 341324
rect 523604 341260 523605 341324
rect 523539 341259 523605 341260
rect 526299 341324 526365 341325
rect 526299 341260 526300 341324
rect 526364 341260 526365 341324
rect 526299 341259 526365 341260
rect 488004 340458 488186 340694
rect 488422 340458 488604 340694
rect 488004 303494 488604 340458
rect 488004 303258 488186 303494
rect 488422 303258 488604 303494
rect 488004 266294 488604 303258
rect 523542 302293 523602 341259
rect 526302 303653 526362 341259
rect 531454 330989 531514 370907
rect 558804 337094 559404 374058
rect 558804 336858 558986 337094
rect 559222 336858 559404 337094
rect 531451 330988 531517 330989
rect 531451 330924 531452 330988
rect 531516 330924 531517 330988
rect 531451 330923 531517 330924
rect 526299 303652 526365 303653
rect 526299 303588 526300 303652
rect 526364 303588 526365 303652
rect 526299 303587 526365 303588
rect 523539 302292 523605 302293
rect 523539 302228 523540 302292
rect 523604 302228 523605 302292
rect 523539 302227 523605 302228
rect 524275 302292 524341 302293
rect 524275 302228 524276 302292
rect 524340 302228 524341 302292
rect 524275 302227 524341 302228
rect 488004 266058 488186 266294
rect 488422 266058 488604 266294
rect 488004 229094 488604 266058
rect 524278 264621 524338 302227
rect 526302 264621 526362 303587
rect 531454 291005 531514 330923
rect 558804 299894 559404 336858
rect 558804 299658 558986 299894
rect 559222 299658 559404 299894
rect 531451 291004 531517 291005
rect 531451 290940 531452 291004
rect 531516 290940 531517 291004
rect 531451 290939 531517 290940
rect 524275 264620 524341 264621
rect 524275 264556 524276 264620
rect 524340 264556 524341 264620
rect 524275 264555 524341 264556
rect 526299 264620 526365 264621
rect 526299 264556 526300 264620
rect 526364 264556 526365 264620
rect 526299 264555 526365 264556
rect 531454 251021 531514 290939
rect 558804 262694 559404 299658
rect 558804 262458 558986 262694
rect 559222 262458 559404 262694
rect 531451 251020 531517 251021
rect 531451 250956 531452 251020
rect 531516 250956 531517 251020
rect 531451 250955 531517 250956
rect 531454 248430 531514 250955
rect 531454 248370 531882 248430
rect 488004 228858 488186 229094
rect 488422 228858 488604 229094
rect 488004 191894 488604 228858
rect 488004 191658 488186 191894
rect 488422 191658 488604 191894
rect 488004 154694 488604 191658
rect 488004 154458 488186 154694
rect 488422 154458 488604 154694
rect 488004 117494 488604 154458
rect 488004 117258 488186 117494
rect 488422 117258 488604 117494
rect 488004 80294 488604 117258
rect 488004 80058 488186 80294
rect 488422 80058 488604 80294
rect 488004 43094 488604 80058
rect 488004 42858 488186 43094
rect 488422 42858 488604 43094
rect 488004 5894 488604 42858
rect 488004 5658 488186 5894
rect 488422 5658 488604 5894
rect 488004 -1746 488604 5658
rect 488004 -1982 488186 -1746
rect 488422 -1982 488604 -1746
rect 488004 -2164 488604 -1982
rect 521604 225494 522204 240008
rect 521604 225258 521786 225494
rect 522022 225258 522204 225494
rect 521604 188294 522204 225258
rect 521604 188058 521786 188294
rect 522022 188058 522204 188294
rect 521604 151094 522204 188058
rect 521604 150858 521786 151094
rect 522022 150858 522204 151094
rect 521604 113894 522204 150858
rect 521604 113658 521786 113894
rect 522022 113658 522204 113894
rect 521604 76694 522204 113658
rect 521604 76458 521786 76694
rect 522022 76458 522204 76694
rect 521604 39494 522204 76458
rect 521604 39258 521786 39494
rect 522022 39258 522204 39494
rect 521604 2294 522204 39258
rect 521604 2058 521786 2294
rect 522022 2058 522204 2294
rect 521604 -806 522204 2058
rect 521604 -1042 521786 -806
rect 522022 -1042 522204 -806
rect 521604 -2164 522204 -1042
rect 525204 229094 525804 240008
rect 525204 228858 525386 229094
rect 525622 228858 525804 229094
rect 525204 191894 525804 228858
rect 525204 191658 525386 191894
rect 525622 191658 525804 191894
rect 525204 154694 525804 191658
rect 525204 154458 525386 154694
rect 525622 154458 525804 154694
rect 525204 117494 525804 154458
rect 525204 117258 525386 117494
rect 525622 117258 525804 117494
rect 525204 80294 525804 117258
rect 525204 80058 525386 80294
rect 525622 80058 525804 80294
rect 525204 43094 525804 80058
rect 525204 42858 525386 43094
rect 525622 42858 525804 43094
rect 525204 5894 525804 42858
rect 531822 19821 531882 248370
rect 558804 225494 559404 262458
rect 558804 225258 558986 225494
rect 559222 225258 559404 225494
rect 558804 188294 559404 225258
rect 558804 188058 558986 188294
rect 559222 188058 559404 188294
rect 558804 151094 559404 188058
rect 558804 150858 558986 151094
rect 559222 150858 559404 151094
rect 558804 113894 559404 150858
rect 558804 113658 558986 113894
rect 559222 113658 559404 113894
rect 558804 76694 559404 113658
rect 558804 76458 558986 76694
rect 559222 76458 559404 76694
rect 558804 39494 559404 76458
rect 558804 39258 558986 39494
rect 559222 39258 559404 39494
rect 531819 19820 531885 19821
rect 531819 19756 531820 19820
rect 531884 19756 531885 19820
rect 531819 19755 531885 19756
rect 525204 5658 525386 5894
rect 525622 5658 525804 5894
rect 525204 -1746 525804 5658
rect 525204 -1982 525386 -1746
rect 525622 -1982 525804 -1746
rect 525204 -2164 525804 -1982
rect 558804 2294 559404 39258
rect 558804 2058 558986 2294
rect 559222 2058 559404 2294
rect 558804 -806 559404 2058
rect 558804 -1042 558986 -806
rect 559222 -1042 559404 -806
rect 558804 -2164 559404 -1042
rect 562404 705918 563004 706100
rect 562404 705682 562586 705918
rect 562822 705682 563004 705918
rect 562404 675494 563004 705682
rect 586560 705918 587160 706100
rect 586560 705682 586742 705918
rect 586978 705682 587160 705918
rect 562404 675258 562586 675494
rect 562822 675258 563004 675494
rect 562404 638294 563004 675258
rect 562404 638058 562586 638294
rect 562822 638058 563004 638294
rect 562404 601094 563004 638058
rect 562404 600858 562586 601094
rect 562822 600858 563004 601094
rect 562404 563894 563004 600858
rect 562404 563658 562586 563894
rect 562822 563658 563004 563894
rect 562404 526694 563004 563658
rect 562404 526458 562586 526694
rect 562822 526458 563004 526694
rect 562404 489494 563004 526458
rect 562404 489258 562586 489494
rect 562822 489258 563004 489494
rect 562404 452294 563004 489258
rect 562404 452058 562586 452294
rect 562822 452058 563004 452294
rect 562404 415094 563004 452058
rect 562404 414858 562586 415094
rect 562822 414858 563004 415094
rect 562404 377894 563004 414858
rect 562404 377658 562586 377894
rect 562822 377658 563004 377894
rect 562404 340694 563004 377658
rect 562404 340458 562586 340694
rect 562822 340458 563004 340694
rect 562404 303494 563004 340458
rect 562404 303258 562586 303494
rect 562822 303258 563004 303494
rect 562404 266294 563004 303258
rect 562404 266058 562586 266294
rect 562822 266058 563004 266294
rect 562404 229094 563004 266058
rect 562404 228858 562586 229094
rect 562822 228858 563004 229094
rect 562404 191894 563004 228858
rect 562404 191658 562586 191894
rect 562822 191658 563004 191894
rect 562404 154694 563004 191658
rect 562404 154458 562586 154694
rect 562822 154458 563004 154694
rect 562404 117494 563004 154458
rect 562404 117258 562586 117494
rect 562822 117258 563004 117494
rect 562404 80294 563004 117258
rect 562404 80058 562586 80294
rect 562822 80058 563004 80294
rect 562404 43094 563004 80058
rect 562404 42858 562586 43094
rect 562822 42858 563004 43094
rect 562404 5894 563004 42858
rect 562404 5658 562586 5894
rect 562822 5658 563004 5894
rect 562404 -1746 563004 5658
rect 585620 704978 586220 705160
rect 585620 704742 585802 704978
rect 586038 704742 586220 704978
rect 585620 671894 586220 704742
rect 585620 671658 585802 671894
rect 586038 671658 586220 671894
rect 585620 634694 586220 671658
rect 585620 634458 585802 634694
rect 586038 634458 586220 634694
rect 585620 597494 586220 634458
rect 585620 597258 585802 597494
rect 586038 597258 586220 597494
rect 585620 560294 586220 597258
rect 585620 560058 585802 560294
rect 586038 560058 586220 560294
rect 585620 523094 586220 560058
rect 585620 522858 585802 523094
rect 586038 522858 586220 523094
rect 585620 485894 586220 522858
rect 585620 485658 585802 485894
rect 586038 485658 586220 485894
rect 585620 448694 586220 485658
rect 585620 448458 585802 448694
rect 586038 448458 586220 448694
rect 585620 411494 586220 448458
rect 585620 411258 585802 411494
rect 586038 411258 586220 411494
rect 585620 374294 586220 411258
rect 585620 374058 585802 374294
rect 586038 374058 586220 374294
rect 585620 337094 586220 374058
rect 585620 336858 585802 337094
rect 586038 336858 586220 337094
rect 585620 299894 586220 336858
rect 585620 299658 585802 299894
rect 586038 299658 586220 299894
rect 585620 262694 586220 299658
rect 585620 262458 585802 262694
rect 586038 262458 586220 262694
rect 585620 225494 586220 262458
rect 585620 225258 585802 225494
rect 586038 225258 586220 225494
rect 585620 188294 586220 225258
rect 585620 188058 585802 188294
rect 586038 188058 586220 188294
rect 585620 151094 586220 188058
rect 585620 150858 585802 151094
rect 586038 150858 586220 151094
rect 585620 113894 586220 150858
rect 585620 113658 585802 113894
rect 586038 113658 586220 113894
rect 585620 76694 586220 113658
rect 585620 76458 585802 76694
rect 586038 76458 586220 76694
rect 585620 39494 586220 76458
rect 585620 39258 585802 39494
rect 586038 39258 586220 39494
rect 585620 2294 586220 39258
rect 585620 2058 585802 2294
rect 586038 2058 586220 2294
rect 585620 -806 586220 2058
rect 585620 -1042 585802 -806
rect 586038 -1042 586220 -806
rect 585620 -1224 586220 -1042
rect 586560 675494 587160 705682
rect 586560 675258 586742 675494
rect 586978 675258 587160 675494
rect 586560 638294 587160 675258
rect 586560 638058 586742 638294
rect 586978 638058 587160 638294
rect 586560 601094 587160 638058
rect 586560 600858 586742 601094
rect 586978 600858 587160 601094
rect 586560 563894 587160 600858
rect 586560 563658 586742 563894
rect 586978 563658 587160 563894
rect 586560 526694 587160 563658
rect 586560 526458 586742 526694
rect 586978 526458 587160 526694
rect 586560 489494 587160 526458
rect 586560 489258 586742 489494
rect 586978 489258 587160 489494
rect 586560 452294 587160 489258
rect 586560 452058 586742 452294
rect 586978 452058 587160 452294
rect 586560 415094 587160 452058
rect 586560 414858 586742 415094
rect 586978 414858 587160 415094
rect 586560 377894 587160 414858
rect 586560 377658 586742 377894
rect 586978 377658 587160 377894
rect 586560 340694 587160 377658
rect 586560 340458 586742 340694
rect 586978 340458 587160 340694
rect 586560 303494 587160 340458
rect 586560 303258 586742 303494
rect 586978 303258 587160 303494
rect 586560 266294 587160 303258
rect 586560 266058 586742 266294
rect 586978 266058 587160 266294
rect 586560 229094 587160 266058
rect 586560 228858 586742 229094
rect 586978 228858 587160 229094
rect 586560 191894 587160 228858
rect 586560 191658 586742 191894
rect 586978 191658 587160 191894
rect 586560 154694 587160 191658
rect 586560 154458 586742 154694
rect 586978 154458 587160 154694
rect 586560 117494 587160 154458
rect 586560 117258 586742 117494
rect 586978 117258 587160 117494
rect 586560 80294 587160 117258
rect 586560 80058 586742 80294
rect 586978 80058 587160 80294
rect 586560 43094 587160 80058
rect 586560 42858 586742 43094
rect 586978 42858 587160 43094
rect 586560 5894 587160 42858
rect 586560 5658 586742 5894
rect 586978 5658 587160 5894
rect 562404 -1982 562586 -1746
rect 562822 -1982 563004 -1746
rect 562404 -2164 563004 -1982
rect 586560 -1746 587160 5658
rect 586560 -1982 586742 -1746
rect 586978 -1982 587160 -1746
rect 586560 -2164 587160 -1982
<< via4 >>
rect -3054 705682 -2818 705918
rect -3054 675258 -2818 675494
rect -3054 638058 -2818 638294
rect -3054 600858 -2818 601094
rect -3054 563658 -2818 563894
rect -3054 526458 -2818 526694
rect -3054 489258 -2818 489494
rect -3054 452058 -2818 452294
rect -3054 414858 -2818 415094
rect -3054 377658 -2818 377894
rect -3054 340458 -2818 340694
rect -3054 303258 -2818 303494
rect -3054 266058 -2818 266294
rect -3054 228858 -2818 229094
rect -3054 191658 -2818 191894
rect -3054 154458 -2818 154694
rect -3054 117258 -2818 117494
rect -3054 80058 -2818 80294
rect -3054 42858 -2818 43094
rect -3054 5658 -2818 5894
rect -2114 704742 -1878 704978
rect -2114 671658 -1878 671894
rect -2114 634458 -1878 634694
rect -2114 597258 -1878 597494
rect -2114 560058 -1878 560294
rect -2114 522858 -1878 523094
rect -2114 485658 -1878 485894
rect -2114 448458 -1878 448694
rect -2114 411258 -1878 411494
rect -2114 374058 -1878 374294
rect -2114 336858 -1878 337094
rect -2114 299658 -1878 299894
rect -2114 262458 -1878 262694
rect -2114 225258 -1878 225494
rect -2114 188058 -1878 188294
rect -2114 150858 -1878 151094
rect -2114 113658 -1878 113894
rect -2114 76458 -1878 76694
rect -2114 39258 -1878 39494
rect -2114 2058 -1878 2294
rect -2114 -1042 -1878 -806
rect 986 704742 1222 704978
rect 986 671658 1222 671894
rect 986 634458 1222 634694
rect 986 597258 1222 597494
rect 986 560058 1222 560294
rect 986 522858 1222 523094
rect 986 485658 1222 485894
rect 986 448458 1222 448694
rect 986 411258 1222 411494
rect 986 374058 1222 374294
rect 986 336858 1222 337094
rect 986 299658 1222 299894
rect 986 262458 1222 262694
rect 986 225258 1222 225494
rect 986 188058 1222 188294
rect 986 150858 1222 151094
rect 986 113658 1222 113894
rect 986 76458 1222 76694
rect 986 39258 1222 39494
rect 986 2058 1222 2294
rect 986 -1042 1222 -806
rect -3054 -1982 -2818 -1746
rect 4586 705682 4822 705918
rect 4586 675258 4822 675494
rect 4586 638058 4822 638294
rect 4586 600858 4822 601094
rect 4586 563658 4822 563894
rect 4586 526458 4822 526694
rect 4586 489258 4822 489494
rect 4586 452058 4822 452294
rect 4586 414858 4822 415094
rect 4586 377658 4822 377894
rect 4586 340458 4822 340694
rect 4586 303258 4822 303494
rect 4586 266058 4822 266294
rect 4586 228858 4822 229094
rect 4586 191658 4822 191894
rect 4586 154458 4822 154694
rect 4586 117258 4822 117494
rect 4586 80058 4822 80294
rect 4586 42858 4822 43094
rect 4586 5658 4822 5894
rect 4586 -1982 4822 -1746
rect 38186 704742 38422 704978
rect 38186 671658 38422 671894
rect 38186 634458 38422 634694
rect 38186 597258 38422 597494
rect 38186 560058 38422 560294
rect 38186 522858 38422 523094
rect 38186 485658 38422 485894
rect 38186 448458 38422 448694
rect 38186 411258 38422 411494
rect 38186 374058 38422 374294
rect 38186 336858 38422 337094
rect 38186 299658 38422 299894
rect 38186 262458 38422 262694
rect 38186 225258 38422 225494
rect 38186 188058 38422 188294
rect 38186 150858 38422 151094
rect 38186 113658 38422 113894
rect 38186 76458 38422 76694
rect 38186 39258 38422 39494
rect 38186 2058 38422 2294
rect 38186 -1042 38422 -806
rect 41786 705682 42022 705918
rect 41786 675258 42022 675494
rect 41786 638058 42022 638294
rect 41786 600858 42022 601094
rect 41786 563658 42022 563894
rect 41786 526458 42022 526694
rect 41786 489258 42022 489494
rect 41786 452058 42022 452294
rect 41786 414858 42022 415094
rect 41786 377658 42022 377894
rect 41786 340458 42022 340694
rect 41786 303258 42022 303494
rect 41786 266058 42022 266294
rect 41786 228858 42022 229094
rect 41786 191658 42022 191894
rect 41786 154458 42022 154694
rect 41786 117258 42022 117494
rect 41786 80058 42022 80294
rect 41786 42858 42022 43094
rect 41786 5658 42022 5894
rect 41786 -1982 42022 -1746
rect 75386 704742 75622 704978
rect 75386 671658 75622 671894
rect 75386 634458 75622 634694
rect 75386 597258 75622 597494
rect 75386 560058 75622 560294
rect 75386 522858 75622 523094
rect 75386 485658 75622 485894
rect 75386 448458 75622 448694
rect 75386 411258 75622 411494
rect 75386 374058 75622 374294
rect 75386 336858 75622 337094
rect 75386 299658 75622 299894
rect 75386 262458 75622 262694
rect 75386 225258 75622 225494
rect 75386 188058 75622 188294
rect 75386 150858 75622 151094
rect 75386 113658 75622 113894
rect 75386 76458 75622 76694
rect 75386 39258 75622 39494
rect 75386 2058 75622 2294
rect 75386 -1042 75622 -806
rect 78986 705682 79222 705918
rect 78986 675258 79222 675494
rect 78986 638058 79222 638294
rect 78986 600858 79222 601094
rect 78986 563658 79222 563894
rect 78986 526458 79222 526694
rect 78986 489258 79222 489494
rect 78986 452058 79222 452294
rect 78986 414858 79222 415094
rect 78986 377658 79222 377894
rect 78986 340458 79222 340694
rect 78986 303258 79222 303494
rect 78986 266058 79222 266294
rect 78986 228858 79222 229094
rect 78986 191658 79222 191894
rect 78986 154458 79222 154694
rect 78986 117258 79222 117494
rect 78986 80058 79222 80294
rect 78986 42858 79222 43094
rect 78986 5658 79222 5894
rect 78986 -1982 79222 -1746
rect 112586 704742 112822 704978
rect 112586 671658 112822 671894
rect 112586 634458 112822 634694
rect 112586 597258 112822 597494
rect 112586 560058 112822 560294
rect 112586 522858 112822 523094
rect 112586 485658 112822 485894
rect 112586 448458 112822 448694
rect 112586 411258 112822 411494
rect 112586 374058 112822 374294
rect 112586 336858 112822 337094
rect 112586 299658 112822 299894
rect 112586 262458 112822 262694
rect 112586 225258 112822 225494
rect 112586 188058 112822 188294
rect 112586 150858 112822 151094
rect 112586 113658 112822 113894
rect 112586 76458 112822 76694
rect 112586 39258 112822 39494
rect 112586 2058 112822 2294
rect 112586 -1042 112822 -806
rect 116186 705682 116422 705918
rect 116186 675258 116422 675494
rect 116186 638058 116422 638294
rect 116186 600858 116422 601094
rect 116186 563658 116422 563894
rect 116186 526458 116422 526694
rect 116186 489258 116422 489494
rect 116186 452058 116422 452294
rect 116186 414858 116422 415094
rect 116186 377658 116422 377894
rect 116186 340458 116422 340694
rect 116186 303258 116422 303494
rect 116186 266058 116422 266294
rect 116186 228858 116422 229094
rect 116186 191658 116422 191894
rect 116186 154458 116422 154694
rect 116186 117258 116422 117494
rect 116186 80058 116422 80294
rect 116186 42858 116422 43094
rect 116186 5658 116422 5894
rect 116186 -1982 116422 -1746
rect 149786 704742 150022 704978
rect 149786 671658 150022 671894
rect 149786 634458 150022 634694
rect 149786 597258 150022 597494
rect 149786 560058 150022 560294
rect 149786 522858 150022 523094
rect 149786 485658 150022 485894
rect 149786 448458 150022 448694
rect 149786 411258 150022 411494
rect 149786 374058 150022 374294
rect 149786 336858 150022 337094
rect 149786 299658 150022 299894
rect 149786 262458 150022 262694
rect 149786 225258 150022 225494
rect 149786 188058 150022 188294
rect 149786 150858 150022 151094
rect 149786 113658 150022 113894
rect 149786 76458 150022 76694
rect 149786 39258 150022 39494
rect 149786 2058 150022 2294
rect 149786 -1042 150022 -806
rect 153386 705682 153622 705918
rect 153386 675258 153622 675494
rect 153386 638058 153622 638294
rect 153386 600858 153622 601094
rect 153386 563658 153622 563894
rect 153386 526458 153622 526694
rect 153386 489258 153622 489494
rect 153386 452058 153622 452294
rect 153386 414858 153622 415094
rect 153386 377658 153622 377894
rect 153386 340458 153622 340694
rect 153386 303258 153622 303494
rect 153386 266058 153622 266294
rect 153386 228858 153622 229094
rect 153386 191658 153622 191894
rect 153386 154458 153622 154694
rect 153386 117258 153622 117494
rect 153386 80058 153622 80294
rect 153386 42858 153622 43094
rect 153386 5658 153622 5894
rect 153386 -1982 153622 -1746
rect 186986 704742 187222 704978
rect 186986 671658 187222 671894
rect 186986 634458 187222 634694
rect 186986 597258 187222 597494
rect 186986 560058 187222 560294
rect 186986 522858 187222 523094
rect 186986 485658 187222 485894
rect 186986 448458 187222 448694
rect 186986 411258 187222 411494
rect 186986 374058 187222 374294
rect 186986 336858 187222 337094
rect 186986 299658 187222 299894
rect 186986 262458 187222 262694
rect 186986 225258 187222 225494
rect 186986 188058 187222 188294
rect 186986 150858 187222 151094
rect 186986 113658 187222 113894
rect 186986 76458 187222 76694
rect 186986 39258 187222 39494
rect 186986 2058 187222 2294
rect 186986 -1042 187222 -806
rect 190586 705682 190822 705918
rect 190586 675258 190822 675494
rect 190586 638058 190822 638294
rect 190586 600858 190822 601094
rect 190586 563658 190822 563894
rect 190586 526458 190822 526694
rect 190586 489258 190822 489494
rect 190586 452058 190822 452294
rect 190586 414858 190822 415094
rect 190586 377658 190822 377894
rect 190586 340458 190822 340694
rect 190586 303258 190822 303494
rect 190586 266058 190822 266294
rect 190586 228858 190822 229094
rect 190586 191658 190822 191894
rect 190586 154458 190822 154694
rect 190586 117258 190822 117494
rect 190586 80058 190822 80294
rect 190586 42858 190822 43094
rect 190586 5658 190822 5894
rect 190586 -1982 190822 -1746
rect 224186 704742 224422 704978
rect 224186 671658 224422 671894
rect 224186 634458 224422 634694
rect 224186 597258 224422 597494
rect 224186 560058 224422 560294
rect 224186 522858 224422 523094
rect 224186 485658 224422 485894
rect 224186 448458 224422 448694
rect 224186 411258 224422 411494
rect 224186 374058 224422 374294
rect 224186 336858 224422 337094
rect 224186 299658 224422 299894
rect 224186 262458 224422 262694
rect 224186 225258 224422 225494
rect 224186 188058 224422 188294
rect 224186 150858 224422 151094
rect 224186 113658 224422 113894
rect 224186 76458 224422 76694
rect 224186 39258 224422 39494
rect 224186 2058 224422 2294
rect 224186 -1042 224422 -806
rect 227786 705682 228022 705918
rect 227786 675258 228022 675494
rect 227786 638058 228022 638294
rect 227786 600858 228022 601094
rect 227786 563658 228022 563894
rect 227786 526458 228022 526694
rect 227786 489258 228022 489494
rect 227786 452058 228022 452294
rect 227786 414858 228022 415094
rect 227786 377658 228022 377894
rect 227786 340458 228022 340694
rect 227786 303258 228022 303494
rect 227786 266058 228022 266294
rect 227786 228858 228022 229094
rect 227786 191658 228022 191894
rect 227786 154458 228022 154694
rect 227786 117258 228022 117494
rect 227786 80058 228022 80294
rect 227786 42858 228022 43094
rect 227786 5658 228022 5894
rect 227786 -1982 228022 -1746
rect 261386 704742 261622 704978
rect 261386 671658 261622 671894
rect 261386 634458 261622 634694
rect 261386 597258 261622 597494
rect 261386 560058 261622 560294
rect 261386 522858 261622 523094
rect 261386 485658 261622 485894
rect 261386 448458 261622 448694
rect 261386 411258 261622 411494
rect 261386 374058 261622 374294
rect 261386 336858 261622 337094
rect 261386 299658 261622 299894
rect 261386 262458 261622 262694
rect 261386 225258 261622 225494
rect 261386 188058 261622 188294
rect 261386 150858 261622 151094
rect 261386 113658 261622 113894
rect 261386 76458 261622 76694
rect 261386 39258 261622 39494
rect 261386 2058 261622 2294
rect 261386 -1042 261622 -806
rect 264986 705682 265222 705918
rect 264986 675258 265222 675494
rect 264986 638058 265222 638294
rect 264986 600858 265222 601094
rect 264986 563658 265222 563894
rect 264986 526458 265222 526694
rect 298586 704742 298822 704978
rect 298586 671658 298822 671894
rect 298586 634458 298822 634694
rect 298586 597258 298822 597494
rect 298586 560058 298822 560294
rect 298586 522858 298822 523094
rect 264986 489258 265222 489494
rect 264986 452058 265222 452294
rect 264986 414858 265222 415094
rect 302186 705682 302422 705918
rect 302186 675258 302422 675494
rect 302186 638058 302422 638294
rect 302186 600858 302422 601094
rect 302186 563658 302422 563894
rect 302186 526458 302422 526694
rect 298586 485658 298822 485894
rect 298586 448458 298822 448694
rect 298586 411258 298822 411494
rect 335786 704742 336022 704978
rect 335786 671658 336022 671894
rect 335786 634458 336022 634694
rect 335786 597258 336022 597494
rect 335786 560058 336022 560294
rect 335786 522858 336022 523094
rect 302186 489258 302422 489494
rect 302186 452058 302422 452294
rect 264986 377658 265222 377894
rect 302186 414858 302422 415094
rect 298586 374058 298822 374294
rect 302186 377658 302422 377894
rect 264986 340458 265222 340694
rect 264986 303258 265222 303494
rect 298586 336858 298822 337094
rect 298586 299658 298822 299894
rect 264986 266058 265222 266294
rect 302186 340458 302422 340694
rect 302186 303258 302422 303494
rect 298586 262458 298822 262694
rect 264986 228858 265222 229094
rect 335786 485658 336022 485894
rect 335786 448458 336022 448694
rect 335786 411258 336022 411494
rect 335786 374058 336022 374294
rect 335786 336858 336022 337094
rect 335786 299658 336022 299894
rect 302186 266058 302422 266294
rect 298586 225258 298822 225494
rect 335786 262458 336022 262694
rect 302186 228858 302422 229094
rect 335786 225258 336022 225494
rect 264986 191658 265222 191894
rect 264986 154458 265222 154694
rect 264986 117258 265222 117494
rect 264986 80058 265222 80294
rect 264986 42858 265222 43094
rect 298586 188058 298822 188294
rect 298586 150858 298822 151094
rect 298586 113658 298822 113894
rect 298586 76458 298822 76694
rect 298586 39258 298822 39494
rect 264986 5658 265222 5894
rect 264986 -1982 265222 -1746
rect 298586 2058 298822 2294
rect 298586 -1042 298822 -806
rect 302186 191658 302422 191894
rect 302186 154458 302422 154694
rect 302186 117258 302422 117494
rect 335786 188058 336022 188294
rect 335786 150858 336022 151094
rect 335786 113658 336022 113894
rect 302186 80058 302422 80294
rect 302186 42858 302422 43094
rect 302186 5658 302422 5894
rect 302186 -1982 302422 -1746
rect 335786 76458 336022 76694
rect 335786 39258 336022 39494
rect 335786 2058 336022 2294
rect 335786 -1042 336022 -806
rect 339386 705682 339622 705918
rect 339386 675258 339622 675494
rect 339386 638058 339622 638294
rect 339386 600858 339622 601094
rect 339386 563658 339622 563894
rect 339386 526458 339622 526694
rect 339386 489258 339622 489494
rect 339386 452058 339622 452294
rect 339386 414858 339622 415094
rect 339386 377658 339622 377894
rect 339386 340458 339622 340694
rect 339386 303258 339622 303494
rect 339386 266058 339622 266294
rect 339386 228858 339622 229094
rect 339386 191658 339622 191894
rect 339386 154458 339622 154694
rect 339386 117258 339622 117494
rect 339386 80058 339622 80294
rect 339386 42858 339622 43094
rect 339386 5658 339622 5894
rect 339386 -1982 339622 -1746
rect 372986 704742 373222 704978
rect 372986 671658 373222 671894
rect 372986 634458 373222 634694
rect 372986 597258 373222 597494
rect 372986 560058 373222 560294
rect 372986 522858 373222 523094
rect 372986 485658 373222 485894
rect 372986 448458 373222 448694
rect 372986 411258 373222 411494
rect 372986 374058 373222 374294
rect 372986 336858 373222 337094
rect 372986 299658 373222 299894
rect 372986 262458 373222 262694
rect 372986 225258 373222 225494
rect 372986 188058 373222 188294
rect 372986 150858 373222 151094
rect 372986 113658 373222 113894
rect 372986 76458 373222 76694
rect 372986 39258 373222 39494
rect 372986 2058 373222 2294
rect 372986 -1042 373222 -806
rect 376586 705682 376822 705918
rect 376586 675258 376822 675494
rect 376586 638058 376822 638294
rect 376586 600858 376822 601094
rect 376586 563658 376822 563894
rect 376586 526458 376822 526694
rect 376586 489258 376822 489494
rect 376586 452058 376822 452294
rect 376586 414858 376822 415094
rect 376586 377658 376822 377894
rect 376586 340458 376822 340694
rect 376586 303258 376822 303494
rect 376586 266058 376822 266294
rect 376586 228858 376822 229094
rect 376586 191658 376822 191894
rect 376586 154458 376822 154694
rect 376586 117258 376822 117494
rect 376586 80058 376822 80294
rect 376586 42858 376822 43094
rect 376586 5658 376822 5894
rect 376586 -1982 376822 -1746
rect 410186 704742 410422 704978
rect 410186 671658 410422 671894
rect 410186 634458 410422 634694
rect 410186 597258 410422 597494
rect 410186 560058 410422 560294
rect 410186 522858 410422 523094
rect 410186 485658 410422 485894
rect 410186 448458 410422 448694
rect 410186 411258 410422 411494
rect 410186 374058 410422 374294
rect 410186 336858 410422 337094
rect 410186 299658 410422 299894
rect 410186 262458 410422 262694
rect 410186 225258 410422 225494
rect 410186 188058 410422 188294
rect 410186 150858 410422 151094
rect 410186 113658 410422 113894
rect 410186 76458 410422 76694
rect 410186 39258 410422 39494
rect 410186 2058 410422 2294
rect 410186 -1042 410422 -806
rect 413786 705682 414022 705918
rect 413786 675258 414022 675494
rect 413786 638058 414022 638294
rect 413786 600858 414022 601094
rect 413786 563658 414022 563894
rect 413786 526458 414022 526694
rect 413786 489258 414022 489494
rect 413786 452058 414022 452294
rect 413786 414858 414022 415094
rect 413786 377658 414022 377894
rect 413786 340458 414022 340694
rect 413786 303258 414022 303494
rect 413786 266058 414022 266294
rect 413786 228858 414022 229094
rect 413786 191658 414022 191894
rect 413786 154458 414022 154694
rect 413786 117258 414022 117494
rect 413786 80058 414022 80294
rect 413786 42858 414022 43094
rect 413786 5658 414022 5894
rect 413786 -1982 414022 -1746
rect 447386 704742 447622 704978
rect 447386 671658 447622 671894
rect 447386 634458 447622 634694
rect 447386 597258 447622 597494
rect 447386 560058 447622 560294
rect 447386 522858 447622 523094
rect 447386 485658 447622 485894
rect 447386 448458 447622 448694
rect 447386 411258 447622 411494
rect 447386 374058 447622 374294
rect 447386 336858 447622 337094
rect 447386 299658 447622 299894
rect 447386 262458 447622 262694
rect 447386 225258 447622 225494
rect 447386 188058 447622 188294
rect 447386 150858 447622 151094
rect 447386 113658 447622 113894
rect 447386 76458 447622 76694
rect 447386 39258 447622 39494
rect 447386 2058 447622 2294
rect 447386 -1042 447622 -806
rect 450986 705682 451222 705918
rect 450986 675258 451222 675494
rect 450986 638058 451222 638294
rect 450986 600858 451222 601094
rect 450986 563658 451222 563894
rect 450986 526458 451222 526694
rect 450986 489258 451222 489494
rect 450986 452058 451222 452294
rect 450986 414858 451222 415094
rect 450986 377658 451222 377894
rect 450986 340458 451222 340694
rect 450986 303258 451222 303494
rect 450986 266058 451222 266294
rect 450986 228858 451222 229094
rect 450986 191658 451222 191894
rect 450986 154458 451222 154694
rect 450986 117258 451222 117494
rect 450986 80058 451222 80294
rect 450986 42858 451222 43094
rect 450986 5658 451222 5894
rect 450986 -1982 451222 -1746
rect 484586 704742 484822 704978
rect 484586 671658 484822 671894
rect 484586 634458 484822 634694
rect 484586 597258 484822 597494
rect 484586 560058 484822 560294
rect 484586 522858 484822 523094
rect 484586 485658 484822 485894
rect 484586 448458 484822 448694
rect 484586 411258 484822 411494
rect 484586 374058 484822 374294
rect 484586 336858 484822 337094
rect 484586 299658 484822 299894
rect 484586 262458 484822 262694
rect 484586 225258 484822 225494
rect 484586 188058 484822 188294
rect 484586 150858 484822 151094
rect 484586 113658 484822 113894
rect 484586 76458 484822 76694
rect 484586 39258 484822 39494
rect 484586 2058 484822 2294
rect 484586 -1042 484822 -806
rect 488186 705682 488422 705918
rect 488186 675258 488422 675494
rect 488186 638058 488422 638294
rect 488186 600858 488422 601094
rect 488186 563658 488422 563894
rect 488186 526458 488422 526694
rect 488186 489258 488422 489494
rect 488186 452058 488422 452294
rect 521786 704742 522022 704978
rect 521786 671658 522022 671894
rect 521786 634458 522022 634694
rect 521786 597258 522022 597494
rect 521786 560058 522022 560294
rect 521786 522858 522022 523094
rect 521786 485658 522022 485894
rect 521786 448458 522022 448694
rect 525386 705682 525622 705918
rect 525386 675258 525622 675494
rect 525386 638058 525622 638294
rect 525386 600858 525622 601094
rect 525386 563658 525622 563894
rect 525386 526458 525622 526694
rect 525386 489258 525622 489494
rect 525386 452058 525622 452294
rect 558986 704742 559222 704978
rect 558986 671658 559222 671894
rect 558986 634458 559222 634694
rect 558986 597258 559222 597494
rect 558986 560058 559222 560294
rect 558986 522858 559222 523094
rect 558986 485658 559222 485894
rect 558986 448458 559222 448694
rect 488186 414858 488422 415094
rect 558986 411258 559222 411494
rect 488186 377658 488422 377894
rect 558986 374058 559222 374294
rect 488186 340458 488422 340694
rect 488186 303258 488422 303494
rect 558986 336858 559222 337094
rect 488186 266058 488422 266294
rect 558986 299658 559222 299894
rect 558986 262458 559222 262694
rect 488186 228858 488422 229094
rect 488186 191658 488422 191894
rect 488186 154458 488422 154694
rect 488186 117258 488422 117494
rect 488186 80058 488422 80294
rect 488186 42858 488422 43094
rect 488186 5658 488422 5894
rect 488186 -1982 488422 -1746
rect 521786 225258 522022 225494
rect 521786 188058 522022 188294
rect 521786 150858 522022 151094
rect 521786 113658 522022 113894
rect 521786 76458 522022 76694
rect 521786 39258 522022 39494
rect 521786 2058 522022 2294
rect 521786 -1042 522022 -806
rect 525386 228858 525622 229094
rect 525386 191658 525622 191894
rect 525386 154458 525622 154694
rect 525386 117258 525622 117494
rect 525386 80058 525622 80294
rect 525386 42858 525622 43094
rect 558986 225258 559222 225494
rect 558986 188058 559222 188294
rect 558986 150858 559222 151094
rect 558986 113658 559222 113894
rect 558986 76458 559222 76694
rect 558986 39258 559222 39494
rect 525386 5658 525622 5894
rect 525386 -1982 525622 -1746
rect 558986 2058 559222 2294
rect 558986 -1042 559222 -806
rect 562586 705682 562822 705918
rect 586742 705682 586978 705918
rect 562586 675258 562822 675494
rect 562586 638058 562822 638294
rect 562586 600858 562822 601094
rect 562586 563658 562822 563894
rect 562586 526458 562822 526694
rect 562586 489258 562822 489494
rect 562586 452058 562822 452294
rect 562586 414858 562822 415094
rect 562586 377658 562822 377894
rect 562586 340458 562822 340694
rect 562586 303258 562822 303494
rect 562586 266058 562822 266294
rect 562586 228858 562822 229094
rect 562586 191658 562822 191894
rect 562586 154458 562822 154694
rect 562586 117258 562822 117494
rect 562586 80058 562822 80294
rect 562586 42858 562822 43094
rect 562586 5658 562822 5894
rect 585802 704742 586038 704978
rect 585802 671658 586038 671894
rect 585802 634458 586038 634694
rect 585802 597258 586038 597494
rect 585802 560058 586038 560294
rect 585802 522858 586038 523094
rect 585802 485658 586038 485894
rect 585802 448458 586038 448694
rect 585802 411258 586038 411494
rect 585802 374058 586038 374294
rect 585802 336858 586038 337094
rect 585802 299658 586038 299894
rect 585802 262458 586038 262694
rect 585802 225258 586038 225494
rect 585802 188058 586038 188294
rect 585802 150858 586038 151094
rect 585802 113658 586038 113894
rect 585802 76458 586038 76694
rect 585802 39258 586038 39494
rect 585802 2058 586038 2294
rect 585802 -1042 586038 -806
rect 586742 675258 586978 675494
rect 586742 638058 586978 638294
rect 586742 600858 586978 601094
rect 586742 563658 586978 563894
rect 586742 526458 586978 526694
rect 586742 489258 586978 489494
rect 586742 452058 586978 452294
rect 586742 414858 586978 415094
rect 586742 377658 586978 377894
rect 586742 340458 586978 340694
rect 586742 303258 586978 303494
rect 586742 266058 586978 266294
rect 586742 228858 586978 229094
rect 586742 191658 586978 191894
rect 586742 154458 586978 154694
rect 586742 117258 586978 117494
rect 586742 80058 586978 80294
rect 586742 42858 586978 43094
rect 586742 5658 586978 5894
rect 562586 -1982 562822 -1746
rect 586742 -1982 586978 -1746
<< metal5 >>
rect -3236 705918 587160 706100
rect -3236 705682 -3054 705918
rect -2818 705682 4586 705918
rect 4822 705682 41786 705918
rect 42022 705682 78986 705918
rect 79222 705682 116186 705918
rect 116422 705682 153386 705918
rect 153622 705682 190586 705918
rect 190822 705682 227786 705918
rect 228022 705682 264986 705918
rect 265222 705682 302186 705918
rect 302422 705682 339386 705918
rect 339622 705682 376586 705918
rect 376822 705682 413786 705918
rect 414022 705682 450986 705918
rect 451222 705682 488186 705918
rect 488422 705682 525386 705918
rect 525622 705682 562586 705918
rect 562822 705682 586742 705918
rect 586978 705682 587160 705918
rect -3236 705500 587160 705682
rect -2296 704978 586220 705160
rect -2296 704742 -2114 704978
rect -1878 704742 986 704978
rect 1222 704742 38186 704978
rect 38422 704742 75386 704978
rect 75622 704742 112586 704978
rect 112822 704742 149786 704978
rect 150022 704742 186986 704978
rect 187222 704742 224186 704978
rect 224422 704742 261386 704978
rect 261622 704742 298586 704978
rect 298822 704742 335786 704978
rect 336022 704742 372986 704978
rect 373222 704742 410186 704978
rect 410422 704742 447386 704978
rect 447622 704742 484586 704978
rect 484822 704742 521786 704978
rect 522022 704742 558986 704978
rect 559222 704742 585802 704978
rect 586038 704742 586220 704978
rect -2296 704560 586220 704742
rect -3236 675494 587160 675676
rect -3236 675258 -3054 675494
rect -2818 675258 4586 675494
rect 4822 675258 41786 675494
rect 42022 675258 78986 675494
rect 79222 675258 116186 675494
rect 116422 675258 153386 675494
rect 153622 675258 190586 675494
rect 190822 675258 227786 675494
rect 228022 675258 264986 675494
rect 265222 675258 302186 675494
rect 302422 675258 339386 675494
rect 339622 675258 376586 675494
rect 376822 675258 413786 675494
rect 414022 675258 450986 675494
rect 451222 675258 488186 675494
rect 488422 675258 525386 675494
rect 525622 675258 562586 675494
rect 562822 675258 586742 675494
rect 586978 675258 587160 675494
rect -3236 675076 587160 675258
rect -3236 671894 587160 672076
rect -3236 671658 -2114 671894
rect -1878 671658 986 671894
rect 1222 671658 38186 671894
rect 38422 671658 75386 671894
rect 75622 671658 112586 671894
rect 112822 671658 149786 671894
rect 150022 671658 186986 671894
rect 187222 671658 224186 671894
rect 224422 671658 261386 671894
rect 261622 671658 298586 671894
rect 298822 671658 335786 671894
rect 336022 671658 372986 671894
rect 373222 671658 410186 671894
rect 410422 671658 447386 671894
rect 447622 671658 484586 671894
rect 484822 671658 521786 671894
rect 522022 671658 558986 671894
rect 559222 671658 585802 671894
rect 586038 671658 587160 671894
rect -3236 671476 587160 671658
rect -3236 638294 587160 638476
rect -3236 638058 -3054 638294
rect -2818 638058 4586 638294
rect 4822 638058 41786 638294
rect 42022 638058 78986 638294
rect 79222 638058 116186 638294
rect 116422 638058 153386 638294
rect 153622 638058 190586 638294
rect 190822 638058 227786 638294
rect 228022 638058 264986 638294
rect 265222 638058 302186 638294
rect 302422 638058 339386 638294
rect 339622 638058 376586 638294
rect 376822 638058 413786 638294
rect 414022 638058 450986 638294
rect 451222 638058 488186 638294
rect 488422 638058 525386 638294
rect 525622 638058 562586 638294
rect 562822 638058 586742 638294
rect 586978 638058 587160 638294
rect -3236 637876 587160 638058
rect -3236 634694 587160 634876
rect -3236 634458 -2114 634694
rect -1878 634458 986 634694
rect 1222 634458 38186 634694
rect 38422 634458 75386 634694
rect 75622 634458 112586 634694
rect 112822 634458 149786 634694
rect 150022 634458 186986 634694
rect 187222 634458 224186 634694
rect 224422 634458 261386 634694
rect 261622 634458 298586 634694
rect 298822 634458 335786 634694
rect 336022 634458 372986 634694
rect 373222 634458 410186 634694
rect 410422 634458 447386 634694
rect 447622 634458 484586 634694
rect 484822 634458 521786 634694
rect 522022 634458 558986 634694
rect 559222 634458 585802 634694
rect 586038 634458 587160 634694
rect -3236 634276 587160 634458
rect -3236 601094 587160 601276
rect -3236 600858 -3054 601094
rect -2818 600858 4586 601094
rect 4822 600858 41786 601094
rect 42022 600858 78986 601094
rect 79222 600858 116186 601094
rect 116422 600858 153386 601094
rect 153622 600858 190586 601094
rect 190822 600858 227786 601094
rect 228022 600858 264986 601094
rect 265222 600858 302186 601094
rect 302422 600858 339386 601094
rect 339622 600858 376586 601094
rect 376822 600858 413786 601094
rect 414022 600858 450986 601094
rect 451222 600858 488186 601094
rect 488422 600858 525386 601094
rect 525622 600858 562586 601094
rect 562822 600858 586742 601094
rect 586978 600858 587160 601094
rect -3236 600676 587160 600858
rect -3236 597494 587160 597676
rect -3236 597258 -2114 597494
rect -1878 597258 986 597494
rect 1222 597258 38186 597494
rect 38422 597258 75386 597494
rect 75622 597258 112586 597494
rect 112822 597258 149786 597494
rect 150022 597258 186986 597494
rect 187222 597258 224186 597494
rect 224422 597258 261386 597494
rect 261622 597258 298586 597494
rect 298822 597258 335786 597494
rect 336022 597258 372986 597494
rect 373222 597258 410186 597494
rect 410422 597258 447386 597494
rect 447622 597258 484586 597494
rect 484822 597258 521786 597494
rect 522022 597258 558986 597494
rect 559222 597258 585802 597494
rect 586038 597258 587160 597494
rect -3236 597076 587160 597258
rect -3236 563894 587160 564076
rect -3236 563658 -3054 563894
rect -2818 563658 4586 563894
rect 4822 563658 41786 563894
rect 42022 563658 78986 563894
rect 79222 563658 116186 563894
rect 116422 563658 153386 563894
rect 153622 563658 190586 563894
rect 190822 563658 227786 563894
rect 228022 563658 264986 563894
rect 265222 563658 302186 563894
rect 302422 563658 339386 563894
rect 339622 563658 376586 563894
rect 376822 563658 413786 563894
rect 414022 563658 450986 563894
rect 451222 563658 488186 563894
rect 488422 563658 525386 563894
rect 525622 563658 562586 563894
rect 562822 563658 586742 563894
rect 586978 563658 587160 563894
rect -3236 563476 587160 563658
rect -3236 560294 587160 560476
rect -3236 560058 -2114 560294
rect -1878 560058 986 560294
rect 1222 560058 38186 560294
rect 38422 560058 75386 560294
rect 75622 560058 112586 560294
rect 112822 560058 149786 560294
rect 150022 560058 186986 560294
rect 187222 560058 224186 560294
rect 224422 560058 261386 560294
rect 261622 560058 298586 560294
rect 298822 560058 335786 560294
rect 336022 560058 372986 560294
rect 373222 560058 410186 560294
rect 410422 560058 447386 560294
rect 447622 560058 484586 560294
rect 484822 560058 521786 560294
rect 522022 560058 558986 560294
rect 559222 560058 585802 560294
rect 586038 560058 587160 560294
rect -3236 559876 587160 560058
rect -3236 526694 587160 526876
rect -3236 526458 -3054 526694
rect -2818 526458 4586 526694
rect 4822 526458 41786 526694
rect 42022 526458 78986 526694
rect 79222 526458 116186 526694
rect 116422 526458 153386 526694
rect 153622 526458 190586 526694
rect 190822 526458 227786 526694
rect 228022 526458 264986 526694
rect 265222 526458 302186 526694
rect 302422 526458 339386 526694
rect 339622 526458 376586 526694
rect 376822 526458 413786 526694
rect 414022 526458 450986 526694
rect 451222 526458 488186 526694
rect 488422 526458 525386 526694
rect 525622 526458 562586 526694
rect 562822 526458 586742 526694
rect 586978 526458 587160 526694
rect -3236 526276 587160 526458
rect -3236 523094 587160 523276
rect -3236 522858 -2114 523094
rect -1878 522858 986 523094
rect 1222 522858 38186 523094
rect 38422 522858 75386 523094
rect 75622 522858 112586 523094
rect 112822 522858 149786 523094
rect 150022 522858 186986 523094
rect 187222 522858 224186 523094
rect 224422 522858 261386 523094
rect 261622 522858 298586 523094
rect 298822 522858 335786 523094
rect 336022 522858 372986 523094
rect 373222 522858 410186 523094
rect 410422 522858 447386 523094
rect 447622 522858 484586 523094
rect 484822 522858 521786 523094
rect 522022 522858 558986 523094
rect 559222 522858 585802 523094
rect 586038 522858 587160 523094
rect -3236 522676 587160 522858
rect -3236 489494 587160 489676
rect -3236 489258 -3054 489494
rect -2818 489258 4586 489494
rect 4822 489258 41786 489494
rect 42022 489258 78986 489494
rect 79222 489258 116186 489494
rect 116422 489258 153386 489494
rect 153622 489258 190586 489494
rect 190822 489258 227786 489494
rect 228022 489258 264986 489494
rect 265222 489258 302186 489494
rect 302422 489258 339386 489494
rect 339622 489258 376586 489494
rect 376822 489258 413786 489494
rect 414022 489258 450986 489494
rect 451222 489258 488186 489494
rect 488422 489258 525386 489494
rect 525622 489258 562586 489494
rect 562822 489258 586742 489494
rect 586978 489258 587160 489494
rect -3236 489076 587160 489258
rect -3236 485894 587160 486076
rect -3236 485658 -2114 485894
rect -1878 485658 986 485894
rect 1222 485658 38186 485894
rect 38422 485658 75386 485894
rect 75622 485658 112586 485894
rect 112822 485658 149786 485894
rect 150022 485658 186986 485894
rect 187222 485658 224186 485894
rect 224422 485658 261386 485894
rect 261622 485658 298586 485894
rect 298822 485658 335786 485894
rect 336022 485658 372986 485894
rect 373222 485658 410186 485894
rect 410422 485658 447386 485894
rect 447622 485658 484586 485894
rect 484822 485658 521786 485894
rect 522022 485658 558986 485894
rect 559222 485658 585802 485894
rect 586038 485658 587160 485894
rect -3236 485476 587160 485658
rect -3236 452294 587160 452476
rect -3236 452058 -3054 452294
rect -2818 452058 4586 452294
rect 4822 452058 41786 452294
rect 42022 452058 78986 452294
rect 79222 452058 116186 452294
rect 116422 452058 153386 452294
rect 153622 452058 190586 452294
rect 190822 452058 227786 452294
rect 228022 452058 264986 452294
rect 265222 452058 302186 452294
rect 302422 452058 339386 452294
rect 339622 452058 376586 452294
rect 376822 452058 413786 452294
rect 414022 452058 450986 452294
rect 451222 452058 488186 452294
rect 488422 452058 525386 452294
rect 525622 452058 562586 452294
rect 562822 452058 586742 452294
rect 586978 452058 587160 452294
rect -3236 451876 587160 452058
rect -3236 448694 587160 448876
rect -3236 448458 -2114 448694
rect -1878 448458 986 448694
rect 1222 448458 38186 448694
rect 38422 448458 75386 448694
rect 75622 448458 112586 448694
rect 112822 448458 149786 448694
rect 150022 448458 186986 448694
rect 187222 448458 224186 448694
rect 224422 448458 261386 448694
rect 261622 448458 298586 448694
rect 298822 448458 335786 448694
rect 336022 448458 372986 448694
rect 373222 448458 410186 448694
rect 410422 448458 447386 448694
rect 447622 448458 484586 448694
rect 484822 448458 521786 448694
rect 522022 448458 558986 448694
rect 559222 448458 585802 448694
rect 586038 448458 587160 448694
rect -3236 448276 587160 448458
rect -3236 415094 587160 415276
rect -3236 414858 -3054 415094
rect -2818 414858 4586 415094
rect 4822 414858 41786 415094
rect 42022 414858 78986 415094
rect 79222 414858 116186 415094
rect 116422 414858 153386 415094
rect 153622 414858 190586 415094
rect 190822 414858 227786 415094
rect 228022 414858 264986 415094
rect 265222 414858 302186 415094
rect 302422 414858 339386 415094
rect 339622 414858 376586 415094
rect 376822 414858 413786 415094
rect 414022 414858 450986 415094
rect 451222 414858 488186 415094
rect 488422 414858 562586 415094
rect 562822 414858 586742 415094
rect 586978 414858 587160 415094
rect -3236 414676 587160 414858
rect -3236 411494 587160 411676
rect -3236 411258 -2114 411494
rect -1878 411258 986 411494
rect 1222 411258 38186 411494
rect 38422 411258 75386 411494
rect 75622 411258 112586 411494
rect 112822 411258 149786 411494
rect 150022 411258 186986 411494
rect 187222 411258 224186 411494
rect 224422 411258 261386 411494
rect 261622 411258 298586 411494
rect 298822 411258 335786 411494
rect 336022 411258 372986 411494
rect 373222 411258 410186 411494
rect 410422 411258 447386 411494
rect 447622 411258 484586 411494
rect 484822 411258 558986 411494
rect 559222 411258 585802 411494
rect 586038 411258 587160 411494
rect -3236 411076 587160 411258
rect -3236 377894 587160 378076
rect -3236 377658 -3054 377894
rect -2818 377658 4586 377894
rect 4822 377658 41786 377894
rect 42022 377658 78986 377894
rect 79222 377658 116186 377894
rect 116422 377658 153386 377894
rect 153622 377658 190586 377894
rect 190822 377658 227786 377894
rect 228022 377658 264986 377894
rect 265222 377658 302186 377894
rect 302422 377658 339386 377894
rect 339622 377658 376586 377894
rect 376822 377658 413786 377894
rect 414022 377658 450986 377894
rect 451222 377658 488186 377894
rect 488422 377658 562586 377894
rect 562822 377658 586742 377894
rect 586978 377658 587160 377894
rect -3236 377476 587160 377658
rect -3236 374294 587160 374476
rect -3236 374058 -2114 374294
rect -1878 374058 986 374294
rect 1222 374058 38186 374294
rect 38422 374058 75386 374294
rect 75622 374058 112586 374294
rect 112822 374058 149786 374294
rect 150022 374058 186986 374294
rect 187222 374058 224186 374294
rect 224422 374058 261386 374294
rect 261622 374058 298586 374294
rect 298822 374058 335786 374294
rect 336022 374058 372986 374294
rect 373222 374058 410186 374294
rect 410422 374058 447386 374294
rect 447622 374058 484586 374294
rect 484822 374058 558986 374294
rect 559222 374058 585802 374294
rect 586038 374058 587160 374294
rect -3236 373876 587160 374058
rect -3236 340694 587160 340876
rect -3236 340458 -3054 340694
rect -2818 340458 4586 340694
rect 4822 340458 41786 340694
rect 42022 340458 78986 340694
rect 79222 340458 116186 340694
rect 116422 340458 153386 340694
rect 153622 340458 190586 340694
rect 190822 340458 227786 340694
rect 228022 340458 264986 340694
rect 265222 340458 302186 340694
rect 302422 340458 339386 340694
rect 339622 340458 376586 340694
rect 376822 340458 413786 340694
rect 414022 340458 450986 340694
rect 451222 340458 488186 340694
rect 488422 340458 562586 340694
rect 562822 340458 586742 340694
rect 586978 340458 587160 340694
rect -3236 340276 587160 340458
rect -3236 337094 587160 337276
rect -3236 336858 -2114 337094
rect -1878 336858 986 337094
rect 1222 336858 38186 337094
rect 38422 336858 75386 337094
rect 75622 336858 112586 337094
rect 112822 336858 149786 337094
rect 150022 336858 186986 337094
rect 187222 336858 224186 337094
rect 224422 336858 261386 337094
rect 261622 336858 298586 337094
rect 298822 336858 335786 337094
rect 336022 336858 372986 337094
rect 373222 336858 410186 337094
rect 410422 336858 447386 337094
rect 447622 336858 484586 337094
rect 484822 336858 558986 337094
rect 559222 336858 585802 337094
rect 586038 336858 587160 337094
rect -3236 336676 587160 336858
rect -3236 303494 587160 303676
rect -3236 303258 -3054 303494
rect -2818 303258 4586 303494
rect 4822 303258 41786 303494
rect 42022 303258 78986 303494
rect 79222 303258 116186 303494
rect 116422 303258 153386 303494
rect 153622 303258 190586 303494
rect 190822 303258 227786 303494
rect 228022 303258 264986 303494
rect 265222 303258 302186 303494
rect 302422 303258 339386 303494
rect 339622 303258 376586 303494
rect 376822 303258 413786 303494
rect 414022 303258 450986 303494
rect 451222 303258 488186 303494
rect 488422 303258 562586 303494
rect 562822 303258 586742 303494
rect 586978 303258 587160 303494
rect -3236 303076 587160 303258
rect -3236 299894 587160 300076
rect -3236 299658 -2114 299894
rect -1878 299658 986 299894
rect 1222 299658 38186 299894
rect 38422 299658 75386 299894
rect 75622 299658 112586 299894
rect 112822 299658 149786 299894
rect 150022 299658 186986 299894
rect 187222 299658 224186 299894
rect 224422 299658 261386 299894
rect 261622 299658 298586 299894
rect 298822 299658 335786 299894
rect 336022 299658 372986 299894
rect 373222 299658 410186 299894
rect 410422 299658 447386 299894
rect 447622 299658 484586 299894
rect 484822 299658 558986 299894
rect 559222 299658 585802 299894
rect 586038 299658 587160 299894
rect -3236 299476 587160 299658
rect -3236 266294 587160 266476
rect -3236 266058 -3054 266294
rect -2818 266058 4586 266294
rect 4822 266058 41786 266294
rect 42022 266058 78986 266294
rect 79222 266058 116186 266294
rect 116422 266058 153386 266294
rect 153622 266058 190586 266294
rect 190822 266058 227786 266294
rect 228022 266058 264986 266294
rect 265222 266058 302186 266294
rect 302422 266058 339386 266294
rect 339622 266058 376586 266294
rect 376822 266058 413786 266294
rect 414022 266058 450986 266294
rect 451222 266058 488186 266294
rect 488422 266058 562586 266294
rect 562822 266058 586742 266294
rect 586978 266058 587160 266294
rect -3236 265876 587160 266058
rect -3236 262694 587160 262876
rect -3236 262458 -2114 262694
rect -1878 262458 986 262694
rect 1222 262458 38186 262694
rect 38422 262458 75386 262694
rect 75622 262458 112586 262694
rect 112822 262458 149786 262694
rect 150022 262458 186986 262694
rect 187222 262458 224186 262694
rect 224422 262458 261386 262694
rect 261622 262458 298586 262694
rect 298822 262458 335786 262694
rect 336022 262458 372986 262694
rect 373222 262458 410186 262694
rect 410422 262458 447386 262694
rect 447622 262458 484586 262694
rect 484822 262458 558986 262694
rect 559222 262458 585802 262694
rect 586038 262458 587160 262694
rect -3236 262276 587160 262458
rect -3236 229094 587160 229276
rect -3236 228858 -3054 229094
rect -2818 228858 4586 229094
rect 4822 228858 41786 229094
rect 42022 228858 78986 229094
rect 79222 228858 116186 229094
rect 116422 228858 153386 229094
rect 153622 228858 190586 229094
rect 190822 228858 227786 229094
rect 228022 228858 264986 229094
rect 265222 228858 302186 229094
rect 302422 228858 339386 229094
rect 339622 228858 376586 229094
rect 376822 228858 413786 229094
rect 414022 228858 450986 229094
rect 451222 228858 488186 229094
rect 488422 228858 525386 229094
rect 525622 228858 562586 229094
rect 562822 228858 586742 229094
rect 586978 228858 587160 229094
rect -3236 228676 587160 228858
rect -3236 225494 587160 225676
rect -3236 225258 -2114 225494
rect -1878 225258 986 225494
rect 1222 225258 38186 225494
rect 38422 225258 75386 225494
rect 75622 225258 112586 225494
rect 112822 225258 149786 225494
rect 150022 225258 186986 225494
rect 187222 225258 224186 225494
rect 224422 225258 261386 225494
rect 261622 225258 298586 225494
rect 298822 225258 335786 225494
rect 336022 225258 372986 225494
rect 373222 225258 410186 225494
rect 410422 225258 447386 225494
rect 447622 225258 484586 225494
rect 484822 225258 521786 225494
rect 522022 225258 558986 225494
rect 559222 225258 585802 225494
rect 586038 225258 587160 225494
rect -3236 225076 587160 225258
rect -3236 191894 587160 192076
rect -3236 191658 -3054 191894
rect -2818 191658 4586 191894
rect 4822 191658 41786 191894
rect 42022 191658 78986 191894
rect 79222 191658 116186 191894
rect 116422 191658 153386 191894
rect 153622 191658 190586 191894
rect 190822 191658 227786 191894
rect 228022 191658 264986 191894
rect 265222 191658 302186 191894
rect 302422 191658 339386 191894
rect 339622 191658 376586 191894
rect 376822 191658 413786 191894
rect 414022 191658 450986 191894
rect 451222 191658 488186 191894
rect 488422 191658 525386 191894
rect 525622 191658 562586 191894
rect 562822 191658 586742 191894
rect 586978 191658 587160 191894
rect -3236 191476 587160 191658
rect -3236 188294 587160 188476
rect -3236 188058 -2114 188294
rect -1878 188058 986 188294
rect 1222 188058 38186 188294
rect 38422 188058 75386 188294
rect 75622 188058 112586 188294
rect 112822 188058 149786 188294
rect 150022 188058 186986 188294
rect 187222 188058 224186 188294
rect 224422 188058 261386 188294
rect 261622 188058 298586 188294
rect 298822 188058 335786 188294
rect 336022 188058 372986 188294
rect 373222 188058 410186 188294
rect 410422 188058 447386 188294
rect 447622 188058 484586 188294
rect 484822 188058 521786 188294
rect 522022 188058 558986 188294
rect 559222 188058 585802 188294
rect 586038 188058 587160 188294
rect -3236 187876 587160 188058
rect -3236 154694 587160 154876
rect -3236 154458 -3054 154694
rect -2818 154458 4586 154694
rect 4822 154458 41786 154694
rect 42022 154458 78986 154694
rect 79222 154458 116186 154694
rect 116422 154458 153386 154694
rect 153622 154458 190586 154694
rect 190822 154458 227786 154694
rect 228022 154458 264986 154694
rect 265222 154458 302186 154694
rect 302422 154458 339386 154694
rect 339622 154458 376586 154694
rect 376822 154458 413786 154694
rect 414022 154458 450986 154694
rect 451222 154458 488186 154694
rect 488422 154458 525386 154694
rect 525622 154458 562586 154694
rect 562822 154458 586742 154694
rect 586978 154458 587160 154694
rect -3236 154276 587160 154458
rect -3236 151094 587160 151276
rect -3236 150858 -2114 151094
rect -1878 150858 986 151094
rect 1222 150858 38186 151094
rect 38422 150858 75386 151094
rect 75622 150858 112586 151094
rect 112822 150858 149786 151094
rect 150022 150858 186986 151094
rect 187222 150858 224186 151094
rect 224422 150858 261386 151094
rect 261622 150858 298586 151094
rect 298822 150858 335786 151094
rect 336022 150858 372986 151094
rect 373222 150858 410186 151094
rect 410422 150858 447386 151094
rect 447622 150858 484586 151094
rect 484822 150858 521786 151094
rect 522022 150858 558986 151094
rect 559222 150858 585802 151094
rect 586038 150858 587160 151094
rect -3236 150676 587160 150858
rect -3236 117494 587160 117676
rect -3236 117258 -3054 117494
rect -2818 117258 4586 117494
rect 4822 117258 41786 117494
rect 42022 117258 78986 117494
rect 79222 117258 116186 117494
rect 116422 117258 153386 117494
rect 153622 117258 190586 117494
rect 190822 117258 227786 117494
rect 228022 117258 264986 117494
rect 265222 117258 302186 117494
rect 302422 117258 339386 117494
rect 339622 117258 376586 117494
rect 376822 117258 413786 117494
rect 414022 117258 450986 117494
rect 451222 117258 488186 117494
rect 488422 117258 525386 117494
rect 525622 117258 562586 117494
rect 562822 117258 586742 117494
rect 586978 117258 587160 117494
rect -3236 117076 587160 117258
rect -3236 113894 587160 114076
rect -3236 113658 -2114 113894
rect -1878 113658 986 113894
rect 1222 113658 38186 113894
rect 38422 113658 75386 113894
rect 75622 113658 112586 113894
rect 112822 113658 149786 113894
rect 150022 113658 186986 113894
rect 187222 113658 224186 113894
rect 224422 113658 261386 113894
rect 261622 113658 298586 113894
rect 298822 113658 335786 113894
rect 336022 113658 372986 113894
rect 373222 113658 410186 113894
rect 410422 113658 447386 113894
rect 447622 113658 484586 113894
rect 484822 113658 521786 113894
rect 522022 113658 558986 113894
rect 559222 113658 585802 113894
rect 586038 113658 587160 113894
rect -3236 113476 587160 113658
rect -3236 80294 587160 80476
rect -3236 80058 -3054 80294
rect -2818 80058 4586 80294
rect 4822 80058 41786 80294
rect 42022 80058 78986 80294
rect 79222 80058 116186 80294
rect 116422 80058 153386 80294
rect 153622 80058 190586 80294
rect 190822 80058 227786 80294
rect 228022 80058 264986 80294
rect 265222 80058 302186 80294
rect 302422 80058 339386 80294
rect 339622 80058 376586 80294
rect 376822 80058 413786 80294
rect 414022 80058 450986 80294
rect 451222 80058 488186 80294
rect 488422 80058 525386 80294
rect 525622 80058 562586 80294
rect 562822 80058 586742 80294
rect 586978 80058 587160 80294
rect -3236 79876 587160 80058
rect -3236 76694 587160 76876
rect -3236 76458 -2114 76694
rect -1878 76458 986 76694
rect 1222 76458 38186 76694
rect 38422 76458 75386 76694
rect 75622 76458 112586 76694
rect 112822 76458 149786 76694
rect 150022 76458 186986 76694
rect 187222 76458 224186 76694
rect 224422 76458 261386 76694
rect 261622 76458 298586 76694
rect 298822 76458 335786 76694
rect 336022 76458 372986 76694
rect 373222 76458 410186 76694
rect 410422 76458 447386 76694
rect 447622 76458 484586 76694
rect 484822 76458 521786 76694
rect 522022 76458 558986 76694
rect 559222 76458 585802 76694
rect 586038 76458 587160 76694
rect -3236 76276 587160 76458
rect -3236 43094 587160 43276
rect -3236 42858 -3054 43094
rect -2818 42858 4586 43094
rect 4822 42858 41786 43094
rect 42022 42858 78986 43094
rect 79222 42858 116186 43094
rect 116422 42858 153386 43094
rect 153622 42858 190586 43094
rect 190822 42858 227786 43094
rect 228022 42858 264986 43094
rect 265222 42858 302186 43094
rect 302422 42858 339386 43094
rect 339622 42858 376586 43094
rect 376822 42858 413786 43094
rect 414022 42858 450986 43094
rect 451222 42858 488186 43094
rect 488422 42858 525386 43094
rect 525622 42858 562586 43094
rect 562822 42858 586742 43094
rect 586978 42858 587160 43094
rect -3236 42676 587160 42858
rect -3236 39494 587160 39676
rect -3236 39258 -2114 39494
rect -1878 39258 986 39494
rect 1222 39258 38186 39494
rect 38422 39258 75386 39494
rect 75622 39258 112586 39494
rect 112822 39258 149786 39494
rect 150022 39258 186986 39494
rect 187222 39258 224186 39494
rect 224422 39258 261386 39494
rect 261622 39258 298586 39494
rect 298822 39258 335786 39494
rect 336022 39258 372986 39494
rect 373222 39258 410186 39494
rect 410422 39258 447386 39494
rect 447622 39258 484586 39494
rect 484822 39258 521786 39494
rect 522022 39258 558986 39494
rect 559222 39258 585802 39494
rect 586038 39258 587160 39494
rect -3236 39076 587160 39258
rect -3236 5894 587160 6076
rect -3236 5658 -3054 5894
rect -2818 5658 4586 5894
rect 4822 5658 41786 5894
rect 42022 5658 78986 5894
rect 79222 5658 116186 5894
rect 116422 5658 153386 5894
rect 153622 5658 190586 5894
rect 190822 5658 227786 5894
rect 228022 5658 264986 5894
rect 265222 5658 302186 5894
rect 302422 5658 339386 5894
rect 339622 5658 376586 5894
rect 376822 5658 413786 5894
rect 414022 5658 450986 5894
rect 451222 5658 488186 5894
rect 488422 5658 525386 5894
rect 525622 5658 562586 5894
rect 562822 5658 586742 5894
rect 586978 5658 587160 5894
rect -3236 5476 587160 5658
rect -3236 2294 587160 2476
rect -3236 2058 -2114 2294
rect -1878 2058 986 2294
rect 1222 2058 38186 2294
rect 38422 2058 75386 2294
rect 75622 2058 112586 2294
rect 112822 2058 149786 2294
rect 150022 2058 186986 2294
rect 187222 2058 224186 2294
rect 224422 2058 261386 2294
rect 261622 2058 298586 2294
rect 298822 2058 335786 2294
rect 336022 2058 372986 2294
rect 373222 2058 410186 2294
rect 410422 2058 447386 2294
rect 447622 2058 484586 2294
rect 484822 2058 521786 2294
rect 522022 2058 558986 2294
rect 559222 2058 585802 2294
rect 586038 2058 587160 2294
rect -3236 1876 587160 2058
rect -2296 -806 586220 -624
rect -2296 -1042 -2114 -806
rect -1878 -1042 986 -806
rect 1222 -1042 38186 -806
rect 38422 -1042 75386 -806
rect 75622 -1042 112586 -806
rect 112822 -1042 149786 -806
rect 150022 -1042 186986 -806
rect 187222 -1042 224186 -806
rect 224422 -1042 261386 -806
rect 261622 -1042 298586 -806
rect 298822 -1042 335786 -806
rect 336022 -1042 372986 -806
rect 373222 -1042 410186 -806
rect 410422 -1042 447386 -806
rect 447622 -1042 484586 -806
rect 484822 -1042 521786 -806
rect 522022 -1042 558986 -806
rect 559222 -1042 585802 -806
rect 586038 -1042 586220 -806
rect -2296 -1224 586220 -1042
rect -3236 -1746 587160 -1564
rect -3236 -1982 -3054 -1746
rect -2818 -1982 4586 -1746
rect 4822 -1982 41786 -1746
rect 42022 -1982 78986 -1746
rect 79222 -1982 116186 -1746
rect 116422 -1982 153386 -1746
rect 153622 -1982 190586 -1746
rect 190822 -1982 227786 -1746
rect 228022 -1982 264986 -1746
rect 265222 -1982 302186 -1746
rect 302422 -1982 339386 -1746
rect 339622 -1982 376586 -1746
rect 376822 -1982 413786 -1746
rect 414022 -1982 450986 -1746
rect 451222 -1982 488186 -1746
rect 488422 -1982 525386 -1746
rect 525622 -1982 562586 -1746
rect 562822 -1982 586742 -1746
rect 586978 -1982 587160 -1746
rect -3236 -2164 587160 -1982
use mux16x1_project  mprj1
timestamp 0
transform 1 0 520000 0 1 400000
box 0 552 10000 22000
use mux16x1_project  mprj2
timestamp 0
transform 1 0 520000 0 1 360000
box 0 552 10000 22000
use mux16x1_project  mprj3
timestamp 0
transform 1 0 520000 0 1 320000
box 0 552 10000 22000
use mux16x1_project  mprj4
timestamp 0
transform 1 0 520000 0 1 280000
box 0 552 10000 22000
use mux16x1_project  mprj5
timestamp 0
transform 1 0 520000 0 1 240000
box 0 552 10000 22000
use sky130_osu_ring_oscillator_mpr2aa_8_b0r1  ro1
timestamp 0
transform 1 0 292001 0 1 490002
box -1 -2 16356 1789
use sky130_osu_ring_oscillator_mpr2ca_8_b0r1  ro3
timestamp 0
transform 1 0 292005 0 1 450000
box 0 0 17146 1776
use sky130_osu_ring_oscillator_mpr2ct_8_b0r1  ro4
timestamp 0
transform 1 0 292688 0 1 430000
box -677 0 17094 1776
use sky130_osu_ring_oscillator_mpr2ea_8_b0r1  ro5
timestamp 0
transform 1 0 292655 0 1 410000
box -645 0 16230 1776
use sky130_osu_ring_oscillator_mpr2et_8_b0r1  ro6
timestamp 0
transform 1 0 293101 0 1 390000
box -1093 0 18018 1776
use sky130_osu_ring_oscillator_mpr2xa_8_b0r1  ro7
timestamp 0
transform 1 0 292560 0 1 369999
box -550 1 15260 1777
use sky130_osu_ring_oscillator_mpr2ca_8_b0r2  ro11
timestamp 0
transform 1 0 292591 0 1 290000
box -591 0 16585 1776
use sky130_osu_ring_oscillator_mpr2ct_8_b0r2  ro12
timestamp 0
transform 1 0 292686 0 1 270000
box -677 0 17094 1776
use sky130_osu_ring_oscillator_mpr2ea_8_b0r2  ro13
timestamp 0
transform 1 0 292654 0 1 250000
box -646 0 16230 1776
use sky130_osu_ring_oscillator_mpr2et_8_b0r2  ro14
timestamp 0
transform 1 0 293101 0 1 230000
box -1093 0 18018 1776
use sky130_osu_ring_oscillator_mpr2xa_8_b0r2  ro15
timestamp 0
transform 1 0 292559 0 1 209999
box -550 1 15260 1777
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal4 s -2296 -1224 -1696 705160 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -2296 -1224 586220 -624 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -2296 704560 586220 705160 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 585620 -1224 586220 705160 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 804 -2164 1404 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 38004 -2164 38604 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 75204 -2164 75804 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 112404 -2164 113004 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 149604 -2164 150204 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 186804 -2164 187404 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 224004 -2164 224604 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 261204 -2164 261804 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 298404 -2164 299004 208377 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 298404 212781 299004 368377 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 298404 372781 299004 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 335604 -2164 336204 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 372804 -2164 373404 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 410004 -2164 410604 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 447204 -2164 447804 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 484404 -2164 485004 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 521604 -2164 522204 240008 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 521604 421752 522204 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s 558804 -2164 559404 706100 0 FreeSans 3840 90 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 1876 587160 2476 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 39076 587160 39676 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 76276 587160 76876 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 113476 587160 114076 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 150676 587160 151276 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 187876 587160 188476 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 225076 587160 225676 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 262276 587160 262876 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 299476 587160 300076 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 336676 587160 337276 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 373876 587160 374476 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 411076 587160 411676 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 448276 587160 448876 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 485476 587160 486076 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 522676 587160 523276 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 559876 587160 560476 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 597076 587160 597676 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 634276 587160 634876 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal5 s -3236 671476 587160 672076 0 FreeSans 2560 0 0 0 vccd1
port 143 nsew power bidirectional
flabel metal4 s -3236 -2164 -2636 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 -2164 587160 -1564 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 705500 587160 706100 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 586560 -2164 587160 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 4404 -2164 5004 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 41604 -2164 42204 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 78804 -2164 79404 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 116004 -2164 116604 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 153204 -2164 153804 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 190404 -2164 191004 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 227604 -2164 228204 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 264804 -2164 265404 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 302004 -2164 302604 208377 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 302004 212781 302604 368377 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 302004 372781 302604 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 339204 -2164 339804 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 376404 -2164 377004 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 413604 -2164 414204 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 450804 -2164 451404 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 488004 -2164 488604 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 525204 -2164 525804 240008 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 525204 421752 525804 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal4 s 562404 -2164 563004 706100 0 FreeSans 3840 90 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 5476 587160 6076 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 42676 587160 43276 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 79876 587160 80476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 117076 587160 117676 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 154276 587160 154876 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 191476 587160 192076 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 228676 587160 229276 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 265876 587160 266476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 303076 587160 303676 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 340276 587160 340876 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 377476 587160 378076 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 414676 587160 415276 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 451876 587160 452476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 489076 587160 489676 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 526276 587160 526876 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 563476 587160 564076 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 600676 587160 601276 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 637876 587160 638476 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal5 s -3236 675076 587160 675676 0 FreeSans 2560 0 0 0 vssd1
port 144 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 145 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 146 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 147 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 148 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 149 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 150 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 151 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 152 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 153 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 154 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 155 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 156 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 157 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 158 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 159 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 160 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 161 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 162 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 163 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 164 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 165 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 166 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 167 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 168 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 169 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 170 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 171 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 172 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 173 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 174 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 175 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 176 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 177 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 178 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 179 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 180 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 181 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 182 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 183 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 184 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 185 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 186 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 187 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 188 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 189 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 190 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 191 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 192 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 193 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 194 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 195 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 196 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 197 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 198 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 199 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 200 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 201 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 202 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 203 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 204 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 205 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 206 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 207 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 208 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 209 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 210 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 211 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 212 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 213 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 214 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 215 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 216 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 217 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 218 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 219 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 220 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 221 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 222 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 223 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 224 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 225 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 226 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 227 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 228 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 229 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 230 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 231 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 232 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 233 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 234 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 235 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 236 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 237 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 238 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 239 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 240 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 241 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 242 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 243 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 244 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 245 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 246 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 247 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 248 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 249 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 250 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
