magic
tech sky130A
magscale 1 2
timestamp 1716047795
<< error_s >>
rect 1776 1756 1785 1786
rect 1804 1756 1813 1758
rect 2729 1640 2754 1647
rect 2757 1627 2782 1647
<< nwell >>
rect 1 1749 474 1750
rect 1 1120 3713 1749
rect 1 1115 616 1120
rect 1 1087 558 1115
rect 1 820 150 1087
rect 204 1035 260 1036
rect 446 850 558 1087
rect 2521 1086 2747 1120
rect 2523 744 2737 1086
rect 2759 800 2827 870
rect 3519 793 3549 828
rect 3668 744 3713 1120
<< ndiff >>
rect 3604 442 3638 476
<< locali >>
rect 1 2173 3714 2493
rect 3439 1722 3544 1758
rect 3440 1690 3441 1722
rect 3605 1461 3639 1495
rect 3286 1407 3322 1408
rect 1 1087 3713 1407
rect 2521 1086 2747 1087
rect 3284 1085 3329 1087
rect 3677 1086 3713 1087
rect 3604 998 3638 1032
rect 3440 772 3441 805
rect 3439 733 3538 772
rect 621 575 642 578
rect 621 549 660 575
rect 1081 549 1120 575
rect 1448 549 1487 572
rect 1816 549 1855 575
rect 2186 549 2226 573
rect 2521 572 2559 575
rect 2520 549 2559 572
rect 185 544 2559 549
rect 150 320 2559 544
rect 0 0 3713 320
<< viali >>
rect 3320 1879 3366 1925
rect 3604 1743 3638 1777
rect 3321 591 3367 637
rect 3604 442 3638 476
<< metal1 >>
rect 1 2173 3714 2493
rect 1751 1756 1785 2173
rect 1905 1934 1981 1943
rect 1905 1878 1914 1934
rect 1970 1878 1981 1934
rect 3320 1931 3366 1937
rect 3314 1925 3372 1931
rect 3314 1916 3320 1925
rect 3082 1909 3320 1916
rect 3094 1903 3320 1909
rect 1905 1869 1981 1878
rect 3048 1882 3320 1903
rect 3048 1869 3094 1882
rect 3314 1879 3320 1882
rect 3366 1879 3372 1925
rect 3314 1870 3372 1879
rect 3320 1867 3366 1870
rect 3127 1847 3192 1854
rect 3127 1829 3134 1847
rect 1965 1795 3134 1829
rect 3186 1795 3192 1847
rect 3127 1789 3192 1795
rect 1751 1755 1806 1756
rect 1751 1721 1841 1755
rect 2967 1709 2973 1767
rect 3025 1709 3031 1767
rect 3423 1762 3440 1794
rect 3438 1760 3440 1762
rect 1633 1694 1703 1700
rect 1633 1636 1639 1694
rect 1697 1681 1703 1694
rect 2757 1691 2825 1697
rect 2757 1681 2763 1691
rect 1697 1676 1706 1681
rect 2754 1676 2763 1681
rect 1697 1647 2763 1676
rect 1697 1640 2754 1647
rect 1697 1636 1703 1640
rect 1633 1630 1703 1636
rect 2757 1633 2763 1647
rect 2821 1681 2825 1691
rect 2821 1647 2854 1681
rect 2821 1633 2825 1647
rect 2757 1627 2825 1633
rect 2145 1405 2194 1407
rect 4 1085 3716 1405
rect 2646 953 2714 959
rect 2646 895 2652 953
rect 2710 895 2714 953
rect 2646 889 2714 895
rect 2664 698 2698 889
rect 2759 864 2827 870
rect 2759 806 2765 864
rect 2823 806 2827 864
rect 2759 800 2827 806
rect 2967 790 3031 796
rect 2967 772 2973 790
rect 2961 738 2973 772
rect 3025 738 3031 790
rect 2967 732 3031 738
rect 3122 716 3192 722
rect 3122 698 3128 716
rect 2664 664 3128 698
rect 3122 658 3128 664
rect 3186 658 3192 716
rect 3122 652 3192 658
rect 3321 645 3367 649
rect 3315 637 3373 645
rect 3315 624 3321 637
rect 3048 623 3082 624
rect 3094 623 3321 624
rect 3048 591 3321 623
rect 3367 591 3373 637
rect 3048 590 3373 591
rect 3315 583 3373 590
rect 621 575 642 576
rect 621 549 660 575
rect 1081 549 1120 575
rect 1448 549 1487 572
rect 1816 549 1855 576
rect 2521 572 2559 581
rect 3321 579 3367 583
rect 2520 549 2559 572
rect 185 544 2559 549
rect 150 521 2559 544
rect 150 465 565 521
rect 621 465 2559 521
rect 150 320 2559 465
rect 0 0 3714 320
<< via1 >>
rect 1914 1878 1970 1934
rect 3134 1795 3186 1847
rect 2973 1709 3025 1767
rect 1639 1636 1697 1694
rect 2763 1633 2821 1691
rect 2652 895 2710 953
rect 2765 806 2823 864
rect 2973 738 3025 790
rect 3128 658 3186 716
rect 565 465 621 521
<< metal2 >>
rect 1905 1934 1980 1943
rect 1905 1878 1914 1934
rect 1970 1878 1980 1934
rect 1905 1869 1980 1878
rect 3127 1847 3192 1854
rect 3127 1841 3134 1847
rect 2904 1807 3134 1841
rect 1630 1694 1706 1703
rect 1630 1636 1639 1694
rect 1697 1636 1706 1694
rect 1630 1627 1706 1636
rect 2757 1691 2825 1697
rect 2757 1633 2763 1691
rect 2821 1633 2825 1691
rect 2757 1627 2825 1633
rect 1871 1086 2698 1124
rect 1871 1036 1909 1086
rect 204 1035 260 1036
rect 1468 1035 1524 1036
rect 1860 1035 1916 1036
rect 2060 1035 2116 1036
rect 1871 1003 1909 1035
rect 2660 959 2698 1086
rect 2646 953 2714 959
rect 692 923 748 924
rect 1228 923 1284 924
rect 2646 895 2652 953
rect 2710 895 2714 953
rect 2646 889 2714 895
rect 2664 888 2698 889
rect 2774 870 2808 1627
rect 2759 864 2827 870
rect 980 810 1036 812
rect 2759 806 2765 864
rect 2823 806 2827 864
rect 2759 800 2827 806
rect 2904 772 2936 1807
rect 3127 1795 3134 1807
rect 3186 1795 3192 1847
rect 3127 1789 3192 1795
rect 2967 1709 2973 1767
rect 3025 1709 3031 1767
rect 2967 1702 3031 1709
rect 2973 1667 3007 1702
rect 2973 1632 3008 1667
rect 2973 1597 3168 1632
rect 2967 790 3031 796
rect 2967 772 2973 790
rect 564 527 598 766
rect 2904 738 2973 772
rect 3025 738 3031 790
rect 2967 732 3031 738
rect 3133 722 3168 1597
rect 3122 716 3192 722
rect 2252 699 2308 700
rect 3122 658 3128 716
rect 3186 658 3192 716
rect 3122 652 3192 658
rect 559 521 627 527
rect 559 465 565 521
rect 621 465 627 521
rect 559 459 627 465
<< via2 >>
rect 1914 1878 1970 1934
rect 1639 1636 1697 1694
<< metal3 >>
rect 1635 1703 1700 2472
rect 1905 1937 1980 1943
rect 1905 1934 2106 1937
rect 1905 1878 1914 1934
rect 1970 1878 2106 1934
rect 1905 1877 2106 1878
rect 1905 1869 1980 1877
rect 1630 1694 1706 1703
rect 1630 1636 1639 1694
rect 1697 1636 1706 1694
rect 1630 1627 1706 1636
rect 2046 1399 2106 1877
rect 79 1185 2106 1399
rect 1 1140 2106 1185
rect 1 1087 169 1140
rect 79 803 139 1087
rect 199 965 265 1032
rect 694 920 754 1140
rect 687 881 754 920
rect 687 852 751 881
rect 981 808 1041 1140
rect 1463 964 1530 1032
rect 1856 1025 1920 1032
rect 2056 1025 2120 1036
rect 1223 853 1288 920
rect 79 743 345 803
rect 975 745 1041 808
rect 975 740 1039 745
rect 2247 628 2312 700
use scs130hd_mpr2et_8  scs130hd_mpr2et_8_0
timestamp 1713287902
transform 1 0 150 0 1 559
box -48 -48 2440 592
use sky130_osu_sc_12T_hs__fill_2  sky130_osu_sc_12T_hs__fill_2_0
timestamp 1714057206
transform 1 0 2174 0 -1 2234
box -7 0 161 897
use sky130_osu_sc_12T_hs__fill_8  sky130_osu_sc_12T_hs__fill_8_0
timestamp 1714057206
transform 1 0 2345 0 -1 2234
box -9 0 179 897
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1714057206
transform 1 0 3286 0 1 260
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_2
timestamp 1714057206
transform 1 0 3483 0 1 260
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1714057206
transform 1 0 3484 0 -1 2233
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1714057206
transform 1 0 3286 0 -1 2233
box -10 0 199 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1714057206
transform 1 0 2737 0 1 259
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1714057206
transform 1 0 1614 0 -1 2234
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1714057206
transform 1 0 2737 0 -1 2234
box -10 0 552 902
<< labels >>
rlabel metal2 2793 835 2793 835 1 sel
port 9 n
rlabel metal1 78 291 78 291 1 vssd1
port 6 n
rlabel metal1 46 291 46 291 1 vssd1
port 6 n
rlabel metal1 43 2204 43 2204 1 vssd1
port 6 n
rlabel metal1 45 2202 45 2202 1 vssd1
port 6 n
rlabel metal1 1965 1795 1985 1829 1 in
port 10 n
rlabel metal1 55 1251 55 1251 1 vccd1
port 5 n
rlabel metal1 45 1251 45 1251 1 vccd1
port 5 n
rlabel viali 3604 442 3638 476 1 Y1
port 12 n
rlabel viali 3604 1743 3638 1777 1 Y0
port 11 n
<< end >>
