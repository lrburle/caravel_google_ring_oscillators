magic
tech sky130A
magscale 1 2
timestamp 1697204803
<< error_p >>
rect 1329 478 1472 480
rect 270 464 371 475
rect 557 474 821 475
rect 821 464 876 474
rect 979 468 988 477
rect 1026 468 1035 477
rect 1329 475 1451 478
rect 1301 474 1318 475
rect 1131 468 1301 474
rect 255 462 270 464
rect 249 460 255 462
rect 878 460 883 462
rect 245 455 249 460
rect 883 455 890 460
rect 970 459 979 468
rect 1035 465 1131 468
rect 1472 464 1580 478
rect 1330 456 1346 463
rect 1348 456 1364 463
rect 890 448 902 455
rect 1320 454 1332 456
rect 1342 454 1354 456
rect 1360 454 1364 456
rect 1548 454 1564 463
rect 1580 462 1598 464
rect 1599 458 1606 461
rect 1606 454 1612 458
rect 1320 449 1364 454
rect 1507 449 1544 450
rect 1612 449 1615 454
rect 1316 447 1318 449
rect 1320 447 1452 449
rect 371 446 725 447
rect 351 444 369 446
rect 811 444 824 446
rect 903 444 906 446
rect 1314 444 1452 447
rect 295 441 351 444
rect 169 433 181 441
rect 191 433 203 441
rect 267 435 351 441
rect 824 435 834 444
rect 267 434 295 435
rect 165 430 167 433
rect 267 432 286 434
rect 835 432 838 434
rect 207 429 211 430
rect 157 418 165 429
rect 168 427 203 429
rect 166 418 168 424
rect 157 417 166 418
rect 165 413 166 417
rect 164 412 165 413
rect 162 407 164 410
rect 37 405 102 406
rect 29 397 37 405
rect 102 397 106 405
rect 28 391 29 397
rect 157 395 165 407
rect 169 397 171 427
rect 200 426 203 427
rect 202 420 203 426
rect 207 422 215 429
rect 211 421 219 422
rect 243 421 244 431
rect 267 421 282 432
rect 541 422 578 424
rect 219 420 225 421
rect 242 420 243 421
rect 267 420 274 421
rect 225 410 287 420
rect 295 413 301 419
rect 341 413 347 419
rect 541 418 567 422
rect 578 418 583 422
rect 838 421 851 432
rect 814 420 828 421
rect 535 413 541 418
rect 583 413 592 418
rect 289 410 295 413
rect 296 411 353 413
rect 592 412 593 413
rect 430 411 433 412
rect 451 411 454 412
rect 533 411 534 412
rect 593 411 596 412
rect 296 410 304 411
rect 267 409 304 410
rect 169 395 203 397
rect 158 392 160 395
rect 154 379 158 391
rect 169 383 181 391
rect 194 386 203 395
rect 241 393 242 396
rect 267 392 272 409
rect 289 407 304 409
rect 347 407 353 411
rect 426 408 430 411
rect 454 408 459 411
rect 596 409 597 411
rect 788 410 814 420
rect 828 418 835 420
rect 906 418 927 444
rect 1308 437 1452 444
rect 1468 447 1569 449
rect 1468 437 1580 447
rect 1269 431 1330 437
rect 1234 428 1269 431
rect 1047 422 1234 428
rect 1320 427 1330 431
rect 835 413 850 418
rect 825 412 850 413
rect 859 412 863 413
rect 821 411 825 412
rect 835 411 872 412
rect 597 408 600 409
rect 295 405 304 407
rect 295 392 300 405
rect 348 396 367 399
rect 402 396 426 408
rect 459 400 477 408
rect 532 400 533 408
rect 204 389 214 391
rect 214 388 217 389
rect 219 386 228 388
rect 192 383 194 386
rect 228 384 239 386
rect 240 384 241 392
rect 267 384 273 392
rect 191 380 192 383
rect 239 379 273 384
rect 105 365 106 379
rect 55 356 64 365
rect 102 361 111 365
rect 102 356 116 361
rect 46 353 55 356
rect 46 352 49 353
rect 39 349 48 352
rect 27 348 48 349
rect 27 346 45 348
rect 85 346 91 352
rect 105 347 120 356
rect 145 349 154 378
rect 27 341 39 346
rect 23 339 26 341
rect 27 340 28 341
rect 33 340 39 341
rect 91 340 97 346
rect 104 345 116 347
rect 143 345 145 349
rect 183 348 191 379
rect 240 367 241 379
rect 267 376 295 379
rect 267 374 297 376
rect 267 372 298 374
rect 299 372 300 392
rect 367 387 429 396
rect 477 393 485 400
rect 531 392 532 399
rect 600 395 604 408
rect 780 407 788 410
rect 818 409 821 411
rect 814 408 818 409
rect 809 406 814 408
rect 835 406 850 411
rect 859 410 863 411
rect 872 410 873 411
rect 929 410 934 416
rect 970 412 979 421
rect 1035 419 1047 422
rect 1035 412 1044 419
rect 1314 413 1330 427
rect 1353 413 1354 437
rect 1359 432 1380 437
rect 1364 431 1380 432
rect 1497 430 1503 437
rect 1549 430 1555 437
rect 1569 431 1580 437
rect 1615 431 1624 449
rect 1364 413 1380 429
rect 1497 426 1505 430
rect 1503 424 1505 426
rect 1413 415 1441 419
rect 1443 415 1454 419
rect 863 406 868 410
rect 873 406 875 409
rect 934 406 937 410
rect 775 405 779 406
rect 850 405 853 406
rect 875 405 876 406
rect 771 403 775 405
rect 381 384 395 387
rect 417 386 418 387
rect 429 384 449 387
rect 530 384 531 391
rect 603 384 604 391
rect 652 384 658 390
rect 698 389 704 390
rect 735 389 771 403
rect 855 400 859 403
rect 870 401 874 404
rect 979 403 988 412
rect 1012 402 1015 404
rect 1026 403 1035 412
rect 1320 411 1354 413
rect 1363 412 1364 413
rect 1359 411 1364 412
rect 1409 411 1413 415
rect 1320 409 1364 411
rect 1407 410 1409 411
rect 1316 406 1317 408
rect 1090 402 1099 404
rect 1007 400 1012 402
rect 698 388 735 389
rect 698 384 704 388
rect 790 387 796 393
rect 836 387 842 393
rect 858 390 859 400
rect 1005 399 1007 400
rect 1101 399 1107 402
rect 876 396 880 399
rect 944 396 946 399
rect 880 387 890 396
rect 369 372 377 384
rect 381 382 415 384
rect 267 369 328 372
rect 267 358 273 369
rect 295 367 328 369
rect 289 366 328 367
rect 347 366 353 367
rect 289 362 353 366
rect 289 361 375 362
rect 241 355 242 358
rect 267 354 276 358
rect 295 355 301 361
rect 341 358 375 361
rect 341 355 347 358
rect 359 354 375 358
rect 381 354 383 382
rect 412 380 415 382
rect 267 350 282 354
rect 369 350 383 354
rect 413 350 415 380
rect 419 372 427 384
rect 449 375 512 384
rect 646 379 652 384
rect 664 382 700 384
rect 664 379 669 382
rect 605 378 652 379
rect 666 378 669 379
rect 704 378 710 384
rect 784 381 790 387
rect 842 381 848 387
rect 605 377 648 378
rect 529 375 530 377
rect 551 375 605 377
rect 485 363 500 375
rect 512 374 551 375
rect 529 370 530 374
rect 661 370 664 377
rect 788 374 790 375
rect 182 345 183 347
rect 242 346 243 350
rect 102 340 104 345
rect 248 344 254 350
rect 267 344 286 350
rect 294 344 300 350
rect 142 340 143 344
rect 101 338 102 340
rect 141 338 142 340
rect 15 325 23 337
rect 27 335 45 337
rect 100 336 101 337
rect 180 336 182 344
rect 242 338 248 344
rect 267 338 306 344
rect 308 338 320 346
rect 379 342 380 346
rect 381 345 398 350
rect 389 340 396 345
rect 398 344 402 345
rect 417 344 419 346
rect 485 345 500 361
rect 527 347 529 369
rect 402 341 421 344
rect 526 341 538 346
rect 548 341 560 346
rect 601 345 603 369
rect 652 345 661 369
rect 784 366 788 374
rect 697 345 700 350
rect 738 349 773 351
rect 784 349 786 366
rect 808 350 809 370
rect 856 369 858 385
rect 890 383 895 387
rect 946 383 958 396
rect 1107 392 1120 399
rect 1330 397 1346 409
rect 1348 397 1364 409
rect 1403 406 1407 409
rect 1399 402 1403 406
rect 1454 402 1467 415
rect 1503 408 1506 424
rect 1505 402 1506 408
rect 1509 408 1510 430
rect 1548 426 1555 430
rect 1576 428 1578 431
rect 1548 424 1549 426
rect 1569 425 1570 427
rect 1509 404 1511 408
rect 1542 404 1543 407
rect 1547 406 1549 424
rect 1578 420 1582 428
rect 1583 416 1584 418
rect 1584 411 1586 416
rect 1624 414 1632 431
rect 1586 406 1589 410
rect 1509 402 1513 404
rect 1547 403 1548 406
rect 1589 404 1590 406
rect 1395 399 1398 402
rect 1467 400 1470 402
rect 1393 394 1395 399
rect 1470 398 1472 400
rect 1228 393 1265 394
rect 1228 392 1253 393
rect 1265 392 1266 393
rect 1122 389 1126 392
rect 1193 389 1220 392
rect 1268 389 1275 392
rect 1320 390 1321 393
rect 1275 384 1286 389
rect 1321 386 1323 390
rect 1356 388 1357 393
rect 1391 392 1393 394
rect 1472 393 1474 398
rect 1500 396 1506 402
rect 1513 400 1519 402
rect 1520 398 1526 400
rect 1546 398 1552 402
rect 1590 401 1591 404
rect 1591 399 1592 401
rect 1526 397 1552 398
rect 1389 389 1391 392
rect 1286 383 1290 384
rect 958 380 959 383
rect 1290 379 1297 383
rect 853 358 855 361
rect 847 354 852 357
rect 844 352 847 354
rect 842 351 844 352
rect 728 347 738 349
rect 773 347 790 349
rect 717 345 728 347
rect 651 341 652 344
rect 695 341 697 345
rect 705 342 717 345
rect 784 341 786 347
rect 808 345 809 347
rect 876 345 892 361
rect 900 351 932 379
rect 960 372 966 379
rect 1297 378 1299 379
rect 1299 374 1315 378
rect 1315 373 1320 374
rect 1323 373 1331 385
rect 970 361 978 368
rect 978 359 985 361
rect 985 355 1001 359
rect 1004 355 1005 370
rect 1320 368 1336 373
rect 1357 370 1361 386
rect 1387 384 1389 389
rect 1474 385 1477 392
rect 1494 390 1500 396
rect 1526 392 1570 397
rect 1592 396 1594 399
rect 1552 390 1558 392
rect 1594 389 1597 396
rect 1386 383 1387 384
rect 1597 383 1600 389
rect 1632 384 1633 414
rect 1740 392 1756 395
rect 1668 384 1691 392
rect 1756 384 1763 392
rect 1385 381 1386 383
rect 1384 380 1385 381
rect 1600 380 1601 383
rect 1383 378 1384 379
rect 1380 374 1383 378
rect 1378 373 1380 374
rect 1601 373 1602 379
rect 1630 373 1632 383
rect 1660 379 1668 384
rect 1763 379 1770 384
rect 1650 373 1660 379
rect 1763 377 1772 379
rect 1361 368 1362 369
rect 1375 368 1378 373
rect 1499 368 1500 370
rect 1331 364 1332 367
rect 1336 365 1373 368
rect 1063 362 1094 363
rect 1054 361 1063 362
rect 1094 361 1101 362
rect 1361 361 1362 365
rect 1025 358 1054 361
rect 1101 358 1116 361
rect 1023 357 1025 358
rect 1013 355 1023 357
rect 1116 355 1133 358
rect 1333 356 1334 358
rect 1362 356 1364 361
rect 1367 356 1376 365
rect 1414 356 1423 365
rect 1498 363 1499 368
rect 1358 355 1367 356
rect 1001 352 1367 355
rect 932 350 934 351
rect 809 341 813 345
rect 863 341 876 345
rect 934 344 942 350
rect 1003 349 1013 352
rect 1143 351 1151 352
rect 1151 347 1169 351
rect 1334 347 1335 350
rect 1364 347 1365 350
rect 996 345 1001 347
rect 267 336 322 338
rect 396 336 402 340
rect 416 339 417 341
rect 15 303 23 315
rect 27 306 29 335
rect 99 334 100 335
rect 140 334 141 335
rect 267 334 324 336
rect 402 334 403 336
rect 415 335 416 338
rect 421 337 590 341
rect 649 338 651 341
rect 646 337 652 338
rect 692 337 695 341
rect 522 335 524 337
rect 526 336 527 337
rect 590 336 652 337
rect 94 330 100 334
rect 139 330 140 334
rect 179 330 180 334
rect 235 330 242 334
rect 267 333 332 334
rect 80 329 100 330
rect 80 319 94 329
rect 136 320 139 330
rect 177 319 179 330
rect 232 320 235 330
rect 64 307 80 319
rect 27 303 30 306
rect 61 303 64 307
rect 111 300 120 309
rect 132 307 136 319
rect 176 316 177 319
rect 231 316 232 319
rect 26 298 28 299
rect 33 298 39 300
rect 27 294 39 298
rect 91 294 97 300
rect 103 298 111 300
rect 130 299 132 307
rect 172 300 176 316
rect 226 300 231 316
rect 244 305 247 333
rect 294 332 320 333
rect 318 302 320 332
rect 324 322 332 333
rect 403 320 423 334
rect 471 320 485 335
rect 514 322 522 334
rect 526 332 560 334
rect 294 300 320 302
rect 324 300 332 312
rect 374 300 380 320
rect 403 300 410 320
rect 423 318 435 320
rect 469 318 471 320
rect 423 316 469 318
rect 526 300 528 332
rect 558 328 560 332
rect 559 307 560 328
rect 564 322 572 334
rect 646 332 652 336
rect 690 332 692 336
rect 704 332 710 338
rect 784 335 790 341
rect 813 337 828 341
rect 828 336 829 337
rect 842 336 876 341
rect 942 340 948 344
rect 992 342 996 345
rect 600 322 601 330
rect 644 322 647 332
rect 652 326 658 332
rect 684 322 690 332
rect 698 326 704 332
rect 787 324 788 332
rect 790 329 796 335
rect 829 334 848 336
rect 564 313 565 322
rect 594 311 600 321
rect 639 311 644 322
rect 582 307 594 311
rect 638 308 639 311
rect 677 308 684 322
rect 827 313 830 333
rect 836 329 842 334
rect 860 329 876 336
rect 948 335 959 340
rect 987 339 991 341
rect 984 338 987 339
rect 980 335 984 338
rect 1004 336 1007 341
rect 1169 338 1214 347
rect 1260 343 1273 344
rect 1239 341 1257 343
rect 1278 341 1301 343
rect 1237 340 1249 341
rect 1301 340 1310 341
rect 1310 339 1311 340
rect 1335 339 1336 347
rect 1230 338 1237 339
rect 959 328 990 335
rect 1007 332 1011 336
rect 1214 332 1237 338
rect 1311 335 1318 339
rect 1318 332 1324 335
rect 1336 332 1337 338
rect 1011 329 1084 332
rect 1214 330 1236 332
rect 936 321 990 328
rect 1001 322 1201 329
rect 1222 323 1230 330
rect 1236 328 1241 330
rect 1001 321 1035 322
rect 676 307 677 308
rect 565 306 566 307
rect 581 306 582 307
rect 560 300 581 306
rect 632 300 638 307
rect 102 296 111 298
rect 27 291 37 294
rect 39 291 45 294
rect 90 293 91 294
rect 100 293 111 296
rect 47 292 95 293
rect 98 292 100 293
rect 47 291 98 292
rect 102 291 111 293
rect 37 288 45 291
rect 37 283 41 288
rect 90 281 91 291
rect 126 286 130 299
rect 169 287 172 299
rect 222 287 226 299
rect 242 292 248 298
rect 271 297 275 300
rect 565 299 566 300
rect 122 282 126 286
rect 168 282 169 286
rect 220 283 222 287
rect 248 286 254 292
rect 120 281 122 282
rect 264 281 271 297
rect 300 292 306 298
rect 373 296 374 299
rect 402 296 403 299
rect 632 298 635 300
rect 634 297 635 298
rect 628 296 634 297
rect 294 286 300 292
rect 308 288 320 296
rect 524 294 525 296
rect 368 282 372 294
rect 398 282 401 291
rect 525 282 527 290
rect 566 283 567 290
rect 627 288 634 296
rect 621 281 634 288
rect 661 281 676 306
rect 788 300 790 313
rect 823 285 827 311
rect 936 309 968 321
rect 990 317 1035 321
rect 1068 317 1201 322
rect 1001 313 1201 317
rect 1215 316 1222 323
rect 1212 313 1215 316
rect 1241 313 1280 328
rect 1324 327 1337 332
rect 1365 328 1368 344
rect 1423 342 1432 356
rect 1494 355 1498 363
rect 1493 352 1494 355
rect 1487 344 1491 347
rect 1494 344 1500 350
rect 1552 344 1558 350
rect 1589 347 1650 373
rect 1769 372 1772 377
rect 1768 363 1772 372
rect 1661 350 1671 351
rect 1673 350 1684 351
rect 1653 347 1661 350
rect 1684 347 1706 350
rect 1768 347 1769 363
rect 1783 356 1792 365
rect 1830 356 1839 365
rect 1774 347 1783 356
rect 1839 347 1848 356
rect 1589 345 1653 347
rect 1583 344 1589 345
rect 1597 344 1598 345
rect 1628 344 1630 345
rect 1643 344 1653 345
rect 1474 342 1486 343
rect 1432 340 1436 342
rect 1454 341 1474 342
rect 1448 340 1454 341
rect 1474 336 1476 341
rect 1500 338 1506 344
rect 1534 340 1535 342
rect 1472 333 1474 336
rect 1471 332 1472 333
rect 1324 323 1339 327
rect 1337 322 1340 323
rect 1286 313 1298 319
rect 1001 312 1035 313
rect 1068 312 1308 313
rect 1337 312 1339 322
rect 1340 321 1341 322
rect 1341 316 1350 321
rect 1368 317 1370 327
rect 1459 323 1471 332
rect 1453 322 1459 323
rect 1425 321 1441 322
rect 1449 321 1453 322
rect 1518 321 1533 340
rect 1546 338 1552 344
rect 1583 342 1643 344
rect 1572 336 1643 342
rect 1706 336 1795 347
rect 1568 332 1572 336
rect 1560 327 1568 332
rect 1583 327 1643 336
rect 1397 316 1420 321
rect 1548 317 1583 327
rect 1593 321 1596 327
rect 1592 317 1593 321
rect 1628 319 1630 327
rect 1763 322 1768 330
rect 1795 327 1811 336
rect 1350 312 1356 316
rect 996 310 1000 312
rect 933 307 936 309
rect 991 307 995 309
rect 1084 308 1308 312
rect 1356 310 1362 312
rect 1387 310 1397 316
rect 1511 313 1514 317
rect 1521 316 1580 317
rect 1362 309 1363 310
rect 1100 307 1308 308
rect 918 298 933 307
rect 981 303 991 307
rect 1100 304 1316 307
rect 1213 303 1222 304
rect 1296 303 1318 304
rect 1339 303 1342 309
rect 1363 308 1367 309
rect 909 293 918 298
rect 1222 293 1240 303
rect 904 291 909 293
rect 1240 291 1244 293
rect 869 290 875 291
rect 902 290 904 291
rect 851 285 902 290
rect 915 285 921 291
rect 965 286 968 290
rect 1245 286 1253 290
rect 42 277 43 281
rect 43 274 44 277
rect 90 273 92 281
rect 108 273 120 281
rect 167 279 168 281
rect 219 279 220 281
rect 166 273 167 279
rect 218 274 219 279
rect 261 273 264 281
rect 367 278 368 281
rect 366 274 367 277
rect 395 275 397 281
rect 567 278 568 281
rect 528 273 532 278
rect 619 273 628 281
rect 657 273 665 281
rect 44 258 52 273
rect 90 266 94 273
rect 106 269 108 273
rect 165 269 166 273
rect 216 269 217 273
rect 92 258 94 266
rect 103 260 106 269
rect 163 260 165 269
rect 214 265 216 268
rect 210 261 216 265
rect 52 250 56 258
rect 94 252 95 258
rect 102 256 103 260
rect 162 256 163 260
rect 210 256 214 261
rect 256 260 261 273
rect 101 250 102 255
rect 160 250 162 255
rect 210 250 212 256
rect 253 255 256 259
rect 306 255 322 265
rect 324 255 340 265
rect 360 258 366 273
rect 249 250 253 255
rect 293 250 300 255
rect 345 249 353 255
rect 358 252 360 258
rect 388 252 395 273
rect 529 268 533 273
rect 568 268 574 273
rect 387 250 388 252
rect 402 249 418 265
rect 518 263 584 268
rect 604 265 619 273
rect 518 262 574 263
rect 509 255 518 262
rect 529 259 533 262
rect 425 249 444 250
rect 450 249 452 250
rect 57 245 58 248
rect 58 240 60 244
rect 95 240 96 244
rect 98 241 101 249
rect 158 241 160 249
rect 60 235 62 239
rect 98 235 100 241
rect 156 235 158 239
rect 63 226 66 234
rect 97 231 99 234
rect 100 231 114 235
rect 97 227 114 231
rect 66 216 71 226
rect 71 212 72 216
rect 98 215 114 227
rect 148 231 156 235
rect 194 233 210 249
rect 244 242 249 249
rect 289 242 293 249
rect 345 248 356 249
rect 386 248 402 249
rect 452 248 453 249
rect 501 248 509 255
rect 532 252 533 258
rect 568 252 574 262
rect 584 255 588 262
rect 602 260 619 265
rect 650 260 657 273
rect 659 270 665 273
rect 790 273 792 285
rect 802 281 814 285
rect 830 283 851 285
rect 821 282 830 283
rect 816 281 823 282
rect 802 277 816 281
rect 602 259 604 260
rect 602 256 603 259
rect 648 258 650 260
rect 647 257 648 258
rect 588 253 592 255
rect 601 253 602 254
rect 647 253 650 257
rect 680 253 692 256
rect 574 250 575 252
rect 529 249 531 250
rect 588 249 599 253
rect 646 249 647 253
rect 680 249 696 253
rect 698 249 714 265
rect 716 249 732 265
rect 790 261 798 273
rect 802 272 818 273
rect 802 271 812 272
rect 734 249 743 253
rect 793 251 794 255
rect 518 248 528 249
rect 345 247 357 248
rect 352 245 357 247
rect 244 233 248 242
rect 148 215 164 231
rect 194 215 210 231
rect 244 228 260 231
rect 239 222 260 228
rect 280 228 289 242
rect 352 233 356 245
rect 384 240 402 248
rect 382 235 384 239
rect 386 233 402 240
rect 425 239 437 247
rect 440 240 518 248
rect 575 240 577 248
rect 586 244 601 249
rect 646 247 651 249
rect 680 248 697 249
rect 702 248 714 249
rect 280 226 291 228
rect 300 226 312 232
rect 352 226 353 233
rect 380 229 382 233
rect 269 224 291 226
rect 301 224 312 226
rect 351 224 356 226
rect 263 222 268 224
rect 233 216 239 222
rect 244 215 260 222
rect 278 220 280 224
rect 285 222 291 224
rect 312 222 316 224
rect 291 216 297 222
rect 300 219 312 220
rect 100 212 104 215
rect 72 195 80 212
rect 104 195 111 212
rect 114 199 130 215
rect 132 199 148 215
rect 210 213 218 215
rect 236 213 244 215
rect 310 213 312 219
rect 316 213 324 220
rect 349 219 351 224
rect 352 219 356 224
rect 349 215 356 219
rect 349 213 351 215
rect 210 199 226 213
rect 228 199 244 213
rect 291 198 354 213
rect 378 201 380 227
rect 386 215 402 231
rect 413 223 421 235
rect 425 234 446 235
rect 484 234 490 240
rect 425 233 443 234
rect 402 204 406 208
rect 413 204 421 213
rect 425 204 427 233
rect 578 229 580 237
rect 586 235 608 244
rect 586 233 601 235
rect 638 233 651 247
rect 676 245 678 248
rect 682 247 696 248
rect 680 244 696 247
rect 732 246 748 249
rect 730 244 748 246
rect 638 231 646 233
rect 668 232 676 244
rect 678 242 714 244
rect 678 234 698 242
rect 711 241 714 242
rect 712 234 714 241
rect 718 240 726 244
rect 730 240 752 244
rect 732 235 752 240
rect 790 239 798 251
rect 802 241 804 271
rect 821 267 823 281
rect 863 279 869 285
rect 921 279 927 285
rect 960 282 965 286
rect 1253 282 1258 286
rect 1252 273 1260 282
rect 1264 275 1266 280
rect 1296 275 1316 303
rect 1318 297 1351 303
rect 1339 291 1342 297
rect 1351 296 1357 297
rect 1370 296 1372 309
rect 1382 308 1387 310
rect 1503 309 1511 313
rect 1521 309 1548 316
rect 1558 310 1559 315
rect 1686 314 1689 315
rect 1706 314 1710 315
rect 1680 313 1686 314
rect 1710 313 1716 314
rect 1426 297 1438 298
rect 1375 296 1397 297
rect 1357 295 1397 296
rect 1418 295 1438 297
rect 1458 295 1521 309
rect 1370 291 1372 295
rect 1426 290 1521 295
rect 1427 288 1458 290
rect 1496 288 1497 290
rect 1556 288 1558 306
rect 1590 304 1592 313
rect 1627 304 1628 313
rect 1676 312 1680 313
rect 1663 309 1676 312
rect 1717 309 1723 312
rect 1755 309 1763 322
rect 1811 313 1835 327
rect 1840 314 1841 340
rect 1835 312 1837 313
rect 1837 309 1840 312
rect 1658 308 1663 309
rect 1723 308 1726 309
rect 1589 301 1590 303
rect 1625 301 1627 303
rect 1629 301 1658 308
rect 1726 306 1739 308
rect 1754 307 1755 309
rect 1794 307 1795 309
rect 1726 301 1754 306
rect 1583 290 1629 301
rect 1738 296 1759 301
rect 1789 296 1794 306
rect 1573 288 1583 290
rect 1264 273 1316 275
rect 836 267 837 273
rect 1298 271 1316 273
rect 947 270 950 271
rect 923 268 958 270
rect 821 241 825 267
rect 919 266 923 268
rect 837 253 839 266
rect 890 249 919 266
rect 921 253 925 258
rect 931 253 947 268
rect 926 252 947 253
rect 958 265 1118 268
rect 802 239 836 241
rect 821 236 825 239
rect 580 219 583 229
rect 583 210 585 219
rect 586 215 601 231
rect 638 215 652 231
rect 675 222 676 229
rect 585 206 586 210
rect 402 203 427 204
rect 456 203 459 204
rect 402 201 459 203
rect 402 199 418 201
rect 586 200 587 204
rect 80 187 83 195
rect 111 189 116 195
rect 116 186 120 189
rect 310 186 312 198
rect 315 186 349 198
rect 354 197 356 198
rect 463 197 490 200
rect 587 198 588 200
rect 602 199 618 213
rect 620 199 636 213
rect 668 210 676 222
rect 680 215 698 234
rect 732 233 748 235
rect 732 215 748 231
rect 778 215 793 231
rect 795 216 797 233
rect 802 227 814 235
rect 824 227 836 235
rect 838 231 839 249
rect 925 246 935 252
rect 958 249 1124 265
rect 1186 249 1202 265
rect 1204 249 1220 265
rect 1264 261 1276 269
rect 1286 261 1298 269
rect 1264 251 1266 261
rect 1316 257 1320 271
rect 1342 269 1344 286
rect 1344 260 1345 269
rect 1372 260 1375 286
rect 1414 284 1460 286
rect 1555 285 1573 288
rect 1461 284 1463 285
rect 1554 284 1573 285
rect 1586 284 1587 288
rect 1414 281 1428 284
rect 1403 274 1422 281
rect 1403 273 1414 274
rect 1382 265 1403 273
rect 1378 259 1403 265
rect 1378 253 1382 259
rect 1414 252 1422 264
rect 1426 255 1428 281
rect 1497 279 1498 284
rect 1545 281 1556 284
rect 1533 277 1545 281
rect 1464 268 1465 277
rect 1498 268 1499 277
rect 1529 276 1533 277
rect 1520 273 1529 276
rect 1504 269 1520 273
rect 1501 268 1504 269
rect 1467 261 1500 268
rect 1459 255 1460 260
rect 1466 258 1500 261
rect 1554 260 1556 281
rect 1585 278 1586 284
rect 1583 268 1585 277
rect 1625 270 1627 290
rect 1675 286 1738 296
rect 1739 290 1759 296
rect 1759 288 1764 290
rect 1666 285 1675 286
rect 1660 283 1666 285
rect 1764 284 1771 288
rect 1785 286 1789 296
rect 1784 285 1785 286
rect 1771 283 1783 284
rect 1582 262 1583 267
rect 1623 261 1625 268
rect 1426 254 1430 255
rect 1457 254 1460 255
rect 1426 252 1460 254
rect 1376 249 1377 251
rect 1422 249 1423 251
rect 1459 250 1460 252
rect 1464 252 1472 258
rect 1499 257 1500 258
rect 1500 252 1501 257
rect 1553 252 1554 259
rect 1567 252 1573 258
rect 1581 257 1582 261
rect 1622 259 1623 261
rect 1630 259 1660 283
rect 1771 278 1784 283
rect 1829 279 1832 309
rect 1837 308 1841 309
rect 1840 301 1842 308
rect 1841 297 1842 301
rect 1840 291 1842 297
rect 1835 287 1840 291
rect 1841 281 1842 288
rect 1773 265 1784 278
rect 1839 277 1841 281
rect 1836 275 1839 277
rect 1579 253 1581 257
rect 1613 252 1619 258
rect 1621 257 1630 259
rect 1620 252 1630 257
rect 1464 251 1467 252
rect 1468 249 1469 251
rect 930 244 935 246
rect 1055 244 1064 249
rect 1102 244 1111 249
rect 842 243 851 244
rect 840 239 848 243
rect 851 240 866 243
rect 866 239 869 240
rect 863 233 869 239
rect 921 233 927 239
rect 935 235 944 244
rect 1046 235 1055 244
rect 1111 235 1120 244
rect 1037 233 1044 234
rect 869 231 875 233
rect 680 213 714 215
rect 727 213 732 215
rect 825 213 828 227
rect 838 215 844 231
rect 869 227 890 231
rect 915 227 921 233
rect 1031 232 1037 233
rect 1088 232 1092 234
rect 1124 233 1140 249
rect 1170 233 1186 249
rect 1197 244 1203 249
rect 1197 243 1212 244
rect 1191 237 1197 243
rect 1220 239 1236 249
rect 1243 243 1249 249
rect 1196 232 1197 234
rect 1229 232 1234 239
rect 1249 237 1255 243
rect 1267 241 1268 249
rect 1029 231 1031 232
rect 1028 228 1029 231
rect 1093 230 1095 231
rect 874 215 890 227
rect 941 219 968 222
rect 924 215 941 219
rect 968 215 976 219
rect 680 210 732 213
rect 793 210 799 213
rect 828 212 832 213
rect 680 198 684 206
rect 716 199 732 210
rect 794 203 811 210
rect 828 203 838 212
rect 794 199 810 203
rect 811 201 816 203
rect 820 201 832 203
rect 816 200 832 201
rect 812 199 832 200
rect 890 199 906 215
rect 976 213 979 215
rect 1044 213 1050 219
rect 1053 213 1055 220
rect 1095 213 1096 219
rect 1124 215 1140 231
rect 1170 215 1186 231
rect 1188 220 1197 232
rect 979 204 999 213
rect 1028 208 1029 210
rect 1038 207 1044 213
rect 1096 207 1102 213
rect 1117 204 1124 215
rect 999 200 1007 204
rect 356 192 377 197
rect 377 188 393 192
rect 425 189 437 197
rect 588 195 589 197
rect 484 188 490 194
rect 515 188 570 194
rect 589 191 590 195
rect 590 188 592 189
rect 599 188 608 197
rect 678 188 684 197
rect 736 188 742 194
rect 743 188 752 197
rect 797 192 800 199
rect 83 182 85 186
rect 120 181 128 186
rect 346 183 347 186
rect 393 182 418 188
rect 490 182 496 188
rect 536 182 542 188
rect 312 181 314 182
rect 85 178 87 181
rect 128 178 133 181
rect 302 180 312 181
rect 291 179 312 180
rect 418 179 422 182
rect 543 179 552 188
rect 590 186 599 188
rect 590 183 605 186
rect 590 179 599 183
rect 605 181 609 183
rect 684 182 696 188
rect 730 182 743 188
rect 799 185 800 192
rect 609 180 612 181
rect 133 177 135 178
rect 300 177 319 179
rect 88 174 89 177
rect 135 174 139 177
rect 89 168 92 174
rect 139 172 143 174
rect 143 170 146 172
rect 233 170 239 176
rect 291 170 297 176
rect 300 174 337 177
rect 344 174 345 177
rect 311 170 337 174
rect 340 170 344 172
rect 376 170 377 171
rect 146 167 150 170
rect 92 161 96 167
rect 150 161 160 167
rect 163 161 175 165
rect 239 164 245 170
rect 285 164 291 170
rect 337 167 377 170
rect 337 164 376 167
rect 422 166 439 179
rect 543 178 544 179
rect 612 177 619 180
rect 687 179 696 182
rect 734 179 743 182
rect 793 180 800 185
rect 828 183 832 199
rect 870 188 879 197
rect 935 188 944 197
rect 1007 195 1018 200
rect 1111 199 1124 204
rect 1186 210 1195 215
rect 1196 210 1197 220
rect 1186 204 1197 210
rect 1200 204 1202 232
rect 1268 231 1270 232
rect 1266 226 1270 231
rect 1319 231 1320 249
rect 1362 234 1378 249
rect 1454 248 1459 249
rect 1426 240 1438 248
rect 1448 240 1460 248
rect 1362 233 1380 234
rect 1378 231 1380 233
rect 1186 199 1202 204
rect 1251 214 1312 226
rect 1319 220 1332 231
rect 1318 215 1332 220
rect 1362 218 1380 231
rect 1447 228 1454 240
rect 1470 237 1471 240
rect 1501 237 1502 246
rect 1552 240 1553 249
rect 1561 246 1567 252
rect 1619 249 1625 252
rect 1674 249 1690 265
rect 1770 261 1784 265
rect 1832 261 1834 275
rect 1835 261 1841 267
rect 1770 259 1789 261
rect 1770 252 1773 259
rect 1783 255 1789 259
rect 1829 255 1835 261
rect 1770 249 1771 252
rect 1834 251 1835 255
rect 1617 246 1625 249
rect 1617 245 1619 246
rect 1620 241 1621 243
rect 1621 238 1623 241
rect 1471 230 1472 234
rect 1502 230 1503 236
rect 1440 222 1447 228
rect 1439 221 1440 222
rect 1362 215 1378 218
rect 1412 215 1439 221
rect 1251 200 1316 214
rect 1282 199 1298 200
rect 1300 199 1316 200
rect 1343 199 1344 201
rect 1378 199 1394 215
rect 1472 208 1476 226
rect 1503 220 1504 229
rect 1552 228 1554 235
rect 1617 231 1618 235
rect 1623 232 1626 238
rect 1658 233 1674 249
rect 1708 243 1736 249
rect 1702 235 1736 243
rect 1698 232 1700 235
rect 1708 231 1736 235
rect 1754 233 1770 249
rect 1831 240 1835 249
rect 1829 235 1831 240
rect 1554 222 1555 228
rect 1617 223 1634 231
rect 1504 207 1509 220
rect 1556 215 1564 221
rect 1618 217 1634 223
rect 1690 220 1698 231
rect 1687 219 1698 220
rect 1702 229 1736 231
rect 1618 215 1628 217
rect 1564 214 1566 215
rect 1476 201 1477 207
rect 1509 200 1511 207
rect 1566 206 1580 214
rect 1618 207 1619 215
rect 1634 209 1639 217
rect 1687 211 1696 219
rect 1615 206 1619 207
rect 1561 205 1594 206
rect 1615 205 1625 206
rect 1561 200 1567 205
rect 1111 197 1117 199
rect 1188 198 1202 199
rect 1314 198 1317 199
rect 1196 197 1249 198
rect 1029 195 1030 197
rect 1111 195 1120 197
rect 793 179 799 180
rect 839 179 845 185
rect 879 179 888 188
rect 926 179 935 188
rect 1018 187 1032 195
rect 1106 188 1120 195
rect 1191 191 1255 197
rect 1318 191 1333 197
rect 1340 195 1341 197
rect 1336 191 1340 194
rect 1382 193 1383 194
rect 1106 187 1111 188
rect 1032 186 1035 187
rect 545 175 546 177
rect 547 168 550 174
rect 619 172 634 177
rect 787 173 793 179
rect 845 174 851 179
rect 899 175 911 179
rect 952 175 968 185
rect 1030 183 1031 186
rect 1035 183 1074 186
rect 1104 184 1111 187
rect 1197 186 1212 191
rect 1243 188 1252 191
rect 1197 185 1203 186
rect 1243 185 1249 188
rect 1031 180 1074 183
rect 1035 178 1074 180
rect 1097 180 1104 184
rect 1106 180 1111 184
rect 1252 180 1275 188
rect 1333 186 1346 191
rect 1382 188 1390 193
rect 1478 192 1479 197
rect 1512 191 1515 197
rect 1567 194 1573 200
rect 1578 199 1594 205
rect 1596 199 1612 205
rect 1619 200 1625 205
rect 1639 203 1642 209
rect 1678 202 1687 211
rect 1613 194 1619 200
rect 1644 197 1646 201
rect 1332 183 1334 186
rect 1346 182 1354 186
rect 1383 185 1390 188
rect 1479 187 1480 191
rect 1392 183 1393 185
rect 1480 182 1481 185
rect 1515 182 1518 191
rect 1601 186 1604 188
rect 1646 184 1654 197
rect 1674 195 1678 199
rect 1690 197 1698 209
rect 1702 199 1704 229
rect 1733 228 1736 229
rect 1740 220 1783 232
rect 1734 217 1783 220
rect 1804 217 1829 235
rect 1734 211 1743 217
rect 1754 215 1770 217
rect 1783 215 1829 217
rect 1743 205 1752 211
rect 1746 204 1752 205
rect 1770 209 1804 215
rect 1747 200 1750 204
rect 1770 199 1786 209
rect 1804 203 1821 209
rect 1807 199 1813 203
rect 1821 201 1827 203
rect 1827 199 1831 201
rect 1853 199 1859 205
rect 1702 198 1717 199
rect 1702 197 1721 198
rect 1678 191 1683 195
rect 1718 193 1736 197
rect 1753 194 1759 197
rect 1801 194 1807 199
rect 1702 191 1736 193
rect 1759 192 1807 194
rect 1859 193 1865 199
rect 1683 190 1719 191
rect 1702 185 1714 190
rect 1769 185 1780 190
rect 1780 184 1782 185
rect 1654 182 1655 184
rect 1097 179 1111 180
rect 1084 178 1097 179
rect 1104 176 1106 179
rect 1275 176 1286 180
rect 1329 178 1330 180
rect 895 174 977 175
rect 845 173 911 174
rect 888 172 911 173
rect 634 167 646 172
rect 888 170 895 172
rect 899 171 911 172
rect 977 170 980 173
rect 1096 172 1103 175
rect 1286 172 1298 176
rect 1326 174 1328 177
rect 1298 170 1305 172
rect 1321 170 1325 172
rect 884 169 888 170
rect 877 167 884 169
rect 914 168 915 170
rect 980 169 982 170
rect 336 162 407 164
rect 160 160 175 161
rect 337 160 407 162
rect 439 160 443 166
rect 550 164 552 167
rect 163 157 175 160
rect 99 153 104 157
rect 176 155 179 157
rect 328 153 336 160
rect 338 158 348 160
rect 338 153 342 158
rect 104 137 125 153
rect 169 151 193 153
rect 173 146 193 151
rect 328 148 338 153
rect 335 146 338 148
rect 125 136 127 137
rect 131 130 132 133
rect 129 119 136 128
rect 173 121 175 146
rect 179 141 187 146
rect 193 140 199 146
rect 332 142 335 146
rect 199 135 205 140
rect 327 137 335 142
rect 327 136 333 137
rect 205 133 208 135
rect 141 119 175 121
rect 179 119 187 131
rect 208 129 209 133
rect 321 130 327 136
rect 331 133 332 135
rect 330 129 331 132
rect 340 130 342 153
rect 372 156 427 160
rect 372 142 395 156
rect 403 154 427 156
rect 447 154 448 156
rect 408 149 427 154
rect 448 149 452 154
rect 552 151 559 164
rect 646 163 676 167
rect 895 165 911 167
rect 646 155 688 163
rect 415 142 427 149
rect 452 142 458 149
rect 559 146 562 151
rect 640 150 689 151
rect 372 136 379 142
rect 372 134 385 136
rect 372 130 374 134
rect 379 130 385 134
rect 390 132 399 141
rect 418 137 427 142
rect 458 137 461 142
rect 329 126 330 128
rect 373 126 374 130
rect 392 127 408 132
rect 421 130 427 137
rect 461 130 467 137
rect 562 136 599 146
rect 640 143 654 150
rect 670 149 689 150
rect 686 144 689 149
rect 639 140 640 142
rect 599 134 605 136
rect 637 135 639 140
rect 605 133 610 134
rect 636 133 637 135
rect 426 128 427 130
rect 467 127 469 130
rect 610 129 626 133
rect 626 128 628 129
rect 209 121 211 126
rect 328 121 329 126
rect 394 123 397 127
rect 399 123 408 127
rect 400 121 401 123
rect 136 117 137 119
rect 140 117 141 119
rect 327 117 328 119
rect 401 118 402 121
rect 136 101 140 117
rect 176 115 179 117
rect 141 107 153 115
rect 163 107 175 115
rect 211 101 215 117
rect 400 103 402 116
rect 429 113 441 126
rect 469 113 481 127
rect 631 126 637 128
rect 637 124 645 126
rect 642 122 646 124
rect 642 117 649 122
rect 686 119 688 144
rect 689 138 690 143
rect 692 139 700 151
rect 845 135 873 136
rect 909 135 911 165
rect 915 155 923 167
rect 982 153 984 169
rect 1305 168 1311 170
rect 1318 168 1321 170
rect 1038 161 1044 167
rect 1096 161 1102 167
rect 1302 164 1322 168
rect 1354 164 1375 182
rect 1380 179 1391 181
rect 1302 162 1318 164
rect 1297 161 1302 162
rect 1322 161 1330 164
rect 1044 155 1050 161
rect 1090 155 1096 161
rect 1290 158 1297 161
rect 1330 160 1333 161
rect 1375 160 1380 164
rect 1285 157 1290 158
rect 1333 157 1339 160
rect 1380 157 1384 160
rect 1388 157 1390 179
rect 1391 178 1392 179
rect 1394 178 1402 181
rect 1392 175 1402 178
rect 1394 170 1402 175
rect 1481 174 1482 182
rect 1518 178 1521 182
rect 1482 170 1483 174
rect 1511 170 1523 178
rect 1533 170 1545 178
rect 1608 170 1621 182
rect 1394 169 1403 170
rect 1399 167 1403 169
rect 1394 157 1402 159
rect 1403 157 1426 167
rect 1483 165 1490 170
rect 1507 168 1510 170
rect 1523 166 1524 170
rect 1530 166 1536 170
rect 1484 164 1490 165
rect 1499 164 1507 166
rect 1511 164 1557 166
rect 1478 158 1484 164
rect 1511 158 1513 164
rect 1536 158 1542 164
rect 1543 158 1557 164
rect 1276 154 1285 157
rect 1271 152 1276 154
rect 690 134 691 135
rect 865 133 873 135
rect 877 133 911 135
rect 915 133 923 145
rect 982 135 984 151
rect 1255 147 1271 152
rect 1239 142 1255 147
rect 1339 146 1357 157
rect 1384 148 1428 157
rect 1482 154 1484 155
rect 1480 150 1482 154
rect 1366 147 1428 148
rect 1384 146 1428 147
rect 1339 143 1358 146
rect 1332 142 1366 143
rect 1384 142 1453 146
rect 1543 143 1545 158
rect 1549 154 1564 158
rect 1552 146 1564 154
rect 1621 153 1640 170
rect 1655 156 1689 182
rect 1784 164 1807 182
rect 1643 147 1653 150
rect 1654 147 1666 156
rect 1689 155 1691 156
rect 1691 150 1731 155
rect 1753 150 1765 155
rect 1731 148 1765 150
rect 1731 147 1779 148
rect 1801 147 1807 153
rect 1859 147 1865 153
rect 1228 139 1239 142
rect 1322 139 1330 142
rect 1339 141 1358 142
rect 691 129 692 133
rect 654 117 688 119
rect 692 117 700 129
rect 787 127 793 133
rect 845 127 851 133
rect 877 129 884 133
rect 993 132 999 138
rect 1039 132 1045 138
rect 1085 132 1228 139
rect 1300 132 1322 139
rect 1356 133 1358 141
rect 1359 134 1365 139
rect 1378 135 1453 142
rect 980 129 982 132
rect 877 128 889 129
rect 793 121 799 127
rect 839 121 845 127
rect 877 126 892 128
rect 899 126 911 129
rect 979 128 980 129
rect 978 126 979 128
rect 987 126 993 132
rect 1045 126 1051 132
rect 1052 130 1073 132
rect 1295 130 1300 132
rect 1289 128 1295 130
rect 1358 129 1359 133
rect 1367 130 1370 132
rect 1056 126 1091 128
rect 877 121 889 126
rect 892 121 914 126
rect 976 124 978 126
rect 914 117 927 121
rect 927 116 932 117
rect 941 116 991 124
rect 1044 123 1056 126
rect 1035 121 1044 123
rect 1096 121 1098 126
rect 1279 125 1287 128
rect 1359 127 1360 128
rect 1272 123 1279 125
rect 1034 117 1035 121
rect 1265 120 1272 123
rect 1360 121 1362 123
rect 1260 119 1265 120
rect 1254 117 1260 119
rect 690 113 692 116
rect 932 115 991 116
rect 941 113 991 115
rect 135 95 136 99
rect 215 98 216 101
rect 397 97 400 103
rect 135 71 137 95
rect 215 71 216 95
rect 327 90 330 97
rect 321 88 330 90
rect 321 84 327 88
rect 330 84 354 88
rect 379 84 385 90
rect 395 89 397 97
rect 327 78 354 84
rect 373 78 379 84
rect 389 83 395 88
rect 399 83 408 85
rect 441 84 466 113
rect 481 107 488 113
rect 654 107 666 113
rect 676 107 688 113
rect 918 107 941 113
rect 488 105 694 107
rect 907 105 918 107
rect 635 83 636 101
rect 137 67 140 71
rect 330 67 354 78
rect 389 76 408 83
rect 467 80 471 83
rect 471 77 476 80
rect 389 71 404 76
rect 476 72 520 77
rect 388 67 404 71
rect 520 69 540 72
rect 634 71 636 83
rect 694 95 853 105
rect 865 95 907 105
rect 1031 102 1034 115
rect 1098 102 1101 117
rect 1249 115 1254 117
rect 1246 114 1249 115
rect 1241 113 1246 114
rect 1235 111 1241 113
rect 1362 111 1367 121
rect 1376 119 1383 125
rect 1384 123 1453 135
rect 1480 133 1481 139
rect 1544 133 1545 142
rect 1549 134 1557 144
rect 1564 143 1568 146
rect 1629 143 1654 147
rect 1751 145 1764 147
rect 1552 132 1557 134
rect 1568 133 1579 143
rect 1384 119 1428 123
rect 1383 112 1391 119
rect 1428 112 1436 119
rect 1453 117 1459 123
rect 1482 120 1483 123
rect 1484 118 1499 128
rect 1459 114 1463 117
rect 1216 109 1235 111
rect 1179 105 1216 109
rect 1102 101 1179 105
rect 1367 101 1380 111
rect 1391 101 1421 112
rect 1436 104 1446 112
rect 1463 104 1467 114
rect 1478 112 1499 118
rect 1525 123 1536 128
rect 1525 122 1549 123
rect 1525 120 1545 122
rect 1579 120 1584 133
rect 1629 129 1678 143
rect 1703 139 1749 145
rect 1767 144 1769 147
rect 1779 145 1799 147
rect 1807 145 1826 147
rect 1750 141 1765 143
rect 1695 135 1703 139
rect 1629 128 1674 129
rect 1525 118 1536 120
rect 1611 119 1629 128
rect 1650 124 1674 128
rect 1678 128 1684 129
rect 1686 128 1695 135
rect 1678 127 1686 128
rect 1684 126 1688 127
rect 1650 118 1681 124
rect 1688 123 1696 126
rect 1696 121 1706 123
rect 1707 119 1710 120
rect 1525 112 1542 118
rect 1583 112 1584 117
rect 1594 112 1609 118
rect 1484 106 1490 112
rect 1530 106 1536 112
rect 1574 104 1594 112
rect 1650 110 1674 118
rect 1713 117 1718 119
rect 694 93 865 95
rect 694 83 696 93
rect 987 85 993 86
rect 965 83 993 85
rect 694 75 700 83
rect 959 80 976 83
rect 987 80 993 83
rect 941 77 959 80
rect 695 71 700 75
rect 922 74 941 77
rect 993 74 999 80
rect 1025 77 1031 101
rect 1095 96 1096 98
rect 1101 96 1179 101
rect 1062 94 1096 96
rect 1100 94 1108 96
rect 1100 92 1105 94
rect 1052 89 1061 90
rect 1045 80 1051 86
rect 1084 82 1096 90
rect 1101 84 1105 92
rect 1039 74 1045 80
rect 1103 77 1105 84
rect 1380 83 1426 101
rect 1446 88 1490 104
rect 1510 88 1511 101
rect 1535 88 1574 104
rect 1583 101 1584 104
rect 1456 87 1527 88
rect 1535 87 1564 88
rect 1456 84 1564 87
rect 1462 83 1467 84
rect 1380 82 1428 83
rect 907 72 922 74
rect 711 71 751 72
rect 905 71 907 72
rect 550 69 711 71
rect 751 69 780 71
rect 634 67 637 69
rect 693 67 700 69
rect 140 59 148 67
rect 208 59 215 66
rect 148 58 208 59
rect 372 51 388 67
rect 637 56 643 67
rect 690 59 693 66
rect 780 63 841 69
rect 851 63 901 71
rect 1101 68 1103 77
rect 682 56 690 59
rect 643 54 684 56
rect 1025 54 1038 65
rect 1079 57 1101 68
rect 1380 67 1426 82
rect 1430 78 1433 80
rect 1433 77 1435 78
rect 1435 74 1442 77
rect 1462 75 1476 83
rect 1510 75 1511 84
rect 1582 78 1583 94
rect 1609 87 1674 110
rect 1719 115 1725 117
rect 1719 109 1727 115
rect 1731 111 1733 113
rect 1763 111 1765 141
rect 1769 131 1777 143
rect 1807 141 1813 145
rect 1853 141 1859 147
rect 1877 134 1888 143
rect 1731 109 1765 111
rect 1769 109 1777 121
rect 1888 119 1891 133
rect 1891 117 1892 119
rect 1727 105 1730 107
rect 1731 97 1743 105
rect 1753 97 1765 105
rect 1892 102 1895 117
rect 1731 89 1740 97
rect 1894 89 1895 102
rect 1595 82 1607 87
rect 1586 78 1595 82
rect 1442 72 1448 74
rect 1460 71 1476 75
rect 1451 67 1476 71
rect 1510 67 1512 71
rect 1444 63 1469 67
rect 1039 54 1079 57
rect 650 51 666 54
rect 668 51 684 54
rect 1444 51 1460 63
rect 1469 60 1477 63
rect 1477 59 1486 60
rect 1512 56 1517 67
rect 1544 61 1586 78
rect 1650 70 1674 87
rect 1541 60 1544 61
rect 1535 59 1541 60
rect 1573 59 1580 61
rect 1569 56 1573 59
rect 1517 52 1538 56
rect 1560 52 1569 56
rect 1710 47 1734 70
rect 1740 67 1779 89
rect 1779 62 1788 67
rect 1885 63 1894 84
rect 1884 62 1885 63
rect 1788 56 1805 62
rect 1880 57 1884 62
rect 1877 56 1880 57
rect 1805 52 1877 56
rect 66 -2 116 47
rect 146 -2 212 47
rect 242 -2 308 47
rect 338 -2 404 47
rect 434 -2 484 47
rect 554 -2 604 47
rect 634 -2 700 47
rect 730 -2 796 47
rect 826 -2 892 47
rect 922 -2 972 47
rect 1042 -2 1092 47
rect 1122 -2 1188 47
rect 1218 -2 1284 47
rect 1314 -2 1380 47
rect 1410 -2 1460 47
rect 1530 -2 1580 47
rect 1610 -2 1676 47
rect 1706 -2 1772 47
rect 1802 -2 1852 47
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 51 38 1868 183
rect 33 -17 67 17
rect 521 -17 555 17
rect 1009 -17 1043 17
rect 1497 -17 1531 17
<< nmos >>
rect 116 48 146 177
rect 212 48 242 177
rect 308 48 338 177
rect 404 48 434 177
rect 604 48 634 177
rect 700 48 730 177
rect 796 48 826 177
rect 892 48 922 177
rect 1092 48 1122 177
rect 1188 48 1218 177
rect 1284 48 1314 177
rect 1380 48 1410 177
rect 1580 48 1610 177
rect 1676 48 1706 177
rect 1772 48 1802 177
<< scnmos >>
rect 116 47 146 48
rect 212 47 242 48
rect 308 47 338 48
rect 404 47 434 48
rect 604 47 634 48
rect 700 47 730 48
rect 796 47 826 48
rect 892 47 922 48
rect 1092 47 1122 48
rect 1188 47 1218 48
rect 1284 47 1314 48
rect 1380 47 1410 48
rect 1580 47 1610 48
rect 1676 47 1706 48
rect 1772 47 1802 48
<< pmos >>
rect 116 297 146 497
rect 212 297 242 497
rect 308 297 338 497
rect 404 297 434 497
rect 604 297 634 497
rect 700 297 730 497
rect 796 297 826 497
rect 892 297 922 497
rect 1092 297 1122 497
rect 1188 297 1218 497
rect 1284 297 1314 497
rect 1380 297 1410 497
rect 1580 297 1610 497
rect 1676 297 1706 497
rect 1772 297 1802 497
<< ndiff >>
rect 58 101 116 177
rect 58 67 66 101
rect 100 67 116 101
rect 58 47 116 67
rect 146 101 212 177
rect 146 67 162 101
rect 196 67 212 101
rect 146 47 212 67
rect 242 101 308 177
rect 242 67 258 101
rect 292 67 308 101
rect 242 47 308 67
rect 338 101 404 177
rect 338 67 354 101
rect 388 67 404 101
rect 338 47 404 67
rect 434 101 492 177
rect 434 67 450 101
rect 484 67 492 101
rect 434 47 492 67
rect 546 101 604 177
rect 546 67 554 101
rect 588 67 604 101
rect 546 47 604 67
rect 634 101 700 177
rect 634 67 650 101
rect 684 67 700 101
rect 634 47 700 67
rect 730 101 796 177
rect 730 67 746 101
rect 780 67 796 101
rect 730 47 796 67
rect 826 47 892 177
rect 922 169 980 177
rect 922 135 934 169
rect 968 135 980 169
rect 922 47 980 135
rect 1034 101 1092 177
rect 1034 67 1042 101
rect 1076 67 1092 101
rect 1034 47 1092 67
rect 1122 47 1188 177
rect 1218 101 1284 177
rect 1218 67 1234 101
rect 1268 67 1284 101
rect 1218 47 1284 67
rect 1314 47 1380 177
rect 1410 101 1468 177
rect 1410 67 1426 101
rect 1460 67 1468 101
rect 1410 47 1468 67
rect 1522 101 1580 177
rect 1522 67 1530 101
rect 1564 67 1580 101
rect 1522 47 1580 67
rect 1610 101 1676 177
rect 1610 67 1626 101
rect 1660 67 1676 101
rect 1610 47 1676 67
rect 1706 47 1772 177
rect 1802 101 1860 177
rect 1802 67 1818 101
rect 1852 67 1860 101
rect 1802 47 1860 67
<< pdiff >>
rect 58 379 116 497
rect 58 345 66 379
rect 100 345 116 379
rect 58 297 116 345
rect 146 297 212 497
rect 242 477 308 497
rect 242 443 258 477
rect 292 443 308 477
rect 242 297 308 443
rect 338 297 404 497
rect 434 379 492 497
rect 434 345 450 379
rect 484 345 492 379
rect 434 297 492 345
rect 546 379 604 497
rect 546 345 554 379
rect 588 345 604 379
rect 546 297 604 345
rect 634 297 700 497
rect 730 477 796 497
rect 730 443 746 477
rect 780 443 796 477
rect 730 297 796 443
rect 826 379 892 497
rect 826 345 842 379
rect 876 345 892 379
rect 826 297 892 345
rect 922 477 980 497
rect 922 443 938 477
rect 972 443 980 477
rect 922 297 980 443
rect 1034 379 1092 497
rect 1034 345 1042 379
rect 1076 345 1092 379
rect 1034 297 1092 345
rect 1122 477 1188 497
rect 1122 443 1138 477
rect 1172 443 1188 477
rect 1122 297 1188 443
rect 1218 379 1284 497
rect 1218 345 1234 379
rect 1268 345 1284 379
rect 1218 297 1284 345
rect 1314 447 1380 497
rect 1314 413 1330 447
rect 1364 413 1380 447
rect 1314 297 1380 413
rect 1410 379 1468 497
rect 1410 345 1426 379
rect 1460 345 1468 379
rect 1410 297 1468 345
rect 1522 447 1580 497
rect 1522 413 1530 447
rect 1564 413 1580 447
rect 1522 297 1580 413
rect 1610 477 1676 497
rect 1610 443 1626 477
rect 1660 443 1676 477
rect 1610 297 1676 443
rect 1706 379 1772 497
rect 1706 345 1722 379
rect 1756 345 1772 379
rect 1706 297 1772 345
rect 1802 477 1860 497
rect 1802 443 1818 477
rect 1852 443 1860 477
rect 1802 297 1860 443
<< ndiffc >>
rect 66 67 100 101
rect 162 67 196 101
rect 258 67 292 101
rect 354 67 388 101
rect 450 67 484 101
rect 554 67 588 101
rect 650 67 684 101
rect 746 67 780 101
rect 934 135 968 169
rect 1042 67 1076 101
rect 1234 67 1268 101
rect 1426 67 1460 101
rect 1530 67 1564 101
rect 1626 67 1660 101
rect 1818 67 1852 101
<< pdiffc >>
rect 66 345 100 379
rect 258 443 292 477
rect 450 345 484 379
rect 554 345 588 379
rect 746 443 780 477
rect 842 345 876 379
rect 938 443 972 477
rect 1042 345 1076 379
rect 1138 443 1172 477
rect 1234 345 1268 379
rect 1330 413 1364 447
rect 1426 345 1460 379
rect 1530 413 1564 447
rect 1626 443 1660 477
rect 1722 345 1756 379
rect 1818 443 1852 477
<< poly >>
rect 116 497 146 523
rect 212 497 242 523
rect 308 497 338 523
rect 404 497 434 523
rect 604 497 634 523
rect 700 497 730 523
rect 796 497 826 523
rect 892 497 922 523
rect 1092 497 1122 523
rect 1188 497 1218 523
rect 1284 497 1314 523
rect 1380 497 1410 523
rect 1580 497 1610 523
rect 1676 497 1706 523
rect 1772 497 1802 523
rect 116 265 146 297
rect 212 265 242 297
rect 308 265 338 297
rect 404 265 434 297
rect 604 265 634 297
rect 700 265 730 297
rect 796 265 826 297
rect 892 265 922 297
rect 1092 265 1122 297
rect 1188 265 1218 297
rect 1284 265 1314 297
rect 1380 265 1410 297
rect 1580 265 1610 297
rect 1676 265 1706 297
rect 1772 265 1802 297
rect 104 249 158 265
rect 104 215 114 249
rect 148 215 158 249
rect 104 199 158 215
rect 200 249 254 265
rect 200 215 210 249
rect 244 215 254 249
rect 200 199 254 215
rect 296 249 350 265
rect 296 215 306 249
rect 340 215 350 249
rect 296 199 350 215
rect 392 249 446 265
rect 392 215 402 249
rect 436 215 446 249
rect 392 199 446 215
rect 592 249 646 265
rect 592 215 602 249
rect 636 215 646 249
rect 592 199 646 215
rect 688 249 742 265
rect 688 215 698 249
rect 732 215 742 249
rect 688 199 742 215
rect 784 249 838 265
rect 784 215 794 249
rect 828 215 838 249
rect 784 199 838 215
rect 880 249 934 265
rect 880 215 890 249
rect 924 215 934 249
rect 880 199 934 215
rect 1080 249 1134 265
rect 1080 215 1090 249
rect 1124 215 1134 249
rect 1080 199 1134 215
rect 1176 249 1230 265
rect 1176 215 1186 249
rect 1220 215 1230 249
rect 1176 199 1230 215
rect 1272 249 1326 265
rect 1272 215 1282 249
rect 1316 215 1326 249
rect 1272 199 1326 215
rect 1368 249 1422 265
rect 1368 215 1378 249
rect 1412 215 1422 249
rect 1368 199 1422 215
rect 1568 249 1622 265
rect 1568 215 1578 249
rect 1612 215 1622 249
rect 1568 199 1622 215
rect 1664 249 1718 265
rect 1664 215 1674 249
rect 1708 215 1718 249
rect 1664 199 1718 215
rect 1760 249 1814 265
rect 1760 215 1770 249
rect 1804 215 1814 249
rect 1760 199 1814 215
rect 116 177 146 199
rect 212 177 242 199
rect 308 177 338 199
rect 404 177 434 199
rect 604 177 634 199
rect 700 177 730 199
rect 796 177 826 199
rect 892 177 922 199
rect 1092 177 1122 199
rect 1188 177 1218 199
rect 1284 177 1314 199
rect 1380 177 1410 199
rect 1580 177 1610 199
rect 1676 177 1706 199
rect 1772 177 1802 199
rect 116 21 146 47
rect 212 21 242 47
rect 308 21 338 47
rect 404 21 434 47
rect 604 21 634 47
rect 700 21 730 47
rect 796 21 826 47
rect 892 21 922 47
rect 1092 21 1122 47
rect 1188 21 1218 47
rect 1284 21 1314 47
rect 1380 21 1410 47
rect 1580 21 1610 47
rect 1676 21 1706 47
rect 1772 21 1802 47
<< polycont >>
rect 114 215 148 249
rect 210 215 244 249
rect 306 215 340 249
rect 402 215 436 249
rect 602 215 636 249
rect 698 215 732 249
rect 794 215 828 249
rect 890 215 924 249
rect 1090 215 1124 249
rect 1186 215 1220 249
rect 1282 215 1316 249
rect 1378 215 1412 249
rect 1578 215 1612 249
rect 1674 215 1708 249
rect 1770 215 1804 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 258 477 292 527
tri 168 427 169 429 se
tri 166 418 168 424 se
rect 168 418 169 427
tri 165 413 166 418 se
rect 166 413 169 418
tri 164 412 165 413 se
rect 165 412 169 413
tri 162 406 164 410 se
rect 164 406 169 412
tri 37 405 102 406 se
tri 29 397 37 405 se
rect 37 397 102 405
tri 102 397 106 405 sw
tri 160 397 162 405 se
rect 162 397 169 406
tri 28 391 29 397 se
rect 29 391 106 397
tri 158 392 160 397 se
rect 160 395 169 397
rect 258 427 292 443
rect 746 477 780 527
rect 746 427 780 443
rect 938 477 972 527
rect 938 427 972 443
rect 1138 477 1172 527
rect 1626 477 1660 527
rect 1138 427 1172 443
tri 1320 454 1322 456 se
rect 1322 454 1360 456
tri 1360 454 1361 456 sw
rect 1320 447 1361 454
tri 1361 447 1364 453 sw
rect 1320 444 1330 447
tri 541 418 567 424 se
tri 567 422 578 424 sw
rect 567 418 578 422
tri 578 418 583 422 sw
tri 535 413 541 418 se
rect 541 413 583 418
tri 583 413 592 418 sw
rect 1509 447 1569 454
rect 1509 438 1530 447
tri 1413 415 1441 419 se
rect 1441 415 1443 419
tri 1443 415 1454 419 sw
rect 535 412 592 413
tri 592 412 593 413 sw
tri 825 412 836 413 se
tri 836 412 848 413 sw
tri 430 411 433 412 se
rect 433 411 451 412
tri 451 411 454 412 sw
tri 533 411 534 412 se
rect 534 411 593 412
tri 593 411 596 412 sw
tri 821 411 825 412 se
rect 825 411 848 412
tri 848 411 872 412 sw
tri 426 408 430 411 se
rect 430 408 454 411
tri 454 408 459 411 sw
rect 533 409 596 411
tri 596 409 597 411 sw
tri 818 409 821 411 se
rect 821 410 872 411
tri 872 410 873 411 sw
rect 821 409 873 410
rect 1354 412 1363 413
tri 1363 412 1364 413 nw
rect 1354 411 1359 412
tri 1359 411 1363 412 nw
tri 1409 411 1413 415 se
rect 1413 411 1454 415
tri 1354 410 1359 411 nw
tri 1407 410 1409 411 se
rect 1409 410 1454 411
tri 1320 409 1354 410 ne
rect 533 408 597 409
tri 597 408 600 409 sw
tri 814 408 818 409 se
rect 818 408 873 409
tri 402 395 426 408 se
rect 426 400 459 408
tri 459 400 477 408 sw
tri 532 400 533 408 se
rect 533 400 600 408
rect 426 395 477 400
rect 160 392 194 395
rect 28 379 106 391
rect 28 345 66 379
rect 100 347 105 379
tri 105 349 106 379 nw
tri 154 379 158 391 se
rect 158 386 194 392
tri 194 386 203 395 nw
tri 395 391 402 395 se
rect 402 393 477 395
tri 477 393 485 400 sw
rect 402 391 485 393
tri 531 392 532 399 se
rect 532 395 600 400
tri 600 395 604 408 sw
rect 532 392 604 395
rect 531 391 604 392
rect 158 383 192 386
tri 192 383 194 386 nw
tri 381 384 395 391 se
rect 395 384 485 391
rect 158 379 191 383
tri 191 380 192 383 nw
tri 145 349 154 378 se
rect 154 349 183 379
rect 100 345 104 347
tri 104 345 105 347 nw
tri 143 345 145 349 se
rect 145 347 183 349
tri 183 348 191 379 nw
rect 415 379 485 384
rect 415 350 450 379
tri 381 348 386 350 ne
rect 386 348 450 350
rect 145 345 182 347
tri 182 345 183 347 nw
tri 386 345 389 348 ne
rect 389 345 450 348
rect 484 345 485 379
tri 530 384 531 391 se
rect 531 384 603 391
tri 603 384 604 391 nw
tri 809 406 814 408 se
rect 814 406 873 408
tri 873 406 875 409 sw
tri 1403 406 1407 409 se
rect 1407 406 1454 410
rect 530 379 603 384
tri 529 370 530 377 se
rect 530 370 554 379
tri 27 340 28 345 se
rect 28 340 102 345
tri 102 340 104 345 nw
rect 143 344 182 345
tri 142 340 143 344 se
rect 143 340 180 344
rect 27 337 101 340
tri 101 338 102 340 nw
tri 141 338 142 340 se
rect 142 338 180 340
rect 61 335 100 337
tri 100 336 101 337 nw
rect 61 334 99 335
tri 99 334 100 335 nw
tri 140 334 141 335 se
rect 141 334 180 338
tri 180 336 182 344 nw
tri 389 340 396 345 ne
rect 396 340 485 345
tri 527 347 529 369 se
rect 529 347 554 370
rect 527 345 554 347
rect 588 369 603 379
tri 664 379 666 384 se
tri 661 370 664 377 se
rect 664 370 666 379
rect 588 345 601 369
tri 601 345 603 369 nw
tri 652 345 661 369 se
rect 661 350 666 370
rect 843 405 875 406
tri 875 405 876 406 sw
rect 843 379 876 405
tri 1012 402 1015 404 se
rect 1015 402 1090 404
tri 1090 402 1099 404 sw
tri 1399 402 1403 406 se
rect 1403 402 1454 406
tri 1454 402 1467 415 sw
rect 1564 425 1569 447
rect 1626 427 1660 443
rect 1818 477 1852 527
rect 1818 427 1852 443
tri 1569 425 1570 427 sw
rect 1564 413 1570 425
rect 1543 404 1570 413
tri 1509 402 1513 404 ne
rect 1513 402 1570 404
tri 1007 400 1012 402 se
rect 1012 400 1101 402
rect 661 345 697 350
tri 697 345 700 350 nw
tri 808 350 809 370 se
rect 809 350 842 372
rect 808 347 842 350
tri 808 345 809 347 ne
rect 809 345 842 347
tri 1005 399 1007 400 se
rect 1007 399 1101 400
tri 1101 399 1107 402 sw
tri 1395 399 1398 402 se
rect 1398 400 1467 402
tri 1467 400 1470 402 sw
tri 1513 400 1519 402 ne
rect 1519 400 1570 402
rect 1398 399 1470 400
rect 1005 392 1107 399
tri 1107 392 1120 399 sw
tri 1393 394 1395 399 se
rect 1395 398 1470 399
tri 1470 398 1472 400 sw
tri 1520 398 1526 400 ne
rect 1526 398 1570 400
rect 1395 394 1472 398
tri 1228 392 1253 394 se
tri 1253 393 1265 394 sw
rect 1253 392 1265 393
tri 1265 392 1266 393 sw
tri 1391 392 1393 394 se
rect 1393 393 1472 394
tri 1472 393 1474 398 sw
rect 1393 392 1474 393
tri 1526 392 1549 398 ne
rect 1549 397 1570 398
tri 1549 392 1570 397 nw
rect 1005 389 1122 392
tri 1122 389 1126 392 sw
tri 1193 389 1220 392 se
rect 1220 389 1268 392
tri 1268 389 1275 392 sw
tri 1389 389 1391 392 se
rect 1391 389 1474 392
rect 1005 384 1275 389
tri 1275 384 1286 389 sw
tri 1387 384 1389 389 se
rect 1389 385 1474 389
tri 1474 385 1477 392 sw
rect 1389 384 1477 385
tri 1668 384 1691 392 se
rect 1691 384 1756 392
tri 1756 384 1763 392 sw
rect 1005 383 1286 384
tri 1286 383 1290 384 sw
tri 1386 383 1387 384 se
rect 1387 383 1477 384
rect 1005 379 1290 383
tri 1290 379 1297 383 sw
tri 1385 381 1386 383 se
rect 1386 381 1477 383
tri 1384 380 1385 381 se
rect 1385 380 1477 381
rect 1384 379 1477 380
tri 1660 379 1668 384 se
rect 1668 379 1763 384
tri 396 336 402 340 ne
rect 402 336 485 340
tri 402 334 403 336 ne
rect 403 335 485 336
rect 403 334 471 335
rect 61 330 94 334
tri 94 330 99 334 nw
tri 139 330 140 334 se
rect 140 330 179 334
tri 179 330 180 334 nw
tri 235 330 242 334 se
rect 242 330 286 334
rect 61 319 80 330
tri 80 319 94 330 nw
tri 136 320 139 330 se
rect 139 320 177 330
rect 136 319 177 320
tri 177 319 179 330 nw
tri 232 320 235 330 se
rect 235 320 286 330
rect 61 307 64 319
tri 64 307 80 319 nw
tri 132 307 136 319 se
rect 136 316 176 319
tri 176 316 177 319 nw
tri 231 316 232 319 se
rect 232 316 286 320
rect 136 307 172 316
tri 61 303 64 307 nw
tri 130 299 132 307 se
rect 132 299 172 307
tri 172 300 176 316 nw
tri 226 300 231 316 se
rect 231 300 286 316
tri 403 320 423 334 ne
rect 423 320 471 334
tri 471 320 485 335 nw
tri 526 336 527 340 se
rect 527 336 601 345
tri 651 341 652 344 se
rect 652 341 695 345
tri 695 341 697 345 nw
tri 809 341 813 345 ne
rect 813 341 863 345
tri 863 341 876 345 nw
tri 1004 349 1005 370 se
rect 1005 349 1042 379
rect 1004 345 1042 349
rect 1076 345 1234 379
rect 1268 378 1297 379
tri 1297 378 1299 379 sw
tri 1383 378 1384 379 se
rect 1384 378 1426 379
rect 1268 374 1299 378
tri 1299 374 1315 378 sw
tri 1380 374 1383 378 se
rect 1383 374 1426 378
rect 1268 373 1315 374
tri 1315 373 1320 374 sw
tri 1378 373 1380 374 se
rect 1380 373 1426 374
rect 1268 368 1320 373
tri 1320 368 1336 373 sw
tri 1375 368 1378 373 se
rect 1378 368 1426 373
rect 1268 365 1336 368
tri 1336 365 1356 368 sw
tri 1356 365 1373 368 se
rect 1373 365 1426 368
rect 1268 345 1426 365
rect 1460 345 1477 379
tri 1650 373 1660 379 se
rect 1660 373 1722 379
tri 1589 345 1650 373 se
rect 1650 345 1722 373
rect 1756 377 1763 379
tri 1763 377 1770 384 sw
rect 1756 372 1769 377
tri 1769 373 1770 377 nw
rect 1756 345 1768 372
rect 1004 344 1477 345
rect 1004 343 1260 344
tri 1260 343 1265 344 nw
tri 1265 343 1273 344 ne
rect 1273 343 1477 344
rect 1004 341 1249 343
tri 1249 341 1257 343 nw
tri 1278 341 1301 343 ne
rect 1301 341 1476 343
tri 1476 342 1477 343 nw
tri 1583 342 1589 345 se
rect 1589 342 1768 345
tri 649 336 651 341 se
rect 651 336 692 341
tri 692 337 695 341 nw
tri 813 337 828 341 ne
rect 828 337 848 341
tri 828 336 829 337 ne
rect 829 336 848 337
tri 848 336 863 341 nw
tri 1004 336 1007 341 ne
rect 1007 339 1237 341
tri 1237 340 1249 341 nw
tri 1301 340 1310 341 ne
rect 1310 340 1474 341
tri 1310 339 1311 340 ne
rect 1311 339 1474 340
rect 1007 336 1230 339
rect 526 334 601 336
tri 423 316 435 320 ne
rect 435 318 469 320
tri 469 318 471 320 nw
tri 435 316 469 318 nw
rect 560 330 601 334
tri 647 332 649 336 se
rect 649 332 690 336
tri 690 332 692 336 nw
tri 829 334 839 336 ne
tri 839 334 848 336 nw
tri 1007 332 1011 336 ne
rect 1011 332 1230 336
tri 1230 332 1237 339 nw
tri 1311 335 1318 339 ne
rect 1318 336 1474 339
tri 1474 336 1476 341 nw
tri 1572 336 1583 342 se
rect 1583 336 1768 342
tri 1768 336 1769 372 nw
rect 1318 335 1472 336
tri 1318 332 1324 335 ne
rect 1324 333 1472 335
tri 1472 333 1474 336 nw
rect 1324 332 1471 333
tri 1471 332 1472 333 nw
tri 1568 332 1572 336 se
rect 1572 332 1768 336
rect 560 321 600 330
tri 600 322 601 330 nw
tri 644 322 647 332 se
rect 647 322 684 332
tri 684 322 690 332 nw
tri 1011 322 1084 332 ne
rect 1084 323 1222 332
tri 1222 323 1230 332 nw
tri 1324 323 1337 332 ne
rect 1337 323 1459 332
tri 1459 323 1471 332 nw
tri 1560 323 1568 332 se
rect 1568 330 1768 332
rect 1568 323 1763 330
rect 1084 322 1215 323
rect 560 311 594 321
tri 594 311 600 321 nw
tri 639 311 644 322 se
rect 644 311 677 322
rect 560 307 582 311
tri 582 307 594 311 nw
tri 638 308 639 311 se
rect 639 308 677 311
tri 677 308 684 322 nw
tri 1084 308 1189 322 ne
rect 1189 316 1215 322
tri 1215 316 1222 323 nw
tri 1337 322 1340 323 ne
rect 1340 322 1453 323
tri 1453 322 1459 323 nw
tri 1559 322 1560 323 se
rect 1560 322 1763 323
tri 1763 322 1768 330 nw
tri 1340 321 1341 322 ne
rect 1341 321 1425 322
tri 1425 321 1429 322 nw
tri 1429 321 1441 322 ne
rect 1441 321 1449 322
tri 1449 321 1453 322 nw
tri 1341 316 1350 321 ne
rect 1350 316 1397 321
tri 1397 316 1420 321 nw
rect 1189 312 1212 316
tri 1212 312 1215 316 nw
tri 1350 312 1356 316 ne
rect 1356 312 1387 316
rect 1189 309 1209 312
tri 1209 309 1212 312 nw
tri 1356 310 1362 312 ne
rect 1362 310 1387 312
tri 1387 310 1397 316 nw
tri 1558 310 1559 315 se
rect 1559 310 1755 322
tri 1362 309 1363 310 ne
rect 1363 309 1382 310
rect 1189 308 1205 309
tri 1205 308 1209 309 nw
tri 1363 308 1367 309 ne
rect 1367 308 1382 309
tri 1382 308 1387 310 nw
rect 1558 309 1755 310
tri 1755 309 1763 322 nw
rect 560 306 581 307
tri 581 306 582 307 nw
rect 638 306 676 308
tri 676 307 677 308 nw
tri 1189 307 1199 308 ne
rect 1199 307 1202 308
tri 1202 307 1205 308 nw
tri 560 300 581 306 nw
tri 635 300 638 306 se
rect 638 300 661 306
tri 126 286 130 299 se
rect 130 286 169 299
tri 169 287 172 299 nw
tri 222 287 226 299 se
rect 226 297 271 300
tri 271 297 275 300 nw
tri 634 297 635 299 se
rect 635 297 661 300
rect 226 287 264 297
tri 122 282 126 286 se
rect 126 282 168 286
tri 168 282 169 286 nw
tri 220 283 222 287 se
rect 222 283 264 287
tri 120 281 122 282 se
rect 122 281 168 282
rect 220 281 264 283
tri 264 281 271 297 nw
tri 628 281 634 297 se
rect 634 281 661 297
tri 661 281 676 306 nw
tri 108 273 120 281 se
rect 120 279 167 281
tri 167 279 168 281 nw
tri 219 279 220 281 se
rect 220 279 261 281
rect 120 273 166 279
tri 166 273 167 279 nw
tri 218 274 219 279 se
rect 219 274 261 279
rect 218 273 261 274
tri 261 273 264 281 nw
tri 619 273 628 281 se
rect 628 273 657 281
tri 657 273 661 281 nw
tri 106 269 108 273 se
rect 108 269 165 273
tri 165 269 166 273 nw
tri 216 269 217 273 se
rect 217 269 256 273
tri 103 260 106 269 se
rect 106 260 163 269
tri 163 260 165 269 nw
tri 214 261 216 268 se
rect 216 261 256 269
tri 102 256 103 260 se
rect 103 256 162 260
tri 162 256 163 260 nw
tri 212 256 214 260 se
rect 214 259 256 261
tri 256 260 261 273 nw
tri 604 260 619 273 se
rect 619 260 650 273
tri 650 260 657 273 nw
tri 793 266 796 273 se
rect 796 266 802 273
tri 603 259 604 260 se
rect 604 259 648 260
rect 214 256 253 259
rect 102 255 162 256
rect 212 255 253 256
tri 253 255 256 259 nw
tri 602 256 603 259 se
rect 603 258 648 259
tri 648 258 650 260 nw
rect 603 256 647 258
tri 101 250 102 255 se
rect 102 250 160 255
tri 160 250 162 255 nw
tri 210 250 212 255 se
rect 212 250 249 255
tri 249 250 253 255 nw
tri 293 250 300 255 se
rect 300 250 345 255
rect 101 249 160 250
tri 98 241 101 249 se
rect 101 241 114 249
tri 98 235 100 241 ne
rect 100 235 114 241
tri 100 215 114 235 ne
rect 148 239 158 249
tri 158 241 160 249 nw
rect 210 249 249 250
rect 293 249 345 250
rect 148 235 156 239
tri 156 235 158 239 nw
tri 148 216 156 235 nw
tri 244 242 249 249 nw
tri 289 242 293 249 se
rect 293 242 306 249
tri 280 226 289 242 se
rect 289 226 306 242
tri 210 213 218 215 ne
rect 218 213 236 215
tri 236 213 244 215 nw
tri 278 220 280 226 se
rect 280 220 306 226
rect 340 247 345 249
tri 345 247 353 255 sw
tri 601 253 602 254 se
rect 602 253 647 256
tri 647 253 648 258 nw
tri 425 249 444 250 se
rect 444 249 450 250
tri 450 249 452 250 sw
rect 601 249 646 253
tri 646 249 647 253 nw
rect 793 249 802 266
tri 836 267 837 273 sw
rect 1264 271 1298 273
tri 1298 271 1316 307 sw
rect 1558 306 1754 309
tri 1754 307 1755 309 nw
tri 1794 307 1795 309 se
tri 1556 286 1558 306 se
rect 1558 296 1738 306
tri 1738 296 1754 306 nw
tri 1789 296 1794 306 se
rect 1794 296 1795 307
rect 1558 286 1675 296
tri 1675 286 1738 296 nw
tri 1785 286 1789 296 se
rect 1789 286 1795 296
tri 1414 281 1426 286 se
tri 1403 273 1414 281 se
rect 1414 273 1426 281
tri 923 268 938 270 se
tri 938 268 958 270 sw
rect 1264 268 1316 271
rect 836 253 837 267
tri 919 266 923 268 se
rect 923 266 958 268
tri 837 253 839 266 sw
rect 836 249 839 253
rect 340 219 352 247
tri 352 226 353 247 nw
rect 436 248 452 249
tri 452 248 453 249 sw
rect 436 247 453 248
tri 453 247 456 248 sw
rect 436 240 456 247
tri 456 240 459 247 sw
rect 436 235 459 240
rect 340 215 350 219
tri 350 215 352 219 nw
rect 312 214 350 215
rect 312 212 349 214
tri 349 212 350 214 nw
rect 312 186 315 212
tri 315 186 349 212 nw
rect 402 208 425 215
tri 402 204 406 208 ne
rect 406 204 425 208
tri 406 201 425 204 ne
rect 601 215 602 249
rect 636 247 646 249
tri 696 248 697 249 se
rect 697 248 698 249
tri 691 247 696 248 se
rect 696 247 698 248
rect 636 215 638 247
tri 638 215 646 247 nw
tri 680 244 691 247 se
rect 691 244 698 247
rect 601 213 638 215
rect 714 213 727 215
tri 727 213 732 215 nw
rect 793 215 794 249
rect 836 239 838 249
rect 828 215 838 239
tri 838 215 839 249 nw
tri 890 249 919 266 se
rect 919 249 958 266
tri 958 249 1118 268 sw
tri 1264 251 1266 268 ne
rect 1266 257 1316 268
tri 1316 257 1320 271 sw
tri 1382 259 1403 273 se
rect 1403 259 1426 273
rect 1266 249 1320 257
rect 924 222 1090 249
rect 924 219 941 222
tri 941 219 953 222 nw
tri 953 219 968 222 ne
rect 968 219 1047 222
tri 924 215 941 219 nw
tri 968 215 976 219 ne
rect 976 215 1047 219
rect 793 213 838 215
tri 976 213 979 215 ne
rect 979 213 1047 215
tri 714 210 727 213 nw
tri 793 210 799 213 ne
rect 799 212 838 213
rect 799 210 831 212
tri 799 203 811 210 ne
rect 811 203 831 210
tri 831 203 838 212 nw
tri 979 204 999 213 ne
rect 999 204 1047 213
tri 811 201 816 203 ne
rect 816 201 820 203
tri 816 200 820 201 ne
tri 820 200 831 203 nw
tri 999 200 1007 204 ne
rect 1007 200 1047 204
tri 1007 195 1018 200 ne
rect 1018 195 1047 200
tri 1018 187 1032 195 ne
rect 1032 188 1047 195
rect 1081 215 1090 222
rect 1081 204 1117 215
tri 1117 204 1124 215 nw
tri 1220 239 1229 249 sw
tri 1267 241 1268 249 ne
rect 1220 232 1229 239
tri 1229 232 1234 239 sw
rect 1268 232 1282 249
tri 1268 222 1270 232 ne
rect 1270 222 1282 232
tri 1270 216 1273 222 ne
tri 1186 204 1195 215 ne
rect 1195 204 1200 215
rect 1081 195 1111 204
tri 1111 195 1117 204 nw
tri 1195 198 1200 204 ne
rect 1273 215 1282 222
rect 1316 220 1319 249
tri 1319 222 1320 249 nw
tri 1378 253 1382 259 se
rect 1382 253 1426 259
rect 1378 252 1426 253
rect 1556 285 1666 286
tri 1666 285 1675 286 nw
tri 1784 285 1785 286 se
rect 1785 285 1795 286
tri 1554 260 1556 285 se
rect 1556 283 1660 285
tri 1660 283 1666 285 nw
rect 1556 260 1630 283
rect 1554 259 1630 260
tri 1630 259 1660 283 nw
tri 1773 259 1784 283 se
rect 1784 275 1795 285
tri 1829 279 1832 309 sw
rect 1829 275 1832 279
rect 1784 260 1832 275
tri 1832 260 1834 275 sw
rect 1784 259 1834 260
rect 1378 249 1459 252
tri 1459 250 1460 252 nw
tri 1553 252 1554 259 se
rect 1554 252 1621 259
tri 1621 252 1630 259 nw
tri 1771 252 1773 259 se
rect 1773 252 1834 259
rect 1553 249 1619 252
tri 1619 249 1621 252 nw
tri 1770 249 1771 252 se
rect 1771 251 1834 252
tri 1834 251 1835 259 sw
rect 1771 249 1835 251
rect 1316 215 1318 220
tri 1318 215 1319 220 nw
rect 1412 240 1454 249
tri 1454 240 1459 249 nw
tri 1552 240 1553 249 se
rect 1553 240 1578 249
rect 1412 228 1447 240
tri 1447 228 1454 240 nw
rect 1552 235 1578 240
rect 1612 239 1617 249
tri 1617 245 1619 249 nw
tri 1552 228 1554 235 ne
rect 1554 228 1578 235
rect 1412 222 1440 228
tri 1440 222 1447 228 nw
tri 1554 222 1555 228 ne
rect 1412 221 1439 222
tri 1439 221 1440 222 nw
rect 1555 221 1578 228
tri 1412 215 1439 221 nw
tri 1556 215 1564 221 ne
rect 1564 215 1578 221
rect 1614 223 1617 239
tri 1617 223 1618 235 sw
tri 1273 214 1274 215 ne
rect 1274 214 1318 215
tri 1564 214 1566 215 ne
rect 1566 214 1580 215
tri 1566 205 1580 214 ne
rect 1614 207 1618 223
tri 1708 231 1736 249 sw
rect 1804 240 1831 249
tri 1831 240 1835 249 nw
rect 1804 235 1829 240
tri 1829 235 1831 240 nw
tri 1804 215 1829 235 nw
tri 1618 207 1619 215 sw
rect 1614 205 1615 207
tri 1615 205 1619 207 nw
rect 1674 199 1702 215
tri 1674 195 1678 199 ne
rect 1678 197 1702 199
rect 1678 195 1718 197
rect 1081 188 1106 195
rect 1032 187 1106 188
tri 1106 187 1111 195 nw
tri 1678 191 1683 195 ne
rect 1683 191 1718 195
tri 1718 191 1736 197 nw
tri 1683 190 1717 191 ne
tri 1717 190 1718 191 nw
tri 1032 186 1035 187 ne
rect 1035 186 1104 187
tri 1035 178 1074 186 ne
rect 1074 184 1104 186
tri 1104 184 1106 187 nw
rect 1074 179 1097 184
tri 1097 179 1104 184 nw
rect 1074 178 1084 179
tri 1084 178 1097 179 nw
tri 895 173 903 175 se
tri 903 174 977 175 sw
rect 903 173 977 174
tri 888 170 895 173 se
rect 895 170 977 173
tri 977 170 980 173 sw
tri 884 169 888 170 se
rect 888 169 980 170
tri 980 169 982 170 sw
tri 877 167 884 169 se
rect 884 167 934 169
tri 338 153 340 160 se
tri 175 146 193 153 sw
tri 335 146 338 153 se
rect 338 146 340 153
rect 175 140 193 146
tri 193 140 199 146 sw
rect 175 135 199 140
tri 199 135 205 140 sw
tri 332 137 335 146 se
rect 335 137 340 146
rect 175 133 205 135
tri 205 133 208 135 sw
tri 331 133 332 135 se
rect 332 133 340 137
rect 175 129 208 133
tri 208 129 209 133 sw
rect 175 121 209 129
tri 330 129 331 132 se
rect 331 129 340 133
tri 329 126 330 128 se
rect 330 126 340 129
tri 374 142 395 160 sw
tri 640 143 654 151 se
rect 374 135 395 142
tri 639 140 640 142 se
rect 640 140 654 143
tri 395 135 397 140 sw
tri 637 135 639 140 se
rect 639 135 654 140
rect 374 133 397 135
tri 397 133 398 135 sw
tri 636 133 637 135 se
rect 637 133 654 135
rect 374 129 398 133
tri 398 129 399 133 sw
rect 374 127 399 129
tri 399 127 400 128 sw
rect 374 126 400 127
tri 209 121 211 126 sw
rect 175 119 211 121
tri 328 121 329 126 se
rect 329 121 400 126
tri 400 121 401 126 sw
tri 140 117 141 119 se
rect 141 117 211 119
tri 327 117 328 119 se
rect 328 118 401 121
tri 401 118 402 121 sw
rect 328 117 402 118
rect 636 117 654 133
tri 688 144 689 151 sw
rect 688 138 689 144
tri 689 138 690 143 sw
rect 688 134 690 138
tri 690 134 691 135 sw
rect 688 129 691 134
rect 911 135 934 167
rect 968 135 982 169
rect 911 133 982 135
tri 1390 179 1391 181 sw
rect 1390 178 1391 179
tri 1391 178 1392 179 sw
rect 1390 175 1392 178
tri 1392 175 1394 178 sw
rect 1390 170 1394 175
tri 1394 170 1399 175 sw
rect 1390 167 1399 170
tri 1399 167 1403 170 sw
rect 1390 147 1403 167
rect 1356 146 1403 147
tri 1403 146 1426 167 sw
tri 1356 133 1358 146 ne
rect 1358 133 1426 146
tri 691 129 692 133 sw
tri 877 129 884 133 ne
rect 884 132 982 133
rect 884 129 980 132
tri 980 129 982 132 nw
tri 1358 129 1359 133 ne
rect 688 126 692 129
tri 884 128 887 129 ne
rect 887 128 979 129
tri 979 128 980 129 nw
rect 1359 128 1426 133
tri 692 126 693 128 sw
tri 887 126 892 128 ne
rect 892 126 978 128
tri 978 126 979 128 nw
tri 1056 126 1062 128 se
rect 688 121 693 126
tri 693 121 694 126 sw
tri 892 121 914 126 ne
rect 914 123 976 126
tri 976 123 978 126 nw
tri 1044 123 1056 126 se
rect 1056 123 1062 126
rect 914 121 966 123
tri 966 121 976 123 nw
tri 1035 121 1044 123 se
rect 1044 121 1062 123
rect 688 117 694 121
tri 914 117 927 121 ne
rect 927 117 953 121
tri 953 117 966 121 nw
tri 1034 117 1035 121 se
rect 1035 117 1062 121
rect 66 101 100 117
tri 136 101 140 117 se
rect 140 101 211 117
tri 211 101 215 117 sw
rect 258 101 292 117
tri 135 95 136 99 se
rect 136 95 162 101
tri 135 71 137 95 ne
rect 137 71 162 95
tri 137 67 140 71 ne
rect 140 67 162 71
rect 196 98 215 101
tri 215 98 216 101 sw
rect 196 95 216 98
rect 196 67 215 95
tri 215 71 216 95 nw
rect 66 17 100 67
tri 140 59 148 67 ne
rect 148 66 215 67
rect 148 59 208 66
tri 208 59 215 66 nw
rect 327 116 402 117
rect 327 103 400 116
tri 400 103 402 116 nw
rect 327 101 397 103
rect 327 97 354 101
tri 327 88 330 97 ne
rect 330 88 354 97
tri 330 67 354 88 ne
rect 388 97 397 101
tri 397 97 400 103 nw
rect 450 101 484 117
rect 388 88 395 97
tri 395 89 397 97 nw
rect 388 71 389 88
tri 389 71 395 88 nw
tri 388 67 389 71 nw
tri 148 58 208 59 ne
rect 258 17 292 67
rect 450 17 484 67
rect 554 101 588 117
rect 636 101 694 117
rect 746 101 780 117
tri 927 116 932 117 ne
rect 932 116 948 117
tri 948 116 953 117 nw
tri 932 115 945 116 ne
tri 945 115 948 116 nw
tri 1031 102 1034 115 se
rect 1034 102 1062 117
rect 1031 101 1062 102
tri 1359 127 1360 128 ne
tri 1096 121 1098 126 sw
rect 1360 123 1426 128
tri 1426 123 1453 146 sw
tri 1545 158 1552 166 sw
rect 1545 146 1552 158
tri 1552 146 1564 158 sw
rect 1545 143 1564 146
tri 1564 143 1568 146 sw
rect 1545 133 1568 143
tri 1568 133 1579 143 sw
rect 1545 132 1579 133
tri 1360 121 1362 123 ne
rect 1362 121 1453 123
rect 1096 102 1098 121
tri 1098 102 1101 117 sw
tri 635 71 636 101 se
rect 636 71 650 101
tri 635 67 637 71 ne
rect 637 67 650 71
rect 684 75 694 101
tri 694 75 696 101 sw
rect 684 71 695 75
tri 695 71 696 75 nw
rect 684 67 693 71
tri 693 67 695 71 nw
rect 554 17 588 67
tri 637 56 643 67 ne
rect 643 66 693 67
rect 643 59 690 66
tri 690 59 693 66 nw
rect 643 56 682 59
tri 682 56 690 59 nw
tri 643 54 676 56 ne
tri 676 54 682 56 nw
rect 746 17 780 67
tri 1025 77 1031 101 se
rect 1031 77 1042 101
rect 1096 94 1101 102
rect 1234 101 1268 117
tri 1362 111 1367 121 ne
rect 1367 117 1453 121
tri 1453 117 1459 123 sw
rect 1511 120 1579 132
tri 1579 120 1584 133 sw
rect 1511 117 1584 120
rect 1367 114 1459 117
tri 1459 114 1463 117 sw
rect 1367 111 1463 114
tri 1367 101 1380 111 ne
rect 1380 102 1463 111
tri 1463 102 1467 114 sw
rect 1380 101 1467 102
rect 1511 101 1583 117
tri 1583 101 1584 117 nw
rect 1626 101 1660 117
rect 1025 67 1042 77
rect 1076 84 1101 94
tri 1101 84 1105 101 sw
rect 1076 77 1103 84
tri 1103 77 1105 84 nw
rect 1076 68 1101 77
tri 1101 68 1103 77 nw
rect 1076 67 1079 68
rect 1025 65 1079 67
tri 1025 54 1038 65 ne
rect 1038 57 1079 65
tri 1079 57 1101 68 nw
tri 1380 67 1426 101 ne
rect 1460 75 1462 101
tri 1462 75 1467 101 nw
tri 1510 75 1511 101 se
rect 1511 75 1530 101
tri 1460 67 1462 75 nw
rect 1510 71 1530 75
tri 1510 67 1512 71 ne
rect 1512 67 1530 71
rect 1564 94 1583 101
rect 1564 70 1582 94
tri 1582 71 1583 94 nw
rect 1564 67 1580 70
tri 1580 68 1582 70 nw
rect 1038 54 1039 57
tri 1039 54 1079 57 nw
rect 1234 17 1268 67
tri 1512 56 1517 67 ne
rect 1517 59 1573 67
tri 1573 59 1580 67 nw
rect 1765 134 1877 143
tri 1877 134 1888 143 sw
rect 1765 119 1888 134
tri 1888 119 1891 133 sw
rect 1765 117 1891 119
tri 1891 117 1892 119 sw
rect 1765 109 1892 117
rect 1731 102 1892 109
tri 1892 102 1895 117 sw
rect 1731 101 1894 102
tri 1731 89 1740 101 ne
rect 1740 89 1818 101
tri 1740 67 1779 89 ne
rect 1779 67 1818 89
rect 1852 84 1894 101
tri 1894 89 1895 102 nw
rect 1852 67 1885 84
rect 1517 56 1569 59
tri 1569 56 1573 59 nw
tri 1517 52 1538 56 ne
rect 1538 52 1560 56
tri 1560 52 1569 56 nw
rect 1626 17 1660 67
tri 1779 62 1788 67 ne
rect 1788 63 1885 67
tri 1885 63 1894 84 nw
rect 1788 62 1884 63
tri 1884 62 1885 63 nw
tri 1788 56 1805 62 ne
rect 1805 57 1880 62
tri 1880 57 1884 62 nw
rect 1805 56 1877 57
tri 1877 56 1880 57 nw
tri 1805 52 1866 56 ne
tri 1866 52 1877 56 nw
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 169 395 203 429
rect 1320 413 1330 444
rect 1330 413 1354 444
rect 1320 410 1354 413
rect 381 350 415 384
rect 27 303 61 337
rect 666 350 700 384
rect 809 379 843 406
rect 1509 413 1530 438
rect 1530 413 1543 438
rect 1509 404 1543 413
rect 809 372 842 379
rect 842 372 843 379
rect 286 300 320 334
rect 526 300 560 334
rect 1264 273 1298 307
rect 802 249 836 273
rect 278 215 306 220
rect 306 215 312 220
rect 425 215 436 235
rect 436 215 459 235
rect 278 186 312 215
rect 425 201 459 215
rect 680 215 698 244
rect 698 215 714 244
rect 680 210 714 215
rect 802 239 828 249
rect 828 239 836 249
rect 1047 188 1081 222
rect 1200 215 1220 232
rect 1220 215 1234 232
rect 1200 198 1234 215
rect 1426 252 1460 286
rect 1795 275 1829 309
rect 1580 215 1612 239
rect 1612 215 1614 239
rect 1580 205 1614 215
rect 1702 215 1708 231
rect 1708 215 1736 231
rect 1702 197 1736 215
rect 141 119 175 153
rect 340 126 374 160
rect 654 117 688 151
rect 877 133 911 167
rect 1356 147 1390 181
rect 1062 101 1096 128
rect 1511 132 1545 166
rect 1062 94 1076 101
rect 1076 94 1096 101
rect 1731 109 1765 143
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
tri 1507 449 1544 450 se
tri 1544 449 1545 450 sw
tri 1316 445 1318 449 se
rect 1318 445 1355 449
tri 1355 445 1357 449 sw
tri 1503 445 1507 449 se
rect 1507 445 1545 449
tri 1545 445 1550 449 sw
rect 1316 444 1357 445
tri 1357 444 1358 445 sw
tri 165 430 167 433 se
rect 167 430 204 433
tri 204 430 207 433 sw
rect 165 429 207 430
rect 165 395 169 429
rect 203 422 207 429
tri 207 422 211 430 sw
rect 203 421 211 422
tri 211 421 219 422 sw
rect 203 420 219 421
tri 219 420 225 421 sw
tri 814 420 825 421 se
tri 825 420 828 421 sw
rect 203 410 225 420
tri 225 410 287 420 sw
rect 203 409 287 410
tri 287 409 295 410 sw
rect 203 395 295 409
rect 165 393 295 395
tri 165 391 167 393 ne
rect 167 391 295 393
tri 204 389 214 391 ne
rect 214 389 295 391
tri 214 388 217 389 ne
rect 217 388 295 389
tri 219 386 228 388 ne
rect 228 386 295 388
tri 228 384 239 386 ne
rect 239 384 295 386
tri 239 379 268 384 ne
rect 268 379 295 384
tri 268 369 295 379 ne
tri 788 410 814 420 se
rect 814 418 828 420
tri 828 418 835 420 sw
rect 814 410 835 418
tri 780 407 788 410 se
rect 788 407 835 410
tri 779 406 780 407 se
rect 780 406 835 407
tri 835 406 850 418 sw
rect 1316 410 1320 444
rect 1354 442 1358 444
tri 1358 442 1359 444 sw
rect 1354 410 1359 442
rect 1316 408 1359 410
rect 1503 438 1549 445
rect 1503 430 1509 438
tri 1503 408 1505 430 ne
tri 1316 406 1317 408 ne
rect 1317 406 1358 408
tri 1358 406 1359 408 nw
tri 775 405 779 406 se
rect 779 405 809 406
tri 771 403 775 405 se
rect 775 403 809 405
tri 735 389 771 403 se
rect 771 389 809 403
tri 702 388 735 389 se
rect 735 388 809 389
tri 377 386 379 388 se
rect 379 386 417 388
tri 417 386 418 388 sw
rect 664 387 809 388
rect 843 405 850 406
tri 850 405 853 406 sw
rect 843 403 853 405
tri 853 403 855 405 sw
tri 1317 403 1320 406 ne
rect 1320 404 1358 406
rect 843 400 855 403
tri 855 400 859 403 sw
rect 377 384 419 386
tri 663 385 664 386 se
rect 664 385 790 387
rect 663 384 790 385
rect 377 350 381 384
rect 415 350 419 384
rect 377 348 419 350
tri 377 346 379 348 ne
rect 379 346 419 348
tri 23 339 26 341 se
rect 26 339 39 341
rect 23 337 39 339
rect 23 303 27 337
rect 23 302 39 303
tri 23 299 26 302 ne
rect 26 299 39 302
tri 26 298 28 299 ne
rect 28 298 39 299
tri 28 296 33 298 ne
rect 33 296 39 298
tri 34 294 36 296 ne
rect 36 294 39 296
tri 379 342 380 346 ne
rect 380 342 417 346
tri 417 342 419 346 nw
rect 704 351 790 384
rect 843 385 858 400
tri 858 390 859 400 nw
rect 1320 402 1357 404
tri 1357 403 1358 404 nw
rect 1505 404 1509 430
rect 1543 430 1549 438
tri 1549 430 1550 445 nw
rect 1543 406 1548 430
tri 1548 406 1549 430 nw
rect 1543 404 1547 406
rect 1505 403 1547 404
tri 1547 403 1548 406 nw
tri 1505 402 1506 403 ne
rect 1320 393 1356 402
tri 1356 397 1357 402 nw
rect 1506 396 1547 403
tri 1320 390 1321 393 ne
rect 1321 390 1356 393
tri 1321 386 1323 390 ne
rect 1323 388 1356 390
tri 1356 388 1357 393 sw
rect 843 372 856 385
rect 380 338 416 342
tri 416 339 417 342 nw
rect 300 336 322 338
tri 322 336 324 338 sw
rect 300 334 324 336
rect 320 300 324 334
rect 380 334 415 338
tri 415 335 416 338 nw
tri 522 335 524 338 se
rect 524 336 562 338
tri 562 336 564 338 sw
rect 524 335 564 336
rect 380 320 410 334
tri 410 320 415 334 nw
rect 522 334 564 335
tri 36 291 37 294 ne
rect 37 291 90 294
rect 300 298 324 300
tri 374 300 380 320 se
rect 380 300 403 320
tri 403 300 410 320 nw
rect 522 300 526 334
rect 560 313 564 334
rect 704 349 738 351
tri 738 349 749 351 nw
tri 749 349 773 351 ne
rect 773 349 790 351
rect 704 347 728 349
tri 728 347 738 349 nw
tri 773 347 790 349 ne
rect 704 345 717 347
tri 717 345 728 347 nw
rect 704 342 705 345
tri 705 342 717 345 nw
rect 842 362 856 372
tri 856 369 858 385 nw
rect 1323 385 1357 388
tri 1323 369 1331 385 ne
rect 1331 370 1357 385
tri 1357 370 1361 386 sw
rect 1331 367 1361 370
tri 1331 364 1332 367 ne
rect 1332 363 1361 367
tri 1063 362 1079 363 se
tri 1079 362 1094 363 sw
tri 1332 362 1333 363 ne
rect 842 361 855 362
tri 855 361 856 362 nw
tri 1054 361 1063 362 se
rect 1063 361 1094 362
tri 1094 361 1101 362 sw
rect 1333 361 1361 363
tri 1361 361 1362 369 sw
rect 842 358 853 361
tri 853 358 855 361 nw
tri 1025 358 1054 361 se
rect 1054 358 1101 361
tri 1101 358 1116 361 sw
rect 1333 358 1362 361
rect 842 357 852 358
tri 852 357 853 358 nw
tri 1023 357 1025 358 se
rect 1025 357 1116 358
rect 842 354 847 357
tri 847 354 852 357 nw
tri 1013 354 1023 357 se
rect 1023 354 1116 357
tri 1116 354 1133 358 sw
tri 1333 356 1334 358 ne
rect 842 352 844 354
tri 844 352 847 354 nw
tri 842 351 844 352 nw
tri 1003 349 1013 354 se
rect 1013 352 1133 354
tri 1133 352 1143 354 sw
rect 1334 352 1362 358
tri 1362 352 1364 361 sw
rect 1013 351 1143 352
tri 1143 351 1151 352 sw
rect 1013 349 1151 351
tri 1001 347 1003 349 se
rect 1003 347 1151 349
tri 1151 347 1169 351 sw
rect 1334 350 1364 352
tri 1334 347 1335 350 ne
rect 1335 347 1364 350
tri 1364 347 1365 350 sw
tri 996 345 1001 347 se
rect 1001 345 1169 347
tri 992 342 996 345 se
rect 996 342 1169 345
tri 991 341 992 342 se
rect 992 341 1169 342
tri 987 339 991 341 se
rect 991 339 1169 341
tri 984 338 987 339 se
rect 987 338 1169 339
tri 1169 338 1214 347 sw
tri 1335 339 1336 347 ne
rect 1336 338 1365 347
tri 1661 350 1671 351 se
rect 1671 350 1673 351
tri 1673 350 1684 351 sw
tri 1653 347 1661 350 se
rect 1661 347 1684 350
tri 1684 347 1706 350 sw
tri 1643 344 1653 347 se
rect 1653 344 1706 347
tri 980 335 984 338 se
rect 984 335 1214 338
tri 971 330 980 335 se
rect 980 331 1214 335
rect 980 330 1039 331
tri 1039 330 1048 331 nw
tri 1048 330 1061 331 ne
rect 1061 330 1214 331
tri 1214 330 1236 338 sw
tri 1336 331 1337 338 ne
tri 968 328 971 330 se
rect 971 329 1035 330
tri 1035 329 1039 330 nw
tri 1061 329 1068 330 ne
rect 1068 329 1236 330
rect 971 328 1001 329
tri 564 313 565 328 sw
rect 560 300 565 313
tri 936 309 968 328 se
rect 968 312 1001 328
tri 1001 312 1035 329 nw
tri 1068 312 1201 329 ne
rect 1201 328 1236 329
tri 1236 328 1241 330 sw
rect 1337 328 1365 338
tri 1365 328 1368 344 sw
rect 1201 312 1241 328
tri 1241 312 1280 328 sw
rect 1337 327 1368 328
tri 1583 327 1643 344 se
rect 1643 336 1706 344
tri 1706 336 1795 347 sw
rect 1643 327 1795 336
tri 1795 327 1811 336 sw
tri 1337 312 1339 327 ne
rect 1339 317 1368 327
tri 1368 317 1370 327 sw
tri 1548 317 1583 327 se
rect 1583 317 1811 327
rect 968 310 996 312
tri 996 310 1000 312 nw
tri 1202 310 1208 312 ne
rect 1208 311 1280 312
tri 1280 311 1300 312 sw
rect 1208 310 1300 311
rect 968 309 995 310
tri 995 309 996 310 nw
tri 1208 309 1209 310 ne
rect 1209 309 1300 310
tri 1300 309 1301 311 sw
rect 1339 309 1370 317
tri 1521 309 1548 317 se
rect 1548 315 1811 317
rect 1548 314 1686 315
tri 1686 314 1689 315 nw
tri 1706 314 1710 315 ne
rect 1710 314 1811 315
rect 1548 313 1680 314
tri 1680 313 1686 314 nw
tri 1710 313 1716 314 ne
rect 1716 313 1811 314
tri 1811 313 1835 327 sw
rect 1548 312 1676 313
tri 1676 312 1680 313 nw
tri 1716 312 1717 313 ne
rect 1717 312 1783 313
rect 1548 309 1663 312
tri 1663 309 1676 312 nw
tri 1717 309 1723 312 ne
rect 1723 309 1783 312
tri 1835 312 1837 313 sw
tri 933 307 936 309 se
rect 936 307 991 309
tri 991 307 995 309 nw
tri 1209 307 1213 309 ne
rect 1213 308 1301 309
tri 1301 308 1302 309 sw
rect 1213 307 1302 308
rect 374 299 403 300
rect 300 296 322 298
tri 322 296 324 298 nw
tri 373 296 374 299 se
rect 374 296 402 299
tri 402 296 403 299 nw
rect 522 299 565 300
tri 565 299 566 307 sw
rect 522 298 566 299
tri 918 298 933 307 se
rect 933 303 981 307
tri 981 303 991 307 nw
tri 1213 303 1222 307 ne
rect 1222 303 1264 307
rect 933 298 968 303
tri 522 296 524 298 ne
rect 524 296 566 298
tri 372 295 373 296 se
rect 373 295 402 296
tri 37 283 41 291 ne
rect 41 283 90 291
tri 90 283 91 291 sw
rect 41 282 91 283
tri 41 281 42 282 ne
rect 42 281 91 282
tri 368 282 372 294 se
rect 372 291 401 295
tri 401 294 402 295 nw
tri 524 294 525 296 ne
rect 372 282 398 291
tri 398 282 401 291 nw
rect 525 290 566 296
tri 909 293 918 298 se
rect 918 293 968 298
tri 904 291 909 293 se
rect 909 291 968 293
tri 902 290 904 291 se
rect 904 290 968 291
tri 968 290 981 303 nw
tri 1222 293 1240 303 ne
rect 1240 293 1264 303
tri 1240 291 1244 293 ne
rect 1244 291 1264 293
tri 1244 290 1245 291 ne
rect 1245 290 1264 291
tri 525 282 527 290 ne
rect 527 283 566 290
tri 566 283 567 290 sw
tri 851 285 902 290 se
rect 902 286 965 290
tri 965 286 968 290 nw
tri 1245 286 1253 290 ne
rect 1253 286 1264 290
rect 902 285 960 286
tri 830 283 851 285 se
rect 851 283 869 285
rect 527 282 567 283
tri 821 282 830 283 se
rect 830 282 869 283
rect 368 281 397 282
tri 397 281 398 282 nw
tri 527 281 528 282 ne
tri 42 277 43 281 ne
rect 43 278 91 281
tri 91 278 92 281 sw
rect 43 277 92 278
tri 367 278 368 281 se
rect 368 278 395 281
tri 43 274 44 277 ne
rect 44 273 92 277
tri 366 274 367 277 se
rect 367 274 395 278
tri 395 275 397 281 nw
rect 528 278 567 282
tri 816 281 821 282 se
rect 821 281 869 282
tri 567 278 568 281 sw
rect 528 275 568 278
tri 806 277 816 281 se
rect 816 277 869 281
rect 366 273 395 274
tri 528 273 529 275 ne
rect 529 273 568 275
tri 798 275 800 277 se
rect 800 275 869 277
rect 798 273 869 275
tri 44 258 52 273 ne
rect 52 258 92 273
tri 92 258 94 273 sw
tri 360 258 366 273 se
rect 366 258 388 273
tri 52 250 56 258 ne
rect 56 252 94 258
tri 94 252 95 258 sw
rect 56 248 95 252
tri 358 252 360 258 se
rect 360 252 388 258
tri 388 252 395 273 nw
tri 529 259 533 273 ne
tri 532 252 533 258 se
rect 533 252 568 273
tri 568 252 574 273 sw
tri 357 249 358 250 se
rect 358 249 387 252
tri 387 250 388 252 nw
rect 532 250 574 252
tri 574 250 575 252 sw
tri 529 249 531 250 se
rect 531 249 575 250
rect 357 248 386 249
tri 386 248 387 249 nw
tri 518 248 528 249 se
rect 528 248 575 249
tri 57 245 58 248 ne
rect 58 244 95 248
tri 356 245 357 248 se
rect 357 245 384 248
tri 58 240 60 244 ne
rect 60 240 95 244
tri 95 240 96 244 sw
rect 60 239 96 240
tri 354 240 356 244 se
rect 356 240 384 245
tri 384 240 386 248 nw
tri 440 240 518 248 se
rect 518 240 575 248
tri 575 240 577 248 sw
rect 354 239 384 240
rect 437 239 490 240
tri 60 235 62 239 ne
rect 62 235 96 239
tri 352 235 354 239 se
rect 354 235 382 239
tri 382 235 384 239 nw
tri 421 237 423 239 se
rect 423 237 490 239
rect 421 235 490 237
tri 62 234 63 235 ne
rect 63 234 96 235
tri 96 234 97 235 sw
tri 63 226 66 234 ne
rect 66 227 97 234
tri 97 227 99 234 sw
rect 66 226 99 227
rect 352 233 382 235
rect 352 227 380 233
tri 380 229 382 233 nw
tri 66 216 71 226 ne
rect 71 222 99 226
tri 269 224 287 226 se
rect 287 224 301 226
tri 301 224 312 226 sw
tri 351 224 352 226 se
rect 352 224 378 227
tri 99 222 100 224 sw
tri 263 222 268 224 se
rect 268 222 312 224
tri 312 222 316 224 sw
rect 71 216 100 222
rect 291 220 316 222
tri 71 212 72 216 ne
rect 72 212 100 216
tri 100 212 104 220 sw
tri 72 195 80 212 ne
rect 80 195 104 212
tri 104 195 111 212 sw
tri 80 187 83 195 ne
rect 83 189 111 195
tri 111 189 116 195 sw
rect 83 186 116 189
tri 116 186 120 189 sw
rect 312 186 316 220
tri 349 201 351 224 se
rect 351 201 378 224
tri 378 201 380 227 nw
rect 421 201 425 235
rect 459 201 490 235
tri 348 196 349 197 se
rect 349 196 378 201
rect 421 200 490 201
rect 421 199 460 200
tri 421 197 423 199 ne
rect 423 197 460 199
tri 460 197 463 200 nw
tri 463 197 490 200 ne
rect 348 191 378 196
tri 347 188 348 191 se
rect 348 188 377 191
tri 377 188 378 191 nw
rect 542 238 577 240
tri 676 245 678 248 se
rect 678 245 715 248
tri 715 245 718 248 sw
rect 676 244 718 245
tri 577 238 578 239 sw
rect 542 229 578 238
tri 578 229 580 237 sw
rect 542 219 580 229
tri 580 219 583 229 sw
tri 675 220 676 229 se
tri 675 219 676 220 ne
rect 542 210 583 219
tri 583 210 585 219 sw
rect 676 210 680 244
rect 714 240 718 244
rect 798 239 802 273
rect 836 244 869 273
rect 836 243 842 244
tri 842 243 847 244 nw
tri 847 243 851 244 ne
rect 851 243 869 244
rect 836 239 840 243
tri 840 240 842 243 nw
tri 851 240 866 243 ne
rect 866 240 869 243
tri 866 239 869 240 ne
rect 798 237 840 239
tri 798 235 800 237 ne
rect 800 235 838 237
tri 838 235 840 237 nw
rect 921 282 960 285
tri 960 282 965 286 nw
tri 1253 282 1258 286 ne
rect 1258 282 1264 286
rect 921 273 952 282
tri 952 274 960 282 nw
tri 1258 280 1260 282 ne
rect 921 271 950 273
tri 950 271 952 273 nw
rect 1260 273 1264 282
rect 1298 273 1302 307
tri 1339 291 1342 309 ne
rect 1342 291 1370 309
tri 1370 291 1372 309 sw
rect 1260 271 1302 273
rect 921 269 947 271
tri 947 269 950 271 nw
tri 1260 269 1262 271 ne
rect 1262 269 1300 271
tri 1300 269 1302 271 nw
rect 1342 286 1372 291
tri 1458 290 1521 309 se
rect 1521 308 1658 309
tri 1658 308 1663 309 nw
tri 1723 308 1726 309 ne
rect 1726 308 1783 309
rect 1521 301 1629 308
tri 1629 301 1658 308 nw
tri 1726 301 1739 308 ne
rect 1739 301 1783 308
rect 1521 290 1583 301
tri 1583 290 1629 301 nw
tri 1739 290 1759 301 ne
rect 1759 290 1783 301
tri 1422 288 1424 290 se
rect 1424 288 1573 290
tri 1573 288 1583 290 nw
tri 1759 288 1764 290 ne
rect 1764 288 1783 290
rect 1422 286 1555 288
tri 1342 269 1344 286 ne
rect 1344 269 1372 286
rect 921 252 931 269
tri 931 252 947 269 nw
tri 1344 260 1345 269 ne
rect 1345 260 1372 269
tri 1372 260 1375 286 sw
rect 1345 252 1375 260
rect 1422 252 1426 286
rect 1460 284 1555 286
tri 1555 284 1573 288 nw
tri 1764 284 1771 288 ne
rect 1771 284 1783 288
rect 1460 281 1545 284
tri 1545 281 1555 284 nw
rect 1460 277 1533 281
tri 1533 277 1545 281 nw
tri 1771 278 1783 284 ne
rect 1460 276 1529 277
tri 1529 276 1533 277 nw
rect 1460 273 1520 276
tri 1520 273 1529 276 nw
rect 1835 308 1837 312
tri 1837 308 1840 312 sw
rect 1835 301 1840 308
tri 1840 301 1842 308 sw
rect 1835 288 1842 301
rect 1835 281 1841 288
tri 1841 281 1842 288 nw
rect 1835 277 1839 281
tri 1839 277 1841 281 nw
rect 1835 275 1836 277
tri 1836 275 1839 277 nw
rect 1460 269 1504 273
tri 1504 269 1520 273 nw
rect 1460 268 1501 269
tri 1501 268 1504 269 nw
rect 1460 258 1467 268
tri 1467 258 1500 268 nw
tri 1835 274 1836 275 nw
rect 1460 252 1464 258
tri 921 242 931 252 nw
tri 1345 251 1346 252 ne
rect 1346 251 1375 252
tri 1375 251 1376 252 sw
rect 1422 251 1464 252
tri 1464 251 1467 258 nw
rect 1346 249 1376 251
tri 1376 249 1377 251 sw
tri 1422 249 1423 251 ne
rect 1423 249 1461 251
tri 1196 234 1197 235 se
tri 1037 233 1044 234 se
rect 1044 233 1088 234
tri 1031 232 1037 233 se
rect 1037 232 1088 233
tri 1088 232 1092 234 sw
tri 1029 231 1031 232 se
rect 1031 231 1092 232
tri 1092 231 1093 232 sw
rect 542 206 585 210
tri 585 206 586 210 sw
rect 676 208 684 210
tri 676 206 678 208 ne
rect 678 206 684 208
rect 542 200 586 206
tri 586 200 587 204 sw
rect 542 198 587 200
tri 587 198 588 200 sw
rect 542 195 588 198
tri 588 195 589 197 sw
rect 542 191 589 195
tri 589 191 590 195 sw
rect 542 188 590 191
tri 590 188 592 189 sw
tri 1028 228 1029 231 se
rect 1029 230 1093 231
tri 1093 230 1095 231 sw
rect 1029 228 1095 230
rect 1028 222 1095 228
rect 1028 213 1047 222
rect 1081 213 1095 222
rect 1028 210 1044 213
tri 1028 208 1029 210 ne
rect 1029 197 1044 210
tri 1029 195 1030 197 ne
tri 83 182 85 186 ne
rect 85 181 120 186
tri 120 181 128 186 sw
tri 85 178 87 181 ne
rect 87 178 128 181
tri 128 178 133 181 sw
tri 87 177 88 178 ne
rect 88 177 133 178
tri 133 177 135 178 sw
tri 88 174 89 177 ne
rect 89 174 135 177
tri 135 174 139 177 sw
tri 89 168 92 174 ne
rect 92 172 139 174
tri 139 172 143 174 sw
rect 92 170 143 172
tri 143 170 146 172 sw
rect 291 184 316 186
rect 291 182 314 184
tri 314 182 316 184 nw
tri 346 183 347 186 se
rect 347 183 377 188
tri 539 186 540 188 ne
rect 540 186 592 188
tri 592 186 597 188 sw
rect 1030 186 1044 197
rect 1196 196 1197 234
rect 1346 238 1377 249
rect 1424 248 1461 249
tri 1461 248 1464 251 nw
tri 1619 243 1620 244 sw
rect 1619 241 1620 243
tri 1620 241 1621 243 sw
tri 1377 238 1378 239 sw
rect 1346 218 1378 238
tri 1378 218 1380 234 sw
rect 1346 204 1380 218
rect 1619 238 1621 241
tri 1621 238 1623 241 sw
rect 1619 232 1623 238
tri 1623 232 1626 238 sw
rect 1619 217 1626 232
tri 1698 232 1700 235 se
rect 1700 232 1737 235
tri 1737 232 1740 235 sw
rect 1698 231 1740 232
tri 1626 217 1634 231 sw
rect 1619 209 1634 217
tri 1634 209 1639 217 sw
tri 1380 204 1381 205 sw
tri 1344 201 1346 203 se
rect 1346 201 1381 204
tri 1343 199 1344 201 se
rect 1344 200 1381 201
tri 1381 200 1382 201 sw
rect 1619 203 1639 209
tri 1639 203 1642 209 sw
rect 1619 201 1642 203
tri 1642 201 1644 203 sw
rect 1619 200 1644 201
rect 1344 199 1382 200
tri 1588 199 1590 200 ne
rect 1590 199 1644 200
tri 1196 195 1197 196 ne
tri 1341 197 1343 199 se
rect 1343 197 1382 199
tri 1340 195 1341 197 se
rect 1341 195 1382 197
tri 1336 189 1340 194 se
rect 1340 189 1382 195
rect 1336 188 1382 189
tri 1382 188 1383 194 sw
tri 1590 188 1601 199 ne
rect 1601 197 1644 199
tri 1644 197 1646 201 sw
rect 1698 197 1702 231
rect 1736 217 1740 231
tri 1740 217 1783 232 sw
rect 1736 209 1783 217
tri 1783 209 1804 217 sw
rect 1736 203 1804 209
tri 1804 203 1821 209 sw
rect 1736 201 1821 203
tri 1821 201 1827 203 sw
rect 1736 199 1827 201
tri 1827 199 1831 201 sw
rect 1736 197 1807 199
rect 1601 188 1646 197
tri 540 183 542 186 ne
rect 542 183 597 186
tri 597 183 605 186 sw
tri 1030 183 1031 186 ne
rect 1031 183 1044 186
rect 291 181 312 182
tri 312 181 314 182 nw
tri 345 181 346 182 se
rect 346 181 377 183
rect 291 180 302 181
tri 302 180 312 181 nw
tri 291 179 302 180 nw
tri 344 174 345 177 se
rect 345 174 377 181
rect 542 181 605 183
tri 605 181 609 183 sw
tri 542 180 543 181 ne
rect 543 180 609 181
tri 609 180 612 181 sw
tri 1031 180 1037 183 ne
rect 1037 180 1044 183
tri 543 178 544 180 ne
rect 544 178 612 180
rect 545 177 612 178
tri 612 177 619 180 sw
tri 545 175 546 177 ne
rect 546 175 619 177
tri 546 174 547 175 ne
rect 547 174 619 175
tri 343 170 344 172 se
rect 344 171 377 174
rect 344 170 376 171
rect 92 167 146 170
tri 146 167 150 170 sw
tri 92 161 96 167 ne
rect 96 161 150 167
tri 150 161 160 167 sw
tri 342 164 343 167 se
rect 343 164 376 170
tri 376 167 377 171 nw
tri 547 168 550 174 ne
rect 550 172 619 174
tri 619 172 634 177 sw
rect 550 167 634 172
tri 634 167 646 172 sw
tri 550 164 552 167 ne
rect 552 164 646 167
tri 336 162 339 164 se
rect 339 162 376 164
tri 376 162 378 164 sw
rect 96 160 160 161
tri 160 160 163 161 sw
rect 336 160 378 162
tri 96 157 99 160 ne
rect 99 157 163 160
tri 163 157 175 160 sw
tri 99 153 104 157 ne
rect 104 155 176 157
tri 176 155 179 157 sw
rect 104 153 179 155
tri 104 137 125 153 ne
rect 125 137 141 153
tri 125 136 127 137 ne
rect 127 136 141 137
tri 127 133 130 136 ne
rect 130 133 141 136
tri 131 130 132 133 ne
rect 132 128 141 133
tri 133 119 136 128 ne
rect 136 119 141 128
rect 175 119 179 153
rect 336 136 340 160
rect 374 136 378 160
tri 552 151 559 164 ne
rect 559 155 646 164
tri 646 155 676 167 sw
rect 559 153 690 155
tri 690 153 692 155 sw
rect 559 151 692 153
tri 559 146 562 151 ne
rect 562 146 654 151
tri 562 136 599 146 ne
rect 599 136 654 146
tri 136 117 137 119 ne
rect 137 117 179 119
tri 137 115 139 117 ne
rect 139 115 176 117
tri 176 115 179 117 nw
tri 599 134 605 136 ne
rect 605 134 654 136
tri 605 133 610 134 ne
rect 610 133 654 134
tri 610 129 626 133 ne
rect 626 129 654 133
tri 626 128 628 129 ne
rect 628 128 654 129
tri 631 126 637 128 ne
rect 637 126 654 128
tri 637 124 645 126 ne
rect 645 124 654 126
tri 645 122 646 124 ne
rect 646 122 654 124
tri 646 117 649 122 ne
rect 649 117 654 122
rect 688 117 692 151
tri 1037 178 1044 180 ne
tri 845 173 895 174 sw
rect 845 172 895 173
tri 895 172 899 173 sw
rect 845 171 899 172
tri 899 171 901 172 sw
rect 845 170 913 171
tri 913 170 914 171 sw
rect 845 168 914 170
tri 914 168 915 170 sw
rect 845 167 915 168
rect 845 136 877 167
tri 845 135 871 136 ne
rect 871 135 877 136
tri 871 133 873 135 ne
rect 873 133 877 135
rect 911 133 915 167
tri 1334 186 1336 188 se
rect 1336 186 1383 188
tri 1332 183 1334 186 se
rect 1334 185 1383 186
tri 1383 185 1386 188 sw
tri 1601 186 1604 188 ne
rect 1604 186 1646 188
rect 1334 183 1392 185
tri 1392 183 1393 185 sw
tri 1330 181 1332 183 se
rect 1332 182 1393 183
tri 1393 182 1394 183 sw
tri 1604 182 1608 186 ne
rect 1608 184 1646 186
tri 1646 184 1654 197 sw
rect 1698 195 1807 197
tri 1698 193 1700 195 ne
rect 1700 193 1807 195
tri 1711 190 1719 193 ne
rect 1719 190 1807 193
tri 1769 185 1780 190 ne
rect 1780 185 1807 190
tri 1780 184 1782 185 ne
rect 1782 184 1807 185
rect 1608 182 1654 184
tri 1654 182 1655 184 sw
tri 1782 182 1784 184 ne
rect 1784 182 1807 184
rect 1332 181 1394 182
tri 1329 178 1330 180 se
rect 1330 178 1356 181
tri 1328 177 1329 178 se
rect 1329 177 1356 178
tri 1326 174 1328 177 se
rect 1328 174 1356 177
tri 1325 172 1326 173 se
rect 1326 172 1356 174
tri 1321 170 1325 172 se
rect 1325 170 1356 172
tri 1318 168 1321 170 se
rect 1321 168 1356 170
tri 1302 162 1318 168 se
rect 1318 162 1356 168
tri 1297 161 1302 162 se
rect 1302 161 1356 162
tri 1290 158 1297 161 se
rect 1297 158 1356 161
tri 1285 157 1290 158 se
rect 1290 157 1356 158
tri 1276 154 1285 157 se
rect 1285 154 1356 157
tri 1271 152 1276 154 se
rect 1276 152 1356 154
tri 1255 147 1271 152 se
rect 1271 147 1356 152
rect 1390 155 1394 181
tri 1608 170 1621 182 ne
rect 1621 170 1655 182
tri 1507 168 1510 170 se
rect 1510 168 1547 170
tri 1547 168 1549 170 sw
rect 1507 166 1549 168
rect 1507 164 1511 166
tri 1394 155 1395 157 sw
rect 1390 147 1395 155
tri 1482 154 1484 155 se
tri 1239 142 1255 147 se
rect 1255 146 1395 147
rect 1255 143 1392 146
rect 1255 142 1332 143
tri 1332 142 1336 143 nw
tri 1336 142 1366 143 ne
rect 1366 142 1392 143
tri 1392 142 1395 146 nw
tri 1480 150 1482 154 se
rect 1482 150 1484 154
tri 1228 139 1239 142 se
rect 1239 139 1322 142
tri 1322 139 1330 142 nw
rect 1480 139 1484 150
rect 873 131 915 133
tri 1085 132 1228 139 se
rect 1228 132 1300 139
tri 1300 132 1322 139 nw
tri 1480 133 1481 139 ne
tri 873 129 875 131 ne
rect 875 129 913 131
tri 913 129 915 131 nw
tri 649 116 650 117 ne
rect 650 116 692 117
rect 650 115 690 116
tri 650 113 652 115 ne
rect 652 113 690 115
tri 690 113 692 116 nw
tri 1052 130 1061 132 se
rect 1061 130 1295 132
tri 1295 130 1300 132 nw
rect 1481 130 1484 139
rect 1545 134 1549 166
tri 1621 153 1640 170 ne
rect 1640 156 1655 170
tri 1655 156 1689 182 sw
tri 1784 164 1807 182 ne
rect 1640 155 1689 156
tri 1689 155 1691 156 sw
rect 1640 153 1691 155
tri 1640 150 1643 153 ne
rect 1643 150 1691 153
tri 1691 150 1731 155 sw
tri 1643 144 1653 150 ne
rect 1653 147 1731 150
tri 1731 147 1756 150 sw
rect 1653 144 1767 147
tri 1767 144 1769 147 sw
tri 1653 143 1654 144 ne
rect 1654 143 1769 144
tri 1549 134 1552 143 sw
rect 1545 132 1552 134
rect 1045 128 1289 130
tri 1289 128 1295 130 nw
tri 1481 129 1482 130 ne
rect 1045 94 1062 128
rect 1096 125 1279 128
tri 1279 125 1287 128 nw
rect 1096 123 1272 125
tri 1272 123 1279 125 nw
rect 1482 123 1484 130
rect 1096 120 1265 123
tri 1265 120 1272 123 nw
tri 1482 120 1483 123 ne
rect 1483 120 1484 123
rect 1096 119 1260 120
tri 1260 119 1265 120 nw
tri 1483 119 1484 120 ne
rect 1096 117 1254 119
tri 1254 117 1260 119 nw
rect 1096 115 1249 117
tri 1249 115 1254 117 nw
rect 1096 114 1246 115
tri 1246 114 1249 115 nw
rect 1096 113 1241 114
tri 1241 113 1246 114 nw
rect 1096 111 1235 113
tri 1235 111 1241 113 nw
rect 1536 126 1552 132
tri 1654 129 1678 143 ne
rect 1678 129 1731 143
tri 1678 127 1684 129 ne
rect 1684 127 1731 129
tri 1684 126 1688 127 ne
rect 1688 126 1731 127
rect 1536 123 1549 126
tri 1549 123 1552 126 nw
tri 1688 123 1696 126 ne
rect 1696 123 1731 126
tri 1536 122 1549 123 nw
tri 1696 121 1706 123 ne
rect 1706 121 1731 123
tri 1706 120 1707 121 ne
rect 1707 120 1731 121
tri 1707 119 1710 120 ne
rect 1710 119 1731 120
tri 1713 117 1718 119 ne
rect 1718 117 1731 119
tri 1719 115 1725 117 ne
rect 1725 115 1731 117
tri 1725 113 1727 115 ne
rect 1096 109 1216 111
tri 1216 109 1235 111 nw
rect 1727 109 1731 115
rect 1765 109 1769 143
rect 1096 105 1179 109
tri 1179 105 1216 109 nw
rect 1727 107 1769 109
tri 1727 105 1730 107 ne
rect 1730 105 1767 107
tri 1767 105 1769 107 nw
rect 1096 96 1102 105
tri 1102 96 1179 105 nw
rect 1096 94 1100 96
rect 1045 92 1100 94
tri 1100 92 1102 96 nw
rect 1045 90 1098 92
tri 1098 90 1100 92 nw
rect 1045 89 1052 90
tri 1052 89 1061 90 nw
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< via1 >>
rect 295 361 347 413
rect 39 337 91 346
rect 39 303 61 337
rect 61 303 91 337
rect 39 294 91 303
rect 248 334 300 344
rect 652 350 666 384
rect 666 350 700 384
rect 700 350 704 384
rect 790 372 809 387
rect 809 372 842 387
rect 248 300 286 334
rect 286 300 300 334
rect 248 292 300 300
rect 652 332 704 350
rect 790 335 842 372
rect 1500 344 1552 396
rect 1783 309 1835 313
rect 239 220 291 222
rect 239 186 278 220
rect 278 186 291 220
rect 490 188 542 240
rect 684 210 714 240
rect 714 210 736 240
rect 869 233 921 285
rect 1783 275 1795 309
rect 1795 275 1829 309
rect 1829 275 1835 309
rect 1783 261 1835 275
rect 684 188 736 210
rect 239 170 291 186
rect 1044 188 1047 213
rect 1047 188 1081 213
rect 1081 188 1096 213
rect 1197 232 1249 243
rect 1197 198 1200 232
rect 1200 198 1234 232
rect 1234 198 1249 232
rect 1567 239 1619 252
rect 1567 205 1580 239
rect 1580 205 1614 239
rect 1614 205 1619 239
rect 1567 200 1619 205
rect 1197 191 1249 198
rect 327 126 340 136
rect 340 126 374 136
rect 374 126 379 136
rect 327 84 379 126
rect 793 127 845 179
rect 1044 161 1096 188
rect 993 80 1045 132
rect 1484 132 1511 164
rect 1511 132 1536 164
rect 1807 147 1859 199
rect 1484 112 1536 132
<< metal2 >>
tri 1329 475 1451 480 se
tri 1451 478 1472 480 sw
rect 1451 475 1472 478
tri 270 464 371 475 se
rect 371 474 557 475
tri 557 474 821 475 sw
tri 1301 474 1318 475 se
rect 1318 474 1472 475
rect 371 464 821 474
tri 821 464 876 474 sw
tri 1131 468 1301 474 se
rect 1301 468 1472 474
tri 255 462 270 464 se
rect 270 462 876 464
tri 876 462 878 464 sw
tri 249 460 255 462 se
rect 255 460 878 462
tri 878 460 883 462 sw
tri 245 455 249 460 se
rect 249 455 883 460
tri 883 455 890 460 sw
rect 245 448 890 455
tri 890 448 902 455 sw
rect 245 447 902 448
tri 902 447 903 448 sw
tri 244 446 245 447 se
rect 245 446 371 447
tri 371 446 381 447 nw
tri 381 446 725 447 ne
rect 725 446 903 447
rect 244 444 351 446
tri 351 444 369 446 nw
tri 811 444 824 446 ne
rect 824 444 903 446
tri 903 444 906 446 sw
rect 244 435 295 444
tri 295 435 351 444 nw
tri 824 435 834 444 ne
rect 834 435 906 444
rect 244 434 286 435
tri 286 434 295 435 nw
tri 834 434 835 435 ne
rect 835 434 906 435
rect 244 432 282 434
tri 282 432 286 434 nw
tri 835 432 838 434 ne
rect 838 432 906 434
tri 243 421 244 431 se
rect 244 421 274 432
tri 274 421 282 432 nw
tri 838 421 851 432 ne
rect 851 421 906 432
tri 242 413 243 421 se
rect 243 413 273 421
tri 273 418 274 421 nw
tri 851 413 859 421 ne
rect 859 418 906 421
tri 906 418 927 444 sw
rect 859 416 927 418
tri 927 416 929 418 sw
rect 859 413 929 416
tri 241 393 242 396 se
rect 242 393 272 413
tri 272 410 273 413 nw
tri 240 373 241 392 se
tri 240 367 241 373 ne
rect 241 370 272 393
tri 272 370 273 392 sw
rect 241 358 273 370
tri 859 410 863 413 ne
rect 863 410 929 413
tri 929 410 934 416 sw
tri 1035 465 1131 468 se
rect 1131 465 1472 468
rect 1035 464 1472 465
tri 1472 464 1580 478 sw
rect 1035 462 1580 464
tri 1580 462 1598 464 sw
rect 1035 461 1598 462
tri 1598 461 1599 462 sw
rect 1035 458 1599 461
tri 1599 458 1606 461 sw
rect 1035 454 1606 458
tri 1606 454 1612 458 sw
rect 1035 449 1612 454
tri 1612 449 1615 454 sw
rect 1035 437 1327 449
tri 1327 437 1452 449 nw
tri 1468 437 1569 449 ne
rect 1569 437 1615 449
rect 1035 431 1269 437
tri 1269 431 1327 437 nw
tri 1569 431 1576 437 ne
rect 1576 431 1615 437
tri 1615 431 1624 449 sw
rect 1035 428 1234 431
tri 1234 428 1269 431 nw
tri 1576 428 1578 431 ne
rect 1578 428 1624 431
rect 1035 422 1047 428
tri 1047 422 1234 428 nw
tri 1035 419 1047 422 nw
tri 1578 420 1582 428 ne
rect 1582 419 1624 428
tri 1582 418 1583 419 ne
rect 1583 418 1624 419
tri 1583 416 1584 418 ne
rect 1584 416 1624 418
tri 1584 411 1586 416 ne
rect 1586 414 1624 416
tri 1624 414 1632 431 sw
rect 1586 410 1632 414
tri 863 406 868 410 ne
rect 868 406 934 410
tri 934 406 937 410 sw
tri 1586 406 1589 410 ne
rect 1589 406 1632 410
tri 868 404 870 406 ne
rect 870 404 937 406
tri 870 401 874 404 ne
rect 874 401 937 404
tri 874 399 876 401 ne
rect 876 399 937 401
tri 937 399 944 406 sw
tri 1589 404 1590 406 ne
rect 1590 404 1632 406
tri 1632 404 1633 414 sw
tri 1590 401 1591 404 ne
rect 1591 401 1632 404
tri 1591 399 1592 401 ne
rect 1592 399 1632 401
rect 347 396 348 399
tri 348 396 367 399 sw
tri 876 396 880 399 ne
rect 880 396 944 399
tri 944 396 946 399 sw
tri 1592 396 1594 399 ne
rect 1594 396 1632 399
rect 347 387 367 396
tri 367 387 429 396 sw
tri 880 387 890 396 ne
rect 890 387 946 396
rect 347 384 429 387
tri 429 384 449 387 sw
rect 347 375 449 384
tri 449 375 512 384 sw
tri 605 377 648 379 se
rect 648 377 652 379
tri 551 375 605 377 se
rect 605 375 652 377
rect 347 374 512 375
tri 512 374 529 375 sw
tri 529 374 551 375 se
rect 551 374 652 375
rect 347 362 652 374
tri 347 358 359 362 ne
rect 359 358 652 362
tri 48 352 49 353 se
rect 49 352 55 353
tri 45 348 48 352 se
rect 48 348 55 352
rect 45 346 55 348
tri 241 355 242 358 ne
rect 242 354 273 358
tri 273 354 276 358 sw
tri 359 354 369 358 ne
rect 369 354 652 358
rect 242 350 276 354
tri 276 350 282 354 sw
tri 369 350 381 354 ne
rect 381 350 652 354
tri 242 346 243 350 ne
rect 243 345 282 350
tri 282 345 286 350 sw
tri 381 345 398 350 ne
rect 398 345 652 350
rect 243 344 286 345
tri 398 344 402 345 ne
rect 402 344 652 345
tri 243 338 244 344 ne
rect 244 333 248 344
tri 244 305 247 333 ne
rect 247 301 248 333
tri 247 300 248 301 ne
rect 91 298 103 300
tri 103 299 104 300 nw
rect 91 296 102 298
tri 102 297 103 298 nw
rect 91 294 100 296
tri 46 293 47 294 ne
rect 47 293 100 294
tri 100 293 102 296 nw
tri 47 291 95 293 ne
rect 95 292 98 293
tri 98 292 100 293 nw
tri 402 341 421 344 ne
rect 421 341 652 344
tri 421 337 590 341 ne
rect 590 337 652 341
tri 590 336 652 337 ne
tri 788 374 790 375 se
tri 784 366 788 374 se
rect 788 366 790 374
tri 784 341 786 366 ne
rect 786 339 790 366
tri 786 337 787 339 ne
rect 787 335 790 339
tri 890 383 895 387 ne
rect 895 383 946 387
tri 946 383 958 396 sw
tri 895 379 899 383 ne
rect 899 380 958 383
tri 958 380 959 383 sw
rect 899 379 959 380
tri 959 379 960 380 sw
tri 900 351 932 379 ne
rect 932 372 960 379
tri 960 372 966 379 sw
rect 932 368 966 372
tri 966 368 970 372 sw
tri 1499 368 1500 370 se
rect 932 361 970 368
tri 970 361 978 368 sw
tri 1498 363 1499 368 se
rect 1499 363 1500 368
rect 932 359 978 361
tri 978 359 985 361 sw
rect 932 355 985 359
tri 985 355 1001 359 sw
rect 932 352 1001 355
tri 1001 352 1367 355 sw
rect 932 351 1367 352
tri 932 350 934 351 ne
rect 934 350 1367 351
tri 934 344 942 350 ne
rect 942 344 1367 350
tri 942 340 948 344 ne
rect 948 340 1367 344
tri 948 335 959 340 ne
rect 959 335 1367 340
rect 787 333 830 335
rect 787 332 827 333
tri 787 324 788 332 ne
rect 788 313 827 332
tri 827 313 830 333 nw
tri 959 321 990 335 ne
rect 990 321 1367 335
tri 990 317 1008 321 ne
rect 1008 317 1367 321
tri 1008 313 1100 317 ne
rect 1100 313 1367 317
tri 788 300 790 313 ne
rect 790 311 827 313
tri 95 291 98 292 nw
rect 790 285 823 311
tri 823 285 827 311 nw
tri 1100 304 1308 313 ne
rect 1308 304 1367 313
tri 1308 303 1318 304 ne
rect 1318 303 1367 304
tri 1318 297 1351 303 ne
rect 1351 300 1367 303
tri 1494 355 1498 363 se
rect 1498 355 1500 363
tri 1493 352 1494 355 se
rect 1494 352 1500 355
tri 1492 350 1493 351 se
rect 1493 350 1500 352
tri 1423 342 1432 348 sw
tri 1491 347 1492 348 se
rect 1492 347 1500 350
tri 1487 344 1491 347 se
rect 1491 344 1500 347
tri 1594 389 1597 396 ne
rect 1597 389 1632 396
tri 1597 383 1600 389 ne
rect 1600 383 1632 389
tri 1632 384 1633 404 nw
tri 1600 380 1601 383 ne
rect 1601 379 1630 383
tri 1601 372 1602 379 ne
tri 1598 352 1602 372 se
rect 1602 352 1630 379
tri 1630 352 1632 383 nw
rect 1598 350 1630 352
tri 1597 344 1598 347 se
rect 1598 344 1628 350
tri 1486 343 1487 344 se
rect 1487 343 1535 344
tri 1474 342 1486 343 se
rect 1486 342 1535 343
tri 1535 342 1537 344 nw
rect 1423 340 1432 342
tri 1432 340 1436 342 sw
tri 1454 341 1474 342 se
rect 1474 341 1534 342
tri 1448 340 1454 341 se
rect 1454 340 1534 341
tri 1534 340 1535 342 nw
tri 1596 340 1597 342 se
rect 1597 340 1628 344
rect 1423 321 1518 340
tri 1518 321 1533 340 nw
tri 1593 321 1596 339 se
rect 1596 321 1628 340
rect 1423 317 1514 321
tri 1514 317 1518 321 nw
tri 1592 317 1593 321 se
rect 1593 317 1628 321
tri 1628 319 1630 350 nw
rect 1423 313 1511 317
tri 1511 313 1514 317 nw
rect 1592 313 1628 317
rect 1423 303 1503 313
tri 1503 304 1511 313 nw
tri 1590 304 1592 313 se
rect 1592 304 1627 313
tri 1627 304 1628 313 nw
tri 1839 347 1840 348 sw
rect 1839 314 1840 347
tri 1840 314 1841 340 sw
rect 1590 303 1627 304
rect 1423 300 1499 303
rect 1351 297 1499 300
tri 1499 298 1503 303 nw
tri 1589 298 1590 303 se
rect 1590 298 1625 303
rect 1589 297 1625 298
tri 1351 296 1357 297 ne
rect 1357 296 1375 297
tri 1357 295 1375 296 ne
tri 1375 295 1397 297 nw
tri 1418 295 1427 297 ne
rect 1427 295 1496 297
tri 1427 288 1458 295 ne
rect 1458 288 1496 295
tri 1496 290 1498 297 nw
tri 1587 290 1588 296 se
rect 1588 290 1625 297
tri 1496 288 1497 290 sw
tri 1458 285 1461 288 ne
rect 1461 285 1497 288
tri 790 269 792 285 ne
rect 792 282 823 285
rect 792 268 821 282
tri 518 262 572 268 se
tri 572 263 584 268 sw
tri 792 264 793 268 ne
rect 572 262 584 263
tri 509 255 518 262 se
rect 518 255 584 262
tri 584 255 588 262 sw
rect 793 255 821 268
tri 821 267 823 282 nw
tri 501 240 509 255 se
rect 509 244 588 255
tri 588 244 592 255 sw
tri 793 247 794 255 ne
rect 794 244 821 255
rect 509 240 543 244
tri 291 198 354 213 sw
rect 291 197 354 198
tri 354 197 356 198 sw
rect 291 192 356 197
tri 356 192 377 197 sw
rect 291 188 377 192
tri 377 188 393 192 sw
rect 542 194 543 240
tri 794 240 795 244 ne
rect 795 236 821 244
tri 821 236 825 267 sw
rect 795 233 825 236
tri 1461 284 1463 285 ne
rect 1463 279 1497 285
tri 1586 284 1587 288 se
rect 1587 284 1625 290
tri 1497 279 1498 284 sw
rect 1463 278 1498 279
rect 1464 277 1498 278
tri 1585 278 1586 284 se
rect 1586 278 1625 284
tri 1464 268 1465 277 ne
rect 1465 268 1498 277
tri 1498 268 1499 277 sw
rect 1465 267 1499 268
tri 1583 268 1585 277 se
rect 1585 268 1625 278
tri 1625 270 1627 303 nw
rect 1839 300 1841 314
rect 1466 261 1499 267
tri 1582 262 1583 267 se
rect 1583 262 1623 268
rect 1582 261 1623 262
tri 1623 261 1625 268 nw
rect 1835 297 1841 300
tri 1841 297 1842 304 sw
rect 1835 291 1840 297
tri 1840 291 1842 297 nw
tri 1835 287 1840 291 nw
tri 1466 258 1467 261 ne
tri 921 253 925 258 sw
rect 921 246 925 253
rect 1467 257 1499 261
tri 1499 257 1500 261 sw
tri 1581 257 1582 261 se
rect 1582 257 1622 261
tri 1622 257 1623 261 nw
tri 1467 252 1468 257 ne
rect 1468 252 1500 257
tri 1500 252 1501 257 sw
tri 1579 253 1581 257 se
rect 1581 253 1620 257
rect 1579 252 1620 253
tri 925 246 930 252 sw
rect 1468 251 1501 252
tri 1468 249 1469 251 ne
rect 921 244 930 246
tri 930 244 931 246 sw
tri 795 216 797 233 ne
rect 797 213 825 233
tri 825 213 828 233 sw
tri 797 192 799 213 ne
rect 291 182 393 188
tri 393 182 418 188 sw
rect 799 183 828 213
tri 828 183 832 213 sw
tri 1053 213 1055 220 se
rect 1469 243 1501 251
tri 1469 242 1470 243 ne
rect 1470 240 1501 243
tri 1470 237 1471 240 ne
rect 1471 237 1501 240
tri 1501 237 1502 246 sw
rect 1471 234 1502 237
tri 1471 230 1472 234 ne
rect 1472 230 1502 234
tri 1502 230 1503 236 sw
rect 1472 226 1503 230
rect 1249 200 1251 226
tri 1251 200 1312 226 sw
tri 1472 208 1476 226 ne
rect 1476 220 1503 226
tri 1503 220 1504 229 sw
rect 1476 207 1504 220
tri 1504 207 1509 220 sw
tri 1476 201 1477 207 ne
rect 1477 200 1509 207
tri 1509 200 1511 207 sw
rect 1619 251 1620 252
tri 1620 251 1622 257 nw
tri 1619 249 1620 251 nw
rect 1249 199 1312 200
tri 1312 199 1314 200 sw
rect 1477 199 1511 200
rect 1249 198 1314 199
tri 1314 198 1317 199 sw
tri 1477 198 1478 199 ne
rect 1478 198 1511 199
tri 1511 198 1512 199 sw
rect 1249 197 1317 198
tri 1317 197 1318 198 sw
rect 1478 197 1512 198
rect 1249 191 1318 197
tri 1318 191 1333 197 sw
tri 1478 192 1479 197 ne
rect 1479 191 1512 197
tri 1512 191 1515 197 sw
tri 1244 188 1252 191 ne
rect 1252 188 1333 191
rect 799 182 832 183
rect 291 179 418 182
tri 418 179 422 182 sw
tri 799 180 800 182 ne
rect 800 179 832 182
tri 303 178 305 179 ne
rect 305 178 422 179
tri 305 177 311 178 ne
rect 311 177 422 178
tri 311 170 337 177 ne
rect 337 170 422 177
tri 337 160 376 170 ne
rect 376 166 422 170
tri 422 166 439 179 sw
rect 376 160 439 166
tri 439 160 443 166 sw
tri 376 158 388 160 ne
rect 388 158 443 160
tri 388 156 403 158 ne
rect 403 156 443 158
tri 443 156 447 160 sw
tri 403 154 408 156 ne
rect 408 154 447 156
tri 447 154 448 156 sw
tri 408 149 415 154 ne
rect 415 149 448 154
tri 448 149 452 154 sw
tri 415 142 418 149 ne
rect 418 142 452 149
tri 452 142 458 149 sw
tri 418 137 421 142 ne
rect 421 137 458 142
tri 458 137 461 142 sw
rect 421 136 461 137
tri 421 130 426 136 ne
rect 426 130 461 136
tri 461 130 467 137 sw
tri 426 128 428 130 ne
rect 428 127 467 130
tri 467 127 469 130 sw
rect 1096 180 1106 188
tri 1106 180 1107 188 nw
tri 1252 180 1275 188 ne
rect 1275 186 1333 188
tri 1333 186 1346 191 sw
tri 1479 187 1480 191 ne
rect 1275 182 1346 186
tri 1346 182 1354 186 sw
rect 1480 185 1515 191
tri 1480 182 1481 185 ne
rect 1481 182 1515 185
tri 1515 182 1518 191 sw
rect 1275 180 1354 182
rect 1096 176 1104 180
tri 1104 176 1106 180 nw
tri 1275 176 1286 180 ne
rect 1286 176 1354 180
rect 1096 175 1103 176
tri 1103 175 1104 176 nw
tri 1096 172 1103 175 nw
tri 1286 172 1298 176 ne
rect 1298 172 1354 176
tri 1298 170 1305 172 ne
rect 1305 170 1354 172
tri 1305 168 1311 170 ne
rect 1311 168 1354 170
tri 1311 164 1322 168 ne
rect 1322 164 1354 168
tri 1354 164 1375 182 sw
tri 1481 174 1482 182 ne
rect 1482 174 1518 182
tri 1518 174 1521 182 sw
tri 1482 170 1483 174 ne
rect 1483 170 1521 174
tri 1521 170 1523 174 sw
tri 1684 170 1687 174 se
tri 1483 165 1484 170 ne
rect 1484 166 1523 170
tri 1523 166 1524 170 sw
rect 1484 164 1524 166
tri 1677 164 1684 170 se
rect 1684 164 1687 170
tri 1322 161 1330 164 ne
rect 1330 161 1375 164
tri 1330 160 1333 161 ne
rect 1333 160 1375 161
tri 1375 160 1380 164 sw
tri 1333 157 1339 160 ne
rect 1339 157 1380 160
tri 1380 157 1384 160 sw
tri 1339 141 1357 157 ne
rect 1357 141 1384 157
tri 1357 139 1359 141 ne
rect 1359 139 1384 141
tri 1359 134 1365 139 ne
rect 1365 134 1384 139
tri 1365 132 1367 134 ne
rect 1367 132 1384 134
tri 428 126 429 127 ne
rect 429 126 469 127
tri 429 113 441 126 ne
rect 441 113 469 126
tri 469 113 481 127 sw
tri 941 113 991 124 se
rect 991 113 993 124
tri 441 84 466 113 ne
rect 466 107 481 113
tri 481 107 488 113 sw
tri 918 107 941 113 se
rect 941 107 993 113
rect 466 105 488 107
tri 488 105 694 107 sw
tri 907 105 918 107 se
rect 918 105 993 107
rect 466 93 694 105
tri 694 93 853 105 sw
tri 865 95 907 105 se
rect 907 95 993 105
tri 853 93 865 95 se
rect 865 93 993 95
rect 466 85 993 93
rect 466 84 976 85
tri 466 83 467 84 ne
rect 467 83 976 84
tri 976 83 990 85 nw
tri 467 80 471 83 ne
rect 471 80 959 83
tri 959 80 976 83 nw
tri 1367 130 1370 132 ne
rect 1370 130 1384 132
tri 1371 125 1376 130 ne
rect 1376 125 1384 130
tri 1376 119 1383 125 ne
rect 1383 119 1384 125
tri 1384 119 1428 157 sw
tri 1383 112 1391 119 ne
rect 1391 112 1428 119
tri 1428 112 1436 119 sw
tri 1672 160 1677 164 se
rect 1677 160 1687 164
tri 1667 157 1672 160 se
rect 1672 157 1687 160
tri 1666 156 1667 157 se
rect 1667 156 1687 157
tri 1654 147 1666 156 se
rect 1666 155 1687 156
tri 1743 205 1746 206 sw
rect 1743 204 1746 205
tri 1746 204 1747 205 sw
rect 1743 200 1747 204
tri 1747 200 1750 204 sw
rect 1743 197 1750 200
tri 1750 197 1753 200 sw
rect 1743 194 1753 197
tri 1753 194 1759 197 sw
rect 1743 192 1759 194
tri 1759 192 1807 194 sw
rect 1743 155 1807 192
rect 1666 148 1807 155
rect 1666 147 1764 148
tri 1764 147 1770 148 nw
tri 1770 147 1779 148 ne
rect 1779 147 1807 148
tri 1629 128 1654 147 se
rect 1654 145 1751 147
tri 1751 145 1764 147 nw
tri 1779 145 1799 147 ne
rect 1799 145 1810 147
tri 1810 145 1826 147 nw
rect 1654 139 1703 145
tri 1703 139 1749 145 nw
rect 1654 135 1695 139
tri 1695 135 1703 139 nw
rect 1654 128 1686 135
tri 1686 128 1695 135 nw
tri 1611 119 1629 128 se
rect 1629 127 1684 128
tri 1684 127 1686 128 nw
rect 1629 124 1681 127
tri 1681 124 1684 127 nw
rect 1629 119 1674 124
tri 1609 118 1610 119 se
rect 1610 118 1674 119
tri 1674 118 1681 124 nw
tri 1594 112 1609 118 se
rect 1609 112 1665 118
tri 1391 87 1421 112 ne
rect 1421 104 1436 112
tri 1436 104 1446 112 sw
tri 1574 104 1594 112 se
rect 1594 110 1665 112
tri 1665 110 1674 118 nw
rect 1594 104 1609 110
rect 1421 88 1446 104
tri 1446 88 1490 104 sw
tri 1535 88 1574 104 se
rect 1574 88 1609 104
rect 1421 87 1490 88
tri 1490 87 1527 88 sw
rect 1535 87 1609 88
tri 1609 87 1665 110 nw
tri 1421 83 1426 87 ne
rect 1426 83 1595 87
tri 1426 82 1428 83 ne
rect 1428 82 1595 83
tri 1595 82 1607 87 nw
tri 1428 80 1430 82 ne
rect 1430 80 1586 82
tri 471 77 476 80 ne
rect 476 77 941 80
tri 941 77 959 80 nw
tri 1430 78 1433 80 ne
rect 1433 78 1586 80
tri 1586 78 1595 82 nw
tri 1433 77 1435 78 ne
rect 1435 77 1544 78
tri 476 72 520 77 ne
rect 520 74 922 77
tri 922 74 941 77 nw
tri 1435 74 1442 77 ne
rect 1442 74 1544 77
rect 520 72 907 74
tri 907 72 922 74 nw
tri 1442 72 1448 74 ne
rect 1448 72 1544 74
tri 520 69 540 72 ne
rect 540 71 711 72
tri 711 71 736 72 nw
tri 736 71 751 72 ne
rect 751 71 905 72
tri 905 71 907 72 nw
tri 1448 71 1449 72 ne
rect 1449 71 1544 72
rect 540 69 550 71
tri 550 69 711 71 nw
tri 751 69 780 71 ne
rect 780 69 851 71
tri 780 63 841 69 ne
rect 841 63 851 69
tri 851 63 901 71 nw
tri 1451 63 1469 71 ne
rect 1469 63 1544 71
tri 1469 60 1477 63 ne
rect 1477 61 1544 63
tri 1544 61 1586 78 nw
rect 1477 60 1541 61
tri 1541 60 1544 61 nw
tri 1477 59 1486 60 ne
rect 1486 59 1535 60
tri 1535 59 1541 60 nw
<< via2 >>
rect 979 412 1035 468
rect 55 346 111 356
rect 55 300 91 346
rect 91 300 111 346
rect 1367 300 1423 356
rect 1783 313 1839 356
rect 543 188 599 244
rect 687 240 743 244
rect 687 188 736 240
rect 736 188 743 240
rect 1783 300 1835 313
rect 1835 300 1839 313
rect 879 233 921 244
rect 921 233 935 244
rect 879 188 935 233
rect 1055 213 1111 244
rect 1055 188 1096 213
rect 1096 188 1111 213
rect 343 84 379 132
rect 379 84 399 132
rect 343 76 399 84
rect 1687 155 1743 211
<< metal3 >>
rect 974 470 1040 473
rect 733 468 1040 470
rect 733 412 979 468
rect 1035 412 1040 468
rect 733 410 1040 412
rect 50 356 116 361
rect 50 300 55 356
rect 111 300 116 356
rect 50 215 116 300
rect 538 244 604 329
rect 733 249 793 410
rect 974 407 1040 410
rect 1362 356 1428 361
rect 1362 300 1367 356
rect 1423 300 1428 356
rect 338 132 404 217
rect 538 188 543 244
rect 599 188 604 244
rect 538 183 604 188
rect 682 244 793 249
rect 682 188 687 244
rect 743 188 793 244
rect 682 186 793 188
rect 874 244 940 249
rect 874 188 879 244
rect 935 188 940 244
rect 682 183 748 186
rect 338 76 343 132
rect 399 76 404 132
rect 874 103 940 188
rect 1050 244 1116 249
rect 1050 188 1055 244
rect 1111 188 1116 244
rect 1362 215 1428 300
rect 1778 356 1844 441
rect 1778 300 1783 356
rect 1839 300 1844 356
rect 1778 295 1844 300
rect 1050 103 1116 188
rect 1682 211 1748 216
rect 1682 177 1687 211
rect 1674 155 1687 177
rect 1743 155 1748 211
rect 338 71 404 76
rect 1674 70 1748 155
rect 1674 47 1710 70
<< labels >>
flabel nwell s 33 527 67 561 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 521 527 555 561 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 1009 527 1043 561 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 1497 527 1531 561 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel pwell s 33 -17 67 17 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 521 -17 555 17 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 1009 -17 1043 17 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 1497 -17 1531 17 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel comment s 3 -8 3 -8 0 FreeSans 100 0 0 0 scs130hd_mpr2ea_8
flabel metal3 s 338 71 404 217 0 FreeSans 100 0 0 0 R1
port 3 nsew
flabel metal3 s 1050 103 1116 249 0 FreeSans 100 0 0 0 B1
port 4 nsew
flabel metal3 s 538 183 604 329 0 FreeSans 100 0 0 0 R3
port 5 nsew
flabel metal3 s 1362 215 1428 361 0 FreeSans 100 0 0 0 R0
port 6 nsew
flabel metal3 s 1682 70 1748 216 0 FreeSans 100 0 0 0 A0
port 7 nsew
flabel metal3 s 50 215 116 361 0 FreeSans 100 0 0 0 R2
port 8 nsew
flabel metal3 s 874 103 940 249 0 FreeSans 100 0 0 0 A1
port 9 nsew
flabel metal3 s 1778 295 1844 441 0 FreeSans 100 0 0 0 B0
port 10 nsew
flabel metal1 s 31 -17 65 17 0 FreeSans 100 0 0 0 vgnd
port 11 nsew
flabel metal1 s 31 527 65 561 0 FreeSans 100 0 0 0 vpwr
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 1932 544
<< end >>
