magic
tech sky130A
magscale 1 2
timestamp 1701356954
<< obsli1 >>
rect 1104 2159 8832 19601
<< obsm1 >>
rect 934 2128 8992 19632
<< metal2 >>
rect 1214 21200 1270 22000
rect 3698 21200 3754 22000
rect 6182 21200 6238 22000
rect 8666 21200 8722 22000
<< obsm2 >>
rect 938 21144 1158 21298
rect 1326 21144 3642 21298
rect 3810 21144 6126 21298
rect 6294 21144 8610 21298
rect 8778 21144 8986 21298
rect 938 711 8986 21144
<< metal3 >>
rect 0 20952 800 21072
rect 0 19592 800 19712
rect 0 18232 800 18352
rect 0 16872 800 16992
rect 0 15512 800 15632
rect 0 14152 800 14272
rect 0 12792 800 12912
rect 0 11432 800 11552
rect 9200 10888 10000 11008
rect 0 10072 800 10192
rect 0 8712 800 8832
rect 0 7352 800 7472
rect 0 5992 800 6112
rect 0 4632 800 4752
rect 0 3272 800 3392
rect 0 1912 800 2032
rect 0 552 800 672
<< obsm3 >>
rect 880 20872 9200 21045
rect 800 19792 9200 20872
rect 880 19512 9200 19792
rect 800 18432 9200 19512
rect 880 18152 9200 18432
rect 800 17072 9200 18152
rect 880 16792 9200 17072
rect 800 15712 9200 16792
rect 880 15432 9200 15712
rect 800 14352 9200 15432
rect 880 14072 9200 14352
rect 800 12992 9200 14072
rect 880 12712 9200 12992
rect 800 11632 9200 12712
rect 880 11352 9200 11632
rect 800 11088 9200 11352
rect 800 10808 9120 11088
rect 800 10272 9200 10808
rect 880 9992 9200 10272
rect 800 8912 9200 9992
rect 880 8632 9200 8912
rect 800 7552 9200 8632
rect 880 7272 9200 7552
rect 800 6192 9200 7272
rect 880 5912 9200 6192
rect 800 4832 9200 5912
rect 880 4552 9200 4832
rect 800 3472 9200 4552
rect 880 3192 9200 3472
rect 800 2112 9200 3192
rect 880 1832 9200 2112
rect 800 752 9200 1832
rect 880 582 9200 752
<< metal4 >>
rect 1910 2128 2230 19632
rect 2876 2128 3196 19632
rect 3842 2128 4162 19632
rect 4808 2128 5128 19632
rect 5774 2128 6094 19632
rect 6740 2128 7060 19632
rect 7706 2128 8026 19632
rect 8672 2128 8992 19632
<< labels >>
rlabel metal3 s 0 20952 800 21072 6 data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 data_in[11]
port 3 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 data_in[12]
port 4 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 data_in[13]
port 5 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 data_in[14]
port 6 nsew signal input
rlabel metal3 s 0 552 800 672 6 data_in[15]
port 7 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 data_in[1]
port 8 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 data_in[2]
port 9 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 data_in[3]
port 10 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 data_in[4]
port 11 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 data_in[5]
port 12 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 data_in[6]
port 13 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 data_in[7]
port 14 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 data_in[8]
port 15 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 data_in[9]
port 16 nsew signal input
rlabel metal2 s 1214 21200 1270 22000 6 select[0]
port 17 nsew signal input
rlabel metal2 s 3698 21200 3754 22000 6 select[1]
port 18 nsew signal input
rlabel metal2 s 6182 21200 6238 22000 6 select[2]
port 19 nsew signal input
rlabel metal2 s 8666 21200 8722 22000 6 select[3]
port 20 nsew signal input
rlabel metal4 s 1910 2128 2230 19632 6 vccd1
port 21 nsew power bidirectional
rlabel metal4 s 3842 2128 4162 19632 6 vccd1
port 21 nsew power bidirectional
rlabel metal4 s 5774 2128 6094 19632 6 vccd1
port 21 nsew power bidirectional
rlabel metal4 s 7706 2128 8026 19632 6 vccd1
port 21 nsew power bidirectional
rlabel metal4 s 2876 2128 3196 19632 6 vssd1
port 22 nsew ground bidirectional
rlabel metal4 s 4808 2128 5128 19632 6 vssd1
port 22 nsew ground bidirectional
rlabel metal4 s 6740 2128 7060 19632 6 vssd1
port 22 nsew ground bidirectional
rlabel metal4 s 8672 2128 8992 19632 6 vssd1
port 22 nsew ground bidirectional
rlabel metal3 s 9200 10888 10000 11008 6 y
port 23 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 10000 22000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 354194
string GDS_FILE /import/yukari1/lrburle/google_ring_oscillator/caravel/openlane/mux16x1_project/runs/23_11_30_09_08/results/signoff/mux16x1_project.magic.gds
string GDS_START 123234
<< end >>

