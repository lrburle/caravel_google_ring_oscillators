VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 141.925 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
    LAYER met4 ;
      RECT 138.725 -0.23 139.055 1.175 ;
      RECT 1.945 -0.23 2.275 0.945 ;
      RECT 1.945 -0.23 139.055 0.07 ;
      RECT 130.59 1.41 135.835 1.74 ;
      RECT 117.56 1.405 117.9 1.74 ;
      RECT 117.56 1.415 135.835 1.735 ;
      RECT 134.525 0.455 134.98 0.94 ;
      RECT 134.52 0.455 134.98 0.885 ;
      RECT 129.975 0.45 130.515 0.86 ;
      RECT 116.715 0.47 117.045 0.8 ;
      RECT 116.715 0.475 117.24 0.795 ;
      RECT 116.715 0.475 134.98 0.775 ;
      RECT 117.43 0.455 134.98 0.775 ;
      RECT 129.805 0.45 130.845 0.775 ;
      RECT 102.995 1.41 108.24 1.74 ;
      RECT 89.965 1.405 90.305 1.74 ;
      RECT 89.965 1.415 108.24 1.735 ;
      RECT 106.93 0.455 107.385 0.94 ;
      RECT 106.925 0.455 107.385 0.885 ;
      RECT 102.38 0.45 102.92 0.86 ;
      RECT 89.12 0.47 89.45 0.8 ;
      RECT 89.12 0.475 89.645 0.795 ;
      RECT 89.12 0.475 107.385 0.775 ;
      RECT 89.835 0.455 107.385 0.775 ;
      RECT 102.21 0.45 103.25 0.775 ;
      RECT 75.4 1.41 80.645 1.74 ;
      RECT 62.37 1.405 62.71 1.74 ;
      RECT 62.37 1.415 80.645 1.735 ;
      RECT 79.335 0.455 79.79 0.94 ;
      RECT 79.33 0.455 79.79 0.885 ;
      RECT 74.785 0.45 75.325 0.86 ;
      RECT 61.525 0.47 61.855 0.8 ;
      RECT 61.525 0.475 62.05 0.795 ;
      RECT 61.525 0.475 79.79 0.775 ;
      RECT 62.24 0.455 79.79 0.775 ;
      RECT 74.615 0.45 75.655 0.775 ;
      RECT 47.805 1.41 53.05 1.74 ;
      RECT 34.775 1.405 35.115 1.74 ;
      RECT 34.775 1.415 53.05 1.735 ;
      RECT 51.74 0.455 52.195 0.94 ;
      RECT 51.735 0.455 52.195 0.885 ;
      RECT 47.19 0.45 47.73 0.86 ;
      RECT 33.93 0.47 34.26 0.8 ;
      RECT 33.93 0.475 34.455 0.795 ;
      RECT 33.93 0.475 52.195 0.775 ;
      RECT 34.645 0.455 52.195 0.775 ;
      RECT 47.02 0.45 48.06 0.775 ;
      RECT 20.21 1.41 25.455 1.74 ;
      RECT 7.18 1.405 7.52 1.74 ;
      RECT 7.18 1.415 25.455 1.735 ;
      RECT 24.145 0.455 24.6 0.94 ;
      RECT 24.14 0.455 24.6 0.885 ;
      RECT 19.595 0.45 20.135 0.86 ;
      RECT 6.335 0.47 6.665 0.8 ;
      RECT 6.335 0.475 6.86 0.795 ;
      RECT 6.335 0.475 24.6 0.775 ;
      RECT 7.05 0.455 24.6 0.775 ;
      RECT 19.425 0.45 20.465 0.775 ;
      RECT 120.16 2.14 130.005 2.475 ;
      RECT 92.565 2.14 102.41 2.475 ;
      RECT 64.97 2.14 74.815 2.475 ;
      RECT 37.375 2.14 47.22 2.475 ;
      RECT 9.78 2.14 19.625 2.475 ;
    LAYER via3 ;
      RECT 138.79 0.905 138.99 1.105 ;
      RECT 135.57 1.475 135.77 1.675 ;
      RECT 134.715 0.605 134.915 0.805 ;
      RECT 131.435 1.475 131.635 1.675 ;
      RECT 130.175 0.545 130.375 0.745 ;
      RECT 129.73 2.205 129.93 2.405 ;
      RECT 120.225 2.205 120.425 2.405 ;
      RECT 117.635 1.475 117.835 1.675 ;
      RECT 116.78 0.535 116.98 0.735 ;
      RECT 107.975 1.475 108.175 1.675 ;
      RECT 107.12 0.605 107.32 0.805 ;
      RECT 103.84 1.475 104.04 1.675 ;
      RECT 102.58 0.545 102.78 0.745 ;
      RECT 102.135 2.205 102.335 2.405 ;
      RECT 92.63 2.205 92.83 2.405 ;
      RECT 90.04 1.475 90.24 1.675 ;
      RECT 89.185 0.535 89.385 0.735 ;
      RECT 80.38 1.475 80.58 1.675 ;
      RECT 79.525 0.605 79.725 0.805 ;
      RECT 76.245 1.475 76.445 1.675 ;
      RECT 74.985 0.545 75.185 0.745 ;
      RECT 74.54 2.205 74.74 2.405 ;
      RECT 65.035 2.205 65.235 2.405 ;
      RECT 62.445 1.475 62.645 1.675 ;
      RECT 61.59 0.535 61.79 0.735 ;
      RECT 52.785 1.475 52.985 1.675 ;
      RECT 51.93 0.605 52.13 0.805 ;
      RECT 48.65 1.475 48.85 1.675 ;
      RECT 47.39 0.545 47.59 0.745 ;
      RECT 46.945 2.205 47.145 2.405 ;
      RECT 37.44 2.205 37.64 2.405 ;
      RECT 34.85 1.475 35.05 1.675 ;
      RECT 33.995 0.535 34.195 0.735 ;
      RECT 25.19 1.475 25.39 1.675 ;
      RECT 24.335 0.605 24.535 0.805 ;
      RECT 21.055 1.475 21.255 1.675 ;
      RECT 19.795 0.545 19.995 0.745 ;
      RECT 19.35 2.205 19.55 2.405 ;
      RECT 9.845 2.205 10.045 2.405 ;
      RECT 7.255 1.475 7.455 1.675 ;
      RECT 6.4 0.535 6.6 0.735 ;
      RECT 2.01 0.68 2.21 0.88 ;
    LAYER met3 ;
      RECT 129.65 2.14 129.99 2.495 ;
      RECT 133.67 0.35 134.04 2.47 ;
      RECT 129.655 2.1 134.04 2.47 ;
      RECT 129.655 1.16 130.005 2.47 ;
      RECT 129.655 1.16 130.025 1.53 ;
      RECT 127.36 1.475 127.69 2.205 ;
      RECT 127.36 1.475 128.32 1.805 ;
      RECT 127.99 -0.18 128.32 1.805 ;
      RECT 127.97 -0.18 128.34 0.19 ;
      RECT 114.29 1.47 114.755 1.84 ;
      RECT 114.42 -0.17 114.755 1.84 ;
      RECT 123.72 0.515 124.05 1.245 ;
      RECT 122.84 -0.17 123.17 1.245 ;
      RECT 126.88 0.35 127.21 1.08 ;
      RECT 126.84 0.235 127.02 0.885 ;
      RECT 122.84 0.515 127.21 0.85 ;
      RECT 122.84 -0.09 123.175 0.85 ;
      RECT 122.835 -0.09 123.175 0.245 ;
      RECT 114.42 -0.17 114.925 0.245 ;
      RECT 114.42 -0.17 123.17 0.13 ;
      RECT 123.34 2.035 123.67 2.365 ;
      RECT 122.135 2.05 123.67 2.35 ;
      RECT 122.135 0.93 122.435 2.35 ;
      RECT 121.88 0.915 122.21 1.245 ;
      RECT 120.165 0.355 120.485 2.495 ;
      RECT 120.16 0.355 120.49 2.48 ;
      RECT 102.055 2.14 102.395 2.495 ;
      RECT 106.075 0.35 106.445 2.47 ;
      RECT 102.06 2.1 106.445 2.47 ;
      RECT 102.06 1.16 102.41 2.47 ;
      RECT 102.06 1.16 102.43 1.53 ;
      RECT 99.765 1.475 100.095 2.205 ;
      RECT 99.765 1.475 100.725 1.805 ;
      RECT 100.395 -0.18 100.725 1.805 ;
      RECT 100.375 -0.18 100.745 0.19 ;
      RECT 86.695 1.47 87.16 1.84 ;
      RECT 86.825 -0.17 87.16 1.84 ;
      RECT 96.125 0.515 96.455 1.245 ;
      RECT 95.245 -0.17 95.575 1.245 ;
      RECT 99.285 0.35 99.615 1.08 ;
      RECT 99.245 0.235 99.425 0.885 ;
      RECT 95.245 0.515 99.615 0.85 ;
      RECT 95.245 -0.09 95.58 0.85 ;
      RECT 95.24 -0.09 95.58 0.245 ;
      RECT 86.825 -0.17 87.33 0.245 ;
      RECT 86.825 -0.17 95.575 0.13 ;
      RECT 95.745 2.035 96.075 2.365 ;
      RECT 94.54 2.05 96.075 2.35 ;
      RECT 94.54 0.93 94.84 2.35 ;
      RECT 94.285 0.915 94.615 1.245 ;
      RECT 92.57 0.355 92.89 2.495 ;
      RECT 92.565 0.355 92.895 2.48 ;
      RECT 74.46 2.14 74.8 2.495 ;
      RECT 78.48 0.35 78.85 2.47 ;
      RECT 74.465 2.1 78.85 2.47 ;
      RECT 74.465 1.16 74.815 2.47 ;
      RECT 74.465 1.16 74.835 1.53 ;
      RECT 72.17 1.475 72.5 2.205 ;
      RECT 72.17 1.475 73.13 1.805 ;
      RECT 72.8 -0.18 73.13 1.805 ;
      RECT 72.78 -0.18 73.15 0.19 ;
      RECT 59.1 1.47 59.565 1.84 ;
      RECT 59.23 -0.17 59.565 1.84 ;
      RECT 68.53 0.515 68.86 1.245 ;
      RECT 67.65 -0.17 67.98 1.245 ;
      RECT 71.69 0.35 72.02 1.08 ;
      RECT 71.65 0.235 71.83 0.885 ;
      RECT 67.65 0.515 72.02 0.85 ;
      RECT 67.65 -0.09 67.985 0.85 ;
      RECT 67.645 -0.09 67.985 0.245 ;
      RECT 59.23 -0.17 59.735 0.245 ;
      RECT 59.23 -0.17 67.98 0.13 ;
      RECT 68.15 2.035 68.48 2.365 ;
      RECT 66.945 2.05 68.48 2.35 ;
      RECT 66.945 0.93 67.245 2.35 ;
      RECT 66.69 0.915 67.02 1.245 ;
      RECT 64.975 0.355 65.295 2.495 ;
      RECT 64.97 0.355 65.3 2.48 ;
      RECT 46.865 2.14 47.205 2.495 ;
      RECT 50.885 0.35 51.255 2.47 ;
      RECT 46.87 2.1 51.255 2.47 ;
      RECT 46.87 1.16 47.22 2.47 ;
      RECT 46.87 1.16 47.24 1.53 ;
      RECT 44.575 1.475 44.905 2.205 ;
      RECT 44.575 1.475 45.535 1.805 ;
      RECT 45.205 -0.18 45.535 1.805 ;
      RECT 45.185 -0.18 45.555 0.19 ;
      RECT 31.505 1.47 31.97 1.84 ;
      RECT 31.635 -0.17 31.97 1.84 ;
      RECT 40.935 0.515 41.265 1.245 ;
      RECT 40.055 -0.17 40.385 1.245 ;
      RECT 44.095 0.35 44.425 1.08 ;
      RECT 44.055 0.235 44.235 0.885 ;
      RECT 40.055 0.515 44.425 0.85 ;
      RECT 40.055 -0.09 40.39 0.85 ;
      RECT 40.05 -0.09 40.39 0.245 ;
      RECT 31.635 -0.17 32.14 0.245 ;
      RECT 31.635 -0.17 40.385 0.13 ;
      RECT 40.555 2.035 40.885 2.365 ;
      RECT 39.35 2.05 40.885 2.35 ;
      RECT 39.35 0.93 39.65 2.35 ;
      RECT 39.095 0.915 39.425 1.245 ;
      RECT 37.38 0.355 37.7 2.495 ;
      RECT 37.375 0.355 37.705 2.48 ;
      RECT 19.27 2.14 19.61 2.495 ;
      RECT 23.29 0.35 23.66 2.47 ;
      RECT 19.275 2.1 23.66 2.47 ;
      RECT 19.275 1.16 19.625 2.47 ;
      RECT 19.275 1.16 19.645 1.53 ;
      RECT 16.98 1.475 17.31 2.205 ;
      RECT 16.98 1.475 17.94 1.805 ;
      RECT 17.61 -0.18 17.94 1.805 ;
      RECT 17.59 -0.18 17.96 0.19 ;
      RECT 3.91 1.47 4.375 1.84 ;
      RECT 4.04 -0.17 4.375 1.84 ;
      RECT 13.34 0.515 13.67 1.245 ;
      RECT 12.46 -0.17 12.79 1.245 ;
      RECT 16.5 0.35 16.83 1.08 ;
      RECT 16.46 0.235 16.64 0.885 ;
      RECT 12.46 0.515 16.83 0.85 ;
      RECT 12.46 -0.09 12.795 0.85 ;
      RECT 12.455 -0.09 12.795 0.245 ;
      RECT 4.04 -0.17 4.545 0.245 ;
      RECT 4.04 -0.17 12.79 0.13 ;
      RECT 12.96 2.035 13.29 2.365 ;
      RECT 11.755 2.05 13.29 2.35 ;
      RECT 11.755 0.93 12.055 2.35 ;
      RECT 11.5 0.915 11.83 1.245 ;
      RECT 9.785 0.355 10.105 2.495 ;
      RECT 9.78 0.355 10.11 2.48 ;
      RECT 138.685 0.8 139.055 1.515 ;
      RECT 135.37 1.335 135.91 1.805 ;
      RECT 134.525 0.455 135.065 0.92 ;
      RECT 131.235 1.335 131.775 1.8 ;
      RECT 129.975 0.395 130.515 0.86 ;
      RECT 125.28 1.075 125.61 1.805 ;
      RECT 121.16 0.915 121.49 1.645 ;
      RECT 118.72 1.075 119.05 1.805 ;
      RECT 117.375 1.33 117.915 1.795 ;
      RECT 116.23 0.45 117.43 0.855 ;
      RECT 107.775 1.335 108.315 1.805 ;
      RECT 106.93 0.455 107.47 0.92 ;
      RECT 103.64 1.335 104.18 1.8 ;
      RECT 102.38 0.395 102.92 0.86 ;
      RECT 97.685 1.075 98.015 1.805 ;
      RECT 93.565 0.915 93.895 1.645 ;
      RECT 91.125 1.075 91.455 1.805 ;
      RECT 89.78 1.33 90.32 1.795 ;
      RECT 88.635 0.45 89.835 0.855 ;
      RECT 80.18 1.335 80.72 1.805 ;
      RECT 79.335 0.455 79.875 0.92 ;
      RECT 76.045 1.335 76.585 1.8 ;
      RECT 74.785 0.395 75.325 0.86 ;
      RECT 70.09 1.075 70.42 1.805 ;
      RECT 65.97 0.915 66.3 1.645 ;
      RECT 63.53 1.075 63.86 1.805 ;
      RECT 62.185 1.33 62.725 1.795 ;
      RECT 61.04 0.45 62.24 0.855 ;
      RECT 52.585 1.335 53.125 1.805 ;
      RECT 51.74 0.455 52.28 0.92 ;
      RECT 48.45 1.335 48.99 1.8 ;
      RECT 47.19 0.395 47.73 0.86 ;
      RECT 42.495 1.075 42.825 1.805 ;
      RECT 38.375 0.915 38.705 1.645 ;
      RECT 35.935 1.075 36.265 1.805 ;
      RECT 34.59 1.33 35.13 1.795 ;
      RECT 33.445 0.45 34.645 0.855 ;
      RECT 24.99 1.335 25.53 1.805 ;
      RECT 24.145 0.455 24.685 0.92 ;
      RECT 20.855 1.335 21.395 1.8 ;
      RECT 19.595 0.395 20.135 0.86 ;
      RECT 14.9 1.075 15.23 1.805 ;
      RECT 10.78 0.915 11.11 1.645 ;
      RECT 8.34 1.075 8.67 1.805 ;
      RECT 6.995 1.33 7.535 1.795 ;
      RECT 5.85 0.45 7.05 0.855 ;
      RECT 1.875 0.53 2.36 1.04 ;
    LAYER via2 ;
      RECT 138.77 0.885 138.97 1.085 ;
      RECT 135.55 1.455 135.75 1.655 ;
      RECT 134.695 0.585 134.895 0.785 ;
      RECT 133.755 0.435 133.955 0.635 ;
      RECT 131.415 1.455 131.615 1.655 ;
      RECT 130.155 0.525 130.355 0.725 ;
      RECT 129.74 1.245 129.94 1.445 ;
      RECT 128.055 -0.095 128.255 0.105 ;
      RECT 127.425 1.54 127.625 1.74 ;
      RECT 126.945 0.815 127.145 1.015 ;
      RECT 125.345 1.54 125.545 1.74 ;
      RECT 123.785 0.98 123.985 1.18 ;
      RECT 123.405 2.1 123.605 2.3 ;
      RECT 122.905 0.98 123.105 1.18 ;
      RECT 121.945 0.98 122.145 1.18 ;
      RECT 121.225 0.98 121.425 1.18 ;
      RECT 120.225 0.42 120.425 0.62 ;
      RECT 118.785 1.54 118.985 1.74 ;
      RECT 117.615 1.455 117.815 1.655 ;
      RECT 116.76 0.515 116.96 0.715 ;
      RECT 114.375 1.555 114.575 1.755 ;
      RECT 107.955 1.455 108.155 1.655 ;
      RECT 107.1 0.585 107.3 0.785 ;
      RECT 106.16 0.435 106.36 0.635 ;
      RECT 103.82 1.455 104.02 1.655 ;
      RECT 102.56 0.525 102.76 0.725 ;
      RECT 102.145 1.245 102.345 1.445 ;
      RECT 100.46 -0.095 100.66 0.105 ;
      RECT 99.83 1.54 100.03 1.74 ;
      RECT 99.35 0.815 99.55 1.015 ;
      RECT 97.75 1.54 97.95 1.74 ;
      RECT 96.19 0.98 96.39 1.18 ;
      RECT 95.81 2.1 96.01 2.3 ;
      RECT 95.31 0.98 95.51 1.18 ;
      RECT 94.35 0.98 94.55 1.18 ;
      RECT 93.63 0.98 93.83 1.18 ;
      RECT 92.63 0.42 92.83 0.62 ;
      RECT 91.19 1.54 91.39 1.74 ;
      RECT 90.02 1.455 90.22 1.655 ;
      RECT 89.165 0.515 89.365 0.715 ;
      RECT 86.78 1.555 86.98 1.755 ;
      RECT 80.36 1.455 80.56 1.655 ;
      RECT 79.505 0.585 79.705 0.785 ;
      RECT 78.565 0.435 78.765 0.635 ;
      RECT 76.225 1.455 76.425 1.655 ;
      RECT 74.965 0.525 75.165 0.725 ;
      RECT 74.55 1.245 74.75 1.445 ;
      RECT 72.865 -0.095 73.065 0.105 ;
      RECT 72.235 1.54 72.435 1.74 ;
      RECT 71.755 0.815 71.955 1.015 ;
      RECT 70.155 1.54 70.355 1.74 ;
      RECT 68.595 0.98 68.795 1.18 ;
      RECT 68.215 2.1 68.415 2.3 ;
      RECT 67.715 0.98 67.915 1.18 ;
      RECT 66.755 0.98 66.955 1.18 ;
      RECT 66.035 0.98 66.235 1.18 ;
      RECT 65.035 0.42 65.235 0.62 ;
      RECT 63.595 1.54 63.795 1.74 ;
      RECT 62.425 1.455 62.625 1.655 ;
      RECT 61.57 0.515 61.77 0.715 ;
      RECT 59.185 1.555 59.385 1.755 ;
      RECT 52.765 1.455 52.965 1.655 ;
      RECT 51.91 0.585 52.11 0.785 ;
      RECT 50.97 0.435 51.17 0.635 ;
      RECT 48.63 1.455 48.83 1.655 ;
      RECT 47.37 0.525 47.57 0.725 ;
      RECT 46.955 1.245 47.155 1.445 ;
      RECT 45.27 -0.095 45.47 0.105 ;
      RECT 44.64 1.54 44.84 1.74 ;
      RECT 44.16 0.815 44.36 1.015 ;
      RECT 42.56 1.54 42.76 1.74 ;
      RECT 41 0.98 41.2 1.18 ;
      RECT 40.62 2.1 40.82 2.3 ;
      RECT 40.12 0.98 40.32 1.18 ;
      RECT 39.16 0.98 39.36 1.18 ;
      RECT 38.44 0.98 38.64 1.18 ;
      RECT 37.44 0.42 37.64 0.62 ;
      RECT 36 1.54 36.2 1.74 ;
      RECT 34.83 1.455 35.03 1.655 ;
      RECT 33.975 0.515 34.175 0.715 ;
      RECT 31.59 1.555 31.79 1.755 ;
      RECT 25.17 1.455 25.37 1.655 ;
      RECT 24.315 0.585 24.515 0.785 ;
      RECT 23.375 0.435 23.575 0.635 ;
      RECT 21.035 1.455 21.235 1.655 ;
      RECT 19.775 0.525 19.975 0.725 ;
      RECT 19.36 1.245 19.56 1.445 ;
      RECT 17.675 -0.095 17.875 0.105 ;
      RECT 17.045 1.54 17.245 1.74 ;
      RECT 16.565 0.815 16.765 1.015 ;
      RECT 14.965 1.54 15.165 1.74 ;
      RECT 13.405 0.98 13.605 1.18 ;
      RECT 13.025 2.1 13.225 2.3 ;
      RECT 12.525 0.98 12.725 1.18 ;
      RECT 11.565 0.98 11.765 1.18 ;
      RECT 10.845 0.98 11.045 1.18 ;
      RECT 9.845 0.42 10.045 0.62 ;
      RECT 8.405 1.54 8.605 1.74 ;
      RECT 7.235 1.455 7.435 1.655 ;
      RECT 6.38 0.515 6.58 0.715 ;
      RECT 3.995 1.555 4.195 1.755 ;
      RECT 2.01 0.68 2.21 0.88 ;
    LAYER met2 ;
      RECT 133.67 0.35 134.04 0.72 ;
      RECT 134.185 0.365 134.445 0.69 ;
      RECT 133.67 0.395 134.445 0.655 ;
      RECT 124.455 0.955 124.69 1.215 ;
      RECT 127.6 0.735 127.765 0.995 ;
      RECT 127.505 0.725 127.52 0.995 ;
      RECT 126.105 0.295 126.145 0.435 ;
      RECT 127.52 0.73 127.6 0.995 ;
      RECT 127.465 0.725 127.505 0.961 ;
      RECT 127.451 0.725 127.465 0.961 ;
      RECT 127.365 0.73 127.451 0.963 ;
      RECT 127.32 0.737 127.365 0.965 ;
      RECT 127.29 0.737 127.32 0.967 ;
      RECT 127.265 0.732 127.29 0.969 ;
      RECT 127.235 0.728 127.265 0.978 ;
      RECT 127.225 0.725 127.235 0.99 ;
      RECT 127.22 0.725 127.225 0.998 ;
      RECT 127.215 0.725 127.22 1.003 ;
      RECT 127.205 0.724 127.215 1.013 ;
      RECT 127.2 0.723 127.205 1.023 ;
      RECT 127.185 0.722 127.2 1.028 ;
      RECT 127.157 0.719 127.185 1.055 ;
      RECT 127.071 0.711 127.157 1.055 ;
      RECT 126.985 0.7 127.071 1.055 ;
      RECT 126.945 0.685 126.985 1.055 ;
      RECT 126.905 0.659 126.945 1.055 ;
      RECT 126.9 0.641 126.905 0.867 ;
      RECT 126.89 0.637 126.9 0.857 ;
      RECT 126.875 0.627 126.89 0.844 ;
      RECT 126.855 0.611 126.875 0.829 ;
      RECT 126.84 0.596 126.855 0.814 ;
      RECT 126.83 0.585 126.84 0.804 ;
      RECT 126.805 0.569 126.83 0.793 ;
      RECT 126.8 0.556 126.805 0.783 ;
      RECT 126.795 0.552 126.8 0.778 ;
      RECT 126.74 0.538 126.795 0.756 ;
      RECT 126.701 0.519 126.74 0.72 ;
      RECT 126.615 0.493 126.701 0.673 ;
      RECT 126.611 0.475 126.615 0.639 ;
      RECT 126.525 0.456 126.611 0.617 ;
      RECT 126.52 0.438 126.525 0.595 ;
      RECT 126.515 0.436 126.52 0.593 ;
      RECT 126.505 0.435 126.515 0.588 ;
      RECT 126.445 0.422 126.505 0.574 ;
      RECT 126.4 0.4 126.445 0.553 ;
      RECT 126.34 0.377 126.4 0.532 ;
      RECT 126.276 0.352 126.34 0.507 ;
      RECT 126.19 0.322 126.276 0.476 ;
      RECT 126.175 0.302 126.19 0.455 ;
      RECT 126.145 0.297 126.175 0.446 ;
      RECT 126.092 0.295 126.105 0.435 ;
      RECT 126.006 0.295 126.092 0.437 ;
      RECT 125.92 0.295 126.006 0.439 ;
      RECT 125.9 0.295 125.92 0.443 ;
      RECT 125.855 0.297 125.9 0.454 ;
      RECT 125.815 0.307 125.855 0.47 ;
      RECT 125.811 0.316 125.815 0.478 ;
      RECT 125.725 0.336 125.811 0.494 ;
      RECT 125.715 0.355 125.725 0.512 ;
      RECT 125.71 0.357 125.715 0.515 ;
      RECT 125.7 0.361 125.71 0.518 ;
      RECT 125.68 0.366 125.7 0.528 ;
      RECT 125.65 0.376 125.68 0.548 ;
      RECT 125.645 0.383 125.65 0.562 ;
      RECT 125.635 0.387 125.645 0.569 ;
      RECT 125.62 0.395 125.635 0.58 ;
      RECT 125.61 0.405 125.62 0.591 ;
      RECT 125.6 0.412 125.61 0.599 ;
      RECT 125.575 0.425 125.6 0.614 ;
      RECT 125.511 0.461 125.575 0.653 ;
      RECT 125.425 0.524 125.511 0.717 ;
      RECT 125.39 0.575 125.425 0.77 ;
      RECT 125.385 0.592 125.39 0.787 ;
      RECT 125.37 0.601 125.385 0.794 ;
      RECT 125.35 0.616 125.37 0.808 ;
      RECT 125.345 0.627 125.35 0.818 ;
      RECT 125.325 0.64 125.345 0.828 ;
      RECT 125.32 0.65 125.325 0.838 ;
      RECT 125.305 0.655 125.32 0.847 ;
      RECT 125.295 0.665 125.305 0.858 ;
      RECT 125.265 0.682 125.295 0.875 ;
      RECT 125.255 0.7 125.265 0.893 ;
      RECT 125.24 0.711 125.255 0.904 ;
      RECT 125.2 0.735 125.24 0.92 ;
      RECT 125.165 0.769 125.2 0.937 ;
      RECT 125.135 0.792 125.165 0.949 ;
      RECT 125.12 0.802 125.135 0.958 ;
      RECT 125.08 0.812 125.12 0.969 ;
      RECT 125.06 0.823 125.08 0.981 ;
      RECT 125.055 0.827 125.06 0.988 ;
      RECT 125.04 0.831 125.055 0.993 ;
      RECT 125.03 0.836 125.04 0.998 ;
      RECT 125.025 0.839 125.03 1.001 ;
      RECT 124.995 0.845 125.025 1.008 ;
      RECT 124.96 0.855 124.995 1.022 ;
      RECT 124.9 0.87 124.96 1.042 ;
      RECT 124.845 0.89 124.9 1.066 ;
      RECT 124.816 0.905 124.845 1.084 ;
      RECT 124.73 0.925 124.816 1.109 ;
      RECT 124.725 0.94 124.73 1.129 ;
      RECT 124.715 0.943 124.725 1.13 ;
      RECT 124.69 0.95 124.715 1.215 ;
      RECT 127.385 1.443 127.665 1.78 ;
      RECT 127.385 1.453 127.67 1.738 ;
      RECT 127.385 1.462 127.675 1.635 ;
      RECT 127.385 1.477 127.68 1.503 ;
      RECT 127.385 1.305 127.645 1.78 ;
      RECT 125.105 2.185 125.115 2.375 ;
      RECT 123.365 2.06 123.645 2.34 ;
      RECT 126.41 1 126.415 1.485 ;
      RECT 126.305 1 126.365 1.26 ;
      RECT 126.63 1.97 126.635 2.045 ;
      RECT 126.62 1.837 126.63 2.08 ;
      RECT 126.61 1.672 126.62 2.101 ;
      RECT 126.605 1.542 126.61 2.117 ;
      RECT 126.595 1.432 126.605 2.133 ;
      RECT 126.59 1.331 126.595 2.15 ;
      RECT 126.585 1.313 126.59 2.16 ;
      RECT 126.58 1.295 126.585 2.17 ;
      RECT 126.57 1.27 126.58 2.185 ;
      RECT 126.565 1.25 126.57 2.2 ;
      RECT 126.545 1 126.565 2.225 ;
      RECT 126.53 1 126.545 2.258 ;
      RECT 126.5 1 126.53 2.28 ;
      RECT 126.48 1 126.5 2.294 ;
      RECT 126.46 1 126.48 1.81 ;
      RECT 126.475 1.877 126.48 2.299 ;
      RECT 126.47 1.907 126.475 2.301 ;
      RECT 126.465 1.92 126.47 2.304 ;
      RECT 126.46 1.93 126.465 2.308 ;
      RECT 126.455 1 126.46 1.728 ;
      RECT 126.455 1.94 126.46 2.31 ;
      RECT 126.45 1 126.455 1.705 ;
      RECT 126.44 1.962 126.455 2.31 ;
      RECT 126.435 1 126.45 1.65 ;
      RECT 126.43 1.987 126.44 2.31 ;
      RECT 126.43 1 126.435 1.595 ;
      RECT 126.42 1 126.43 1.543 ;
      RECT 126.425 2 126.43 2.311 ;
      RECT 126.42 2.012 126.425 2.312 ;
      RECT 126.415 1 126.42 1.503 ;
      RECT 126.415 2.025 126.42 2.313 ;
      RECT 126.4 2.04 126.415 2.314 ;
      RECT 126.405 1 126.41 1.465 ;
      RECT 126.4 1 126.405 1.43 ;
      RECT 126.395 1 126.4 1.405 ;
      RECT 126.39 2.067 126.4 2.316 ;
      RECT 126.385 1 126.395 1.363 ;
      RECT 126.385 2.085 126.39 2.317 ;
      RECT 126.38 1 126.385 1.323 ;
      RECT 126.38 2.092 126.385 2.318 ;
      RECT 126.375 1 126.38 1.295 ;
      RECT 126.37 2.11 126.38 2.319 ;
      RECT 126.365 1 126.375 1.275 ;
      RECT 126.36 2.13 126.37 2.321 ;
      RECT 126.35 2.147 126.36 2.322 ;
      RECT 126.315 2.17 126.35 2.325 ;
      RECT 126.26 2.188 126.315 2.331 ;
      RECT 126.174 2.196 126.26 2.34 ;
      RECT 126.088 2.207 126.174 2.351 ;
      RECT 126.002 2.217 126.088 2.362 ;
      RECT 125.916 2.227 126.002 2.374 ;
      RECT 125.83 2.237 125.916 2.385 ;
      RECT 125.81 2.243 125.83 2.391 ;
      RECT 125.73 2.245 125.81 2.395 ;
      RECT 125.725 2.244 125.73 2.4 ;
      RECT 125.717 2.243 125.725 2.4 ;
      RECT 125.631 2.239 125.717 2.398 ;
      RECT 125.545 2.231 125.631 2.395 ;
      RECT 125.459 2.222 125.545 2.391 ;
      RECT 125.373 2.214 125.459 2.388 ;
      RECT 125.287 2.206 125.373 2.384 ;
      RECT 125.201 2.197 125.287 2.381 ;
      RECT 125.115 2.189 125.201 2.377 ;
      RECT 125.06 2.182 125.105 2.375 ;
      RECT 124.975 2.175 125.06 2.373 ;
      RECT 124.901 2.167 124.975 2.369 ;
      RECT 124.815 2.159 124.901 2.366 ;
      RECT 124.812 2.155 124.815 2.364 ;
      RECT 124.726 2.151 124.812 2.363 ;
      RECT 124.64 2.143 124.726 2.36 ;
      RECT 124.555 2.138 124.64 2.357 ;
      RECT 124.469 2.135 124.555 2.354 ;
      RECT 124.383 2.133 124.469 2.351 ;
      RECT 124.297 2.13 124.383 2.348 ;
      RECT 124.211 2.127 124.297 2.345 ;
      RECT 124.125 2.124 124.211 2.342 ;
      RECT 124.049 2.122 124.125 2.339 ;
      RECT 123.963 2.119 124.049 2.336 ;
      RECT 123.877 2.116 123.963 2.334 ;
      RECT 123.791 2.114 123.877 2.331 ;
      RECT 123.705 2.111 123.791 2.328 ;
      RECT 123.645 2.102 123.705 2.326 ;
      RECT 126.155 1.72 126.23 1.98 ;
      RECT 126.135 1.7 126.14 1.98 ;
      RECT 125.455 1.485 125.56 1.78 ;
      RECT 119.9 1.46 119.97 1.72 ;
      RECT 125.795 1.335 125.8 1.706 ;
      RECT 125.785 1.39 125.79 1.706 ;
      RECT 126.09 0.56 126.15 0.82 ;
      RECT 126.145 1.715 126.155 1.98 ;
      RECT 126.14 1.705 126.145 1.98 ;
      RECT 126.06 1.652 126.135 1.98 ;
      RECT 126.085 0.56 126.09 0.84 ;
      RECT 126.075 0.56 126.085 0.86 ;
      RECT 126.06 0.56 126.075 0.89 ;
      RECT 126.045 0.56 126.06 0.933 ;
      RECT 126.04 1.595 126.06 1.98 ;
      RECT 126.03 0.56 126.045 0.97 ;
      RECT 126.025 1.575 126.04 1.98 ;
      RECT 126.025 0.56 126.03 0.993 ;
      RECT 126.015 0.56 126.025 1.018 ;
      RECT 125.985 1.542 126.025 1.98 ;
      RECT 125.99 0.56 126.015 1.068 ;
      RECT 125.985 0.56 125.99 1.123 ;
      RECT 125.98 0.56 125.985 1.165 ;
      RECT 125.97 1.505 125.985 1.98 ;
      RECT 125.975 0.56 125.98 1.208 ;
      RECT 125.97 0.56 125.975 1.273 ;
      RECT 125.965 0.56 125.97 1.295 ;
      RECT 125.965 1.493 125.97 1.845 ;
      RECT 125.96 0.56 125.965 1.363 ;
      RECT 125.96 1.485 125.965 1.828 ;
      RECT 125.955 0.56 125.96 1.408 ;
      RECT 125.95 1.467 125.96 1.805 ;
      RECT 125.95 0.56 125.955 1.445 ;
      RECT 125.94 0.56 125.95 1.785 ;
      RECT 125.935 0.56 125.94 1.768 ;
      RECT 125.93 0.56 125.935 1.753 ;
      RECT 125.925 0.56 125.93 1.738 ;
      RECT 125.905 0.56 125.925 1.728 ;
      RECT 125.9 0.56 125.905 1.718 ;
      RECT 125.89 0.56 125.9 1.714 ;
      RECT 125.885 0.837 125.89 1.713 ;
      RECT 125.88 0.86 125.885 1.712 ;
      RECT 125.875 0.89 125.88 1.711 ;
      RECT 125.87 0.917 125.875 1.71 ;
      RECT 125.865 0.945 125.87 1.71 ;
      RECT 125.86 0.972 125.865 1.71 ;
      RECT 125.855 0.992 125.86 1.71 ;
      RECT 125.85 1.02 125.855 1.71 ;
      RECT 125.84 1.062 125.85 1.71 ;
      RECT 125.83 1.107 125.84 1.709 ;
      RECT 125.825 1.16 125.83 1.708 ;
      RECT 125.82 1.192 125.825 1.707 ;
      RECT 125.815 1.212 125.82 1.706 ;
      RECT 125.81 1.25 125.815 1.706 ;
      RECT 125.805 1.272 125.81 1.706 ;
      RECT 125.8 1.297 125.805 1.706 ;
      RECT 125.79 1.362 125.795 1.706 ;
      RECT 125.775 1.422 125.785 1.706 ;
      RECT 125.76 1.432 125.775 1.706 ;
      RECT 125.74 1.442 125.76 1.706 ;
      RECT 125.71 1.447 125.74 1.703 ;
      RECT 125.65 1.457 125.71 1.7 ;
      RECT 125.63 1.466 125.65 1.705 ;
      RECT 125.605 1.472 125.63 1.718 ;
      RECT 125.585 1.477 125.605 1.733 ;
      RECT 125.56 1.482 125.585 1.78 ;
      RECT 125.431 1.484 125.455 1.78 ;
      RECT 125.345 1.479 125.431 1.78 ;
      RECT 125.305 1.476 125.345 1.78 ;
      RECT 125.255 1.478 125.305 1.76 ;
      RECT 125.225 1.482 125.255 1.76 ;
      RECT 125.146 1.492 125.225 1.76 ;
      RECT 125.06 1.507 125.146 1.761 ;
      RECT 125.01 1.517 125.06 1.762 ;
      RECT 125.002 1.52 125.01 1.762 ;
      RECT 124.916 1.522 125.002 1.763 ;
      RECT 124.83 1.526 124.916 1.763 ;
      RECT 124.744 1.53 124.83 1.764 ;
      RECT 124.658 1.533 124.744 1.765 ;
      RECT 124.572 1.537 124.658 1.765 ;
      RECT 124.486 1.541 124.572 1.766 ;
      RECT 124.4 1.544 124.486 1.767 ;
      RECT 124.314 1.548 124.4 1.767 ;
      RECT 124.228 1.552 124.314 1.768 ;
      RECT 124.142 1.556 124.228 1.769 ;
      RECT 124.056 1.559 124.142 1.769 ;
      RECT 123.97 1.563 124.056 1.77 ;
      RECT 123.94 1.565 123.97 1.77 ;
      RECT 123.854 1.568 123.94 1.771 ;
      RECT 123.768 1.572 123.854 1.772 ;
      RECT 123.682 1.576 123.768 1.773 ;
      RECT 123.596 1.579 123.682 1.773 ;
      RECT 123.51 1.583 123.596 1.774 ;
      RECT 123.475 1.588 123.51 1.775 ;
      RECT 123.42 1.598 123.475 1.782 ;
      RECT 123.395 1.61 123.42 1.792 ;
      RECT 123.36 1.623 123.395 1.8 ;
      RECT 123.32 1.64 123.36 1.823 ;
      RECT 123.3 1.653 123.32 1.85 ;
      RECT 123.27 1.665 123.3 1.878 ;
      RECT 123.265 1.673 123.27 1.898 ;
      RECT 123.26 1.676 123.265 1.908 ;
      RECT 123.21 1.688 123.26 1.942 ;
      RECT 123.2 1.703 123.21 1.975 ;
      RECT 123.19 1.709 123.2 1.988 ;
      RECT 123.18 1.716 123.19 2 ;
      RECT 123.155 1.729 123.18 2.018 ;
      RECT 123.14 1.744 123.155 2.04 ;
      RECT 123.13 1.752 123.14 2.056 ;
      RECT 123.115 1.761 123.13 2.071 ;
      RECT 123.105 1.771 123.115 2.085 ;
      RECT 123.086 1.784 123.105 2.102 ;
      RECT 123 1.829 123.086 2.167 ;
      RECT 122.985 1.874 123 2.225 ;
      RECT 122.98 1.883 122.985 2.238 ;
      RECT 122.97 1.89 122.98 2.243 ;
      RECT 122.965 1.895 122.97 2.247 ;
      RECT 122.945 1.905 122.965 2.254 ;
      RECT 122.92 1.925 122.945 2.268 ;
      RECT 122.885 1.95 122.92 2.288 ;
      RECT 122.87 1.973 122.885 2.303 ;
      RECT 122.86 1.983 122.87 2.308 ;
      RECT 122.85 1.991 122.86 2.315 ;
      RECT 122.84 2 122.85 2.321 ;
      RECT 122.82 2.012 122.84 2.323 ;
      RECT 122.81 2.025 122.82 2.325 ;
      RECT 122.785 2.04 122.81 2.328 ;
      RECT 122.765 2.057 122.785 2.332 ;
      RECT 122.725 2.085 122.765 2.338 ;
      RECT 122.66 2.132 122.725 2.347 ;
      RECT 122.645 2.165 122.66 2.355 ;
      RECT 122.64 2.172 122.645 2.357 ;
      RECT 122.59 2.197 122.64 2.362 ;
      RECT 122.575 2.221 122.59 2.369 ;
      RECT 122.525 2.226 122.575 2.37 ;
      RECT 122.439 2.23 122.525 2.37 ;
      RECT 122.353 2.23 122.439 2.37 ;
      RECT 122.267 2.23 122.353 2.371 ;
      RECT 122.181 2.23 122.267 2.371 ;
      RECT 122.095 2.23 122.181 2.371 ;
      RECT 122.029 2.23 122.095 2.371 ;
      RECT 121.943 2.23 122.029 2.372 ;
      RECT 121.857 2.23 121.943 2.372 ;
      RECT 121.771 2.231 121.857 2.373 ;
      RECT 121.685 2.231 121.771 2.373 ;
      RECT 121.599 2.231 121.685 2.373 ;
      RECT 121.513 2.231 121.599 2.374 ;
      RECT 121.427 2.231 121.513 2.374 ;
      RECT 121.341 2.232 121.427 2.375 ;
      RECT 121.255 2.232 121.341 2.375 ;
      RECT 121.235 2.232 121.255 2.375 ;
      RECT 121.149 2.232 121.235 2.375 ;
      RECT 121.063 2.232 121.149 2.375 ;
      RECT 120.977 2.233 121.063 2.375 ;
      RECT 120.891 2.233 120.977 2.375 ;
      RECT 120.805 2.233 120.891 2.375 ;
      RECT 120.719 2.234 120.805 2.375 ;
      RECT 120.633 2.234 120.719 2.375 ;
      RECT 120.547 2.234 120.633 2.375 ;
      RECT 120.461 2.234 120.547 2.375 ;
      RECT 120.375 2.235 120.461 2.375 ;
      RECT 120.325 2.232 120.375 2.375 ;
      RECT 120.315 2.23 120.325 2.374 ;
      RECT 120.311 2.23 120.315 2.373 ;
      RECT 120.225 2.225 120.311 2.368 ;
      RECT 120.203 2.218 120.225 2.362 ;
      RECT 120.117 2.209 120.203 2.356 ;
      RECT 120.031 2.196 120.117 2.347 ;
      RECT 119.945 2.182 120.031 2.337 ;
      RECT 119.9 2.172 119.945 2.33 ;
      RECT 119.88 1.46 119.9 1.738 ;
      RECT 119.88 2.165 119.9 2.326 ;
      RECT 119.85 1.46 119.88 1.76 ;
      RECT 119.84 2.132 119.88 2.323 ;
      RECT 119.835 1.46 119.85 1.78 ;
      RECT 119.835 2.097 119.84 2.321 ;
      RECT 119.83 1.46 119.835 1.905 ;
      RECT 119.83 2.057 119.835 2.321 ;
      RECT 119.82 1.46 119.83 2.321 ;
      RECT 119.745 1.46 119.82 2.315 ;
      RECT 119.715 1.46 119.745 2.305 ;
      RECT 119.71 1.46 119.715 2.297 ;
      RECT 119.705 1.502 119.71 2.29 ;
      RECT 119.695 1.571 119.705 2.281 ;
      RECT 119.69 1.641 119.695 2.233 ;
      RECT 119.685 1.705 119.69 2.13 ;
      RECT 119.68 1.74 119.685 2.085 ;
      RECT 119.678 1.777 119.68 1.977 ;
      RECT 119.675 1.785 119.678 1.97 ;
      RECT 119.67 1.85 119.675 1.913 ;
      RECT 123.745 0.94 124.025 1.22 ;
      RECT 123.735 0.94 124.025 1.083 ;
      RECT 123.69 0.805 123.95 1.065 ;
      RECT 123.69 0.92 124.005 1.065 ;
      RECT 123.69 0.89 124 1.065 ;
      RECT 123.69 0.877 123.99 1.065 ;
      RECT 123.69 0.867 123.985 1.065 ;
      RECT 119.665 0.85 119.925 1.11 ;
      RECT 123.435 0.4 123.695 0.66 ;
      RECT 123.425 0.425 123.695 0.62 ;
      RECT 123.42 0.425 123.425 0.619 ;
      RECT 123.35 0.42 123.42 0.611 ;
      RECT 123.265 0.407 123.35 0.594 ;
      RECT 123.261 0.399 123.265 0.584 ;
      RECT 123.175 0.392 123.261 0.574 ;
      RECT 123.166 0.384 123.175 0.564 ;
      RECT 123.08 0.377 123.166 0.552 ;
      RECT 123.06 0.368 123.08 0.538 ;
      RECT 123.005 0.363 123.06 0.53 ;
      RECT 122.995 0.357 123.005 0.524 ;
      RECT 122.975 0.355 122.995 0.52 ;
      RECT 122.967 0.354 122.975 0.516 ;
      RECT 122.881 0.346 122.967 0.505 ;
      RECT 122.795 0.332 122.881 0.485 ;
      RECT 122.735 0.32 122.795 0.47 ;
      RECT 122.725 0.315 122.735 0.465 ;
      RECT 122.675 0.315 122.725 0.467 ;
      RECT 122.628 0.317 122.675 0.471 ;
      RECT 122.542 0.324 122.628 0.476 ;
      RECT 122.456 0.332 122.542 0.482 ;
      RECT 122.37 0.341 122.456 0.488 ;
      RECT 122.311 0.347 122.37 0.493 ;
      RECT 122.225 0.352 122.311 0.499 ;
      RECT 122.15 0.357 122.225 0.505 ;
      RECT 122.111 0.359 122.15 0.51 ;
      RECT 122.025 0.356 122.111 0.515 ;
      RECT 121.94 0.354 122.025 0.522 ;
      RECT 121.908 0.353 121.94 0.525 ;
      RECT 121.822 0.352 121.908 0.526 ;
      RECT 121.736 0.351 121.822 0.527 ;
      RECT 121.65 0.35 121.736 0.527 ;
      RECT 121.564 0.349 121.65 0.528 ;
      RECT 121.478 0.348 121.564 0.529 ;
      RECT 121.392 0.347 121.478 0.53 ;
      RECT 121.306 0.346 121.392 0.53 ;
      RECT 121.22 0.345 121.306 0.531 ;
      RECT 121.17 0.345 121.22 0.532 ;
      RECT 121.156 0.346 121.17 0.532 ;
      RECT 121.07 0.353 121.156 0.533 ;
      RECT 120.996 0.364 121.07 0.534 ;
      RECT 120.91 0.373 120.996 0.535 ;
      RECT 120.875 0.38 120.91 0.55 ;
      RECT 120.85 0.383 120.875 0.58 ;
      RECT 120.825 0.392 120.85 0.609 ;
      RECT 120.815 0.403 120.825 0.629 ;
      RECT 120.805 0.411 120.815 0.643 ;
      RECT 120.8 0.417 120.805 0.653 ;
      RECT 120.775 0.434 120.8 0.67 ;
      RECT 120.76 0.456 120.775 0.698 ;
      RECT 120.73 0.482 120.76 0.728 ;
      RECT 120.71 0.511 120.73 0.758 ;
      RECT 120.705 0.526 120.71 0.775 ;
      RECT 120.685 0.541 120.705 0.79 ;
      RECT 120.675 0.559 120.685 0.808 ;
      RECT 120.665 0.57 120.675 0.823 ;
      RECT 120.615 0.602 120.665 0.849 ;
      RECT 120.61 0.632 120.615 0.869 ;
      RECT 120.6 0.645 120.61 0.875 ;
      RECT 120.591 0.655 120.6 0.883 ;
      RECT 120.58 0.666 120.591 0.891 ;
      RECT 120.575 0.676 120.58 0.897 ;
      RECT 120.56 0.697 120.575 0.904 ;
      RECT 120.545 0.727 120.56 0.912 ;
      RECT 120.51 0.757 120.545 0.918 ;
      RECT 120.485 0.775 120.51 0.925 ;
      RECT 120.435 0.783 120.485 0.934 ;
      RECT 120.41 0.788 120.435 0.943 ;
      RECT 120.355 0.794 120.41 0.953 ;
      RECT 120.35 0.799 120.355 0.961 ;
      RECT 120.336 0.802 120.35 0.963 ;
      RECT 120.25 0.814 120.336 0.975 ;
      RECT 120.24 0.826 120.25 0.988 ;
      RECT 120.155 0.839 120.24 1 ;
      RECT 120.111 0.856 120.155 1.014 ;
      RECT 120.025 0.873 120.111 1.03 ;
      RECT 119.995 0.887 120.025 1.044 ;
      RECT 119.985 0.892 119.995 1.049 ;
      RECT 119.925 0.895 119.985 1.058 ;
      RECT 122.815 1.165 123.075 1.425 ;
      RECT 122.815 1.165 123.095 1.278 ;
      RECT 122.815 1.165 123.12 1.245 ;
      RECT 122.815 1.165 123.125 1.225 ;
      RECT 122.865 0.94 123.145 1.22 ;
      RECT 122.42 1.675 122.68 1.935 ;
      RECT 122.41 1.532 122.605 1.873 ;
      RECT 122.405 1.64 122.62 1.865 ;
      RECT 122.4 1.69 122.68 1.855 ;
      RECT 122.39 1.767 122.68 1.84 ;
      RECT 122.41 1.615 122.62 1.873 ;
      RECT 122.42 1.49 122.605 1.935 ;
      RECT 122.42 1.385 122.585 1.935 ;
      RECT 122.43 1.372 122.585 1.935 ;
      RECT 122.43 1.33 122.575 1.935 ;
      RECT 122.435 1.255 122.575 1.935 ;
      RECT 122.465 0.905 122.575 1.935 ;
      RECT 122.47 0.635 122.595 1.258 ;
      RECT 122.44 1.21 122.595 1.258 ;
      RECT 122.455 1.012 122.575 1.935 ;
      RECT 122.445 1.122 122.595 1.258 ;
      RECT 122.47 0.635 122.61 1.115 ;
      RECT 122.47 0.635 122.63 0.99 ;
      RECT 122.435 0.635 122.695 0.895 ;
      RECT 121.905 0.94 122.185 1.22 ;
      RECT 121.89 0.94 122.185 1.2 ;
      RECT 119.945 1.805 120.205 2.065 ;
      RECT 121.73 1.66 121.99 1.92 ;
      RECT 121.71 1.68 121.99 1.895 ;
      RECT 121.667 1.68 121.71 1.894 ;
      RECT 121.581 1.681 121.667 1.891 ;
      RECT 121.495 1.682 121.581 1.887 ;
      RECT 121.42 1.684 121.495 1.884 ;
      RECT 121.397 1.685 121.42 1.882 ;
      RECT 121.311 1.686 121.397 1.88 ;
      RECT 121.225 1.687 121.311 1.877 ;
      RECT 121.201 1.688 121.225 1.875 ;
      RECT 121.115 1.69 121.201 1.872 ;
      RECT 121.03 1.692 121.115 1.873 ;
      RECT 120.973 1.693 121.03 1.879 ;
      RECT 120.887 1.695 120.973 1.889 ;
      RECT 120.801 1.698 120.887 1.902 ;
      RECT 120.715 1.7 120.801 1.914 ;
      RECT 120.701 1.701 120.715 1.921 ;
      RECT 120.615 1.702 120.701 1.929 ;
      RECT 120.575 1.704 120.615 1.938 ;
      RECT 120.566 1.705 120.575 1.941 ;
      RECT 120.48 1.713 120.566 1.947 ;
      RECT 120.46 1.722 120.48 1.955 ;
      RECT 120.375 1.737 120.46 1.963 ;
      RECT 120.315 1.76 120.375 1.974 ;
      RECT 120.305 1.772 120.315 1.979 ;
      RECT 120.265 1.782 120.305 1.983 ;
      RECT 120.21 1.799 120.265 1.991 ;
      RECT 120.205 1.809 120.21 1.995 ;
      RECT 121.271 0.94 121.33 1.337 ;
      RECT 121.185 0.94 121.39 1.328 ;
      RECT 121.18 0.97 121.39 1.323 ;
      RECT 121.146 0.97 121.39 1.321 ;
      RECT 121.06 0.97 121.39 1.315 ;
      RECT 121.015 0.97 121.41 1.293 ;
      RECT 121.015 0.97 121.43 1.248 ;
      RECT 120.975 0.97 121.43 1.238 ;
      RECT 121.185 0.94 121.465 1.22 ;
      RECT 120.92 0.94 121.18 1.2 ;
      RECT 120.105 0.42 120.365 0.68 ;
      RECT 120.185 0.38 120.465 0.66 ;
      RECT 118.745 1.5 119.025 1.78 ;
      RECT 118.715 1.462 118.97 1.765 ;
      RECT 118.71 1.463 118.97 1.763 ;
      RECT 118.705 1.464 118.97 1.757 ;
      RECT 118.7 1.467 118.97 1.75 ;
      RECT 118.695 1.5 119.025 1.743 ;
      RECT 118.665 1.47 118.97 1.73 ;
      RECT 118.665 1.497 118.99 1.73 ;
      RECT 118.665 1.487 118.985 1.73 ;
      RECT 118.665 1.472 118.98 1.73 ;
      RECT 118.745 1.459 118.96 1.78 ;
      RECT 118.831 1.457 118.96 1.78 ;
      RECT 118.917 1.455 118.945 1.78 ;
      RECT 106.075 0.35 106.445 0.72 ;
      RECT 106.59 0.365 106.85 0.69 ;
      RECT 106.075 0.395 106.85 0.655 ;
      RECT 96.86 0.955 97.095 1.215 ;
      RECT 100.005 0.735 100.17 0.995 ;
      RECT 99.91 0.725 99.925 0.995 ;
      RECT 98.51 0.295 98.55 0.435 ;
      RECT 99.925 0.73 100.005 0.995 ;
      RECT 99.87 0.725 99.91 0.961 ;
      RECT 99.856 0.725 99.87 0.961 ;
      RECT 99.77 0.73 99.856 0.963 ;
      RECT 99.725 0.737 99.77 0.965 ;
      RECT 99.695 0.737 99.725 0.967 ;
      RECT 99.67 0.732 99.695 0.969 ;
      RECT 99.64 0.728 99.67 0.978 ;
      RECT 99.63 0.725 99.64 0.99 ;
      RECT 99.625 0.725 99.63 0.998 ;
      RECT 99.62 0.725 99.625 1.003 ;
      RECT 99.61 0.724 99.62 1.013 ;
      RECT 99.605 0.723 99.61 1.023 ;
      RECT 99.59 0.722 99.605 1.028 ;
      RECT 99.562 0.719 99.59 1.055 ;
      RECT 99.476 0.711 99.562 1.055 ;
      RECT 99.39 0.7 99.476 1.055 ;
      RECT 99.35 0.685 99.39 1.055 ;
      RECT 99.31 0.659 99.35 1.055 ;
      RECT 99.305 0.641 99.31 0.867 ;
      RECT 99.295 0.637 99.305 0.857 ;
      RECT 99.28 0.627 99.295 0.844 ;
      RECT 99.26 0.611 99.28 0.829 ;
      RECT 99.245 0.596 99.26 0.814 ;
      RECT 99.235 0.585 99.245 0.804 ;
      RECT 99.21 0.569 99.235 0.793 ;
      RECT 99.205 0.556 99.21 0.783 ;
      RECT 99.2 0.552 99.205 0.778 ;
      RECT 99.145 0.538 99.2 0.756 ;
      RECT 99.106 0.519 99.145 0.72 ;
      RECT 99.02 0.493 99.106 0.673 ;
      RECT 99.016 0.475 99.02 0.639 ;
      RECT 98.93 0.456 99.016 0.617 ;
      RECT 98.925 0.438 98.93 0.595 ;
      RECT 98.92 0.436 98.925 0.593 ;
      RECT 98.91 0.435 98.92 0.588 ;
      RECT 98.85 0.422 98.91 0.574 ;
      RECT 98.805 0.4 98.85 0.553 ;
      RECT 98.745 0.377 98.805 0.532 ;
      RECT 98.681 0.352 98.745 0.507 ;
      RECT 98.595 0.322 98.681 0.476 ;
      RECT 98.58 0.302 98.595 0.455 ;
      RECT 98.55 0.297 98.58 0.446 ;
      RECT 98.497 0.295 98.51 0.435 ;
      RECT 98.411 0.295 98.497 0.437 ;
      RECT 98.325 0.295 98.411 0.439 ;
      RECT 98.305 0.295 98.325 0.443 ;
      RECT 98.26 0.297 98.305 0.454 ;
      RECT 98.22 0.307 98.26 0.47 ;
      RECT 98.216 0.316 98.22 0.478 ;
      RECT 98.13 0.336 98.216 0.494 ;
      RECT 98.12 0.355 98.13 0.512 ;
      RECT 98.115 0.357 98.12 0.515 ;
      RECT 98.105 0.361 98.115 0.518 ;
      RECT 98.085 0.366 98.105 0.528 ;
      RECT 98.055 0.376 98.085 0.548 ;
      RECT 98.05 0.383 98.055 0.562 ;
      RECT 98.04 0.387 98.05 0.569 ;
      RECT 98.025 0.395 98.04 0.58 ;
      RECT 98.015 0.405 98.025 0.591 ;
      RECT 98.005 0.412 98.015 0.599 ;
      RECT 97.98 0.425 98.005 0.614 ;
      RECT 97.916 0.461 97.98 0.653 ;
      RECT 97.83 0.524 97.916 0.717 ;
      RECT 97.795 0.575 97.83 0.77 ;
      RECT 97.79 0.592 97.795 0.787 ;
      RECT 97.775 0.601 97.79 0.794 ;
      RECT 97.755 0.616 97.775 0.808 ;
      RECT 97.75 0.627 97.755 0.818 ;
      RECT 97.73 0.64 97.75 0.828 ;
      RECT 97.725 0.65 97.73 0.838 ;
      RECT 97.71 0.655 97.725 0.847 ;
      RECT 97.7 0.665 97.71 0.858 ;
      RECT 97.67 0.682 97.7 0.875 ;
      RECT 97.66 0.7 97.67 0.893 ;
      RECT 97.645 0.711 97.66 0.904 ;
      RECT 97.605 0.735 97.645 0.92 ;
      RECT 97.57 0.769 97.605 0.937 ;
      RECT 97.54 0.792 97.57 0.949 ;
      RECT 97.525 0.802 97.54 0.958 ;
      RECT 97.485 0.812 97.525 0.969 ;
      RECT 97.465 0.823 97.485 0.981 ;
      RECT 97.46 0.827 97.465 0.988 ;
      RECT 97.445 0.831 97.46 0.993 ;
      RECT 97.435 0.836 97.445 0.998 ;
      RECT 97.43 0.839 97.435 1.001 ;
      RECT 97.4 0.845 97.43 1.008 ;
      RECT 97.365 0.855 97.4 1.022 ;
      RECT 97.305 0.87 97.365 1.042 ;
      RECT 97.25 0.89 97.305 1.066 ;
      RECT 97.221 0.905 97.25 1.084 ;
      RECT 97.135 0.925 97.221 1.109 ;
      RECT 97.13 0.94 97.135 1.129 ;
      RECT 97.12 0.943 97.13 1.13 ;
      RECT 97.095 0.95 97.12 1.215 ;
      RECT 99.79 1.443 100.07 1.78 ;
      RECT 99.79 1.453 100.075 1.738 ;
      RECT 99.79 1.462 100.08 1.635 ;
      RECT 99.79 1.477 100.085 1.503 ;
      RECT 99.79 1.305 100.05 1.78 ;
      RECT 97.51 2.185 97.52 2.375 ;
      RECT 95.77 2.06 96.05 2.34 ;
      RECT 98.815 1 98.82 1.485 ;
      RECT 98.71 1 98.77 1.26 ;
      RECT 99.035 1.97 99.04 2.045 ;
      RECT 99.025 1.837 99.035 2.08 ;
      RECT 99.015 1.672 99.025 2.101 ;
      RECT 99.01 1.542 99.015 2.117 ;
      RECT 99 1.432 99.01 2.133 ;
      RECT 98.995 1.331 99 2.15 ;
      RECT 98.99 1.313 98.995 2.16 ;
      RECT 98.985 1.295 98.99 2.17 ;
      RECT 98.975 1.27 98.985 2.185 ;
      RECT 98.97 1.25 98.975 2.2 ;
      RECT 98.95 1 98.97 2.225 ;
      RECT 98.935 1 98.95 2.258 ;
      RECT 98.905 1 98.935 2.28 ;
      RECT 98.885 1 98.905 2.294 ;
      RECT 98.865 1 98.885 1.81 ;
      RECT 98.88 1.877 98.885 2.299 ;
      RECT 98.875 1.907 98.88 2.301 ;
      RECT 98.87 1.92 98.875 2.304 ;
      RECT 98.865 1.93 98.87 2.308 ;
      RECT 98.86 1 98.865 1.728 ;
      RECT 98.86 1.94 98.865 2.31 ;
      RECT 98.855 1 98.86 1.705 ;
      RECT 98.845 1.962 98.86 2.31 ;
      RECT 98.84 1 98.855 1.65 ;
      RECT 98.835 1.987 98.845 2.31 ;
      RECT 98.835 1 98.84 1.595 ;
      RECT 98.825 1 98.835 1.543 ;
      RECT 98.83 2 98.835 2.311 ;
      RECT 98.825 2.012 98.83 2.312 ;
      RECT 98.82 1 98.825 1.503 ;
      RECT 98.82 2.025 98.825 2.313 ;
      RECT 98.805 2.04 98.82 2.314 ;
      RECT 98.81 1 98.815 1.465 ;
      RECT 98.805 1 98.81 1.43 ;
      RECT 98.8 1 98.805 1.405 ;
      RECT 98.795 2.067 98.805 2.316 ;
      RECT 98.79 1 98.8 1.363 ;
      RECT 98.79 2.085 98.795 2.317 ;
      RECT 98.785 1 98.79 1.323 ;
      RECT 98.785 2.092 98.79 2.318 ;
      RECT 98.78 1 98.785 1.295 ;
      RECT 98.775 2.11 98.785 2.319 ;
      RECT 98.77 1 98.78 1.275 ;
      RECT 98.765 2.13 98.775 2.321 ;
      RECT 98.755 2.147 98.765 2.322 ;
      RECT 98.72 2.17 98.755 2.325 ;
      RECT 98.665 2.188 98.72 2.331 ;
      RECT 98.579 2.196 98.665 2.34 ;
      RECT 98.493 2.207 98.579 2.351 ;
      RECT 98.407 2.217 98.493 2.362 ;
      RECT 98.321 2.227 98.407 2.374 ;
      RECT 98.235 2.237 98.321 2.385 ;
      RECT 98.215 2.243 98.235 2.391 ;
      RECT 98.135 2.245 98.215 2.395 ;
      RECT 98.13 2.244 98.135 2.4 ;
      RECT 98.122 2.243 98.13 2.4 ;
      RECT 98.036 2.239 98.122 2.398 ;
      RECT 97.95 2.231 98.036 2.395 ;
      RECT 97.864 2.222 97.95 2.391 ;
      RECT 97.778 2.214 97.864 2.388 ;
      RECT 97.692 2.206 97.778 2.384 ;
      RECT 97.606 2.197 97.692 2.381 ;
      RECT 97.52 2.189 97.606 2.377 ;
      RECT 97.465 2.182 97.51 2.375 ;
      RECT 97.38 2.175 97.465 2.373 ;
      RECT 97.306 2.167 97.38 2.369 ;
      RECT 97.22 2.159 97.306 2.366 ;
      RECT 97.217 2.155 97.22 2.364 ;
      RECT 97.131 2.151 97.217 2.363 ;
      RECT 97.045 2.143 97.131 2.36 ;
      RECT 96.96 2.138 97.045 2.357 ;
      RECT 96.874 2.135 96.96 2.354 ;
      RECT 96.788 2.133 96.874 2.351 ;
      RECT 96.702 2.13 96.788 2.348 ;
      RECT 96.616 2.127 96.702 2.345 ;
      RECT 96.53 2.124 96.616 2.342 ;
      RECT 96.454 2.122 96.53 2.339 ;
      RECT 96.368 2.119 96.454 2.336 ;
      RECT 96.282 2.116 96.368 2.334 ;
      RECT 96.196 2.114 96.282 2.331 ;
      RECT 96.11 2.111 96.196 2.328 ;
      RECT 96.05 2.102 96.11 2.326 ;
      RECT 98.56 1.72 98.635 1.98 ;
      RECT 98.54 1.7 98.545 1.98 ;
      RECT 97.86 1.485 97.965 1.78 ;
      RECT 92.305 1.46 92.375 1.72 ;
      RECT 98.2 1.335 98.205 1.706 ;
      RECT 98.19 1.39 98.195 1.706 ;
      RECT 98.495 0.56 98.555 0.82 ;
      RECT 98.55 1.715 98.56 1.98 ;
      RECT 98.545 1.705 98.55 1.98 ;
      RECT 98.465 1.652 98.54 1.98 ;
      RECT 98.49 0.56 98.495 0.84 ;
      RECT 98.48 0.56 98.49 0.86 ;
      RECT 98.465 0.56 98.48 0.89 ;
      RECT 98.45 0.56 98.465 0.933 ;
      RECT 98.445 1.595 98.465 1.98 ;
      RECT 98.435 0.56 98.45 0.97 ;
      RECT 98.43 1.575 98.445 1.98 ;
      RECT 98.43 0.56 98.435 0.993 ;
      RECT 98.42 0.56 98.43 1.018 ;
      RECT 98.39 1.542 98.43 1.98 ;
      RECT 98.395 0.56 98.42 1.068 ;
      RECT 98.39 0.56 98.395 1.123 ;
      RECT 98.385 0.56 98.39 1.165 ;
      RECT 98.375 1.505 98.39 1.98 ;
      RECT 98.38 0.56 98.385 1.208 ;
      RECT 98.375 0.56 98.38 1.273 ;
      RECT 98.37 0.56 98.375 1.295 ;
      RECT 98.37 1.493 98.375 1.845 ;
      RECT 98.365 0.56 98.37 1.363 ;
      RECT 98.365 1.485 98.37 1.828 ;
      RECT 98.36 0.56 98.365 1.408 ;
      RECT 98.355 1.467 98.365 1.805 ;
      RECT 98.355 0.56 98.36 1.445 ;
      RECT 98.345 0.56 98.355 1.785 ;
      RECT 98.34 0.56 98.345 1.768 ;
      RECT 98.335 0.56 98.34 1.753 ;
      RECT 98.33 0.56 98.335 1.738 ;
      RECT 98.31 0.56 98.33 1.728 ;
      RECT 98.305 0.56 98.31 1.718 ;
      RECT 98.295 0.56 98.305 1.714 ;
      RECT 98.29 0.837 98.295 1.713 ;
      RECT 98.285 0.86 98.29 1.712 ;
      RECT 98.28 0.89 98.285 1.711 ;
      RECT 98.275 0.917 98.28 1.71 ;
      RECT 98.27 0.945 98.275 1.71 ;
      RECT 98.265 0.972 98.27 1.71 ;
      RECT 98.26 0.992 98.265 1.71 ;
      RECT 98.255 1.02 98.26 1.71 ;
      RECT 98.245 1.062 98.255 1.71 ;
      RECT 98.235 1.107 98.245 1.709 ;
      RECT 98.23 1.16 98.235 1.708 ;
      RECT 98.225 1.192 98.23 1.707 ;
      RECT 98.22 1.212 98.225 1.706 ;
      RECT 98.215 1.25 98.22 1.706 ;
      RECT 98.21 1.272 98.215 1.706 ;
      RECT 98.205 1.297 98.21 1.706 ;
      RECT 98.195 1.362 98.2 1.706 ;
      RECT 98.18 1.422 98.19 1.706 ;
      RECT 98.165 1.432 98.18 1.706 ;
      RECT 98.145 1.442 98.165 1.706 ;
      RECT 98.115 1.447 98.145 1.703 ;
      RECT 98.055 1.457 98.115 1.7 ;
      RECT 98.035 1.466 98.055 1.705 ;
      RECT 98.01 1.472 98.035 1.718 ;
      RECT 97.99 1.477 98.01 1.733 ;
      RECT 97.965 1.482 97.99 1.78 ;
      RECT 97.836 1.484 97.86 1.78 ;
      RECT 97.75 1.479 97.836 1.78 ;
      RECT 97.71 1.476 97.75 1.78 ;
      RECT 97.66 1.478 97.71 1.76 ;
      RECT 97.63 1.482 97.66 1.76 ;
      RECT 97.551 1.492 97.63 1.76 ;
      RECT 97.465 1.507 97.551 1.761 ;
      RECT 97.415 1.517 97.465 1.762 ;
      RECT 97.407 1.52 97.415 1.762 ;
      RECT 97.321 1.522 97.407 1.763 ;
      RECT 97.235 1.526 97.321 1.763 ;
      RECT 97.149 1.53 97.235 1.764 ;
      RECT 97.063 1.533 97.149 1.765 ;
      RECT 96.977 1.537 97.063 1.765 ;
      RECT 96.891 1.541 96.977 1.766 ;
      RECT 96.805 1.544 96.891 1.767 ;
      RECT 96.719 1.548 96.805 1.767 ;
      RECT 96.633 1.552 96.719 1.768 ;
      RECT 96.547 1.556 96.633 1.769 ;
      RECT 96.461 1.559 96.547 1.769 ;
      RECT 96.375 1.563 96.461 1.77 ;
      RECT 96.345 1.565 96.375 1.77 ;
      RECT 96.259 1.568 96.345 1.771 ;
      RECT 96.173 1.572 96.259 1.772 ;
      RECT 96.087 1.576 96.173 1.773 ;
      RECT 96.001 1.579 96.087 1.773 ;
      RECT 95.915 1.583 96.001 1.774 ;
      RECT 95.88 1.588 95.915 1.775 ;
      RECT 95.825 1.598 95.88 1.782 ;
      RECT 95.8 1.61 95.825 1.792 ;
      RECT 95.765 1.623 95.8 1.8 ;
      RECT 95.725 1.64 95.765 1.823 ;
      RECT 95.705 1.653 95.725 1.85 ;
      RECT 95.675 1.665 95.705 1.878 ;
      RECT 95.67 1.673 95.675 1.898 ;
      RECT 95.665 1.676 95.67 1.908 ;
      RECT 95.615 1.688 95.665 1.942 ;
      RECT 95.605 1.703 95.615 1.975 ;
      RECT 95.595 1.709 95.605 1.988 ;
      RECT 95.585 1.716 95.595 2 ;
      RECT 95.56 1.729 95.585 2.018 ;
      RECT 95.545 1.744 95.56 2.04 ;
      RECT 95.535 1.752 95.545 2.056 ;
      RECT 95.52 1.761 95.535 2.071 ;
      RECT 95.51 1.771 95.52 2.085 ;
      RECT 95.491 1.784 95.51 2.102 ;
      RECT 95.405 1.829 95.491 2.167 ;
      RECT 95.39 1.874 95.405 2.225 ;
      RECT 95.385 1.883 95.39 2.238 ;
      RECT 95.375 1.89 95.385 2.243 ;
      RECT 95.37 1.895 95.375 2.247 ;
      RECT 95.35 1.905 95.37 2.254 ;
      RECT 95.325 1.925 95.35 2.268 ;
      RECT 95.29 1.95 95.325 2.288 ;
      RECT 95.275 1.973 95.29 2.303 ;
      RECT 95.265 1.983 95.275 2.308 ;
      RECT 95.255 1.991 95.265 2.315 ;
      RECT 95.245 2 95.255 2.321 ;
      RECT 95.225 2.012 95.245 2.323 ;
      RECT 95.215 2.025 95.225 2.325 ;
      RECT 95.19 2.04 95.215 2.328 ;
      RECT 95.17 2.057 95.19 2.332 ;
      RECT 95.13 2.085 95.17 2.338 ;
      RECT 95.065 2.132 95.13 2.347 ;
      RECT 95.05 2.165 95.065 2.355 ;
      RECT 95.045 2.172 95.05 2.357 ;
      RECT 94.995 2.197 95.045 2.362 ;
      RECT 94.98 2.221 94.995 2.369 ;
      RECT 94.93 2.226 94.98 2.37 ;
      RECT 94.844 2.23 94.93 2.37 ;
      RECT 94.758 2.23 94.844 2.37 ;
      RECT 94.672 2.23 94.758 2.371 ;
      RECT 94.586 2.23 94.672 2.371 ;
      RECT 94.5 2.23 94.586 2.371 ;
      RECT 94.434 2.23 94.5 2.371 ;
      RECT 94.348 2.23 94.434 2.372 ;
      RECT 94.262 2.23 94.348 2.372 ;
      RECT 94.176 2.231 94.262 2.373 ;
      RECT 94.09 2.231 94.176 2.373 ;
      RECT 94.004 2.231 94.09 2.373 ;
      RECT 93.918 2.231 94.004 2.374 ;
      RECT 93.832 2.231 93.918 2.374 ;
      RECT 93.746 2.232 93.832 2.375 ;
      RECT 93.66 2.232 93.746 2.375 ;
      RECT 93.64 2.232 93.66 2.375 ;
      RECT 93.554 2.232 93.64 2.375 ;
      RECT 93.468 2.232 93.554 2.375 ;
      RECT 93.382 2.233 93.468 2.375 ;
      RECT 93.296 2.233 93.382 2.375 ;
      RECT 93.21 2.233 93.296 2.375 ;
      RECT 93.124 2.234 93.21 2.375 ;
      RECT 93.038 2.234 93.124 2.375 ;
      RECT 92.952 2.234 93.038 2.375 ;
      RECT 92.866 2.234 92.952 2.375 ;
      RECT 92.78 2.235 92.866 2.375 ;
      RECT 92.73 2.232 92.78 2.375 ;
      RECT 92.72 2.23 92.73 2.374 ;
      RECT 92.716 2.23 92.72 2.373 ;
      RECT 92.63 2.225 92.716 2.368 ;
      RECT 92.608 2.218 92.63 2.362 ;
      RECT 92.522 2.209 92.608 2.356 ;
      RECT 92.436 2.196 92.522 2.347 ;
      RECT 92.35 2.182 92.436 2.337 ;
      RECT 92.305 2.172 92.35 2.33 ;
      RECT 92.285 1.46 92.305 1.738 ;
      RECT 92.285 2.165 92.305 2.326 ;
      RECT 92.255 1.46 92.285 1.76 ;
      RECT 92.245 2.132 92.285 2.323 ;
      RECT 92.24 1.46 92.255 1.78 ;
      RECT 92.24 2.097 92.245 2.321 ;
      RECT 92.235 1.46 92.24 1.905 ;
      RECT 92.235 2.057 92.24 2.321 ;
      RECT 92.225 1.46 92.235 2.321 ;
      RECT 92.15 1.46 92.225 2.315 ;
      RECT 92.12 1.46 92.15 2.305 ;
      RECT 92.115 1.46 92.12 2.297 ;
      RECT 92.11 1.502 92.115 2.29 ;
      RECT 92.1 1.571 92.11 2.281 ;
      RECT 92.095 1.641 92.1 2.233 ;
      RECT 92.09 1.705 92.095 2.13 ;
      RECT 92.085 1.74 92.09 2.085 ;
      RECT 92.083 1.777 92.085 1.977 ;
      RECT 92.08 1.785 92.083 1.97 ;
      RECT 92.075 1.85 92.08 1.913 ;
      RECT 96.15 0.94 96.43 1.22 ;
      RECT 96.14 0.94 96.43 1.083 ;
      RECT 96.095 0.805 96.355 1.065 ;
      RECT 96.095 0.92 96.41 1.065 ;
      RECT 96.095 0.89 96.405 1.065 ;
      RECT 96.095 0.877 96.395 1.065 ;
      RECT 96.095 0.867 96.39 1.065 ;
      RECT 92.07 0.85 92.33 1.11 ;
      RECT 95.84 0.4 96.1 0.66 ;
      RECT 95.83 0.425 96.1 0.62 ;
      RECT 95.825 0.425 95.83 0.619 ;
      RECT 95.755 0.42 95.825 0.611 ;
      RECT 95.67 0.407 95.755 0.594 ;
      RECT 95.666 0.399 95.67 0.584 ;
      RECT 95.58 0.392 95.666 0.574 ;
      RECT 95.571 0.384 95.58 0.564 ;
      RECT 95.485 0.377 95.571 0.552 ;
      RECT 95.465 0.368 95.485 0.538 ;
      RECT 95.41 0.363 95.465 0.53 ;
      RECT 95.4 0.357 95.41 0.524 ;
      RECT 95.38 0.355 95.4 0.52 ;
      RECT 95.372 0.354 95.38 0.516 ;
      RECT 95.286 0.346 95.372 0.505 ;
      RECT 95.2 0.332 95.286 0.485 ;
      RECT 95.14 0.32 95.2 0.47 ;
      RECT 95.13 0.315 95.14 0.465 ;
      RECT 95.08 0.315 95.13 0.467 ;
      RECT 95.033 0.317 95.08 0.471 ;
      RECT 94.947 0.324 95.033 0.476 ;
      RECT 94.861 0.332 94.947 0.482 ;
      RECT 94.775 0.341 94.861 0.488 ;
      RECT 94.716 0.347 94.775 0.493 ;
      RECT 94.63 0.352 94.716 0.499 ;
      RECT 94.555 0.357 94.63 0.505 ;
      RECT 94.516 0.359 94.555 0.51 ;
      RECT 94.43 0.356 94.516 0.515 ;
      RECT 94.345 0.354 94.43 0.522 ;
      RECT 94.313 0.353 94.345 0.525 ;
      RECT 94.227 0.352 94.313 0.526 ;
      RECT 94.141 0.351 94.227 0.527 ;
      RECT 94.055 0.35 94.141 0.527 ;
      RECT 93.969 0.349 94.055 0.528 ;
      RECT 93.883 0.348 93.969 0.529 ;
      RECT 93.797 0.347 93.883 0.53 ;
      RECT 93.711 0.346 93.797 0.53 ;
      RECT 93.625 0.345 93.711 0.531 ;
      RECT 93.575 0.345 93.625 0.532 ;
      RECT 93.561 0.346 93.575 0.532 ;
      RECT 93.475 0.353 93.561 0.533 ;
      RECT 93.401 0.364 93.475 0.534 ;
      RECT 93.315 0.373 93.401 0.535 ;
      RECT 93.28 0.38 93.315 0.55 ;
      RECT 93.255 0.383 93.28 0.58 ;
      RECT 93.23 0.392 93.255 0.609 ;
      RECT 93.22 0.403 93.23 0.629 ;
      RECT 93.21 0.411 93.22 0.643 ;
      RECT 93.205 0.417 93.21 0.653 ;
      RECT 93.18 0.434 93.205 0.67 ;
      RECT 93.165 0.456 93.18 0.698 ;
      RECT 93.135 0.482 93.165 0.728 ;
      RECT 93.115 0.511 93.135 0.758 ;
      RECT 93.11 0.526 93.115 0.775 ;
      RECT 93.09 0.541 93.11 0.79 ;
      RECT 93.08 0.559 93.09 0.808 ;
      RECT 93.07 0.57 93.08 0.823 ;
      RECT 93.02 0.602 93.07 0.849 ;
      RECT 93.015 0.632 93.02 0.869 ;
      RECT 93.005 0.645 93.015 0.875 ;
      RECT 92.996 0.655 93.005 0.883 ;
      RECT 92.985 0.666 92.996 0.891 ;
      RECT 92.98 0.676 92.985 0.897 ;
      RECT 92.965 0.697 92.98 0.904 ;
      RECT 92.95 0.727 92.965 0.912 ;
      RECT 92.915 0.757 92.95 0.918 ;
      RECT 92.89 0.775 92.915 0.925 ;
      RECT 92.84 0.783 92.89 0.934 ;
      RECT 92.815 0.788 92.84 0.943 ;
      RECT 92.76 0.794 92.815 0.953 ;
      RECT 92.755 0.799 92.76 0.961 ;
      RECT 92.741 0.802 92.755 0.963 ;
      RECT 92.655 0.814 92.741 0.975 ;
      RECT 92.645 0.826 92.655 0.988 ;
      RECT 92.56 0.839 92.645 1 ;
      RECT 92.516 0.856 92.56 1.014 ;
      RECT 92.43 0.873 92.516 1.03 ;
      RECT 92.4 0.887 92.43 1.044 ;
      RECT 92.39 0.892 92.4 1.049 ;
      RECT 92.33 0.895 92.39 1.058 ;
      RECT 95.22 1.165 95.48 1.425 ;
      RECT 95.22 1.165 95.5 1.278 ;
      RECT 95.22 1.165 95.525 1.245 ;
      RECT 95.22 1.165 95.53 1.225 ;
      RECT 95.27 0.94 95.55 1.22 ;
      RECT 94.825 1.675 95.085 1.935 ;
      RECT 94.815 1.532 95.01 1.873 ;
      RECT 94.81 1.64 95.025 1.865 ;
      RECT 94.805 1.69 95.085 1.855 ;
      RECT 94.795 1.767 95.085 1.84 ;
      RECT 94.815 1.615 95.025 1.873 ;
      RECT 94.825 1.49 95.01 1.935 ;
      RECT 94.825 1.385 94.99 1.935 ;
      RECT 94.835 1.372 94.99 1.935 ;
      RECT 94.835 1.33 94.98 1.935 ;
      RECT 94.84 1.255 94.98 1.935 ;
      RECT 94.87 0.905 94.98 1.935 ;
      RECT 94.875 0.635 95 1.258 ;
      RECT 94.845 1.21 95 1.258 ;
      RECT 94.86 1.012 94.98 1.935 ;
      RECT 94.85 1.122 95 1.258 ;
      RECT 94.875 0.635 95.015 1.115 ;
      RECT 94.875 0.635 95.035 0.99 ;
      RECT 94.84 0.635 95.1 0.895 ;
      RECT 94.31 0.94 94.59 1.22 ;
      RECT 94.295 0.94 94.59 1.2 ;
      RECT 92.35 1.805 92.61 2.065 ;
      RECT 94.135 1.66 94.395 1.92 ;
      RECT 94.115 1.68 94.395 1.895 ;
      RECT 94.072 1.68 94.115 1.894 ;
      RECT 93.986 1.681 94.072 1.891 ;
      RECT 93.9 1.682 93.986 1.887 ;
      RECT 93.825 1.684 93.9 1.884 ;
      RECT 93.802 1.685 93.825 1.882 ;
      RECT 93.716 1.686 93.802 1.88 ;
      RECT 93.63 1.687 93.716 1.877 ;
      RECT 93.606 1.688 93.63 1.875 ;
      RECT 93.52 1.69 93.606 1.872 ;
      RECT 93.435 1.692 93.52 1.873 ;
      RECT 93.378 1.693 93.435 1.879 ;
      RECT 93.292 1.695 93.378 1.889 ;
      RECT 93.206 1.698 93.292 1.902 ;
      RECT 93.12 1.7 93.206 1.914 ;
      RECT 93.106 1.701 93.12 1.921 ;
      RECT 93.02 1.702 93.106 1.929 ;
      RECT 92.98 1.704 93.02 1.938 ;
      RECT 92.971 1.705 92.98 1.941 ;
      RECT 92.885 1.713 92.971 1.947 ;
      RECT 92.865 1.722 92.885 1.955 ;
      RECT 92.78 1.737 92.865 1.963 ;
      RECT 92.72 1.76 92.78 1.974 ;
      RECT 92.71 1.772 92.72 1.979 ;
      RECT 92.67 1.782 92.71 1.983 ;
      RECT 92.615 1.799 92.67 1.991 ;
      RECT 92.61 1.809 92.615 1.995 ;
      RECT 93.676 0.94 93.735 1.337 ;
      RECT 93.59 0.94 93.795 1.328 ;
      RECT 93.585 0.97 93.795 1.323 ;
      RECT 93.551 0.97 93.795 1.321 ;
      RECT 93.465 0.97 93.795 1.315 ;
      RECT 93.42 0.97 93.815 1.293 ;
      RECT 93.42 0.97 93.835 1.248 ;
      RECT 93.38 0.97 93.835 1.238 ;
      RECT 93.59 0.94 93.87 1.22 ;
      RECT 93.325 0.94 93.585 1.2 ;
      RECT 92.51 0.42 92.77 0.68 ;
      RECT 92.59 0.38 92.87 0.66 ;
      RECT 91.15 1.5 91.43 1.78 ;
      RECT 91.12 1.462 91.375 1.765 ;
      RECT 91.115 1.463 91.375 1.763 ;
      RECT 91.11 1.464 91.375 1.757 ;
      RECT 91.105 1.467 91.375 1.75 ;
      RECT 91.1 1.5 91.43 1.743 ;
      RECT 91.07 1.47 91.375 1.73 ;
      RECT 91.07 1.497 91.395 1.73 ;
      RECT 91.07 1.487 91.39 1.73 ;
      RECT 91.07 1.472 91.385 1.73 ;
      RECT 91.15 1.459 91.365 1.78 ;
      RECT 91.236 1.457 91.365 1.78 ;
      RECT 91.322 1.455 91.35 1.78 ;
      RECT 78.48 0.35 78.85 0.72 ;
      RECT 78.995 0.365 79.255 0.69 ;
      RECT 78.48 0.395 79.255 0.655 ;
      RECT 69.265 0.955 69.5 1.215 ;
      RECT 72.41 0.735 72.575 0.995 ;
      RECT 72.315 0.725 72.33 0.995 ;
      RECT 70.915 0.295 70.955 0.435 ;
      RECT 72.33 0.73 72.41 0.995 ;
      RECT 72.275 0.725 72.315 0.961 ;
      RECT 72.261 0.725 72.275 0.961 ;
      RECT 72.175 0.73 72.261 0.963 ;
      RECT 72.13 0.737 72.175 0.965 ;
      RECT 72.1 0.737 72.13 0.967 ;
      RECT 72.075 0.732 72.1 0.969 ;
      RECT 72.045 0.728 72.075 0.978 ;
      RECT 72.035 0.725 72.045 0.99 ;
      RECT 72.03 0.725 72.035 0.998 ;
      RECT 72.025 0.725 72.03 1.003 ;
      RECT 72.015 0.724 72.025 1.013 ;
      RECT 72.01 0.723 72.015 1.023 ;
      RECT 71.995 0.722 72.01 1.028 ;
      RECT 71.967 0.719 71.995 1.055 ;
      RECT 71.881 0.711 71.967 1.055 ;
      RECT 71.795 0.7 71.881 1.055 ;
      RECT 71.755 0.685 71.795 1.055 ;
      RECT 71.715 0.659 71.755 1.055 ;
      RECT 71.71 0.641 71.715 0.867 ;
      RECT 71.7 0.637 71.71 0.857 ;
      RECT 71.685 0.627 71.7 0.844 ;
      RECT 71.665 0.611 71.685 0.829 ;
      RECT 71.65 0.596 71.665 0.814 ;
      RECT 71.64 0.585 71.65 0.804 ;
      RECT 71.615 0.569 71.64 0.793 ;
      RECT 71.61 0.556 71.615 0.783 ;
      RECT 71.605 0.552 71.61 0.778 ;
      RECT 71.55 0.538 71.605 0.756 ;
      RECT 71.511 0.519 71.55 0.72 ;
      RECT 71.425 0.493 71.511 0.673 ;
      RECT 71.421 0.475 71.425 0.639 ;
      RECT 71.335 0.456 71.421 0.617 ;
      RECT 71.33 0.438 71.335 0.595 ;
      RECT 71.325 0.436 71.33 0.593 ;
      RECT 71.315 0.435 71.325 0.588 ;
      RECT 71.255 0.422 71.315 0.574 ;
      RECT 71.21 0.4 71.255 0.553 ;
      RECT 71.15 0.377 71.21 0.532 ;
      RECT 71.086 0.352 71.15 0.507 ;
      RECT 71 0.322 71.086 0.476 ;
      RECT 70.985 0.302 71 0.455 ;
      RECT 70.955 0.297 70.985 0.446 ;
      RECT 70.902 0.295 70.915 0.435 ;
      RECT 70.816 0.295 70.902 0.437 ;
      RECT 70.73 0.295 70.816 0.439 ;
      RECT 70.71 0.295 70.73 0.443 ;
      RECT 70.665 0.297 70.71 0.454 ;
      RECT 70.625 0.307 70.665 0.47 ;
      RECT 70.621 0.316 70.625 0.478 ;
      RECT 70.535 0.336 70.621 0.494 ;
      RECT 70.525 0.355 70.535 0.512 ;
      RECT 70.52 0.357 70.525 0.515 ;
      RECT 70.51 0.361 70.52 0.518 ;
      RECT 70.49 0.366 70.51 0.528 ;
      RECT 70.46 0.376 70.49 0.548 ;
      RECT 70.455 0.383 70.46 0.562 ;
      RECT 70.445 0.387 70.455 0.569 ;
      RECT 70.43 0.395 70.445 0.58 ;
      RECT 70.42 0.405 70.43 0.591 ;
      RECT 70.41 0.412 70.42 0.599 ;
      RECT 70.385 0.425 70.41 0.614 ;
      RECT 70.321 0.461 70.385 0.653 ;
      RECT 70.235 0.524 70.321 0.717 ;
      RECT 70.2 0.575 70.235 0.77 ;
      RECT 70.195 0.592 70.2 0.787 ;
      RECT 70.18 0.601 70.195 0.794 ;
      RECT 70.16 0.616 70.18 0.808 ;
      RECT 70.155 0.627 70.16 0.818 ;
      RECT 70.135 0.64 70.155 0.828 ;
      RECT 70.13 0.65 70.135 0.838 ;
      RECT 70.115 0.655 70.13 0.847 ;
      RECT 70.105 0.665 70.115 0.858 ;
      RECT 70.075 0.682 70.105 0.875 ;
      RECT 70.065 0.7 70.075 0.893 ;
      RECT 70.05 0.711 70.065 0.904 ;
      RECT 70.01 0.735 70.05 0.92 ;
      RECT 69.975 0.769 70.01 0.937 ;
      RECT 69.945 0.792 69.975 0.949 ;
      RECT 69.93 0.802 69.945 0.958 ;
      RECT 69.89 0.812 69.93 0.969 ;
      RECT 69.87 0.823 69.89 0.981 ;
      RECT 69.865 0.827 69.87 0.988 ;
      RECT 69.85 0.831 69.865 0.993 ;
      RECT 69.84 0.836 69.85 0.998 ;
      RECT 69.835 0.839 69.84 1.001 ;
      RECT 69.805 0.845 69.835 1.008 ;
      RECT 69.77 0.855 69.805 1.022 ;
      RECT 69.71 0.87 69.77 1.042 ;
      RECT 69.655 0.89 69.71 1.066 ;
      RECT 69.626 0.905 69.655 1.084 ;
      RECT 69.54 0.925 69.626 1.109 ;
      RECT 69.535 0.94 69.54 1.129 ;
      RECT 69.525 0.943 69.535 1.13 ;
      RECT 69.5 0.95 69.525 1.215 ;
      RECT 72.195 1.443 72.475 1.78 ;
      RECT 72.195 1.453 72.48 1.738 ;
      RECT 72.195 1.462 72.485 1.635 ;
      RECT 72.195 1.477 72.49 1.503 ;
      RECT 72.195 1.305 72.455 1.78 ;
      RECT 69.915 2.185 69.925 2.375 ;
      RECT 68.175 2.06 68.455 2.34 ;
      RECT 71.22 1 71.225 1.485 ;
      RECT 71.115 1 71.175 1.26 ;
      RECT 71.44 1.97 71.445 2.045 ;
      RECT 71.43 1.837 71.44 2.08 ;
      RECT 71.42 1.672 71.43 2.101 ;
      RECT 71.415 1.542 71.42 2.117 ;
      RECT 71.405 1.432 71.415 2.133 ;
      RECT 71.4 1.331 71.405 2.15 ;
      RECT 71.395 1.313 71.4 2.16 ;
      RECT 71.39 1.295 71.395 2.17 ;
      RECT 71.38 1.27 71.39 2.185 ;
      RECT 71.375 1.25 71.38 2.2 ;
      RECT 71.355 1 71.375 2.225 ;
      RECT 71.34 1 71.355 2.258 ;
      RECT 71.31 1 71.34 2.28 ;
      RECT 71.29 1 71.31 2.294 ;
      RECT 71.27 1 71.29 1.81 ;
      RECT 71.285 1.877 71.29 2.299 ;
      RECT 71.28 1.907 71.285 2.301 ;
      RECT 71.275 1.92 71.28 2.304 ;
      RECT 71.27 1.93 71.275 2.308 ;
      RECT 71.265 1 71.27 1.728 ;
      RECT 71.265 1.94 71.27 2.31 ;
      RECT 71.26 1 71.265 1.705 ;
      RECT 71.25 1.962 71.265 2.31 ;
      RECT 71.245 1 71.26 1.65 ;
      RECT 71.24 1.987 71.25 2.31 ;
      RECT 71.24 1 71.245 1.595 ;
      RECT 71.23 1 71.24 1.543 ;
      RECT 71.235 2 71.24 2.311 ;
      RECT 71.23 2.012 71.235 2.312 ;
      RECT 71.225 1 71.23 1.503 ;
      RECT 71.225 2.025 71.23 2.313 ;
      RECT 71.21 2.04 71.225 2.314 ;
      RECT 71.215 1 71.22 1.465 ;
      RECT 71.21 1 71.215 1.43 ;
      RECT 71.205 1 71.21 1.405 ;
      RECT 71.2 2.067 71.21 2.316 ;
      RECT 71.195 1 71.205 1.363 ;
      RECT 71.195 2.085 71.2 2.317 ;
      RECT 71.19 1 71.195 1.323 ;
      RECT 71.19 2.092 71.195 2.318 ;
      RECT 71.185 1 71.19 1.295 ;
      RECT 71.18 2.11 71.19 2.319 ;
      RECT 71.175 1 71.185 1.275 ;
      RECT 71.17 2.13 71.18 2.321 ;
      RECT 71.16 2.147 71.17 2.322 ;
      RECT 71.125 2.17 71.16 2.325 ;
      RECT 71.07 2.188 71.125 2.331 ;
      RECT 70.984 2.196 71.07 2.34 ;
      RECT 70.898 2.207 70.984 2.351 ;
      RECT 70.812 2.217 70.898 2.362 ;
      RECT 70.726 2.227 70.812 2.374 ;
      RECT 70.64 2.237 70.726 2.385 ;
      RECT 70.62 2.243 70.64 2.391 ;
      RECT 70.54 2.245 70.62 2.395 ;
      RECT 70.535 2.244 70.54 2.4 ;
      RECT 70.527 2.243 70.535 2.4 ;
      RECT 70.441 2.239 70.527 2.398 ;
      RECT 70.355 2.231 70.441 2.395 ;
      RECT 70.269 2.222 70.355 2.391 ;
      RECT 70.183 2.214 70.269 2.388 ;
      RECT 70.097 2.206 70.183 2.384 ;
      RECT 70.011 2.197 70.097 2.381 ;
      RECT 69.925 2.189 70.011 2.377 ;
      RECT 69.87 2.182 69.915 2.375 ;
      RECT 69.785 2.175 69.87 2.373 ;
      RECT 69.711 2.167 69.785 2.369 ;
      RECT 69.625 2.159 69.711 2.366 ;
      RECT 69.622 2.155 69.625 2.364 ;
      RECT 69.536 2.151 69.622 2.363 ;
      RECT 69.45 2.143 69.536 2.36 ;
      RECT 69.365 2.138 69.45 2.357 ;
      RECT 69.279 2.135 69.365 2.354 ;
      RECT 69.193 2.133 69.279 2.351 ;
      RECT 69.107 2.13 69.193 2.348 ;
      RECT 69.021 2.127 69.107 2.345 ;
      RECT 68.935 2.124 69.021 2.342 ;
      RECT 68.859 2.122 68.935 2.339 ;
      RECT 68.773 2.119 68.859 2.336 ;
      RECT 68.687 2.116 68.773 2.334 ;
      RECT 68.601 2.114 68.687 2.331 ;
      RECT 68.515 2.111 68.601 2.328 ;
      RECT 68.455 2.102 68.515 2.326 ;
      RECT 70.965 1.72 71.04 1.98 ;
      RECT 70.945 1.7 70.95 1.98 ;
      RECT 70.265 1.485 70.37 1.78 ;
      RECT 64.71 1.46 64.78 1.72 ;
      RECT 70.605 1.335 70.61 1.706 ;
      RECT 70.595 1.39 70.6 1.706 ;
      RECT 70.9 0.56 70.96 0.82 ;
      RECT 70.955 1.715 70.965 1.98 ;
      RECT 70.95 1.705 70.955 1.98 ;
      RECT 70.87 1.652 70.945 1.98 ;
      RECT 70.895 0.56 70.9 0.84 ;
      RECT 70.885 0.56 70.895 0.86 ;
      RECT 70.87 0.56 70.885 0.89 ;
      RECT 70.855 0.56 70.87 0.933 ;
      RECT 70.85 1.595 70.87 1.98 ;
      RECT 70.84 0.56 70.855 0.97 ;
      RECT 70.835 1.575 70.85 1.98 ;
      RECT 70.835 0.56 70.84 0.993 ;
      RECT 70.825 0.56 70.835 1.018 ;
      RECT 70.795 1.542 70.835 1.98 ;
      RECT 70.8 0.56 70.825 1.068 ;
      RECT 70.795 0.56 70.8 1.123 ;
      RECT 70.79 0.56 70.795 1.165 ;
      RECT 70.78 1.505 70.795 1.98 ;
      RECT 70.785 0.56 70.79 1.208 ;
      RECT 70.78 0.56 70.785 1.273 ;
      RECT 70.775 0.56 70.78 1.295 ;
      RECT 70.775 1.493 70.78 1.845 ;
      RECT 70.77 0.56 70.775 1.363 ;
      RECT 70.77 1.485 70.775 1.828 ;
      RECT 70.765 0.56 70.77 1.408 ;
      RECT 70.76 1.467 70.77 1.805 ;
      RECT 70.76 0.56 70.765 1.445 ;
      RECT 70.75 0.56 70.76 1.785 ;
      RECT 70.745 0.56 70.75 1.768 ;
      RECT 70.74 0.56 70.745 1.753 ;
      RECT 70.735 0.56 70.74 1.738 ;
      RECT 70.715 0.56 70.735 1.728 ;
      RECT 70.71 0.56 70.715 1.718 ;
      RECT 70.7 0.56 70.71 1.714 ;
      RECT 70.695 0.837 70.7 1.713 ;
      RECT 70.69 0.86 70.695 1.712 ;
      RECT 70.685 0.89 70.69 1.711 ;
      RECT 70.68 0.917 70.685 1.71 ;
      RECT 70.675 0.945 70.68 1.71 ;
      RECT 70.67 0.972 70.675 1.71 ;
      RECT 70.665 0.992 70.67 1.71 ;
      RECT 70.66 1.02 70.665 1.71 ;
      RECT 70.65 1.062 70.66 1.71 ;
      RECT 70.64 1.107 70.65 1.709 ;
      RECT 70.635 1.16 70.64 1.708 ;
      RECT 70.63 1.192 70.635 1.707 ;
      RECT 70.625 1.212 70.63 1.706 ;
      RECT 70.62 1.25 70.625 1.706 ;
      RECT 70.615 1.272 70.62 1.706 ;
      RECT 70.61 1.297 70.615 1.706 ;
      RECT 70.6 1.362 70.605 1.706 ;
      RECT 70.585 1.422 70.595 1.706 ;
      RECT 70.57 1.432 70.585 1.706 ;
      RECT 70.55 1.442 70.57 1.706 ;
      RECT 70.52 1.447 70.55 1.703 ;
      RECT 70.46 1.457 70.52 1.7 ;
      RECT 70.44 1.466 70.46 1.705 ;
      RECT 70.415 1.472 70.44 1.718 ;
      RECT 70.395 1.477 70.415 1.733 ;
      RECT 70.37 1.482 70.395 1.78 ;
      RECT 70.241 1.484 70.265 1.78 ;
      RECT 70.155 1.479 70.241 1.78 ;
      RECT 70.115 1.476 70.155 1.78 ;
      RECT 70.065 1.478 70.115 1.76 ;
      RECT 70.035 1.482 70.065 1.76 ;
      RECT 69.956 1.492 70.035 1.76 ;
      RECT 69.87 1.507 69.956 1.761 ;
      RECT 69.82 1.517 69.87 1.762 ;
      RECT 69.812 1.52 69.82 1.762 ;
      RECT 69.726 1.522 69.812 1.763 ;
      RECT 69.64 1.526 69.726 1.763 ;
      RECT 69.554 1.53 69.64 1.764 ;
      RECT 69.468 1.533 69.554 1.765 ;
      RECT 69.382 1.537 69.468 1.765 ;
      RECT 69.296 1.541 69.382 1.766 ;
      RECT 69.21 1.544 69.296 1.767 ;
      RECT 69.124 1.548 69.21 1.767 ;
      RECT 69.038 1.552 69.124 1.768 ;
      RECT 68.952 1.556 69.038 1.769 ;
      RECT 68.866 1.559 68.952 1.769 ;
      RECT 68.78 1.563 68.866 1.77 ;
      RECT 68.75 1.565 68.78 1.77 ;
      RECT 68.664 1.568 68.75 1.771 ;
      RECT 68.578 1.572 68.664 1.772 ;
      RECT 68.492 1.576 68.578 1.773 ;
      RECT 68.406 1.579 68.492 1.773 ;
      RECT 68.32 1.583 68.406 1.774 ;
      RECT 68.285 1.588 68.32 1.775 ;
      RECT 68.23 1.598 68.285 1.782 ;
      RECT 68.205 1.61 68.23 1.792 ;
      RECT 68.17 1.623 68.205 1.8 ;
      RECT 68.13 1.64 68.17 1.823 ;
      RECT 68.11 1.653 68.13 1.85 ;
      RECT 68.08 1.665 68.11 1.878 ;
      RECT 68.075 1.673 68.08 1.898 ;
      RECT 68.07 1.676 68.075 1.908 ;
      RECT 68.02 1.688 68.07 1.942 ;
      RECT 68.01 1.703 68.02 1.975 ;
      RECT 68 1.709 68.01 1.988 ;
      RECT 67.99 1.716 68 2 ;
      RECT 67.965 1.729 67.99 2.018 ;
      RECT 67.95 1.744 67.965 2.04 ;
      RECT 67.94 1.752 67.95 2.056 ;
      RECT 67.925 1.761 67.94 2.071 ;
      RECT 67.915 1.771 67.925 2.085 ;
      RECT 67.896 1.784 67.915 2.102 ;
      RECT 67.81 1.829 67.896 2.167 ;
      RECT 67.795 1.874 67.81 2.225 ;
      RECT 67.79 1.883 67.795 2.238 ;
      RECT 67.78 1.89 67.79 2.243 ;
      RECT 67.775 1.895 67.78 2.247 ;
      RECT 67.755 1.905 67.775 2.254 ;
      RECT 67.73 1.925 67.755 2.268 ;
      RECT 67.695 1.95 67.73 2.288 ;
      RECT 67.68 1.973 67.695 2.303 ;
      RECT 67.67 1.983 67.68 2.308 ;
      RECT 67.66 1.991 67.67 2.315 ;
      RECT 67.65 2 67.66 2.321 ;
      RECT 67.63 2.012 67.65 2.323 ;
      RECT 67.62 2.025 67.63 2.325 ;
      RECT 67.595 2.04 67.62 2.328 ;
      RECT 67.575 2.057 67.595 2.332 ;
      RECT 67.535 2.085 67.575 2.338 ;
      RECT 67.47 2.132 67.535 2.347 ;
      RECT 67.455 2.165 67.47 2.355 ;
      RECT 67.45 2.172 67.455 2.357 ;
      RECT 67.4 2.197 67.45 2.362 ;
      RECT 67.385 2.221 67.4 2.369 ;
      RECT 67.335 2.226 67.385 2.37 ;
      RECT 67.249 2.23 67.335 2.37 ;
      RECT 67.163 2.23 67.249 2.37 ;
      RECT 67.077 2.23 67.163 2.371 ;
      RECT 66.991 2.23 67.077 2.371 ;
      RECT 66.905 2.23 66.991 2.371 ;
      RECT 66.839 2.23 66.905 2.371 ;
      RECT 66.753 2.23 66.839 2.372 ;
      RECT 66.667 2.23 66.753 2.372 ;
      RECT 66.581 2.231 66.667 2.373 ;
      RECT 66.495 2.231 66.581 2.373 ;
      RECT 66.409 2.231 66.495 2.373 ;
      RECT 66.323 2.231 66.409 2.374 ;
      RECT 66.237 2.231 66.323 2.374 ;
      RECT 66.151 2.232 66.237 2.375 ;
      RECT 66.065 2.232 66.151 2.375 ;
      RECT 66.045 2.232 66.065 2.375 ;
      RECT 65.959 2.232 66.045 2.375 ;
      RECT 65.873 2.232 65.959 2.375 ;
      RECT 65.787 2.233 65.873 2.375 ;
      RECT 65.701 2.233 65.787 2.375 ;
      RECT 65.615 2.233 65.701 2.375 ;
      RECT 65.529 2.234 65.615 2.375 ;
      RECT 65.443 2.234 65.529 2.375 ;
      RECT 65.357 2.234 65.443 2.375 ;
      RECT 65.271 2.234 65.357 2.375 ;
      RECT 65.185 2.235 65.271 2.375 ;
      RECT 65.135 2.232 65.185 2.375 ;
      RECT 65.125 2.23 65.135 2.374 ;
      RECT 65.121 2.23 65.125 2.373 ;
      RECT 65.035 2.225 65.121 2.368 ;
      RECT 65.013 2.218 65.035 2.362 ;
      RECT 64.927 2.209 65.013 2.356 ;
      RECT 64.841 2.196 64.927 2.347 ;
      RECT 64.755 2.182 64.841 2.337 ;
      RECT 64.71 2.172 64.755 2.33 ;
      RECT 64.69 1.46 64.71 1.738 ;
      RECT 64.69 2.165 64.71 2.326 ;
      RECT 64.66 1.46 64.69 1.76 ;
      RECT 64.65 2.132 64.69 2.323 ;
      RECT 64.645 1.46 64.66 1.78 ;
      RECT 64.645 2.097 64.65 2.321 ;
      RECT 64.64 1.46 64.645 1.905 ;
      RECT 64.64 2.057 64.645 2.321 ;
      RECT 64.63 1.46 64.64 2.321 ;
      RECT 64.555 1.46 64.63 2.315 ;
      RECT 64.525 1.46 64.555 2.305 ;
      RECT 64.52 1.46 64.525 2.297 ;
      RECT 64.515 1.502 64.52 2.29 ;
      RECT 64.505 1.571 64.515 2.281 ;
      RECT 64.5 1.641 64.505 2.233 ;
      RECT 64.495 1.705 64.5 2.13 ;
      RECT 64.49 1.74 64.495 2.085 ;
      RECT 64.488 1.777 64.49 1.977 ;
      RECT 64.485 1.785 64.488 1.97 ;
      RECT 64.48 1.85 64.485 1.913 ;
      RECT 68.555 0.94 68.835 1.22 ;
      RECT 68.545 0.94 68.835 1.083 ;
      RECT 68.5 0.805 68.76 1.065 ;
      RECT 68.5 0.92 68.815 1.065 ;
      RECT 68.5 0.89 68.81 1.065 ;
      RECT 68.5 0.877 68.8 1.065 ;
      RECT 68.5 0.867 68.795 1.065 ;
      RECT 64.475 0.85 64.735 1.11 ;
      RECT 68.245 0.4 68.505 0.66 ;
      RECT 68.235 0.425 68.505 0.62 ;
      RECT 68.23 0.425 68.235 0.619 ;
      RECT 68.16 0.42 68.23 0.611 ;
      RECT 68.075 0.407 68.16 0.594 ;
      RECT 68.071 0.399 68.075 0.584 ;
      RECT 67.985 0.392 68.071 0.574 ;
      RECT 67.976 0.384 67.985 0.564 ;
      RECT 67.89 0.377 67.976 0.552 ;
      RECT 67.87 0.368 67.89 0.538 ;
      RECT 67.815 0.363 67.87 0.53 ;
      RECT 67.805 0.357 67.815 0.524 ;
      RECT 67.785 0.355 67.805 0.52 ;
      RECT 67.777 0.354 67.785 0.516 ;
      RECT 67.691 0.346 67.777 0.505 ;
      RECT 67.605 0.332 67.691 0.485 ;
      RECT 67.545 0.32 67.605 0.47 ;
      RECT 67.535 0.315 67.545 0.465 ;
      RECT 67.485 0.315 67.535 0.467 ;
      RECT 67.438 0.317 67.485 0.471 ;
      RECT 67.352 0.324 67.438 0.476 ;
      RECT 67.266 0.332 67.352 0.482 ;
      RECT 67.18 0.341 67.266 0.488 ;
      RECT 67.121 0.347 67.18 0.493 ;
      RECT 67.035 0.352 67.121 0.499 ;
      RECT 66.96 0.357 67.035 0.505 ;
      RECT 66.921 0.359 66.96 0.51 ;
      RECT 66.835 0.356 66.921 0.515 ;
      RECT 66.75 0.354 66.835 0.522 ;
      RECT 66.718 0.353 66.75 0.525 ;
      RECT 66.632 0.352 66.718 0.526 ;
      RECT 66.546 0.351 66.632 0.527 ;
      RECT 66.46 0.35 66.546 0.527 ;
      RECT 66.374 0.349 66.46 0.528 ;
      RECT 66.288 0.348 66.374 0.529 ;
      RECT 66.202 0.347 66.288 0.53 ;
      RECT 66.116 0.346 66.202 0.53 ;
      RECT 66.03 0.345 66.116 0.531 ;
      RECT 65.98 0.345 66.03 0.532 ;
      RECT 65.966 0.346 65.98 0.532 ;
      RECT 65.88 0.353 65.966 0.533 ;
      RECT 65.806 0.364 65.88 0.534 ;
      RECT 65.72 0.373 65.806 0.535 ;
      RECT 65.685 0.38 65.72 0.55 ;
      RECT 65.66 0.383 65.685 0.58 ;
      RECT 65.635 0.392 65.66 0.609 ;
      RECT 65.625 0.403 65.635 0.629 ;
      RECT 65.615 0.411 65.625 0.643 ;
      RECT 65.61 0.417 65.615 0.653 ;
      RECT 65.585 0.434 65.61 0.67 ;
      RECT 65.57 0.456 65.585 0.698 ;
      RECT 65.54 0.482 65.57 0.728 ;
      RECT 65.52 0.511 65.54 0.758 ;
      RECT 65.515 0.526 65.52 0.775 ;
      RECT 65.495 0.541 65.515 0.79 ;
      RECT 65.485 0.559 65.495 0.808 ;
      RECT 65.475 0.57 65.485 0.823 ;
      RECT 65.425 0.602 65.475 0.849 ;
      RECT 65.42 0.632 65.425 0.869 ;
      RECT 65.41 0.645 65.42 0.875 ;
      RECT 65.401 0.655 65.41 0.883 ;
      RECT 65.39 0.666 65.401 0.891 ;
      RECT 65.385 0.676 65.39 0.897 ;
      RECT 65.37 0.697 65.385 0.904 ;
      RECT 65.355 0.727 65.37 0.912 ;
      RECT 65.32 0.757 65.355 0.918 ;
      RECT 65.295 0.775 65.32 0.925 ;
      RECT 65.245 0.783 65.295 0.934 ;
      RECT 65.22 0.788 65.245 0.943 ;
      RECT 65.165 0.794 65.22 0.953 ;
      RECT 65.16 0.799 65.165 0.961 ;
      RECT 65.146 0.802 65.16 0.963 ;
      RECT 65.06 0.814 65.146 0.975 ;
      RECT 65.05 0.826 65.06 0.988 ;
      RECT 64.965 0.839 65.05 1 ;
      RECT 64.921 0.856 64.965 1.014 ;
      RECT 64.835 0.873 64.921 1.03 ;
      RECT 64.805 0.887 64.835 1.044 ;
      RECT 64.795 0.892 64.805 1.049 ;
      RECT 64.735 0.895 64.795 1.058 ;
      RECT 67.625 1.165 67.885 1.425 ;
      RECT 67.625 1.165 67.905 1.278 ;
      RECT 67.625 1.165 67.93 1.245 ;
      RECT 67.625 1.165 67.935 1.225 ;
      RECT 67.675 0.94 67.955 1.22 ;
      RECT 67.23 1.675 67.49 1.935 ;
      RECT 67.22 1.532 67.415 1.873 ;
      RECT 67.215 1.64 67.43 1.865 ;
      RECT 67.21 1.69 67.49 1.855 ;
      RECT 67.2 1.767 67.49 1.84 ;
      RECT 67.22 1.615 67.43 1.873 ;
      RECT 67.23 1.49 67.415 1.935 ;
      RECT 67.23 1.385 67.395 1.935 ;
      RECT 67.24 1.372 67.395 1.935 ;
      RECT 67.24 1.33 67.385 1.935 ;
      RECT 67.245 1.255 67.385 1.935 ;
      RECT 67.275 0.905 67.385 1.935 ;
      RECT 67.28 0.635 67.405 1.258 ;
      RECT 67.25 1.21 67.405 1.258 ;
      RECT 67.265 1.012 67.385 1.935 ;
      RECT 67.255 1.122 67.405 1.258 ;
      RECT 67.28 0.635 67.42 1.115 ;
      RECT 67.28 0.635 67.44 0.99 ;
      RECT 67.245 0.635 67.505 0.895 ;
      RECT 66.715 0.94 66.995 1.22 ;
      RECT 66.7 0.94 66.995 1.2 ;
      RECT 64.755 1.805 65.015 2.065 ;
      RECT 66.54 1.66 66.8 1.92 ;
      RECT 66.52 1.68 66.8 1.895 ;
      RECT 66.477 1.68 66.52 1.894 ;
      RECT 66.391 1.681 66.477 1.891 ;
      RECT 66.305 1.682 66.391 1.887 ;
      RECT 66.23 1.684 66.305 1.884 ;
      RECT 66.207 1.685 66.23 1.882 ;
      RECT 66.121 1.686 66.207 1.88 ;
      RECT 66.035 1.687 66.121 1.877 ;
      RECT 66.011 1.688 66.035 1.875 ;
      RECT 65.925 1.69 66.011 1.872 ;
      RECT 65.84 1.692 65.925 1.873 ;
      RECT 65.783 1.693 65.84 1.879 ;
      RECT 65.697 1.695 65.783 1.889 ;
      RECT 65.611 1.698 65.697 1.902 ;
      RECT 65.525 1.7 65.611 1.914 ;
      RECT 65.511 1.701 65.525 1.921 ;
      RECT 65.425 1.702 65.511 1.929 ;
      RECT 65.385 1.704 65.425 1.938 ;
      RECT 65.376 1.705 65.385 1.941 ;
      RECT 65.29 1.713 65.376 1.947 ;
      RECT 65.27 1.722 65.29 1.955 ;
      RECT 65.185 1.737 65.27 1.963 ;
      RECT 65.125 1.76 65.185 1.974 ;
      RECT 65.115 1.772 65.125 1.979 ;
      RECT 65.075 1.782 65.115 1.983 ;
      RECT 65.02 1.799 65.075 1.991 ;
      RECT 65.015 1.809 65.02 1.995 ;
      RECT 66.081 0.94 66.14 1.337 ;
      RECT 65.995 0.94 66.2 1.328 ;
      RECT 65.99 0.97 66.2 1.323 ;
      RECT 65.956 0.97 66.2 1.321 ;
      RECT 65.87 0.97 66.2 1.315 ;
      RECT 65.825 0.97 66.22 1.293 ;
      RECT 65.825 0.97 66.24 1.248 ;
      RECT 65.785 0.97 66.24 1.238 ;
      RECT 65.995 0.94 66.275 1.22 ;
      RECT 65.73 0.94 65.99 1.2 ;
      RECT 64.915 0.42 65.175 0.68 ;
      RECT 64.995 0.38 65.275 0.66 ;
      RECT 63.555 1.5 63.835 1.78 ;
      RECT 63.525 1.462 63.78 1.765 ;
      RECT 63.52 1.463 63.78 1.763 ;
      RECT 63.515 1.464 63.78 1.757 ;
      RECT 63.51 1.467 63.78 1.75 ;
      RECT 63.505 1.5 63.835 1.743 ;
      RECT 63.475 1.47 63.78 1.73 ;
      RECT 63.475 1.497 63.8 1.73 ;
      RECT 63.475 1.487 63.795 1.73 ;
      RECT 63.475 1.472 63.79 1.73 ;
      RECT 63.555 1.459 63.77 1.78 ;
      RECT 63.641 1.457 63.77 1.78 ;
      RECT 63.727 1.455 63.755 1.78 ;
      RECT 50.885 0.35 51.255 0.72 ;
      RECT 51.4 0.365 51.66 0.69 ;
      RECT 50.885 0.395 51.66 0.655 ;
      RECT 41.67 0.955 41.905 1.215 ;
      RECT 44.815 0.735 44.98 0.995 ;
      RECT 44.72 0.725 44.735 0.995 ;
      RECT 43.32 0.295 43.36 0.435 ;
      RECT 44.735 0.73 44.815 0.995 ;
      RECT 44.68 0.725 44.72 0.961 ;
      RECT 44.666 0.725 44.68 0.961 ;
      RECT 44.58 0.73 44.666 0.963 ;
      RECT 44.535 0.737 44.58 0.965 ;
      RECT 44.505 0.737 44.535 0.967 ;
      RECT 44.48 0.732 44.505 0.969 ;
      RECT 44.45 0.728 44.48 0.978 ;
      RECT 44.44 0.725 44.45 0.99 ;
      RECT 44.435 0.725 44.44 0.998 ;
      RECT 44.43 0.725 44.435 1.003 ;
      RECT 44.42 0.724 44.43 1.013 ;
      RECT 44.415 0.723 44.42 1.023 ;
      RECT 44.4 0.722 44.415 1.028 ;
      RECT 44.372 0.719 44.4 1.055 ;
      RECT 44.286 0.711 44.372 1.055 ;
      RECT 44.2 0.7 44.286 1.055 ;
      RECT 44.16 0.685 44.2 1.055 ;
      RECT 44.12 0.659 44.16 1.055 ;
      RECT 44.115 0.641 44.12 0.867 ;
      RECT 44.105 0.637 44.115 0.857 ;
      RECT 44.09 0.627 44.105 0.844 ;
      RECT 44.07 0.611 44.09 0.829 ;
      RECT 44.055 0.596 44.07 0.814 ;
      RECT 44.045 0.585 44.055 0.804 ;
      RECT 44.02 0.569 44.045 0.793 ;
      RECT 44.015 0.556 44.02 0.783 ;
      RECT 44.01 0.552 44.015 0.778 ;
      RECT 43.955 0.538 44.01 0.756 ;
      RECT 43.916 0.519 43.955 0.72 ;
      RECT 43.83 0.493 43.916 0.673 ;
      RECT 43.826 0.475 43.83 0.639 ;
      RECT 43.74 0.456 43.826 0.617 ;
      RECT 43.735 0.438 43.74 0.595 ;
      RECT 43.73 0.436 43.735 0.593 ;
      RECT 43.72 0.435 43.73 0.588 ;
      RECT 43.66 0.422 43.72 0.574 ;
      RECT 43.615 0.4 43.66 0.553 ;
      RECT 43.555 0.377 43.615 0.532 ;
      RECT 43.491 0.352 43.555 0.507 ;
      RECT 43.405 0.322 43.491 0.476 ;
      RECT 43.39 0.302 43.405 0.455 ;
      RECT 43.36 0.297 43.39 0.446 ;
      RECT 43.307 0.295 43.32 0.435 ;
      RECT 43.221 0.295 43.307 0.437 ;
      RECT 43.135 0.295 43.221 0.439 ;
      RECT 43.115 0.295 43.135 0.443 ;
      RECT 43.07 0.297 43.115 0.454 ;
      RECT 43.03 0.307 43.07 0.47 ;
      RECT 43.026 0.316 43.03 0.478 ;
      RECT 42.94 0.336 43.026 0.494 ;
      RECT 42.93 0.355 42.94 0.512 ;
      RECT 42.925 0.357 42.93 0.515 ;
      RECT 42.915 0.361 42.925 0.518 ;
      RECT 42.895 0.366 42.915 0.528 ;
      RECT 42.865 0.376 42.895 0.548 ;
      RECT 42.86 0.383 42.865 0.562 ;
      RECT 42.85 0.387 42.86 0.569 ;
      RECT 42.835 0.395 42.85 0.58 ;
      RECT 42.825 0.405 42.835 0.591 ;
      RECT 42.815 0.412 42.825 0.599 ;
      RECT 42.79 0.425 42.815 0.614 ;
      RECT 42.726 0.461 42.79 0.653 ;
      RECT 42.64 0.524 42.726 0.717 ;
      RECT 42.605 0.575 42.64 0.77 ;
      RECT 42.6 0.592 42.605 0.787 ;
      RECT 42.585 0.601 42.6 0.794 ;
      RECT 42.565 0.616 42.585 0.808 ;
      RECT 42.56 0.627 42.565 0.818 ;
      RECT 42.54 0.64 42.56 0.828 ;
      RECT 42.535 0.65 42.54 0.838 ;
      RECT 42.52 0.655 42.535 0.847 ;
      RECT 42.51 0.665 42.52 0.858 ;
      RECT 42.48 0.682 42.51 0.875 ;
      RECT 42.47 0.7 42.48 0.893 ;
      RECT 42.455 0.711 42.47 0.904 ;
      RECT 42.415 0.735 42.455 0.92 ;
      RECT 42.38 0.769 42.415 0.937 ;
      RECT 42.35 0.792 42.38 0.949 ;
      RECT 42.335 0.802 42.35 0.958 ;
      RECT 42.295 0.812 42.335 0.969 ;
      RECT 42.275 0.823 42.295 0.981 ;
      RECT 42.27 0.827 42.275 0.988 ;
      RECT 42.255 0.831 42.27 0.993 ;
      RECT 42.245 0.836 42.255 0.998 ;
      RECT 42.24 0.839 42.245 1.001 ;
      RECT 42.21 0.845 42.24 1.008 ;
      RECT 42.175 0.855 42.21 1.022 ;
      RECT 42.115 0.87 42.175 1.042 ;
      RECT 42.06 0.89 42.115 1.066 ;
      RECT 42.031 0.905 42.06 1.084 ;
      RECT 41.945 0.925 42.031 1.109 ;
      RECT 41.94 0.94 41.945 1.129 ;
      RECT 41.93 0.943 41.94 1.13 ;
      RECT 41.905 0.95 41.93 1.215 ;
      RECT 44.6 1.443 44.88 1.78 ;
      RECT 44.6 1.453 44.885 1.738 ;
      RECT 44.6 1.462 44.89 1.635 ;
      RECT 44.6 1.477 44.895 1.503 ;
      RECT 44.6 1.305 44.86 1.78 ;
      RECT 42.32 2.185 42.33 2.375 ;
      RECT 40.58 2.06 40.86 2.34 ;
      RECT 43.625 1 43.63 1.485 ;
      RECT 43.52 1 43.58 1.26 ;
      RECT 43.845 1.97 43.85 2.045 ;
      RECT 43.835 1.837 43.845 2.08 ;
      RECT 43.825 1.672 43.835 2.101 ;
      RECT 43.82 1.542 43.825 2.117 ;
      RECT 43.81 1.432 43.82 2.133 ;
      RECT 43.805 1.331 43.81 2.15 ;
      RECT 43.8 1.313 43.805 2.16 ;
      RECT 43.795 1.295 43.8 2.17 ;
      RECT 43.785 1.27 43.795 2.185 ;
      RECT 43.78 1.25 43.785 2.2 ;
      RECT 43.76 1 43.78 2.225 ;
      RECT 43.745 1 43.76 2.258 ;
      RECT 43.715 1 43.745 2.28 ;
      RECT 43.695 1 43.715 2.294 ;
      RECT 43.675 1 43.695 1.81 ;
      RECT 43.69 1.877 43.695 2.299 ;
      RECT 43.685 1.907 43.69 2.301 ;
      RECT 43.68 1.92 43.685 2.304 ;
      RECT 43.675 1.93 43.68 2.308 ;
      RECT 43.67 1 43.675 1.728 ;
      RECT 43.67 1.94 43.675 2.31 ;
      RECT 43.665 1 43.67 1.705 ;
      RECT 43.655 1.962 43.67 2.31 ;
      RECT 43.65 1 43.665 1.65 ;
      RECT 43.645 1.987 43.655 2.31 ;
      RECT 43.645 1 43.65 1.595 ;
      RECT 43.635 1 43.645 1.543 ;
      RECT 43.64 2 43.645 2.311 ;
      RECT 43.635 2.012 43.64 2.312 ;
      RECT 43.63 1 43.635 1.503 ;
      RECT 43.63 2.025 43.635 2.313 ;
      RECT 43.615 2.04 43.63 2.314 ;
      RECT 43.62 1 43.625 1.465 ;
      RECT 43.615 1 43.62 1.43 ;
      RECT 43.61 1 43.615 1.405 ;
      RECT 43.605 2.067 43.615 2.316 ;
      RECT 43.6 1 43.61 1.363 ;
      RECT 43.6 2.085 43.605 2.317 ;
      RECT 43.595 1 43.6 1.323 ;
      RECT 43.595 2.092 43.6 2.318 ;
      RECT 43.59 1 43.595 1.295 ;
      RECT 43.585 2.11 43.595 2.319 ;
      RECT 43.58 1 43.59 1.275 ;
      RECT 43.575 2.13 43.585 2.321 ;
      RECT 43.565 2.147 43.575 2.322 ;
      RECT 43.53 2.17 43.565 2.325 ;
      RECT 43.475 2.188 43.53 2.331 ;
      RECT 43.389 2.196 43.475 2.34 ;
      RECT 43.303 2.207 43.389 2.351 ;
      RECT 43.217 2.217 43.303 2.362 ;
      RECT 43.131 2.227 43.217 2.374 ;
      RECT 43.045 2.237 43.131 2.385 ;
      RECT 43.025 2.243 43.045 2.391 ;
      RECT 42.945 2.245 43.025 2.395 ;
      RECT 42.94 2.244 42.945 2.4 ;
      RECT 42.932 2.243 42.94 2.4 ;
      RECT 42.846 2.239 42.932 2.398 ;
      RECT 42.76 2.231 42.846 2.395 ;
      RECT 42.674 2.222 42.76 2.391 ;
      RECT 42.588 2.214 42.674 2.388 ;
      RECT 42.502 2.206 42.588 2.384 ;
      RECT 42.416 2.197 42.502 2.381 ;
      RECT 42.33 2.189 42.416 2.377 ;
      RECT 42.275 2.182 42.32 2.375 ;
      RECT 42.19 2.175 42.275 2.373 ;
      RECT 42.116 2.167 42.19 2.369 ;
      RECT 42.03 2.159 42.116 2.366 ;
      RECT 42.027 2.155 42.03 2.364 ;
      RECT 41.941 2.151 42.027 2.363 ;
      RECT 41.855 2.143 41.941 2.36 ;
      RECT 41.77 2.138 41.855 2.357 ;
      RECT 41.684 2.135 41.77 2.354 ;
      RECT 41.598 2.133 41.684 2.351 ;
      RECT 41.512 2.13 41.598 2.348 ;
      RECT 41.426 2.127 41.512 2.345 ;
      RECT 41.34 2.124 41.426 2.342 ;
      RECT 41.264 2.122 41.34 2.339 ;
      RECT 41.178 2.119 41.264 2.336 ;
      RECT 41.092 2.116 41.178 2.334 ;
      RECT 41.006 2.114 41.092 2.331 ;
      RECT 40.92 2.111 41.006 2.328 ;
      RECT 40.86 2.102 40.92 2.326 ;
      RECT 43.37 1.72 43.445 1.98 ;
      RECT 43.35 1.7 43.355 1.98 ;
      RECT 42.67 1.485 42.775 1.78 ;
      RECT 37.115 1.46 37.185 1.72 ;
      RECT 43.01 1.335 43.015 1.706 ;
      RECT 43 1.39 43.005 1.706 ;
      RECT 43.305 0.56 43.365 0.82 ;
      RECT 43.36 1.715 43.37 1.98 ;
      RECT 43.355 1.705 43.36 1.98 ;
      RECT 43.275 1.652 43.35 1.98 ;
      RECT 43.3 0.56 43.305 0.84 ;
      RECT 43.29 0.56 43.3 0.86 ;
      RECT 43.275 0.56 43.29 0.89 ;
      RECT 43.26 0.56 43.275 0.933 ;
      RECT 43.255 1.595 43.275 1.98 ;
      RECT 43.245 0.56 43.26 0.97 ;
      RECT 43.24 1.575 43.255 1.98 ;
      RECT 43.24 0.56 43.245 0.993 ;
      RECT 43.23 0.56 43.24 1.018 ;
      RECT 43.2 1.542 43.24 1.98 ;
      RECT 43.205 0.56 43.23 1.068 ;
      RECT 43.2 0.56 43.205 1.123 ;
      RECT 43.195 0.56 43.2 1.165 ;
      RECT 43.185 1.505 43.2 1.98 ;
      RECT 43.19 0.56 43.195 1.208 ;
      RECT 43.185 0.56 43.19 1.273 ;
      RECT 43.18 0.56 43.185 1.295 ;
      RECT 43.18 1.493 43.185 1.845 ;
      RECT 43.175 0.56 43.18 1.363 ;
      RECT 43.175 1.485 43.18 1.828 ;
      RECT 43.17 0.56 43.175 1.408 ;
      RECT 43.165 1.467 43.175 1.805 ;
      RECT 43.165 0.56 43.17 1.445 ;
      RECT 43.155 0.56 43.165 1.785 ;
      RECT 43.15 0.56 43.155 1.768 ;
      RECT 43.145 0.56 43.15 1.753 ;
      RECT 43.14 0.56 43.145 1.738 ;
      RECT 43.12 0.56 43.14 1.728 ;
      RECT 43.115 0.56 43.12 1.718 ;
      RECT 43.105 0.56 43.115 1.714 ;
      RECT 43.1 0.837 43.105 1.713 ;
      RECT 43.095 0.86 43.1 1.712 ;
      RECT 43.09 0.89 43.095 1.711 ;
      RECT 43.085 0.917 43.09 1.71 ;
      RECT 43.08 0.945 43.085 1.71 ;
      RECT 43.075 0.972 43.08 1.71 ;
      RECT 43.07 0.992 43.075 1.71 ;
      RECT 43.065 1.02 43.07 1.71 ;
      RECT 43.055 1.062 43.065 1.71 ;
      RECT 43.045 1.107 43.055 1.709 ;
      RECT 43.04 1.16 43.045 1.708 ;
      RECT 43.035 1.192 43.04 1.707 ;
      RECT 43.03 1.212 43.035 1.706 ;
      RECT 43.025 1.25 43.03 1.706 ;
      RECT 43.02 1.272 43.025 1.706 ;
      RECT 43.015 1.297 43.02 1.706 ;
      RECT 43.005 1.362 43.01 1.706 ;
      RECT 42.99 1.422 43 1.706 ;
      RECT 42.975 1.432 42.99 1.706 ;
      RECT 42.955 1.442 42.975 1.706 ;
      RECT 42.925 1.447 42.955 1.703 ;
      RECT 42.865 1.457 42.925 1.7 ;
      RECT 42.845 1.466 42.865 1.705 ;
      RECT 42.82 1.472 42.845 1.718 ;
      RECT 42.8 1.477 42.82 1.733 ;
      RECT 42.775 1.482 42.8 1.78 ;
      RECT 42.646 1.484 42.67 1.78 ;
      RECT 42.56 1.479 42.646 1.78 ;
      RECT 42.52 1.476 42.56 1.78 ;
      RECT 42.47 1.478 42.52 1.76 ;
      RECT 42.44 1.482 42.47 1.76 ;
      RECT 42.361 1.492 42.44 1.76 ;
      RECT 42.275 1.507 42.361 1.761 ;
      RECT 42.225 1.517 42.275 1.762 ;
      RECT 42.217 1.52 42.225 1.762 ;
      RECT 42.131 1.522 42.217 1.763 ;
      RECT 42.045 1.526 42.131 1.763 ;
      RECT 41.959 1.53 42.045 1.764 ;
      RECT 41.873 1.533 41.959 1.765 ;
      RECT 41.787 1.537 41.873 1.765 ;
      RECT 41.701 1.541 41.787 1.766 ;
      RECT 41.615 1.544 41.701 1.767 ;
      RECT 41.529 1.548 41.615 1.767 ;
      RECT 41.443 1.552 41.529 1.768 ;
      RECT 41.357 1.556 41.443 1.769 ;
      RECT 41.271 1.559 41.357 1.769 ;
      RECT 41.185 1.563 41.271 1.77 ;
      RECT 41.155 1.565 41.185 1.77 ;
      RECT 41.069 1.568 41.155 1.771 ;
      RECT 40.983 1.572 41.069 1.772 ;
      RECT 40.897 1.576 40.983 1.773 ;
      RECT 40.811 1.579 40.897 1.773 ;
      RECT 40.725 1.583 40.811 1.774 ;
      RECT 40.69 1.588 40.725 1.775 ;
      RECT 40.635 1.598 40.69 1.782 ;
      RECT 40.61 1.61 40.635 1.792 ;
      RECT 40.575 1.623 40.61 1.8 ;
      RECT 40.535 1.64 40.575 1.823 ;
      RECT 40.515 1.653 40.535 1.85 ;
      RECT 40.485 1.665 40.515 1.878 ;
      RECT 40.48 1.673 40.485 1.898 ;
      RECT 40.475 1.676 40.48 1.908 ;
      RECT 40.425 1.688 40.475 1.942 ;
      RECT 40.415 1.703 40.425 1.975 ;
      RECT 40.405 1.709 40.415 1.988 ;
      RECT 40.395 1.716 40.405 2 ;
      RECT 40.37 1.729 40.395 2.018 ;
      RECT 40.355 1.744 40.37 2.04 ;
      RECT 40.345 1.752 40.355 2.056 ;
      RECT 40.33 1.761 40.345 2.071 ;
      RECT 40.32 1.771 40.33 2.085 ;
      RECT 40.301 1.784 40.32 2.102 ;
      RECT 40.215 1.829 40.301 2.167 ;
      RECT 40.2 1.874 40.215 2.225 ;
      RECT 40.195 1.883 40.2 2.238 ;
      RECT 40.185 1.89 40.195 2.243 ;
      RECT 40.18 1.895 40.185 2.247 ;
      RECT 40.16 1.905 40.18 2.254 ;
      RECT 40.135 1.925 40.16 2.268 ;
      RECT 40.1 1.95 40.135 2.288 ;
      RECT 40.085 1.973 40.1 2.303 ;
      RECT 40.075 1.983 40.085 2.308 ;
      RECT 40.065 1.991 40.075 2.315 ;
      RECT 40.055 2 40.065 2.321 ;
      RECT 40.035 2.012 40.055 2.323 ;
      RECT 40.025 2.025 40.035 2.325 ;
      RECT 40 2.04 40.025 2.328 ;
      RECT 39.98 2.057 40 2.332 ;
      RECT 39.94 2.085 39.98 2.338 ;
      RECT 39.875 2.132 39.94 2.347 ;
      RECT 39.86 2.165 39.875 2.355 ;
      RECT 39.855 2.172 39.86 2.357 ;
      RECT 39.805 2.197 39.855 2.362 ;
      RECT 39.79 2.221 39.805 2.369 ;
      RECT 39.74 2.226 39.79 2.37 ;
      RECT 39.654 2.23 39.74 2.37 ;
      RECT 39.568 2.23 39.654 2.37 ;
      RECT 39.482 2.23 39.568 2.371 ;
      RECT 39.396 2.23 39.482 2.371 ;
      RECT 39.31 2.23 39.396 2.371 ;
      RECT 39.244 2.23 39.31 2.371 ;
      RECT 39.158 2.23 39.244 2.372 ;
      RECT 39.072 2.23 39.158 2.372 ;
      RECT 38.986 2.231 39.072 2.373 ;
      RECT 38.9 2.231 38.986 2.373 ;
      RECT 38.814 2.231 38.9 2.373 ;
      RECT 38.728 2.231 38.814 2.374 ;
      RECT 38.642 2.231 38.728 2.374 ;
      RECT 38.556 2.232 38.642 2.375 ;
      RECT 38.47 2.232 38.556 2.375 ;
      RECT 38.45 2.232 38.47 2.375 ;
      RECT 38.364 2.232 38.45 2.375 ;
      RECT 38.278 2.232 38.364 2.375 ;
      RECT 38.192 2.233 38.278 2.375 ;
      RECT 38.106 2.233 38.192 2.375 ;
      RECT 38.02 2.233 38.106 2.375 ;
      RECT 37.934 2.234 38.02 2.375 ;
      RECT 37.848 2.234 37.934 2.375 ;
      RECT 37.762 2.234 37.848 2.375 ;
      RECT 37.676 2.234 37.762 2.375 ;
      RECT 37.59 2.235 37.676 2.375 ;
      RECT 37.54 2.232 37.59 2.375 ;
      RECT 37.53 2.23 37.54 2.374 ;
      RECT 37.526 2.23 37.53 2.373 ;
      RECT 37.44 2.225 37.526 2.368 ;
      RECT 37.418 2.218 37.44 2.362 ;
      RECT 37.332 2.209 37.418 2.356 ;
      RECT 37.246 2.196 37.332 2.347 ;
      RECT 37.16 2.182 37.246 2.337 ;
      RECT 37.115 2.172 37.16 2.33 ;
      RECT 37.095 1.46 37.115 1.738 ;
      RECT 37.095 2.165 37.115 2.326 ;
      RECT 37.065 1.46 37.095 1.76 ;
      RECT 37.055 2.132 37.095 2.323 ;
      RECT 37.05 1.46 37.065 1.78 ;
      RECT 37.05 2.097 37.055 2.321 ;
      RECT 37.045 1.46 37.05 1.905 ;
      RECT 37.045 2.057 37.05 2.321 ;
      RECT 37.035 1.46 37.045 2.321 ;
      RECT 36.96 1.46 37.035 2.315 ;
      RECT 36.93 1.46 36.96 2.305 ;
      RECT 36.925 1.46 36.93 2.297 ;
      RECT 36.92 1.502 36.925 2.29 ;
      RECT 36.91 1.571 36.92 2.281 ;
      RECT 36.905 1.641 36.91 2.233 ;
      RECT 36.9 1.705 36.905 2.13 ;
      RECT 36.895 1.74 36.9 2.085 ;
      RECT 36.893 1.777 36.895 1.977 ;
      RECT 36.89 1.785 36.893 1.97 ;
      RECT 36.885 1.85 36.89 1.913 ;
      RECT 40.96 0.94 41.24 1.22 ;
      RECT 40.95 0.94 41.24 1.083 ;
      RECT 40.905 0.805 41.165 1.065 ;
      RECT 40.905 0.92 41.22 1.065 ;
      RECT 40.905 0.89 41.215 1.065 ;
      RECT 40.905 0.877 41.205 1.065 ;
      RECT 40.905 0.867 41.2 1.065 ;
      RECT 36.88 0.85 37.14 1.11 ;
      RECT 40.65 0.4 40.91 0.66 ;
      RECT 40.64 0.425 40.91 0.62 ;
      RECT 40.635 0.425 40.64 0.619 ;
      RECT 40.565 0.42 40.635 0.611 ;
      RECT 40.48 0.407 40.565 0.594 ;
      RECT 40.476 0.399 40.48 0.584 ;
      RECT 40.39 0.392 40.476 0.574 ;
      RECT 40.381 0.384 40.39 0.564 ;
      RECT 40.295 0.377 40.381 0.552 ;
      RECT 40.275 0.368 40.295 0.538 ;
      RECT 40.22 0.363 40.275 0.53 ;
      RECT 40.21 0.357 40.22 0.524 ;
      RECT 40.19 0.355 40.21 0.52 ;
      RECT 40.182 0.354 40.19 0.516 ;
      RECT 40.096 0.346 40.182 0.505 ;
      RECT 40.01 0.332 40.096 0.485 ;
      RECT 39.95 0.32 40.01 0.47 ;
      RECT 39.94 0.315 39.95 0.465 ;
      RECT 39.89 0.315 39.94 0.467 ;
      RECT 39.843 0.317 39.89 0.471 ;
      RECT 39.757 0.324 39.843 0.476 ;
      RECT 39.671 0.332 39.757 0.482 ;
      RECT 39.585 0.341 39.671 0.488 ;
      RECT 39.526 0.347 39.585 0.493 ;
      RECT 39.44 0.352 39.526 0.499 ;
      RECT 39.365 0.357 39.44 0.505 ;
      RECT 39.326 0.359 39.365 0.51 ;
      RECT 39.24 0.356 39.326 0.515 ;
      RECT 39.155 0.354 39.24 0.522 ;
      RECT 39.123 0.353 39.155 0.525 ;
      RECT 39.037 0.352 39.123 0.526 ;
      RECT 38.951 0.351 39.037 0.527 ;
      RECT 38.865 0.35 38.951 0.527 ;
      RECT 38.779 0.349 38.865 0.528 ;
      RECT 38.693 0.348 38.779 0.529 ;
      RECT 38.607 0.347 38.693 0.53 ;
      RECT 38.521 0.346 38.607 0.53 ;
      RECT 38.435 0.345 38.521 0.531 ;
      RECT 38.385 0.345 38.435 0.532 ;
      RECT 38.371 0.346 38.385 0.532 ;
      RECT 38.285 0.353 38.371 0.533 ;
      RECT 38.211 0.364 38.285 0.534 ;
      RECT 38.125 0.373 38.211 0.535 ;
      RECT 38.09 0.38 38.125 0.55 ;
      RECT 38.065 0.383 38.09 0.58 ;
      RECT 38.04 0.392 38.065 0.609 ;
      RECT 38.03 0.403 38.04 0.629 ;
      RECT 38.02 0.411 38.03 0.643 ;
      RECT 38.015 0.417 38.02 0.653 ;
      RECT 37.99 0.434 38.015 0.67 ;
      RECT 37.975 0.456 37.99 0.698 ;
      RECT 37.945 0.482 37.975 0.728 ;
      RECT 37.925 0.511 37.945 0.758 ;
      RECT 37.92 0.526 37.925 0.775 ;
      RECT 37.9 0.541 37.92 0.79 ;
      RECT 37.89 0.559 37.9 0.808 ;
      RECT 37.88 0.57 37.89 0.823 ;
      RECT 37.83 0.602 37.88 0.849 ;
      RECT 37.825 0.632 37.83 0.869 ;
      RECT 37.815 0.645 37.825 0.875 ;
      RECT 37.806 0.655 37.815 0.883 ;
      RECT 37.795 0.666 37.806 0.891 ;
      RECT 37.79 0.676 37.795 0.897 ;
      RECT 37.775 0.697 37.79 0.904 ;
      RECT 37.76 0.727 37.775 0.912 ;
      RECT 37.725 0.757 37.76 0.918 ;
      RECT 37.7 0.775 37.725 0.925 ;
      RECT 37.65 0.783 37.7 0.934 ;
      RECT 37.625 0.788 37.65 0.943 ;
      RECT 37.57 0.794 37.625 0.953 ;
      RECT 37.565 0.799 37.57 0.961 ;
      RECT 37.551 0.802 37.565 0.963 ;
      RECT 37.465 0.814 37.551 0.975 ;
      RECT 37.455 0.826 37.465 0.988 ;
      RECT 37.37 0.839 37.455 1 ;
      RECT 37.326 0.856 37.37 1.014 ;
      RECT 37.24 0.873 37.326 1.03 ;
      RECT 37.21 0.887 37.24 1.044 ;
      RECT 37.2 0.892 37.21 1.049 ;
      RECT 37.14 0.895 37.2 1.058 ;
      RECT 40.03 1.165 40.29 1.425 ;
      RECT 40.03 1.165 40.31 1.278 ;
      RECT 40.03 1.165 40.335 1.245 ;
      RECT 40.03 1.165 40.34 1.225 ;
      RECT 40.08 0.94 40.36 1.22 ;
      RECT 39.635 1.675 39.895 1.935 ;
      RECT 39.625 1.532 39.82 1.873 ;
      RECT 39.62 1.64 39.835 1.865 ;
      RECT 39.615 1.69 39.895 1.855 ;
      RECT 39.605 1.767 39.895 1.84 ;
      RECT 39.625 1.615 39.835 1.873 ;
      RECT 39.635 1.49 39.82 1.935 ;
      RECT 39.635 1.385 39.8 1.935 ;
      RECT 39.645 1.372 39.8 1.935 ;
      RECT 39.645 1.33 39.79 1.935 ;
      RECT 39.65 1.255 39.79 1.935 ;
      RECT 39.68 0.905 39.79 1.935 ;
      RECT 39.685 0.635 39.81 1.258 ;
      RECT 39.655 1.21 39.81 1.258 ;
      RECT 39.67 1.012 39.79 1.935 ;
      RECT 39.66 1.122 39.81 1.258 ;
      RECT 39.685 0.635 39.825 1.115 ;
      RECT 39.685 0.635 39.845 0.99 ;
      RECT 39.65 0.635 39.91 0.895 ;
      RECT 39.12 0.94 39.4 1.22 ;
      RECT 39.105 0.94 39.4 1.2 ;
      RECT 37.16 1.805 37.42 2.065 ;
      RECT 38.945 1.66 39.205 1.92 ;
      RECT 38.925 1.68 39.205 1.895 ;
      RECT 38.882 1.68 38.925 1.894 ;
      RECT 38.796 1.681 38.882 1.891 ;
      RECT 38.71 1.682 38.796 1.887 ;
      RECT 38.635 1.684 38.71 1.884 ;
      RECT 38.612 1.685 38.635 1.882 ;
      RECT 38.526 1.686 38.612 1.88 ;
      RECT 38.44 1.687 38.526 1.877 ;
      RECT 38.416 1.688 38.44 1.875 ;
      RECT 38.33 1.69 38.416 1.872 ;
      RECT 38.245 1.692 38.33 1.873 ;
      RECT 38.188 1.693 38.245 1.879 ;
      RECT 38.102 1.695 38.188 1.889 ;
      RECT 38.016 1.698 38.102 1.902 ;
      RECT 37.93 1.7 38.016 1.914 ;
      RECT 37.916 1.701 37.93 1.921 ;
      RECT 37.83 1.702 37.916 1.929 ;
      RECT 37.79 1.704 37.83 1.938 ;
      RECT 37.781 1.705 37.79 1.941 ;
      RECT 37.695 1.713 37.781 1.947 ;
      RECT 37.675 1.722 37.695 1.955 ;
      RECT 37.59 1.737 37.675 1.963 ;
      RECT 37.53 1.76 37.59 1.974 ;
      RECT 37.52 1.772 37.53 1.979 ;
      RECT 37.48 1.782 37.52 1.983 ;
      RECT 37.425 1.799 37.48 1.991 ;
      RECT 37.42 1.809 37.425 1.995 ;
      RECT 38.486 0.94 38.545 1.337 ;
      RECT 38.4 0.94 38.605 1.328 ;
      RECT 38.395 0.97 38.605 1.323 ;
      RECT 38.361 0.97 38.605 1.321 ;
      RECT 38.275 0.97 38.605 1.315 ;
      RECT 38.23 0.97 38.625 1.293 ;
      RECT 38.23 0.97 38.645 1.248 ;
      RECT 38.19 0.97 38.645 1.238 ;
      RECT 38.4 0.94 38.68 1.22 ;
      RECT 38.135 0.94 38.395 1.2 ;
      RECT 37.32 0.42 37.58 0.68 ;
      RECT 37.4 0.38 37.68 0.66 ;
      RECT 35.96 1.5 36.24 1.78 ;
      RECT 35.93 1.462 36.185 1.765 ;
      RECT 35.925 1.463 36.185 1.763 ;
      RECT 35.92 1.464 36.185 1.757 ;
      RECT 35.915 1.467 36.185 1.75 ;
      RECT 35.91 1.5 36.24 1.743 ;
      RECT 35.88 1.47 36.185 1.73 ;
      RECT 35.88 1.497 36.205 1.73 ;
      RECT 35.88 1.487 36.2 1.73 ;
      RECT 35.88 1.472 36.195 1.73 ;
      RECT 35.96 1.459 36.175 1.78 ;
      RECT 36.046 1.457 36.175 1.78 ;
      RECT 36.132 1.455 36.16 1.78 ;
      RECT 23.29 0.35 23.66 0.72 ;
      RECT 23.805 0.365 24.065 0.69 ;
      RECT 23.29 0.395 24.065 0.655 ;
      RECT 14.075 0.955 14.31 1.215 ;
      RECT 17.22 0.735 17.385 0.995 ;
      RECT 17.125 0.725 17.14 0.995 ;
      RECT 15.725 0.295 15.765 0.435 ;
      RECT 17.14 0.73 17.22 0.995 ;
      RECT 17.085 0.725 17.125 0.961 ;
      RECT 17.071 0.725 17.085 0.961 ;
      RECT 16.985 0.73 17.071 0.963 ;
      RECT 16.94 0.737 16.985 0.965 ;
      RECT 16.91 0.737 16.94 0.967 ;
      RECT 16.885 0.732 16.91 0.969 ;
      RECT 16.855 0.728 16.885 0.978 ;
      RECT 16.845 0.725 16.855 0.99 ;
      RECT 16.84 0.725 16.845 0.998 ;
      RECT 16.835 0.725 16.84 1.003 ;
      RECT 16.825 0.724 16.835 1.013 ;
      RECT 16.82 0.723 16.825 1.023 ;
      RECT 16.805 0.722 16.82 1.028 ;
      RECT 16.777 0.719 16.805 1.055 ;
      RECT 16.691 0.711 16.777 1.055 ;
      RECT 16.605 0.7 16.691 1.055 ;
      RECT 16.565 0.685 16.605 1.055 ;
      RECT 16.525 0.659 16.565 1.055 ;
      RECT 16.52 0.641 16.525 0.867 ;
      RECT 16.51 0.637 16.52 0.857 ;
      RECT 16.495 0.627 16.51 0.844 ;
      RECT 16.475 0.611 16.495 0.829 ;
      RECT 16.46 0.596 16.475 0.814 ;
      RECT 16.45 0.585 16.46 0.804 ;
      RECT 16.425 0.569 16.45 0.793 ;
      RECT 16.42 0.556 16.425 0.783 ;
      RECT 16.415 0.552 16.42 0.778 ;
      RECT 16.36 0.538 16.415 0.756 ;
      RECT 16.321 0.519 16.36 0.72 ;
      RECT 16.235 0.493 16.321 0.673 ;
      RECT 16.231 0.475 16.235 0.639 ;
      RECT 16.145 0.456 16.231 0.617 ;
      RECT 16.14 0.438 16.145 0.595 ;
      RECT 16.135 0.436 16.14 0.593 ;
      RECT 16.125 0.435 16.135 0.588 ;
      RECT 16.065 0.422 16.125 0.574 ;
      RECT 16.02 0.4 16.065 0.553 ;
      RECT 15.96 0.377 16.02 0.532 ;
      RECT 15.896 0.352 15.96 0.507 ;
      RECT 15.81 0.322 15.896 0.476 ;
      RECT 15.795 0.302 15.81 0.455 ;
      RECT 15.765 0.297 15.795 0.446 ;
      RECT 15.712 0.295 15.725 0.435 ;
      RECT 15.626 0.295 15.712 0.437 ;
      RECT 15.54 0.295 15.626 0.439 ;
      RECT 15.52 0.295 15.54 0.443 ;
      RECT 15.475 0.297 15.52 0.454 ;
      RECT 15.435 0.307 15.475 0.47 ;
      RECT 15.431 0.316 15.435 0.478 ;
      RECT 15.345 0.336 15.431 0.494 ;
      RECT 15.335 0.355 15.345 0.512 ;
      RECT 15.33 0.357 15.335 0.515 ;
      RECT 15.32 0.361 15.33 0.518 ;
      RECT 15.3 0.366 15.32 0.528 ;
      RECT 15.27 0.376 15.3 0.548 ;
      RECT 15.265 0.383 15.27 0.562 ;
      RECT 15.255 0.387 15.265 0.569 ;
      RECT 15.24 0.395 15.255 0.58 ;
      RECT 15.23 0.405 15.24 0.591 ;
      RECT 15.22 0.412 15.23 0.599 ;
      RECT 15.195 0.425 15.22 0.614 ;
      RECT 15.131 0.461 15.195 0.653 ;
      RECT 15.045 0.524 15.131 0.717 ;
      RECT 15.01 0.575 15.045 0.77 ;
      RECT 15.005 0.592 15.01 0.787 ;
      RECT 14.99 0.601 15.005 0.794 ;
      RECT 14.97 0.616 14.99 0.808 ;
      RECT 14.965 0.627 14.97 0.818 ;
      RECT 14.945 0.64 14.965 0.828 ;
      RECT 14.94 0.65 14.945 0.838 ;
      RECT 14.925 0.655 14.94 0.847 ;
      RECT 14.915 0.665 14.925 0.858 ;
      RECT 14.885 0.682 14.915 0.875 ;
      RECT 14.875 0.7 14.885 0.893 ;
      RECT 14.86 0.711 14.875 0.904 ;
      RECT 14.82 0.735 14.86 0.92 ;
      RECT 14.785 0.769 14.82 0.937 ;
      RECT 14.755 0.792 14.785 0.949 ;
      RECT 14.74 0.802 14.755 0.958 ;
      RECT 14.7 0.812 14.74 0.969 ;
      RECT 14.68 0.823 14.7 0.981 ;
      RECT 14.675 0.827 14.68 0.988 ;
      RECT 14.66 0.831 14.675 0.993 ;
      RECT 14.65 0.836 14.66 0.998 ;
      RECT 14.645 0.839 14.65 1.001 ;
      RECT 14.615 0.845 14.645 1.008 ;
      RECT 14.58 0.855 14.615 1.022 ;
      RECT 14.52 0.87 14.58 1.042 ;
      RECT 14.465 0.89 14.52 1.066 ;
      RECT 14.436 0.905 14.465 1.084 ;
      RECT 14.35 0.925 14.436 1.109 ;
      RECT 14.345 0.94 14.35 1.129 ;
      RECT 14.335 0.943 14.345 1.13 ;
      RECT 14.31 0.95 14.335 1.215 ;
      RECT 17.005 1.443 17.285 1.78 ;
      RECT 17.005 1.453 17.29 1.738 ;
      RECT 17.005 1.462 17.295 1.635 ;
      RECT 17.005 1.477 17.3 1.503 ;
      RECT 17.005 1.305 17.265 1.78 ;
      RECT 14.725 2.185 14.735 2.375 ;
      RECT 12.985 2.06 13.265 2.34 ;
      RECT 16.03 1 16.035 1.485 ;
      RECT 15.925 1 15.985 1.26 ;
      RECT 16.25 1.97 16.255 2.045 ;
      RECT 16.24 1.837 16.25 2.08 ;
      RECT 16.23 1.672 16.24 2.101 ;
      RECT 16.225 1.542 16.23 2.117 ;
      RECT 16.215 1.432 16.225 2.133 ;
      RECT 16.21 1.331 16.215 2.15 ;
      RECT 16.205 1.313 16.21 2.16 ;
      RECT 16.2 1.295 16.205 2.17 ;
      RECT 16.19 1.27 16.2 2.185 ;
      RECT 16.185 1.25 16.19 2.2 ;
      RECT 16.165 1 16.185 2.225 ;
      RECT 16.15 1 16.165 2.258 ;
      RECT 16.12 1 16.15 2.28 ;
      RECT 16.1 1 16.12 2.294 ;
      RECT 16.08 1 16.1 1.81 ;
      RECT 16.095 1.877 16.1 2.299 ;
      RECT 16.09 1.907 16.095 2.301 ;
      RECT 16.085 1.92 16.09 2.304 ;
      RECT 16.08 1.93 16.085 2.308 ;
      RECT 16.075 1 16.08 1.728 ;
      RECT 16.075 1.94 16.08 2.31 ;
      RECT 16.07 1 16.075 1.705 ;
      RECT 16.06 1.962 16.075 2.31 ;
      RECT 16.055 1 16.07 1.65 ;
      RECT 16.05 1.987 16.06 2.31 ;
      RECT 16.05 1 16.055 1.595 ;
      RECT 16.04 1 16.05 1.543 ;
      RECT 16.045 2 16.05 2.311 ;
      RECT 16.04 2.012 16.045 2.312 ;
      RECT 16.035 1 16.04 1.503 ;
      RECT 16.035 2.025 16.04 2.313 ;
      RECT 16.02 2.04 16.035 2.314 ;
      RECT 16.025 1 16.03 1.465 ;
      RECT 16.02 1 16.025 1.43 ;
      RECT 16.015 1 16.02 1.405 ;
      RECT 16.01 2.067 16.02 2.316 ;
      RECT 16.005 1 16.015 1.363 ;
      RECT 16.005 2.085 16.01 2.317 ;
      RECT 16 1 16.005 1.323 ;
      RECT 16 2.092 16.005 2.318 ;
      RECT 15.995 1 16 1.295 ;
      RECT 15.99 2.11 16 2.319 ;
      RECT 15.985 1 15.995 1.275 ;
      RECT 15.98 2.13 15.99 2.321 ;
      RECT 15.97 2.147 15.98 2.322 ;
      RECT 15.935 2.17 15.97 2.325 ;
      RECT 15.88 2.188 15.935 2.331 ;
      RECT 15.794 2.196 15.88 2.34 ;
      RECT 15.708 2.207 15.794 2.351 ;
      RECT 15.622 2.217 15.708 2.362 ;
      RECT 15.536 2.227 15.622 2.374 ;
      RECT 15.45 2.237 15.536 2.385 ;
      RECT 15.43 2.243 15.45 2.391 ;
      RECT 15.35 2.245 15.43 2.395 ;
      RECT 15.345 2.244 15.35 2.4 ;
      RECT 15.337 2.243 15.345 2.4 ;
      RECT 15.251 2.239 15.337 2.398 ;
      RECT 15.165 2.231 15.251 2.395 ;
      RECT 15.079 2.222 15.165 2.391 ;
      RECT 14.993 2.214 15.079 2.388 ;
      RECT 14.907 2.206 14.993 2.384 ;
      RECT 14.821 2.197 14.907 2.381 ;
      RECT 14.735 2.189 14.821 2.377 ;
      RECT 14.68 2.182 14.725 2.375 ;
      RECT 14.595 2.175 14.68 2.373 ;
      RECT 14.521 2.167 14.595 2.369 ;
      RECT 14.435 2.159 14.521 2.366 ;
      RECT 14.432 2.155 14.435 2.364 ;
      RECT 14.346 2.151 14.432 2.363 ;
      RECT 14.26 2.143 14.346 2.36 ;
      RECT 14.175 2.138 14.26 2.357 ;
      RECT 14.089 2.135 14.175 2.354 ;
      RECT 14.003 2.133 14.089 2.351 ;
      RECT 13.917 2.13 14.003 2.348 ;
      RECT 13.831 2.127 13.917 2.345 ;
      RECT 13.745 2.124 13.831 2.342 ;
      RECT 13.669 2.122 13.745 2.339 ;
      RECT 13.583 2.119 13.669 2.336 ;
      RECT 13.497 2.116 13.583 2.334 ;
      RECT 13.411 2.114 13.497 2.331 ;
      RECT 13.325 2.111 13.411 2.328 ;
      RECT 13.265 2.102 13.325 2.326 ;
      RECT 15.775 1.72 15.85 1.98 ;
      RECT 15.755 1.7 15.76 1.98 ;
      RECT 15.075 1.485 15.18 1.78 ;
      RECT 9.52 1.46 9.59 1.72 ;
      RECT 15.415 1.335 15.42 1.706 ;
      RECT 15.405 1.39 15.41 1.706 ;
      RECT 15.71 0.56 15.77 0.82 ;
      RECT 15.765 1.715 15.775 1.98 ;
      RECT 15.76 1.705 15.765 1.98 ;
      RECT 15.68 1.652 15.755 1.98 ;
      RECT 15.705 0.56 15.71 0.84 ;
      RECT 15.695 0.56 15.705 0.86 ;
      RECT 15.68 0.56 15.695 0.89 ;
      RECT 15.665 0.56 15.68 0.933 ;
      RECT 15.66 1.595 15.68 1.98 ;
      RECT 15.65 0.56 15.665 0.97 ;
      RECT 15.645 1.575 15.66 1.98 ;
      RECT 15.645 0.56 15.65 0.993 ;
      RECT 15.635 0.56 15.645 1.018 ;
      RECT 15.605 1.542 15.645 1.98 ;
      RECT 15.61 0.56 15.635 1.068 ;
      RECT 15.605 0.56 15.61 1.123 ;
      RECT 15.6 0.56 15.605 1.165 ;
      RECT 15.59 1.505 15.605 1.98 ;
      RECT 15.595 0.56 15.6 1.208 ;
      RECT 15.59 0.56 15.595 1.273 ;
      RECT 15.585 0.56 15.59 1.295 ;
      RECT 15.585 1.493 15.59 1.845 ;
      RECT 15.58 0.56 15.585 1.363 ;
      RECT 15.58 1.485 15.585 1.828 ;
      RECT 15.575 0.56 15.58 1.408 ;
      RECT 15.57 1.467 15.58 1.805 ;
      RECT 15.57 0.56 15.575 1.445 ;
      RECT 15.56 0.56 15.57 1.785 ;
      RECT 15.555 0.56 15.56 1.768 ;
      RECT 15.55 0.56 15.555 1.753 ;
      RECT 15.545 0.56 15.55 1.738 ;
      RECT 15.525 0.56 15.545 1.728 ;
      RECT 15.52 0.56 15.525 1.718 ;
      RECT 15.51 0.56 15.52 1.714 ;
      RECT 15.505 0.837 15.51 1.713 ;
      RECT 15.5 0.86 15.505 1.712 ;
      RECT 15.495 0.89 15.5 1.711 ;
      RECT 15.49 0.917 15.495 1.71 ;
      RECT 15.485 0.945 15.49 1.71 ;
      RECT 15.48 0.972 15.485 1.71 ;
      RECT 15.475 0.992 15.48 1.71 ;
      RECT 15.47 1.02 15.475 1.71 ;
      RECT 15.46 1.062 15.47 1.71 ;
      RECT 15.45 1.107 15.46 1.709 ;
      RECT 15.445 1.16 15.45 1.708 ;
      RECT 15.44 1.192 15.445 1.707 ;
      RECT 15.435 1.212 15.44 1.706 ;
      RECT 15.43 1.25 15.435 1.706 ;
      RECT 15.425 1.272 15.43 1.706 ;
      RECT 15.42 1.297 15.425 1.706 ;
      RECT 15.41 1.362 15.415 1.706 ;
      RECT 15.395 1.422 15.405 1.706 ;
      RECT 15.38 1.432 15.395 1.706 ;
      RECT 15.36 1.442 15.38 1.706 ;
      RECT 15.33 1.447 15.36 1.703 ;
      RECT 15.27 1.457 15.33 1.7 ;
      RECT 15.25 1.466 15.27 1.705 ;
      RECT 15.225 1.472 15.25 1.718 ;
      RECT 15.205 1.477 15.225 1.733 ;
      RECT 15.18 1.482 15.205 1.78 ;
      RECT 15.051 1.484 15.075 1.78 ;
      RECT 14.965 1.479 15.051 1.78 ;
      RECT 14.925 1.476 14.965 1.78 ;
      RECT 14.875 1.478 14.925 1.76 ;
      RECT 14.845 1.482 14.875 1.76 ;
      RECT 14.766 1.492 14.845 1.76 ;
      RECT 14.68 1.507 14.766 1.761 ;
      RECT 14.63 1.517 14.68 1.762 ;
      RECT 14.622 1.52 14.63 1.762 ;
      RECT 14.536 1.522 14.622 1.763 ;
      RECT 14.45 1.526 14.536 1.763 ;
      RECT 14.364 1.53 14.45 1.764 ;
      RECT 14.278 1.533 14.364 1.765 ;
      RECT 14.192 1.537 14.278 1.765 ;
      RECT 14.106 1.541 14.192 1.766 ;
      RECT 14.02 1.544 14.106 1.767 ;
      RECT 13.934 1.548 14.02 1.767 ;
      RECT 13.848 1.552 13.934 1.768 ;
      RECT 13.762 1.556 13.848 1.769 ;
      RECT 13.676 1.559 13.762 1.769 ;
      RECT 13.59 1.563 13.676 1.77 ;
      RECT 13.56 1.565 13.59 1.77 ;
      RECT 13.474 1.568 13.56 1.771 ;
      RECT 13.388 1.572 13.474 1.772 ;
      RECT 13.302 1.576 13.388 1.773 ;
      RECT 13.216 1.579 13.302 1.773 ;
      RECT 13.13 1.583 13.216 1.774 ;
      RECT 13.095 1.588 13.13 1.775 ;
      RECT 13.04 1.598 13.095 1.782 ;
      RECT 13.015 1.61 13.04 1.792 ;
      RECT 12.98 1.623 13.015 1.8 ;
      RECT 12.94 1.64 12.98 1.823 ;
      RECT 12.92 1.653 12.94 1.85 ;
      RECT 12.89 1.665 12.92 1.878 ;
      RECT 12.885 1.673 12.89 1.898 ;
      RECT 12.88 1.676 12.885 1.908 ;
      RECT 12.83 1.688 12.88 1.942 ;
      RECT 12.82 1.703 12.83 1.975 ;
      RECT 12.81 1.709 12.82 1.988 ;
      RECT 12.8 1.716 12.81 2 ;
      RECT 12.775 1.729 12.8 2.018 ;
      RECT 12.76 1.744 12.775 2.04 ;
      RECT 12.75 1.752 12.76 2.056 ;
      RECT 12.735 1.761 12.75 2.071 ;
      RECT 12.725 1.771 12.735 2.085 ;
      RECT 12.706 1.784 12.725 2.102 ;
      RECT 12.62 1.829 12.706 2.167 ;
      RECT 12.605 1.874 12.62 2.225 ;
      RECT 12.6 1.883 12.605 2.238 ;
      RECT 12.59 1.89 12.6 2.243 ;
      RECT 12.585 1.895 12.59 2.247 ;
      RECT 12.565 1.905 12.585 2.254 ;
      RECT 12.54 1.925 12.565 2.268 ;
      RECT 12.505 1.95 12.54 2.288 ;
      RECT 12.49 1.973 12.505 2.303 ;
      RECT 12.48 1.983 12.49 2.308 ;
      RECT 12.47 1.991 12.48 2.315 ;
      RECT 12.46 2 12.47 2.321 ;
      RECT 12.44 2.012 12.46 2.323 ;
      RECT 12.43 2.025 12.44 2.325 ;
      RECT 12.405 2.04 12.43 2.328 ;
      RECT 12.385 2.057 12.405 2.332 ;
      RECT 12.345 2.085 12.385 2.338 ;
      RECT 12.28 2.132 12.345 2.347 ;
      RECT 12.265 2.165 12.28 2.355 ;
      RECT 12.26 2.172 12.265 2.357 ;
      RECT 12.21 2.197 12.26 2.362 ;
      RECT 12.195 2.221 12.21 2.369 ;
      RECT 12.145 2.226 12.195 2.37 ;
      RECT 12.059 2.23 12.145 2.37 ;
      RECT 11.973 2.23 12.059 2.37 ;
      RECT 11.887 2.23 11.973 2.371 ;
      RECT 11.801 2.23 11.887 2.371 ;
      RECT 11.715 2.23 11.801 2.371 ;
      RECT 11.649 2.23 11.715 2.371 ;
      RECT 11.563 2.23 11.649 2.372 ;
      RECT 11.477 2.23 11.563 2.372 ;
      RECT 11.391 2.231 11.477 2.373 ;
      RECT 11.305 2.231 11.391 2.373 ;
      RECT 11.219 2.231 11.305 2.373 ;
      RECT 11.133 2.231 11.219 2.374 ;
      RECT 11.047 2.231 11.133 2.374 ;
      RECT 10.961 2.232 11.047 2.375 ;
      RECT 10.875 2.232 10.961 2.375 ;
      RECT 10.855 2.232 10.875 2.375 ;
      RECT 10.769 2.232 10.855 2.375 ;
      RECT 10.683 2.232 10.769 2.375 ;
      RECT 10.597 2.233 10.683 2.375 ;
      RECT 10.511 2.233 10.597 2.375 ;
      RECT 10.425 2.233 10.511 2.375 ;
      RECT 10.339 2.234 10.425 2.375 ;
      RECT 10.253 2.234 10.339 2.375 ;
      RECT 10.167 2.234 10.253 2.375 ;
      RECT 10.081 2.234 10.167 2.375 ;
      RECT 9.995 2.235 10.081 2.375 ;
      RECT 9.945 2.232 9.995 2.375 ;
      RECT 9.935 2.23 9.945 2.374 ;
      RECT 9.931 2.23 9.935 2.373 ;
      RECT 9.845 2.225 9.931 2.368 ;
      RECT 9.823 2.218 9.845 2.362 ;
      RECT 9.737 2.209 9.823 2.356 ;
      RECT 9.651 2.196 9.737 2.347 ;
      RECT 9.565 2.182 9.651 2.337 ;
      RECT 9.52 2.172 9.565 2.33 ;
      RECT 9.5 1.46 9.52 1.738 ;
      RECT 9.5 2.165 9.52 2.326 ;
      RECT 9.47 1.46 9.5 1.76 ;
      RECT 9.46 2.132 9.5 2.323 ;
      RECT 9.455 1.46 9.47 1.78 ;
      RECT 9.455 2.097 9.46 2.321 ;
      RECT 9.45 1.46 9.455 1.905 ;
      RECT 9.45 2.057 9.455 2.321 ;
      RECT 9.44 1.46 9.45 2.321 ;
      RECT 9.365 1.46 9.44 2.315 ;
      RECT 9.335 1.46 9.365 2.305 ;
      RECT 9.33 1.46 9.335 2.297 ;
      RECT 9.325 1.502 9.33 2.29 ;
      RECT 9.315 1.571 9.325 2.281 ;
      RECT 9.31 1.641 9.315 2.233 ;
      RECT 9.305 1.705 9.31 2.13 ;
      RECT 9.3 1.74 9.305 2.085 ;
      RECT 9.298 1.777 9.3 1.977 ;
      RECT 9.295 1.785 9.298 1.97 ;
      RECT 9.29 1.85 9.295 1.913 ;
      RECT 13.365 0.94 13.645 1.22 ;
      RECT 13.355 0.94 13.645 1.083 ;
      RECT 13.31 0.805 13.57 1.065 ;
      RECT 13.31 0.92 13.625 1.065 ;
      RECT 13.31 0.89 13.62 1.065 ;
      RECT 13.31 0.877 13.61 1.065 ;
      RECT 13.31 0.867 13.605 1.065 ;
      RECT 9.285 0.85 9.545 1.11 ;
      RECT 13.055 0.4 13.315 0.66 ;
      RECT 13.045 0.425 13.315 0.62 ;
      RECT 13.04 0.425 13.045 0.619 ;
      RECT 12.97 0.42 13.04 0.611 ;
      RECT 12.885 0.407 12.97 0.594 ;
      RECT 12.881 0.399 12.885 0.584 ;
      RECT 12.795 0.392 12.881 0.574 ;
      RECT 12.786 0.384 12.795 0.564 ;
      RECT 12.7 0.377 12.786 0.552 ;
      RECT 12.68 0.368 12.7 0.538 ;
      RECT 12.625 0.363 12.68 0.53 ;
      RECT 12.615 0.357 12.625 0.524 ;
      RECT 12.595 0.355 12.615 0.52 ;
      RECT 12.587 0.354 12.595 0.516 ;
      RECT 12.501 0.346 12.587 0.505 ;
      RECT 12.415 0.332 12.501 0.485 ;
      RECT 12.355 0.32 12.415 0.47 ;
      RECT 12.345 0.315 12.355 0.465 ;
      RECT 12.295 0.315 12.345 0.467 ;
      RECT 12.248 0.317 12.295 0.471 ;
      RECT 12.162 0.324 12.248 0.476 ;
      RECT 12.076 0.332 12.162 0.482 ;
      RECT 11.99 0.341 12.076 0.488 ;
      RECT 11.931 0.347 11.99 0.493 ;
      RECT 11.845 0.352 11.931 0.499 ;
      RECT 11.77 0.357 11.845 0.505 ;
      RECT 11.731 0.359 11.77 0.51 ;
      RECT 11.645 0.356 11.731 0.515 ;
      RECT 11.56 0.354 11.645 0.522 ;
      RECT 11.528 0.353 11.56 0.525 ;
      RECT 11.442 0.352 11.528 0.526 ;
      RECT 11.356 0.351 11.442 0.527 ;
      RECT 11.27 0.35 11.356 0.527 ;
      RECT 11.184 0.349 11.27 0.528 ;
      RECT 11.098 0.348 11.184 0.529 ;
      RECT 11.012 0.347 11.098 0.53 ;
      RECT 10.926 0.346 11.012 0.53 ;
      RECT 10.84 0.345 10.926 0.531 ;
      RECT 10.79 0.345 10.84 0.532 ;
      RECT 10.776 0.346 10.79 0.532 ;
      RECT 10.69 0.353 10.776 0.533 ;
      RECT 10.616 0.364 10.69 0.534 ;
      RECT 10.53 0.373 10.616 0.535 ;
      RECT 10.495 0.38 10.53 0.55 ;
      RECT 10.47 0.383 10.495 0.58 ;
      RECT 10.445 0.392 10.47 0.609 ;
      RECT 10.435 0.403 10.445 0.629 ;
      RECT 10.425 0.411 10.435 0.643 ;
      RECT 10.42 0.417 10.425 0.653 ;
      RECT 10.395 0.434 10.42 0.67 ;
      RECT 10.38 0.456 10.395 0.698 ;
      RECT 10.35 0.482 10.38 0.728 ;
      RECT 10.33 0.511 10.35 0.758 ;
      RECT 10.325 0.526 10.33 0.775 ;
      RECT 10.305 0.541 10.325 0.79 ;
      RECT 10.295 0.559 10.305 0.808 ;
      RECT 10.285 0.57 10.295 0.823 ;
      RECT 10.235 0.602 10.285 0.849 ;
      RECT 10.23 0.632 10.235 0.869 ;
      RECT 10.22 0.645 10.23 0.875 ;
      RECT 10.211 0.655 10.22 0.883 ;
      RECT 10.2 0.666 10.211 0.891 ;
      RECT 10.195 0.676 10.2 0.897 ;
      RECT 10.18 0.697 10.195 0.904 ;
      RECT 10.165 0.727 10.18 0.912 ;
      RECT 10.13 0.757 10.165 0.918 ;
      RECT 10.105 0.775 10.13 0.925 ;
      RECT 10.055 0.783 10.105 0.934 ;
      RECT 10.03 0.788 10.055 0.943 ;
      RECT 9.975 0.794 10.03 0.953 ;
      RECT 9.97 0.799 9.975 0.961 ;
      RECT 9.956 0.802 9.97 0.963 ;
      RECT 9.87 0.814 9.956 0.975 ;
      RECT 9.86 0.826 9.87 0.988 ;
      RECT 9.775 0.839 9.86 1 ;
      RECT 9.731 0.856 9.775 1.014 ;
      RECT 9.645 0.873 9.731 1.03 ;
      RECT 9.615 0.887 9.645 1.044 ;
      RECT 9.605 0.892 9.615 1.049 ;
      RECT 9.545 0.895 9.605 1.058 ;
      RECT 12.435 1.165 12.695 1.425 ;
      RECT 12.435 1.165 12.715 1.278 ;
      RECT 12.435 1.165 12.74 1.245 ;
      RECT 12.435 1.165 12.745 1.225 ;
      RECT 12.485 0.94 12.765 1.22 ;
      RECT 12.04 1.675 12.3 1.935 ;
      RECT 12.03 1.532 12.225 1.873 ;
      RECT 12.025 1.64 12.24 1.865 ;
      RECT 12.02 1.69 12.3 1.855 ;
      RECT 12.01 1.767 12.3 1.84 ;
      RECT 12.03 1.615 12.24 1.873 ;
      RECT 12.04 1.49 12.225 1.935 ;
      RECT 12.04 1.385 12.205 1.935 ;
      RECT 12.05 1.372 12.205 1.935 ;
      RECT 12.05 1.33 12.195 1.935 ;
      RECT 12.055 1.255 12.195 1.935 ;
      RECT 12.085 0.905 12.195 1.935 ;
      RECT 12.09 0.635 12.215 1.258 ;
      RECT 12.06 1.21 12.215 1.258 ;
      RECT 12.075 1.012 12.195 1.935 ;
      RECT 12.065 1.122 12.215 1.258 ;
      RECT 12.09 0.635 12.23 1.115 ;
      RECT 12.09 0.635 12.25 0.99 ;
      RECT 12.055 0.635 12.315 0.895 ;
      RECT 11.525 0.94 11.805 1.22 ;
      RECT 11.51 0.94 11.805 1.2 ;
      RECT 9.565 1.805 9.825 2.065 ;
      RECT 11.35 1.66 11.61 1.92 ;
      RECT 11.33 1.68 11.61 1.895 ;
      RECT 11.287 1.68 11.33 1.894 ;
      RECT 11.201 1.681 11.287 1.891 ;
      RECT 11.115 1.682 11.201 1.887 ;
      RECT 11.04 1.684 11.115 1.884 ;
      RECT 11.017 1.685 11.04 1.882 ;
      RECT 10.931 1.686 11.017 1.88 ;
      RECT 10.845 1.687 10.931 1.877 ;
      RECT 10.821 1.688 10.845 1.875 ;
      RECT 10.735 1.69 10.821 1.872 ;
      RECT 10.65 1.692 10.735 1.873 ;
      RECT 10.593 1.693 10.65 1.879 ;
      RECT 10.507 1.695 10.593 1.889 ;
      RECT 10.421 1.698 10.507 1.902 ;
      RECT 10.335 1.7 10.421 1.914 ;
      RECT 10.321 1.701 10.335 1.921 ;
      RECT 10.235 1.702 10.321 1.929 ;
      RECT 10.195 1.704 10.235 1.938 ;
      RECT 10.186 1.705 10.195 1.941 ;
      RECT 10.1 1.713 10.186 1.947 ;
      RECT 10.08 1.722 10.1 1.955 ;
      RECT 9.995 1.737 10.08 1.963 ;
      RECT 9.935 1.76 9.995 1.974 ;
      RECT 9.925 1.772 9.935 1.979 ;
      RECT 9.885 1.782 9.925 1.983 ;
      RECT 9.83 1.799 9.885 1.991 ;
      RECT 9.825 1.809 9.83 1.995 ;
      RECT 10.891 0.94 10.95 1.337 ;
      RECT 10.805 0.94 11.01 1.328 ;
      RECT 10.8 0.97 11.01 1.323 ;
      RECT 10.766 0.97 11.01 1.321 ;
      RECT 10.68 0.97 11.01 1.315 ;
      RECT 10.635 0.97 11.03 1.293 ;
      RECT 10.635 0.97 11.05 1.248 ;
      RECT 10.595 0.97 11.05 1.238 ;
      RECT 10.805 0.94 11.085 1.22 ;
      RECT 10.54 0.94 10.8 1.2 ;
      RECT 9.725 0.42 9.985 0.68 ;
      RECT 9.805 0.38 10.085 0.66 ;
      RECT 8.365 1.5 8.645 1.78 ;
      RECT 8.335 1.462 8.59 1.765 ;
      RECT 8.33 1.463 8.59 1.763 ;
      RECT 8.325 1.464 8.59 1.757 ;
      RECT 8.32 1.467 8.59 1.75 ;
      RECT 8.315 1.5 8.645 1.743 ;
      RECT 8.285 1.47 8.59 1.73 ;
      RECT 8.285 1.497 8.61 1.73 ;
      RECT 8.285 1.487 8.605 1.73 ;
      RECT 8.285 1.472 8.6 1.73 ;
      RECT 8.365 1.459 8.58 1.78 ;
      RECT 8.451 1.457 8.58 1.78 ;
      RECT 8.537 1.455 8.565 1.78 ;
      RECT 138.685 0.8 139.055 1.175 ;
      RECT 135.465 1.37 135.815 1.74 ;
      RECT 134.655 0.5 134.935 0.87 ;
      RECT 131.33 1.37 131.68 1.74 ;
      RECT 130.115 0.44 130.395 0.81 ;
      RECT 129.655 1.16 130.025 1.53 ;
      RECT 127.97 -0.18 128.34 0.19 ;
      RECT 117.53 1.37 117.88 1.74 ;
      RECT 116.72 0.43 117 0.8 ;
      RECT 114.29 1.47 114.66 1.84 ;
      RECT 107.87 1.37 108.22 1.74 ;
      RECT 107.06 0.5 107.34 0.87 ;
      RECT 103.735 1.37 104.085 1.74 ;
      RECT 102.52 0.44 102.8 0.81 ;
      RECT 102.06 1.16 102.43 1.53 ;
      RECT 100.375 -0.18 100.745 0.19 ;
      RECT 89.935 1.37 90.285 1.74 ;
      RECT 89.125 0.43 89.405 0.8 ;
      RECT 86.695 1.47 87.065 1.84 ;
      RECT 80.275 1.37 80.625 1.74 ;
      RECT 79.465 0.5 79.745 0.87 ;
      RECT 76.14 1.37 76.49 1.74 ;
      RECT 74.925 0.44 75.205 0.81 ;
      RECT 74.465 1.16 74.835 1.53 ;
      RECT 72.78 -0.18 73.15 0.19 ;
      RECT 62.34 1.37 62.69 1.74 ;
      RECT 61.53 0.43 61.81 0.8 ;
      RECT 59.1 1.47 59.47 1.84 ;
      RECT 52.68 1.37 53.03 1.74 ;
      RECT 51.87 0.5 52.15 0.87 ;
      RECT 48.545 1.37 48.895 1.74 ;
      RECT 47.33 0.44 47.61 0.81 ;
      RECT 46.87 1.16 47.24 1.53 ;
      RECT 45.185 -0.18 45.555 0.19 ;
      RECT 34.745 1.37 35.095 1.74 ;
      RECT 33.935 0.43 34.215 0.8 ;
      RECT 31.505 1.47 31.875 1.84 ;
      RECT 25.085 1.37 25.435 1.74 ;
      RECT 24.275 0.5 24.555 0.87 ;
      RECT 20.95 1.37 21.3 1.74 ;
      RECT 19.735 0.44 20.015 0.81 ;
      RECT 19.275 1.16 19.645 1.53 ;
      RECT 17.59 -0.18 17.96 0.19 ;
      RECT 7.15 1.37 7.5 1.74 ;
      RECT 6.34 0.43 6.62 0.8 ;
      RECT 3.91 1.47 4.28 1.84 ;
      RECT 1.925 0.595 2.295 0.965 ;
    LAYER via1 ;
      RECT 138.785 0.9 138.935 1.05 ;
      RECT 135.565 1.47 135.715 1.62 ;
      RECT 134.71 0.6 134.86 0.75 ;
      RECT 134.24 0.45 134.39 0.6 ;
      RECT 131.43 1.47 131.58 1.62 ;
      RECT 130.17 0.54 130.32 0.69 ;
      RECT 129.755 1.26 129.905 1.41 ;
      RECT 128.08 -0.07 128.23 0.08 ;
      RECT 127.56 0.79 127.71 0.94 ;
      RECT 127.44 1.36 127.59 1.51 ;
      RECT 126.36 1.055 126.51 1.205 ;
      RECT 126.025 1.775 126.175 1.925 ;
      RECT 125.945 0.615 126.095 0.765 ;
      RECT 124.51 1.01 124.66 1.16 ;
      RECT 123.745 0.86 123.895 1.01 ;
      RECT 123.49 0.455 123.64 0.605 ;
      RECT 122.87 1.22 123.02 1.37 ;
      RECT 122.49 0.69 122.64 0.84 ;
      RECT 122.475 1.73 122.625 1.88 ;
      RECT 121.945 0.995 122.095 1.145 ;
      RECT 121.785 1.715 121.935 1.865 ;
      RECT 120.975 0.995 121.125 1.145 ;
      RECT 120.16 0.475 120.31 0.625 ;
      RECT 120 1.86 120.15 2.01 ;
      RECT 119.765 1.515 119.915 1.665 ;
      RECT 119.72 0.905 119.87 1.055 ;
      RECT 118.72 1.525 118.87 1.675 ;
      RECT 117.63 1.47 117.78 1.62 ;
      RECT 116.775 0.53 116.925 0.68 ;
      RECT 114.41 1.57 114.56 1.72 ;
      RECT 107.97 1.47 108.12 1.62 ;
      RECT 107.115 0.6 107.265 0.75 ;
      RECT 106.645 0.45 106.795 0.6 ;
      RECT 103.835 1.47 103.985 1.62 ;
      RECT 102.575 0.54 102.725 0.69 ;
      RECT 102.16 1.26 102.31 1.41 ;
      RECT 100.485 -0.07 100.635 0.08 ;
      RECT 99.965 0.79 100.115 0.94 ;
      RECT 99.845 1.36 99.995 1.51 ;
      RECT 98.765 1.055 98.915 1.205 ;
      RECT 98.43 1.775 98.58 1.925 ;
      RECT 98.35 0.615 98.5 0.765 ;
      RECT 96.915 1.01 97.065 1.16 ;
      RECT 96.15 0.86 96.3 1.01 ;
      RECT 95.895 0.455 96.045 0.605 ;
      RECT 95.275 1.22 95.425 1.37 ;
      RECT 94.895 0.69 95.045 0.84 ;
      RECT 94.88 1.73 95.03 1.88 ;
      RECT 94.35 0.995 94.5 1.145 ;
      RECT 94.19 1.715 94.34 1.865 ;
      RECT 93.38 0.995 93.53 1.145 ;
      RECT 92.565 0.475 92.715 0.625 ;
      RECT 92.405 1.86 92.555 2.01 ;
      RECT 92.17 1.515 92.32 1.665 ;
      RECT 92.125 0.905 92.275 1.055 ;
      RECT 91.125 1.525 91.275 1.675 ;
      RECT 90.035 1.47 90.185 1.62 ;
      RECT 89.18 0.53 89.33 0.68 ;
      RECT 86.815 1.57 86.965 1.72 ;
      RECT 80.375 1.47 80.525 1.62 ;
      RECT 79.52 0.6 79.67 0.75 ;
      RECT 79.05 0.45 79.2 0.6 ;
      RECT 76.24 1.47 76.39 1.62 ;
      RECT 74.98 0.54 75.13 0.69 ;
      RECT 74.565 1.26 74.715 1.41 ;
      RECT 72.89 -0.07 73.04 0.08 ;
      RECT 72.37 0.79 72.52 0.94 ;
      RECT 72.25 1.36 72.4 1.51 ;
      RECT 71.17 1.055 71.32 1.205 ;
      RECT 70.835 1.775 70.985 1.925 ;
      RECT 70.755 0.615 70.905 0.765 ;
      RECT 69.32 1.01 69.47 1.16 ;
      RECT 68.555 0.86 68.705 1.01 ;
      RECT 68.3 0.455 68.45 0.605 ;
      RECT 67.68 1.22 67.83 1.37 ;
      RECT 67.3 0.69 67.45 0.84 ;
      RECT 67.285 1.73 67.435 1.88 ;
      RECT 66.755 0.995 66.905 1.145 ;
      RECT 66.595 1.715 66.745 1.865 ;
      RECT 65.785 0.995 65.935 1.145 ;
      RECT 64.97 0.475 65.12 0.625 ;
      RECT 64.81 1.86 64.96 2.01 ;
      RECT 64.575 1.515 64.725 1.665 ;
      RECT 64.53 0.905 64.68 1.055 ;
      RECT 63.53 1.525 63.68 1.675 ;
      RECT 62.44 1.47 62.59 1.62 ;
      RECT 61.585 0.53 61.735 0.68 ;
      RECT 59.22 1.57 59.37 1.72 ;
      RECT 52.78 1.47 52.93 1.62 ;
      RECT 51.925 0.6 52.075 0.75 ;
      RECT 51.455 0.45 51.605 0.6 ;
      RECT 48.645 1.47 48.795 1.62 ;
      RECT 47.385 0.54 47.535 0.69 ;
      RECT 46.97 1.26 47.12 1.41 ;
      RECT 45.295 -0.07 45.445 0.08 ;
      RECT 44.775 0.79 44.925 0.94 ;
      RECT 44.655 1.36 44.805 1.51 ;
      RECT 43.575 1.055 43.725 1.205 ;
      RECT 43.24 1.775 43.39 1.925 ;
      RECT 43.16 0.615 43.31 0.765 ;
      RECT 41.725 1.01 41.875 1.16 ;
      RECT 40.96 0.86 41.11 1.01 ;
      RECT 40.705 0.455 40.855 0.605 ;
      RECT 40.085 1.22 40.235 1.37 ;
      RECT 39.705 0.69 39.855 0.84 ;
      RECT 39.69 1.73 39.84 1.88 ;
      RECT 39.16 0.995 39.31 1.145 ;
      RECT 39 1.715 39.15 1.865 ;
      RECT 38.19 0.995 38.34 1.145 ;
      RECT 37.375 0.475 37.525 0.625 ;
      RECT 37.215 1.86 37.365 2.01 ;
      RECT 36.98 1.515 37.13 1.665 ;
      RECT 36.935 0.905 37.085 1.055 ;
      RECT 35.935 1.525 36.085 1.675 ;
      RECT 34.845 1.47 34.995 1.62 ;
      RECT 33.99 0.53 34.14 0.68 ;
      RECT 31.625 1.57 31.775 1.72 ;
      RECT 25.185 1.47 25.335 1.62 ;
      RECT 24.33 0.6 24.48 0.75 ;
      RECT 23.86 0.45 24.01 0.6 ;
      RECT 21.05 1.47 21.2 1.62 ;
      RECT 19.79 0.54 19.94 0.69 ;
      RECT 19.375 1.26 19.525 1.41 ;
      RECT 17.7 -0.07 17.85 0.08 ;
      RECT 17.18 0.79 17.33 0.94 ;
      RECT 17.06 1.36 17.21 1.51 ;
      RECT 15.98 1.055 16.13 1.205 ;
      RECT 15.645 1.775 15.795 1.925 ;
      RECT 15.565 0.615 15.715 0.765 ;
      RECT 14.13 1.01 14.28 1.16 ;
      RECT 13.365 0.86 13.515 1.01 ;
      RECT 13.11 0.455 13.26 0.605 ;
      RECT 12.49 1.22 12.64 1.37 ;
      RECT 12.11 0.69 12.26 0.84 ;
      RECT 12.095 1.73 12.245 1.88 ;
      RECT 11.565 0.995 11.715 1.145 ;
      RECT 11.405 1.715 11.555 1.865 ;
      RECT 10.595 0.995 10.745 1.145 ;
      RECT 9.78 0.475 9.93 0.625 ;
      RECT 9.62 1.86 9.77 2.01 ;
      RECT 9.385 1.515 9.535 1.665 ;
      RECT 9.34 0.905 9.49 1.055 ;
      RECT 8.34 1.525 8.49 1.675 ;
      RECT 7.25 1.47 7.4 1.62 ;
      RECT 6.395 0.53 6.545 0.68 ;
      RECT 4.03 1.57 4.18 1.72 ;
      RECT 2.035 0.705 2.185 0.855 ;
    LAYER met1 ;
      RECT 0 2.48 141.925 2.96 ;
      RECT 2.455 1.67 2.63 2.96 ;
      RECT 2.395 1.67 2.685 1.9 ;
      RECT 128.16 1.885 128.465 2.115 ;
      RECT 136.3 1.915 139.715 2.09 ;
      RECT 139.54 1.065 139.715 2.09 ;
      RECT 128.16 1.915 139.715 2.085 ;
      RECT 139.485 1.065 139.815 1.315 ;
      RECT 136.745 1.075 137.035 1.315 ;
      RECT 132.295 1.045 132.555 1.28 ;
      RECT 132.295 1.075 137.035 1.245 ;
      RECT 135.48 1.415 135.8 1.675 ;
      RECT 135.465 1.46 135.8 1.63 ;
      RECT 134.185 0.395 134.48 0.685 ;
      RECT 134.15 0.395 134.48 0.655 ;
      RECT 131.345 1.415 131.665 1.675 ;
      RECT 131.33 1.46 131.665 1.63 ;
      RECT 129.67 1.205 129.99 1.465 ;
      RECT 129.655 1.205 130.01 1.44 ;
      RECT 126.97 0.965 127.155 1.175 ;
      RECT 126.96 0.97 127.17 1.168 ;
      RECT 126.96 0.97 127.256 1.145 ;
      RECT 126.96 0.97 127.315 1.12 ;
      RECT 126.96 0.97 127.37 1.1 ;
      RECT 126.96 0.97 127.38 1.088 ;
      RECT 126.96 0.97 127.575 1.027 ;
      RECT 126.96 0.97 127.605 1.01 ;
      RECT 126.96 0.97 127.625 1 ;
      RECT 127.505 0.735 127.765 0.995 ;
      RECT 127.49 0.825 127.505 1.042 ;
      RECT 127.025 0.957 127.765 0.995 ;
      RECT 127.476 0.836 127.49 1.048 ;
      RECT 127.065 0.95 127.765 0.995 ;
      RECT 127.39 0.876 127.476 1.067 ;
      RECT 127.315 0.937 127.765 0.995 ;
      RECT 127.385 0.912 127.39 1.084 ;
      RECT 127.37 0.922 127.765 0.995 ;
      RECT 127.38 0.917 127.385 1.086 ;
      RECT 127.675 1.422 127.68 1.514 ;
      RECT 127.67 1.4 127.675 1.531 ;
      RECT 127.665 1.39 127.67 1.543 ;
      RECT 127.655 1.381 127.665 1.553 ;
      RECT 127.65 1.376 127.655 1.561 ;
      RECT 127.645 1.372 127.65 1.564 ;
      RECT 127.611 1.305 127.645 1.575 ;
      RECT 127.525 1.305 127.611 1.61 ;
      RECT 127.445 1.305 127.525 1.658 ;
      RECT 127.385 1.305 127.445 1.683 ;
      RECT 127.325 1.405 127.385 1.69 ;
      RECT 127.29 1.43 127.325 1.696 ;
      RECT 127.265 1.445 127.29 1.7 ;
      RECT 127.251 1.454 127.265 1.702 ;
      RECT 127.165 1.481 127.251 1.708 ;
      RECT 127.1 1.522 127.165 1.717 ;
      RECT 127.085 1.542 127.1 1.722 ;
      RECT 127.055 1.552 127.085 1.725 ;
      RECT 127.05 1.562 127.055 1.728 ;
      RECT 127.02 1.567 127.05 1.73 ;
      RECT 127 1.572 127.02 1.734 ;
      RECT 126.915 1.575 127 1.741 ;
      RECT 126.9 1.572 126.915 1.747 ;
      RECT 126.89 1.569 126.9 1.749 ;
      RECT 126.87 1.566 126.89 1.751 ;
      RECT 126.85 1.562 126.87 1.752 ;
      RECT 126.835 1.558 126.85 1.754 ;
      RECT 126.825 1.555 126.835 1.755 ;
      RECT 126.785 1.549 126.825 1.753 ;
      RECT 126.775 1.544 126.785 1.751 ;
      RECT 126.76 1.541 126.775 1.747 ;
      RECT 126.735 1.536 126.76 1.74 ;
      RECT 126.685 1.527 126.735 1.728 ;
      RECT 126.615 1.513 126.685 1.71 ;
      RECT 126.557 1.498 126.615 1.692 ;
      RECT 126.471 1.481 126.557 1.672 ;
      RECT 126.385 1.46 126.471 1.647 ;
      RECT 126.335 1.445 126.385 1.628 ;
      RECT 126.331 1.439 126.335 1.62 ;
      RECT 126.245 1.429 126.331 1.607 ;
      RECT 126.21 1.414 126.245 1.59 ;
      RECT 126.195 1.407 126.21 1.583 ;
      RECT 126.135 1.395 126.195 1.571 ;
      RECT 126.115 1.382 126.135 1.559 ;
      RECT 126.075 1.373 126.115 1.551 ;
      RECT 126.07 1.365 126.075 1.544 ;
      RECT 125.99 1.355 126.07 1.53 ;
      RECT 125.975 1.342 125.99 1.515 ;
      RECT 125.97 1.34 125.975 1.513 ;
      RECT 125.891 1.328 125.97 1.5 ;
      RECT 125.805 1.303 125.891 1.475 ;
      RECT 125.79 1.272 125.805 1.46 ;
      RECT 125.775 1.247 125.79 1.456 ;
      RECT 125.76 1.24 125.775 1.452 ;
      RECT 125.585 1.245 125.59 1.448 ;
      RECT 125.58 1.25 125.585 1.443 ;
      RECT 125.59 1.24 125.76 1.45 ;
      RECT 126.305 1 126.41 1.26 ;
      RECT 127.12 0.525 127.125 0.75 ;
      RECT 127.25 0.525 127.305 0.735 ;
      RECT 127.305 0.53 127.315 0.728 ;
      RECT 127.211 0.525 127.25 0.738 ;
      RECT 127.125 0.525 127.211 0.745 ;
      RECT 127.105 0.53 127.12 0.751 ;
      RECT 127.095 0.57 127.105 0.753 ;
      RECT 127.065 0.58 127.095 0.755 ;
      RECT 127.06 0.585 127.065 0.757 ;
      RECT 127.035 0.59 127.06 0.759 ;
      RECT 127.02 0.595 127.035 0.761 ;
      RECT 127.005 0.597 127.02 0.763 ;
      RECT 127 0.602 127.005 0.765 ;
      RECT 126.95 0.61 127 0.768 ;
      RECT 126.925 0.619 126.95 0.773 ;
      RECT 126.915 0.626 126.925 0.778 ;
      RECT 126.91 0.629 126.915 0.782 ;
      RECT 126.89 0.632 126.91 0.791 ;
      RECT 126.86 0.64 126.89 0.811 ;
      RECT 126.831 0.653 126.86 0.833 ;
      RECT 126.745 0.687 126.831 0.877 ;
      RECT 126.74 0.713 126.745 0.915 ;
      RECT 126.735 0.717 126.74 0.924 ;
      RECT 126.7 0.73 126.735 0.957 ;
      RECT 126.69 0.744 126.7 0.995 ;
      RECT 126.685 0.748 126.69 1.008 ;
      RECT 126.68 0.752 126.685 1.013 ;
      RECT 126.67 0.76 126.68 1.025 ;
      RECT 126.665 0.767 126.67 1.04 ;
      RECT 126.64 0.78 126.665 1.065 ;
      RECT 126.6 0.809 126.64 1.12 ;
      RECT 126.585 0.834 126.6 1.175 ;
      RECT 126.575 0.845 126.585 1.198 ;
      RECT 126.57 0.852 126.575 1.21 ;
      RECT 126.565 0.856 126.57 1.218 ;
      RECT 126.51 0.884 126.565 1.26 ;
      RECT 126.49 0.92 126.51 1.26 ;
      RECT 126.475 0.935 126.49 1.26 ;
      RECT 126.42 0.967 126.475 1.26 ;
      RECT 126.41 0.997 126.42 1.26 ;
      RECT 126.02 0.612 126.205 0.85 ;
      RECT 126.005 0.614 126.215 0.845 ;
      RECT 125.89 0.56 126.15 0.82 ;
      RECT 125.885 0.597 126.15 0.774 ;
      RECT 125.88 0.607 126.15 0.771 ;
      RECT 125.875 0.647 126.215 0.765 ;
      RECT 125.87 0.68 126.215 0.755 ;
      RECT 125.88 0.622 126.23 0.693 ;
      RECT 126.177 1.72 126.19 2.25 ;
      RECT 126.091 1.72 126.19 2.249 ;
      RECT 126.091 1.72 126.195 2.248 ;
      RECT 126.005 1.72 126.195 2.246 ;
      RECT 126 1.72 126.195 2.243 ;
      RECT 126 1.72 126.205 2.241 ;
      RECT 125.995 2.012 126.205 2.238 ;
      RECT 125.995 2.022 126.21 2.235 ;
      RECT 125.995 2.09 126.215 2.231 ;
      RECT 125.985 2.095 126.215 2.23 ;
      RECT 125.985 2.187 126.22 2.227 ;
      RECT 125.97 1.72 126.23 1.98 ;
      RECT 125.2 0.71 125.245 2.245 ;
      RECT 125.4 0.71 125.43 0.925 ;
      RECT 123.775 0.45 123.895 0.66 ;
      RECT 123.435 0.4 123.695 0.66 ;
      RECT 123.435 0.445 123.73 0.65 ;
      RECT 125.44 0.726 125.445 0.78 ;
      RECT 125.435 0.719 125.44 0.913 ;
      RECT 125.43 0.713 125.435 0.92 ;
      RECT 125.385 0.71 125.4 0.933 ;
      RECT 125.38 0.71 125.385 0.955 ;
      RECT 125.375 0.71 125.38 1.003 ;
      RECT 125.37 0.71 125.375 1.023 ;
      RECT 125.36 0.71 125.37 1.13 ;
      RECT 125.355 0.71 125.36 1.193 ;
      RECT 125.35 0.71 125.355 1.25 ;
      RECT 125.345 0.71 125.35 1.258 ;
      RECT 125.33 0.71 125.345 1.365 ;
      RECT 125.32 0.71 125.33 1.5 ;
      RECT 125.31 0.71 125.32 1.61 ;
      RECT 125.3 0.71 125.31 1.667 ;
      RECT 125.295 0.71 125.3 1.707 ;
      RECT 125.29 0.71 125.295 1.743 ;
      RECT 125.28 0.71 125.29 1.783 ;
      RECT 125.275 0.71 125.28 1.825 ;
      RECT 125.255 0.71 125.275 1.89 ;
      RECT 125.26 2.035 125.265 2.215 ;
      RECT 125.255 2.017 125.26 2.223 ;
      RECT 125.25 0.71 125.255 1.953 ;
      RECT 125.25 1.997 125.255 2.23 ;
      RECT 125.245 0.71 125.25 2.24 ;
      RECT 125.19 0.71 125.2 1.01 ;
      RECT 125.195 1.257 125.2 2.245 ;
      RECT 125.19 1.322 125.195 2.245 ;
      RECT 125.185 0.711 125.19 1 ;
      RECT 125.18 1.387 125.19 2.245 ;
      RECT 125.175 0.712 125.185 0.99 ;
      RECT 125.165 1.5 125.18 2.245 ;
      RECT 125.17 0.713 125.175 0.98 ;
      RECT 125.15 0.714 125.17 0.958 ;
      RECT 125.155 1.597 125.165 2.245 ;
      RECT 125.15 1.672 125.155 2.245 ;
      RECT 125.14 0.713 125.15 0.935 ;
      RECT 125.145 1.715 125.15 2.245 ;
      RECT 125.14 1.742 125.145 2.245 ;
      RECT 125.13 0.711 125.14 0.923 ;
      RECT 125.135 1.785 125.14 2.245 ;
      RECT 125.13 1.812 125.135 2.245 ;
      RECT 125.12 0.71 125.13 0.91 ;
      RECT 125.125 1.827 125.13 2.245 ;
      RECT 125.085 1.885 125.125 2.245 ;
      RECT 125.115 0.709 125.12 0.895 ;
      RECT 125.11 0.707 125.115 0.888 ;
      RECT 125.1 0.704 125.11 0.878 ;
      RECT 125.095 0.701 125.1 0.863 ;
      RECT 125.08 0.697 125.095 0.856 ;
      RECT 125.075 1.94 125.085 2.245 ;
      RECT 125.075 0.694 125.08 0.851 ;
      RECT 125.06 0.69 125.075 0.845 ;
      RECT 125.07 1.957 125.075 2.245 ;
      RECT 125.06 2.02 125.07 2.245 ;
      RECT 124.98 0.675 125.06 0.825 ;
      RECT 125.055 2.027 125.06 2.24 ;
      RECT 125.05 2.035 125.055 2.23 ;
      RECT 124.97 0.661 124.98 0.809 ;
      RECT 124.955 0.657 124.97 0.807 ;
      RECT 124.945 0.652 124.955 0.803 ;
      RECT 124.92 0.645 124.945 0.795 ;
      RECT 124.915 0.64 124.92 0.79 ;
      RECT 124.905 0.64 124.915 0.788 ;
      RECT 124.895 0.638 124.905 0.786 ;
      RECT 124.865 0.63 124.895 0.78 ;
      RECT 124.85 0.622 124.865 0.773 ;
      RECT 124.83 0.617 124.85 0.766 ;
      RECT 124.825 0.613 124.83 0.761 ;
      RECT 124.795 0.606 124.825 0.755 ;
      RECT 124.77 0.597 124.795 0.745 ;
      RECT 124.74 0.59 124.77 0.737 ;
      RECT 124.715 0.58 124.74 0.728 ;
      RECT 124.7 0.572 124.715 0.722 ;
      RECT 124.675 0.567 124.7 0.717 ;
      RECT 124.665 0.563 124.675 0.712 ;
      RECT 124.645 0.558 124.665 0.707 ;
      RECT 124.61 0.553 124.645 0.7 ;
      RECT 124.55 0.548 124.61 0.693 ;
      RECT 124.537 0.544 124.55 0.691 ;
      RECT 124.451 0.539 124.537 0.688 ;
      RECT 124.365 0.529 124.451 0.684 ;
      RECT 124.324 0.522 124.365 0.681 ;
      RECT 124.238 0.515 124.324 0.678 ;
      RECT 124.152 0.505 124.238 0.674 ;
      RECT 124.066 0.495 124.152 0.669 ;
      RECT 123.98 0.485 124.066 0.665 ;
      RECT 123.97 0.47 123.98 0.663 ;
      RECT 123.96 0.455 123.97 0.663 ;
      RECT 123.895 0.45 123.96 0.662 ;
      RECT 123.73 0.447 123.775 0.655 ;
      RECT 124.975 1.352 124.98 1.543 ;
      RECT 124.97 1.347 124.975 1.55 ;
      RECT 124.956 1.345 124.97 1.556 ;
      RECT 124.87 1.345 124.956 1.558 ;
      RECT 124.866 1.345 124.87 1.561 ;
      RECT 124.78 1.345 124.866 1.579 ;
      RECT 124.77 1.35 124.78 1.598 ;
      RECT 124.76 1.405 124.77 1.602 ;
      RECT 124.735 1.42 124.76 1.609 ;
      RECT 124.695 1.44 124.735 1.622 ;
      RECT 124.69 1.452 124.695 1.632 ;
      RECT 124.675 1.458 124.69 1.637 ;
      RECT 124.67 1.463 124.675 1.641 ;
      RECT 124.65 1.47 124.67 1.646 ;
      RECT 124.58 1.495 124.65 1.663 ;
      RECT 124.54 1.523 124.58 1.683 ;
      RECT 124.535 1.533 124.54 1.691 ;
      RECT 124.515 1.54 124.535 1.693 ;
      RECT 124.51 1.547 124.515 1.696 ;
      RECT 124.48 1.555 124.51 1.699 ;
      RECT 124.475 1.56 124.48 1.703 ;
      RECT 124.401 1.564 124.475 1.711 ;
      RECT 124.315 1.573 124.401 1.727 ;
      RECT 124.311 1.578 124.315 1.736 ;
      RECT 124.225 1.583 124.311 1.746 ;
      RECT 124.185 1.591 124.225 1.758 ;
      RECT 124.135 1.597 124.185 1.765 ;
      RECT 124.05 1.606 124.135 1.78 ;
      RECT 123.975 1.617 124.05 1.798 ;
      RECT 123.94 1.624 123.975 1.808 ;
      RECT 123.865 1.632 123.94 1.813 ;
      RECT 123.81 1.641 123.865 1.813 ;
      RECT 123.785 1.646 123.81 1.811 ;
      RECT 123.775 1.649 123.785 1.809 ;
      RECT 123.74 1.651 123.775 1.807 ;
      RECT 123.71 1.653 123.74 1.803 ;
      RECT 123.665 1.652 123.71 1.799 ;
      RECT 123.645 1.647 123.665 1.796 ;
      RECT 123.595 1.632 123.645 1.793 ;
      RECT 123.585 1.617 123.595 1.788 ;
      RECT 123.535 1.602 123.585 1.778 ;
      RECT 123.485 1.577 123.535 1.758 ;
      RECT 123.475 1.562 123.485 1.74 ;
      RECT 123.47 1.56 123.475 1.734 ;
      RECT 123.45 1.555 123.47 1.729 ;
      RECT 123.445 1.547 123.45 1.723 ;
      RECT 123.43 1.541 123.445 1.716 ;
      RECT 123.425 1.536 123.43 1.708 ;
      RECT 123.405 1.531 123.425 1.7 ;
      RECT 123.39 1.524 123.405 1.693 ;
      RECT 123.375 1.518 123.39 1.684 ;
      RECT 123.37 1.512 123.375 1.677 ;
      RECT 123.325 1.487 123.37 1.663 ;
      RECT 123.31 1.457 123.325 1.645 ;
      RECT 123.295 1.44 123.31 1.636 ;
      RECT 123.27 1.42 123.295 1.624 ;
      RECT 123.23 1.39 123.27 1.604 ;
      RECT 123.22 1.36 123.23 1.589 ;
      RECT 123.205 1.35 123.22 1.582 ;
      RECT 123.15 1.315 123.205 1.561 ;
      RECT 123.135 1.278 123.15 1.54 ;
      RECT 123.125 1.265 123.135 1.532 ;
      RECT 123.075 1.235 123.125 1.514 ;
      RECT 123.06 1.165 123.075 1.495 ;
      RECT 123.015 1.165 123.06 1.478 ;
      RECT 122.99 1.165 123.015 1.46 ;
      RECT 122.98 1.165 122.99 1.453 ;
      RECT 122.901 1.165 122.98 1.446 ;
      RECT 122.815 1.165 122.901 1.438 ;
      RECT 122.8 1.197 122.815 1.433 ;
      RECT 122.725 1.207 122.8 1.429 ;
      RECT 122.705 1.217 122.725 1.424 ;
      RECT 122.68 1.217 122.705 1.421 ;
      RECT 122.67 1.207 122.68 1.42 ;
      RECT 122.66 1.18 122.67 1.419 ;
      RECT 122.62 1.175 122.66 1.417 ;
      RECT 122.575 1.175 122.62 1.413 ;
      RECT 122.55 1.175 122.575 1.408 ;
      RECT 122.5 1.175 122.55 1.395 ;
      RECT 122.46 1.18 122.47 1.38 ;
      RECT 122.47 1.175 122.5 1.385 ;
      RECT 124.455 0.955 124.715 1.215 ;
      RECT 124.45 0.977 124.715 1.173 ;
      RECT 123.69 0.805 123.91 1.17 ;
      RECT 123.672 0.892 123.91 1.169 ;
      RECT 123.655 0.897 123.91 1.166 ;
      RECT 123.655 0.897 123.93 1.165 ;
      RECT 123.625 0.907 123.93 1.163 ;
      RECT 123.62 0.922 123.93 1.159 ;
      RECT 123.62 0.922 123.935 1.158 ;
      RECT 123.615 0.98 123.935 1.156 ;
      RECT 123.615 0.98 123.945 1.153 ;
      RECT 123.61 1.045 123.945 1.148 ;
      RECT 123.69 0.805 123.95 1.065 ;
      RECT 122.435 0.635 122.695 0.895 ;
      RECT 122.435 0.678 122.781 0.869 ;
      RECT 122.435 0.678 122.825 0.868 ;
      RECT 122.435 0.678 122.845 0.866 ;
      RECT 122.435 0.678 122.945 0.865 ;
      RECT 122.435 0.678 122.965 0.863 ;
      RECT 122.435 0.678 122.975 0.858 ;
      RECT 122.845 0.645 123.035 0.855 ;
      RECT 122.845 0.647 123.04 0.853 ;
      RECT 122.835 0.652 123.045 0.845 ;
      RECT 122.781 0.676 123.045 0.845 ;
      RECT 122.825 0.67 122.835 0.867 ;
      RECT 122.835 0.65 123.04 0.853 ;
      RECT 121.79 1.71 121.995 1.94 ;
      RECT 121.73 1.66 121.785 1.92 ;
      RECT 121.79 1.66 121.99 1.94 ;
      RECT 122.76 1.975 122.765 2.002 ;
      RECT 122.75 1.885 122.76 2.007 ;
      RECT 122.745 1.807 122.75 2.013 ;
      RECT 122.735 1.797 122.745 2.02 ;
      RECT 122.73 1.787 122.735 2.026 ;
      RECT 122.72 1.782 122.73 2.028 ;
      RECT 122.705 1.774 122.72 2.036 ;
      RECT 122.69 1.765 122.705 2.048 ;
      RECT 122.68 1.757 122.69 2.058 ;
      RECT 122.645 1.675 122.68 2.076 ;
      RECT 122.61 1.675 122.645 2.095 ;
      RECT 122.595 1.675 122.61 2.103 ;
      RECT 122.54 1.675 122.595 2.103 ;
      RECT 122.506 1.675 122.54 2.094 ;
      RECT 122.42 1.675 122.506 2.07 ;
      RECT 122.41 1.735 122.42 2.052 ;
      RECT 122.37 1.737 122.41 2.043 ;
      RECT 122.365 1.739 122.37 2.033 ;
      RECT 122.345 1.741 122.365 2.028 ;
      RECT 122.335 1.744 122.345 2.023 ;
      RECT 122.325 1.745 122.335 2.018 ;
      RECT 122.301 1.746 122.325 2.01 ;
      RECT 122.215 1.751 122.301 1.988 ;
      RECT 122.16 1.75 122.215 1.961 ;
      RECT 122.145 1.743 122.16 1.948 ;
      RECT 122.11 1.738 122.145 1.944 ;
      RECT 122.055 1.73 122.11 1.943 ;
      RECT 121.995 1.717 122.055 1.941 ;
      RECT 121.785 1.66 121.79 1.928 ;
      RECT 121.86 1.03 122.045 1.24 ;
      RECT 121.85 1.035 122.06 1.233 ;
      RECT 121.89 0.94 122.15 1.2 ;
      RECT 121.845 1.097 122.15 1.123 ;
      RECT 121.19 0.89 121.195 1.69 ;
      RECT 121.135 0.94 121.165 1.69 ;
      RECT 121.125 0.94 121.13 1.25 ;
      RECT 121.11 0.94 121.115 1.245 ;
      RECT 120.655 0.985 120.67 1.2 ;
      RECT 120.585 0.985 120.67 1.195 ;
      RECT 121.85 0.565 121.92 0.775 ;
      RECT 121.92 0.572 121.93 0.77 ;
      RECT 121.816 0.565 121.85 0.782 ;
      RECT 121.73 0.565 121.816 0.806 ;
      RECT 121.72 0.57 121.73 0.825 ;
      RECT 121.715 0.582 121.72 0.828 ;
      RECT 121.7 0.597 121.715 0.832 ;
      RECT 121.695 0.615 121.7 0.836 ;
      RECT 121.655 0.625 121.695 0.845 ;
      RECT 121.64 0.632 121.655 0.857 ;
      RECT 121.625 0.637 121.64 0.862 ;
      RECT 121.61 0.64 121.625 0.867 ;
      RECT 121.6 0.642 121.61 0.871 ;
      RECT 121.565 0.649 121.6 0.879 ;
      RECT 121.53 0.657 121.565 0.893 ;
      RECT 121.52 0.663 121.53 0.902 ;
      RECT 121.515 0.665 121.52 0.904 ;
      RECT 121.495 0.668 121.515 0.91 ;
      RECT 121.465 0.675 121.495 0.921 ;
      RECT 121.455 0.681 121.465 0.928 ;
      RECT 121.43 0.684 121.455 0.935 ;
      RECT 121.42 0.688 121.43 0.943 ;
      RECT 121.415 0.689 121.42 0.965 ;
      RECT 121.41 0.69 121.415 0.98 ;
      RECT 121.405 0.691 121.41 0.995 ;
      RECT 121.4 0.692 121.405 1.01 ;
      RECT 121.395 0.693 121.4 1.04 ;
      RECT 121.385 0.695 121.395 1.073 ;
      RECT 121.37 0.699 121.385 1.12 ;
      RECT 121.36 0.702 121.37 1.165 ;
      RECT 121.355 0.705 121.36 1.193 ;
      RECT 121.345 0.707 121.355 1.22 ;
      RECT 121.34 0.71 121.345 1.255 ;
      RECT 121.31 0.715 121.34 1.313 ;
      RECT 121.305 0.72 121.31 1.398 ;
      RECT 121.3 0.722 121.305 1.433 ;
      RECT 121.295 0.724 121.3 1.515 ;
      RECT 121.29 0.726 121.295 1.603 ;
      RECT 121.28 0.728 121.29 1.685 ;
      RECT 121.265 0.742 121.28 1.69 ;
      RECT 121.23 0.787 121.265 1.69 ;
      RECT 121.22 0.827 121.23 1.69 ;
      RECT 121.205 0.855 121.22 1.69 ;
      RECT 121.2 0.872 121.205 1.69 ;
      RECT 121.195 0.88 121.2 1.69 ;
      RECT 121.185 0.895 121.19 1.69 ;
      RECT 121.18 0.902 121.185 1.69 ;
      RECT 121.17 0.922 121.18 1.69 ;
      RECT 121.165 0.935 121.17 1.69 ;
      RECT 121.13 0.94 121.135 1.275 ;
      RECT 121.115 1.33 121.135 1.69 ;
      RECT 121.115 0.94 121.125 1.248 ;
      RECT 121.11 1.37 121.115 1.69 ;
      RECT 121.06 0.94 121.11 1.243 ;
      RECT 121.105 1.407 121.11 1.69 ;
      RECT 121.095 1.43 121.105 1.69 ;
      RECT 121.09 1.475 121.095 1.69 ;
      RECT 121.08 1.485 121.09 1.683 ;
      RECT 121.006 0.94 121.06 1.237 ;
      RECT 120.92 0.94 121.006 1.23 ;
      RECT 120.871 0.987 120.92 1.223 ;
      RECT 120.785 0.995 120.871 1.216 ;
      RECT 120.77 0.992 120.785 1.211 ;
      RECT 120.756 0.985 120.77 1.21 ;
      RECT 120.67 0.985 120.756 1.205 ;
      RECT 120.575 0.99 120.585 1.19 ;
      RECT 120.165 0.42 120.18 0.82 ;
      RECT 120.36 0.42 120.365 0.68 ;
      RECT 120.105 0.42 120.15 0.68 ;
      RECT 120.56 1.725 120.565 1.93 ;
      RECT 120.555 1.715 120.56 1.935 ;
      RECT 120.55 1.702 120.555 1.94 ;
      RECT 120.545 1.682 120.55 1.94 ;
      RECT 120.52 1.635 120.545 1.94 ;
      RECT 120.485 1.55 120.52 1.94 ;
      RECT 120.48 1.487 120.485 1.94 ;
      RECT 120.475 1.472 120.48 1.94 ;
      RECT 120.46 1.432 120.475 1.94 ;
      RECT 120.455 1.407 120.46 1.94 ;
      RECT 120.445 1.39 120.455 1.94 ;
      RECT 120.41 1.312 120.445 1.94 ;
      RECT 120.405 1.255 120.41 1.94 ;
      RECT 120.4 1.242 120.405 1.94 ;
      RECT 120.39 1.22 120.4 1.94 ;
      RECT 120.38 1.185 120.39 1.94 ;
      RECT 120.37 1.155 120.38 1.94 ;
      RECT 120.36 1.07 120.37 1.583 ;
      RECT 120.367 1.715 120.37 1.94 ;
      RECT 120.365 1.725 120.367 1.94 ;
      RECT 120.355 1.735 120.365 1.935 ;
      RECT 120.35 0.42 120.36 0.815 ;
      RECT 120.355 0.947 120.36 1.558 ;
      RECT 120.35 0.845 120.355 1.541 ;
      RECT 120.34 0.42 120.35 1.517 ;
      RECT 120.335 0.42 120.34 1.488 ;
      RECT 120.33 0.42 120.335 1.478 ;
      RECT 120.31 0.42 120.33 1.44 ;
      RECT 120.305 0.42 120.31 1.398 ;
      RECT 120.3 0.42 120.305 1.378 ;
      RECT 120.27 0.42 120.3 1.328 ;
      RECT 120.26 0.42 120.27 1.275 ;
      RECT 120.255 0.42 120.26 1.248 ;
      RECT 120.25 0.42 120.255 1.233 ;
      RECT 120.24 0.42 120.25 1.21 ;
      RECT 120.23 0.42 120.24 1.185 ;
      RECT 120.225 0.42 120.23 1.125 ;
      RECT 120.215 0.42 120.225 1.063 ;
      RECT 120.21 0.42 120.215 0.983 ;
      RECT 120.205 0.42 120.21 0.948 ;
      RECT 120.2 0.42 120.205 0.923 ;
      RECT 120.195 0.42 120.2 0.908 ;
      RECT 120.19 0.42 120.195 0.878 ;
      RECT 120.185 0.42 120.19 0.855 ;
      RECT 120.18 0.42 120.185 0.828 ;
      RECT 120.15 0.42 120.165 0.815 ;
      RECT 119.305 1.955 119.49 2.165 ;
      RECT 119.295 1.96 119.505 2.158 ;
      RECT 119.295 1.96 119.525 2.13 ;
      RECT 119.295 1.96 119.54 2.109 ;
      RECT 119.295 1.96 119.555 2.107 ;
      RECT 119.295 1.96 119.565 2.106 ;
      RECT 119.295 1.96 119.595 2.103 ;
      RECT 119.945 1.805 120.205 2.065 ;
      RECT 119.905 1.852 120.205 2.048 ;
      RECT 119.896 1.86 119.905 2.051 ;
      RECT 119.49 1.953 120.205 2.048 ;
      RECT 119.81 1.878 119.896 2.058 ;
      RECT 119.505 1.95 120.205 2.048 ;
      RECT 119.751 1.9 119.81 2.07 ;
      RECT 119.525 1.946 120.205 2.048 ;
      RECT 119.665 1.912 119.751 2.081 ;
      RECT 119.54 1.942 120.205 2.048 ;
      RECT 119.61 1.925 119.665 2.093 ;
      RECT 119.555 1.94 120.205 2.048 ;
      RECT 119.595 1.931 119.61 2.099 ;
      RECT 119.565 1.936 120.205 2.048 ;
      RECT 119.71 1.46 119.97 1.72 ;
      RECT 119.71 1.48 120.08 1.69 ;
      RECT 119.71 1.485 120.09 1.685 ;
      RECT 119.901 0.899 119.98 1.13 ;
      RECT 119.815 0.902 120.03 1.125 ;
      RECT 119.81 0.902 120.03 1.12 ;
      RECT 119.81 0.907 120.04 1.118 ;
      RECT 119.785 0.907 120.04 1.115 ;
      RECT 119.785 0.915 120.05 1.113 ;
      RECT 119.665 0.85 119.925 1.11 ;
      RECT 119.665 0.897 119.975 1.11 ;
      RECT 118.92 1.47 118.925 1.73 ;
      RECT 118.75 1.24 118.755 1.73 ;
      RECT 118.635 1.48 118.64 1.705 ;
      RECT 119.345 0.575 119.35 0.785 ;
      RECT 119.35 0.58 119.365 0.78 ;
      RECT 119.285 0.575 119.345 0.793 ;
      RECT 119.27 0.575 119.285 0.803 ;
      RECT 119.22 0.575 119.27 0.82 ;
      RECT 119.2 0.575 119.22 0.843 ;
      RECT 119.185 0.575 119.2 0.855 ;
      RECT 119.165 0.575 119.185 0.865 ;
      RECT 119.155 0.58 119.165 0.874 ;
      RECT 119.15 0.59 119.155 0.879 ;
      RECT 119.145 0.602 119.15 0.883 ;
      RECT 119.135 0.625 119.145 0.888 ;
      RECT 119.13 0.64 119.135 0.892 ;
      RECT 119.125 0.657 119.13 0.895 ;
      RECT 119.12 0.665 119.125 0.898 ;
      RECT 119.11 0.67 119.12 0.902 ;
      RECT 119.105 0.677 119.11 0.907 ;
      RECT 119.095 0.682 119.105 0.911 ;
      RECT 119.07 0.694 119.095 0.922 ;
      RECT 119.05 0.711 119.07 0.938 ;
      RECT 119.025 0.728 119.05 0.96 ;
      RECT 118.99 0.751 119.025 1.018 ;
      RECT 118.97 0.773 118.99 1.08 ;
      RECT 118.965 0.783 118.97 1.115 ;
      RECT 118.955 0.79 118.965 1.153 ;
      RECT 118.95 0.797 118.955 1.173 ;
      RECT 118.945 0.808 118.95 1.21 ;
      RECT 118.94 0.816 118.945 1.275 ;
      RECT 118.93 0.827 118.94 1.328 ;
      RECT 118.925 0.845 118.93 1.398 ;
      RECT 118.92 0.855 118.925 1.435 ;
      RECT 118.915 0.865 118.92 1.73 ;
      RECT 118.91 0.877 118.915 1.73 ;
      RECT 118.905 0.887 118.91 1.73 ;
      RECT 118.895 0.897 118.905 1.73 ;
      RECT 118.885 0.92 118.895 1.73 ;
      RECT 118.87 0.955 118.885 1.73 ;
      RECT 118.83 1.017 118.87 1.73 ;
      RECT 118.825 1.07 118.83 1.73 ;
      RECT 118.8 1.105 118.825 1.73 ;
      RECT 118.785 1.15 118.8 1.73 ;
      RECT 118.78 1.172 118.785 1.73 ;
      RECT 118.77 1.185 118.78 1.73 ;
      RECT 118.76 1.21 118.77 1.73 ;
      RECT 118.755 1.232 118.76 1.73 ;
      RECT 118.73 1.27 118.75 1.73 ;
      RECT 118.69 1.327 118.73 1.73 ;
      RECT 118.685 1.377 118.69 1.73 ;
      RECT 118.68 1.395 118.685 1.73 ;
      RECT 118.675 1.407 118.68 1.73 ;
      RECT 118.665 1.425 118.675 1.73 ;
      RECT 118.655 1.445 118.665 1.705 ;
      RECT 118.65 1.462 118.655 1.705 ;
      RECT 118.64 1.475 118.65 1.705 ;
      RECT 118.61 1.485 118.635 1.705 ;
      RECT 118.6 1.492 118.61 1.705 ;
      RECT 118.585 1.502 118.6 1.7 ;
      RECT 117.545 1.415 117.865 1.675 ;
      RECT 117.41 1.46 117.865 1.63 ;
      RECT 111.07 1.515 111.445 1.765 ;
      RECT 111.17 0.73 111.345 1.765 ;
      RECT 111.17 0.73 117.095 0.905 ;
      RECT 116.69 0.475 117.01 0.905 ;
      RECT 116.69 0.505 117.09 0.675 ;
      RECT 114.355 1.515 114.65 1.805 ;
      RECT 114.325 1.515 114.65 1.775 ;
      RECT 100.565 1.885 100.87 2.115 ;
      RECT 108.705 1.915 112.12 2.09 ;
      RECT 111.945 1.065 112.12 2.09 ;
      RECT 100.565 1.915 112.12 2.085 ;
      RECT 111.89 1.065 112.22 1.315 ;
      RECT 109.15 1.075 109.44 1.315 ;
      RECT 104.7 1.045 104.96 1.28 ;
      RECT 104.7 1.075 109.44 1.245 ;
      RECT 107.885 1.415 108.205 1.675 ;
      RECT 107.87 1.46 108.205 1.63 ;
      RECT 106.59 0.395 106.885 0.685 ;
      RECT 106.555 0.395 106.885 0.655 ;
      RECT 103.75 1.415 104.07 1.675 ;
      RECT 103.735 1.46 104.07 1.63 ;
      RECT 102.075 1.205 102.395 1.465 ;
      RECT 102.06 1.205 102.415 1.44 ;
      RECT 99.375 0.965 99.56 1.175 ;
      RECT 99.365 0.97 99.575 1.168 ;
      RECT 99.365 0.97 99.661 1.145 ;
      RECT 99.365 0.97 99.72 1.12 ;
      RECT 99.365 0.97 99.775 1.1 ;
      RECT 99.365 0.97 99.785 1.088 ;
      RECT 99.365 0.97 99.98 1.027 ;
      RECT 99.365 0.97 100.01 1.01 ;
      RECT 99.365 0.97 100.03 1 ;
      RECT 99.91 0.735 100.17 0.995 ;
      RECT 99.895 0.825 99.91 1.042 ;
      RECT 99.43 0.957 100.17 0.995 ;
      RECT 99.881 0.836 99.895 1.048 ;
      RECT 99.47 0.95 100.17 0.995 ;
      RECT 99.795 0.876 99.881 1.067 ;
      RECT 99.72 0.937 100.17 0.995 ;
      RECT 99.79 0.912 99.795 1.084 ;
      RECT 99.775 0.922 100.17 0.995 ;
      RECT 99.785 0.917 99.79 1.086 ;
      RECT 100.08 1.422 100.085 1.514 ;
      RECT 100.075 1.4 100.08 1.531 ;
      RECT 100.07 1.39 100.075 1.543 ;
      RECT 100.06 1.381 100.07 1.553 ;
      RECT 100.055 1.376 100.06 1.561 ;
      RECT 100.05 1.372 100.055 1.564 ;
      RECT 100.016 1.305 100.05 1.575 ;
      RECT 99.93 1.305 100.016 1.61 ;
      RECT 99.85 1.305 99.93 1.658 ;
      RECT 99.79 1.305 99.85 1.683 ;
      RECT 99.73 1.405 99.79 1.69 ;
      RECT 99.695 1.43 99.73 1.696 ;
      RECT 99.67 1.445 99.695 1.7 ;
      RECT 99.656 1.454 99.67 1.702 ;
      RECT 99.57 1.481 99.656 1.708 ;
      RECT 99.505 1.522 99.57 1.717 ;
      RECT 99.49 1.542 99.505 1.722 ;
      RECT 99.46 1.552 99.49 1.725 ;
      RECT 99.455 1.562 99.46 1.728 ;
      RECT 99.425 1.567 99.455 1.73 ;
      RECT 99.405 1.572 99.425 1.734 ;
      RECT 99.32 1.575 99.405 1.741 ;
      RECT 99.305 1.572 99.32 1.747 ;
      RECT 99.295 1.569 99.305 1.749 ;
      RECT 99.275 1.566 99.295 1.751 ;
      RECT 99.255 1.562 99.275 1.752 ;
      RECT 99.24 1.558 99.255 1.754 ;
      RECT 99.23 1.555 99.24 1.755 ;
      RECT 99.19 1.549 99.23 1.753 ;
      RECT 99.18 1.544 99.19 1.751 ;
      RECT 99.165 1.541 99.18 1.747 ;
      RECT 99.14 1.536 99.165 1.74 ;
      RECT 99.09 1.527 99.14 1.728 ;
      RECT 99.02 1.513 99.09 1.71 ;
      RECT 98.962 1.498 99.02 1.692 ;
      RECT 98.876 1.481 98.962 1.672 ;
      RECT 98.79 1.46 98.876 1.647 ;
      RECT 98.74 1.445 98.79 1.628 ;
      RECT 98.736 1.439 98.74 1.62 ;
      RECT 98.65 1.429 98.736 1.607 ;
      RECT 98.615 1.414 98.65 1.59 ;
      RECT 98.6 1.407 98.615 1.583 ;
      RECT 98.54 1.395 98.6 1.571 ;
      RECT 98.52 1.382 98.54 1.559 ;
      RECT 98.48 1.373 98.52 1.551 ;
      RECT 98.475 1.365 98.48 1.544 ;
      RECT 98.395 1.355 98.475 1.53 ;
      RECT 98.38 1.342 98.395 1.515 ;
      RECT 98.375 1.34 98.38 1.513 ;
      RECT 98.296 1.328 98.375 1.5 ;
      RECT 98.21 1.303 98.296 1.475 ;
      RECT 98.195 1.272 98.21 1.46 ;
      RECT 98.18 1.247 98.195 1.456 ;
      RECT 98.165 1.24 98.18 1.452 ;
      RECT 97.99 1.245 97.995 1.448 ;
      RECT 97.985 1.25 97.99 1.443 ;
      RECT 97.995 1.24 98.165 1.45 ;
      RECT 98.71 1 98.815 1.26 ;
      RECT 99.525 0.525 99.53 0.75 ;
      RECT 99.655 0.525 99.71 0.735 ;
      RECT 99.71 0.53 99.72 0.728 ;
      RECT 99.616 0.525 99.655 0.738 ;
      RECT 99.53 0.525 99.616 0.745 ;
      RECT 99.51 0.53 99.525 0.751 ;
      RECT 99.5 0.57 99.51 0.753 ;
      RECT 99.47 0.58 99.5 0.755 ;
      RECT 99.465 0.585 99.47 0.757 ;
      RECT 99.44 0.59 99.465 0.759 ;
      RECT 99.425 0.595 99.44 0.761 ;
      RECT 99.41 0.597 99.425 0.763 ;
      RECT 99.405 0.602 99.41 0.765 ;
      RECT 99.355 0.61 99.405 0.768 ;
      RECT 99.33 0.619 99.355 0.773 ;
      RECT 99.32 0.626 99.33 0.778 ;
      RECT 99.315 0.629 99.32 0.782 ;
      RECT 99.295 0.632 99.315 0.791 ;
      RECT 99.265 0.64 99.295 0.811 ;
      RECT 99.236 0.653 99.265 0.833 ;
      RECT 99.15 0.687 99.236 0.877 ;
      RECT 99.145 0.713 99.15 0.915 ;
      RECT 99.14 0.717 99.145 0.924 ;
      RECT 99.105 0.73 99.14 0.957 ;
      RECT 99.095 0.744 99.105 0.995 ;
      RECT 99.09 0.748 99.095 1.008 ;
      RECT 99.085 0.752 99.09 1.013 ;
      RECT 99.075 0.76 99.085 1.025 ;
      RECT 99.07 0.767 99.075 1.04 ;
      RECT 99.045 0.78 99.07 1.065 ;
      RECT 99.005 0.809 99.045 1.12 ;
      RECT 98.99 0.834 99.005 1.175 ;
      RECT 98.98 0.845 98.99 1.198 ;
      RECT 98.975 0.852 98.98 1.21 ;
      RECT 98.97 0.856 98.975 1.218 ;
      RECT 98.915 0.884 98.97 1.26 ;
      RECT 98.895 0.92 98.915 1.26 ;
      RECT 98.88 0.935 98.895 1.26 ;
      RECT 98.825 0.967 98.88 1.26 ;
      RECT 98.815 0.997 98.825 1.26 ;
      RECT 98.425 0.612 98.61 0.85 ;
      RECT 98.41 0.614 98.62 0.845 ;
      RECT 98.295 0.56 98.555 0.82 ;
      RECT 98.29 0.597 98.555 0.774 ;
      RECT 98.285 0.607 98.555 0.771 ;
      RECT 98.28 0.647 98.62 0.765 ;
      RECT 98.275 0.68 98.62 0.755 ;
      RECT 98.285 0.622 98.635 0.693 ;
      RECT 98.582 1.72 98.595 2.25 ;
      RECT 98.496 1.72 98.595 2.249 ;
      RECT 98.496 1.72 98.6 2.248 ;
      RECT 98.41 1.72 98.6 2.246 ;
      RECT 98.405 1.72 98.6 2.243 ;
      RECT 98.405 1.72 98.61 2.241 ;
      RECT 98.4 2.012 98.61 2.238 ;
      RECT 98.4 2.022 98.615 2.235 ;
      RECT 98.4 2.09 98.62 2.231 ;
      RECT 98.39 2.095 98.62 2.23 ;
      RECT 98.39 2.187 98.625 2.227 ;
      RECT 98.375 1.72 98.635 1.98 ;
      RECT 97.605 0.71 97.65 2.245 ;
      RECT 97.805 0.71 97.835 0.925 ;
      RECT 96.18 0.45 96.3 0.66 ;
      RECT 95.84 0.4 96.1 0.66 ;
      RECT 95.84 0.445 96.135 0.65 ;
      RECT 97.845 0.726 97.85 0.78 ;
      RECT 97.84 0.719 97.845 0.913 ;
      RECT 97.835 0.713 97.84 0.92 ;
      RECT 97.79 0.71 97.805 0.933 ;
      RECT 97.785 0.71 97.79 0.955 ;
      RECT 97.78 0.71 97.785 1.003 ;
      RECT 97.775 0.71 97.78 1.023 ;
      RECT 97.765 0.71 97.775 1.13 ;
      RECT 97.76 0.71 97.765 1.193 ;
      RECT 97.755 0.71 97.76 1.25 ;
      RECT 97.75 0.71 97.755 1.258 ;
      RECT 97.735 0.71 97.75 1.365 ;
      RECT 97.725 0.71 97.735 1.5 ;
      RECT 97.715 0.71 97.725 1.61 ;
      RECT 97.705 0.71 97.715 1.667 ;
      RECT 97.7 0.71 97.705 1.707 ;
      RECT 97.695 0.71 97.7 1.743 ;
      RECT 97.685 0.71 97.695 1.783 ;
      RECT 97.68 0.71 97.685 1.825 ;
      RECT 97.66 0.71 97.68 1.89 ;
      RECT 97.665 2.035 97.67 2.215 ;
      RECT 97.66 2.017 97.665 2.223 ;
      RECT 97.655 0.71 97.66 1.953 ;
      RECT 97.655 1.997 97.66 2.23 ;
      RECT 97.65 0.71 97.655 2.24 ;
      RECT 97.595 0.71 97.605 1.01 ;
      RECT 97.6 1.257 97.605 2.245 ;
      RECT 97.595 1.322 97.6 2.245 ;
      RECT 97.59 0.711 97.595 1 ;
      RECT 97.585 1.387 97.595 2.245 ;
      RECT 97.58 0.712 97.59 0.99 ;
      RECT 97.57 1.5 97.585 2.245 ;
      RECT 97.575 0.713 97.58 0.98 ;
      RECT 97.555 0.714 97.575 0.958 ;
      RECT 97.56 1.597 97.57 2.245 ;
      RECT 97.555 1.672 97.56 2.245 ;
      RECT 97.545 0.713 97.555 0.935 ;
      RECT 97.55 1.715 97.555 2.245 ;
      RECT 97.545 1.742 97.55 2.245 ;
      RECT 97.535 0.711 97.545 0.923 ;
      RECT 97.54 1.785 97.545 2.245 ;
      RECT 97.535 1.812 97.54 2.245 ;
      RECT 97.525 0.71 97.535 0.91 ;
      RECT 97.53 1.827 97.535 2.245 ;
      RECT 97.49 1.885 97.53 2.245 ;
      RECT 97.52 0.709 97.525 0.895 ;
      RECT 97.515 0.707 97.52 0.888 ;
      RECT 97.505 0.704 97.515 0.878 ;
      RECT 97.5 0.701 97.505 0.863 ;
      RECT 97.485 0.697 97.5 0.856 ;
      RECT 97.48 1.94 97.49 2.245 ;
      RECT 97.48 0.694 97.485 0.851 ;
      RECT 97.465 0.69 97.48 0.845 ;
      RECT 97.475 1.957 97.48 2.245 ;
      RECT 97.465 2.02 97.475 2.245 ;
      RECT 97.385 0.675 97.465 0.825 ;
      RECT 97.46 2.027 97.465 2.24 ;
      RECT 97.455 2.035 97.46 2.23 ;
      RECT 97.375 0.661 97.385 0.809 ;
      RECT 97.36 0.657 97.375 0.807 ;
      RECT 97.35 0.652 97.36 0.803 ;
      RECT 97.325 0.645 97.35 0.795 ;
      RECT 97.32 0.64 97.325 0.79 ;
      RECT 97.31 0.64 97.32 0.788 ;
      RECT 97.3 0.638 97.31 0.786 ;
      RECT 97.27 0.63 97.3 0.78 ;
      RECT 97.255 0.622 97.27 0.773 ;
      RECT 97.235 0.617 97.255 0.766 ;
      RECT 97.23 0.613 97.235 0.761 ;
      RECT 97.2 0.606 97.23 0.755 ;
      RECT 97.175 0.597 97.2 0.745 ;
      RECT 97.145 0.59 97.175 0.737 ;
      RECT 97.12 0.58 97.145 0.728 ;
      RECT 97.105 0.572 97.12 0.722 ;
      RECT 97.08 0.567 97.105 0.717 ;
      RECT 97.07 0.563 97.08 0.712 ;
      RECT 97.05 0.558 97.07 0.707 ;
      RECT 97.015 0.553 97.05 0.7 ;
      RECT 96.955 0.548 97.015 0.693 ;
      RECT 96.942 0.544 96.955 0.691 ;
      RECT 96.856 0.539 96.942 0.688 ;
      RECT 96.77 0.529 96.856 0.684 ;
      RECT 96.729 0.522 96.77 0.681 ;
      RECT 96.643 0.515 96.729 0.678 ;
      RECT 96.557 0.505 96.643 0.674 ;
      RECT 96.471 0.495 96.557 0.669 ;
      RECT 96.385 0.485 96.471 0.665 ;
      RECT 96.375 0.47 96.385 0.663 ;
      RECT 96.365 0.455 96.375 0.663 ;
      RECT 96.3 0.45 96.365 0.662 ;
      RECT 96.135 0.447 96.18 0.655 ;
      RECT 97.38 1.352 97.385 1.543 ;
      RECT 97.375 1.347 97.38 1.55 ;
      RECT 97.361 1.345 97.375 1.556 ;
      RECT 97.275 1.345 97.361 1.558 ;
      RECT 97.271 1.345 97.275 1.561 ;
      RECT 97.185 1.345 97.271 1.579 ;
      RECT 97.175 1.35 97.185 1.598 ;
      RECT 97.165 1.405 97.175 1.602 ;
      RECT 97.14 1.42 97.165 1.609 ;
      RECT 97.1 1.44 97.14 1.622 ;
      RECT 97.095 1.452 97.1 1.632 ;
      RECT 97.08 1.458 97.095 1.637 ;
      RECT 97.075 1.463 97.08 1.641 ;
      RECT 97.055 1.47 97.075 1.646 ;
      RECT 96.985 1.495 97.055 1.663 ;
      RECT 96.945 1.523 96.985 1.683 ;
      RECT 96.94 1.533 96.945 1.691 ;
      RECT 96.92 1.54 96.94 1.693 ;
      RECT 96.915 1.547 96.92 1.696 ;
      RECT 96.885 1.555 96.915 1.699 ;
      RECT 96.88 1.56 96.885 1.703 ;
      RECT 96.806 1.564 96.88 1.711 ;
      RECT 96.72 1.573 96.806 1.727 ;
      RECT 96.716 1.578 96.72 1.736 ;
      RECT 96.63 1.583 96.716 1.746 ;
      RECT 96.59 1.591 96.63 1.758 ;
      RECT 96.54 1.597 96.59 1.765 ;
      RECT 96.455 1.606 96.54 1.78 ;
      RECT 96.38 1.617 96.455 1.798 ;
      RECT 96.345 1.624 96.38 1.808 ;
      RECT 96.27 1.632 96.345 1.813 ;
      RECT 96.215 1.641 96.27 1.813 ;
      RECT 96.19 1.646 96.215 1.811 ;
      RECT 96.18 1.649 96.19 1.809 ;
      RECT 96.145 1.651 96.18 1.807 ;
      RECT 96.115 1.653 96.145 1.803 ;
      RECT 96.07 1.652 96.115 1.799 ;
      RECT 96.05 1.647 96.07 1.796 ;
      RECT 96 1.632 96.05 1.793 ;
      RECT 95.99 1.617 96 1.788 ;
      RECT 95.94 1.602 95.99 1.778 ;
      RECT 95.89 1.577 95.94 1.758 ;
      RECT 95.88 1.562 95.89 1.74 ;
      RECT 95.875 1.56 95.88 1.734 ;
      RECT 95.855 1.555 95.875 1.729 ;
      RECT 95.85 1.547 95.855 1.723 ;
      RECT 95.835 1.541 95.85 1.716 ;
      RECT 95.83 1.536 95.835 1.708 ;
      RECT 95.81 1.531 95.83 1.7 ;
      RECT 95.795 1.524 95.81 1.693 ;
      RECT 95.78 1.518 95.795 1.684 ;
      RECT 95.775 1.512 95.78 1.677 ;
      RECT 95.73 1.487 95.775 1.663 ;
      RECT 95.715 1.457 95.73 1.645 ;
      RECT 95.7 1.44 95.715 1.636 ;
      RECT 95.675 1.42 95.7 1.624 ;
      RECT 95.635 1.39 95.675 1.604 ;
      RECT 95.625 1.36 95.635 1.589 ;
      RECT 95.61 1.35 95.625 1.582 ;
      RECT 95.555 1.315 95.61 1.561 ;
      RECT 95.54 1.278 95.555 1.54 ;
      RECT 95.53 1.265 95.54 1.532 ;
      RECT 95.48 1.235 95.53 1.514 ;
      RECT 95.465 1.165 95.48 1.495 ;
      RECT 95.42 1.165 95.465 1.478 ;
      RECT 95.395 1.165 95.42 1.46 ;
      RECT 95.385 1.165 95.395 1.453 ;
      RECT 95.306 1.165 95.385 1.446 ;
      RECT 95.22 1.165 95.306 1.438 ;
      RECT 95.205 1.197 95.22 1.433 ;
      RECT 95.13 1.207 95.205 1.429 ;
      RECT 95.11 1.217 95.13 1.424 ;
      RECT 95.085 1.217 95.11 1.421 ;
      RECT 95.075 1.207 95.085 1.42 ;
      RECT 95.065 1.18 95.075 1.419 ;
      RECT 95.025 1.175 95.065 1.417 ;
      RECT 94.98 1.175 95.025 1.413 ;
      RECT 94.955 1.175 94.98 1.408 ;
      RECT 94.905 1.175 94.955 1.395 ;
      RECT 94.865 1.18 94.875 1.38 ;
      RECT 94.875 1.175 94.905 1.385 ;
      RECT 96.86 0.955 97.12 1.215 ;
      RECT 96.855 0.977 97.12 1.173 ;
      RECT 96.095 0.805 96.315 1.17 ;
      RECT 96.077 0.892 96.315 1.169 ;
      RECT 96.06 0.897 96.315 1.166 ;
      RECT 96.06 0.897 96.335 1.165 ;
      RECT 96.03 0.907 96.335 1.163 ;
      RECT 96.025 0.922 96.335 1.159 ;
      RECT 96.025 0.922 96.34 1.158 ;
      RECT 96.02 0.98 96.34 1.156 ;
      RECT 96.02 0.98 96.35 1.153 ;
      RECT 96.015 1.045 96.35 1.148 ;
      RECT 96.095 0.805 96.355 1.065 ;
      RECT 94.84 0.635 95.1 0.895 ;
      RECT 94.84 0.678 95.186 0.869 ;
      RECT 94.84 0.678 95.23 0.868 ;
      RECT 94.84 0.678 95.25 0.866 ;
      RECT 94.84 0.678 95.35 0.865 ;
      RECT 94.84 0.678 95.37 0.863 ;
      RECT 94.84 0.678 95.38 0.858 ;
      RECT 95.25 0.645 95.44 0.855 ;
      RECT 95.25 0.647 95.445 0.853 ;
      RECT 95.24 0.652 95.45 0.845 ;
      RECT 95.186 0.676 95.45 0.845 ;
      RECT 95.23 0.67 95.24 0.867 ;
      RECT 95.24 0.65 95.445 0.853 ;
      RECT 94.195 1.71 94.4 1.94 ;
      RECT 94.135 1.66 94.19 1.92 ;
      RECT 94.195 1.66 94.395 1.94 ;
      RECT 95.165 1.975 95.17 2.002 ;
      RECT 95.155 1.885 95.165 2.007 ;
      RECT 95.15 1.807 95.155 2.013 ;
      RECT 95.14 1.797 95.15 2.02 ;
      RECT 95.135 1.787 95.14 2.026 ;
      RECT 95.125 1.782 95.135 2.028 ;
      RECT 95.11 1.774 95.125 2.036 ;
      RECT 95.095 1.765 95.11 2.048 ;
      RECT 95.085 1.757 95.095 2.058 ;
      RECT 95.05 1.675 95.085 2.076 ;
      RECT 95.015 1.675 95.05 2.095 ;
      RECT 95 1.675 95.015 2.103 ;
      RECT 94.945 1.675 95 2.103 ;
      RECT 94.911 1.675 94.945 2.094 ;
      RECT 94.825 1.675 94.911 2.07 ;
      RECT 94.815 1.735 94.825 2.052 ;
      RECT 94.775 1.737 94.815 2.043 ;
      RECT 94.77 1.739 94.775 2.033 ;
      RECT 94.75 1.741 94.77 2.028 ;
      RECT 94.74 1.744 94.75 2.023 ;
      RECT 94.73 1.745 94.74 2.018 ;
      RECT 94.706 1.746 94.73 2.01 ;
      RECT 94.62 1.751 94.706 1.988 ;
      RECT 94.565 1.75 94.62 1.961 ;
      RECT 94.55 1.743 94.565 1.948 ;
      RECT 94.515 1.738 94.55 1.944 ;
      RECT 94.46 1.73 94.515 1.943 ;
      RECT 94.4 1.717 94.46 1.941 ;
      RECT 94.19 1.66 94.195 1.928 ;
      RECT 94.265 1.03 94.45 1.24 ;
      RECT 94.255 1.035 94.465 1.233 ;
      RECT 94.295 0.94 94.555 1.2 ;
      RECT 94.25 1.097 94.555 1.123 ;
      RECT 93.595 0.89 93.6 1.69 ;
      RECT 93.54 0.94 93.57 1.69 ;
      RECT 93.53 0.94 93.535 1.25 ;
      RECT 93.515 0.94 93.52 1.245 ;
      RECT 93.06 0.985 93.075 1.2 ;
      RECT 92.99 0.985 93.075 1.195 ;
      RECT 94.255 0.565 94.325 0.775 ;
      RECT 94.325 0.572 94.335 0.77 ;
      RECT 94.221 0.565 94.255 0.782 ;
      RECT 94.135 0.565 94.221 0.806 ;
      RECT 94.125 0.57 94.135 0.825 ;
      RECT 94.12 0.582 94.125 0.828 ;
      RECT 94.105 0.597 94.12 0.832 ;
      RECT 94.1 0.615 94.105 0.836 ;
      RECT 94.06 0.625 94.1 0.845 ;
      RECT 94.045 0.632 94.06 0.857 ;
      RECT 94.03 0.637 94.045 0.862 ;
      RECT 94.015 0.64 94.03 0.867 ;
      RECT 94.005 0.642 94.015 0.871 ;
      RECT 93.97 0.649 94.005 0.879 ;
      RECT 93.935 0.657 93.97 0.893 ;
      RECT 93.925 0.663 93.935 0.902 ;
      RECT 93.92 0.665 93.925 0.904 ;
      RECT 93.9 0.668 93.92 0.91 ;
      RECT 93.87 0.675 93.9 0.921 ;
      RECT 93.86 0.681 93.87 0.928 ;
      RECT 93.835 0.684 93.86 0.935 ;
      RECT 93.825 0.688 93.835 0.943 ;
      RECT 93.82 0.689 93.825 0.965 ;
      RECT 93.815 0.69 93.82 0.98 ;
      RECT 93.81 0.691 93.815 0.995 ;
      RECT 93.805 0.692 93.81 1.01 ;
      RECT 93.8 0.693 93.805 1.04 ;
      RECT 93.79 0.695 93.8 1.073 ;
      RECT 93.775 0.699 93.79 1.12 ;
      RECT 93.765 0.702 93.775 1.165 ;
      RECT 93.76 0.705 93.765 1.193 ;
      RECT 93.75 0.707 93.76 1.22 ;
      RECT 93.745 0.71 93.75 1.255 ;
      RECT 93.715 0.715 93.745 1.313 ;
      RECT 93.71 0.72 93.715 1.398 ;
      RECT 93.705 0.722 93.71 1.433 ;
      RECT 93.7 0.724 93.705 1.515 ;
      RECT 93.695 0.726 93.7 1.603 ;
      RECT 93.685 0.728 93.695 1.685 ;
      RECT 93.67 0.742 93.685 1.69 ;
      RECT 93.635 0.787 93.67 1.69 ;
      RECT 93.625 0.827 93.635 1.69 ;
      RECT 93.61 0.855 93.625 1.69 ;
      RECT 93.605 0.872 93.61 1.69 ;
      RECT 93.6 0.88 93.605 1.69 ;
      RECT 93.59 0.895 93.595 1.69 ;
      RECT 93.585 0.902 93.59 1.69 ;
      RECT 93.575 0.922 93.585 1.69 ;
      RECT 93.57 0.935 93.575 1.69 ;
      RECT 93.535 0.94 93.54 1.275 ;
      RECT 93.52 1.33 93.54 1.69 ;
      RECT 93.52 0.94 93.53 1.248 ;
      RECT 93.515 1.37 93.52 1.69 ;
      RECT 93.465 0.94 93.515 1.243 ;
      RECT 93.51 1.407 93.515 1.69 ;
      RECT 93.5 1.43 93.51 1.69 ;
      RECT 93.495 1.475 93.5 1.69 ;
      RECT 93.485 1.485 93.495 1.683 ;
      RECT 93.411 0.94 93.465 1.237 ;
      RECT 93.325 0.94 93.411 1.23 ;
      RECT 93.276 0.987 93.325 1.223 ;
      RECT 93.19 0.995 93.276 1.216 ;
      RECT 93.175 0.992 93.19 1.211 ;
      RECT 93.161 0.985 93.175 1.21 ;
      RECT 93.075 0.985 93.161 1.205 ;
      RECT 92.98 0.99 92.99 1.19 ;
      RECT 92.57 0.42 92.585 0.82 ;
      RECT 92.765 0.42 92.77 0.68 ;
      RECT 92.51 0.42 92.555 0.68 ;
      RECT 92.965 1.725 92.97 1.93 ;
      RECT 92.96 1.715 92.965 1.935 ;
      RECT 92.955 1.702 92.96 1.94 ;
      RECT 92.95 1.682 92.955 1.94 ;
      RECT 92.925 1.635 92.95 1.94 ;
      RECT 92.89 1.55 92.925 1.94 ;
      RECT 92.885 1.487 92.89 1.94 ;
      RECT 92.88 1.472 92.885 1.94 ;
      RECT 92.865 1.432 92.88 1.94 ;
      RECT 92.86 1.407 92.865 1.94 ;
      RECT 92.85 1.39 92.86 1.94 ;
      RECT 92.815 1.312 92.85 1.94 ;
      RECT 92.81 1.255 92.815 1.94 ;
      RECT 92.805 1.242 92.81 1.94 ;
      RECT 92.795 1.22 92.805 1.94 ;
      RECT 92.785 1.185 92.795 1.94 ;
      RECT 92.775 1.155 92.785 1.94 ;
      RECT 92.765 1.07 92.775 1.583 ;
      RECT 92.772 1.715 92.775 1.94 ;
      RECT 92.77 1.725 92.772 1.94 ;
      RECT 92.76 1.735 92.77 1.935 ;
      RECT 92.755 0.42 92.765 0.815 ;
      RECT 92.76 0.947 92.765 1.558 ;
      RECT 92.755 0.845 92.76 1.541 ;
      RECT 92.745 0.42 92.755 1.517 ;
      RECT 92.74 0.42 92.745 1.488 ;
      RECT 92.735 0.42 92.74 1.478 ;
      RECT 92.715 0.42 92.735 1.44 ;
      RECT 92.71 0.42 92.715 1.398 ;
      RECT 92.705 0.42 92.71 1.378 ;
      RECT 92.675 0.42 92.705 1.328 ;
      RECT 92.665 0.42 92.675 1.275 ;
      RECT 92.66 0.42 92.665 1.248 ;
      RECT 92.655 0.42 92.66 1.233 ;
      RECT 92.645 0.42 92.655 1.21 ;
      RECT 92.635 0.42 92.645 1.185 ;
      RECT 92.63 0.42 92.635 1.125 ;
      RECT 92.62 0.42 92.63 1.063 ;
      RECT 92.615 0.42 92.62 0.983 ;
      RECT 92.61 0.42 92.615 0.948 ;
      RECT 92.605 0.42 92.61 0.923 ;
      RECT 92.6 0.42 92.605 0.908 ;
      RECT 92.595 0.42 92.6 0.878 ;
      RECT 92.59 0.42 92.595 0.855 ;
      RECT 92.585 0.42 92.59 0.828 ;
      RECT 92.555 0.42 92.57 0.815 ;
      RECT 91.71 1.955 91.895 2.165 ;
      RECT 91.7 1.96 91.91 2.158 ;
      RECT 91.7 1.96 91.93 2.13 ;
      RECT 91.7 1.96 91.945 2.109 ;
      RECT 91.7 1.96 91.96 2.107 ;
      RECT 91.7 1.96 91.97 2.106 ;
      RECT 91.7 1.96 92 2.103 ;
      RECT 92.35 1.805 92.61 2.065 ;
      RECT 92.31 1.852 92.61 2.048 ;
      RECT 92.301 1.86 92.31 2.051 ;
      RECT 91.895 1.953 92.61 2.048 ;
      RECT 92.215 1.878 92.301 2.058 ;
      RECT 91.91 1.95 92.61 2.048 ;
      RECT 92.156 1.9 92.215 2.07 ;
      RECT 91.93 1.946 92.61 2.048 ;
      RECT 92.07 1.912 92.156 2.081 ;
      RECT 91.945 1.942 92.61 2.048 ;
      RECT 92.015 1.925 92.07 2.093 ;
      RECT 91.96 1.94 92.61 2.048 ;
      RECT 92 1.931 92.015 2.099 ;
      RECT 91.97 1.936 92.61 2.048 ;
      RECT 92.115 1.46 92.375 1.72 ;
      RECT 92.115 1.48 92.485 1.69 ;
      RECT 92.115 1.485 92.495 1.685 ;
      RECT 92.306 0.899 92.385 1.13 ;
      RECT 92.22 0.902 92.435 1.125 ;
      RECT 92.215 0.902 92.435 1.12 ;
      RECT 92.215 0.907 92.445 1.118 ;
      RECT 92.19 0.907 92.445 1.115 ;
      RECT 92.19 0.915 92.455 1.113 ;
      RECT 92.07 0.85 92.33 1.11 ;
      RECT 92.07 0.897 92.38 1.11 ;
      RECT 91.325 1.47 91.33 1.73 ;
      RECT 91.155 1.24 91.16 1.73 ;
      RECT 91.04 1.48 91.045 1.705 ;
      RECT 91.75 0.575 91.755 0.785 ;
      RECT 91.755 0.58 91.77 0.78 ;
      RECT 91.69 0.575 91.75 0.793 ;
      RECT 91.675 0.575 91.69 0.803 ;
      RECT 91.625 0.575 91.675 0.82 ;
      RECT 91.605 0.575 91.625 0.843 ;
      RECT 91.59 0.575 91.605 0.855 ;
      RECT 91.57 0.575 91.59 0.865 ;
      RECT 91.56 0.58 91.57 0.874 ;
      RECT 91.555 0.59 91.56 0.879 ;
      RECT 91.55 0.602 91.555 0.883 ;
      RECT 91.54 0.625 91.55 0.888 ;
      RECT 91.535 0.64 91.54 0.892 ;
      RECT 91.53 0.657 91.535 0.895 ;
      RECT 91.525 0.665 91.53 0.898 ;
      RECT 91.515 0.67 91.525 0.902 ;
      RECT 91.51 0.677 91.515 0.907 ;
      RECT 91.5 0.682 91.51 0.911 ;
      RECT 91.475 0.694 91.5 0.922 ;
      RECT 91.455 0.711 91.475 0.938 ;
      RECT 91.43 0.728 91.455 0.96 ;
      RECT 91.395 0.751 91.43 1.018 ;
      RECT 91.375 0.773 91.395 1.08 ;
      RECT 91.37 0.783 91.375 1.115 ;
      RECT 91.36 0.79 91.37 1.153 ;
      RECT 91.355 0.797 91.36 1.173 ;
      RECT 91.35 0.808 91.355 1.21 ;
      RECT 91.345 0.816 91.35 1.275 ;
      RECT 91.335 0.827 91.345 1.328 ;
      RECT 91.33 0.845 91.335 1.398 ;
      RECT 91.325 0.855 91.33 1.435 ;
      RECT 91.32 0.865 91.325 1.73 ;
      RECT 91.315 0.877 91.32 1.73 ;
      RECT 91.31 0.887 91.315 1.73 ;
      RECT 91.3 0.897 91.31 1.73 ;
      RECT 91.29 0.92 91.3 1.73 ;
      RECT 91.275 0.955 91.29 1.73 ;
      RECT 91.235 1.017 91.275 1.73 ;
      RECT 91.23 1.07 91.235 1.73 ;
      RECT 91.205 1.105 91.23 1.73 ;
      RECT 91.19 1.15 91.205 1.73 ;
      RECT 91.185 1.172 91.19 1.73 ;
      RECT 91.175 1.185 91.185 1.73 ;
      RECT 91.165 1.21 91.175 1.73 ;
      RECT 91.16 1.232 91.165 1.73 ;
      RECT 91.135 1.27 91.155 1.73 ;
      RECT 91.095 1.327 91.135 1.73 ;
      RECT 91.09 1.377 91.095 1.73 ;
      RECT 91.085 1.395 91.09 1.73 ;
      RECT 91.08 1.407 91.085 1.73 ;
      RECT 91.07 1.425 91.08 1.73 ;
      RECT 91.06 1.445 91.07 1.705 ;
      RECT 91.055 1.462 91.06 1.705 ;
      RECT 91.045 1.475 91.055 1.705 ;
      RECT 91.015 1.485 91.04 1.705 ;
      RECT 91.005 1.492 91.015 1.705 ;
      RECT 90.99 1.502 91.005 1.7 ;
      RECT 89.95 1.415 90.27 1.675 ;
      RECT 89.815 1.46 90.27 1.63 ;
      RECT 83.49 1.515 83.865 1.765 ;
      RECT 83.59 0.73 83.765 1.765 ;
      RECT 83.59 0.73 89.515 0.905 ;
      RECT 89.095 0.475 89.415 0.905 ;
      RECT 89.095 0.505 89.495 0.675 ;
      RECT 86.76 1.515 87.055 1.805 ;
      RECT 86.73 1.515 87.055 1.775 ;
      RECT 72.97 1.885 73.275 2.115 ;
      RECT 81.11 1.915 84.525 2.09 ;
      RECT 84.35 1.065 84.525 2.09 ;
      RECT 72.97 1.915 84.525 2.085 ;
      RECT 84.295 1.065 84.625 1.315 ;
      RECT 81.555 1.075 81.845 1.315 ;
      RECT 77.105 1.045 77.365 1.28 ;
      RECT 77.105 1.075 81.845 1.245 ;
      RECT 80.29 1.415 80.61 1.675 ;
      RECT 80.275 1.46 80.61 1.63 ;
      RECT 78.995 0.395 79.29 0.685 ;
      RECT 78.96 0.395 79.29 0.655 ;
      RECT 76.155 1.415 76.475 1.675 ;
      RECT 76.14 1.46 76.475 1.63 ;
      RECT 74.48 1.205 74.8 1.465 ;
      RECT 74.465 1.205 74.82 1.44 ;
      RECT 71.78 0.965 71.965 1.175 ;
      RECT 71.77 0.97 71.98 1.168 ;
      RECT 71.77 0.97 72.066 1.145 ;
      RECT 71.77 0.97 72.125 1.12 ;
      RECT 71.77 0.97 72.18 1.1 ;
      RECT 71.77 0.97 72.19 1.088 ;
      RECT 71.77 0.97 72.385 1.027 ;
      RECT 71.77 0.97 72.415 1.01 ;
      RECT 71.77 0.97 72.435 1 ;
      RECT 72.315 0.735 72.575 0.995 ;
      RECT 72.3 0.825 72.315 1.042 ;
      RECT 71.835 0.957 72.575 0.995 ;
      RECT 72.286 0.836 72.3 1.048 ;
      RECT 71.875 0.95 72.575 0.995 ;
      RECT 72.2 0.876 72.286 1.067 ;
      RECT 72.125 0.937 72.575 0.995 ;
      RECT 72.195 0.912 72.2 1.084 ;
      RECT 72.18 0.922 72.575 0.995 ;
      RECT 72.19 0.917 72.195 1.086 ;
      RECT 72.485 1.422 72.49 1.514 ;
      RECT 72.48 1.4 72.485 1.531 ;
      RECT 72.475 1.39 72.48 1.543 ;
      RECT 72.465 1.381 72.475 1.553 ;
      RECT 72.46 1.376 72.465 1.561 ;
      RECT 72.455 1.372 72.46 1.564 ;
      RECT 72.421 1.305 72.455 1.575 ;
      RECT 72.335 1.305 72.421 1.61 ;
      RECT 72.255 1.305 72.335 1.658 ;
      RECT 72.195 1.305 72.255 1.683 ;
      RECT 72.135 1.405 72.195 1.69 ;
      RECT 72.1 1.43 72.135 1.696 ;
      RECT 72.075 1.445 72.1 1.7 ;
      RECT 72.061 1.454 72.075 1.702 ;
      RECT 71.975 1.481 72.061 1.708 ;
      RECT 71.91 1.522 71.975 1.717 ;
      RECT 71.895 1.542 71.91 1.722 ;
      RECT 71.865 1.552 71.895 1.725 ;
      RECT 71.86 1.562 71.865 1.728 ;
      RECT 71.83 1.567 71.86 1.73 ;
      RECT 71.81 1.572 71.83 1.734 ;
      RECT 71.725 1.575 71.81 1.741 ;
      RECT 71.71 1.572 71.725 1.747 ;
      RECT 71.7 1.569 71.71 1.749 ;
      RECT 71.68 1.566 71.7 1.751 ;
      RECT 71.66 1.562 71.68 1.752 ;
      RECT 71.645 1.558 71.66 1.754 ;
      RECT 71.635 1.555 71.645 1.755 ;
      RECT 71.595 1.549 71.635 1.753 ;
      RECT 71.585 1.544 71.595 1.751 ;
      RECT 71.57 1.541 71.585 1.747 ;
      RECT 71.545 1.536 71.57 1.74 ;
      RECT 71.495 1.527 71.545 1.728 ;
      RECT 71.425 1.513 71.495 1.71 ;
      RECT 71.367 1.498 71.425 1.692 ;
      RECT 71.281 1.481 71.367 1.672 ;
      RECT 71.195 1.46 71.281 1.647 ;
      RECT 71.145 1.445 71.195 1.628 ;
      RECT 71.141 1.439 71.145 1.62 ;
      RECT 71.055 1.429 71.141 1.607 ;
      RECT 71.02 1.414 71.055 1.59 ;
      RECT 71.005 1.407 71.02 1.583 ;
      RECT 70.945 1.395 71.005 1.571 ;
      RECT 70.925 1.382 70.945 1.559 ;
      RECT 70.885 1.373 70.925 1.551 ;
      RECT 70.88 1.365 70.885 1.544 ;
      RECT 70.8 1.355 70.88 1.53 ;
      RECT 70.785 1.342 70.8 1.515 ;
      RECT 70.78 1.34 70.785 1.513 ;
      RECT 70.701 1.328 70.78 1.5 ;
      RECT 70.615 1.303 70.701 1.475 ;
      RECT 70.6 1.272 70.615 1.46 ;
      RECT 70.585 1.247 70.6 1.456 ;
      RECT 70.57 1.24 70.585 1.452 ;
      RECT 70.395 1.245 70.4 1.448 ;
      RECT 70.39 1.25 70.395 1.443 ;
      RECT 70.4 1.24 70.57 1.45 ;
      RECT 71.115 1 71.22 1.26 ;
      RECT 71.93 0.525 71.935 0.75 ;
      RECT 72.06 0.525 72.115 0.735 ;
      RECT 72.115 0.53 72.125 0.728 ;
      RECT 72.021 0.525 72.06 0.738 ;
      RECT 71.935 0.525 72.021 0.745 ;
      RECT 71.915 0.53 71.93 0.751 ;
      RECT 71.905 0.57 71.915 0.753 ;
      RECT 71.875 0.58 71.905 0.755 ;
      RECT 71.87 0.585 71.875 0.757 ;
      RECT 71.845 0.59 71.87 0.759 ;
      RECT 71.83 0.595 71.845 0.761 ;
      RECT 71.815 0.597 71.83 0.763 ;
      RECT 71.81 0.602 71.815 0.765 ;
      RECT 71.76 0.61 71.81 0.768 ;
      RECT 71.735 0.619 71.76 0.773 ;
      RECT 71.725 0.626 71.735 0.778 ;
      RECT 71.72 0.629 71.725 0.782 ;
      RECT 71.7 0.632 71.72 0.791 ;
      RECT 71.67 0.64 71.7 0.811 ;
      RECT 71.641 0.653 71.67 0.833 ;
      RECT 71.555 0.687 71.641 0.877 ;
      RECT 71.55 0.713 71.555 0.915 ;
      RECT 71.545 0.717 71.55 0.924 ;
      RECT 71.51 0.73 71.545 0.957 ;
      RECT 71.5 0.744 71.51 0.995 ;
      RECT 71.495 0.748 71.5 1.008 ;
      RECT 71.49 0.752 71.495 1.013 ;
      RECT 71.48 0.76 71.49 1.025 ;
      RECT 71.475 0.767 71.48 1.04 ;
      RECT 71.45 0.78 71.475 1.065 ;
      RECT 71.41 0.809 71.45 1.12 ;
      RECT 71.395 0.834 71.41 1.175 ;
      RECT 71.385 0.845 71.395 1.198 ;
      RECT 71.38 0.852 71.385 1.21 ;
      RECT 71.375 0.856 71.38 1.218 ;
      RECT 71.32 0.884 71.375 1.26 ;
      RECT 71.3 0.92 71.32 1.26 ;
      RECT 71.285 0.935 71.3 1.26 ;
      RECT 71.23 0.967 71.285 1.26 ;
      RECT 71.22 0.997 71.23 1.26 ;
      RECT 70.83 0.612 71.015 0.85 ;
      RECT 70.815 0.614 71.025 0.845 ;
      RECT 70.7 0.56 70.96 0.82 ;
      RECT 70.695 0.597 70.96 0.774 ;
      RECT 70.69 0.607 70.96 0.771 ;
      RECT 70.685 0.647 71.025 0.765 ;
      RECT 70.68 0.68 71.025 0.755 ;
      RECT 70.69 0.622 71.04 0.693 ;
      RECT 70.987 1.72 71 2.25 ;
      RECT 70.901 1.72 71 2.249 ;
      RECT 70.901 1.72 71.005 2.248 ;
      RECT 70.815 1.72 71.005 2.246 ;
      RECT 70.81 1.72 71.005 2.243 ;
      RECT 70.81 1.72 71.015 2.241 ;
      RECT 70.805 2.012 71.015 2.238 ;
      RECT 70.805 2.022 71.02 2.235 ;
      RECT 70.805 2.09 71.025 2.231 ;
      RECT 70.795 2.095 71.025 2.23 ;
      RECT 70.795 2.187 71.03 2.227 ;
      RECT 70.78 1.72 71.04 1.98 ;
      RECT 70.01 0.71 70.055 2.245 ;
      RECT 70.21 0.71 70.24 0.925 ;
      RECT 68.585 0.45 68.705 0.66 ;
      RECT 68.245 0.4 68.505 0.66 ;
      RECT 68.245 0.445 68.54 0.65 ;
      RECT 70.25 0.726 70.255 0.78 ;
      RECT 70.245 0.719 70.25 0.913 ;
      RECT 70.24 0.713 70.245 0.92 ;
      RECT 70.195 0.71 70.21 0.933 ;
      RECT 70.19 0.71 70.195 0.955 ;
      RECT 70.185 0.71 70.19 1.003 ;
      RECT 70.18 0.71 70.185 1.023 ;
      RECT 70.17 0.71 70.18 1.13 ;
      RECT 70.165 0.71 70.17 1.193 ;
      RECT 70.16 0.71 70.165 1.25 ;
      RECT 70.155 0.71 70.16 1.258 ;
      RECT 70.14 0.71 70.155 1.365 ;
      RECT 70.13 0.71 70.14 1.5 ;
      RECT 70.12 0.71 70.13 1.61 ;
      RECT 70.11 0.71 70.12 1.667 ;
      RECT 70.105 0.71 70.11 1.707 ;
      RECT 70.1 0.71 70.105 1.743 ;
      RECT 70.09 0.71 70.1 1.783 ;
      RECT 70.085 0.71 70.09 1.825 ;
      RECT 70.065 0.71 70.085 1.89 ;
      RECT 70.07 2.035 70.075 2.215 ;
      RECT 70.065 2.017 70.07 2.223 ;
      RECT 70.06 0.71 70.065 1.953 ;
      RECT 70.06 1.997 70.065 2.23 ;
      RECT 70.055 0.71 70.06 2.24 ;
      RECT 70 0.71 70.01 1.01 ;
      RECT 70.005 1.257 70.01 2.245 ;
      RECT 70 1.322 70.005 2.245 ;
      RECT 69.995 0.711 70 1 ;
      RECT 69.99 1.387 70 2.245 ;
      RECT 69.985 0.712 69.995 0.99 ;
      RECT 69.975 1.5 69.99 2.245 ;
      RECT 69.98 0.713 69.985 0.98 ;
      RECT 69.96 0.714 69.98 0.958 ;
      RECT 69.965 1.597 69.975 2.245 ;
      RECT 69.96 1.672 69.965 2.245 ;
      RECT 69.95 0.713 69.96 0.935 ;
      RECT 69.955 1.715 69.96 2.245 ;
      RECT 69.95 1.742 69.955 2.245 ;
      RECT 69.94 0.711 69.95 0.923 ;
      RECT 69.945 1.785 69.95 2.245 ;
      RECT 69.94 1.812 69.945 2.245 ;
      RECT 69.93 0.71 69.94 0.91 ;
      RECT 69.935 1.827 69.94 2.245 ;
      RECT 69.895 1.885 69.935 2.245 ;
      RECT 69.925 0.709 69.93 0.895 ;
      RECT 69.92 0.707 69.925 0.888 ;
      RECT 69.91 0.704 69.92 0.878 ;
      RECT 69.905 0.701 69.91 0.863 ;
      RECT 69.89 0.697 69.905 0.856 ;
      RECT 69.885 1.94 69.895 2.245 ;
      RECT 69.885 0.694 69.89 0.851 ;
      RECT 69.87 0.69 69.885 0.845 ;
      RECT 69.88 1.957 69.885 2.245 ;
      RECT 69.87 2.02 69.88 2.245 ;
      RECT 69.79 0.675 69.87 0.825 ;
      RECT 69.865 2.027 69.87 2.24 ;
      RECT 69.86 2.035 69.865 2.23 ;
      RECT 69.78 0.661 69.79 0.809 ;
      RECT 69.765 0.657 69.78 0.807 ;
      RECT 69.755 0.652 69.765 0.803 ;
      RECT 69.73 0.645 69.755 0.795 ;
      RECT 69.725 0.64 69.73 0.79 ;
      RECT 69.715 0.64 69.725 0.788 ;
      RECT 69.705 0.638 69.715 0.786 ;
      RECT 69.675 0.63 69.705 0.78 ;
      RECT 69.66 0.622 69.675 0.773 ;
      RECT 69.64 0.617 69.66 0.766 ;
      RECT 69.635 0.613 69.64 0.761 ;
      RECT 69.605 0.606 69.635 0.755 ;
      RECT 69.58 0.597 69.605 0.745 ;
      RECT 69.55 0.59 69.58 0.737 ;
      RECT 69.525 0.58 69.55 0.728 ;
      RECT 69.51 0.572 69.525 0.722 ;
      RECT 69.485 0.567 69.51 0.717 ;
      RECT 69.475 0.563 69.485 0.712 ;
      RECT 69.455 0.558 69.475 0.707 ;
      RECT 69.42 0.553 69.455 0.7 ;
      RECT 69.36 0.548 69.42 0.693 ;
      RECT 69.347 0.544 69.36 0.691 ;
      RECT 69.261 0.539 69.347 0.688 ;
      RECT 69.175 0.529 69.261 0.684 ;
      RECT 69.134 0.522 69.175 0.681 ;
      RECT 69.048 0.515 69.134 0.678 ;
      RECT 68.962 0.505 69.048 0.674 ;
      RECT 68.876 0.495 68.962 0.669 ;
      RECT 68.79 0.485 68.876 0.665 ;
      RECT 68.78 0.47 68.79 0.663 ;
      RECT 68.77 0.455 68.78 0.663 ;
      RECT 68.705 0.45 68.77 0.662 ;
      RECT 68.54 0.447 68.585 0.655 ;
      RECT 69.785 1.352 69.79 1.543 ;
      RECT 69.78 1.347 69.785 1.55 ;
      RECT 69.766 1.345 69.78 1.556 ;
      RECT 69.68 1.345 69.766 1.558 ;
      RECT 69.676 1.345 69.68 1.561 ;
      RECT 69.59 1.345 69.676 1.579 ;
      RECT 69.58 1.35 69.59 1.598 ;
      RECT 69.57 1.405 69.58 1.602 ;
      RECT 69.545 1.42 69.57 1.609 ;
      RECT 69.505 1.44 69.545 1.622 ;
      RECT 69.5 1.452 69.505 1.632 ;
      RECT 69.485 1.458 69.5 1.637 ;
      RECT 69.48 1.463 69.485 1.641 ;
      RECT 69.46 1.47 69.48 1.646 ;
      RECT 69.39 1.495 69.46 1.663 ;
      RECT 69.35 1.523 69.39 1.683 ;
      RECT 69.345 1.533 69.35 1.691 ;
      RECT 69.325 1.54 69.345 1.693 ;
      RECT 69.32 1.547 69.325 1.696 ;
      RECT 69.29 1.555 69.32 1.699 ;
      RECT 69.285 1.56 69.29 1.703 ;
      RECT 69.211 1.564 69.285 1.711 ;
      RECT 69.125 1.573 69.211 1.727 ;
      RECT 69.121 1.578 69.125 1.736 ;
      RECT 69.035 1.583 69.121 1.746 ;
      RECT 68.995 1.591 69.035 1.758 ;
      RECT 68.945 1.597 68.995 1.765 ;
      RECT 68.86 1.606 68.945 1.78 ;
      RECT 68.785 1.617 68.86 1.798 ;
      RECT 68.75 1.624 68.785 1.808 ;
      RECT 68.675 1.632 68.75 1.813 ;
      RECT 68.62 1.641 68.675 1.813 ;
      RECT 68.595 1.646 68.62 1.811 ;
      RECT 68.585 1.649 68.595 1.809 ;
      RECT 68.55 1.651 68.585 1.807 ;
      RECT 68.52 1.653 68.55 1.803 ;
      RECT 68.475 1.652 68.52 1.799 ;
      RECT 68.455 1.647 68.475 1.796 ;
      RECT 68.405 1.632 68.455 1.793 ;
      RECT 68.395 1.617 68.405 1.788 ;
      RECT 68.345 1.602 68.395 1.778 ;
      RECT 68.295 1.577 68.345 1.758 ;
      RECT 68.285 1.562 68.295 1.74 ;
      RECT 68.28 1.56 68.285 1.734 ;
      RECT 68.26 1.555 68.28 1.729 ;
      RECT 68.255 1.547 68.26 1.723 ;
      RECT 68.24 1.541 68.255 1.716 ;
      RECT 68.235 1.536 68.24 1.708 ;
      RECT 68.215 1.531 68.235 1.7 ;
      RECT 68.2 1.524 68.215 1.693 ;
      RECT 68.185 1.518 68.2 1.684 ;
      RECT 68.18 1.512 68.185 1.677 ;
      RECT 68.135 1.487 68.18 1.663 ;
      RECT 68.12 1.457 68.135 1.645 ;
      RECT 68.105 1.44 68.12 1.636 ;
      RECT 68.08 1.42 68.105 1.624 ;
      RECT 68.04 1.39 68.08 1.604 ;
      RECT 68.03 1.36 68.04 1.589 ;
      RECT 68.015 1.35 68.03 1.582 ;
      RECT 67.96 1.315 68.015 1.561 ;
      RECT 67.945 1.278 67.96 1.54 ;
      RECT 67.935 1.265 67.945 1.532 ;
      RECT 67.885 1.235 67.935 1.514 ;
      RECT 67.87 1.165 67.885 1.495 ;
      RECT 67.825 1.165 67.87 1.478 ;
      RECT 67.8 1.165 67.825 1.46 ;
      RECT 67.79 1.165 67.8 1.453 ;
      RECT 67.711 1.165 67.79 1.446 ;
      RECT 67.625 1.165 67.711 1.438 ;
      RECT 67.61 1.197 67.625 1.433 ;
      RECT 67.535 1.207 67.61 1.429 ;
      RECT 67.515 1.217 67.535 1.424 ;
      RECT 67.49 1.217 67.515 1.421 ;
      RECT 67.48 1.207 67.49 1.42 ;
      RECT 67.47 1.18 67.48 1.419 ;
      RECT 67.43 1.175 67.47 1.417 ;
      RECT 67.385 1.175 67.43 1.413 ;
      RECT 67.36 1.175 67.385 1.408 ;
      RECT 67.31 1.175 67.36 1.395 ;
      RECT 67.27 1.18 67.28 1.38 ;
      RECT 67.28 1.175 67.31 1.385 ;
      RECT 69.265 0.955 69.525 1.215 ;
      RECT 69.26 0.977 69.525 1.173 ;
      RECT 68.5 0.805 68.72 1.17 ;
      RECT 68.482 0.892 68.72 1.169 ;
      RECT 68.465 0.897 68.72 1.166 ;
      RECT 68.465 0.897 68.74 1.165 ;
      RECT 68.435 0.907 68.74 1.163 ;
      RECT 68.43 0.922 68.74 1.159 ;
      RECT 68.43 0.922 68.745 1.158 ;
      RECT 68.425 0.98 68.745 1.156 ;
      RECT 68.425 0.98 68.755 1.153 ;
      RECT 68.42 1.045 68.755 1.148 ;
      RECT 68.5 0.805 68.76 1.065 ;
      RECT 67.245 0.635 67.505 0.895 ;
      RECT 67.245 0.678 67.591 0.869 ;
      RECT 67.245 0.678 67.635 0.868 ;
      RECT 67.245 0.678 67.655 0.866 ;
      RECT 67.245 0.678 67.755 0.865 ;
      RECT 67.245 0.678 67.775 0.863 ;
      RECT 67.245 0.678 67.785 0.858 ;
      RECT 67.655 0.645 67.845 0.855 ;
      RECT 67.655 0.647 67.85 0.853 ;
      RECT 67.645 0.652 67.855 0.845 ;
      RECT 67.591 0.676 67.855 0.845 ;
      RECT 67.635 0.67 67.645 0.867 ;
      RECT 67.645 0.65 67.85 0.853 ;
      RECT 66.6 1.71 66.805 1.94 ;
      RECT 66.54 1.66 66.595 1.92 ;
      RECT 66.6 1.66 66.8 1.94 ;
      RECT 67.57 1.975 67.575 2.002 ;
      RECT 67.56 1.885 67.57 2.007 ;
      RECT 67.555 1.807 67.56 2.013 ;
      RECT 67.545 1.797 67.555 2.02 ;
      RECT 67.54 1.787 67.545 2.026 ;
      RECT 67.53 1.782 67.54 2.028 ;
      RECT 67.515 1.774 67.53 2.036 ;
      RECT 67.5 1.765 67.515 2.048 ;
      RECT 67.49 1.757 67.5 2.058 ;
      RECT 67.455 1.675 67.49 2.076 ;
      RECT 67.42 1.675 67.455 2.095 ;
      RECT 67.405 1.675 67.42 2.103 ;
      RECT 67.35 1.675 67.405 2.103 ;
      RECT 67.316 1.675 67.35 2.094 ;
      RECT 67.23 1.675 67.316 2.07 ;
      RECT 67.22 1.735 67.23 2.052 ;
      RECT 67.18 1.737 67.22 2.043 ;
      RECT 67.175 1.739 67.18 2.033 ;
      RECT 67.155 1.741 67.175 2.028 ;
      RECT 67.145 1.744 67.155 2.023 ;
      RECT 67.135 1.745 67.145 2.018 ;
      RECT 67.111 1.746 67.135 2.01 ;
      RECT 67.025 1.751 67.111 1.988 ;
      RECT 66.97 1.75 67.025 1.961 ;
      RECT 66.955 1.743 66.97 1.948 ;
      RECT 66.92 1.738 66.955 1.944 ;
      RECT 66.865 1.73 66.92 1.943 ;
      RECT 66.805 1.717 66.865 1.941 ;
      RECT 66.595 1.66 66.6 1.928 ;
      RECT 66.67 1.03 66.855 1.24 ;
      RECT 66.66 1.035 66.87 1.233 ;
      RECT 66.7 0.94 66.96 1.2 ;
      RECT 66.655 1.097 66.96 1.123 ;
      RECT 66 0.89 66.005 1.69 ;
      RECT 65.945 0.94 65.975 1.69 ;
      RECT 65.935 0.94 65.94 1.25 ;
      RECT 65.92 0.94 65.925 1.245 ;
      RECT 65.465 0.985 65.48 1.2 ;
      RECT 65.395 0.985 65.48 1.195 ;
      RECT 66.66 0.565 66.73 0.775 ;
      RECT 66.73 0.572 66.74 0.77 ;
      RECT 66.626 0.565 66.66 0.782 ;
      RECT 66.54 0.565 66.626 0.806 ;
      RECT 66.53 0.57 66.54 0.825 ;
      RECT 66.525 0.582 66.53 0.828 ;
      RECT 66.51 0.597 66.525 0.832 ;
      RECT 66.505 0.615 66.51 0.836 ;
      RECT 66.465 0.625 66.505 0.845 ;
      RECT 66.45 0.632 66.465 0.857 ;
      RECT 66.435 0.637 66.45 0.862 ;
      RECT 66.42 0.64 66.435 0.867 ;
      RECT 66.41 0.642 66.42 0.871 ;
      RECT 66.375 0.649 66.41 0.879 ;
      RECT 66.34 0.657 66.375 0.893 ;
      RECT 66.33 0.663 66.34 0.902 ;
      RECT 66.325 0.665 66.33 0.904 ;
      RECT 66.305 0.668 66.325 0.91 ;
      RECT 66.275 0.675 66.305 0.921 ;
      RECT 66.265 0.681 66.275 0.928 ;
      RECT 66.24 0.684 66.265 0.935 ;
      RECT 66.23 0.688 66.24 0.943 ;
      RECT 66.225 0.689 66.23 0.965 ;
      RECT 66.22 0.69 66.225 0.98 ;
      RECT 66.215 0.691 66.22 0.995 ;
      RECT 66.21 0.692 66.215 1.01 ;
      RECT 66.205 0.693 66.21 1.04 ;
      RECT 66.195 0.695 66.205 1.073 ;
      RECT 66.18 0.699 66.195 1.12 ;
      RECT 66.17 0.702 66.18 1.165 ;
      RECT 66.165 0.705 66.17 1.193 ;
      RECT 66.155 0.707 66.165 1.22 ;
      RECT 66.15 0.71 66.155 1.255 ;
      RECT 66.12 0.715 66.15 1.313 ;
      RECT 66.115 0.72 66.12 1.398 ;
      RECT 66.11 0.722 66.115 1.433 ;
      RECT 66.105 0.724 66.11 1.515 ;
      RECT 66.1 0.726 66.105 1.603 ;
      RECT 66.09 0.728 66.1 1.685 ;
      RECT 66.075 0.742 66.09 1.69 ;
      RECT 66.04 0.787 66.075 1.69 ;
      RECT 66.03 0.827 66.04 1.69 ;
      RECT 66.015 0.855 66.03 1.69 ;
      RECT 66.01 0.872 66.015 1.69 ;
      RECT 66.005 0.88 66.01 1.69 ;
      RECT 65.995 0.895 66 1.69 ;
      RECT 65.99 0.902 65.995 1.69 ;
      RECT 65.98 0.922 65.99 1.69 ;
      RECT 65.975 0.935 65.98 1.69 ;
      RECT 65.94 0.94 65.945 1.275 ;
      RECT 65.925 1.33 65.945 1.69 ;
      RECT 65.925 0.94 65.935 1.248 ;
      RECT 65.92 1.37 65.925 1.69 ;
      RECT 65.87 0.94 65.92 1.243 ;
      RECT 65.915 1.407 65.92 1.69 ;
      RECT 65.905 1.43 65.915 1.69 ;
      RECT 65.9 1.475 65.905 1.69 ;
      RECT 65.89 1.485 65.9 1.683 ;
      RECT 65.816 0.94 65.87 1.237 ;
      RECT 65.73 0.94 65.816 1.23 ;
      RECT 65.681 0.987 65.73 1.223 ;
      RECT 65.595 0.995 65.681 1.216 ;
      RECT 65.58 0.992 65.595 1.211 ;
      RECT 65.566 0.985 65.58 1.21 ;
      RECT 65.48 0.985 65.566 1.205 ;
      RECT 65.385 0.99 65.395 1.19 ;
      RECT 64.975 0.42 64.99 0.82 ;
      RECT 65.17 0.42 65.175 0.68 ;
      RECT 64.915 0.42 64.96 0.68 ;
      RECT 65.37 1.725 65.375 1.93 ;
      RECT 65.365 1.715 65.37 1.935 ;
      RECT 65.36 1.702 65.365 1.94 ;
      RECT 65.355 1.682 65.36 1.94 ;
      RECT 65.33 1.635 65.355 1.94 ;
      RECT 65.295 1.55 65.33 1.94 ;
      RECT 65.29 1.487 65.295 1.94 ;
      RECT 65.285 1.472 65.29 1.94 ;
      RECT 65.27 1.432 65.285 1.94 ;
      RECT 65.265 1.407 65.27 1.94 ;
      RECT 65.255 1.39 65.265 1.94 ;
      RECT 65.22 1.312 65.255 1.94 ;
      RECT 65.215 1.255 65.22 1.94 ;
      RECT 65.21 1.242 65.215 1.94 ;
      RECT 65.2 1.22 65.21 1.94 ;
      RECT 65.19 1.185 65.2 1.94 ;
      RECT 65.18 1.155 65.19 1.94 ;
      RECT 65.17 1.07 65.18 1.583 ;
      RECT 65.177 1.715 65.18 1.94 ;
      RECT 65.175 1.725 65.177 1.94 ;
      RECT 65.165 1.735 65.175 1.935 ;
      RECT 65.16 0.42 65.17 0.815 ;
      RECT 65.165 0.947 65.17 1.558 ;
      RECT 65.16 0.845 65.165 1.541 ;
      RECT 65.15 0.42 65.16 1.517 ;
      RECT 65.145 0.42 65.15 1.488 ;
      RECT 65.14 0.42 65.145 1.478 ;
      RECT 65.12 0.42 65.14 1.44 ;
      RECT 65.115 0.42 65.12 1.398 ;
      RECT 65.11 0.42 65.115 1.378 ;
      RECT 65.08 0.42 65.11 1.328 ;
      RECT 65.07 0.42 65.08 1.275 ;
      RECT 65.065 0.42 65.07 1.248 ;
      RECT 65.06 0.42 65.065 1.233 ;
      RECT 65.05 0.42 65.06 1.21 ;
      RECT 65.04 0.42 65.05 1.185 ;
      RECT 65.035 0.42 65.04 1.125 ;
      RECT 65.025 0.42 65.035 1.063 ;
      RECT 65.02 0.42 65.025 0.983 ;
      RECT 65.015 0.42 65.02 0.948 ;
      RECT 65.01 0.42 65.015 0.923 ;
      RECT 65.005 0.42 65.01 0.908 ;
      RECT 65 0.42 65.005 0.878 ;
      RECT 64.995 0.42 65 0.855 ;
      RECT 64.99 0.42 64.995 0.828 ;
      RECT 64.96 0.42 64.975 0.815 ;
      RECT 64.115 1.955 64.3 2.165 ;
      RECT 64.105 1.96 64.315 2.158 ;
      RECT 64.105 1.96 64.335 2.13 ;
      RECT 64.105 1.96 64.35 2.109 ;
      RECT 64.105 1.96 64.365 2.107 ;
      RECT 64.105 1.96 64.375 2.106 ;
      RECT 64.105 1.96 64.405 2.103 ;
      RECT 64.755 1.805 65.015 2.065 ;
      RECT 64.715 1.852 65.015 2.048 ;
      RECT 64.706 1.86 64.715 2.051 ;
      RECT 64.3 1.953 65.015 2.048 ;
      RECT 64.62 1.878 64.706 2.058 ;
      RECT 64.315 1.95 65.015 2.048 ;
      RECT 64.561 1.9 64.62 2.07 ;
      RECT 64.335 1.946 65.015 2.048 ;
      RECT 64.475 1.912 64.561 2.081 ;
      RECT 64.35 1.942 65.015 2.048 ;
      RECT 64.42 1.925 64.475 2.093 ;
      RECT 64.365 1.94 65.015 2.048 ;
      RECT 64.405 1.931 64.42 2.099 ;
      RECT 64.375 1.936 65.015 2.048 ;
      RECT 64.52 1.46 64.78 1.72 ;
      RECT 64.52 1.48 64.89 1.69 ;
      RECT 64.52 1.485 64.9 1.685 ;
      RECT 64.711 0.899 64.79 1.13 ;
      RECT 64.625 0.902 64.84 1.125 ;
      RECT 64.62 0.902 64.84 1.12 ;
      RECT 64.62 0.907 64.85 1.118 ;
      RECT 64.595 0.907 64.85 1.115 ;
      RECT 64.595 0.915 64.86 1.113 ;
      RECT 64.475 0.85 64.735 1.11 ;
      RECT 64.475 0.897 64.785 1.11 ;
      RECT 63.73 1.47 63.735 1.73 ;
      RECT 63.56 1.24 63.565 1.73 ;
      RECT 63.445 1.48 63.45 1.705 ;
      RECT 64.155 0.575 64.16 0.785 ;
      RECT 64.16 0.58 64.175 0.78 ;
      RECT 64.095 0.575 64.155 0.793 ;
      RECT 64.08 0.575 64.095 0.803 ;
      RECT 64.03 0.575 64.08 0.82 ;
      RECT 64.01 0.575 64.03 0.843 ;
      RECT 63.995 0.575 64.01 0.855 ;
      RECT 63.975 0.575 63.995 0.865 ;
      RECT 63.965 0.58 63.975 0.874 ;
      RECT 63.96 0.59 63.965 0.879 ;
      RECT 63.955 0.602 63.96 0.883 ;
      RECT 63.945 0.625 63.955 0.888 ;
      RECT 63.94 0.64 63.945 0.892 ;
      RECT 63.935 0.657 63.94 0.895 ;
      RECT 63.93 0.665 63.935 0.898 ;
      RECT 63.92 0.67 63.93 0.902 ;
      RECT 63.915 0.677 63.92 0.907 ;
      RECT 63.905 0.682 63.915 0.911 ;
      RECT 63.88 0.694 63.905 0.922 ;
      RECT 63.86 0.711 63.88 0.938 ;
      RECT 63.835 0.728 63.86 0.96 ;
      RECT 63.8 0.751 63.835 1.018 ;
      RECT 63.78 0.773 63.8 1.08 ;
      RECT 63.775 0.783 63.78 1.115 ;
      RECT 63.765 0.79 63.775 1.153 ;
      RECT 63.76 0.797 63.765 1.173 ;
      RECT 63.755 0.808 63.76 1.21 ;
      RECT 63.75 0.816 63.755 1.275 ;
      RECT 63.74 0.827 63.75 1.328 ;
      RECT 63.735 0.845 63.74 1.398 ;
      RECT 63.73 0.855 63.735 1.435 ;
      RECT 63.725 0.865 63.73 1.73 ;
      RECT 63.72 0.877 63.725 1.73 ;
      RECT 63.715 0.887 63.72 1.73 ;
      RECT 63.705 0.897 63.715 1.73 ;
      RECT 63.695 0.92 63.705 1.73 ;
      RECT 63.68 0.955 63.695 1.73 ;
      RECT 63.64 1.017 63.68 1.73 ;
      RECT 63.635 1.07 63.64 1.73 ;
      RECT 63.61 1.105 63.635 1.73 ;
      RECT 63.595 1.15 63.61 1.73 ;
      RECT 63.59 1.172 63.595 1.73 ;
      RECT 63.58 1.185 63.59 1.73 ;
      RECT 63.57 1.21 63.58 1.73 ;
      RECT 63.565 1.232 63.57 1.73 ;
      RECT 63.54 1.27 63.56 1.73 ;
      RECT 63.5 1.327 63.54 1.73 ;
      RECT 63.495 1.377 63.5 1.73 ;
      RECT 63.49 1.395 63.495 1.73 ;
      RECT 63.485 1.407 63.49 1.73 ;
      RECT 63.475 1.425 63.485 1.73 ;
      RECT 63.465 1.445 63.475 1.705 ;
      RECT 63.46 1.462 63.465 1.705 ;
      RECT 63.45 1.475 63.46 1.705 ;
      RECT 63.42 1.485 63.445 1.705 ;
      RECT 63.41 1.492 63.42 1.705 ;
      RECT 63.395 1.502 63.41 1.7 ;
      RECT 62.355 1.415 62.675 1.675 ;
      RECT 62.22 1.46 62.675 1.63 ;
      RECT 55.91 1.515 56.285 1.765 ;
      RECT 56.01 0.73 56.185 1.765 ;
      RECT 56.01 0.73 61.935 0.905 ;
      RECT 61.5 0.475 61.82 0.905 ;
      RECT 61.5 0.505 61.9 0.675 ;
      RECT 59.165 1.515 59.46 1.805 ;
      RECT 59.135 1.515 59.46 1.775 ;
      RECT 45.375 1.885 45.68 2.115 ;
      RECT 53.515 1.915 56.93 2.09 ;
      RECT 56.755 1.065 56.93 2.09 ;
      RECT 45.375 1.915 56.93 2.085 ;
      RECT 56.7 1.065 57.03 1.315 ;
      RECT 53.96 1.075 54.25 1.315 ;
      RECT 49.51 1.045 49.77 1.28 ;
      RECT 49.51 1.075 54.25 1.245 ;
      RECT 52.695 1.415 53.015 1.675 ;
      RECT 52.68 1.46 53.015 1.63 ;
      RECT 51.4 0.395 51.695 0.685 ;
      RECT 51.365 0.395 51.695 0.655 ;
      RECT 48.56 1.415 48.88 1.675 ;
      RECT 48.545 1.46 48.88 1.63 ;
      RECT 46.885 1.205 47.205 1.465 ;
      RECT 46.87 1.205 47.225 1.44 ;
      RECT 44.185 0.965 44.37 1.175 ;
      RECT 44.175 0.97 44.385 1.168 ;
      RECT 44.175 0.97 44.471 1.145 ;
      RECT 44.175 0.97 44.53 1.12 ;
      RECT 44.175 0.97 44.585 1.1 ;
      RECT 44.175 0.97 44.595 1.088 ;
      RECT 44.175 0.97 44.79 1.027 ;
      RECT 44.175 0.97 44.82 1.01 ;
      RECT 44.175 0.97 44.84 1 ;
      RECT 44.72 0.735 44.98 0.995 ;
      RECT 44.705 0.825 44.72 1.042 ;
      RECT 44.24 0.957 44.98 0.995 ;
      RECT 44.691 0.836 44.705 1.048 ;
      RECT 44.28 0.95 44.98 0.995 ;
      RECT 44.605 0.876 44.691 1.067 ;
      RECT 44.53 0.937 44.98 0.995 ;
      RECT 44.6 0.912 44.605 1.084 ;
      RECT 44.585 0.922 44.98 0.995 ;
      RECT 44.595 0.917 44.6 1.086 ;
      RECT 44.89 1.422 44.895 1.514 ;
      RECT 44.885 1.4 44.89 1.531 ;
      RECT 44.88 1.39 44.885 1.543 ;
      RECT 44.87 1.381 44.88 1.553 ;
      RECT 44.865 1.376 44.87 1.561 ;
      RECT 44.86 1.372 44.865 1.564 ;
      RECT 44.826 1.305 44.86 1.575 ;
      RECT 44.74 1.305 44.826 1.61 ;
      RECT 44.66 1.305 44.74 1.658 ;
      RECT 44.6 1.305 44.66 1.683 ;
      RECT 44.54 1.405 44.6 1.69 ;
      RECT 44.505 1.43 44.54 1.696 ;
      RECT 44.48 1.445 44.505 1.7 ;
      RECT 44.466 1.454 44.48 1.702 ;
      RECT 44.38 1.481 44.466 1.708 ;
      RECT 44.315 1.522 44.38 1.717 ;
      RECT 44.3 1.542 44.315 1.722 ;
      RECT 44.27 1.552 44.3 1.725 ;
      RECT 44.265 1.562 44.27 1.728 ;
      RECT 44.235 1.567 44.265 1.73 ;
      RECT 44.215 1.572 44.235 1.734 ;
      RECT 44.13 1.575 44.215 1.741 ;
      RECT 44.115 1.572 44.13 1.747 ;
      RECT 44.105 1.569 44.115 1.749 ;
      RECT 44.085 1.566 44.105 1.751 ;
      RECT 44.065 1.562 44.085 1.752 ;
      RECT 44.05 1.558 44.065 1.754 ;
      RECT 44.04 1.555 44.05 1.755 ;
      RECT 44 1.549 44.04 1.753 ;
      RECT 43.99 1.544 44 1.751 ;
      RECT 43.975 1.541 43.99 1.747 ;
      RECT 43.95 1.536 43.975 1.74 ;
      RECT 43.9 1.527 43.95 1.728 ;
      RECT 43.83 1.513 43.9 1.71 ;
      RECT 43.772 1.498 43.83 1.692 ;
      RECT 43.686 1.481 43.772 1.672 ;
      RECT 43.6 1.46 43.686 1.647 ;
      RECT 43.55 1.445 43.6 1.628 ;
      RECT 43.546 1.439 43.55 1.62 ;
      RECT 43.46 1.429 43.546 1.607 ;
      RECT 43.425 1.414 43.46 1.59 ;
      RECT 43.41 1.407 43.425 1.583 ;
      RECT 43.35 1.395 43.41 1.571 ;
      RECT 43.33 1.382 43.35 1.559 ;
      RECT 43.29 1.373 43.33 1.551 ;
      RECT 43.285 1.365 43.29 1.544 ;
      RECT 43.205 1.355 43.285 1.53 ;
      RECT 43.19 1.342 43.205 1.515 ;
      RECT 43.185 1.34 43.19 1.513 ;
      RECT 43.106 1.328 43.185 1.5 ;
      RECT 43.02 1.303 43.106 1.475 ;
      RECT 43.005 1.272 43.02 1.46 ;
      RECT 42.99 1.247 43.005 1.456 ;
      RECT 42.975 1.24 42.99 1.452 ;
      RECT 42.8 1.245 42.805 1.448 ;
      RECT 42.795 1.25 42.8 1.443 ;
      RECT 42.805 1.24 42.975 1.45 ;
      RECT 43.52 1 43.625 1.26 ;
      RECT 44.335 0.525 44.34 0.75 ;
      RECT 44.465 0.525 44.52 0.735 ;
      RECT 44.52 0.53 44.53 0.728 ;
      RECT 44.426 0.525 44.465 0.738 ;
      RECT 44.34 0.525 44.426 0.745 ;
      RECT 44.32 0.53 44.335 0.751 ;
      RECT 44.31 0.57 44.32 0.753 ;
      RECT 44.28 0.58 44.31 0.755 ;
      RECT 44.275 0.585 44.28 0.757 ;
      RECT 44.25 0.59 44.275 0.759 ;
      RECT 44.235 0.595 44.25 0.761 ;
      RECT 44.22 0.597 44.235 0.763 ;
      RECT 44.215 0.602 44.22 0.765 ;
      RECT 44.165 0.61 44.215 0.768 ;
      RECT 44.14 0.619 44.165 0.773 ;
      RECT 44.13 0.626 44.14 0.778 ;
      RECT 44.125 0.629 44.13 0.782 ;
      RECT 44.105 0.632 44.125 0.791 ;
      RECT 44.075 0.64 44.105 0.811 ;
      RECT 44.046 0.653 44.075 0.833 ;
      RECT 43.96 0.687 44.046 0.877 ;
      RECT 43.955 0.713 43.96 0.915 ;
      RECT 43.95 0.717 43.955 0.924 ;
      RECT 43.915 0.73 43.95 0.957 ;
      RECT 43.905 0.744 43.915 0.995 ;
      RECT 43.9 0.748 43.905 1.008 ;
      RECT 43.895 0.752 43.9 1.013 ;
      RECT 43.885 0.76 43.895 1.025 ;
      RECT 43.88 0.767 43.885 1.04 ;
      RECT 43.855 0.78 43.88 1.065 ;
      RECT 43.815 0.809 43.855 1.12 ;
      RECT 43.8 0.834 43.815 1.175 ;
      RECT 43.79 0.845 43.8 1.198 ;
      RECT 43.785 0.852 43.79 1.21 ;
      RECT 43.78 0.856 43.785 1.218 ;
      RECT 43.725 0.884 43.78 1.26 ;
      RECT 43.705 0.92 43.725 1.26 ;
      RECT 43.69 0.935 43.705 1.26 ;
      RECT 43.635 0.967 43.69 1.26 ;
      RECT 43.625 0.997 43.635 1.26 ;
      RECT 43.235 0.612 43.42 0.85 ;
      RECT 43.22 0.614 43.43 0.845 ;
      RECT 43.105 0.56 43.365 0.82 ;
      RECT 43.1 0.597 43.365 0.774 ;
      RECT 43.095 0.607 43.365 0.771 ;
      RECT 43.09 0.647 43.43 0.765 ;
      RECT 43.085 0.68 43.43 0.755 ;
      RECT 43.095 0.622 43.445 0.693 ;
      RECT 43.392 1.72 43.405 2.25 ;
      RECT 43.306 1.72 43.405 2.249 ;
      RECT 43.306 1.72 43.41 2.248 ;
      RECT 43.22 1.72 43.41 2.246 ;
      RECT 43.215 1.72 43.41 2.243 ;
      RECT 43.215 1.72 43.42 2.241 ;
      RECT 43.21 2.012 43.42 2.238 ;
      RECT 43.21 2.022 43.425 2.235 ;
      RECT 43.21 2.09 43.43 2.231 ;
      RECT 43.2 2.095 43.43 2.23 ;
      RECT 43.2 2.187 43.435 2.227 ;
      RECT 43.185 1.72 43.445 1.98 ;
      RECT 42.415 0.71 42.46 2.245 ;
      RECT 42.615 0.71 42.645 0.925 ;
      RECT 40.99 0.45 41.11 0.66 ;
      RECT 40.65 0.4 40.91 0.66 ;
      RECT 40.65 0.445 40.945 0.65 ;
      RECT 42.655 0.726 42.66 0.78 ;
      RECT 42.65 0.719 42.655 0.913 ;
      RECT 42.645 0.713 42.65 0.92 ;
      RECT 42.6 0.71 42.615 0.933 ;
      RECT 42.595 0.71 42.6 0.955 ;
      RECT 42.59 0.71 42.595 1.003 ;
      RECT 42.585 0.71 42.59 1.023 ;
      RECT 42.575 0.71 42.585 1.13 ;
      RECT 42.57 0.71 42.575 1.193 ;
      RECT 42.565 0.71 42.57 1.25 ;
      RECT 42.56 0.71 42.565 1.258 ;
      RECT 42.545 0.71 42.56 1.365 ;
      RECT 42.535 0.71 42.545 1.5 ;
      RECT 42.525 0.71 42.535 1.61 ;
      RECT 42.515 0.71 42.525 1.667 ;
      RECT 42.51 0.71 42.515 1.707 ;
      RECT 42.505 0.71 42.51 1.743 ;
      RECT 42.495 0.71 42.505 1.783 ;
      RECT 42.49 0.71 42.495 1.825 ;
      RECT 42.47 0.71 42.49 1.89 ;
      RECT 42.475 2.035 42.48 2.215 ;
      RECT 42.47 2.017 42.475 2.223 ;
      RECT 42.465 0.71 42.47 1.953 ;
      RECT 42.465 1.997 42.47 2.23 ;
      RECT 42.46 0.71 42.465 2.24 ;
      RECT 42.405 0.71 42.415 1.01 ;
      RECT 42.41 1.257 42.415 2.245 ;
      RECT 42.405 1.322 42.41 2.245 ;
      RECT 42.4 0.711 42.405 1 ;
      RECT 42.395 1.387 42.405 2.245 ;
      RECT 42.39 0.712 42.4 0.99 ;
      RECT 42.38 1.5 42.395 2.245 ;
      RECT 42.385 0.713 42.39 0.98 ;
      RECT 42.365 0.714 42.385 0.958 ;
      RECT 42.37 1.597 42.38 2.245 ;
      RECT 42.365 1.672 42.37 2.245 ;
      RECT 42.355 0.713 42.365 0.935 ;
      RECT 42.36 1.715 42.365 2.245 ;
      RECT 42.355 1.742 42.36 2.245 ;
      RECT 42.345 0.711 42.355 0.923 ;
      RECT 42.35 1.785 42.355 2.245 ;
      RECT 42.345 1.812 42.35 2.245 ;
      RECT 42.335 0.71 42.345 0.91 ;
      RECT 42.34 1.827 42.345 2.245 ;
      RECT 42.3 1.885 42.34 2.245 ;
      RECT 42.33 0.709 42.335 0.895 ;
      RECT 42.325 0.707 42.33 0.888 ;
      RECT 42.315 0.704 42.325 0.878 ;
      RECT 42.31 0.701 42.315 0.863 ;
      RECT 42.295 0.697 42.31 0.856 ;
      RECT 42.29 1.94 42.3 2.245 ;
      RECT 42.29 0.694 42.295 0.851 ;
      RECT 42.275 0.69 42.29 0.845 ;
      RECT 42.285 1.957 42.29 2.245 ;
      RECT 42.275 2.02 42.285 2.245 ;
      RECT 42.195 0.675 42.275 0.825 ;
      RECT 42.27 2.027 42.275 2.24 ;
      RECT 42.265 2.035 42.27 2.23 ;
      RECT 42.185 0.661 42.195 0.809 ;
      RECT 42.17 0.657 42.185 0.807 ;
      RECT 42.16 0.652 42.17 0.803 ;
      RECT 42.135 0.645 42.16 0.795 ;
      RECT 42.13 0.64 42.135 0.79 ;
      RECT 42.12 0.64 42.13 0.788 ;
      RECT 42.11 0.638 42.12 0.786 ;
      RECT 42.08 0.63 42.11 0.78 ;
      RECT 42.065 0.622 42.08 0.773 ;
      RECT 42.045 0.617 42.065 0.766 ;
      RECT 42.04 0.613 42.045 0.761 ;
      RECT 42.01 0.606 42.04 0.755 ;
      RECT 41.985 0.597 42.01 0.745 ;
      RECT 41.955 0.59 41.985 0.737 ;
      RECT 41.93 0.58 41.955 0.728 ;
      RECT 41.915 0.572 41.93 0.722 ;
      RECT 41.89 0.567 41.915 0.717 ;
      RECT 41.88 0.563 41.89 0.712 ;
      RECT 41.86 0.558 41.88 0.707 ;
      RECT 41.825 0.553 41.86 0.7 ;
      RECT 41.765 0.548 41.825 0.693 ;
      RECT 41.752 0.544 41.765 0.691 ;
      RECT 41.666 0.539 41.752 0.688 ;
      RECT 41.58 0.529 41.666 0.684 ;
      RECT 41.539 0.522 41.58 0.681 ;
      RECT 41.453 0.515 41.539 0.678 ;
      RECT 41.367 0.505 41.453 0.674 ;
      RECT 41.281 0.495 41.367 0.669 ;
      RECT 41.195 0.485 41.281 0.665 ;
      RECT 41.185 0.47 41.195 0.663 ;
      RECT 41.175 0.455 41.185 0.663 ;
      RECT 41.11 0.45 41.175 0.662 ;
      RECT 40.945 0.447 40.99 0.655 ;
      RECT 42.19 1.352 42.195 1.543 ;
      RECT 42.185 1.347 42.19 1.55 ;
      RECT 42.171 1.345 42.185 1.556 ;
      RECT 42.085 1.345 42.171 1.558 ;
      RECT 42.081 1.345 42.085 1.561 ;
      RECT 41.995 1.345 42.081 1.579 ;
      RECT 41.985 1.35 41.995 1.598 ;
      RECT 41.975 1.405 41.985 1.602 ;
      RECT 41.95 1.42 41.975 1.609 ;
      RECT 41.91 1.44 41.95 1.622 ;
      RECT 41.905 1.452 41.91 1.632 ;
      RECT 41.89 1.458 41.905 1.637 ;
      RECT 41.885 1.463 41.89 1.641 ;
      RECT 41.865 1.47 41.885 1.646 ;
      RECT 41.795 1.495 41.865 1.663 ;
      RECT 41.755 1.523 41.795 1.683 ;
      RECT 41.75 1.533 41.755 1.691 ;
      RECT 41.73 1.54 41.75 1.693 ;
      RECT 41.725 1.547 41.73 1.696 ;
      RECT 41.695 1.555 41.725 1.699 ;
      RECT 41.69 1.56 41.695 1.703 ;
      RECT 41.616 1.564 41.69 1.711 ;
      RECT 41.53 1.573 41.616 1.727 ;
      RECT 41.526 1.578 41.53 1.736 ;
      RECT 41.44 1.583 41.526 1.746 ;
      RECT 41.4 1.591 41.44 1.758 ;
      RECT 41.35 1.597 41.4 1.765 ;
      RECT 41.265 1.606 41.35 1.78 ;
      RECT 41.19 1.617 41.265 1.798 ;
      RECT 41.155 1.624 41.19 1.808 ;
      RECT 41.08 1.632 41.155 1.813 ;
      RECT 41.025 1.641 41.08 1.813 ;
      RECT 41 1.646 41.025 1.811 ;
      RECT 40.99 1.649 41 1.809 ;
      RECT 40.955 1.651 40.99 1.807 ;
      RECT 40.925 1.653 40.955 1.803 ;
      RECT 40.88 1.652 40.925 1.799 ;
      RECT 40.86 1.647 40.88 1.796 ;
      RECT 40.81 1.632 40.86 1.793 ;
      RECT 40.8 1.617 40.81 1.788 ;
      RECT 40.75 1.602 40.8 1.778 ;
      RECT 40.7 1.577 40.75 1.758 ;
      RECT 40.69 1.562 40.7 1.74 ;
      RECT 40.685 1.56 40.69 1.734 ;
      RECT 40.665 1.555 40.685 1.729 ;
      RECT 40.66 1.547 40.665 1.723 ;
      RECT 40.645 1.541 40.66 1.716 ;
      RECT 40.64 1.536 40.645 1.708 ;
      RECT 40.62 1.531 40.64 1.7 ;
      RECT 40.605 1.524 40.62 1.693 ;
      RECT 40.59 1.518 40.605 1.684 ;
      RECT 40.585 1.512 40.59 1.677 ;
      RECT 40.54 1.487 40.585 1.663 ;
      RECT 40.525 1.457 40.54 1.645 ;
      RECT 40.51 1.44 40.525 1.636 ;
      RECT 40.485 1.42 40.51 1.624 ;
      RECT 40.445 1.39 40.485 1.604 ;
      RECT 40.435 1.36 40.445 1.589 ;
      RECT 40.42 1.35 40.435 1.582 ;
      RECT 40.365 1.315 40.42 1.561 ;
      RECT 40.35 1.278 40.365 1.54 ;
      RECT 40.34 1.265 40.35 1.532 ;
      RECT 40.29 1.235 40.34 1.514 ;
      RECT 40.275 1.165 40.29 1.495 ;
      RECT 40.23 1.165 40.275 1.478 ;
      RECT 40.205 1.165 40.23 1.46 ;
      RECT 40.195 1.165 40.205 1.453 ;
      RECT 40.116 1.165 40.195 1.446 ;
      RECT 40.03 1.165 40.116 1.438 ;
      RECT 40.015 1.197 40.03 1.433 ;
      RECT 39.94 1.207 40.015 1.429 ;
      RECT 39.92 1.217 39.94 1.424 ;
      RECT 39.895 1.217 39.92 1.421 ;
      RECT 39.885 1.207 39.895 1.42 ;
      RECT 39.875 1.18 39.885 1.419 ;
      RECT 39.835 1.175 39.875 1.417 ;
      RECT 39.79 1.175 39.835 1.413 ;
      RECT 39.765 1.175 39.79 1.408 ;
      RECT 39.715 1.175 39.765 1.395 ;
      RECT 39.675 1.18 39.685 1.38 ;
      RECT 39.685 1.175 39.715 1.385 ;
      RECT 41.67 0.955 41.93 1.215 ;
      RECT 41.665 0.977 41.93 1.173 ;
      RECT 40.905 0.805 41.125 1.17 ;
      RECT 40.887 0.892 41.125 1.169 ;
      RECT 40.87 0.897 41.125 1.166 ;
      RECT 40.87 0.897 41.145 1.165 ;
      RECT 40.84 0.907 41.145 1.163 ;
      RECT 40.835 0.922 41.145 1.159 ;
      RECT 40.835 0.922 41.15 1.158 ;
      RECT 40.83 0.98 41.15 1.156 ;
      RECT 40.83 0.98 41.16 1.153 ;
      RECT 40.825 1.045 41.16 1.148 ;
      RECT 40.905 0.805 41.165 1.065 ;
      RECT 39.65 0.635 39.91 0.895 ;
      RECT 39.65 0.678 39.996 0.869 ;
      RECT 39.65 0.678 40.04 0.868 ;
      RECT 39.65 0.678 40.06 0.866 ;
      RECT 39.65 0.678 40.16 0.865 ;
      RECT 39.65 0.678 40.18 0.863 ;
      RECT 39.65 0.678 40.19 0.858 ;
      RECT 40.06 0.645 40.25 0.855 ;
      RECT 40.06 0.647 40.255 0.853 ;
      RECT 40.05 0.652 40.26 0.845 ;
      RECT 39.996 0.676 40.26 0.845 ;
      RECT 40.04 0.67 40.05 0.867 ;
      RECT 40.05 0.65 40.255 0.853 ;
      RECT 39.005 1.71 39.21 1.94 ;
      RECT 38.945 1.66 39 1.92 ;
      RECT 39.005 1.66 39.205 1.94 ;
      RECT 39.975 1.975 39.98 2.002 ;
      RECT 39.965 1.885 39.975 2.007 ;
      RECT 39.96 1.807 39.965 2.013 ;
      RECT 39.95 1.797 39.96 2.02 ;
      RECT 39.945 1.787 39.95 2.026 ;
      RECT 39.935 1.782 39.945 2.028 ;
      RECT 39.92 1.774 39.935 2.036 ;
      RECT 39.905 1.765 39.92 2.048 ;
      RECT 39.895 1.757 39.905 2.058 ;
      RECT 39.86 1.675 39.895 2.076 ;
      RECT 39.825 1.675 39.86 2.095 ;
      RECT 39.81 1.675 39.825 2.103 ;
      RECT 39.755 1.675 39.81 2.103 ;
      RECT 39.721 1.675 39.755 2.094 ;
      RECT 39.635 1.675 39.721 2.07 ;
      RECT 39.625 1.735 39.635 2.052 ;
      RECT 39.585 1.737 39.625 2.043 ;
      RECT 39.58 1.739 39.585 2.033 ;
      RECT 39.56 1.741 39.58 2.028 ;
      RECT 39.55 1.744 39.56 2.023 ;
      RECT 39.54 1.745 39.55 2.018 ;
      RECT 39.516 1.746 39.54 2.01 ;
      RECT 39.43 1.751 39.516 1.988 ;
      RECT 39.375 1.75 39.43 1.961 ;
      RECT 39.36 1.743 39.375 1.948 ;
      RECT 39.325 1.738 39.36 1.944 ;
      RECT 39.27 1.73 39.325 1.943 ;
      RECT 39.21 1.717 39.27 1.941 ;
      RECT 39 1.66 39.005 1.928 ;
      RECT 39.075 1.03 39.26 1.24 ;
      RECT 39.065 1.035 39.275 1.233 ;
      RECT 39.105 0.94 39.365 1.2 ;
      RECT 39.06 1.097 39.365 1.123 ;
      RECT 38.405 0.89 38.41 1.69 ;
      RECT 38.35 0.94 38.38 1.69 ;
      RECT 38.34 0.94 38.345 1.25 ;
      RECT 38.325 0.94 38.33 1.245 ;
      RECT 37.87 0.985 37.885 1.2 ;
      RECT 37.8 0.985 37.885 1.195 ;
      RECT 39.065 0.565 39.135 0.775 ;
      RECT 39.135 0.572 39.145 0.77 ;
      RECT 39.031 0.565 39.065 0.782 ;
      RECT 38.945 0.565 39.031 0.806 ;
      RECT 38.935 0.57 38.945 0.825 ;
      RECT 38.93 0.582 38.935 0.828 ;
      RECT 38.915 0.597 38.93 0.832 ;
      RECT 38.91 0.615 38.915 0.836 ;
      RECT 38.87 0.625 38.91 0.845 ;
      RECT 38.855 0.632 38.87 0.857 ;
      RECT 38.84 0.637 38.855 0.862 ;
      RECT 38.825 0.64 38.84 0.867 ;
      RECT 38.815 0.642 38.825 0.871 ;
      RECT 38.78 0.649 38.815 0.879 ;
      RECT 38.745 0.657 38.78 0.893 ;
      RECT 38.735 0.663 38.745 0.902 ;
      RECT 38.73 0.665 38.735 0.904 ;
      RECT 38.71 0.668 38.73 0.91 ;
      RECT 38.68 0.675 38.71 0.921 ;
      RECT 38.67 0.681 38.68 0.928 ;
      RECT 38.645 0.684 38.67 0.935 ;
      RECT 38.635 0.688 38.645 0.943 ;
      RECT 38.63 0.689 38.635 0.965 ;
      RECT 38.625 0.69 38.63 0.98 ;
      RECT 38.62 0.691 38.625 0.995 ;
      RECT 38.615 0.692 38.62 1.01 ;
      RECT 38.61 0.693 38.615 1.04 ;
      RECT 38.6 0.695 38.61 1.073 ;
      RECT 38.585 0.699 38.6 1.12 ;
      RECT 38.575 0.702 38.585 1.165 ;
      RECT 38.57 0.705 38.575 1.193 ;
      RECT 38.56 0.707 38.57 1.22 ;
      RECT 38.555 0.71 38.56 1.255 ;
      RECT 38.525 0.715 38.555 1.313 ;
      RECT 38.52 0.72 38.525 1.398 ;
      RECT 38.515 0.722 38.52 1.433 ;
      RECT 38.51 0.724 38.515 1.515 ;
      RECT 38.505 0.726 38.51 1.603 ;
      RECT 38.495 0.728 38.505 1.685 ;
      RECT 38.48 0.742 38.495 1.69 ;
      RECT 38.445 0.787 38.48 1.69 ;
      RECT 38.435 0.827 38.445 1.69 ;
      RECT 38.42 0.855 38.435 1.69 ;
      RECT 38.415 0.872 38.42 1.69 ;
      RECT 38.41 0.88 38.415 1.69 ;
      RECT 38.4 0.895 38.405 1.69 ;
      RECT 38.395 0.902 38.4 1.69 ;
      RECT 38.385 0.922 38.395 1.69 ;
      RECT 38.38 0.935 38.385 1.69 ;
      RECT 38.345 0.94 38.35 1.275 ;
      RECT 38.33 1.33 38.35 1.69 ;
      RECT 38.33 0.94 38.34 1.248 ;
      RECT 38.325 1.37 38.33 1.69 ;
      RECT 38.275 0.94 38.325 1.243 ;
      RECT 38.32 1.407 38.325 1.69 ;
      RECT 38.31 1.43 38.32 1.69 ;
      RECT 38.305 1.475 38.31 1.69 ;
      RECT 38.295 1.485 38.305 1.683 ;
      RECT 38.221 0.94 38.275 1.237 ;
      RECT 38.135 0.94 38.221 1.23 ;
      RECT 38.086 0.987 38.135 1.223 ;
      RECT 38 0.995 38.086 1.216 ;
      RECT 37.985 0.992 38 1.211 ;
      RECT 37.971 0.985 37.985 1.21 ;
      RECT 37.885 0.985 37.971 1.205 ;
      RECT 37.79 0.99 37.8 1.19 ;
      RECT 37.38 0.42 37.395 0.82 ;
      RECT 37.575 0.42 37.58 0.68 ;
      RECT 37.32 0.42 37.365 0.68 ;
      RECT 37.775 1.725 37.78 1.93 ;
      RECT 37.77 1.715 37.775 1.935 ;
      RECT 37.765 1.702 37.77 1.94 ;
      RECT 37.76 1.682 37.765 1.94 ;
      RECT 37.735 1.635 37.76 1.94 ;
      RECT 37.7 1.55 37.735 1.94 ;
      RECT 37.695 1.487 37.7 1.94 ;
      RECT 37.69 1.472 37.695 1.94 ;
      RECT 37.675 1.432 37.69 1.94 ;
      RECT 37.67 1.407 37.675 1.94 ;
      RECT 37.66 1.39 37.67 1.94 ;
      RECT 37.625 1.312 37.66 1.94 ;
      RECT 37.62 1.255 37.625 1.94 ;
      RECT 37.615 1.242 37.62 1.94 ;
      RECT 37.605 1.22 37.615 1.94 ;
      RECT 37.595 1.185 37.605 1.94 ;
      RECT 37.585 1.155 37.595 1.94 ;
      RECT 37.575 1.07 37.585 1.583 ;
      RECT 37.582 1.715 37.585 1.94 ;
      RECT 37.58 1.725 37.582 1.94 ;
      RECT 37.57 1.735 37.58 1.935 ;
      RECT 37.565 0.42 37.575 0.815 ;
      RECT 37.57 0.947 37.575 1.558 ;
      RECT 37.565 0.845 37.57 1.541 ;
      RECT 37.555 0.42 37.565 1.517 ;
      RECT 37.55 0.42 37.555 1.488 ;
      RECT 37.545 0.42 37.55 1.478 ;
      RECT 37.525 0.42 37.545 1.44 ;
      RECT 37.52 0.42 37.525 1.398 ;
      RECT 37.515 0.42 37.52 1.378 ;
      RECT 37.485 0.42 37.515 1.328 ;
      RECT 37.475 0.42 37.485 1.275 ;
      RECT 37.47 0.42 37.475 1.248 ;
      RECT 37.465 0.42 37.47 1.233 ;
      RECT 37.455 0.42 37.465 1.21 ;
      RECT 37.445 0.42 37.455 1.185 ;
      RECT 37.44 0.42 37.445 1.125 ;
      RECT 37.43 0.42 37.44 1.063 ;
      RECT 37.425 0.42 37.43 0.983 ;
      RECT 37.42 0.42 37.425 0.948 ;
      RECT 37.415 0.42 37.42 0.923 ;
      RECT 37.41 0.42 37.415 0.908 ;
      RECT 37.405 0.42 37.41 0.878 ;
      RECT 37.4 0.42 37.405 0.855 ;
      RECT 37.395 0.42 37.4 0.828 ;
      RECT 37.365 0.42 37.38 0.815 ;
      RECT 36.52 1.955 36.705 2.165 ;
      RECT 36.51 1.96 36.72 2.158 ;
      RECT 36.51 1.96 36.74 2.13 ;
      RECT 36.51 1.96 36.755 2.109 ;
      RECT 36.51 1.96 36.77 2.107 ;
      RECT 36.51 1.96 36.78 2.106 ;
      RECT 36.51 1.96 36.81 2.103 ;
      RECT 37.16 1.805 37.42 2.065 ;
      RECT 37.12 1.852 37.42 2.048 ;
      RECT 37.111 1.86 37.12 2.051 ;
      RECT 36.705 1.953 37.42 2.048 ;
      RECT 37.025 1.878 37.111 2.058 ;
      RECT 36.72 1.95 37.42 2.048 ;
      RECT 36.966 1.9 37.025 2.07 ;
      RECT 36.74 1.946 37.42 2.048 ;
      RECT 36.88 1.912 36.966 2.081 ;
      RECT 36.755 1.942 37.42 2.048 ;
      RECT 36.825 1.925 36.88 2.093 ;
      RECT 36.77 1.94 37.42 2.048 ;
      RECT 36.81 1.931 36.825 2.099 ;
      RECT 36.78 1.936 37.42 2.048 ;
      RECT 36.925 1.46 37.185 1.72 ;
      RECT 36.925 1.48 37.295 1.69 ;
      RECT 36.925 1.485 37.305 1.685 ;
      RECT 37.116 0.899 37.195 1.13 ;
      RECT 37.03 0.902 37.245 1.125 ;
      RECT 37.025 0.902 37.245 1.12 ;
      RECT 37.025 0.907 37.255 1.118 ;
      RECT 37 0.907 37.255 1.115 ;
      RECT 37 0.915 37.265 1.113 ;
      RECT 36.88 0.85 37.14 1.11 ;
      RECT 36.88 0.897 37.19 1.11 ;
      RECT 36.135 1.47 36.14 1.73 ;
      RECT 35.965 1.24 35.97 1.73 ;
      RECT 35.85 1.48 35.855 1.705 ;
      RECT 36.56 0.575 36.565 0.785 ;
      RECT 36.565 0.58 36.58 0.78 ;
      RECT 36.5 0.575 36.56 0.793 ;
      RECT 36.485 0.575 36.5 0.803 ;
      RECT 36.435 0.575 36.485 0.82 ;
      RECT 36.415 0.575 36.435 0.843 ;
      RECT 36.4 0.575 36.415 0.855 ;
      RECT 36.38 0.575 36.4 0.865 ;
      RECT 36.37 0.58 36.38 0.874 ;
      RECT 36.365 0.59 36.37 0.879 ;
      RECT 36.36 0.602 36.365 0.883 ;
      RECT 36.35 0.625 36.36 0.888 ;
      RECT 36.345 0.64 36.35 0.892 ;
      RECT 36.34 0.657 36.345 0.895 ;
      RECT 36.335 0.665 36.34 0.898 ;
      RECT 36.325 0.67 36.335 0.902 ;
      RECT 36.32 0.677 36.325 0.907 ;
      RECT 36.31 0.682 36.32 0.911 ;
      RECT 36.285 0.694 36.31 0.922 ;
      RECT 36.265 0.711 36.285 0.938 ;
      RECT 36.24 0.728 36.265 0.96 ;
      RECT 36.205 0.751 36.24 1.018 ;
      RECT 36.185 0.773 36.205 1.08 ;
      RECT 36.18 0.783 36.185 1.115 ;
      RECT 36.17 0.79 36.18 1.153 ;
      RECT 36.165 0.797 36.17 1.173 ;
      RECT 36.16 0.808 36.165 1.21 ;
      RECT 36.155 0.816 36.16 1.275 ;
      RECT 36.145 0.827 36.155 1.328 ;
      RECT 36.14 0.845 36.145 1.398 ;
      RECT 36.135 0.855 36.14 1.435 ;
      RECT 36.13 0.865 36.135 1.73 ;
      RECT 36.125 0.877 36.13 1.73 ;
      RECT 36.12 0.887 36.125 1.73 ;
      RECT 36.11 0.897 36.12 1.73 ;
      RECT 36.1 0.92 36.11 1.73 ;
      RECT 36.085 0.955 36.1 1.73 ;
      RECT 36.045 1.017 36.085 1.73 ;
      RECT 36.04 1.07 36.045 1.73 ;
      RECT 36.015 1.105 36.04 1.73 ;
      RECT 36 1.15 36.015 1.73 ;
      RECT 35.995 1.172 36 1.73 ;
      RECT 35.985 1.185 35.995 1.73 ;
      RECT 35.975 1.21 35.985 1.73 ;
      RECT 35.97 1.232 35.975 1.73 ;
      RECT 35.945 1.27 35.965 1.73 ;
      RECT 35.905 1.327 35.945 1.73 ;
      RECT 35.9 1.377 35.905 1.73 ;
      RECT 35.895 1.395 35.9 1.73 ;
      RECT 35.89 1.407 35.895 1.73 ;
      RECT 35.88 1.425 35.89 1.73 ;
      RECT 35.87 1.445 35.88 1.705 ;
      RECT 35.865 1.462 35.87 1.705 ;
      RECT 35.855 1.475 35.865 1.705 ;
      RECT 35.825 1.485 35.85 1.705 ;
      RECT 35.815 1.492 35.825 1.705 ;
      RECT 35.8 1.502 35.815 1.7 ;
      RECT 34.76 1.415 35.08 1.675 ;
      RECT 34.625 1.46 35.08 1.63 ;
      RECT 28.32 1.475 28.695 1.725 ;
      RECT 28.415 0.73 28.59 1.725 ;
      RECT 28.415 0.73 34.34 0.905 ;
      RECT 33.905 0.475 34.225 0.905 ;
      RECT 33.905 0.505 34.305 0.675 ;
      RECT 31.57 1.515 31.865 1.805 ;
      RECT 31.54 1.515 31.865 1.775 ;
      RECT 17.78 1.885 18.085 2.115 ;
      RECT 25.92 1.915 29.335 2.09 ;
      RECT 29.16 1.065 29.335 2.09 ;
      RECT 17.78 1.915 29.335 2.085 ;
      RECT 29.105 1.065 29.435 1.315 ;
      RECT 26.365 1.075 26.655 1.315 ;
      RECT 21.915 1.045 22.175 1.28 ;
      RECT 21.915 1.075 26.655 1.245 ;
      RECT 25.1 1.415 25.42 1.675 ;
      RECT 25.085 1.46 25.42 1.63 ;
      RECT 23.805 0.395 24.1 0.685 ;
      RECT 23.77 0.395 24.1 0.655 ;
      RECT 20.965 1.415 21.285 1.675 ;
      RECT 20.95 1.46 21.285 1.63 ;
      RECT 19.29 1.205 19.61 1.465 ;
      RECT 19.275 1.205 19.63 1.44 ;
      RECT 16.59 0.965 16.775 1.175 ;
      RECT 16.58 0.97 16.79 1.168 ;
      RECT 16.58 0.97 16.876 1.145 ;
      RECT 16.58 0.97 16.935 1.12 ;
      RECT 16.58 0.97 16.99 1.1 ;
      RECT 16.58 0.97 17 1.088 ;
      RECT 16.58 0.97 17.195 1.027 ;
      RECT 16.58 0.97 17.225 1.01 ;
      RECT 16.58 0.97 17.245 1 ;
      RECT 17.125 0.735 17.385 0.995 ;
      RECT 17.11 0.825 17.125 1.042 ;
      RECT 16.645 0.957 17.385 0.995 ;
      RECT 17.096 0.836 17.11 1.048 ;
      RECT 16.685 0.95 17.385 0.995 ;
      RECT 17.01 0.876 17.096 1.067 ;
      RECT 16.935 0.937 17.385 0.995 ;
      RECT 17.005 0.912 17.01 1.084 ;
      RECT 16.99 0.922 17.385 0.995 ;
      RECT 17 0.917 17.005 1.086 ;
      RECT 17.295 1.422 17.3 1.514 ;
      RECT 17.29 1.4 17.295 1.531 ;
      RECT 17.285 1.39 17.29 1.543 ;
      RECT 17.275 1.381 17.285 1.553 ;
      RECT 17.27 1.376 17.275 1.561 ;
      RECT 17.265 1.372 17.27 1.564 ;
      RECT 17.231 1.305 17.265 1.575 ;
      RECT 17.145 1.305 17.231 1.61 ;
      RECT 17.065 1.305 17.145 1.658 ;
      RECT 17.005 1.305 17.065 1.683 ;
      RECT 16.945 1.405 17.005 1.69 ;
      RECT 16.91 1.43 16.945 1.696 ;
      RECT 16.885 1.445 16.91 1.7 ;
      RECT 16.871 1.454 16.885 1.702 ;
      RECT 16.785 1.481 16.871 1.708 ;
      RECT 16.72 1.522 16.785 1.717 ;
      RECT 16.705 1.542 16.72 1.722 ;
      RECT 16.675 1.552 16.705 1.725 ;
      RECT 16.67 1.562 16.675 1.728 ;
      RECT 16.64 1.567 16.67 1.73 ;
      RECT 16.62 1.572 16.64 1.734 ;
      RECT 16.535 1.575 16.62 1.741 ;
      RECT 16.52 1.572 16.535 1.747 ;
      RECT 16.51 1.569 16.52 1.749 ;
      RECT 16.49 1.566 16.51 1.751 ;
      RECT 16.47 1.562 16.49 1.752 ;
      RECT 16.455 1.558 16.47 1.754 ;
      RECT 16.445 1.555 16.455 1.755 ;
      RECT 16.405 1.549 16.445 1.753 ;
      RECT 16.395 1.544 16.405 1.751 ;
      RECT 16.38 1.541 16.395 1.747 ;
      RECT 16.355 1.536 16.38 1.74 ;
      RECT 16.305 1.527 16.355 1.728 ;
      RECT 16.235 1.513 16.305 1.71 ;
      RECT 16.177 1.498 16.235 1.692 ;
      RECT 16.091 1.481 16.177 1.672 ;
      RECT 16.005 1.46 16.091 1.647 ;
      RECT 15.955 1.445 16.005 1.628 ;
      RECT 15.951 1.439 15.955 1.62 ;
      RECT 15.865 1.429 15.951 1.607 ;
      RECT 15.83 1.414 15.865 1.59 ;
      RECT 15.815 1.407 15.83 1.583 ;
      RECT 15.755 1.395 15.815 1.571 ;
      RECT 15.735 1.382 15.755 1.559 ;
      RECT 15.695 1.373 15.735 1.551 ;
      RECT 15.69 1.365 15.695 1.544 ;
      RECT 15.61 1.355 15.69 1.53 ;
      RECT 15.595 1.342 15.61 1.515 ;
      RECT 15.59 1.34 15.595 1.513 ;
      RECT 15.511 1.328 15.59 1.5 ;
      RECT 15.425 1.303 15.511 1.475 ;
      RECT 15.41 1.272 15.425 1.46 ;
      RECT 15.395 1.247 15.41 1.456 ;
      RECT 15.38 1.24 15.395 1.452 ;
      RECT 15.205 1.245 15.21 1.448 ;
      RECT 15.2 1.25 15.205 1.443 ;
      RECT 15.21 1.24 15.38 1.45 ;
      RECT 15.925 1 16.03 1.26 ;
      RECT 16.74 0.525 16.745 0.75 ;
      RECT 16.87 0.525 16.925 0.735 ;
      RECT 16.925 0.53 16.935 0.728 ;
      RECT 16.831 0.525 16.87 0.738 ;
      RECT 16.745 0.525 16.831 0.745 ;
      RECT 16.725 0.53 16.74 0.751 ;
      RECT 16.715 0.57 16.725 0.753 ;
      RECT 16.685 0.58 16.715 0.755 ;
      RECT 16.68 0.585 16.685 0.757 ;
      RECT 16.655 0.59 16.68 0.759 ;
      RECT 16.64 0.595 16.655 0.761 ;
      RECT 16.625 0.597 16.64 0.763 ;
      RECT 16.62 0.602 16.625 0.765 ;
      RECT 16.57 0.61 16.62 0.768 ;
      RECT 16.545 0.619 16.57 0.773 ;
      RECT 16.535 0.626 16.545 0.778 ;
      RECT 16.53 0.629 16.535 0.782 ;
      RECT 16.51 0.632 16.53 0.791 ;
      RECT 16.48 0.64 16.51 0.811 ;
      RECT 16.451 0.653 16.48 0.833 ;
      RECT 16.365 0.687 16.451 0.877 ;
      RECT 16.36 0.713 16.365 0.915 ;
      RECT 16.355 0.717 16.36 0.924 ;
      RECT 16.32 0.73 16.355 0.957 ;
      RECT 16.31 0.744 16.32 0.995 ;
      RECT 16.305 0.748 16.31 1.008 ;
      RECT 16.3 0.752 16.305 1.013 ;
      RECT 16.29 0.76 16.3 1.025 ;
      RECT 16.285 0.767 16.29 1.04 ;
      RECT 16.26 0.78 16.285 1.065 ;
      RECT 16.22 0.809 16.26 1.12 ;
      RECT 16.205 0.834 16.22 1.175 ;
      RECT 16.195 0.845 16.205 1.198 ;
      RECT 16.19 0.852 16.195 1.21 ;
      RECT 16.185 0.856 16.19 1.218 ;
      RECT 16.13 0.884 16.185 1.26 ;
      RECT 16.11 0.92 16.13 1.26 ;
      RECT 16.095 0.935 16.11 1.26 ;
      RECT 16.04 0.967 16.095 1.26 ;
      RECT 16.03 0.997 16.04 1.26 ;
      RECT 15.64 0.612 15.825 0.85 ;
      RECT 15.625 0.614 15.835 0.845 ;
      RECT 15.51 0.56 15.77 0.82 ;
      RECT 15.505 0.597 15.77 0.774 ;
      RECT 15.5 0.607 15.77 0.771 ;
      RECT 15.495 0.647 15.835 0.765 ;
      RECT 15.49 0.68 15.835 0.755 ;
      RECT 15.5 0.622 15.85 0.693 ;
      RECT 15.797 1.72 15.81 2.25 ;
      RECT 15.711 1.72 15.81 2.249 ;
      RECT 15.711 1.72 15.815 2.248 ;
      RECT 15.625 1.72 15.815 2.246 ;
      RECT 15.62 1.72 15.815 2.243 ;
      RECT 15.62 1.72 15.825 2.241 ;
      RECT 15.615 2.012 15.825 2.238 ;
      RECT 15.615 2.022 15.83 2.235 ;
      RECT 15.615 2.09 15.835 2.231 ;
      RECT 15.605 2.095 15.835 2.23 ;
      RECT 15.605 2.187 15.84 2.227 ;
      RECT 15.59 1.72 15.85 1.98 ;
      RECT 14.82 0.71 14.865 2.245 ;
      RECT 15.02 0.71 15.05 0.925 ;
      RECT 13.395 0.45 13.515 0.66 ;
      RECT 13.055 0.4 13.315 0.66 ;
      RECT 13.055 0.445 13.35 0.65 ;
      RECT 15.06 0.726 15.065 0.78 ;
      RECT 15.055 0.719 15.06 0.913 ;
      RECT 15.05 0.713 15.055 0.92 ;
      RECT 15.005 0.71 15.02 0.933 ;
      RECT 15 0.71 15.005 0.955 ;
      RECT 14.995 0.71 15 1.003 ;
      RECT 14.99 0.71 14.995 1.023 ;
      RECT 14.98 0.71 14.99 1.13 ;
      RECT 14.975 0.71 14.98 1.193 ;
      RECT 14.97 0.71 14.975 1.25 ;
      RECT 14.965 0.71 14.97 1.258 ;
      RECT 14.95 0.71 14.965 1.365 ;
      RECT 14.94 0.71 14.95 1.5 ;
      RECT 14.93 0.71 14.94 1.61 ;
      RECT 14.92 0.71 14.93 1.667 ;
      RECT 14.915 0.71 14.92 1.707 ;
      RECT 14.91 0.71 14.915 1.743 ;
      RECT 14.9 0.71 14.91 1.783 ;
      RECT 14.895 0.71 14.9 1.825 ;
      RECT 14.875 0.71 14.895 1.89 ;
      RECT 14.88 2.035 14.885 2.215 ;
      RECT 14.875 2.017 14.88 2.223 ;
      RECT 14.87 0.71 14.875 1.953 ;
      RECT 14.87 1.997 14.875 2.23 ;
      RECT 14.865 0.71 14.87 2.24 ;
      RECT 14.81 0.71 14.82 1.01 ;
      RECT 14.815 1.257 14.82 2.245 ;
      RECT 14.81 1.322 14.815 2.245 ;
      RECT 14.805 0.711 14.81 1 ;
      RECT 14.8 1.387 14.81 2.245 ;
      RECT 14.795 0.712 14.805 0.99 ;
      RECT 14.785 1.5 14.8 2.245 ;
      RECT 14.79 0.713 14.795 0.98 ;
      RECT 14.77 0.714 14.79 0.958 ;
      RECT 14.775 1.597 14.785 2.245 ;
      RECT 14.77 1.672 14.775 2.245 ;
      RECT 14.76 0.713 14.77 0.935 ;
      RECT 14.765 1.715 14.77 2.245 ;
      RECT 14.76 1.742 14.765 2.245 ;
      RECT 14.75 0.711 14.76 0.923 ;
      RECT 14.755 1.785 14.76 2.245 ;
      RECT 14.75 1.812 14.755 2.245 ;
      RECT 14.74 0.71 14.75 0.91 ;
      RECT 14.745 1.827 14.75 2.245 ;
      RECT 14.705 1.885 14.745 2.245 ;
      RECT 14.735 0.709 14.74 0.895 ;
      RECT 14.73 0.707 14.735 0.888 ;
      RECT 14.72 0.704 14.73 0.878 ;
      RECT 14.715 0.701 14.72 0.863 ;
      RECT 14.7 0.697 14.715 0.856 ;
      RECT 14.695 1.94 14.705 2.245 ;
      RECT 14.695 0.694 14.7 0.851 ;
      RECT 14.68 0.69 14.695 0.845 ;
      RECT 14.69 1.957 14.695 2.245 ;
      RECT 14.68 2.02 14.69 2.245 ;
      RECT 14.6 0.675 14.68 0.825 ;
      RECT 14.675 2.027 14.68 2.24 ;
      RECT 14.67 2.035 14.675 2.23 ;
      RECT 14.59 0.661 14.6 0.809 ;
      RECT 14.575 0.657 14.59 0.807 ;
      RECT 14.565 0.652 14.575 0.803 ;
      RECT 14.54 0.645 14.565 0.795 ;
      RECT 14.535 0.64 14.54 0.79 ;
      RECT 14.525 0.64 14.535 0.788 ;
      RECT 14.515 0.638 14.525 0.786 ;
      RECT 14.485 0.63 14.515 0.78 ;
      RECT 14.47 0.622 14.485 0.773 ;
      RECT 14.45 0.617 14.47 0.766 ;
      RECT 14.445 0.613 14.45 0.761 ;
      RECT 14.415 0.606 14.445 0.755 ;
      RECT 14.39 0.597 14.415 0.745 ;
      RECT 14.36 0.59 14.39 0.737 ;
      RECT 14.335 0.58 14.36 0.728 ;
      RECT 14.32 0.572 14.335 0.722 ;
      RECT 14.295 0.567 14.32 0.717 ;
      RECT 14.285 0.563 14.295 0.712 ;
      RECT 14.265 0.558 14.285 0.707 ;
      RECT 14.23 0.553 14.265 0.7 ;
      RECT 14.17 0.548 14.23 0.693 ;
      RECT 14.157 0.544 14.17 0.691 ;
      RECT 14.071 0.539 14.157 0.688 ;
      RECT 13.985 0.529 14.071 0.684 ;
      RECT 13.944 0.522 13.985 0.681 ;
      RECT 13.858 0.515 13.944 0.678 ;
      RECT 13.772 0.505 13.858 0.674 ;
      RECT 13.686 0.495 13.772 0.669 ;
      RECT 13.6 0.485 13.686 0.665 ;
      RECT 13.59 0.47 13.6 0.663 ;
      RECT 13.58 0.455 13.59 0.663 ;
      RECT 13.515 0.45 13.58 0.662 ;
      RECT 13.35 0.447 13.395 0.655 ;
      RECT 14.595 1.352 14.6 1.543 ;
      RECT 14.59 1.347 14.595 1.55 ;
      RECT 14.576 1.345 14.59 1.556 ;
      RECT 14.49 1.345 14.576 1.558 ;
      RECT 14.486 1.345 14.49 1.561 ;
      RECT 14.4 1.345 14.486 1.579 ;
      RECT 14.39 1.35 14.4 1.598 ;
      RECT 14.38 1.405 14.39 1.602 ;
      RECT 14.355 1.42 14.38 1.609 ;
      RECT 14.315 1.44 14.355 1.622 ;
      RECT 14.31 1.452 14.315 1.632 ;
      RECT 14.295 1.458 14.31 1.637 ;
      RECT 14.29 1.463 14.295 1.641 ;
      RECT 14.27 1.47 14.29 1.646 ;
      RECT 14.2 1.495 14.27 1.663 ;
      RECT 14.16 1.523 14.2 1.683 ;
      RECT 14.155 1.533 14.16 1.691 ;
      RECT 14.135 1.54 14.155 1.693 ;
      RECT 14.13 1.547 14.135 1.696 ;
      RECT 14.1 1.555 14.13 1.699 ;
      RECT 14.095 1.56 14.1 1.703 ;
      RECT 14.021 1.564 14.095 1.711 ;
      RECT 13.935 1.573 14.021 1.727 ;
      RECT 13.931 1.578 13.935 1.736 ;
      RECT 13.845 1.583 13.931 1.746 ;
      RECT 13.805 1.591 13.845 1.758 ;
      RECT 13.755 1.597 13.805 1.765 ;
      RECT 13.67 1.606 13.755 1.78 ;
      RECT 13.595 1.617 13.67 1.798 ;
      RECT 13.56 1.624 13.595 1.808 ;
      RECT 13.485 1.632 13.56 1.813 ;
      RECT 13.43 1.641 13.485 1.813 ;
      RECT 13.405 1.646 13.43 1.811 ;
      RECT 13.395 1.649 13.405 1.809 ;
      RECT 13.36 1.651 13.395 1.807 ;
      RECT 13.33 1.653 13.36 1.803 ;
      RECT 13.285 1.652 13.33 1.799 ;
      RECT 13.265 1.647 13.285 1.796 ;
      RECT 13.215 1.632 13.265 1.793 ;
      RECT 13.205 1.617 13.215 1.788 ;
      RECT 13.155 1.602 13.205 1.778 ;
      RECT 13.105 1.577 13.155 1.758 ;
      RECT 13.095 1.562 13.105 1.74 ;
      RECT 13.09 1.56 13.095 1.734 ;
      RECT 13.07 1.555 13.09 1.729 ;
      RECT 13.065 1.547 13.07 1.723 ;
      RECT 13.05 1.541 13.065 1.716 ;
      RECT 13.045 1.536 13.05 1.708 ;
      RECT 13.025 1.531 13.045 1.7 ;
      RECT 13.01 1.524 13.025 1.693 ;
      RECT 12.995 1.518 13.01 1.684 ;
      RECT 12.99 1.512 12.995 1.677 ;
      RECT 12.945 1.487 12.99 1.663 ;
      RECT 12.93 1.457 12.945 1.645 ;
      RECT 12.915 1.44 12.93 1.636 ;
      RECT 12.89 1.42 12.915 1.624 ;
      RECT 12.85 1.39 12.89 1.604 ;
      RECT 12.84 1.36 12.85 1.589 ;
      RECT 12.825 1.35 12.84 1.582 ;
      RECT 12.77 1.315 12.825 1.561 ;
      RECT 12.755 1.278 12.77 1.54 ;
      RECT 12.745 1.265 12.755 1.532 ;
      RECT 12.695 1.235 12.745 1.514 ;
      RECT 12.68 1.165 12.695 1.495 ;
      RECT 12.635 1.165 12.68 1.478 ;
      RECT 12.61 1.165 12.635 1.46 ;
      RECT 12.6 1.165 12.61 1.453 ;
      RECT 12.521 1.165 12.6 1.446 ;
      RECT 12.435 1.165 12.521 1.438 ;
      RECT 12.42 1.197 12.435 1.433 ;
      RECT 12.345 1.207 12.42 1.429 ;
      RECT 12.325 1.217 12.345 1.424 ;
      RECT 12.3 1.217 12.325 1.421 ;
      RECT 12.29 1.207 12.3 1.42 ;
      RECT 12.28 1.18 12.29 1.419 ;
      RECT 12.24 1.175 12.28 1.417 ;
      RECT 12.195 1.175 12.24 1.413 ;
      RECT 12.17 1.175 12.195 1.408 ;
      RECT 12.12 1.175 12.17 1.395 ;
      RECT 12.08 1.18 12.09 1.38 ;
      RECT 12.09 1.175 12.12 1.385 ;
      RECT 14.075 0.955 14.335 1.215 ;
      RECT 14.07 0.977 14.335 1.173 ;
      RECT 13.31 0.805 13.53 1.17 ;
      RECT 13.292 0.892 13.53 1.169 ;
      RECT 13.275 0.897 13.53 1.166 ;
      RECT 13.275 0.897 13.55 1.165 ;
      RECT 13.245 0.907 13.55 1.163 ;
      RECT 13.24 0.922 13.55 1.159 ;
      RECT 13.24 0.922 13.555 1.158 ;
      RECT 13.235 0.98 13.555 1.156 ;
      RECT 13.235 0.98 13.565 1.153 ;
      RECT 13.23 1.045 13.565 1.148 ;
      RECT 13.31 0.805 13.57 1.065 ;
      RECT 12.055 0.635 12.315 0.895 ;
      RECT 12.055 0.678 12.401 0.869 ;
      RECT 12.055 0.678 12.445 0.868 ;
      RECT 12.055 0.678 12.465 0.866 ;
      RECT 12.055 0.678 12.565 0.865 ;
      RECT 12.055 0.678 12.585 0.863 ;
      RECT 12.055 0.678 12.595 0.858 ;
      RECT 12.465 0.645 12.655 0.855 ;
      RECT 12.465 0.647 12.66 0.853 ;
      RECT 12.455 0.652 12.665 0.845 ;
      RECT 12.401 0.676 12.665 0.845 ;
      RECT 12.445 0.67 12.455 0.867 ;
      RECT 12.455 0.65 12.66 0.853 ;
      RECT 11.41 1.71 11.615 1.94 ;
      RECT 11.35 1.66 11.405 1.92 ;
      RECT 11.41 1.66 11.61 1.94 ;
      RECT 12.38 1.975 12.385 2.002 ;
      RECT 12.37 1.885 12.38 2.007 ;
      RECT 12.365 1.807 12.37 2.013 ;
      RECT 12.355 1.797 12.365 2.02 ;
      RECT 12.35 1.787 12.355 2.026 ;
      RECT 12.34 1.782 12.35 2.028 ;
      RECT 12.325 1.774 12.34 2.036 ;
      RECT 12.31 1.765 12.325 2.048 ;
      RECT 12.3 1.757 12.31 2.058 ;
      RECT 12.265 1.675 12.3 2.076 ;
      RECT 12.23 1.675 12.265 2.095 ;
      RECT 12.215 1.675 12.23 2.103 ;
      RECT 12.16 1.675 12.215 2.103 ;
      RECT 12.126 1.675 12.16 2.094 ;
      RECT 12.04 1.675 12.126 2.07 ;
      RECT 12.03 1.735 12.04 2.052 ;
      RECT 11.99 1.737 12.03 2.043 ;
      RECT 11.985 1.739 11.99 2.033 ;
      RECT 11.965 1.741 11.985 2.028 ;
      RECT 11.955 1.744 11.965 2.023 ;
      RECT 11.945 1.745 11.955 2.018 ;
      RECT 11.921 1.746 11.945 2.01 ;
      RECT 11.835 1.751 11.921 1.988 ;
      RECT 11.78 1.75 11.835 1.961 ;
      RECT 11.765 1.743 11.78 1.948 ;
      RECT 11.73 1.738 11.765 1.944 ;
      RECT 11.675 1.73 11.73 1.943 ;
      RECT 11.615 1.717 11.675 1.941 ;
      RECT 11.405 1.66 11.41 1.928 ;
      RECT 11.48 1.03 11.665 1.24 ;
      RECT 11.47 1.035 11.68 1.233 ;
      RECT 11.51 0.94 11.77 1.2 ;
      RECT 11.465 1.097 11.77 1.123 ;
      RECT 10.81 0.89 10.815 1.69 ;
      RECT 10.755 0.94 10.785 1.69 ;
      RECT 10.745 0.94 10.75 1.25 ;
      RECT 10.73 0.94 10.735 1.245 ;
      RECT 10.275 0.985 10.29 1.2 ;
      RECT 10.205 0.985 10.29 1.195 ;
      RECT 11.47 0.565 11.54 0.775 ;
      RECT 11.54 0.572 11.55 0.77 ;
      RECT 11.436 0.565 11.47 0.782 ;
      RECT 11.35 0.565 11.436 0.806 ;
      RECT 11.34 0.57 11.35 0.825 ;
      RECT 11.335 0.582 11.34 0.828 ;
      RECT 11.32 0.597 11.335 0.832 ;
      RECT 11.315 0.615 11.32 0.836 ;
      RECT 11.275 0.625 11.315 0.845 ;
      RECT 11.26 0.632 11.275 0.857 ;
      RECT 11.245 0.637 11.26 0.862 ;
      RECT 11.23 0.64 11.245 0.867 ;
      RECT 11.22 0.642 11.23 0.871 ;
      RECT 11.185 0.649 11.22 0.879 ;
      RECT 11.15 0.657 11.185 0.893 ;
      RECT 11.14 0.663 11.15 0.902 ;
      RECT 11.135 0.665 11.14 0.904 ;
      RECT 11.115 0.668 11.135 0.91 ;
      RECT 11.085 0.675 11.115 0.921 ;
      RECT 11.075 0.681 11.085 0.928 ;
      RECT 11.05 0.684 11.075 0.935 ;
      RECT 11.04 0.688 11.05 0.943 ;
      RECT 11.035 0.689 11.04 0.965 ;
      RECT 11.03 0.69 11.035 0.98 ;
      RECT 11.025 0.691 11.03 0.995 ;
      RECT 11.02 0.692 11.025 1.01 ;
      RECT 11.015 0.693 11.02 1.04 ;
      RECT 11.005 0.695 11.015 1.073 ;
      RECT 10.99 0.699 11.005 1.12 ;
      RECT 10.98 0.702 10.99 1.165 ;
      RECT 10.975 0.705 10.98 1.193 ;
      RECT 10.965 0.707 10.975 1.22 ;
      RECT 10.96 0.71 10.965 1.255 ;
      RECT 10.93 0.715 10.96 1.313 ;
      RECT 10.925 0.72 10.93 1.398 ;
      RECT 10.92 0.722 10.925 1.433 ;
      RECT 10.915 0.724 10.92 1.515 ;
      RECT 10.91 0.726 10.915 1.603 ;
      RECT 10.9 0.728 10.91 1.685 ;
      RECT 10.885 0.742 10.9 1.69 ;
      RECT 10.85 0.787 10.885 1.69 ;
      RECT 10.84 0.827 10.85 1.69 ;
      RECT 10.825 0.855 10.84 1.69 ;
      RECT 10.82 0.872 10.825 1.69 ;
      RECT 10.815 0.88 10.82 1.69 ;
      RECT 10.805 0.895 10.81 1.69 ;
      RECT 10.8 0.902 10.805 1.69 ;
      RECT 10.79 0.922 10.8 1.69 ;
      RECT 10.785 0.935 10.79 1.69 ;
      RECT 10.75 0.94 10.755 1.275 ;
      RECT 10.735 1.33 10.755 1.69 ;
      RECT 10.735 0.94 10.745 1.248 ;
      RECT 10.73 1.37 10.735 1.69 ;
      RECT 10.68 0.94 10.73 1.243 ;
      RECT 10.725 1.407 10.73 1.69 ;
      RECT 10.715 1.43 10.725 1.69 ;
      RECT 10.71 1.475 10.715 1.69 ;
      RECT 10.7 1.485 10.71 1.683 ;
      RECT 10.626 0.94 10.68 1.237 ;
      RECT 10.54 0.94 10.626 1.23 ;
      RECT 10.491 0.987 10.54 1.223 ;
      RECT 10.405 0.995 10.491 1.216 ;
      RECT 10.39 0.992 10.405 1.211 ;
      RECT 10.376 0.985 10.39 1.21 ;
      RECT 10.29 0.985 10.376 1.205 ;
      RECT 10.195 0.99 10.205 1.19 ;
      RECT 9.785 0.42 9.8 0.82 ;
      RECT 9.98 0.42 9.985 0.68 ;
      RECT 9.725 0.42 9.77 0.68 ;
      RECT 10.18 1.725 10.185 1.93 ;
      RECT 10.175 1.715 10.18 1.935 ;
      RECT 10.17 1.702 10.175 1.94 ;
      RECT 10.165 1.682 10.17 1.94 ;
      RECT 10.14 1.635 10.165 1.94 ;
      RECT 10.105 1.55 10.14 1.94 ;
      RECT 10.1 1.487 10.105 1.94 ;
      RECT 10.095 1.472 10.1 1.94 ;
      RECT 10.08 1.432 10.095 1.94 ;
      RECT 10.075 1.407 10.08 1.94 ;
      RECT 10.065 1.39 10.075 1.94 ;
      RECT 10.03 1.312 10.065 1.94 ;
      RECT 10.025 1.255 10.03 1.94 ;
      RECT 10.02 1.242 10.025 1.94 ;
      RECT 10.01 1.22 10.02 1.94 ;
      RECT 10 1.185 10.01 1.94 ;
      RECT 9.99 1.155 10 1.94 ;
      RECT 9.98 1.07 9.99 1.583 ;
      RECT 9.987 1.715 9.99 1.94 ;
      RECT 9.985 1.725 9.987 1.94 ;
      RECT 9.975 1.735 9.985 1.935 ;
      RECT 9.97 0.42 9.98 0.815 ;
      RECT 9.975 0.947 9.98 1.558 ;
      RECT 9.97 0.845 9.975 1.541 ;
      RECT 9.96 0.42 9.97 1.517 ;
      RECT 9.955 0.42 9.96 1.488 ;
      RECT 9.95 0.42 9.955 1.478 ;
      RECT 9.93 0.42 9.95 1.44 ;
      RECT 9.925 0.42 9.93 1.398 ;
      RECT 9.92 0.42 9.925 1.378 ;
      RECT 9.89 0.42 9.92 1.328 ;
      RECT 9.88 0.42 9.89 1.275 ;
      RECT 9.875 0.42 9.88 1.248 ;
      RECT 9.87 0.42 9.875 1.233 ;
      RECT 9.86 0.42 9.87 1.21 ;
      RECT 9.85 0.42 9.86 1.185 ;
      RECT 9.845 0.42 9.85 1.125 ;
      RECT 9.835 0.42 9.845 1.063 ;
      RECT 9.83 0.42 9.835 0.983 ;
      RECT 9.825 0.42 9.83 0.948 ;
      RECT 9.82 0.42 9.825 0.923 ;
      RECT 9.815 0.42 9.82 0.908 ;
      RECT 9.81 0.42 9.815 0.878 ;
      RECT 9.805 0.42 9.81 0.855 ;
      RECT 9.8 0.42 9.805 0.828 ;
      RECT 9.77 0.42 9.785 0.815 ;
      RECT 8.925 1.955 9.11 2.165 ;
      RECT 8.915 1.96 9.125 2.158 ;
      RECT 8.915 1.96 9.145 2.13 ;
      RECT 8.915 1.96 9.16 2.109 ;
      RECT 8.915 1.96 9.175 2.107 ;
      RECT 8.915 1.96 9.185 2.106 ;
      RECT 8.915 1.96 9.215 2.103 ;
      RECT 9.565 1.805 9.825 2.065 ;
      RECT 9.525 1.852 9.825 2.048 ;
      RECT 9.516 1.86 9.525 2.051 ;
      RECT 9.11 1.953 9.825 2.048 ;
      RECT 9.43 1.878 9.516 2.058 ;
      RECT 9.125 1.95 9.825 2.048 ;
      RECT 9.371 1.9 9.43 2.07 ;
      RECT 9.145 1.946 9.825 2.048 ;
      RECT 9.285 1.912 9.371 2.081 ;
      RECT 9.16 1.942 9.825 2.048 ;
      RECT 9.23 1.925 9.285 2.093 ;
      RECT 9.175 1.94 9.825 2.048 ;
      RECT 9.215 1.931 9.23 2.099 ;
      RECT 9.185 1.936 9.825 2.048 ;
      RECT 9.33 1.46 9.59 1.72 ;
      RECT 9.33 1.48 9.7 1.69 ;
      RECT 9.33 1.485 9.71 1.685 ;
      RECT 9.521 0.899 9.6 1.13 ;
      RECT 9.435 0.902 9.65 1.125 ;
      RECT 9.43 0.902 9.65 1.12 ;
      RECT 9.43 0.907 9.66 1.118 ;
      RECT 9.405 0.907 9.66 1.115 ;
      RECT 9.405 0.915 9.67 1.113 ;
      RECT 9.285 0.85 9.545 1.11 ;
      RECT 9.285 0.897 9.595 1.11 ;
      RECT 8.54 1.47 8.545 1.73 ;
      RECT 8.37 1.24 8.375 1.73 ;
      RECT 8.255 1.48 8.26 1.705 ;
      RECT 8.965 0.575 8.97 0.785 ;
      RECT 8.97 0.58 8.985 0.78 ;
      RECT 8.905 0.575 8.965 0.793 ;
      RECT 8.89 0.575 8.905 0.803 ;
      RECT 8.84 0.575 8.89 0.82 ;
      RECT 8.82 0.575 8.84 0.843 ;
      RECT 8.805 0.575 8.82 0.855 ;
      RECT 8.785 0.575 8.805 0.865 ;
      RECT 8.775 0.58 8.785 0.874 ;
      RECT 8.77 0.59 8.775 0.879 ;
      RECT 8.765 0.602 8.77 0.883 ;
      RECT 8.755 0.625 8.765 0.888 ;
      RECT 8.75 0.64 8.755 0.892 ;
      RECT 8.745 0.657 8.75 0.895 ;
      RECT 8.74 0.665 8.745 0.898 ;
      RECT 8.73 0.67 8.74 0.902 ;
      RECT 8.725 0.677 8.73 0.907 ;
      RECT 8.715 0.682 8.725 0.911 ;
      RECT 8.69 0.694 8.715 0.922 ;
      RECT 8.67 0.711 8.69 0.938 ;
      RECT 8.645 0.728 8.67 0.96 ;
      RECT 8.61 0.751 8.645 1.018 ;
      RECT 8.59 0.773 8.61 1.08 ;
      RECT 8.585 0.783 8.59 1.115 ;
      RECT 8.575 0.79 8.585 1.153 ;
      RECT 8.57 0.797 8.575 1.173 ;
      RECT 8.565 0.808 8.57 1.21 ;
      RECT 8.56 0.816 8.565 1.275 ;
      RECT 8.55 0.827 8.56 1.328 ;
      RECT 8.545 0.845 8.55 1.398 ;
      RECT 8.54 0.855 8.545 1.435 ;
      RECT 8.535 0.865 8.54 1.73 ;
      RECT 8.53 0.877 8.535 1.73 ;
      RECT 8.525 0.887 8.53 1.73 ;
      RECT 8.515 0.897 8.525 1.73 ;
      RECT 8.505 0.92 8.515 1.73 ;
      RECT 8.49 0.955 8.505 1.73 ;
      RECT 8.45 1.017 8.49 1.73 ;
      RECT 8.445 1.07 8.45 1.73 ;
      RECT 8.42 1.105 8.445 1.73 ;
      RECT 8.405 1.15 8.42 1.73 ;
      RECT 8.4 1.172 8.405 1.73 ;
      RECT 8.39 1.185 8.4 1.73 ;
      RECT 8.38 1.21 8.39 1.73 ;
      RECT 8.375 1.232 8.38 1.73 ;
      RECT 8.35 1.27 8.37 1.73 ;
      RECT 8.31 1.327 8.35 1.73 ;
      RECT 8.305 1.377 8.31 1.73 ;
      RECT 8.3 1.395 8.305 1.73 ;
      RECT 8.295 1.407 8.3 1.73 ;
      RECT 8.285 1.425 8.295 1.73 ;
      RECT 8.275 1.445 8.285 1.705 ;
      RECT 8.27 1.462 8.275 1.705 ;
      RECT 8.26 1.475 8.27 1.705 ;
      RECT 8.23 1.485 8.255 1.705 ;
      RECT 8.22 1.492 8.23 1.705 ;
      RECT 8.205 1.502 8.22 1.7 ;
      RECT 7.165 1.415 7.485 1.675 ;
      RECT 7.03 1.46 7.485 1.63 ;
      RECT 0.115 1.78 0.405 2.02 ;
      RECT 0.175 1.595 0.35 2.02 ;
      RECT 0.18 1.135 0.35 2.02 ;
      RECT 0.18 1.135 6.76 1.305 ;
      RECT 6.59 0.66 6.76 1.305 ;
      RECT 6.31 0.475 6.63 0.735 ;
      RECT 6.31 0.505 6.71 0.735 ;
      RECT 3.975 1.515 4.27 1.805 ;
      RECT 3.945 1.515 4.27 1.775 ;
      RECT 0 -0.24 141.925 0.24 ;
      RECT 138.695 0.845 139.025 1.115 ;
      RECT 134.625 0.545 134.945 0.805 ;
      RECT 130.085 0.485 130.405 0.745 ;
      RECT 107.03 0.545 107.35 0.805 ;
      RECT 102.49 0.485 102.81 0.745 ;
      RECT 79.435 0.545 79.755 0.805 ;
      RECT 74.895 0.485 75.215 0.745 ;
      RECT 51.84 0.545 52.16 0.805 ;
      RECT 47.3 0.485 47.62 0.745 ;
      RECT 24.245 0.545 24.565 0.805 ;
      RECT 19.705 0.485 20.025 0.745 ;
      RECT 1.95 0.65 2.27 0.91 ;
    LAYER mcon ;
      RECT 141.61 -0.085 141.78 0.085 ;
      RECT 141.61 2.635 141.78 2.805 ;
      RECT 141.15 -0.085 141.32 0.085 ;
      RECT 141.15 2.635 141.32 2.805 ;
      RECT 140.69 -0.085 140.86 0.085 ;
      RECT 140.69 2.635 140.86 2.805 ;
      RECT 140.23 -0.085 140.4 0.085 ;
      RECT 140.23 2.635 140.4 2.805 ;
      RECT 139.77 -0.085 139.94 0.085 ;
      RECT 139.77 2.635 139.94 2.805 ;
      RECT 139.565 1.1 139.735 1.27 ;
      RECT 139.31 -0.085 139.48 0.085 ;
      RECT 139.31 2.635 139.48 2.805 ;
      RECT 138.85 -0.085 139.02 0.085 ;
      RECT 138.85 2.635 139.02 2.805 ;
      RECT 138.795 0.895 138.965 1.065 ;
      RECT 138.39 -0.085 138.56 0.085 ;
      RECT 138.39 2.635 138.56 2.805 ;
      RECT 137.93 -0.085 138.1 0.085 ;
      RECT 137.93 2.635 138.1 2.805 ;
      RECT 137.47 -0.085 137.64 0.085 ;
      RECT 137.47 2.635 137.64 2.805 ;
      RECT 137.01 -0.085 137.18 0.085 ;
      RECT 137.01 2.635 137.18 2.805 ;
      RECT 136.805 1.105 136.975 1.275 ;
      RECT 136.55 -0.085 136.72 0.085 ;
      RECT 136.55 2.635 136.72 2.805 ;
      RECT 136.09 -0.085 136.26 0.085 ;
      RECT 136.09 2.635 136.26 2.805 ;
      RECT 135.63 -0.085 135.8 0.085 ;
      RECT 135.63 2.635 135.8 2.805 ;
      RECT 135.56 1.46 135.73 1.63 ;
      RECT 135.17 -0.085 135.34 0.085 ;
      RECT 135.17 2.635 135.34 2.805 ;
      RECT 134.71 -0.085 134.88 0.085 ;
      RECT 134.71 2.635 134.88 2.805 ;
      RECT 134.7 0.575 134.87 0.745 ;
      RECT 134.255 0.455 134.425 0.625 ;
      RECT 134.25 -0.085 134.42 0.085 ;
      RECT 134.25 2.635 134.42 2.805 ;
      RECT 133.79 -0.085 133.96 0.085 ;
      RECT 133.79 2.635 133.96 2.805 ;
      RECT 133.33 -0.085 133.5 0.085 ;
      RECT 133.33 2.635 133.5 2.805 ;
      RECT 132.87 -0.085 133.04 0.085 ;
      RECT 132.87 2.635 133.04 2.805 ;
      RECT 132.41 -0.085 132.58 0.085 ;
      RECT 132.41 2.635 132.58 2.805 ;
      RECT 132.355 1.075 132.525 1.245 ;
      RECT 131.955 -0.085 132.125 0.085 ;
      RECT 131.955 2.635 132.125 2.805 ;
      RECT 131.495 -0.085 131.665 0.085 ;
      RECT 131.495 2.635 131.665 2.805 ;
      RECT 131.425 1.46 131.595 1.63 ;
      RECT 131.035 -0.085 131.205 0.085 ;
      RECT 131.035 2.635 131.205 2.805 ;
      RECT 130.575 -0.085 130.745 0.085 ;
      RECT 130.575 2.635 130.745 2.805 ;
      RECT 130.16 0.515 130.33 0.685 ;
      RECT 130.115 -0.085 130.285 0.085 ;
      RECT 130.115 2.635 130.285 2.805 ;
      RECT 129.745 1.24 129.915 1.41 ;
      RECT 129.655 -0.085 129.825 0.085 ;
      RECT 129.655 2.635 129.825 2.805 ;
      RECT 129.195 -0.085 129.365 0.085 ;
      RECT 129.195 2.635 129.365 2.805 ;
      RECT 128.735 -0.085 128.905 0.085 ;
      RECT 128.735 2.635 128.905 2.805 ;
      RECT 128.275 -0.085 128.445 0.085 ;
      RECT 128.275 2.635 128.445 2.805 ;
      RECT 128.22 1.915 128.39 2.085 ;
      RECT 127.815 -0.085 127.985 0.085 ;
      RECT 127.815 2.635 127.985 2.805 ;
      RECT 127.445 1.375 127.615 1.545 ;
      RECT 127.355 -0.085 127.525 0.085 ;
      RECT 127.355 2.635 127.525 2.805 ;
      RECT 127.125 0.545 127.295 0.715 ;
      RECT 126.98 0.985 127.15 1.155 ;
      RECT 126.895 -0.085 127.065 0.085 ;
      RECT 126.895 2.635 127.065 2.805 ;
      RECT 126.435 -0.085 126.605 0.085 ;
      RECT 126.435 2.635 126.605 2.805 ;
      RECT 126.37 1.025 126.54 1.195 ;
      RECT 126.025 0.66 126.195 0.83 ;
      RECT 126.015 2.02 126.185 2.19 ;
      RECT 125.975 -0.085 126.145 0.085 ;
      RECT 125.975 2.635 126.145 2.805 ;
      RECT 125.6 1.26 125.77 1.43 ;
      RECT 125.515 -0.085 125.685 0.085 ;
      RECT 125.515 2.635 125.685 2.805 ;
      RECT 125.25 0.735 125.42 0.905 ;
      RECT 125.07 2.05 125.24 2.22 ;
      RECT 125.055 -0.085 125.225 0.085 ;
      RECT 125.055 2.635 125.225 2.805 ;
      RECT 124.79 1.365 124.96 1.535 ;
      RECT 124.595 -0.085 124.765 0.085 ;
      RECT 124.595 2.635 124.765 2.805 ;
      RECT 124.47 0.99 124.64 1.16 ;
      RECT 124.135 -0.085 124.305 0.085 ;
      RECT 124.135 2.635 124.305 2.805 ;
      RECT 123.78 0.47 123.95 0.64 ;
      RECT 123.705 0.94 123.875 1.11 ;
      RECT 123.675 -0.085 123.845 0.085 ;
      RECT 123.675 2.635 123.845 2.805 ;
      RECT 123.215 -0.085 123.385 0.085 ;
      RECT 123.215 2.635 123.385 2.805 ;
      RECT 122.855 0.665 123.025 0.835 ;
      RECT 122.755 -0.085 122.925 0.085 ;
      RECT 122.755 2.635 122.925 2.805 ;
      RECT 122.515 1.86 122.685 2.03 ;
      RECT 122.48 1.195 122.65 1.365 ;
      RECT 122.295 -0.085 122.465 0.085 ;
      RECT 122.295 2.635 122.465 2.805 ;
      RECT 121.87 1.05 122.04 1.22 ;
      RECT 121.835 -0.085 122.005 0.085 ;
      RECT 121.835 2.635 122.005 2.805 ;
      RECT 121.8 1.75 121.97 1.92 ;
      RECT 121.74 0.585 121.91 0.755 ;
      RECT 121.375 -0.085 121.545 0.085 ;
      RECT 121.375 2.635 121.545 2.805 ;
      RECT 121.1 1.5 121.27 1.67 ;
      RECT 120.915 -0.085 121.085 0.085 ;
      RECT 120.915 2.635 121.085 2.805 ;
      RECT 120.595 1.005 120.765 1.175 ;
      RECT 120.455 -0.085 120.625 0.085 ;
      RECT 120.455 2.635 120.625 2.805 ;
      RECT 120.375 1.75 120.545 1.92 ;
      RECT 120.17 0.63 120.34 0.8 ;
      RECT 119.995 -0.085 120.165 0.085 ;
      RECT 119.995 2.635 120.165 2.805 ;
      RECT 119.9 1.5 120.07 1.67 ;
      RECT 119.86 0.93 120.03 1.1 ;
      RECT 119.535 -0.085 119.705 0.085 ;
      RECT 119.535 2.635 119.705 2.805 ;
      RECT 119.315 1.975 119.485 2.145 ;
      RECT 119.175 0.595 119.345 0.765 ;
      RECT 119.075 -0.085 119.245 0.085 ;
      RECT 119.075 2.635 119.245 2.805 ;
      RECT 118.615 -0.085 118.785 0.085 ;
      RECT 118.615 2.635 118.785 2.805 ;
      RECT 118.605 1.515 118.775 1.685 ;
      RECT 118.155 -0.085 118.325 0.085 ;
      RECT 118.155 2.635 118.325 2.805 ;
      RECT 117.695 -0.085 117.865 0.085 ;
      RECT 117.695 2.635 117.865 2.805 ;
      RECT 117.625 1.46 117.795 1.63 ;
      RECT 117.235 -0.085 117.405 0.085 ;
      RECT 117.235 2.635 117.405 2.805 ;
      RECT 116.775 -0.085 116.945 0.085 ;
      RECT 116.775 2.635 116.945 2.805 ;
      RECT 116.765 0.505 116.935 0.675 ;
      RECT 116.315 -0.085 116.485 0.085 ;
      RECT 116.315 2.635 116.485 2.805 ;
      RECT 115.855 -0.085 116.025 0.085 ;
      RECT 115.855 2.635 116.025 2.805 ;
      RECT 115.395 -0.085 115.565 0.085 ;
      RECT 115.395 2.635 115.565 2.805 ;
      RECT 114.935 -0.085 115.105 0.085 ;
      RECT 114.935 2.635 115.105 2.805 ;
      RECT 114.475 -0.085 114.645 0.085 ;
      RECT 114.475 2.635 114.645 2.805 ;
      RECT 114.42 1.575 114.59 1.745 ;
      RECT 114.015 -0.085 114.185 0.085 ;
      RECT 114.015 2.635 114.185 2.805 ;
      RECT 113.555 -0.085 113.725 0.085 ;
      RECT 113.555 2.635 113.725 2.805 ;
      RECT 113.095 -0.085 113.265 0.085 ;
      RECT 113.095 2.635 113.265 2.805 ;
      RECT 112.635 -0.085 112.805 0.085 ;
      RECT 112.635 2.635 112.805 2.805 ;
      RECT 112.175 -0.085 112.345 0.085 ;
      RECT 112.175 2.635 112.345 2.805 ;
      RECT 111.97 1.1 112.14 1.27 ;
      RECT 111.715 -0.085 111.885 0.085 ;
      RECT 111.715 2.635 111.885 2.805 ;
      RECT 111.255 -0.085 111.425 0.085 ;
      RECT 111.255 2.635 111.425 2.805 ;
      RECT 111.2 1.555 111.37 1.725 ;
      RECT 110.795 -0.085 110.965 0.085 ;
      RECT 110.795 2.635 110.965 2.805 ;
      RECT 110.335 -0.085 110.505 0.085 ;
      RECT 110.335 2.635 110.505 2.805 ;
      RECT 109.875 -0.085 110.045 0.085 ;
      RECT 109.875 2.635 110.045 2.805 ;
      RECT 109.415 -0.085 109.585 0.085 ;
      RECT 109.415 2.635 109.585 2.805 ;
      RECT 109.21 1.105 109.38 1.275 ;
      RECT 108.955 -0.085 109.125 0.085 ;
      RECT 108.955 2.635 109.125 2.805 ;
      RECT 108.495 -0.085 108.665 0.085 ;
      RECT 108.495 2.635 108.665 2.805 ;
      RECT 108.035 -0.085 108.205 0.085 ;
      RECT 108.035 2.635 108.205 2.805 ;
      RECT 107.965 1.46 108.135 1.63 ;
      RECT 107.575 -0.085 107.745 0.085 ;
      RECT 107.575 2.635 107.745 2.805 ;
      RECT 107.115 -0.085 107.285 0.085 ;
      RECT 107.115 2.635 107.285 2.805 ;
      RECT 107.105 0.575 107.275 0.745 ;
      RECT 106.66 0.455 106.83 0.625 ;
      RECT 106.655 -0.085 106.825 0.085 ;
      RECT 106.655 2.635 106.825 2.805 ;
      RECT 106.195 -0.085 106.365 0.085 ;
      RECT 106.195 2.635 106.365 2.805 ;
      RECT 105.735 -0.085 105.905 0.085 ;
      RECT 105.735 2.635 105.905 2.805 ;
      RECT 105.275 -0.085 105.445 0.085 ;
      RECT 105.275 2.635 105.445 2.805 ;
      RECT 104.815 -0.085 104.985 0.085 ;
      RECT 104.815 2.635 104.985 2.805 ;
      RECT 104.76 1.075 104.93 1.245 ;
      RECT 104.36 -0.085 104.53 0.085 ;
      RECT 104.36 2.635 104.53 2.805 ;
      RECT 103.9 -0.085 104.07 0.085 ;
      RECT 103.9 2.635 104.07 2.805 ;
      RECT 103.83 1.46 104 1.63 ;
      RECT 103.44 -0.085 103.61 0.085 ;
      RECT 103.44 2.635 103.61 2.805 ;
      RECT 102.98 -0.085 103.15 0.085 ;
      RECT 102.98 2.635 103.15 2.805 ;
      RECT 102.565 0.515 102.735 0.685 ;
      RECT 102.52 -0.085 102.69 0.085 ;
      RECT 102.52 2.635 102.69 2.805 ;
      RECT 102.15 1.24 102.32 1.41 ;
      RECT 102.06 -0.085 102.23 0.085 ;
      RECT 102.06 2.635 102.23 2.805 ;
      RECT 101.6 -0.085 101.77 0.085 ;
      RECT 101.6 2.635 101.77 2.805 ;
      RECT 101.14 -0.085 101.31 0.085 ;
      RECT 101.14 2.635 101.31 2.805 ;
      RECT 100.68 -0.085 100.85 0.085 ;
      RECT 100.68 2.635 100.85 2.805 ;
      RECT 100.625 1.915 100.795 2.085 ;
      RECT 100.22 -0.085 100.39 0.085 ;
      RECT 100.22 2.635 100.39 2.805 ;
      RECT 99.85 1.375 100.02 1.545 ;
      RECT 99.76 -0.085 99.93 0.085 ;
      RECT 99.76 2.635 99.93 2.805 ;
      RECT 99.53 0.545 99.7 0.715 ;
      RECT 99.385 0.985 99.555 1.155 ;
      RECT 99.3 -0.085 99.47 0.085 ;
      RECT 99.3 2.635 99.47 2.805 ;
      RECT 98.84 -0.085 99.01 0.085 ;
      RECT 98.84 2.635 99.01 2.805 ;
      RECT 98.775 1.025 98.945 1.195 ;
      RECT 98.43 0.66 98.6 0.83 ;
      RECT 98.42 2.02 98.59 2.19 ;
      RECT 98.38 -0.085 98.55 0.085 ;
      RECT 98.38 2.635 98.55 2.805 ;
      RECT 98.005 1.26 98.175 1.43 ;
      RECT 97.92 -0.085 98.09 0.085 ;
      RECT 97.92 2.635 98.09 2.805 ;
      RECT 97.655 0.735 97.825 0.905 ;
      RECT 97.475 2.05 97.645 2.22 ;
      RECT 97.46 -0.085 97.63 0.085 ;
      RECT 97.46 2.635 97.63 2.805 ;
      RECT 97.195 1.365 97.365 1.535 ;
      RECT 97 -0.085 97.17 0.085 ;
      RECT 97 2.635 97.17 2.805 ;
      RECT 96.875 0.99 97.045 1.16 ;
      RECT 96.54 -0.085 96.71 0.085 ;
      RECT 96.54 2.635 96.71 2.805 ;
      RECT 96.185 0.47 96.355 0.64 ;
      RECT 96.11 0.94 96.28 1.11 ;
      RECT 96.08 -0.085 96.25 0.085 ;
      RECT 96.08 2.635 96.25 2.805 ;
      RECT 95.62 -0.085 95.79 0.085 ;
      RECT 95.62 2.635 95.79 2.805 ;
      RECT 95.26 0.665 95.43 0.835 ;
      RECT 95.16 -0.085 95.33 0.085 ;
      RECT 95.16 2.635 95.33 2.805 ;
      RECT 94.92 1.86 95.09 2.03 ;
      RECT 94.885 1.195 95.055 1.365 ;
      RECT 94.7 -0.085 94.87 0.085 ;
      RECT 94.7 2.635 94.87 2.805 ;
      RECT 94.275 1.05 94.445 1.22 ;
      RECT 94.24 -0.085 94.41 0.085 ;
      RECT 94.24 2.635 94.41 2.805 ;
      RECT 94.205 1.75 94.375 1.92 ;
      RECT 94.145 0.585 94.315 0.755 ;
      RECT 93.78 -0.085 93.95 0.085 ;
      RECT 93.78 2.635 93.95 2.805 ;
      RECT 93.505 1.5 93.675 1.67 ;
      RECT 93.32 -0.085 93.49 0.085 ;
      RECT 93.32 2.635 93.49 2.805 ;
      RECT 93 1.005 93.17 1.175 ;
      RECT 92.86 -0.085 93.03 0.085 ;
      RECT 92.86 2.635 93.03 2.805 ;
      RECT 92.78 1.75 92.95 1.92 ;
      RECT 92.575 0.63 92.745 0.8 ;
      RECT 92.4 -0.085 92.57 0.085 ;
      RECT 92.4 2.635 92.57 2.805 ;
      RECT 92.305 1.5 92.475 1.67 ;
      RECT 92.265 0.93 92.435 1.1 ;
      RECT 91.94 -0.085 92.11 0.085 ;
      RECT 91.94 2.635 92.11 2.805 ;
      RECT 91.72 1.975 91.89 2.145 ;
      RECT 91.58 0.595 91.75 0.765 ;
      RECT 91.48 -0.085 91.65 0.085 ;
      RECT 91.48 2.635 91.65 2.805 ;
      RECT 91.02 -0.085 91.19 0.085 ;
      RECT 91.02 2.635 91.19 2.805 ;
      RECT 91.01 1.515 91.18 1.685 ;
      RECT 90.56 -0.085 90.73 0.085 ;
      RECT 90.56 2.635 90.73 2.805 ;
      RECT 90.1 -0.085 90.27 0.085 ;
      RECT 90.1 2.635 90.27 2.805 ;
      RECT 90.03 1.46 90.2 1.63 ;
      RECT 89.64 -0.085 89.81 0.085 ;
      RECT 89.64 2.635 89.81 2.805 ;
      RECT 89.18 -0.085 89.35 0.085 ;
      RECT 89.18 2.635 89.35 2.805 ;
      RECT 89.17 0.505 89.34 0.675 ;
      RECT 88.72 -0.085 88.89 0.085 ;
      RECT 88.72 2.635 88.89 2.805 ;
      RECT 88.26 -0.085 88.43 0.085 ;
      RECT 88.26 2.635 88.43 2.805 ;
      RECT 87.8 -0.085 87.97 0.085 ;
      RECT 87.8 2.635 87.97 2.805 ;
      RECT 87.34 -0.085 87.51 0.085 ;
      RECT 87.34 2.635 87.51 2.805 ;
      RECT 86.88 -0.085 87.05 0.085 ;
      RECT 86.88 2.635 87.05 2.805 ;
      RECT 86.825 1.575 86.995 1.745 ;
      RECT 86.42 -0.085 86.59 0.085 ;
      RECT 86.42 2.635 86.59 2.805 ;
      RECT 85.96 -0.085 86.13 0.085 ;
      RECT 85.96 2.635 86.13 2.805 ;
      RECT 85.5 -0.085 85.67 0.085 ;
      RECT 85.5 2.635 85.67 2.805 ;
      RECT 85.04 -0.085 85.21 0.085 ;
      RECT 85.04 2.635 85.21 2.805 ;
      RECT 84.58 -0.085 84.75 0.085 ;
      RECT 84.58 2.635 84.75 2.805 ;
      RECT 84.375 1.1 84.545 1.27 ;
      RECT 84.12 -0.085 84.29 0.085 ;
      RECT 84.12 2.635 84.29 2.805 ;
      RECT 83.66 -0.085 83.83 0.085 ;
      RECT 83.66 2.635 83.83 2.805 ;
      RECT 83.605 1.555 83.775 1.725 ;
      RECT 83.2 -0.085 83.37 0.085 ;
      RECT 83.2 2.635 83.37 2.805 ;
      RECT 82.74 -0.085 82.91 0.085 ;
      RECT 82.74 2.635 82.91 2.805 ;
      RECT 82.28 -0.085 82.45 0.085 ;
      RECT 82.28 2.635 82.45 2.805 ;
      RECT 81.82 -0.085 81.99 0.085 ;
      RECT 81.82 2.635 81.99 2.805 ;
      RECT 81.615 1.105 81.785 1.275 ;
      RECT 81.36 -0.085 81.53 0.085 ;
      RECT 81.36 2.635 81.53 2.805 ;
      RECT 80.9 -0.085 81.07 0.085 ;
      RECT 80.9 2.635 81.07 2.805 ;
      RECT 80.44 -0.085 80.61 0.085 ;
      RECT 80.44 2.635 80.61 2.805 ;
      RECT 80.37 1.46 80.54 1.63 ;
      RECT 79.98 -0.085 80.15 0.085 ;
      RECT 79.98 2.635 80.15 2.805 ;
      RECT 79.52 -0.085 79.69 0.085 ;
      RECT 79.52 2.635 79.69 2.805 ;
      RECT 79.51 0.575 79.68 0.745 ;
      RECT 79.065 0.455 79.235 0.625 ;
      RECT 79.06 -0.085 79.23 0.085 ;
      RECT 79.06 2.635 79.23 2.805 ;
      RECT 78.6 -0.085 78.77 0.085 ;
      RECT 78.6 2.635 78.77 2.805 ;
      RECT 78.14 -0.085 78.31 0.085 ;
      RECT 78.14 2.635 78.31 2.805 ;
      RECT 77.68 -0.085 77.85 0.085 ;
      RECT 77.68 2.635 77.85 2.805 ;
      RECT 77.22 -0.085 77.39 0.085 ;
      RECT 77.22 2.635 77.39 2.805 ;
      RECT 77.165 1.075 77.335 1.245 ;
      RECT 76.765 -0.085 76.935 0.085 ;
      RECT 76.765 2.635 76.935 2.805 ;
      RECT 76.305 -0.085 76.475 0.085 ;
      RECT 76.305 2.635 76.475 2.805 ;
      RECT 76.235 1.46 76.405 1.63 ;
      RECT 75.845 -0.085 76.015 0.085 ;
      RECT 75.845 2.635 76.015 2.805 ;
      RECT 75.385 -0.085 75.555 0.085 ;
      RECT 75.385 2.635 75.555 2.805 ;
      RECT 74.97 0.515 75.14 0.685 ;
      RECT 74.925 -0.085 75.095 0.085 ;
      RECT 74.925 2.635 75.095 2.805 ;
      RECT 74.555 1.24 74.725 1.41 ;
      RECT 74.465 -0.085 74.635 0.085 ;
      RECT 74.465 2.635 74.635 2.805 ;
      RECT 74.005 -0.085 74.175 0.085 ;
      RECT 74.005 2.635 74.175 2.805 ;
      RECT 73.545 -0.085 73.715 0.085 ;
      RECT 73.545 2.635 73.715 2.805 ;
      RECT 73.085 -0.085 73.255 0.085 ;
      RECT 73.085 2.635 73.255 2.805 ;
      RECT 73.03 1.915 73.2 2.085 ;
      RECT 72.625 -0.085 72.795 0.085 ;
      RECT 72.625 2.635 72.795 2.805 ;
      RECT 72.255 1.375 72.425 1.545 ;
      RECT 72.165 -0.085 72.335 0.085 ;
      RECT 72.165 2.635 72.335 2.805 ;
      RECT 71.935 0.545 72.105 0.715 ;
      RECT 71.79 0.985 71.96 1.155 ;
      RECT 71.705 -0.085 71.875 0.085 ;
      RECT 71.705 2.635 71.875 2.805 ;
      RECT 71.245 -0.085 71.415 0.085 ;
      RECT 71.245 2.635 71.415 2.805 ;
      RECT 71.18 1.025 71.35 1.195 ;
      RECT 70.835 0.66 71.005 0.83 ;
      RECT 70.825 2.02 70.995 2.19 ;
      RECT 70.785 -0.085 70.955 0.085 ;
      RECT 70.785 2.635 70.955 2.805 ;
      RECT 70.41 1.26 70.58 1.43 ;
      RECT 70.325 -0.085 70.495 0.085 ;
      RECT 70.325 2.635 70.495 2.805 ;
      RECT 70.06 0.735 70.23 0.905 ;
      RECT 69.88 2.05 70.05 2.22 ;
      RECT 69.865 -0.085 70.035 0.085 ;
      RECT 69.865 2.635 70.035 2.805 ;
      RECT 69.6 1.365 69.77 1.535 ;
      RECT 69.405 -0.085 69.575 0.085 ;
      RECT 69.405 2.635 69.575 2.805 ;
      RECT 69.28 0.99 69.45 1.16 ;
      RECT 68.945 -0.085 69.115 0.085 ;
      RECT 68.945 2.635 69.115 2.805 ;
      RECT 68.59 0.47 68.76 0.64 ;
      RECT 68.515 0.94 68.685 1.11 ;
      RECT 68.485 -0.085 68.655 0.085 ;
      RECT 68.485 2.635 68.655 2.805 ;
      RECT 68.025 -0.085 68.195 0.085 ;
      RECT 68.025 2.635 68.195 2.805 ;
      RECT 67.665 0.665 67.835 0.835 ;
      RECT 67.565 -0.085 67.735 0.085 ;
      RECT 67.565 2.635 67.735 2.805 ;
      RECT 67.325 1.86 67.495 2.03 ;
      RECT 67.29 1.195 67.46 1.365 ;
      RECT 67.105 -0.085 67.275 0.085 ;
      RECT 67.105 2.635 67.275 2.805 ;
      RECT 66.68 1.05 66.85 1.22 ;
      RECT 66.645 -0.085 66.815 0.085 ;
      RECT 66.645 2.635 66.815 2.805 ;
      RECT 66.61 1.75 66.78 1.92 ;
      RECT 66.55 0.585 66.72 0.755 ;
      RECT 66.185 -0.085 66.355 0.085 ;
      RECT 66.185 2.635 66.355 2.805 ;
      RECT 65.91 1.5 66.08 1.67 ;
      RECT 65.725 -0.085 65.895 0.085 ;
      RECT 65.725 2.635 65.895 2.805 ;
      RECT 65.405 1.005 65.575 1.175 ;
      RECT 65.265 -0.085 65.435 0.085 ;
      RECT 65.265 2.635 65.435 2.805 ;
      RECT 65.185 1.75 65.355 1.92 ;
      RECT 64.98 0.63 65.15 0.8 ;
      RECT 64.805 -0.085 64.975 0.085 ;
      RECT 64.805 2.635 64.975 2.805 ;
      RECT 64.71 1.5 64.88 1.67 ;
      RECT 64.67 0.93 64.84 1.1 ;
      RECT 64.345 -0.085 64.515 0.085 ;
      RECT 64.345 2.635 64.515 2.805 ;
      RECT 64.125 1.975 64.295 2.145 ;
      RECT 63.985 0.595 64.155 0.765 ;
      RECT 63.885 -0.085 64.055 0.085 ;
      RECT 63.885 2.635 64.055 2.805 ;
      RECT 63.425 -0.085 63.595 0.085 ;
      RECT 63.425 2.635 63.595 2.805 ;
      RECT 63.415 1.515 63.585 1.685 ;
      RECT 62.965 -0.085 63.135 0.085 ;
      RECT 62.965 2.635 63.135 2.805 ;
      RECT 62.505 -0.085 62.675 0.085 ;
      RECT 62.505 2.635 62.675 2.805 ;
      RECT 62.435 1.46 62.605 1.63 ;
      RECT 62.045 -0.085 62.215 0.085 ;
      RECT 62.045 2.635 62.215 2.805 ;
      RECT 61.585 -0.085 61.755 0.085 ;
      RECT 61.585 2.635 61.755 2.805 ;
      RECT 61.575 0.505 61.745 0.675 ;
      RECT 61.125 -0.085 61.295 0.085 ;
      RECT 61.125 2.635 61.295 2.805 ;
      RECT 60.665 -0.085 60.835 0.085 ;
      RECT 60.665 2.635 60.835 2.805 ;
      RECT 60.205 -0.085 60.375 0.085 ;
      RECT 60.205 2.635 60.375 2.805 ;
      RECT 59.745 -0.085 59.915 0.085 ;
      RECT 59.745 2.635 59.915 2.805 ;
      RECT 59.285 -0.085 59.455 0.085 ;
      RECT 59.285 2.635 59.455 2.805 ;
      RECT 59.23 1.575 59.4 1.745 ;
      RECT 58.825 -0.085 58.995 0.085 ;
      RECT 58.825 2.635 58.995 2.805 ;
      RECT 58.365 -0.085 58.535 0.085 ;
      RECT 58.365 2.635 58.535 2.805 ;
      RECT 57.905 -0.085 58.075 0.085 ;
      RECT 57.905 2.635 58.075 2.805 ;
      RECT 57.445 -0.085 57.615 0.085 ;
      RECT 57.445 2.635 57.615 2.805 ;
      RECT 56.985 -0.085 57.155 0.085 ;
      RECT 56.985 2.635 57.155 2.805 ;
      RECT 56.78 1.1 56.95 1.27 ;
      RECT 56.525 -0.085 56.695 0.085 ;
      RECT 56.525 2.635 56.695 2.805 ;
      RECT 56.065 -0.085 56.235 0.085 ;
      RECT 56.065 2.635 56.235 2.805 ;
      RECT 56.01 1.555 56.18 1.725 ;
      RECT 55.605 -0.085 55.775 0.085 ;
      RECT 55.605 2.635 55.775 2.805 ;
      RECT 55.145 -0.085 55.315 0.085 ;
      RECT 55.145 2.635 55.315 2.805 ;
      RECT 54.685 -0.085 54.855 0.085 ;
      RECT 54.685 2.635 54.855 2.805 ;
      RECT 54.225 -0.085 54.395 0.085 ;
      RECT 54.225 2.635 54.395 2.805 ;
      RECT 54.02 1.105 54.19 1.275 ;
      RECT 53.765 -0.085 53.935 0.085 ;
      RECT 53.765 2.635 53.935 2.805 ;
      RECT 53.305 -0.085 53.475 0.085 ;
      RECT 53.305 2.635 53.475 2.805 ;
      RECT 52.845 -0.085 53.015 0.085 ;
      RECT 52.845 2.635 53.015 2.805 ;
      RECT 52.775 1.46 52.945 1.63 ;
      RECT 52.385 -0.085 52.555 0.085 ;
      RECT 52.385 2.635 52.555 2.805 ;
      RECT 51.925 -0.085 52.095 0.085 ;
      RECT 51.925 2.635 52.095 2.805 ;
      RECT 51.915 0.575 52.085 0.745 ;
      RECT 51.47 0.455 51.64 0.625 ;
      RECT 51.465 -0.085 51.635 0.085 ;
      RECT 51.465 2.635 51.635 2.805 ;
      RECT 51.005 -0.085 51.175 0.085 ;
      RECT 51.005 2.635 51.175 2.805 ;
      RECT 50.545 -0.085 50.715 0.085 ;
      RECT 50.545 2.635 50.715 2.805 ;
      RECT 50.085 -0.085 50.255 0.085 ;
      RECT 50.085 2.635 50.255 2.805 ;
      RECT 49.625 -0.085 49.795 0.085 ;
      RECT 49.625 2.635 49.795 2.805 ;
      RECT 49.57 1.075 49.74 1.245 ;
      RECT 49.17 -0.085 49.34 0.085 ;
      RECT 49.17 2.635 49.34 2.805 ;
      RECT 48.71 -0.085 48.88 0.085 ;
      RECT 48.71 2.635 48.88 2.805 ;
      RECT 48.64 1.46 48.81 1.63 ;
      RECT 48.25 -0.085 48.42 0.085 ;
      RECT 48.25 2.635 48.42 2.805 ;
      RECT 47.79 -0.085 47.96 0.085 ;
      RECT 47.79 2.635 47.96 2.805 ;
      RECT 47.375 0.515 47.545 0.685 ;
      RECT 47.33 -0.085 47.5 0.085 ;
      RECT 47.33 2.635 47.5 2.805 ;
      RECT 46.96 1.24 47.13 1.41 ;
      RECT 46.87 -0.085 47.04 0.085 ;
      RECT 46.87 2.635 47.04 2.805 ;
      RECT 46.41 -0.085 46.58 0.085 ;
      RECT 46.41 2.635 46.58 2.805 ;
      RECT 45.95 -0.085 46.12 0.085 ;
      RECT 45.95 2.635 46.12 2.805 ;
      RECT 45.49 -0.085 45.66 0.085 ;
      RECT 45.49 2.635 45.66 2.805 ;
      RECT 45.435 1.915 45.605 2.085 ;
      RECT 45.03 -0.085 45.2 0.085 ;
      RECT 45.03 2.635 45.2 2.805 ;
      RECT 44.66 1.375 44.83 1.545 ;
      RECT 44.57 -0.085 44.74 0.085 ;
      RECT 44.57 2.635 44.74 2.805 ;
      RECT 44.34 0.545 44.51 0.715 ;
      RECT 44.195 0.985 44.365 1.155 ;
      RECT 44.11 -0.085 44.28 0.085 ;
      RECT 44.11 2.635 44.28 2.805 ;
      RECT 43.65 -0.085 43.82 0.085 ;
      RECT 43.65 2.635 43.82 2.805 ;
      RECT 43.585 1.025 43.755 1.195 ;
      RECT 43.24 0.66 43.41 0.83 ;
      RECT 43.23 2.02 43.4 2.19 ;
      RECT 43.19 -0.085 43.36 0.085 ;
      RECT 43.19 2.635 43.36 2.805 ;
      RECT 42.815 1.26 42.985 1.43 ;
      RECT 42.73 -0.085 42.9 0.085 ;
      RECT 42.73 2.635 42.9 2.805 ;
      RECT 42.465 0.735 42.635 0.905 ;
      RECT 42.285 2.05 42.455 2.22 ;
      RECT 42.27 -0.085 42.44 0.085 ;
      RECT 42.27 2.635 42.44 2.805 ;
      RECT 42.005 1.365 42.175 1.535 ;
      RECT 41.81 -0.085 41.98 0.085 ;
      RECT 41.81 2.635 41.98 2.805 ;
      RECT 41.685 0.99 41.855 1.16 ;
      RECT 41.35 -0.085 41.52 0.085 ;
      RECT 41.35 2.635 41.52 2.805 ;
      RECT 40.995 0.47 41.165 0.64 ;
      RECT 40.92 0.94 41.09 1.11 ;
      RECT 40.89 -0.085 41.06 0.085 ;
      RECT 40.89 2.635 41.06 2.805 ;
      RECT 40.43 -0.085 40.6 0.085 ;
      RECT 40.43 2.635 40.6 2.805 ;
      RECT 40.07 0.665 40.24 0.835 ;
      RECT 39.97 -0.085 40.14 0.085 ;
      RECT 39.97 2.635 40.14 2.805 ;
      RECT 39.73 1.86 39.9 2.03 ;
      RECT 39.695 1.195 39.865 1.365 ;
      RECT 39.51 -0.085 39.68 0.085 ;
      RECT 39.51 2.635 39.68 2.805 ;
      RECT 39.085 1.05 39.255 1.22 ;
      RECT 39.05 -0.085 39.22 0.085 ;
      RECT 39.05 2.635 39.22 2.805 ;
      RECT 39.015 1.75 39.185 1.92 ;
      RECT 38.955 0.585 39.125 0.755 ;
      RECT 38.59 -0.085 38.76 0.085 ;
      RECT 38.59 2.635 38.76 2.805 ;
      RECT 38.315 1.5 38.485 1.67 ;
      RECT 38.13 -0.085 38.3 0.085 ;
      RECT 38.13 2.635 38.3 2.805 ;
      RECT 37.81 1.005 37.98 1.175 ;
      RECT 37.67 -0.085 37.84 0.085 ;
      RECT 37.67 2.635 37.84 2.805 ;
      RECT 37.59 1.75 37.76 1.92 ;
      RECT 37.385 0.63 37.555 0.8 ;
      RECT 37.21 -0.085 37.38 0.085 ;
      RECT 37.21 2.635 37.38 2.805 ;
      RECT 37.115 1.5 37.285 1.67 ;
      RECT 37.075 0.93 37.245 1.1 ;
      RECT 36.75 -0.085 36.92 0.085 ;
      RECT 36.75 2.635 36.92 2.805 ;
      RECT 36.53 1.975 36.7 2.145 ;
      RECT 36.39 0.595 36.56 0.765 ;
      RECT 36.29 -0.085 36.46 0.085 ;
      RECT 36.29 2.635 36.46 2.805 ;
      RECT 35.83 -0.085 36 0.085 ;
      RECT 35.83 2.635 36 2.805 ;
      RECT 35.82 1.515 35.99 1.685 ;
      RECT 35.37 -0.085 35.54 0.085 ;
      RECT 35.37 2.635 35.54 2.805 ;
      RECT 34.91 -0.085 35.08 0.085 ;
      RECT 34.91 2.635 35.08 2.805 ;
      RECT 34.84 1.46 35.01 1.63 ;
      RECT 34.45 -0.085 34.62 0.085 ;
      RECT 34.45 2.635 34.62 2.805 ;
      RECT 33.99 -0.085 34.16 0.085 ;
      RECT 33.99 2.635 34.16 2.805 ;
      RECT 33.98 0.505 34.15 0.675 ;
      RECT 33.53 -0.085 33.7 0.085 ;
      RECT 33.53 2.635 33.7 2.805 ;
      RECT 33.07 -0.085 33.24 0.085 ;
      RECT 33.07 2.635 33.24 2.805 ;
      RECT 32.61 -0.085 32.78 0.085 ;
      RECT 32.61 2.635 32.78 2.805 ;
      RECT 32.15 -0.085 32.32 0.085 ;
      RECT 32.15 2.635 32.32 2.805 ;
      RECT 31.69 -0.085 31.86 0.085 ;
      RECT 31.69 2.635 31.86 2.805 ;
      RECT 31.635 1.575 31.805 1.745 ;
      RECT 31.23 -0.085 31.4 0.085 ;
      RECT 31.23 2.635 31.4 2.805 ;
      RECT 30.77 -0.085 30.94 0.085 ;
      RECT 30.77 2.635 30.94 2.805 ;
      RECT 30.31 -0.085 30.48 0.085 ;
      RECT 30.31 2.635 30.48 2.805 ;
      RECT 29.85 -0.085 30.02 0.085 ;
      RECT 29.85 2.635 30.02 2.805 ;
      RECT 29.39 -0.085 29.56 0.085 ;
      RECT 29.39 2.635 29.56 2.805 ;
      RECT 29.185 1.1 29.355 1.27 ;
      RECT 28.93 -0.085 29.1 0.085 ;
      RECT 28.93 2.635 29.1 2.805 ;
      RECT 28.47 -0.085 28.64 0.085 ;
      RECT 28.47 2.635 28.64 2.805 ;
      RECT 28.415 1.515 28.585 1.685 ;
      RECT 28.01 -0.085 28.18 0.085 ;
      RECT 28.01 2.635 28.18 2.805 ;
      RECT 27.55 -0.085 27.72 0.085 ;
      RECT 27.55 2.635 27.72 2.805 ;
      RECT 27.09 -0.085 27.26 0.085 ;
      RECT 27.09 2.635 27.26 2.805 ;
      RECT 26.63 -0.085 26.8 0.085 ;
      RECT 26.63 2.635 26.8 2.805 ;
      RECT 26.425 1.105 26.595 1.275 ;
      RECT 26.17 -0.085 26.34 0.085 ;
      RECT 26.17 2.635 26.34 2.805 ;
      RECT 25.71 -0.085 25.88 0.085 ;
      RECT 25.71 2.635 25.88 2.805 ;
      RECT 25.25 -0.085 25.42 0.085 ;
      RECT 25.25 2.635 25.42 2.805 ;
      RECT 25.18 1.46 25.35 1.63 ;
      RECT 24.79 -0.085 24.96 0.085 ;
      RECT 24.79 2.635 24.96 2.805 ;
      RECT 24.33 -0.085 24.5 0.085 ;
      RECT 24.33 2.635 24.5 2.805 ;
      RECT 24.32 0.575 24.49 0.745 ;
      RECT 23.875 0.455 24.045 0.625 ;
      RECT 23.87 -0.085 24.04 0.085 ;
      RECT 23.87 2.635 24.04 2.805 ;
      RECT 23.41 -0.085 23.58 0.085 ;
      RECT 23.41 2.635 23.58 2.805 ;
      RECT 22.95 -0.085 23.12 0.085 ;
      RECT 22.95 2.635 23.12 2.805 ;
      RECT 22.49 -0.085 22.66 0.085 ;
      RECT 22.49 2.635 22.66 2.805 ;
      RECT 22.03 -0.085 22.2 0.085 ;
      RECT 22.03 2.635 22.2 2.805 ;
      RECT 21.975 1.075 22.145 1.245 ;
      RECT 21.575 -0.085 21.745 0.085 ;
      RECT 21.575 2.635 21.745 2.805 ;
      RECT 21.115 -0.085 21.285 0.085 ;
      RECT 21.115 2.635 21.285 2.805 ;
      RECT 21.045 1.46 21.215 1.63 ;
      RECT 20.655 -0.085 20.825 0.085 ;
      RECT 20.655 2.635 20.825 2.805 ;
      RECT 20.195 -0.085 20.365 0.085 ;
      RECT 20.195 2.635 20.365 2.805 ;
      RECT 19.78 0.515 19.95 0.685 ;
      RECT 19.735 -0.085 19.905 0.085 ;
      RECT 19.735 2.635 19.905 2.805 ;
      RECT 19.365 1.24 19.535 1.41 ;
      RECT 19.275 -0.085 19.445 0.085 ;
      RECT 19.275 2.635 19.445 2.805 ;
      RECT 18.815 -0.085 18.985 0.085 ;
      RECT 18.815 2.635 18.985 2.805 ;
      RECT 18.355 -0.085 18.525 0.085 ;
      RECT 18.355 2.635 18.525 2.805 ;
      RECT 17.895 -0.085 18.065 0.085 ;
      RECT 17.895 2.635 18.065 2.805 ;
      RECT 17.84 1.915 18.01 2.085 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 17.435 2.635 17.605 2.805 ;
      RECT 17.065 1.375 17.235 1.545 ;
      RECT 16.975 -0.085 17.145 0.085 ;
      RECT 16.975 2.635 17.145 2.805 ;
      RECT 16.745 0.545 16.915 0.715 ;
      RECT 16.6 0.985 16.77 1.155 ;
      RECT 16.515 -0.085 16.685 0.085 ;
      RECT 16.515 2.635 16.685 2.805 ;
      RECT 16.055 -0.085 16.225 0.085 ;
      RECT 16.055 2.635 16.225 2.805 ;
      RECT 15.99 1.025 16.16 1.195 ;
      RECT 15.645 0.66 15.815 0.83 ;
      RECT 15.635 2.02 15.805 2.19 ;
      RECT 15.595 -0.085 15.765 0.085 ;
      RECT 15.595 2.635 15.765 2.805 ;
      RECT 15.22 1.26 15.39 1.43 ;
      RECT 15.135 -0.085 15.305 0.085 ;
      RECT 15.135 2.635 15.305 2.805 ;
      RECT 14.87 0.735 15.04 0.905 ;
      RECT 14.69 2.05 14.86 2.22 ;
      RECT 14.675 -0.085 14.845 0.085 ;
      RECT 14.675 2.635 14.845 2.805 ;
      RECT 14.41 1.365 14.58 1.535 ;
      RECT 14.215 -0.085 14.385 0.085 ;
      RECT 14.215 2.635 14.385 2.805 ;
      RECT 14.09 0.99 14.26 1.16 ;
      RECT 13.755 -0.085 13.925 0.085 ;
      RECT 13.755 2.635 13.925 2.805 ;
      RECT 13.4 0.47 13.57 0.64 ;
      RECT 13.325 0.94 13.495 1.11 ;
      RECT 13.295 -0.085 13.465 0.085 ;
      RECT 13.295 2.635 13.465 2.805 ;
      RECT 12.835 -0.085 13.005 0.085 ;
      RECT 12.835 2.635 13.005 2.805 ;
      RECT 12.475 0.665 12.645 0.835 ;
      RECT 12.375 -0.085 12.545 0.085 ;
      RECT 12.375 2.635 12.545 2.805 ;
      RECT 12.135 1.86 12.305 2.03 ;
      RECT 12.1 1.195 12.27 1.365 ;
      RECT 11.915 -0.085 12.085 0.085 ;
      RECT 11.915 2.635 12.085 2.805 ;
      RECT 11.49 1.05 11.66 1.22 ;
      RECT 11.455 -0.085 11.625 0.085 ;
      RECT 11.455 2.635 11.625 2.805 ;
      RECT 11.42 1.75 11.59 1.92 ;
      RECT 11.36 0.585 11.53 0.755 ;
      RECT 10.995 -0.085 11.165 0.085 ;
      RECT 10.995 2.635 11.165 2.805 ;
      RECT 10.72 1.5 10.89 1.67 ;
      RECT 10.535 -0.085 10.705 0.085 ;
      RECT 10.535 2.635 10.705 2.805 ;
      RECT 10.215 1.005 10.385 1.175 ;
      RECT 10.075 -0.085 10.245 0.085 ;
      RECT 10.075 2.635 10.245 2.805 ;
      RECT 9.995 1.75 10.165 1.92 ;
      RECT 9.79 0.63 9.96 0.8 ;
      RECT 9.615 -0.085 9.785 0.085 ;
      RECT 9.615 2.635 9.785 2.805 ;
      RECT 9.52 1.5 9.69 1.67 ;
      RECT 9.48 0.93 9.65 1.1 ;
      RECT 9.155 -0.085 9.325 0.085 ;
      RECT 9.155 2.635 9.325 2.805 ;
      RECT 8.935 1.975 9.105 2.145 ;
      RECT 8.795 0.595 8.965 0.765 ;
      RECT 8.695 -0.085 8.865 0.085 ;
      RECT 8.695 2.635 8.865 2.805 ;
      RECT 8.235 -0.085 8.405 0.085 ;
      RECT 8.235 2.635 8.405 2.805 ;
      RECT 8.225 1.515 8.395 1.685 ;
      RECT 7.775 -0.085 7.945 0.085 ;
      RECT 7.775 2.635 7.945 2.805 ;
      RECT 7.315 -0.085 7.485 0.085 ;
      RECT 7.315 2.635 7.485 2.805 ;
      RECT 7.245 1.46 7.415 1.63 ;
      RECT 6.855 -0.085 7.025 0.085 ;
      RECT 6.855 2.635 7.025 2.805 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 2.635 6.565 2.805 ;
      RECT 6.385 0.505 6.555 0.675 ;
      RECT 5.935 -0.085 6.105 0.085 ;
      RECT 5.935 2.635 6.105 2.805 ;
      RECT 5.475 -0.085 5.645 0.085 ;
      RECT 5.475 2.635 5.645 2.805 ;
      RECT 5.015 -0.085 5.185 0.085 ;
      RECT 5.015 2.635 5.185 2.805 ;
      RECT 4.555 -0.085 4.725 0.085 ;
      RECT 4.555 2.635 4.725 2.805 ;
      RECT 4.095 -0.085 4.265 0.085 ;
      RECT 4.095 2.635 4.265 2.805 ;
      RECT 4.04 1.575 4.21 1.745 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.455 1.7 2.625 1.87 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.025 0.695 2.195 0.865 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.175 1.815 0.345 1.985 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
    LAYER li ;
      RECT 116.32 -0.085 116.595 1.415 ;
      RECT 88.725 -0.085 89 1.415 ;
      RECT 61.13 -0.085 61.405 1.415 ;
      RECT 33.535 -0.085 33.81 1.415 ;
      RECT 5.94 -0.085 6.215 1.415 ;
      RECT 140.865 -0.085 141.095 0.905 ;
      RECT 139.485 -0.085 139.715 0.905 ;
      RECT 138.105 -0.085 138.335 0.905 ;
      RECT 136.725 -0.085 136.955 0.905 ;
      RECT 113.27 -0.085 113.5 0.905 ;
      RECT 111.89 -0.085 112.12 0.905 ;
      RECT 110.51 -0.085 110.74 0.905 ;
      RECT 109.13 -0.085 109.36 0.905 ;
      RECT 85.675 -0.085 85.905 0.905 ;
      RECT 84.295 -0.085 84.525 0.905 ;
      RECT 82.915 -0.085 83.145 0.905 ;
      RECT 81.535 -0.085 81.765 0.905 ;
      RECT 58.08 -0.085 58.31 0.905 ;
      RECT 56.7 -0.085 56.93 0.905 ;
      RECT 55.32 -0.085 55.55 0.905 ;
      RECT 53.94 -0.085 54.17 0.905 ;
      RECT 30.485 -0.085 30.715 0.905 ;
      RECT 29.105 -0.085 29.335 0.905 ;
      RECT 27.725 -0.085 27.955 0.905 ;
      RECT 26.345 -0.085 26.575 0.905 ;
      RECT 135.07 -0.085 135.58 0.62 ;
      RECT 130.935 -0.085 131.445 0.62 ;
      RECT 117.135 -0.085 117.645 0.62 ;
      RECT 107.475 -0.085 107.985 0.62 ;
      RECT 103.34 -0.085 103.85 0.62 ;
      RECT 89.54 -0.085 90.05 0.62 ;
      RECT 79.88 -0.085 80.39 0.62 ;
      RECT 75.745 -0.085 76.255 0.62 ;
      RECT 61.945 -0.085 62.455 0.62 ;
      RECT 52.285 -0.085 52.795 0.62 ;
      RECT 48.15 -0.085 48.66 0.62 ;
      RECT 34.35 -0.085 34.86 0.62 ;
      RECT 24.69 -0.085 25.2 0.62 ;
      RECT 20.555 -0.085 21.065 0.62 ;
      RECT 6.755 -0.085 7.265 0.62 ;
      RECT 2.805 -0.085 3.315 0.62 ;
      RECT 126.6 -0.085 126.77 0.585 ;
      RECT 124.64 -0.085 124.81 0.585 ;
      RECT 122.2 -0.085 122.37 0.585 ;
      RECT 121.24 -0.085 121.41 0.585 ;
      RECT 120.72 -0.085 120.89 0.585 ;
      RECT 119.76 -0.085 119.93 0.585 ;
      RECT 118.8 -0.085 118.97 0.585 ;
      RECT 99.005 -0.085 99.175 0.585 ;
      RECT 97.045 -0.085 97.215 0.585 ;
      RECT 94.605 -0.085 94.775 0.585 ;
      RECT 93.645 -0.085 93.815 0.585 ;
      RECT 93.125 -0.085 93.295 0.585 ;
      RECT 92.165 -0.085 92.335 0.585 ;
      RECT 91.205 -0.085 91.375 0.585 ;
      RECT 71.41 -0.085 71.58 0.585 ;
      RECT 69.45 -0.085 69.62 0.585 ;
      RECT 67.01 -0.085 67.18 0.585 ;
      RECT 66.05 -0.085 66.22 0.585 ;
      RECT 65.53 -0.085 65.7 0.585 ;
      RECT 64.57 -0.085 64.74 0.585 ;
      RECT 63.61 -0.085 63.78 0.585 ;
      RECT 43.815 -0.085 43.985 0.585 ;
      RECT 41.855 -0.085 42.025 0.585 ;
      RECT 39.415 -0.085 39.585 0.585 ;
      RECT 38.455 -0.085 38.625 0.585 ;
      RECT 37.935 -0.085 38.105 0.585 ;
      RECT 36.975 -0.085 37.145 0.585 ;
      RECT 36.015 -0.085 36.185 0.585 ;
      RECT 16.22 -0.085 16.39 0.585 ;
      RECT 14.26 -0.085 14.43 0.585 ;
      RECT 11.82 -0.085 11.99 0.585 ;
      RECT 10.86 -0.085 11.03 0.585 ;
      RECT 10.34 -0.085 10.51 0.585 ;
      RECT 9.38 -0.085 9.55 0.585 ;
      RECT 8.42 -0.085 8.59 0.585 ;
      RECT 132.78 -0.085 133.11 0.485 ;
      RECT 128.645 -0.085 128.975 0.485 ;
      RECT 114.845 -0.085 115.175 0.485 ;
      RECT 105.185 -0.085 105.515 0.485 ;
      RECT 101.05 -0.085 101.38 0.485 ;
      RECT 87.25 -0.085 87.58 0.485 ;
      RECT 77.59 -0.085 77.92 0.485 ;
      RECT 73.455 -0.085 73.785 0.485 ;
      RECT 59.655 -0.085 59.985 0.485 ;
      RECT 49.995 -0.085 50.325 0.485 ;
      RECT 45.86 -0.085 46.19 0.485 ;
      RECT 32.06 -0.085 32.39 0.485 ;
      RECT 22.4 -0.085 22.73 0.485 ;
      RECT 18.265 -0.085 18.595 0.485 ;
      RECT 4.465 -0.085 4.795 0.485 ;
      RECT 0.515 -0.085 0.845 0.485 ;
      RECT 0 -0.085 141.925 0.085 ;
      RECT 0 2.635 141.925 2.805 ;
      RECT 140.885 1.495 141.095 2.805 ;
      RECT 139.505 1.495 139.715 2.805 ;
      RECT 138.125 1.495 138.335 2.805 ;
      RECT 136.745 1.495 136.955 2.805 ;
      RECT 135.4 1.875 135.57 2.805 ;
      RECT 132.86 1.495 133.03 2.805 ;
      RECT 131.265 1.875 131.435 2.805 ;
      RECT 128.725 1.495 128.895 2.805 ;
      RECT 127.56 2.045 127.73 2.805 ;
      RECT 126.6 2.135 126.77 2.805 ;
      RECT 124.16 2.135 124.33 2.805 ;
      RECT 123.16 2.135 123.33 2.805 ;
      RECT 122.2 2.135 122.37 2.805 ;
      RECT 119.76 2.135 119.93 2.805 ;
      RECT 117.465 1.875 117.635 2.805 ;
      RECT 114.925 1.495 115.095 2.805 ;
      RECT 113.29 1.495 113.5 2.805 ;
      RECT 111.91 1.495 112.12 2.805 ;
      RECT 110.53 1.495 110.74 2.805 ;
      RECT 109.15 1.495 109.36 2.805 ;
      RECT 107.805 1.875 107.975 2.805 ;
      RECT 105.265 1.495 105.435 2.805 ;
      RECT 103.67 1.875 103.84 2.805 ;
      RECT 101.13 1.495 101.3 2.805 ;
      RECT 99.965 2.045 100.135 2.805 ;
      RECT 99.005 2.135 99.175 2.805 ;
      RECT 96.565 2.135 96.735 2.805 ;
      RECT 95.565 2.135 95.735 2.805 ;
      RECT 94.605 2.135 94.775 2.805 ;
      RECT 92.165 2.135 92.335 2.805 ;
      RECT 89.87 1.875 90.04 2.805 ;
      RECT 87.33 1.495 87.5 2.805 ;
      RECT 85.695 1.495 85.905 2.805 ;
      RECT 84.315 1.495 84.525 2.805 ;
      RECT 82.935 1.495 83.145 2.805 ;
      RECT 81.555 1.495 81.765 2.805 ;
      RECT 80.21 1.875 80.38 2.805 ;
      RECT 77.67 1.495 77.84 2.805 ;
      RECT 76.075 1.875 76.245 2.805 ;
      RECT 73.535 1.495 73.705 2.805 ;
      RECT 72.37 2.045 72.54 2.805 ;
      RECT 71.41 2.135 71.58 2.805 ;
      RECT 68.97 2.135 69.14 2.805 ;
      RECT 67.97 2.135 68.14 2.805 ;
      RECT 67.01 2.135 67.18 2.805 ;
      RECT 64.57 2.135 64.74 2.805 ;
      RECT 62.275 1.875 62.445 2.805 ;
      RECT 59.735 1.495 59.905 2.805 ;
      RECT 58.1 1.495 58.31 2.805 ;
      RECT 56.72 1.495 56.93 2.805 ;
      RECT 55.34 1.495 55.55 2.805 ;
      RECT 53.96 1.495 54.17 2.805 ;
      RECT 52.615 1.875 52.785 2.805 ;
      RECT 50.075 1.495 50.245 2.805 ;
      RECT 48.48 1.875 48.65 2.805 ;
      RECT 45.94 1.495 46.11 2.805 ;
      RECT 44.775 2.045 44.945 2.805 ;
      RECT 43.815 2.135 43.985 2.805 ;
      RECT 41.375 2.135 41.545 2.805 ;
      RECT 40.375 2.135 40.545 2.805 ;
      RECT 39.415 2.135 39.585 2.805 ;
      RECT 36.975 2.135 37.145 2.805 ;
      RECT 34.68 1.875 34.85 2.805 ;
      RECT 32.14 1.495 32.31 2.805 ;
      RECT 30.505 1.495 30.715 2.805 ;
      RECT 29.125 1.495 29.335 2.805 ;
      RECT 27.745 1.495 27.955 2.805 ;
      RECT 26.365 1.495 26.575 2.805 ;
      RECT 25.02 1.875 25.19 2.805 ;
      RECT 22.48 1.495 22.65 2.805 ;
      RECT 20.885 1.875 21.055 2.805 ;
      RECT 18.345 1.495 18.515 2.805 ;
      RECT 17.18 2.045 17.35 2.805 ;
      RECT 16.22 2.135 16.39 2.805 ;
      RECT 13.78 2.135 13.95 2.805 ;
      RECT 12.78 2.135 12.95 2.805 ;
      RECT 11.82 2.135 11.99 2.805 ;
      RECT 9.38 2.135 9.55 2.805 ;
      RECT 7.085 1.875 7.255 2.805 ;
      RECT 4.545 1.495 4.715 2.805 ;
      RECT 3.135 1.875 3.305 2.805 ;
      RECT 0.595 1.495 0.765 2.805 ;
      RECT 141.265 1.485 141.595 2.465 ;
      RECT 141.365 0.255 141.595 2.465 ;
      RECT 141.265 1.79 141.725 1.94 ;
      RECT 141.265 0.255 141.595 0.885 ;
      RECT 139.885 1.485 140.215 2.465 ;
      RECT 139.985 0.255 140.215 2.465 ;
      RECT 139.985 1.075 141.195 1.315 ;
      RECT 139.885 0.255 140.215 0.885 ;
      RECT 138.505 1.485 138.835 2.465 ;
      RECT 138.605 0.255 138.835 2.465 ;
      RECT 138.605 0.895 138.965 1.065 ;
      RECT 138.505 0.255 138.835 0.885 ;
      RECT 137.125 1.485 137.455 2.465 ;
      RECT 137.225 0.255 137.455 2.465 ;
      RECT 137.225 1.075 138.435 1.315 ;
      RECT 137.125 0.255 137.455 0.885 ;
      RECT 135.805 1.875 136.32 2.285 ;
      RECT 135.98 0.895 136.32 2.285 ;
      RECT 135.09 0.895 136.32 1.065 ;
      RECT 135.8 0.29 136.045 1.065 ;
      RECT 133.2 2.295 135.23 2.465 ;
      RECT 135.06 1.44 135.23 2.465 ;
      RECT 133.2 0.995 133.37 2.465 ;
      RECT 135.06 1.44 135.81 1.63 ;
      RECT 133.175 0.995 133.37 1.325 ;
      RECT 133.88 1.615 134.89 1.785 ;
      RECT 134.7 0.255 134.89 1.785 ;
      RECT 133.88 0.815 134.05 1.785 ;
      RECT 133.54 1.955 134.665 2.125 ;
      RECT 133.54 0.255 133.71 2.125 ;
      RECT 132.695 0.995 132.95 1.325 ;
      RECT 132.78 0.655 132.95 1.325 ;
      RECT 132.78 0.655 133.71 0.825 ;
      RECT 133.535 0.255 133.71 0.825 ;
      RECT 133.535 0.255 134.065 0.62 ;
      RECT 132.355 1.495 132.69 2.465 ;
      RECT 132.355 0.255 132.525 2.465 ;
      RECT 132.355 0.255 132.61 0.825 ;
      RECT 131.67 1.875 132.185 2.285 ;
      RECT 131.845 0.895 132.185 2.285 ;
      RECT 130.955 0.895 132.185 1.065 ;
      RECT 131.665 0.29 131.91 1.065 ;
      RECT 129.065 2.295 131.095 2.465 ;
      RECT 130.925 1.44 131.095 2.465 ;
      RECT 129.065 0.995 129.235 2.465 ;
      RECT 130.925 1.44 131.675 1.63 ;
      RECT 129.04 0.995 129.235 1.325 ;
      RECT 129.745 1.615 130.755 1.785 ;
      RECT 130.565 0.255 130.755 1.785 ;
      RECT 129.745 0.815 129.915 1.785 ;
      RECT 129.405 1.955 130.53 2.125 ;
      RECT 129.405 0.255 129.575 2.125 ;
      RECT 128.56 0.995 128.815 1.325 ;
      RECT 128.645 0.655 128.815 1.325 ;
      RECT 128.645 0.655 129.575 0.825 ;
      RECT 129.4 0.255 129.575 0.825 ;
      RECT 129.4 0.255 129.93 0.62 ;
      RECT 128.22 1.495 128.555 2.465 ;
      RECT 128.22 0.255 128.39 2.465 ;
      RECT 128.22 0.255 128.475 0.825 ;
      RECT 127.125 0.475 127.855 0.715 ;
      RECT 127.667 0.27 127.855 0.715 ;
      RECT 127.495 0.282 127.87 0.709 ;
      RECT 127.41 0.297 127.89 0.694 ;
      RECT 127.41 0.312 127.895 0.684 ;
      RECT 127.365 0.332 127.91 0.676 ;
      RECT 127.342 0.367 127.925 0.63 ;
      RECT 127.256 0.39 127.93 0.59 ;
      RECT 127.256 0.408 127.94 0.56 ;
      RECT 127.125 0.477 127.945 0.523 ;
      RECT 127.17 0.42 127.94 0.56 ;
      RECT 127.256 0.372 127.925 0.63 ;
      RECT 127.342 0.341 127.91 0.676 ;
      RECT 127.365 0.322 127.895 0.684 ;
      RECT 127.41 0.295 127.87 0.709 ;
      RECT 127.495 0.277 127.855 0.715 ;
      RECT 127.581 0.271 127.855 0.715 ;
      RECT 127.667 0.266 127.8 0.715 ;
      RECT 127.753 0.261 127.8 0.715 ;
      RECT 127.445 1.159 127.615 1.545 ;
      RECT 127.44 1.159 127.615 1.54 ;
      RECT 127.415 1.159 127.615 1.505 ;
      RECT 127.415 1.187 127.625 1.495 ;
      RECT 127.395 1.187 127.625 1.455 ;
      RECT 127.39 1.187 127.625 1.428 ;
      RECT 127.39 1.205 127.63 1.42 ;
      RECT 127.335 1.205 127.63 1.355 ;
      RECT 127.335 1.222 127.64 1.338 ;
      RECT 127.325 1.222 127.64 1.278 ;
      RECT 127.325 1.239 127.645 1.275 ;
      RECT 127.32 1.075 127.49 1.253 ;
      RECT 127.32 1.109 127.576 1.253 ;
      RECT 127.315 1.875 127.32 1.888 ;
      RECT 127.31 1.77 127.315 1.893 ;
      RECT 127.285 1.63 127.31 1.908 ;
      RECT 127.25 1.581 127.285 1.94 ;
      RECT 127.245 1.549 127.25 1.96 ;
      RECT 127.24 1.54 127.245 1.96 ;
      RECT 127.16 1.505 127.24 1.96 ;
      RECT 127.097 1.475 127.16 1.96 ;
      RECT 127.011 1.463 127.097 1.96 ;
      RECT 126.925 1.449 127.011 1.96 ;
      RECT 126.845 1.436 126.925 1.946 ;
      RECT 126.81 1.428 126.845 1.926 ;
      RECT 126.8 1.425 126.81 1.917 ;
      RECT 126.77 1.42 126.8 1.904 ;
      RECT 126.72 1.395 126.77 1.88 ;
      RECT 126.706 1.369 126.72 1.862 ;
      RECT 126.62 1.329 126.706 1.838 ;
      RECT 126.575 1.277 126.62 1.807 ;
      RECT 126.565 1.252 126.575 1.794 ;
      RECT 126.56 1.033 126.565 1.055 ;
      RECT 126.555 1.235 126.565 1.79 ;
      RECT 126.555 1.031 126.56 1.145 ;
      RECT 126.545 1.027 126.555 1.786 ;
      RECT 126.501 1.025 126.545 1.774 ;
      RECT 126.415 1.025 126.501 1.745 ;
      RECT 126.385 1.025 126.415 1.718 ;
      RECT 126.37 1.025 126.385 1.706 ;
      RECT 126.33 1.037 126.37 1.691 ;
      RECT 126.31 1.056 126.33 1.67 ;
      RECT 126.3 1.066 126.31 1.654 ;
      RECT 126.29 1.072 126.3 1.643 ;
      RECT 126.27 1.082 126.29 1.626 ;
      RECT 126.265 1.091 126.27 1.613 ;
      RECT 126.26 1.095 126.265 1.563 ;
      RECT 126.25 1.101 126.26 1.48 ;
      RECT 126.245 1.105 126.25 1.394 ;
      RECT 126.24 1.125 126.245 1.331 ;
      RECT 126.235 1.148 126.24 1.278 ;
      RECT 126.23 1.166 126.235 1.223 ;
      RECT 126.84 0.985 127.01 1.245 ;
      RECT 127.01 0.95 127.055 1.231 ;
      RECT 126.971 0.952 127.06 1.214 ;
      RECT 126.86 0.969 127.146 1.185 ;
      RECT 126.86 0.984 127.15 1.157 ;
      RECT 126.86 0.965 127.06 1.214 ;
      RECT 126.885 0.953 127.01 1.245 ;
      RECT 126.971 0.951 127.055 1.231 ;
      RECT 126.025 0.34 126.195 0.83 ;
      RECT 126.025 0.34 126.23 0.81 ;
      RECT 126.16 0.26 126.27 0.77 ;
      RECT 126.141 0.264 126.29 0.74 ;
      RECT 126.055 0.272 126.31 0.723 ;
      RECT 126.055 0.278 126.315 0.713 ;
      RECT 126.055 0.287 126.335 0.701 ;
      RECT 126.03 0.312 126.365 0.679 ;
      RECT 126.03 0.332 126.37 0.659 ;
      RECT 126.025 0.345 126.38 0.639 ;
      RECT 126.025 0.412 126.385 0.62 ;
      RECT 126.025 0.545 126.39 0.607 ;
      RECT 126.02 0.35 126.38 0.44 ;
      RECT 126.03 0.307 126.335 0.701 ;
      RECT 126.141 0.262 126.27 0.77 ;
      RECT 126.015 2.015 126.315 2.27 ;
      RECT 126.1 1.981 126.315 2.27 ;
      RECT 126.1 1.984 126.32 2.13 ;
      RECT 126.035 2.005 126.32 2.13 ;
      RECT 126.07 1.995 126.315 2.27 ;
      RECT 126.065 2 126.32 2.13 ;
      RECT 126.1 1.979 126.301 2.27 ;
      RECT 126.186 1.97 126.301 2.27 ;
      RECT 126.186 1.964 126.215 2.27 ;
      RECT 125.675 1.605 125.685 2.095 ;
      RECT 125.335 1.54 125.345 1.84 ;
      RECT 125.85 1.712 125.855 1.931 ;
      RECT 125.84 1.692 125.85 1.948 ;
      RECT 125.83 1.672 125.84 1.978 ;
      RECT 125.825 1.662 125.83 1.993 ;
      RECT 125.82 1.658 125.825 1.998 ;
      RECT 125.805 1.65 125.82 2.005 ;
      RECT 125.765 1.63 125.805 2.03 ;
      RECT 125.74 1.612 125.765 2.063 ;
      RECT 125.735 1.61 125.74 2.076 ;
      RECT 125.715 1.607 125.735 2.08 ;
      RECT 125.685 1.605 125.715 2.09 ;
      RECT 125.615 1.607 125.675 2.091 ;
      RECT 125.595 1.607 125.615 2.085 ;
      RECT 125.57 1.605 125.595 2.082 ;
      RECT 125.535 1.6 125.57 2.078 ;
      RECT 125.515 1.594 125.535 2.065 ;
      RECT 125.505 1.591 125.515 2.053 ;
      RECT 125.485 1.588 125.505 2.038 ;
      RECT 125.465 1.584 125.485 2.02 ;
      RECT 125.46 1.581 125.465 2.01 ;
      RECT 125.455 1.58 125.46 2.008 ;
      RECT 125.445 1.577 125.455 2 ;
      RECT 125.435 1.571 125.445 1.983 ;
      RECT 125.425 1.565 125.435 1.965 ;
      RECT 125.415 1.559 125.425 1.953 ;
      RECT 125.405 1.553 125.415 1.933 ;
      RECT 125.4 1.549 125.405 1.918 ;
      RECT 125.395 1.547 125.4 1.91 ;
      RECT 125.39 1.545 125.395 1.903 ;
      RECT 125.385 1.543 125.39 1.893 ;
      RECT 125.38 1.541 125.385 1.887 ;
      RECT 125.37 1.54 125.38 1.877 ;
      RECT 125.36 1.54 125.37 1.868 ;
      RECT 125.345 1.54 125.36 1.853 ;
      RECT 125.305 1.54 125.335 1.837 ;
      RECT 125.285 1.542 125.305 1.832 ;
      RECT 125.28 1.547 125.285 1.83 ;
      RECT 125.25 1.555 125.28 1.828 ;
      RECT 125.22 1.57 125.25 1.827 ;
      RECT 125.175 1.592 125.22 1.832 ;
      RECT 125.17 1.607 125.175 1.836 ;
      RECT 125.155 1.612 125.17 1.838 ;
      RECT 125.15 1.616 125.155 1.84 ;
      RECT 125.09 1.639 125.15 1.849 ;
      RECT 125.07 1.665 125.09 1.862 ;
      RECT 125.06 1.672 125.07 1.866 ;
      RECT 125.045 1.679 125.06 1.869 ;
      RECT 125.025 1.689 125.045 1.872 ;
      RECT 125.02 1.697 125.025 1.875 ;
      RECT 124.975 1.702 125.02 1.882 ;
      RECT 124.965 1.705 124.975 1.889 ;
      RECT 124.955 1.705 124.965 1.893 ;
      RECT 124.92 1.707 124.955 1.905 ;
      RECT 124.9 1.71 124.92 1.918 ;
      RECT 124.86 1.713 124.9 1.929 ;
      RECT 124.845 1.715 124.86 1.942 ;
      RECT 124.835 1.715 124.845 1.947 ;
      RECT 124.81 1.716 124.835 1.955 ;
      RECT 124.8 1.718 124.81 1.96 ;
      RECT 124.795 1.719 124.8 1.963 ;
      RECT 124.77 1.717 124.795 1.966 ;
      RECT 124.755 1.715 124.77 1.967 ;
      RECT 124.735 1.712 124.755 1.969 ;
      RECT 124.715 1.707 124.735 1.969 ;
      RECT 124.655 1.702 124.715 1.966 ;
      RECT 124.62 1.677 124.655 1.962 ;
      RECT 124.61 1.654 124.62 1.96 ;
      RECT 124.58 1.631 124.61 1.96 ;
      RECT 124.57 1.61 124.58 1.96 ;
      RECT 124.545 1.592 124.57 1.958 ;
      RECT 124.53 1.57 124.545 1.955 ;
      RECT 124.515 1.552 124.53 1.953 ;
      RECT 124.495 1.542 124.515 1.951 ;
      RECT 124.48 1.537 124.495 1.95 ;
      RECT 124.465 1.535 124.48 1.949 ;
      RECT 124.435 1.536 124.465 1.947 ;
      RECT 124.415 1.539 124.435 1.945 ;
      RECT 124.358 1.543 124.415 1.945 ;
      RECT 124.272 1.552 124.358 1.945 ;
      RECT 124.186 1.563 124.272 1.945 ;
      RECT 124.1 1.574 124.186 1.945 ;
      RECT 124.08 1.581 124.1 1.953 ;
      RECT 124.07 1.584 124.08 1.96 ;
      RECT 124.005 1.589 124.07 1.978 ;
      RECT 123.975 1.596 124.005 2.003 ;
      RECT 123.965 1.599 123.975 2.01 ;
      RECT 123.92 1.603 123.965 2.015 ;
      RECT 123.89 1.608 123.92 2.02 ;
      RECT 123.889 1.61 123.89 2.02 ;
      RECT 123.803 1.616 123.889 2.02 ;
      RECT 123.717 1.627 123.803 2.02 ;
      RECT 123.631 1.639 123.717 2.02 ;
      RECT 123.545 1.65 123.631 2.02 ;
      RECT 123.53 1.657 123.545 2.015 ;
      RECT 123.525 1.659 123.53 2.009 ;
      RECT 123.505 1.67 123.525 2.004 ;
      RECT 123.495 1.688 123.505 1.998 ;
      RECT 123.49 1.7 123.495 1.798 ;
      RECT 125.785 0.453 125.805 0.54 ;
      RECT 125.78 0.388 125.785 0.572 ;
      RECT 125.77 0.355 125.78 0.577 ;
      RECT 125.765 0.335 125.77 0.583 ;
      RECT 125.735 0.335 125.765 0.6 ;
      RECT 125.686 0.335 125.735 0.636 ;
      RECT 125.6 0.335 125.686 0.694 ;
      RECT 125.571 0.345 125.6 0.743 ;
      RECT 125.485 0.387 125.571 0.796 ;
      RECT 125.465 0.425 125.485 0.843 ;
      RECT 125.44 0.442 125.465 0.863 ;
      RECT 125.43 0.456 125.44 0.883 ;
      RECT 125.425 0.462 125.43 0.893 ;
      RECT 125.42 0.466 125.425 0.9 ;
      RECT 125.37 0.486 125.42 0.905 ;
      RECT 125.305 0.53 125.37 0.905 ;
      RECT 125.28 0.58 125.305 0.905 ;
      RECT 125.27 0.61 125.28 0.905 ;
      RECT 125.265 0.637 125.27 0.905 ;
      RECT 125.26 0.655 125.265 0.905 ;
      RECT 125.25 0.697 125.26 0.905 ;
      RECT 125.6 1.255 125.77 1.43 ;
      RECT 125.54 1.083 125.6 1.418 ;
      RECT 125.53 1.076 125.54 1.401 ;
      RECT 125.485 1.255 125.77 1.381 ;
      RECT 125.466 1.255 125.77 1.359 ;
      RECT 125.38 1.255 125.77 1.324 ;
      RECT 125.36 1.075 125.53 1.28 ;
      RECT 125.36 1.222 125.765 1.28 ;
      RECT 125.36 1.17 125.74 1.28 ;
      RECT 125.36 1.125 125.705 1.28 ;
      RECT 125.36 1.107 125.67 1.28 ;
      RECT 125.36 1.097 125.665 1.28 ;
      RECT 125.08 2.055 125.27 2.28 ;
      RECT 125.07 2.056 125.275 2.275 ;
      RECT 125.07 2.058 125.285 2.255 ;
      RECT 125.07 2.062 125.29 2.24 ;
      RECT 125.07 2.049 125.24 2.275 ;
      RECT 125.07 2.052 125.265 2.275 ;
      RECT 125.08 2.048 125.24 2.28 ;
      RECT 125.166 2.046 125.24 2.28 ;
      RECT 124.79 1.297 124.96 1.535 ;
      RECT 124.79 1.297 125.046 1.449 ;
      RECT 124.79 1.297 125.05 1.359 ;
      RECT 124.84 1.07 125.06 1.338 ;
      RECT 124.835 1.087 125.065 1.311 ;
      RECT 124.8 1.245 125.065 1.311 ;
      RECT 124.82 1.095 124.96 1.535 ;
      RECT 124.81 1.177 125.07 1.294 ;
      RECT 124.805 1.225 125.07 1.294 ;
      RECT 124.81 1.135 125.065 1.311 ;
      RECT 124.835 1.072 125.06 1.338 ;
      RECT 124.4 1.047 124.57 1.245 ;
      RECT 124.4 1.047 124.615 1.22 ;
      RECT 124.47 0.99 124.64 1.178 ;
      RECT 124.445 1.005 124.64 1.178 ;
      RECT 124.06 1.051 124.09 1.245 ;
      RECT 124.055 1.023 124.06 1.245 ;
      RECT 124.025 0.997 124.055 1.247 ;
      RECT 124 0.955 124.025 1.25 ;
      RECT 123.99 0.927 124 1.252 ;
      RECT 123.955 0.907 123.99 1.254 ;
      RECT 123.89 0.892 123.955 1.26 ;
      RECT 123.84 0.89 123.89 1.266 ;
      RECT 123.817 0.892 123.84 1.271 ;
      RECT 123.731 0.903 123.817 1.277 ;
      RECT 123.645 0.921 123.731 1.287 ;
      RECT 123.63 0.932 123.645 1.293 ;
      RECT 123.56 0.955 123.63 1.299 ;
      RECT 123.505 0.987 123.56 1.307 ;
      RECT 123.465 1.01 123.505 1.313 ;
      RECT 123.451 1.023 123.465 1.316 ;
      RECT 123.365 1.045 123.451 1.322 ;
      RECT 123.35 1.07 123.365 1.328 ;
      RECT 123.31 1.085 123.35 1.332 ;
      RECT 123.26 1.1 123.31 1.337 ;
      RECT 123.235 1.107 123.26 1.341 ;
      RECT 123.175 1.102 123.235 1.345 ;
      RECT 123.16 1.093 123.175 1.349 ;
      RECT 123.09 1.083 123.16 1.345 ;
      RECT 123.065 1.075 123.085 1.335 ;
      RECT 123.006 1.075 123.065 1.313 ;
      RECT 122.92 1.075 123.006 1.27 ;
      RECT 123.085 1.075 123.09 1.34 ;
      RECT 123.78 0.306 123.95 0.64 ;
      RECT 123.75 0.306 123.95 0.635 ;
      RECT 123.69 0.273 123.75 0.623 ;
      RECT 123.69 0.329 123.96 0.618 ;
      RECT 123.665 0.329 123.96 0.612 ;
      RECT 123.66 0.27 123.69 0.609 ;
      RECT 123.645 0.276 123.78 0.607 ;
      RECT 123.64 0.284 123.865 0.595 ;
      RECT 123.64 0.336 123.975 0.548 ;
      RECT 123.625 0.292 123.865 0.543 ;
      RECT 123.625 0.362 123.985 0.484 ;
      RECT 123.595 0.312 123.95 0.445 ;
      RECT 123.595 0.402 123.995 0.441 ;
      RECT 123.645 0.281 123.865 0.607 ;
      RECT 122.985 0.611 123.04 0.875 ;
      RECT 122.985 0.611 123.105 0.874 ;
      RECT 122.985 0.611 123.13 0.873 ;
      RECT 122.985 0.611 123.195 0.872 ;
      RECT 123.13 0.577 123.21 0.871 ;
      RECT 122.945 0.621 123.355 0.87 ;
      RECT 122.985 0.618 123.355 0.87 ;
      RECT 122.945 0.626 123.36 0.863 ;
      RECT 122.93 0.628 123.36 0.862 ;
      RECT 122.93 0.635 123.365 0.858 ;
      RECT 122.91 0.634 123.36 0.854 ;
      RECT 122.91 0.642 123.37 0.853 ;
      RECT 122.905 0.639 123.365 0.849 ;
      RECT 122.905 0.652 123.38 0.848 ;
      RECT 122.89 0.642 123.37 0.847 ;
      RECT 122.855 0.655 123.38 0.84 ;
      RECT 123.04 0.61 123.35 0.87 ;
      RECT 123.04 0.595 123.3 0.87 ;
      RECT 123.105 0.582 123.235 0.87 ;
      RECT 122.65 1.671 122.665 2.064 ;
      RECT 122.615 1.676 122.665 2.063 ;
      RECT 122.65 1.675 122.71 2.062 ;
      RECT 122.595 1.686 122.71 2.061 ;
      RECT 122.61 1.682 122.71 2.061 ;
      RECT 122.575 1.692 122.785 2.058 ;
      RECT 122.575 1.711 122.83 2.056 ;
      RECT 122.575 1.718 122.835 2.053 ;
      RECT 122.56 1.695 122.785 2.05 ;
      RECT 122.54 1.7 122.785 2.043 ;
      RECT 122.535 1.704 122.785 2.039 ;
      RECT 122.535 1.721 122.845 2.038 ;
      RECT 122.515 1.715 122.83 2.034 ;
      RECT 122.515 1.724 122.85 2.028 ;
      RECT 122.51 1.73 122.85 1.8 ;
      RECT 122.575 1.69 122.71 2.058 ;
      RECT 122.45 1.053 122.65 1.365 ;
      RECT 122.525 1.031 122.65 1.365 ;
      RECT 122.465 1.05 122.655 1.35 ;
      RECT 122.435 1.061 122.655 1.348 ;
      RECT 122.45 1.056 122.66 1.314 ;
      RECT 122.435 1.16 122.665 1.281 ;
      RECT 122.465 1.032 122.65 1.365 ;
      RECT 122.525 1.01 122.625 1.365 ;
      RECT 122.55 1.007 122.625 1.365 ;
      RECT 122.55 1.002 122.57 1.365 ;
      RECT 121.955 1.07 122.13 1.245 ;
      RECT 121.95 1.07 122.13 1.243 ;
      RECT 121.925 1.07 122.13 1.238 ;
      RECT 121.87 1.05 122.04 1.228 ;
      RECT 121.87 1.057 122.105 1.228 ;
      RECT 121.955 1.737 121.97 1.92 ;
      RECT 121.945 1.715 121.955 1.92 ;
      RECT 121.93 1.695 121.945 1.92 ;
      RECT 121.92 1.67 121.93 1.92 ;
      RECT 121.89 1.635 121.92 1.92 ;
      RECT 121.855 1.575 121.89 1.92 ;
      RECT 121.85 1.537 121.855 1.92 ;
      RECT 121.8 1.488 121.85 1.92 ;
      RECT 121.79 1.438 121.8 1.908 ;
      RECT 121.775 1.417 121.79 1.868 ;
      RECT 121.755 1.385 121.775 1.818 ;
      RECT 121.73 1.341 121.755 1.758 ;
      RECT 121.725 1.313 121.73 1.713 ;
      RECT 121.72 1.304 121.725 1.699 ;
      RECT 121.715 1.297 121.72 1.686 ;
      RECT 121.71 1.292 121.715 1.675 ;
      RECT 121.705 1.277 121.71 1.665 ;
      RECT 121.7 1.255 121.705 1.652 ;
      RECT 121.69 1.215 121.7 1.627 ;
      RECT 121.665 1.145 121.69 1.583 ;
      RECT 121.66 1.085 121.665 1.548 ;
      RECT 121.645 1.065 121.66 1.515 ;
      RECT 121.64 1.065 121.645 1.49 ;
      RECT 121.61 1.065 121.64 1.445 ;
      RECT 121.565 1.065 121.61 1.385 ;
      RECT 121.49 1.065 121.565 1.333 ;
      RECT 121.485 1.065 121.49 1.298 ;
      RECT 121.48 1.065 121.485 1.288 ;
      RECT 121.475 1.065 121.48 1.268 ;
      RECT 121.74 0.285 121.91 0.755 ;
      RECT 121.685 0.278 121.88 0.739 ;
      RECT 121.685 0.292 121.915 0.738 ;
      RECT 121.67 0.293 121.915 0.719 ;
      RECT 121.665 0.311 121.915 0.705 ;
      RECT 121.67 0.294 121.92 0.703 ;
      RECT 121.655 0.325 121.92 0.688 ;
      RECT 121.67 0.3 121.925 0.673 ;
      RECT 121.65 0.34 121.925 0.67 ;
      RECT 121.665 0.312 121.93 0.655 ;
      RECT 121.665 0.324 121.935 0.635 ;
      RECT 121.65 0.34 121.94 0.618 ;
      RECT 121.65 0.35 121.945 0.473 ;
      RECT 121.645 0.35 121.945 0.43 ;
      RECT 121.645 0.365 121.95 0.408 ;
      RECT 121.74 0.275 121.88 0.755 ;
      RECT 121.74 0.273 121.85 0.755 ;
      RECT 121.826 0.27 121.85 0.755 ;
      RECT 121.485 1.937 121.49 1.983 ;
      RECT 121.475 1.785 121.485 2.007 ;
      RECT 121.47 1.63 121.475 2.032 ;
      RECT 121.455 1.592 121.47 2.043 ;
      RECT 121.45 1.575 121.455 2.05 ;
      RECT 121.44 1.563 121.45 2.057 ;
      RECT 121.435 1.554 121.44 2.059 ;
      RECT 121.43 1.552 121.435 2.063 ;
      RECT 121.385 1.543 121.43 2.078 ;
      RECT 121.38 1.535 121.385 2.092 ;
      RECT 121.375 1.532 121.38 2.096 ;
      RECT 121.36 1.527 121.375 2.104 ;
      RECT 121.305 1.517 121.36 2.115 ;
      RECT 121.27 1.505 121.305 2.116 ;
      RECT 121.261 1.5 121.27 2.11 ;
      RECT 121.175 1.5 121.261 2.1 ;
      RECT 121.145 1.5 121.175 2.078 ;
      RECT 121.135 1.5 121.14 2.058 ;
      RECT 121.13 1.5 121.135 2.02 ;
      RECT 121.125 1.5 121.13 1.978 ;
      RECT 121.12 1.5 121.125 1.938 ;
      RECT 121.115 1.5 121.12 1.868 ;
      RECT 121.105 1.5 121.115 1.79 ;
      RECT 121.1 1.5 121.105 1.69 ;
      RECT 121.14 1.5 121.145 2.06 ;
      RECT 120.635 1.582 120.725 2.06 ;
      RECT 120.62 1.585 120.74 2.058 ;
      RECT 120.635 1.584 120.74 2.058 ;
      RECT 120.6 1.591 120.765 2.048 ;
      RECT 120.62 1.585 120.765 2.048 ;
      RECT 120.585 1.597 120.765 2.036 ;
      RECT 120.62 1.588 120.815 2.029 ;
      RECT 120.571 1.605 120.815 2.027 ;
      RECT 120.6 1.595 120.825 2.015 ;
      RECT 120.571 1.616 120.855 2.006 ;
      RECT 120.485 1.64 120.855 2 ;
      RECT 120.485 1.653 120.895 1.983 ;
      RECT 120.48 1.675 120.895 1.976 ;
      RECT 120.45 1.69 120.895 1.966 ;
      RECT 120.445 1.701 120.895 1.956 ;
      RECT 120.415 1.714 120.895 1.947 ;
      RECT 120.4 1.732 120.895 1.936 ;
      RECT 120.375 1.745 120.895 1.926 ;
      RECT 120.635 1.581 120.645 2.06 ;
      RECT 120.681 1.005 120.72 1.25 ;
      RECT 120.595 1.005 120.73 1.248 ;
      RECT 120.48 1.03 120.73 1.245 ;
      RECT 120.48 1.03 120.735 1.243 ;
      RECT 120.48 1.03 120.75 1.238 ;
      RECT 120.586 1.005 120.765 1.218 ;
      RECT 120.5 1.013 120.765 1.218 ;
      RECT 120.17 0.365 120.34 0.8 ;
      RECT 120.16 0.399 120.34 0.783 ;
      RECT 120.24 0.335 120.41 0.77 ;
      RECT 120.145 0.41 120.41 0.748 ;
      RECT 120.24 0.345 120.415 0.738 ;
      RECT 120.17 0.397 120.445 0.723 ;
      RECT 120.13 0.423 120.445 0.708 ;
      RECT 120.13 0.465 120.455 0.688 ;
      RECT 120.125 0.49 120.46 0.67 ;
      RECT 120.125 0.5 120.465 0.655 ;
      RECT 120.12 0.437 120.445 0.653 ;
      RECT 120.12 0.51 120.47 0.638 ;
      RECT 120.115 0.447 120.445 0.635 ;
      RECT 120.11 0.531 120.475 0.618 ;
      RECT 120.11 0.563 120.48 0.598 ;
      RECT 120.105 0.477 120.455 0.59 ;
      RECT 120.11 0.462 120.445 0.618 ;
      RECT 120.125 0.432 120.445 0.67 ;
      RECT 119.97 1.019 120.195 1.275 ;
      RECT 119.97 1.052 120.215 1.265 ;
      RECT 119.935 1.052 120.215 1.263 ;
      RECT 119.935 1.065 120.22 1.253 ;
      RECT 119.935 1.085 120.23 1.245 ;
      RECT 119.935 1.182 120.235 1.238 ;
      RECT 119.915 0.93 120.045 1.228 ;
      RECT 119.87 1.085 120.23 1.17 ;
      RECT 119.86 0.93 120.045 1.115 ;
      RECT 119.86 0.962 120.131 1.115 ;
      RECT 119.825 1.492 119.845 1.67 ;
      RECT 119.79 1.445 119.825 1.67 ;
      RECT 119.775 1.385 119.79 1.67 ;
      RECT 119.75 1.332 119.775 1.67 ;
      RECT 119.735 1.285 119.75 1.67 ;
      RECT 119.715 1.262 119.735 1.67 ;
      RECT 119.69 1.227 119.715 1.67 ;
      RECT 119.68 1.073 119.69 1.67 ;
      RECT 119.65 1.068 119.68 1.661 ;
      RECT 119.645 1.065 119.65 1.651 ;
      RECT 119.63 1.065 119.645 1.625 ;
      RECT 119.625 1.065 119.63 1.588 ;
      RECT 119.6 1.065 119.625 1.54 ;
      RECT 119.58 1.065 119.6 1.465 ;
      RECT 119.57 1.065 119.58 1.425 ;
      RECT 119.565 1.065 119.57 1.4 ;
      RECT 119.56 1.065 119.565 1.383 ;
      RECT 119.555 1.065 119.56 1.365 ;
      RECT 119.55 1.066 119.555 1.355 ;
      RECT 119.54 1.068 119.55 1.323 ;
      RECT 119.53 1.07 119.54 1.29 ;
      RECT 119.52 1.073 119.53 1.263 ;
      RECT 119.845 1.5 120.07 1.67 ;
      RECT 119.175 0.312 119.345 0.765 ;
      RECT 119.175 0.312 119.435 0.731 ;
      RECT 119.175 0.312 119.465 0.715 ;
      RECT 119.175 0.312 119.495 0.688 ;
      RECT 119.431 0.29 119.51 0.67 ;
      RECT 119.21 0.297 119.515 0.655 ;
      RECT 119.21 0.305 119.525 0.618 ;
      RECT 119.17 0.332 119.525 0.59 ;
      RECT 119.155 0.345 119.525 0.555 ;
      RECT 119.175 0.32 119.545 0.545 ;
      RECT 119.15 0.385 119.545 0.515 ;
      RECT 119.15 0.415 119.55 0.498 ;
      RECT 119.145 0.445 119.55 0.485 ;
      RECT 119.21 0.294 119.51 0.67 ;
      RECT 119.345 0.291 119.431 0.749 ;
      RECT 119.296 0.292 119.51 0.67 ;
      RECT 119.44 1.952 119.485 2.145 ;
      RECT 119.43 1.922 119.44 2.145 ;
      RECT 119.425 1.907 119.43 2.145 ;
      RECT 119.385 1.817 119.425 2.145 ;
      RECT 119.38 1.73 119.385 2.145 ;
      RECT 119.37 1.7 119.38 2.145 ;
      RECT 119.365 1.66 119.37 2.145 ;
      RECT 119.355 1.622 119.365 2.145 ;
      RECT 119.35 1.587 119.355 2.145 ;
      RECT 119.33 1.54 119.35 2.145 ;
      RECT 119.315 1.465 119.33 2.145 ;
      RECT 119.31 1.42 119.315 2.14 ;
      RECT 119.305 1.4 119.31 2.113 ;
      RECT 119.3 1.38 119.305 2.098 ;
      RECT 119.295 1.355 119.3 2.078 ;
      RECT 119.29 1.333 119.295 2.063 ;
      RECT 119.285 1.311 119.29 2.045 ;
      RECT 119.28 1.29 119.285 2.035 ;
      RECT 119.27 1.262 119.28 2.005 ;
      RECT 119.26 1.225 119.27 1.973 ;
      RECT 119.25 1.185 119.26 1.94 ;
      RECT 119.24 1.163 119.25 1.91 ;
      RECT 119.21 1.115 119.24 1.842 ;
      RECT 119.195 1.075 119.21 1.769 ;
      RECT 119.185 1.075 119.195 1.735 ;
      RECT 119.18 1.075 119.185 1.71 ;
      RECT 119.175 1.075 119.18 1.695 ;
      RECT 119.17 1.075 119.175 1.673 ;
      RECT 119.165 1.075 119.17 1.66 ;
      RECT 119.15 1.075 119.165 1.625 ;
      RECT 119.13 1.075 119.15 1.565 ;
      RECT 119.12 1.075 119.13 1.515 ;
      RECT 119.1 1.075 119.12 1.463 ;
      RECT 119.08 1.075 119.1 1.42 ;
      RECT 119.07 1.075 119.08 1.408 ;
      RECT 119.04 1.075 119.07 1.395 ;
      RECT 119.01 1.096 119.04 1.375 ;
      RECT 119 1.124 119.01 1.355 ;
      RECT 118.985 1.141 119 1.323 ;
      RECT 118.98 1.155 118.985 1.29 ;
      RECT 118.975 1.163 118.98 1.263 ;
      RECT 118.97 1.171 118.975 1.225 ;
      RECT 118.975 1.695 118.98 2.03 ;
      RECT 118.94 1.682 118.975 2.029 ;
      RECT 118.87 1.622 118.94 2.028 ;
      RECT 118.79 1.565 118.87 2.027 ;
      RECT 118.655 1.525 118.79 2.026 ;
      RECT 118.655 1.712 118.99 2.015 ;
      RECT 118.615 1.712 118.99 2.005 ;
      RECT 118.615 1.73 118.995 2 ;
      RECT 118.615 1.82 119 1.99 ;
      RECT 118.61 1.515 118.775 1.97 ;
      RECT 118.605 1.515 118.775 1.713 ;
      RECT 118.605 1.672 118.97 1.713 ;
      RECT 118.605 1.66 118.965 1.713 ;
      RECT 117.87 1.875 118.385 2.285 ;
      RECT 118.045 0.895 118.385 2.285 ;
      RECT 117.155 0.895 118.385 1.065 ;
      RECT 117.865 0.29 118.11 1.065 ;
      RECT 115.265 2.295 117.295 2.465 ;
      RECT 117.125 1.44 117.295 2.465 ;
      RECT 115.265 0.995 115.435 2.465 ;
      RECT 117.125 1.44 117.875 1.63 ;
      RECT 115.24 0.995 115.435 1.325 ;
      RECT 115.945 1.615 116.955 1.785 ;
      RECT 116.765 0.255 116.955 1.785 ;
      RECT 115.945 0.815 116.115 1.785 ;
      RECT 115.605 1.955 116.73 2.125 ;
      RECT 115.605 0.255 115.775 2.125 ;
      RECT 114.76 0.995 115.015 1.325 ;
      RECT 114.845 0.655 115.015 1.325 ;
      RECT 114.845 0.655 115.775 0.825 ;
      RECT 115.6 0.255 115.775 0.825 ;
      RECT 115.6 0.255 116.13 0.62 ;
      RECT 114.42 1.495 114.755 2.465 ;
      RECT 114.42 0.255 114.59 2.465 ;
      RECT 114.42 0.255 114.675 0.825 ;
      RECT 113.67 1.485 114 2.465 ;
      RECT 113.77 0.255 114 2.465 ;
      RECT 113.67 1.815 114.13 1.97 ;
      RECT 113.67 0.255 114 0.885 ;
      RECT 112.29 1.485 112.62 2.465 ;
      RECT 112.39 0.255 112.62 2.465 ;
      RECT 112.39 1.075 113.6 1.315 ;
      RECT 112.29 0.255 112.62 0.885 ;
      RECT 110.91 1.485 111.24 2.465 ;
      RECT 111.01 0.255 111.24 2.465 ;
      RECT 110.91 1.555 111.37 1.725 ;
      RECT 110.91 0.255 111.24 0.885 ;
      RECT 109.53 1.485 109.86 2.465 ;
      RECT 109.63 0.255 109.86 2.465 ;
      RECT 109.63 1.075 110.84 1.315 ;
      RECT 109.53 0.255 109.86 0.885 ;
      RECT 108.21 1.875 108.725 2.285 ;
      RECT 108.385 0.895 108.725 2.285 ;
      RECT 107.495 0.895 108.725 1.065 ;
      RECT 108.205 0.29 108.45 1.065 ;
      RECT 105.605 2.295 107.635 2.465 ;
      RECT 107.465 1.44 107.635 2.465 ;
      RECT 105.605 0.995 105.775 2.465 ;
      RECT 107.465 1.44 108.215 1.63 ;
      RECT 105.58 0.995 105.775 1.325 ;
      RECT 106.285 1.615 107.295 1.785 ;
      RECT 107.105 0.255 107.295 1.785 ;
      RECT 106.285 0.815 106.455 1.785 ;
      RECT 105.945 1.955 107.07 2.125 ;
      RECT 105.945 0.255 106.115 2.125 ;
      RECT 105.1 0.995 105.355 1.325 ;
      RECT 105.185 0.655 105.355 1.325 ;
      RECT 105.185 0.655 106.115 0.825 ;
      RECT 105.94 0.255 106.115 0.825 ;
      RECT 105.94 0.255 106.47 0.62 ;
      RECT 104.76 1.495 105.095 2.465 ;
      RECT 104.76 0.255 104.93 2.465 ;
      RECT 104.76 0.255 105.015 0.825 ;
      RECT 104.075 1.875 104.59 2.285 ;
      RECT 104.25 0.895 104.59 2.285 ;
      RECT 103.36 0.895 104.59 1.065 ;
      RECT 104.07 0.29 104.315 1.065 ;
      RECT 101.47 2.295 103.5 2.465 ;
      RECT 103.33 1.44 103.5 2.465 ;
      RECT 101.47 0.995 101.64 2.465 ;
      RECT 103.33 1.44 104.08 1.63 ;
      RECT 101.445 0.995 101.64 1.325 ;
      RECT 102.15 1.615 103.16 1.785 ;
      RECT 102.97 0.255 103.16 1.785 ;
      RECT 102.15 0.815 102.32 1.785 ;
      RECT 101.81 1.955 102.935 2.125 ;
      RECT 101.81 0.255 101.98 2.125 ;
      RECT 100.965 0.995 101.22 1.325 ;
      RECT 101.05 0.655 101.22 1.325 ;
      RECT 101.05 0.655 101.98 0.825 ;
      RECT 101.805 0.255 101.98 0.825 ;
      RECT 101.805 0.255 102.335 0.62 ;
      RECT 100.625 1.495 100.96 2.465 ;
      RECT 100.625 0.255 100.795 2.465 ;
      RECT 100.625 0.255 100.88 0.825 ;
      RECT 99.53 0.475 100.26 0.715 ;
      RECT 100.072 0.27 100.26 0.715 ;
      RECT 99.9 0.282 100.275 0.709 ;
      RECT 99.815 0.297 100.295 0.694 ;
      RECT 99.815 0.312 100.3 0.684 ;
      RECT 99.77 0.332 100.315 0.676 ;
      RECT 99.747 0.367 100.33 0.63 ;
      RECT 99.661 0.39 100.335 0.59 ;
      RECT 99.661 0.408 100.345 0.56 ;
      RECT 99.53 0.477 100.35 0.523 ;
      RECT 99.575 0.42 100.345 0.56 ;
      RECT 99.661 0.372 100.33 0.63 ;
      RECT 99.747 0.341 100.315 0.676 ;
      RECT 99.77 0.322 100.3 0.684 ;
      RECT 99.815 0.295 100.275 0.709 ;
      RECT 99.9 0.277 100.26 0.715 ;
      RECT 99.986 0.271 100.26 0.715 ;
      RECT 100.072 0.266 100.205 0.715 ;
      RECT 100.158 0.261 100.205 0.715 ;
      RECT 99.85 1.159 100.02 1.545 ;
      RECT 99.845 1.159 100.02 1.54 ;
      RECT 99.82 1.159 100.02 1.505 ;
      RECT 99.82 1.187 100.03 1.495 ;
      RECT 99.8 1.187 100.03 1.455 ;
      RECT 99.795 1.187 100.03 1.428 ;
      RECT 99.795 1.205 100.035 1.42 ;
      RECT 99.74 1.205 100.035 1.355 ;
      RECT 99.74 1.222 100.045 1.338 ;
      RECT 99.73 1.222 100.045 1.278 ;
      RECT 99.73 1.239 100.05 1.275 ;
      RECT 99.725 1.075 99.895 1.253 ;
      RECT 99.725 1.109 99.981 1.253 ;
      RECT 99.72 1.875 99.725 1.888 ;
      RECT 99.715 1.77 99.72 1.893 ;
      RECT 99.69 1.63 99.715 1.908 ;
      RECT 99.655 1.581 99.69 1.94 ;
      RECT 99.65 1.549 99.655 1.96 ;
      RECT 99.645 1.54 99.65 1.96 ;
      RECT 99.565 1.505 99.645 1.96 ;
      RECT 99.502 1.475 99.565 1.96 ;
      RECT 99.416 1.463 99.502 1.96 ;
      RECT 99.33 1.449 99.416 1.96 ;
      RECT 99.25 1.436 99.33 1.946 ;
      RECT 99.215 1.428 99.25 1.926 ;
      RECT 99.205 1.425 99.215 1.917 ;
      RECT 99.175 1.42 99.205 1.904 ;
      RECT 99.125 1.395 99.175 1.88 ;
      RECT 99.111 1.369 99.125 1.862 ;
      RECT 99.025 1.329 99.111 1.838 ;
      RECT 98.98 1.277 99.025 1.807 ;
      RECT 98.97 1.252 98.98 1.794 ;
      RECT 98.965 1.033 98.97 1.055 ;
      RECT 98.96 1.235 98.97 1.79 ;
      RECT 98.96 1.031 98.965 1.145 ;
      RECT 98.95 1.027 98.96 1.786 ;
      RECT 98.906 1.025 98.95 1.774 ;
      RECT 98.82 1.025 98.906 1.745 ;
      RECT 98.79 1.025 98.82 1.718 ;
      RECT 98.775 1.025 98.79 1.706 ;
      RECT 98.735 1.037 98.775 1.691 ;
      RECT 98.715 1.056 98.735 1.67 ;
      RECT 98.705 1.066 98.715 1.654 ;
      RECT 98.695 1.072 98.705 1.643 ;
      RECT 98.675 1.082 98.695 1.626 ;
      RECT 98.67 1.091 98.675 1.613 ;
      RECT 98.665 1.095 98.67 1.563 ;
      RECT 98.655 1.101 98.665 1.48 ;
      RECT 98.65 1.105 98.655 1.394 ;
      RECT 98.645 1.125 98.65 1.331 ;
      RECT 98.64 1.148 98.645 1.278 ;
      RECT 98.635 1.166 98.64 1.223 ;
      RECT 99.245 0.985 99.415 1.245 ;
      RECT 99.415 0.95 99.46 1.231 ;
      RECT 99.376 0.952 99.465 1.214 ;
      RECT 99.265 0.969 99.551 1.185 ;
      RECT 99.265 0.984 99.555 1.157 ;
      RECT 99.265 0.965 99.465 1.214 ;
      RECT 99.29 0.953 99.415 1.245 ;
      RECT 99.376 0.951 99.46 1.231 ;
      RECT 98.43 0.34 98.6 0.83 ;
      RECT 98.43 0.34 98.635 0.81 ;
      RECT 98.565 0.26 98.675 0.77 ;
      RECT 98.546 0.264 98.695 0.74 ;
      RECT 98.46 0.272 98.715 0.723 ;
      RECT 98.46 0.278 98.72 0.713 ;
      RECT 98.46 0.287 98.74 0.701 ;
      RECT 98.435 0.312 98.77 0.679 ;
      RECT 98.435 0.332 98.775 0.659 ;
      RECT 98.43 0.345 98.785 0.639 ;
      RECT 98.43 0.412 98.79 0.62 ;
      RECT 98.43 0.545 98.795 0.607 ;
      RECT 98.425 0.35 98.785 0.44 ;
      RECT 98.435 0.307 98.74 0.701 ;
      RECT 98.546 0.262 98.675 0.77 ;
      RECT 98.42 2.015 98.72 2.27 ;
      RECT 98.505 1.981 98.72 2.27 ;
      RECT 98.505 1.984 98.725 2.13 ;
      RECT 98.44 2.005 98.725 2.13 ;
      RECT 98.475 1.995 98.72 2.27 ;
      RECT 98.47 2 98.725 2.13 ;
      RECT 98.505 1.979 98.706 2.27 ;
      RECT 98.591 1.97 98.706 2.27 ;
      RECT 98.591 1.964 98.62 2.27 ;
      RECT 98.08 1.605 98.09 2.095 ;
      RECT 97.74 1.54 97.75 1.84 ;
      RECT 98.255 1.712 98.26 1.931 ;
      RECT 98.245 1.692 98.255 1.948 ;
      RECT 98.235 1.672 98.245 1.978 ;
      RECT 98.23 1.662 98.235 1.993 ;
      RECT 98.225 1.658 98.23 1.998 ;
      RECT 98.21 1.65 98.225 2.005 ;
      RECT 98.17 1.63 98.21 2.03 ;
      RECT 98.145 1.612 98.17 2.063 ;
      RECT 98.14 1.61 98.145 2.076 ;
      RECT 98.12 1.607 98.14 2.08 ;
      RECT 98.09 1.605 98.12 2.09 ;
      RECT 98.02 1.607 98.08 2.091 ;
      RECT 98 1.607 98.02 2.085 ;
      RECT 97.975 1.605 98 2.082 ;
      RECT 97.94 1.6 97.975 2.078 ;
      RECT 97.92 1.594 97.94 2.065 ;
      RECT 97.91 1.591 97.92 2.053 ;
      RECT 97.89 1.588 97.91 2.038 ;
      RECT 97.87 1.584 97.89 2.02 ;
      RECT 97.865 1.581 97.87 2.01 ;
      RECT 97.86 1.58 97.865 2.008 ;
      RECT 97.85 1.577 97.86 2 ;
      RECT 97.84 1.571 97.85 1.983 ;
      RECT 97.83 1.565 97.84 1.965 ;
      RECT 97.82 1.559 97.83 1.953 ;
      RECT 97.81 1.553 97.82 1.933 ;
      RECT 97.805 1.549 97.81 1.918 ;
      RECT 97.8 1.547 97.805 1.91 ;
      RECT 97.795 1.545 97.8 1.903 ;
      RECT 97.79 1.543 97.795 1.893 ;
      RECT 97.785 1.541 97.79 1.887 ;
      RECT 97.775 1.54 97.785 1.877 ;
      RECT 97.765 1.54 97.775 1.868 ;
      RECT 97.75 1.54 97.765 1.853 ;
      RECT 97.71 1.54 97.74 1.837 ;
      RECT 97.69 1.542 97.71 1.832 ;
      RECT 97.685 1.547 97.69 1.83 ;
      RECT 97.655 1.555 97.685 1.828 ;
      RECT 97.625 1.57 97.655 1.827 ;
      RECT 97.58 1.592 97.625 1.832 ;
      RECT 97.575 1.607 97.58 1.836 ;
      RECT 97.56 1.612 97.575 1.838 ;
      RECT 97.555 1.616 97.56 1.84 ;
      RECT 97.495 1.639 97.555 1.849 ;
      RECT 97.475 1.665 97.495 1.862 ;
      RECT 97.465 1.672 97.475 1.866 ;
      RECT 97.45 1.679 97.465 1.869 ;
      RECT 97.43 1.689 97.45 1.872 ;
      RECT 97.425 1.697 97.43 1.875 ;
      RECT 97.38 1.702 97.425 1.882 ;
      RECT 97.37 1.705 97.38 1.889 ;
      RECT 97.36 1.705 97.37 1.893 ;
      RECT 97.325 1.707 97.36 1.905 ;
      RECT 97.305 1.71 97.325 1.918 ;
      RECT 97.265 1.713 97.305 1.929 ;
      RECT 97.25 1.715 97.265 1.942 ;
      RECT 97.24 1.715 97.25 1.947 ;
      RECT 97.215 1.716 97.24 1.955 ;
      RECT 97.205 1.718 97.215 1.96 ;
      RECT 97.2 1.719 97.205 1.963 ;
      RECT 97.175 1.717 97.2 1.966 ;
      RECT 97.16 1.715 97.175 1.967 ;
      RECT 97.14 1.712 97.16 1.969 ;
      RECT 97.12 1.707 97.14 1.969 ;
      RECT 97.06 1.702 97.12 1.966 ;
      RECT 97.025 1.677 97.06 1.962 ;
      RECT 97.015 1.654 97.025 1.96 ;
      RECT 96.985 1.631 97.015 1.96 ;
      RECT 96.975 1.61 96.985 1.96 ;
      RECT 96.95 1.592 96.975 1.958 ;
      RECT 96.935 1.57 96.95 1.955 ;
      RECT 96.92 1.552 96.935 1.953 ;
      RECT 96.9 1.542 96.92 1.951 ;
      RECT 96.885 1.537 96.9 1.95 ;
      RECT 96.87 1.535 96.885 1.949 ;
      RECT 96.84 1.536 96.87 1.947 ;
      RECT 96.82 1.539 96.84 1.945 ;
      RECT 96.763 1.543 96.82 1.945 ;
      RECT 96.677 1.552 96.763 1.945 ;
      RECT 96.591 1.563 96.677 1.945 ;
      RECT 96.505 1.574 96.591 1.945 ;
      RECT 96.485 1.581 96.505 1.953 ;
      RECT 96.475 1.584 96.485 1.96 ;
      RECT 96.41 1.589 96.475 1.978 ;
      RECT 96.38 1.596 96.41 2.003 ;
      RECT 96.37 1.599 96.38 2.01 ;
      RECT 96.325 1.603 96.37 2.015 ;
      RECT 96.295 1.608 96.325 2.02 ;
      RECT 96.294 1.61 96.295 2.02 ;
      RECT 96.208 1.616 96.294 2.02 ;
      RECT 96.122 1.627 96.208 2.02 ;
      RECT 96.036 1.639 96.122 2.02 ;
      RECT 95.95 1.65 96.036 2.02 ;
      RECT 95.935 1.657 95.95 2.015 ;
      RECT 95.93 1.659 95.935 2.009 ;
      RECT 95.91 1.67 95.93 2.004 ;
      RECT 95.9 1.688 95.91 1.998 ;
      RECT 95.895 1.7 95.9 1.798 ;
      RECT 98.19 0.453 98.21 0.54 ;
      RECT 98.185 0.388 98.19 0.572 ;
      RECT 98.175 0.355 98.185 0.577 ;
      RECT 98.17 0.335 98.175 0.583 ;
      RECT 98.14 0.335 98.17 0.6 ;
      RECT 98.091 0.335 98.14 0.636 ;
      RECT 98.005 0.335 98.091 0.694 ;
      RECT 97.976 0.345 98.005 0.743 ;
      RECT 97.89 0.387 97.976 0.796 ;
      RECT 97.87 0.425 97.89 0.843 ;
      RECT 97.845 0.442 97.87 0.863 ;
      RECT 97.835 0.456 97.845 0.883 ;
      RECT 97.83 0.462 97.835 0.893 ;
      RECT 97.825 0.466 97.83 0.9 ;
      RECT 97.775 0.486 97.825 0.905 ;
      RECT 97.71 0.53 97.775 0.905 ;
      RECT 97.685 0.58 97.71 0.905 ;
      RECT 97.675 0.61 97.685 0.905 ;
      RECT 97.67 0.637 97.675 0.905 ;
      RECT 97.665 0.655 97.67 0.905 ;
      RECT 97.655 0.697 97.665 0.905 ;
      RECT 98.005 1.255 98.175 1.43 ;
      RECT 97.945 1.083 98.005 1.418 ;
      RECT 97.935 1.076 97.945 1.401 ;
      RECT 97.89 1.255 98.175 1.381 ;
      RECT 97.871 1.255 98.175 1.359 ;
      RECT 97.785 1.255 98.175 1.324 ;
      RECT 97.765 1.075 97.935 1.28 ;
      RECT 97.765 1.222 98.17 1.28 ;
      RECT 97.765 1.17 98.145 1.28 ;
      RECT 97.765 1.125 98.11 1.28 ;
      RECT 97.765 1.107 98.075 1.28 ;
      RECT 97.765 1.097 98.07 1.28 ;
      RECT 97.485 2.055 97.675 2.28 ;
      RECT 97.475 2.056 97.68 2.275 ;
      RECT 97.475 2.058 97.69 2.255 ;
      RECT 97.475 2.062 97.695 2.24 ;
      RECT 97.475 2.049 97.645 2.275 ;
      RECT 97.475 2.052 97.67 2.275 ;
      RECT 97.485 2.048 97.645 2.28 ;
      RECT 97.571 2.046 97.645 2.28 ;
      RECT 97.195 1.297 97.365 1.535 ;
      RECT 97.195 1.297 97.451 1.449 ;
      RECT 97.195 1.297 97.455 1.359 ;
      RECT 97.245 1.07 97.465 1.338 ;
      RECT 97.24 1.087 97.47 1.311 ;
      RECT 97.205 1.245 97.47 1.311 ;
      RECT 97.225 1.095 97.365 1.535 ;
      RECT 97.215 1.177 97.475 1.294 ;
      RECT 97.21 1.225 97.475 1.294 ;
      RECT 97.215 1.135 97.47 1.311 ;
      RECT 97.24 1.072 97.465 1.338 ;
      RECT 96.805 1.047 96.975 1.245 ;
      RECT 96.805 1.047 97.02 1.22 ;
      RECT 96.875 0.99 97.045 1.178 ;
      RECT 96.85 1.005 97.045 1.178 ;
      RECT 96.465 1.051 96.495 1.245 ;
      RECT 96.46 1.023 96.465 1.245 ;
      RECT 96.43 0.997 96.46 1.247 ;
      RECT 96.405 0.955 96.43 1.25 ;
      RECT 96.395 0.927 96.405 1.252 ;
      RECT 96.36 0.907 96.395 1.254 ;
      RECT 96.295 0.892 96.36 1.26 ;
      RECT 96.245 0.89 96.295 1.266 ;
      RECT 96.222 0.892 96.245 1.271 ;
      RECT 96.136 0.903 96.222 1.277 ;
      RECT 96.05 0.921 96.136 1.287 ;
      RECT 96.035 0.932 96.05 1.293 ;
      RECT 95.965 0.955 96.035 1.299 ;
      RECT 95.91 0.987 95.965 1.307 ;
      RECT 95.87 1.01 95.91 1.313 ;
      RECT 95.856 1.023 95.87 1.316 ;
      RECT 95.77 1.045 95.856 1.322 ;
      RECT 95.755 1.07 95.77 1.328 ;
      RECT 95.715 1.085 95.755 1.332 ;
      RECT 95.665 1.1 95.715 1.337 ;
      RECT 95.64 1.107 95.665 1.341 ;
      RECT 95.58 1.102 95.64 1.345 ;
      RECT 95.565 1.093 95.58 1.349 ;
      RECT 95.495 1.083 95.565 1.345 ;
      RECT 95.47 1.075 95.49 1.335 ;
      RECT 95.411 1.075 95.47 1.313 ;
      RECT 95.325 1.075 95.411 1.27 ;
      RECT 95.49 1.075 95.495 1.34 ;
      RECT 96.185 0.306 96.355 0.64 ;
      RECT 96.155 0.306 96.355 0.635 ;
      RECT 96.095 0.273 96.155 0.623 ;
      RECT 96.095 0.329 96.365 0.618 ;
      RECT 96.07 0.329 96.365 0.612 ;
      RECT 96.065 0.27 96.095 0.609 ;
      RECT 96.05 0.276 96.185 0.607 ;
      RECT 96.045 0.284 96.27 0.595 ;
      RECT 96.045 0.336 96.38 0.548 ;
      RECT 96.03 0.292 96.27 0.543 ;
      RECT 96.03 0.362 96.39 0.484 ;
      RECT 96 0.312 96.355 0.445 ;
      RECT 96 0.402 96.4 0.441 ;
      RECT 96.05 0.281 96.27 0.607 ;
      RECT 95.39 0.611 95.445 0.875 ;
      RECT 95.39 0.611 95.51 0.874 ;
      RECT 95.39 0.611 95.535 0.873 ;
      RECT 95.39 0.611 95.6 0.872 ;
      RECT 95.535 0.577 95.615 0.871 ;
      RECT 95.35 0.621 95.76 0.87 ;
      RECT 95.39 0.618 95.76 0.87 ;
      RECT 95.35 0.626 95.765 0.863 ;
      RECT 95.335 0.628 95.765 0.862 ;
      RECT 95.335 0.635 95.77 0.858 ;
      RECT 95.315 0.634 95.765 0.854 ;
      RECT 95.315 0.642 95.775 0.853 ;
      RECT 95.31 0.639 95.77 0.849 ;
      RECT 95.31 0.652 95.785 0.848 ;
      RECT 95.295 0.642 95.775 0.847 ;
      RECT 95.26 0.655 95.785 0.84 ;
      RECT 95.445 0.61 95.755 0.87 ;
      RECT 95.445 0.595 95.705 0.87 ;
      RECT 95.51 0.582 95.64 0.87 ;
      RECT 95.055 1.671 95.07 2.064 ;
      RECT 95.02 1.676 95.07 2.063 ;
      RECT 95.055 1.675 95.115 2.062 ;
      RECT 95 1.686 95.115 2.061 ;
      RECT 95.015 1.682 95.115 2.061 ;
      RECT 94.98 1.692 95.19 2.058 ;
      RECT 94.98 1.711 95.235 2.056 ;
      RECT 94.98 1.718 95.24 2.053 ;
      RECT 94.965 1.695 95.19 2.05 ;
      RECT 94.945 1.7 95.19 2.043 ;
      RECT 94.94 1.704 95.19 2.039 ;
      RECT 94.94 1.721 95.25 2.038 ;
      RECT 94.92 1.715 95.235 2.034 ;
      RECT 94.92 1.724 95.255 2.028 ;
      RECT 94.915 1.73 95.255 1.8 ;
      RECT 94.98 1.69 95.115 2.058 ;
      RECT 94.855 1.053 95.055 1.365 ;
      RECT 94.93 1.031 95.055 1.365 ;
      RECT 94.87 1.05 95.06 1.35 ;
      RECT 94.84 1.061 95.06 1.348 ;
      RECT 94.855 1.056 95.065 1.314 ;
      RECT 94.84 1.16 95.07 1.281 ;
      RECT 94.87 1.032 95.055 1.365 ;
      RECT 94.93 1.01 95.03 1.365 ;
      RECT 94.955 1.007 95.03 1.365 ;
      RECT 94.955 1.002 94.975 1.365 ;
      RECT 94.36 1.07 94.535 1.245 ;
      RECT 94.355 1.07 94.535 1.243 ;
      RECT 94.33 1.07 94.535 1.238 ;
      RECT 94.275 1.05 94.445 1.228 ;
      RECT 94.275 1.057 94.51 1.228 ;
      RECT 94.36 1.737 94.375 1.92 ;
      RECT 94.35 1.715 94.36 1.92 ;
      RECT 94.335 1.695 94.35 1.92 ;
      RECT 94.325 1.67 94.335 1.92 ;
      RECT 94.295 1.635 94.325 1.92 ;
      RECT 94.26 1.575 94.295 1.92 ;
      RECT 94.255 1.537 94.26 1.92 ;
      RECT 94.205 1.488 94.255 1.92 ;
      RECT 94.195 1.438 94.205 1.908 ;
      RECT 94.18 1.417 94.195 1.868 ;
      RECT 94.16 1.385 94.18 1.818 ;
      RECT 94.135 1.341 94.16 1.758 ;
      RECT 94.13 1.313 94.135 1.713 ;
      RECT 94.125 1.304 94.13 1.699 ;
      RECT 94.12 1.297 94.125 1.686 ;
      RECT 94.115 1.292 94.12 1.675 ;
      RECT 94.11 1.277 94.115 1.665 ;
      RECT 94.105 1.255 94.11 1.652 ;
      RECT 94.095 1.215 94.105 1.627 ;
      RECT 94.07 1.145 94.095 1.583 ;
      RECT 94.065 1.085 94.07 1.548 ;
      RECT 94.05 1.065 94.065 1.515 ;
      RECT 94.045 1.065 94.05 1.49 ;
      RECT 94.015 1.065 94.045 1.445 ;
      RECT 93.97 1.065 94.015 1.385 ;
      RECT 93.895 1.065 93.97 1.333 ;
      RECT 93.89 1.065 93.895 1.298 ;
      RECT 93.885 1.065 93.89 1.288 ;
      RECT 93.88 1.065 93.885 1.268 ;
      RECT 94.145 0.285 94.315 0.755 ;
      RECT 94.09 0.278 94.285 0.739 ;
      RECT 94.09 0.292 94.32 0.738 ;
      RECT 94.075 0.293 94.32 0.719 ;
      RECT 94.07 0.311 94.32 0.705 ;
      RECT 94.075 0.294 94.325 0.703 ;
      RECT 94.06 0.325 94.325 0.688 ;
      RECT 94.075 0.3 94.33 0.673 ;
      RECT 94.055 0.34 94.33 0.67 ;
      RECT 94.07 0.312 94.335 0.655 ;
      RECT 94.07 0.324 94.34 0.635 ;
      RECT 94.055 0.34 94.345 0.618 ;
      RECT 94.055 0.35 94.35 0.473 ;
      RECT 94.05 0.35 94.35 0.43 ;
      RECT 94.05 0.365 94.355 0.408 ;
      RECT 94.145 0.275 94.285 0.755 ;
      RECT 94.145 0.273 94.255 0.755 ;
      RECT 94.231 0.27 94.255 0.755 ;
      RECT 93.89 1.937 93.895 1.983 ;
      RECT 93.88 1.785 93.89 2.007 ;
      RECT 93.875 1.63 93.88 2.032 ;
      RECT 93.86 1.592 93.875 2.043 ;
      RECT 93.855 1.575 93.86 2.05 ;
      RECT 93.845 1.563 93.855 2.057 ;
      RECT 93.84 1.554 93.845 2.059 ;
      RECT 93.835 1.552 93.84 2.063 ;
      RECT 93.79 1.543 93.835 2.078 ;
      RECT 93.785 1.535 93.79 2.092 ;
      RECT 93.78 1.532 93.785 2.096 ;
      RECT 93.765 1.527 93.78 2.104 ;
      RECT 93.71 1.517 93.765 2.115 ;
      RECT 93.675 1.505 93.71 2.116 ;
      RECT 93.666 1.5 93.675 2.11 ;
      RECT 93.58 1.5 93.666 2.1 ;
      RECT 93.55 1.5 93.58 2.078 ;
      RECT 93.54 1.5 93.545 2.058 ;
      RECT 93.535 1.5 93.54 2.02 ;
      RECT 93.53 1.5 93.535 1.978 ;
      RECT 93.525 1.5 93.53 1.938 ;
      RECT 93.52 1.5 93.525 1.868 ;
      RECT 93.51 1.5 93.52 1.79 ;
      RECT 93.505 1.5 93.51 1.69 ;
      RECT 93.545 1.5 93.55 2.06 ;
      RECT 93.04 1.582 93.13 2.06 ;
      RECT 93.025 1.585 93.145 2.058 ;
      RECT 93.04 1.584 93.145 2.058 ;
      RECT 93.005 1.591 93.17 2.048 ;
      RECT 93.025 1.585 93.17 2.048 ;
      RECT 92.99 1.597 93.17 2.036 ;
      RECT 93.025 1.588 93.22 2.029 ;
      RECT 92.976 1.605 93.22 2.027 ;
      RECT 93.005 1.595 93.23 2.015 ;
      RECT 92.976 1.616 93.26 2.006 ;
      RECT 92.89 1.64 93.26 2 ;
      RECT 92.89 1.653 93.3 1.983 ;
      RECT 92.885 1.675 93.3 1.976 ;
      RECT 92.855 1.69 93.3 1.966 ;
      RECT 92.85 1.701 93.3 1.956 ;
      RECT 92.82 1.714 93.3 1.947 ;
      RECT 92.805 1.732 93.3 1.936 ;
      RECT 92.78 1.745 93.3 1.926 ;
      RECT 93.04 1.581 93.05 2.06 ;
      RECT 93.086 1.005 93.125 1.25 ;
      RECT 93 1.005 93.135 1.248 ;
      RECT 92.885 1.03 93.135 1.245 ;
      RECT 92.885 1.03 93.14 1.243 ;
      RECT 92.885 1.03 93.155 1.238 ;
      RECT 92.991 1.005 93.17 1.218 ;
      RECT 92.905 1.013 93.17 1.218 ;
      RECT 92.575 0.365 92.745 0.8 ;
      RECT 92.565 0.399 92.745 0.783 ;
      RECT 92.645 0.335 92.815 0.77 ;
      RECT 92.55 0.41 92.815 0.748 ;
      RECT 92.645 0.345 92.82 0.738 ;
      RECT 92.575 0.397 92.85 0.723 ;
      RECT 92.535 0.423 92.85 0.708 ;
      RECT 92.535 0.465 92.86 0.688 ;
      RECT 92.53 0.49 92.865 0.67 ;
      RECT 92.53 0.5 92.87 0.655 ;
      RECT 92.525 0.437 92.85 0.653 ;
      RECT 92.525 0.51 92.875 0.638 ;
      RECT 92.52 0.447 92.85 0.635 ;
      RECT 92.515 0.531 92.88 0.618 ;
      RECT 92.515 0.563 92.885 0.598 ;
      RECT 92.51 0.477 92.86 0.59 ;
      RECT 92.515 0.462 92.85 0.618 ;
      RECT 92.53 0.432 92.85 0.67 ;
      RECT 92.375 1.019 92.6 1.275 ;
      RECT 92.375 1.052 92.62 1.265 ;
      RECT 92.34 1.052 92.62 1.263 ;
      RECT 92.34 1.065 92.625 1.253 ;
      RECT 92.34 1.085 92.635 1.245 ;
      RECT 92.34 1.182 92.64 1.238 ;
      RECT 92.32 0.93 92.45 1.228 ;
      RECT 92.275 1.085 92.635 1.17 ;
      RECT 92.265 0.93 92.45 1.115 ;
      RECT 92.265 0.962 92.536 1.115 ;
      RECT 92.23 1.492 92.25 1.67 ;
      RECT 92.195 1.445 92.23 1.67 ;
      RECT 92.18 1.385 92.195 1.67 ;
      RECT 92.155 1.332 92.18 1.67 ;
      RECT 92.14 1.285 92.155 1.67 ;
      RECT 92.12 1.262 92.14 1.67 ;
      RECT 92.095 1.227 92.12 1.67 ;
      RECT 92.085 1.073 92.095 1.67 ;
      RECT 92.055 1.068 92.085 1.661 ;
      RECT 92.05 1.065 92.055 1.651 ;
      RECT 92.035 1.065 92.05 1.625 ;
      RECT 92.03 1.065 92.035 1.588 ;
      RECT 92.005 1.065 92.03 1.54 ;
      RECT 91.985 1.065 92.005 1.465 ;
      RECT 91.975 1.065 91.985 1.425 ;
      RECT 91.97 1.065 91.975 1.4 ;
      RECT 91.965 1.065 91.97 1.383 ;
      RECT 91.96 1.065 91.965 1.365 ;
      RECT 91.955 1.066 91.96 1.355 ;
      RECT 91.945 1.068 91.955 1.323 ;
      RECT 91.935 1.07 91.945 1.29 ;
      RECT 91.925 1.073 91.935 1.263 ;
      RECT 92.25 1.5 92.475 1.67 ;
      RECT 91.58 0.312 91.75 0.765 ;
      RECT 91.58 0.312 91.84 0.731 ;
      RECT 91.58 0.312 91.87 0.715 ;
      RECT 91.58 0.312 91.9 0.688 ;
      RECT 91.836 0.29 91.915 0.67 ;
      RECT 91.615 0.297 91.92 0.655 ;
      RECT 91.615 0.305 91.93 0.618 ;
      RECT 91.575 0.332 91.93 0.59 ;
      RECT 91.56 0.345 91.93 0.555 ;
      RECT 91.58 0.32 91.95 0.545 ;
      RECT 91.555 0.385 91.95 0.515 ;
      RECT 91.555 0.415 91.955 0.498 ;
      RECT 91.55 0.445 91.955 0.485 ;
      RECT 91.615 0.294 91.915 0.67 ;
      RECT 91.75 0.291 91.836 0.749 ;
      RECT 91.701 0.292 91.915 0.67 ;
      RECT 91.845 1.952 91.89 2.145 ;
      RECT 91.835 1.922 91.845 2.145 ;
      RECT 91.83 1.907 91.835 2.145 ;
      RECT 91.79 1.817 91.83 2.145 ;
      RECT 91.785 1.73 91.79 2.145 ;
      RECT 91.775 1.7 91.785 2.145 ;
      RECT 91.77 1.66 91.775 2.145 ;
      RECT 91.76 1.622 91.77 2.145 ;
      RECT 91.755 1.587 91.76 2.145 ;
      RECT 91.735 1.54 91.755 2.145 ;
      RECT 91.72 1.465 91.735 2.145 ;
      RECT 91.715 1.42 91.72 2.14 ;
      RECT 91.71 1.4 91.715 2.113 ;
      RECT 91.705 1.38 91.71 2.098 ;
      RECT 91.7 1.355 91.705 2.078 ;
      RECT 91.695 1.333 91.7 2.063 ;
      RECT 91.69 1.311 91.695 2.045 ;
      RECT 91.685 1.29 91.69 2.035 ;
      RECT 91.675 1.262 91.685 2.005 ;
      RECT 91.665 1.225 91.675 1.973 ;
      RECT 91.655 1.185 91.665 1.94 ;
      RECT 91.645 1.163 91.655 1.91 ;
      RECT 91.615 1.115 91.645 1.842 ;
      RECT 91.6 1.075 91.615 1.769 ;
      RECT 91.59 1.075 91.6 1.735 ;
      RECT 91.585 1.075 91.59 1.71 ;
      RECT 91.58 1.075 91.585 1.695 ;
      RECT 91.575 1.075 91.58 1.673 ;
      RECT 91.57 1.075 91.575 1.66 ;
      RECT 91.555 1.075 91.57 1.625 ;
      RECT 91.535 1.075 91.555 1.565 ;
      RECT 91.525 1.075 91.535 1.515 ;
      RECT 91.505 1.075 91.525 1.463 ;
      RECT 91.485 1.075 91.505 1.42 ;
      RECT 91.475 1.075 91.485 1.408 ;
      RECT 91.445 1.075 91.475 1.395 ;
      RECT 91.415 1.096 91.445 1.375 ;
      RECT 91.405 1.124 91.415 1.355 ;
      RECT 91.39 1.141 91.405 1.323 ;
      RECT 91.385 1.155 91.39 1.29 ;
      RECT 91.38 1.163 91.385 1.263 ;
      RECT 91.375 1.171 91.38 1.225 ;
      RECT 91.38 1.695 91.385 2.03 ;
      RECT 91.345 1.682 91.38 2.029 ;
      RECT 91.275 1.622 91.345 2.028 ;
      RECT 91.195 1.565 91.275 2.027 ;
      RECT 91.06 1.525 91.195 2.026 ;
      RECT 91.06 1.712 91.395 2.015 ;
      RECT 91.02 1.712 91.395 2.005 ;
      RECT 91.02 1.73 91.4 2 ;
      RECT 91.02 1.82 91.405 1.99 ;
      RECT 91.015 1.515 91.18 1.97 ;
      RECT 91.01 1.515 91.18 1.713 ;
      RECT 91.01 1.672 91.375 1.713 ;
      RECT 91.01 1.66 91.37 1.713 ;
      RECT 90.275 1.875 90.79 2.285 ;
      RECT 90.45 0.895 90.79 2.285 ;
      RECT 89.56 0.895 90.79 1.065 ;
      RECT 90.27 0.29 90.515 1.065 ;
      RECT 87.67 2.295 89.7 2.465 ;
      RECT 89.53 1.44 89.7 2.465 ;
      RECT 87.67 0.995 87.84 2.465 ;
      RECT 89.53 1.44 90.28 1.63 ;
      RECT 87.645 0.995 87.84 1.325 ;
      RECT 88.35 1.615 89.36 1.785 ;
      RECT 89.17 0.255 89.36 1.785 ;
      RECT 88.35 0.815 88.52 1.785 ;
      RECT 88.01 1.955 89.135 2.125 ;
      RECT 88.01 0.255 88.18 2.125 ;
      RECT 87.165 0.995 87.42 1.325 ;
      RECT 87.25 0.655 87.42 1.325 ;
      RECT 87.25 0.655 88.18 0.825 ;
      RECT 88.005 0.255 88.18 0.825 ;
      RECT 88.005 0.255 88.535 0.62 ;
      RECT 86.825 1.495 87.16 2.465 ;
      RECT 86.825 0.255 86.995 2.465 ;
      RECT 86.825 0.255 87.08 0.825 ;
      RECT 86.075 1.485 86.405 2.465 ;
      RECT 86.175 0.255 86.405 2.465 ;
      RECT 86.075 1.75 86.535 1.92 ;
      RECT 86.075 0.255 86.405 0.885 ;
      RECT 84.695 1.485 85.025 2.465 ;
      RECT 84.795 0.255 85.025 2.465 ;
      RECT 84.795 1.075 86.005 1.315 ;
      RECT 84.695 0.255 85.025 0.885 ;
      RECT 83.315 1.485 83.645 2.465 ;
      RECT 83.415 0.255 83.645 2.465 ;
      RECT 83.315 1.555 83.775 1.725 ;
      RECT 83.315 0.255 83.645 0.885 ;
      RECT 81.935 1.485 82.265 2.465 ;
      RECT 82.035 0.255 82.265 2.465 ;
      RECT 82.035 1.075 83.245 1.315 ;
      RECT 81.935 0.255 82.265 0.885 ;
      RECT 80.615 1.875 81.13 2.285 ;
      RECT 80.79 0.895 81.13 2.285 ;
      RECT 79.9 0.895 81.13 1.065 ;
      RECT 80.61 0.29 80.855 1.065 ;
      RECT 78.01 2.295 80.04 2.465 ;
      RECT 79.87 1.44 80.04 2.465 ;
      RECT 78.01 0.995 78.18 2.465 ;
      RECT 79.87 1.44 80.62 1.63 ;
      RECT 77.985 0.995 78.18 1.325 ;
      RECT 78.69 1.615 79.7 1.785 ;
      RECT 79.51 0.255 79.7 1.785 ;
      RECT 78.69 0.815 78.86 1.785 ;
      RECT 78.35 1.955 79.475 2.125 ;
      RECT 78.35 0.255 78.52 2.125 ;
      RECT 77.505 0.995 77.76 1.325 ;
      RECT 77.59 0.655 77.76 1.325 ;
      RECT 77.59 0.655 78.52 0.825 ;
      RECT 78.345 0.255 78.52 0.825 ;
      RECT 78.345 0.255 78.875 0.62 ;
      RECT 77.165 1.495 77.5 2.465 ;
      RECT 77.165 0.255 77.335 2.465 ;
      RECT 77.165 0.255 77.42 0.825 ;
      RECT 76.48 1.875 76.995 2.285 ;
      RECT 76.655 0.895 76.995 2.285 ;
      RECT 75.765 0.895 76.995 1.065 ;
      RECT 76.475 0.29 76.72 1.065 ;
      RECT 73.875 2.295 75.905 2.465 ;
      RECT 75.735 1.44 75.905 2.465 ;
      RECT 73.875 0.995 74.045 2.465 ;
      RECT 75.735 1.44 76.485 1.63 ;
      RECT 73.85 0.995 74.045 1.325 ;
      RECT 74.555 1.615 75.565 1.785 ;
      RECT 75.375 0.255 75.565 1.785 ;
      RECT 74.555 0.815 74.725 1.785 ;
      RECT 74.215 1.955 75.34 2.125 ;
      RECT 74.215 0.255 74.385 2.125 ;
      RECT 73.37 0.995 73.625 1.325 ;
      RECT 73.455 0.655 73.625 1.325 ;
      RECT 73.455 0.655 74.385 0.825 ;
      RECT 74.21 0.255 74.385 0.825 ;
      RECT 74.21 0.255 74.74 0.62 ;
      RECT 73.03 1.495 73.365 2.465 ;
      RECT 73.03 0.255 73.2 2.465 ;
      RECT 73.03 0.255 73.285 0.825 ;
      RECT 71.935 0.475 72.665 0.715 ;
      RECT 72.477 0.27 72.665 0.715 ;
      RECT 72.305 0.282 72.68 0.709 ;
      RECT 72.22 0.297 72.7 0.694 ;
      RECT 72.22 0.312 72.705 0.684 ;
      RECT 72.175 0.332 72.72 0.676 ;
      RECT 72.152 0.367 72.735 0.63 ;
      RECT 72.066 0.39 72.74 0.59 ;
      RECT 72.066 0.408 72.75 0.56 ;
      RECT 71.935 0.477 72.755 0.523 ;
      RECT 71.98 0.42 72.75 0.56 ;
      RECT 72.066 0.372 72.735 0.63 ;
      RECT 72.152 0.341 72.72 0.676 ;
      RECT 72.175 0.322 72.705 0.684 ;
      RECT 72.22 0.295 72.68 0.709 ;
      RECT 72.305 0.277 72.665 0.715 ;
      RECT 72.391 0.271 72.665 0.715 ;
      RECT 72.477 0.266 72.61 0.715 ;
      RECT 72.563 0.261 72.61 0.715 ;
      RECT 72.255 1.159 72.425 1.545 ;
      RECT 72.25 1.159 72.425 1.54 ;
      RECT 72.225 1.159 72.425 1.505 ;
      RECT 72.225 1.187 72.435 1.495 ;
      RECT 72.205 1.187 72.435 1.455 ;
      RECT 72.2 1.187 72.435 1.428 ;
      RECT 72.2 1.205 72.44 1.42 ;
      RECT 72.145 1.205 72.44 1.355 ;
      RECT 72.145 1.222 72.45 1.338 ;
      RECT 72.135 1.222 72.45 1.278 ;
      RECT 72.135 1.239 72.455 1.275 ;
      RECT 72.13 1.075 72.3 1.253 ;
      RECT 72.13 1.109 72.386 1.253 ;
      RECT 72.125 1.875 72.13 1.888 ;
      RECT 72.12 1.77 72.125 1.893 ;
      RECT 72.095 1.63 72.12 1.908 ;
      RECT 72.06 1.581 72.095 1.94 ;
      RECT 72.055 1.549 72.06 1.96 ;
      RECT 72.05 1.54 72.055 1.96 ;
      RECT 71.97 1.505 72.05 1.96 ;
      RECT 71.907 1.475 71.97 1.96 ;
      RECT 71.821 1.463 71.907 1.96 ;
      RECT 71.735 1.449 71.821 1.96 ;
      RECT 71.655 1.436 71.735 1.946 ;
      RECT 71.62 1.428 71.655 1.926 ;
      RECT 71.61 1.425 71.62 1.917 ;
      RECT 71.58 1.42 71.61 1.904 ;
      RECT 71.53 1.395 71.58 1.88 ;
      RECT 71.516 1.369 71.53 1.862 ;
      RECT 71.43 1.329 71.516 1.838 ;
      RECT 71.385 1.277 71.43 1.807 ;
      RECT 71.375 1.252 71.385 1.794 ;
      RECT 71.37 1.033 71.375 1.055 ;
      RECT 71.365 1.235 71.375 1.79 ;
      RECT 71.365 1.031 71.37 1.145 ;
      RECT 71.355 1.027 71.365 1.786 ;
      RECT 71.311 1.025 71.355 1.774 ;
      RECT 71.225 1.025 71.311 1.745 ;
      RECT 71.195 1.025 71.225 1.718 ;
      RECT 71.18 1.025 71.195 1.706 ;
      RECT 71.14 1.037 71.18 1.691 ;
      RECT 71.12 1.056 71.14 1.67 ;
      RECT 71.11 1.066 71.12 1.654 ;
      RECT 71.1 1.072 71.11 1.643 ;
      RECT 71.08 1.082 71.1 1.626 ;
      RECT 71.075 1.091 71.08 1.613 ;
      RECT 71.07 1.095 71.075 1.563 ;
      RECT 71.06 1.101 71.07 1.48 ;
      RECT 71.055 1.105 71.06 1.394 ;
      RECT 71.05 1.125 71.055 1.331 ;
      RECT 71.045 1.148 71.05 1.278 ;
      RECT 71.04 1.166 71.045 1.223 ;
      RECT 71.65 0.985 71.82 1.245 ;
      RECT 71.82 0.95 71.865 1.231 ;
      RECT 71.781 0.952 71.87 1.214 ;
      RECT 71.67 0.969 71.956 1.185 ;
      RECT 71.67 0.984 71.96 1.157 ;
      RECT 71.67 0.965 71.87 1.214 ;
      RECT 71.695 0.953 71.82 1.245 ;
      RECT 71.781 0.951 71.865 1.231 ;
      RECT 70.835 0.34 71.005 0.83 ;
      RECT 70.835 0.34 71.04 0.81 ;
      RECT 70.97 0.26 71.08 0.77 ;
      RECT 70.951 0.264 71.1 0.74 ;
      RECT 70.865 0.272 71.12 0.723 ;
      RECT 70.865 0.278 71.125 0.713 ;
      RECT 70.865 0.287 71.145 0.701 ;
      RECT 70.84 0.312 71.175 0.679 ;
      RECT 70.84 0.332 71.18 0.659 ;
      RECT 70.835 0.345 71.19 0.639 ;
      RECT 70.835 0.412 71.195 0.62 ;
      RECT 70.835 0.545 71.2 0.607 ;
      RECT 70.83 0.35 71.19 0.44 ;
      RECT 70.84 0.307 71.145 0.701 ;
      RECT 70.951 0.262 71.08 0.77 ;
      RECT 70.825 2.015 71.125 2.27 ;
      RECT 70.91 1.981 71.125 2.27 ;
      RECT 70.91 1.984 71.13 2.13 ;
      RECT 70.845 2.005 71.13 2.13 ;
      RECT 70.88 1.995 71.125 2.27 ;
      RECT 70.875 2 71.13 2.13 ;
      RECT 70.91 1.979 71.111 2.27 ;
      RECT 70.996 1.97 71.111 2.27 ;
      RECT 70.996 1.964 71.025 2.27 ;
      RECT 70.485 1.605 70.495 2.095 ;
      RECT 70.145 1.54 70.155 1.84 ;
      RECT 70.66 1.712 70.665 1.931 ;
      RECT 70.65 1.692 70.66 1.948 ;
      RECT 70.64 1.672 70.65 1.978 ;
      RECT 70.635 1.662 70.64 1.993 ;
      RECT 70.63 1.658 70.635 1.998 ;
      RECT 70.615 1.65 70.63 2.005 ;
      RECT 70.575 1.63 70.615 2.03 ;
      RECT 70.55 1.612 70.575 2.063 ;
      RECT 70.545 1.61 70.55 2.076 ;
      RECT 70.525 1.607 70.545 2.08 ;
      RECT 70.495 1.605 70.525 2.09 ;
      RECT 70.425 1.607 70.485 2.091 ;
      RECT 70.405 1.607 70.425 2.085 ;
      RECT 70.38 1.605 70.405 2.082 ;
      RECT 70.345 1.6 70.38 2.078 ;
      RECT 70.325 1.594 70.345 2.065 ;
      RECT 70.315 1.591 70.325 2.053 ;
      RECT 70.295 1.588 70.315 2.038 ;
      RECT 70.275 1.584 70.295 2.02 ;
      RECT 70.27 1.581 70.275 2.01 ;
      RECT 70.265 1.58 70.27 2.008 ;
      RECT 70.255 1.577 70.265 2 ;
      RECT 70.245 1.571 70.255 1.983 ;
      RECT 70.235 1.565 70.245 1.965 ;
      RECT 70.225 1.559 70.235 1.953 ;
      RECT 70.215 1.553 70.225 1.933 ;
      RECT 70.21 1.549 70.215 1.918 ;
      RECT 70.205 1.547 70.21 1.91 ;
      RECT 70.2 1.545 70.205 1.903 ;
      RECT 70.195 1.543 70.2 1.893 ;
      RECT 70.19 1.541 70.195 1.887 ;
      RECT 70.18 1.54 70.19 1.877 ;
      RECT 70.17 1.54 70.18 1.868 ;
      RECT 70.155 1.54 70.17 1.853 ;
      RECT 70.115 1.54 70.145 1.837 ;
      RECT 70.095 1.542 70.115 1.832 ;
      RECT 70.09 1.547 70.095 1.83 ;
      RECT 70.06 1.555 70.09 1.828 ;
      RECT 70.03 1.57 70.06 1.827 ;
      RECT 69.985 1.592 70.03 1.832 ;
      RECT 69.98 1.607 69.985 1.836 ;
      RECT 69.965 1.612 69.98 1.838 ;
      RECT 69.96 1.616 69.965 1.84 ;
      RECT 69.9 1.639 69.96 1.849 ;
      RECT 69.88 1.665 69.9 1.862 ;
      RECT 69.87 1.672 69.88 1.866 ;
      RECT 69.855 1.679 69.87 1.869 ;
      RECT 69.835 1.689 69.855 1.872 ;
      RECT 69.83 1.697 69.835 1.875 ;
      RECT 69.785 1.702 69.83 1.882 ;
      RECT 69.775 1.705 69.785 1.889 ;
      RECT 69.765 1.705 69.775 1.893 ;
      RECT 69.73 1.707 69.765 1.905 ;
      RECT 69.71 1.71 69.73 1.918 ;
      RECT 69.67 1.713 69.71 1.929 ;
      RECT 69.655 1.715 69.67 1.942 ;
      RECT 69.645 1.715 69.655 1.947 ;
      RECT 69.62 1.716 69.645 1.955 ;
      RECT 69.61 1.718 69.62 1.96 ;
      RECT 69.605 1.719 69.61 1.963 ;
      RECT 69.58 1.717 69.605 1.966 ;
      RECT 69.565 1.715 69.58 1.967 ;
      RECT 69.545 1.712 69.565 1.969 ;
      RECT 69.525 1.707 69.545 1.969 ;
      RECT 69.465 1.702 69.525 1.966 ;
      RECT 69.43 1.677 69.465 1.962 ;
      RECT 69.42 1.654 69.43 1.96 ;
      RECT 69.39 1.631 69.42 1.96 ;
      RECT 69.38 1.61 69.39 1.96 ;
      RECT 69.355 1.592 69.38 1.958 ;
      RECT 69.34 1.57 69.355 1.955 ;
      RECT 69.325 1.552 69.34 1.953 ;
      RECT 69.305 1.542 69.325 1.951 ;
      RECT 69.29 1.537 69.305 1.95 ;
      RECT 69.275 1.535 69.29 1.949 ;
      RECT 69.245 1.536 69.275 1.947 ;
      RECT 69.225 1.539 69.245 1.945 ;
      RECT 69.168 1.543 69.225 1.945 ;
      RECT 69.082 1.552 69.168 1.945 ;
      RECT 68.996 1.563 69.082 1.945 ;
      RECT 68.91 1.574 68.996 1.945 ;
      RECT 68.89 1.581 68.91 1.953 ;
      RECT 68.88 1.584 68.89 1.96 ;
      RECT 68.815 1.589 68.88 1.978 ;
      RECT 68.785 1.596 68.815 2.003 ;
      RECT 68.775 1.599 68.785 2.01 ;
      RECT 68.73 1.603 68.775 2.015 ;
      RECT 68.7 1.608 68.73 2.02 ;
      RECT 68.699 1.61 68.7 2.02 ;
      RECT 68.613 1.616 68.699 2.02 ;
      RECT 68.527 1.627 68.613 2.02 ;
      RECT 68.441 1.639 68.527 2.02 ;
      RECT 68.355 1.65 68.441 2.02 ;
      RECT 68.34 1.657 68.355 2.015 ;
      RECT 68.335 1.659 68.34 2.009 ;
      RECT 68.315 1.67 68.335 2.004 ;
      RECT 68.305 1.688 68.315 1.998 ;
      RECT 68.3 1.7 68.305 1.798 ;
      RECT 70.595 0.453 70.615 0.54 ;
      RECT 70.59 0.388 70.595 0.572 ;
      RECT 70.58 0.355 70.59 0.577 ;
      RECT 70.575 0.335 70.58 0.583 ;
      RECT 70.545 0.335 70.575 0.6 ;
      RECT 70.496 0.335 70.545 0.636 ;
      RECT 70.41 0.335 70.496 0.694 ;
      RECT 70.381 0.345 70.41 0.743 ;
      RECT 70.295 0.387 70.381 0.796 ;
      RECT 70.275 0.425 70.295 0.843 ;
      RECT 70.25 0.442 70.275 0.863 ;
      RECT 70.24 0.456 70.25 0.883 ;
      RECT 70.235 0.462 70.24 0.893 ;
      RECT 70.23 0.466 70.235 0.9 ;
      RECT 70.18 0.486 70.23 0.905 ;
      RECT 70.115 0.53 70.18 0.905 ;
      RECT 70.09 0.58 70.115 0.905 ;
      RECT 70.08 0.61 70.09 0.905 ;
      RECT 70.075 0.637 70.08 0.905 ;
      RECT 70.07 0.655 70.075 0.905 ;
      RECT 70.06 0.697 70.07 0.905 ;
      RECT 70.41 1.255 70.58 1.43 ;
      RECT 70.35 1.083 70.41 1.418 ;
      RECT 70.34 1.076 70.35 1.401 ;
      RECT 70.295 1.255 70.58 1.381 ;
      RECT 70.276 1.255 70.58 1.359 ;
      RECT 70.19 1.255 70.58 1.324 ;
      RECT 70.17 1.075 70.34 1.28 ;
      RECT 70.17 1.222 70.575 1.28 ;
      RECT 70.17 1.17 70.55 1.28 ;
      RECT 70.17 1.125 70.515 1.28 ;
      RECT 70.17 1.107 70.48 1.28 ;
      RECT 70.17 1.097 70.475 1.28 ;
      RECT 69.89 2.055 70.08 2.28 ;
      RECT 69.88 2.056 70.085 2.275 ;
      RECT 69.88 2.058 70.095 2.255 ;
      RECT 69.88 2.062 70.1 2.24 ;
      RECT 69.88 2.049 70.05 2.275 ;
      RECT 69.88 2.052 70.075 2.275 ;
      RECT 69.89 2.048 70.05 2.28 ;
      RECT 69.976 2.046 70.05 2.28 ;
      RECT 69.6 1.297 69.77 1.535 ;
      RECT 69.6 1.297 69.856 1.449 ;
      RECT 69.6 1.297 69.86 1.359 ;
      RECT 69.65 1.07 69.87 1.338 ;
      RECT 69.645 1.087 69.875 1.311 ;
      RECT 69.61 1.245 69.875 1.311 ;
      RECT 69.63 1.095 69.77 1.535 ;
      RECT 69.62 1.177 69.88 1.294 ;
      RECT 69.615 1.225 69.88 1.294 ;
      RECT 69.62 1.135 69.875 1.311 ;
      RECT 69.645 1.072 69.87 1.338 ;
      RECT 69.21 1.047 69.38 1.245 ;
      RECT 69.21 1.047 69.425 1.22 ;
      RECT 69.28 0.99 69.45 1.178 ;
      RECT 69.255 1.005 69.45 1.178 ;
      RECT 68.87 1.051 68.9 1.245 ;
      RECT 68.865 1.023 68.87 1.245 ;
      RECT 68.835 0.997 68.865 1.247 ;
      RECT 68.81 0.955 68.835 1.25 ;
      RECT 68.8 0.927 68.81 1.252 ;
      RECT 68.765 0.907 68.8 1.254 ;
      RECT 68.7 0.892 68.765 1.26 ;
      RECT 68.65 0.89 68.7 1.266 ;
      RECT 68.627 0.892 68.65 1.271 ;
      RECT 68.541 0.903 68.627 1.277 ;
      RECT 68.455 0.921 68.541 1.287 ;
      RECT 68.44 0.932 68.455 1.293 ;
      RECT 68.37 0.955 68.44 1.299 ;
      RECT 68.315 0.987 68.37 1.307 ;
      RECT 68.275 1.01 68.315 1.313 ;
      RECT 68.261 1.023 68.275 1.316 ;
      RECT 68.175 1.045 68.261 1.322 ;
      RECT 68.16 1.07 68.175 1.328 ;
      RECT 68.12 1.085 68.16 1.332 ;
      RECT 68.07 1.1 68.12 1.337 ;
      RECT 68.045 1.107 68.07 1.341 ;
      RECT 67.985 1.102 68.045 1.345 ;
      RECT 67.97 1.093 67.985 1.349 ;
      RECT 67.9 1.083 67.97 1.345 ;
      RECT 67.875 1.075 67.895 1.335 ;
      RECT 67.816 1.075 67.875 1.313 ;
      RECT 67.73 1.075 67.816 1.27 ;
      RECT 67.895 1.075 67.9 1.34 ;
      RECT 68.59 0.306 68.76 0.64 ;
      RECT 68.56 0.306 68.76 0.635 ;
      RECT 68.5 0.273 68.56 0.623 ;
      RECT 68.5 0.329 68.77 0.618 ;
      RECT 68.475 0.329 68.77 0.612 ;
      RECT 68.47 0.27 68.5 0.609 ;
      RECT 68.455 0.276 68.59 0.607 ;
      RECT 68.45 0.284 68.675 0.595 ;
      RECT 68.45 0.336 68.785 0.548 ;
      RECT 68.435 0.292 68.675 0.543 ;
      RECT 68.435 0.362 68.795 0.484 ;
      RECT 68.405 0.312 68.76 0.445 ;
      RECT 68.405 0.402 68.805 0.441 ;
      RECT 68.455 0.281 68.675 0.607 ;
      RECT 67.795 0.611 67.85 0.875 ;
      RECT 67.795 0.611 67.915 0.874 ;
      RECT 67.795 0.611 67.94 0.873 ;
      RECT 67.795 0.611 68.005 0.872 ;
      RECT 67.94 0.577 68.02 0.871 ;
      RECT 67.755 0.621 68.165 0.87 ;
      RECT 67.795 0.618 68.165 0.87 ;
      RECT 67.755 0.626 68.17 0.863 ;
      RECT 67.74 0.628 68.17 0.862 ;
      RECT 67.74 0.635 68.175 0.858 ;
      RECT 67.72 0.634 68.17 0.854 ;
      RECT 67.72 0.642 68.18 0.853 ;
      RECT 67.715 0.639 68.175 0.849 ;
      RECT 67.715 0.652 68.19 0.848 ;
      RECT 67.7 0.642 68.18 0.847 ;
      RECT 67.665 0.655 68.19 0.84 ;
      RECT 67.85 0.61 68.16 0.87 ;
      RECT 67.85 0.595 68.11 0.87 ;
      RECT 67.915 0.582 68.045 0.87 ;
      RECT 67.46 1.671 67.475 2.064 ;
      RECT 67.425 1.676 67.475 2.063 ;
      RECT 67.46 1.675 67.52 2.062 ;
      RECT 67.405 1.686 67.52 2.061 ;
      RECT 67.42 1.682 67.52 2.061 ;
      RECT 67.385 1.692 67.595 2.058 ;
      RECT 67.385 1.711 67.64 2.056 ;
      RECT 67.385 1.718 67.645 2.053 ;
      RECT 67.37 1.695 67.595 2.05 ;
      RECT 67.35 1.7 67.595 2.043 ;
      RECT 67.345 1.704 67.595 2.039 ;
      RECT 67.345 1.721 67.655 2.038 ;
      RECT 67.325 1.715 67.64 2.034 ;
      RECT 67.325 1.724 67.66 2.028 ;
      RECT 67.32 1.73 67.66 1.8 ;
      RECT 67.385 1.69 67.52 2.058 ;
      RECT 67.26 1.053 67.46 1.365 ;
      RECT 67.335 1.031 67.46 1.365 ;
      RECT 67.275 1.05 67.465 1.35 ;
      RECT 67.245 1.061 67.465 1.348 ;
      RECT 67.26 1.056 67.47 1.314 ;
      RECT 67.245 1.16 67.475 1.281 ;
      RECT 67.275 1.032 67.46 1.365 ;
      RECT 67.335 1.01 67.435 1.365 ;
      RECT 67.36 1.007 67.435 1.365 ;
      RECT 67.36 1.002 67.38 1.365 ;
      RECT 66.765 1.07 66.94 1.245 ;
      RECT 66.76 1.07 66.94 1.243 ;
      RECT 66.735 1.07 66.94 1.238 ;
      RECT 66.68 1.05 66.85 1.228 ;
      RECT 66.68 1.057 66.915 1.228 ;
      RECT 66.765 1.737 66.78 1.92 ;
      RECT 66.755 1.715 66.765 1.92 ;
      RECT 66.74 1.695 66.755 1.92 ;
      RECT 66.73 1.67 66.74 1.92 ;
      RECT 66.7 1.635 66.73 1.92 ;
      RECT 66.665 1.575 66.7 1.92 ;
      RECT 66.66 1.537 66.665 1.92 ;
      RECT 66.61 1.488 66.66 1.92 ;
      RECT 66.6 1.438 66.61 1.908 ;
      RECT 66.585 1.417 66.6 1.868 ;
      RECT 66.565 1.385 66.585 1.818 ;
      RECT 66.54 1.341 66.565 1.758 ;
      RECT 66.535 1.313 66.54 1.713 ;
      RECT 66.53 1.304 66.535 1.699 ;
      RECT 66.525 1.297 66.53 1.686 ;
      RECT 66.52 1.292 66.525 1.675 ;
      RECT 66.515 1.277 66.52 1.665 ;
      RECT 66.51 1.255 66.515 1.652 ;
      RECT 66.5 1.215 66.51 1.627 ;
      RECT 66.475 1.145 66.5 1.583 ;
      RECT 66.47 1.085 66.475 1.548 ;
      RECT 66.455 1.065 66.47 1.515 ;
      RECT 66.45 1.065 66.455 1.49 ;
      RECT 66.42 1.065 66.45 1.445 ;
      RECT 66.375 1.065 66.42 1.385 ;
      RECT 66.3 1.065 66.375 1.333 ;
      RECT 66.295 1.065 66.3 1.298 ;
      RECT 66.29 1.065 66.295 1.288 ;
      RECT 66.285 1.065 66.29 1.268 ;
      RECT 66.55 0.285 66.72 0.755 ;
      RECT 66.495 0.278 66.69 0.739 ;
      RECT 66.495 0.292 66.725 0.738 ;
      RECT 66.48 0.293 66.725 0.719 ;
      RECT 66.475 0.311 66.725 0.705 ;
      RECT 66.48 0.294 66.73 0.703 ;
      RECT 66.465 0.325 66.73 0.688 ;
      RECT 66.48 0.3 66.735 0.673 ;
      RECT 66.46 0.34 66.735 0.67 ;
      RECT 66.475 0.312 66.74 0.655 ;
      RECT 66.475 0.324 66.745 0.635 ;
      RECT 66.46 0.34 66.75 0.618 ;
      RECT 66.46 0.35 66.755 0.473 ;
      RECT 66.455 0.35 66.755 0.43 ;
      RECT 66.455 0.365 66.76 0.408 ;
      RECT 66.55 0.275 66.69 0.755 ;
      RECT 66.55 0.273 66.66 0.755 ;
      RECT 66.636 0.27 66.66 0.755 ;
      RECT 66.295 1.937 66.3 1.983 ;
      RECT 66.285 1.785 66.295 2.007 ;
      RECT 66.28 1.63 66.285 2.032 ;
      RECT 66.265 1.592 66.28 2.043 ;
      RECT 66.26 1.575 66.265 2.05 ;
      RECT 66.25 1.563 66.26 2.057 ;
      RECT 66.245 1.554 66.25 2.059 ;
      RECT 66.24 1.552 66.245 2.063 ;
      RECT 66.195 1.543 66.24 2.078 ;
      RECT 66.19 1.535 66.195 2.092 ;
      RECT 66.185 1.532 66.19 2.096 ;
      RECT 66.17 1.527 66.185 2.104 ;
      RECT 66.115 1.517 66.17 2.115 ;
      RECT 66.08 1.505 66.115 2.116 ;
      RECT 66.071 1.5 66.08 2.11 ;
      RECT 65.985 1.5 66.071 2.1 ;
      RECT 65.955 1.5 65.985 2.078 ;
      RECT 65.945 1.5 65.95 2.058 ;
      RECT 65.94 1.5 65.945 2.02 ;
      RECT 65.935 1.5 65.94 1.978 ;
      RECT 65.93 1.5 65.935 1.938 ;
      RECT 65.925 1.5 65.93 1.868 ;
      RECT 65.915 1.5 65.925 1.79 ;
      RECT 65.91 1.5 65.915 1.69 ;
      RECT 65.95 1.5 65.955 2.06 ;
      RECT 65.445 1.582 65.535 2.06 ;
      RECT 65.43 1.585 65.55 2.058 ;
      RECT 65.445 1.584 65.55 2.058 ;
      RECT 65.41 1.591 65.575 2.048 ;
      RECT 65.43 1.585 65.575 2.048 ;
      RECT 65.395 1.597 65.575 2.036 ;
      RECT 65.43 1.588 65.625 2.029 ;
      RECT 65.381 1.605 65.625 2.027 ;
      RECT 65.41 1.595 65.635 2.015 ;
      RECT 65.381 1.616 65.665 2.006 ;
      RECT 65.295 1.64 65.665 2 ;
      RECT 65.295 1.653 65.705 1.983 ;
      RECT 65.29 1.675 65.705 1.976 ;
      RECT 65.26 1.69 65.705 1.966 ;
      RECT 65.255 1.701 65.705 1.956 ;
      RECT 65.225 1.714 65.705 1.947 ;
      RECT 65.21 1.732 65.705 1.936 ;
      RECT 65.185 1.745 65.705 1.926 ;
      RECT 65.445 1.581 65.455 2.06 ;
      RECT 65.491 1.005 65.53 1.25 ;
      RECT 65.405 1.005 65.54 1.248 ;
      RECT 65.29 1.03 65.54 1.245 ;
      RECT 65.29 1.03 65.545 1.243 ;
      RECT 65.29 1.03 65.56 1.238 ;
      RECT 65.396 1.005 65.575 1.218 ;
      RECT 65.31 1.013 65.575 1.218 ;
      RECT 64.98 0.365 65.15 0.8 ;
      RECT 64.97 0.399 65.15 0.783 ;
      RECT 65.05 0.335 65.22 0.77 ;
      RECT 64.955 0.41 65.22 0.748 ;
      RECT 65.05 0.345 65.225 0.738 ;
      RECT 64.98 0.397 65.255 0.723 ;
      RECT 64.94 0.423 65.255 0.708 ;
      RECT 64.94 0.465 65.265 0.688 ;
      RECT 64.935 0.49 65.27 0.67 ;
      RECT 64.935 0.5 65.275 0.655 ;
      RECT 64.93 0.437 65.255 0.653 ;
      RECT 64.93 0.51 65.28 0.638 ;
      RECT 64.925 0.447 65.255 0.635 ;
      RECT 64.92 0.531 65.285 0.618 ;
      RECT 64.92 0.563 65.29 0.598 ;
      RECT 64.915 0.477 65.265 0.59 ;
      RECT 64.92 0.462 65.255 0.618 ;
      RECT 64.935 0.432 65.255 0.67 ;
      RECT 64.78 1.019 65.005 1.275 ;
      RECT 64.78 1.052 65.025 1.265 ;
      RECT 64.745 1.052 65.025 1.263 ;
      RECT 64.745 1.065 65.03 1.253 ;
      RECT 64.745 1.085 65.04 1.245 ;
      RECT 64.745 1.182 65.045 1.238 ;
      RECT 64.725 0.93 64.855 1.228 ;
      RECT 64.68 1.085 65.04 1.17 ;
      RECT 64.67 0.93 64.855 1.115 ;
      RECT 64.67 0.962 64.941 1.115 ;
      RECT 64.635 1.492 64.655 1.67 ;
      RECT 64.6 1.445 64.635 1.67 ;
      RECT 64.585 1.385 64.6 1.67 ;
      RECT 64.56 1.332 64.585 1.67 ;
      RECT 64.545 1.285 64.56 1.67 ;
      RECT 64.525 1.262 64.545 1.67 ;
      RECT 64.5 1.227 64.525 1.67 ;
      RECT 64.49 1.073 64.5 1.67 ;
      RECT 64.46 1.068 64.49 1.661 ;
      RECT 64.455 1.065 64.46 1.651 ;
      RECT 64.44 1.065 64.455 1.625 ;
      RECT 64.435 1.065 64.44 1.588 ;
      RECT 64.41 1.065 64.435 1.54 ;
      RECT 64.39 1.065 64.41 1.465 ;
      RECT 64.38 1.065 64.39 1.425 ;
      RECT 64.375 1.065 64.38 1.4 ;
      RECT 64.37 1.065 64.375 1.383 ;
      RECT 64.365 1.065 64.37 1.365 ;
      RECT 64.36 1.066 64.365 1.355 ;
      RECT 64.35 1.068 64.36 1.323 ;
      RECT 64.34 1.07 64.35 1.29 ;
      RECT 64.33 1.073 64.34 1.263 ;
      RECT 64.655 1.5 64.88 1.67 ;
      RECT 63.985 0.312 64.155 0.765 ;
      RECT 63.985 0.312 64.245 0.731 ;
      RECT 63.985 0.312 64.275 0.715 ;
      RECT 63.985 0.312 64.305 0.688 ;
      RECT 64.241 0.29 64.32 0.67 ;
      RECT 64.02 0.297 64.325 0.655 ;
      RECT 64.02 0.305 64.335 0.618 ;
      RECT 63.98 0.332 64.335 0.59 ;
      RECT 63.965 0.345 64.335 0.555 ;
      RECT 63.985 0.32 64.355 0.545 ;
      RECT 63.96 0.385 64.355 0.515 ;
      RECT 63.96 0.415 64.36 0.498 ;
      RECT 63.955 0.445 64.36 0.485 ;
      RECT 64.02 0.294 64.32 0.67 ;
      RECT 64.155 0.291 64.241 0.749 ;
      RECT 64.106 0.292 64.32 0.67 ;
      RECT 64.25 1.952 64.295 2.145 ;
      RECT 64.24 1.922 64.25 2.145 ;
      RECT 64.235 1.907 64.24 2.145 ;
      RECT 64.195 1.817 64.235 2.145 ;
      RECT 64.19 1.73 64.195 2.145 ;
      RECT 64.18 1.7 64.19 2.145 ;
      RECT 64.175 1.66 64.18 2.145 ;
      RECT 64.165 1.622 64.175 2.145 ;
      RECT 64.16 1.587 64.165 2.145 ;
      RECT 64.14 1.54 64.16 2.145 ;
      RECT 64.125 1.465 64.14 2.145 ;
      RECT 64.12 1.42 64.125 2.14 ;
      RECT 64.115 1.4 64.12 2.113 ;
      RECT 64.11 1.38 64.115 2.098 ;
      RECT 64.105 1.355 64.11 2.078 ;
      RECT 64.1 1.333 64.105 2.063 ;
      RECT 64.095 1.311 64.1 2.045 ;
      RECT 64.09 1.29 64.095 2.035 ;
      RECT 64.08 1.262 64.09 2.005 ;
      RECT 64.07 1.225 64.08 1.973 ;
      RECT 64.06 1.185 64.07 1.94 ;
      RECT 64.05 1.163 64.06 1.91 ;
      RECT 64.02 1.115 64.05 1.842 ;
      RECT 64.005 1.075 64.02 1.769 ;
      RECT 63.995 1.075 64.005 1.735 ;
      RECT 63.99 1.075 63.995 1.71 ;
      RECT 63.985 1.075 63.99 1.695 ;
      RECT 63.98 1.075 63.985 1.673 ;
      RECT 63.975 1.075 63.98 1.66 ;
      RECT 63.96 1.075 63.975 1.625 ;
      RECT 63.94 1.075 63.96 1.565 ;
      RECT 63.93 1.075 63.94 1.515 ;
      RECT 63.91 1.075 63.93 1.463 ;
      RECT 63.89 1.075 63.91 1.42 ;
      RECT 63.88 1.075 63.89 1.408 ;
      RECT 63.85 1.075 63.88 1.395 ;
      RECT 63.82 1.096 63.85 1.375 ;
      RECT 63.81 1.124 63.82 1.355 ;
      RECT 63.795 1.141 63.81 1.323 ;
      RECT 63.79 1.155 63.795 1.29 ;
      RECT 63.785 1.163 63.79 1.263 ;
      RECT 63.78 1.171 63.785 1.225 ;
      RECT 63.785 1.695 63.79 2.03 ;
      RECT 63.75 1.682 63.785 2.029 ;
      RECT 63.68 1.622 63.75 2.028 ;
      RECT 63.6 1.565 63.68 2.027 ;
      RECT 63.465 1.525 63.6 2.026 ;
      RECT 63.465 1.712 63.8 2.015 ;
      RECT 63.425 1.712 63.8 2.005 ;
      RECT 63.425 1.73 63.805 2 ;
      RECT 63.425 1.82 63.81 1.99 ;
      RECT 63.42 1.515 63.585 1.97 ;
      RECT 63.415 1.515 63.585 1.713 ;
      RECT 63.415 1.672 63.78 1.713 ;
      RECT 63.415 1.66 63.775 1.713 ;
      RECT 62.68 1.875 63.195 2.285 ;
      RECT 62.855 0.895 63.195 2.285 ;
      RECT 61.965 0.895 63.195 1.065 ;
      RECT 62.675 0.29 62.92 1.065 ;
      RECT 60.075 2.295 62.105 2.465 ;
      RECT 61.935 1.44 62.105 2.465 ;
      RECT 60.075 0.995 60.245 2.465 ;
      RECT 61.935 1.44 62.685 1.63 ;
      RECT 60.05 0.995 60.245 1.325 ;
      RECT 60.755 1.615 61.765 1.785 ;
      RECT 61.575 0.255 61.765 1.785 ;
      RECT 60.755 0.815 60.925 1.785 ;
      RECT 60.415 1.955 61.54 2.125 ;
      RECT 60.415 0.255 60.585 2.125 ;
      RECT 59.57 0.995 59.825 1.325 ;
      RECT 59.655 0.655 59.825 1.325 ;
      RECT 59.655 0.655 60.585 0.825 ;
      RECT 60.41 0.255 60.585 0.825 ;
      RECT 60.41 0.255 60.94 0.62 ;
      RECT 59.23 1.495 59.565 2.465 ;
      RECT 59.23 0.255 59.4 2.465 ;
      RECT 59.23 0.255 59.485 0.825 ;
      RECT 58.48 1.485 58.81 2.465 ;
      RECT 58.58 0.255 58.81 2.465 ;
      RECT 58.48 1.735 58.94 1.9 ;
      RECT 58.48 0.255 58.81 0.885 ;
      RECT 57.1 1.485 57.43 2.465 ;
      RECT 57.2 0.255 57.43 2.465 ;
      RECT 57.2 1.075 58.41 1.315 ;
      RECT 57.1 0.255 57.43 0.885 ;
      RECT 55.72 1.485 56.05 2.465 ;
      RECT 55.82 0.255 56.05 2.465 ;
      RECT 55.72 1.555 56.185 1.725 ;
      RECT 55.72 0.255 56.05 0.885 ;
      RECT 54.34 1.485 54.67 2.465 ;
      RECT 54.44 0.255 54.67 2.465 ;
      RECT 54.44 1.075 55.65 1.315 ;
      RECT 54.34 0.255 54.67 0.885 ;
      RECT 53.02 1.875 53.535 2.285 ;
      RECT 53.195 0.895 53.535 2.285 ;
      RECT 52.305 0.895 53.535 1.065 ;
      RECT 53.015 0.29 53.26 1.065 ;
      RECT 50.415 2.295 52.445 2.465 ;
      RECT 52.275 1.44 52.445 2.465 ;
      RECT 50.415 0.995 50.585 2.465 ;
      RECT 52.275 1.44 53.025 1.63 ;
      RECT 50.39 0.995 50.585 1.325 ;
      RECT 51.095 1.615 52.105 1.785 ;
      RECT 51.915 0.255 52.105 1.785 ;
      RECT 51.095 0.815 51.265 1.785 ;
      RECT 50.755 1.955 51.88 2.125 ;
      RECT 50.755 0.255 50.925 2.125 ;
      RECT 49.91 0.995 50.165 1.325 ;
      RECT 49.995 0.655 50.165 1.325 ;
      RECT 49.995 0.655 50.925 0.825 ;
      RECT 50.75 0.255 50.925 0.825 ;
      RECT 50.75 0.255 51.28 0.62 ;
      RECT 49.57 1.495 49.905 2.465 ;
      RECT 49.57 0.255 49.74 2.465 ;
      RECT 49.57 0.255 49.825 0.825 ;
      RECT 48.885 1.875 49.4 2.285 ;
      RECT 49.06 0.895 49.4 2.285 ;
      RECT 48.17 0.895 49.4 1.065 ;
      RECT 48.88 0.29 49.125 1.065 ;
      RECT 46.28 2.295 48.31 2.465 ;
      RECT 48.14 1.44 48.31 2.465 ;
      RECT 46.28 0.995 46.45 2.465 ;
      RECT 48.14 1.44 48.89 1.63 ;
      RECT 46.255 0.995 46.45 1.325 ;
      RECT 46.96 1.615 47.97 1.785 ;
      RECT 47.78 0.255 47.97 1.785 ;
      RECT 46.96 0.815 47.13 1.785 ;
      RECT 46.62 1.955 47.745 2.125 ;
      RECT 46.62 0.255 46.79 2.125 ;
      RECT 45.775 0.995 46.03 1.325 ;
      RECT 45.86 0.655 46.03 1.325 ;
      RECT 45.86 0.655 46.79 0.825 ;
      RECT 46.615 0.255 46.79 0.825 ;
      RECT 46.615 0.255 47.145 0.62 ;
      RECT 45.435 1.495 45.77 2.465 ;
      RECT 45.435 0.255 45.605 2.465 ;
      RECT 45.435 0.255 45.69 0.825 ;
      RECT 44.34 0.475 45.07 0.715 ;
      RECT 44.882 0.27 45.07 0.715 ;
      RECT 44.71 0.282 45.085 0.709 ;
      RECT 44.625 0.297 45.105 0.694 ;
      RECT 44.625 0.312 45.11 0.684 ;
      RECT 44.58 0.332 45.125 0.676 ;
      RECT 44.557 0.367 45.14 0.63 ;
      RECT 44.471 0.39 45.145 0.59 ;
      RECT 44.471 0.408 45.155 0.56 ;
      RECT 44.34 0.477 45.16 0.523 ;
      RECT 44.385 0.42 45.155 0.56 ;
      RECT 44.471 0.372 45.14 0.63 ;
      RECT 44.557 0.341 45.125 0.676 ;
      RECT 44.58 0.322 45.11 0.684 ;
      RECT 44.625 0.295 45.085 0.709 ;
      RECT 44.71 0.277 45.07 0.715 ;
      RECT 44.796 0.271 45.07 0.715 ;
      RECT 44.882 0.266 45.015 0.715 ;
      RECT 44.968 0.261 45.015 0.715 ;
      RECT 44.66 1.159 44.83 1.545 ;
      RECT 44.655 1.159 44.83 1.54 ;
      RECT 44.63 1.159 44.83 1.505 ;
      RECT 44.63 1.187 44.84 1.495 ;
      RECT 44.61 1.187 44.84 1.455 ;
      RECT 44.605 1.187 44.84 1.428 ;
      RECT 44.605 1.205 44.845 1.42 ;
      RECT 44.55 1.205 44.845 1.355 ;
      RECT 44.55 1.222 44.855 1.338 ;
      RECT 44.54 1.222 44.855 1.278 ;
      RECT 44.54 1.239 44.86 1.275 ;
      RECT 44.535 1.075 44.705 1.253 ;
      RECT 44.535 1.109 44.791 1.253 ;
      RECT 44.53 1.875 44.535 1.888 ;
      RECT 44.525 1.77 44.53 1.893 ;
      RECT 44.5 1.63 44.525 1.908 ;
      RECT 44.465 1.581 44.5 1.94 ;
      RECT 44.46 1.549 44.465 1.96 ;
      RECT 44.455 1.54 44.46 1.96 ;
      RECT 44.375 1.505 44.455 1.96 ;
      RECT 44.312 1.475 44.375 1.96 ;
      RECT 44.226 1.463 44.312 1.96 ;
      RECT 44.14 1.449 44.226 1.96 ;
      RECT 44.06 1.436 44.14 1.946 ;
      RECT 44.025 1.428 44.06 1.926 ;
      RECT 44.015 1.425 44.025 1.917 ;
      RECT 43.985 1.42 44.015 1.904 ;
      RECT 43.935 1.395 43.985 1.88 ;
      RECT 43.921 1.369 43.935 1.862 ;
      RECT 43.835 1.329 43.921 1.838 ;
      RECT 43.79 1.277 43.835 1.807 ;
      RECT 43.78 1.252 43.79 1.794 ;
      RECT 43.775 1.033 43.78 1.055 ;
      RECT 43.77 1.235 43.78 1.79 ;
      RECT 43.77 1.031 43.775 1.145 ;
      RECT 43.76 1.027 43.77 1.786 ;
      RECT 43.716 1.025 43.76 1.774 ;
      RECT 43.63 1.025 43.716 1.745 ;
      RECT 43.6 1.025 43.63 1.718 ;
      RECT 43.585 1.025 43.6 1.706 ;
      RECT 43.545 1.037 43.585 1.691 ;
      RECT 43.525 1.056 43.545 1.67 ;
      RECT 43.515 1.066 43.525 1.654 ;
      RECT 43.505 1.072 43.515 1.643 ;
      RECT 43.485 1.082 43.505 1.626 ;
      RECT 43.48 1.091 43.485 1.613 ;
      RECT 43.475 1.095 43.48 1.563 ;
      RECT 43.465 1.101 43.475 1.48 ;
      RECT 43.46 1.105 43.465 1.394 ;
      RECT 43.455 1.125 43.46 1.331 ;
      RECT 43.45 1.148 43.455 1.278 ;
      RECT 43.445 1.166 43.45 1.223 ;
      RECT 44.055 0.985 44.225 1.245 ;
      RECT 44.225 0.95 44.27 1.231 ;
      RECT 44.186 0.952 44.275 1.214 ;
      RECT 44.075 0.969 44.361 1.185 ;
      RECT 44.075 0.984 44.365 1.157 ;
      RECT 44.075 0.965 44.275 1.214 ;
      RECT 44.1 0.953 44.225 1.245 ;
      RECT 44.186 0.951 44.27 1.231 ;
      RECT 43.24 0.34 43.41 0.83 ;
      RECT 43.24 0.34 43.445 0.81 ;
      RECT 43.375 0.26 43.485 0.77 ;
      RECT 43.356 0.264 43.505 0.74 ;
      RECT 43.27 0.272 43.525 0.723 ;
      RECT 43.27 0.278 43.53 0.713 ;
      RECT 43.27 0.287 43.55 0.701 ;
      RECT 43.245 0.312 43.58 0.679 ;
      RECT 43.245 0.332 43.585 0.659 ;
      RECT 43.24 0.345 43.595 0.639 ;
      RECT 43.24 0.412 43.6 0.62 ;
      RECT 43.24 0.545 43.605 0.607 ;
      RECT 43.235 0.35 43.595 0.44 ;
      RECT 43.245 0.307 43.55 0.701 ;
      RECT 43.356 0.262 43.485 0.77 ;
      RECT 43.23 2.015 43.53 2.27 ;
      RECT 43.315 1.981 43.53 2.27 ;
      RECT 43.315 1.984 43.535 2.13 ;
      RECT 43.25 2.005 43.535 2.13 ;
      RECT 43.285 1.995 43.53 2.27 ;
      RECT 43.28 2 43.535 2.13 ;
      RECT 43.315 1.979 43.516 2.27 ;
      RECT 43.401 1.97 43.516 2.27 ;
      RECT 43.401 1.964 43.43 2.27 ;
      RECT 42.89 1.605 42.9 2.095 ;
      RECT 42.55 1.54 42.56 1.84 ;
      RECT 43.065 1.712 43.07 1.931 ;
      RECT 43.055 1.692 43.065 1.948 ;
      RECT 43.045 1.672 43.055 1.978 ;
      RECT 43.04 1.662 43.045 1.993 ;
      RECT 43.035 1.658 43.04 1.998 ;
      RECT 43.02 1.65 43.035 2.005 ;
      RECT 42.98 1.63 43.02 2.03 ;
      RECT 42.955 1.612 42.98 2.063 ;
      RECT 42.95 1.61 42.955 2.076 ;
      RECT 42.93 1.607 42.95 2.08 ;
      RECT 42.9 1.605 42.93 2.09 ;
      RECT 42.83 1.607 42.89 2.091 ;
      RECT 42.81 1.607 42.83 2.085 ;
      RECT 42.785 1.605 42.81 2.082 ;
      RECT 42.75 1.6 42.785 2.078 ;
      RECT 42.73 1.594 42.75 2.065 ;
      RECT 42.72 1.591 42.73 2.053 ;
      RECT 42.7 1.588 42.72 2.038 ;
      RECT 42.68 1.584 42.7 2.02 ;
      RECT 42.675 1.581 42.68 2.01 ;
      RECT 42.67 1.58 42.675 2.008 ;
      RECT 42.66 1.577 42.67 2 ;
      RECT 42.65 1.571 42.66 1.983 ;
      RECT 42.64 1.565 42.65 1.965 ;
      RECT 42.63 1.559 42.64 1.953 ;
      RECT 42.62 1.553 42.63 1.933 ;
      RECT 42.615 1.549 42.62 1.918 ;
      RECT 42.61 1.547 42.615 1.91 ;
      RECT 42.605 1.545 42.61 1.903 ;
      RECT 42.6 1.543 42.605 1.893 ;
      RECT 42.595 1.541 42.6 1.887 ;
      RECT 42.585 1.54 42.595 1.877 ;
      RECT 42.575 1.54 42.585 1.868 ;
      RECT 42.56 1.54 42.575 1.853 ;
      RECT 42.52 1.54 42.55 1.837 ;
      RECT 42.5 1.542 42.52 1.832 ;
      RECT 42.495 1.547 42.5 1.83 ;
      RECT 42.465 1.555 42.495 1.828 ;
      RECT 42.435 1.57 42.465 1.827 ;
      RECT 42.39 1.592 42.435 1.832 ;
      RECT 42.385 1.607 42.39 1.836 ;
      RECT 42.37 1.612 42.385 1.838 ;
      RECT 42.365 1.616 42.37 1.84 ;
      RECT 42.305 1.639 42.365 1.849 ;
      RECT 42.285 1.665 42.305 1.862 ;
      RECT 42.275 1.672 42.285 1.866 ;
      RECT 42.26 1.679 42.275 1.869 ;
      RECT 42.24 1.689 42.26 1.872 ;
      RECT 42.235 1.697 42.24 1.875 ;
      RECT 42.19 1.702 42.235 1.882 ;
      RECT 42.18 1.705 42.19 1.889 ;
      RECT 42.17 1.705 42.18 1.893 ;
      RECT 42.135 1.707 42.17 1.905 ;
      RECT 42.115 1.71 42.135 1.918 ;
      RECT 42.075 1.713 42.115 1.929 ;
      RECT 42.06 1.715 42.075 1.942 ;
      RECT 42.05 1.715 42.06 1.947 ;
      RECT 42.025 1.716 42.05 1.955 ;
      RECT 42.015 1.718 42.025 1.96 ;
      RECT 42.01 1.719 42.015 1.963 ;
      RECT 41.985 1.717 42.01 1.966 ;
      RECT 41.97 1.715 41.985 1.967 ;
      RECT 41.95 1.712 41.97 1.969 ;
      RECT 41.93 1.707 41.95 1.969 ;
      RECT 41.87 1.702 41.93 1.966 ;
      RECT 41.835 1.677 41.87 1.962 ;
      RECT 41.825 1.654 41.835 1.96 ;
      RECT 41.795 1.631 41.825 1.96 ;
      RECT 41.785 1.61 41.795 1.96 ;
      RECT 41.76 1.592 41.785 1.958 ;
      RECT 41.745 1.57 41.76 1.955 ;
      RECT 41.73 1.552 41.745 1.953 ;
      RECT 41.71 1.542 41.73 1.951 ;
      RECT 41.695 1.537 41.71 1.95 ;
      RECT 41.68 1.535 41.695 1.949 ;
      RECT 41.65 1.536 41.68 1.947 ;
      RECT 41.63 1.539 41.65 1.945 ;
      RECT 41.573 1.543 41.63 1.945 ;
      RECT 41.487 1.552 41.573 1.945 ;
      RECT 41.401 1.563 41.487 1.945 ;
      RECT 41.315 1.574 41.401 1.945 ;
      RECT 41.295 1.581 41.315 1.953 ;
      RECT 41.285 1.584 41.295 1.96 ;
      RECT 41.22 1.589 41.285 1.978 ;
      RECT 41.19 1.596 41.22 2.003 ;
      RECT 41.18 1.599 41.19 2.01 ;
      RECT 41.135 1.603 41.18 2.015 ;
      RECT 41.105 1.608 41.135 2.02 ;
      RECT 41.104 1.61 41.105 2.02 ;
      RECT 41.018 1.616 41.104 2.02 ;
      RECT 40.932 1.627 41.018 2.02 ;
      RECT 40.846 1.639 40.932 2.02 ;
      RECT 40.76 1.65 40.846 2.02 ;
      RECT 40.745 1.657 40.76 2.015 ;
      RECT 40.74 1.659 40.745 2.009 ;
      RECT 40.72 1.67 40.74 2.004 ;
      RECT 40.71 1.688 40.72 1.998 ;
      RECT 40.705 1.7 40.71 1.798 ;
      RECT 43 0.453 43.02 0.54 ;
      RECT 42.995 0.388 43 0.572 ;
      RECT 42.985 0.355 42.995 0.577 ;
      RECT 42.98 0.335 42.985 0.583 ;
      RECT 42.95 0.335 42.98 0.6 ;
      RECT 42.901 0.335 42.95 0.636 ;
      RECT 42.815 0.335 42.901 0.694 ;
      RECT 42.786 0.345 42.815 0.743 ;
      RECT 42.7 0.387 42.786 0.796 ;
      RECT 42.68 0.425 42.7 0.843 ;
      RECT 42.655 0.442 42.68 0.863 ;
      RECT 42.645 0.456 42.655 0.883 ;
      RECT 42.64 0.462 42.645 0.893 ;
      RECT 42.635 0.466 42.64 0.9 ;
      RECT 42.585 0.486 42.635 0.905 ;
      RECT 42.52 0.53 42.585 0.905 ;
      RECT 42.495 0.58 42.52 0.905 ;
      RECT 42.485 0.61 42.495 0.905 ;
      RECT 42.48 0.637 42.485 0.905 ;
      RECT 42.475 0.655 42.48 0.905 ;
      RECT 42.465 0.697 42.475 0.905 ;
      RECT 42.815 1.255 42.985 1.43 ;
      RECT 42.755 1.083 42.815 1.418 ;
      RECT 42.745 1.076 42.755 1.401 ;
      RECT 42.7 1.255 42.985 1.381 ;
      RECT 42.681 1.255 42.985 1.359 ;
      RECT 42.595 1.255 42.985 1.324 ;
      RECT 42.575 1.075 42.745 1.28 ;
      RECT 42.575 1.222 42.98 1.28 ;
      RECT 42.575 1.17 42.955 1.28 ;
      RECT 42.575 1.125 42.92 1.28 ;
      RECT 42.575 1.107 42.885 1.28 ;
      RECT 42.575 1.097 42.88 1.28 ;
      RECT 42.295 2.055 42.485 2.28 ;
      RECT 42.285 2.056 42.49 2.275 ;
      RECT 42.285 2.058 42.5 2.255 ;
      RECT 42.285 2.062 42.505 2.24 ;
      RECT 42.285 2.049 42.455 2.275 ;
      RECT 42.285 2.052 42.48 2.275 ;
      RECT 42.295 2.048 42.455 2.28 ;
      RECT 42.381 2.046 42.455 2.28 ;
      RECT 42.005 1.297 42.175 1.535 ;
      RECT 42.005 1.297 42.261 1.449 ;
      RECT 42.005 1.297 42.265 1.359 ;
      RECT 42.055 1.07 42.275 1.338 ;
      RECT 42.05 1.087 42.28 1.311 ;
      RECT 42.015 1.245 42.28 1.311 ;
      RECT 42.035 1.095 42.175 1.535 ;
      RECT 42.025 1.177 42.285 1.294 ;
      RECT 42.02 1.225 42.285 1.294 ;
      RECT 42.025 1.135 42.28 1.311 ;
      RECT 42.05 1.072 42.275 1.338 ;
      RECT 41.615 1.047 41.785 1.245 ;
      RECT 41.615 1.047 41.83 1.22 ;
      RECT 41.685 0.99 41.855 1.178 ;
      RECT 41.66 1.005 41.855 1.178 ;
      RECT 41.275 1.051 41.305 1.245 ;
      RECT 41.27 1.023 41.275 1.245 ;
      RECT 41.24 0.997 41.27 1.247 ;
      RECT 41.215 0.955 41.24 1.25 ;
      RECT 41.205 0.927 41.215 1.252 ;
      RECT 41.17 0.907 41.205 1.254 ;
      RECT 41.105 0.892 41.17 1.26 ;
      RECT 41.055 0.89 41.105 1.266 ;
      RECT 41.032 0.892 41.055 1.271 ;
      RECT 40.946 0.903 41.032 1.277 ;
      RECT 40.86 0.921 40.946 1.287 ;
      RECT 40.845 0.932 40.86 1.293 ;
      RECT 40.775 0.955 40.845 1.299 ;
      RECT 40.72 0.987 40.775 1.307 ;
      RECT 40.68 1.01 40.72 1.313 ;
      RECT 40.666 1.023 40.68 1.316 ;
      RECT 40.58 1.045 40.666 1.322 ;
      RECT 40.565 1.07 40.58 1.328 ;
      RECT 40.525 1.085 40.565 1.332 ;
      RECT 40.475 1.1 40.525 1.337 ;
      RECT 40.45 1.107 40.475 1.341 ;
      RECT 40.39 1.102 40.45 1.345 ;
      RECT 40.375 1.093 40.39 1.349 ;
      RECT 40.305 1.083 40.375 1.345 ;
      RECT 40.28 1.075 40.3 1.335 ;
      RECT 40.221 1.075 40.28 1.313 ;
      RECT 40.135 1.075 40.221 1.27 ;
      RECT 40.3 1.075 40.305 1.34 ;
      RECT 40.995 0.306 41.165 0.64 ;
      RECT 40.965 0.306 41.165 0.635 ;
      RECT 40.905 0.273 40.965 0.623 ;
      RECT 40.905 0.329 41.175 0.618 ;
      RECT 40.88 0.329 41.175 0.612 ;
      RECT 40.875 0.27 40.905 0.609 ;
      RECT 40.86 0.276 40.995 0.607 ;
      RECT 40.855 0.284 41.08 0.595 ;
      RECT 40.855 0.336 41.19 0.548 ;
      RECT 40.84 0.292 41.08 0.543 ;
      RECT 40.84 0.362 41.2 0.484 ;
      RECT 40.81 0.312 41.165 0.445 ;
      RECT 40.81 0.402 41.21 0.441 ;
      RECT 40.86 0.281 41.08 0.607 ;
      RECT 40.2 0.611 40.255 0.875 ;
      RECT 40.2 0.611 40.32 0.874 ;
      RECT 40.2 0.611 40.345 0.873 ;
      RECT 40.2 0.611 40.41 0.872 ;
      RECT 40.345 0.577 40.425 0.871 ;
      RECT 40.16 0.621 40.57 0.87 ;
      RECT 40.2 0.618 40.57 0.87 ;
      RECT 40.16 0.626 40.575 0.863 ;
      RECT 40.145 0.628 40.575 0.862 ;
      RECT 40.145 0.635 40.58 0.858 ;
      RECT 40.125 0.634 40.575 0.854 ;
      RECT 40.125 0.642 40.585 0.853 ;
      RECT 40.12 0.639 40.58 0.849 ;
      RECT 40.12 0.652 40.595 0.848 ;
      RECT 40.105 0.642 40.585 0.847 ;
      RECT 40.07 0.655 40.595 0.84 ;
      RECT 40.255 0.61 40.565 0.87 ;
      RECT 40.255 0.595 40.515 0.87 ;
      RECT 40.32 0.582 40.45 0.87 ;
      RECT 39.865 1.671 39.88 2.064 ;
      RECT 39.83 1.676 39.88 2.063 ;
      RECT 39.865 1.675 39.925 2.062 ;
      RECT 39.81 1.686 39.925 2.061 ;
      RECT 39.825 1.682 39.925 2.061 ;
      RECT 39.79 1.692 40 2.058 ;
      RECT 39.79 1.711 40.045 2.056 ;
      RECT 39.79 1.718 40.05 2.053 ;
      RECT 39.775 1.695 40 2.05 ;
      RECT 39.755 1.7 40 2.043 ;
      RECT 39.75 1.704 40 2.039 ;
      RECT 39.75 1.721 40.06 2.038 ;
      RECT 39.73 1.715 40.045 2.034 ;
      RECT 39.73 1.724 40.065 2.028 ;
      RECT 39.725 1.73 40.065 1.8 ;
      RECT 39.79 1.69 39.925 2.058 ;
      RECT 39.665 1.053 39.865 1.365 ;
      RECT 39.74 1.031 39.865 1.365 ;
      RECT 39.68 1.05 39.87 1.35 ;
      RECT 39.65 1.061 39.87 1.348 ;
      RECT 39.665 1.056 39.875 1.314 ;
      RECT 39.65 1.16 39.88 1.281 ;
      RECT 39.68 1.032 39.865 1.365 ;
      RECT 39.74 1.01 39.84 1.365 ;
      RECT 39.765 1.007 39.84 1.365 ;
      RECT 39.765 1.002 39.785 1.365 ;
      RECT 39.17 1.07 39.345 1.245 ;
      RECT 39.165 1.07 39.345 1.243 ;
      RECT 39.14 1.07 39.345 1.238 ;
      RECT 39.085 1.05 39.255 1.228 ;
      RECT 39.085 1.057 39.32 1.228 ;
      RECT 39.17 1.737 39.185 1.92 ;
      RECT 39.16 1.715 39.17 1.92 ;
      RECT 39.145 1.695 39.16 1.92 ;
      RECT 39.135 1.67 39.145 1.92 ;
      RECT 39.105 1.635 39.135 1.92 ;
      RECT 39.07 1.575 39.105 1.92 ;
      RECT 39.065 1.537 39.07 1.92 ;
      RECT 39.015 1.488 39.065 1.92 ;
      RECT 39.005 1.438 39.015 1.908 ;
      RECT 38.99 1.417 39.005 1.868 ;
      RECT 38.97 1.385 38.99 1.818 ;
      RECT 38.945 1.341 38.97 1.758 ;
      RECT 38.94 1.313 38.945 1.713 ;
      RECT 38.935 1.304 38.94 1.699 ;
      RECT 38.93 1.297 38.935 1.686 ;
      RECT 38.925 1.292 38.93 1.675 ;
      RECT 38.92 1.277 38.925 1.665 ;
      RECT 38.915 1.255 38.92 1.652 ;
      RECT 38.905 1.215 38.915 1.627 ;
      RECT 38.88 1.145 38.905 1.583 ;
      RECT 38.875 1.085 38.88 1.548 ;
      RECT 38.86 1.065 38.875 1.515 ;
      RECT 38.855 1.065 38.86 1.49 ;
      RECT 38.825 1.065 38.855 1.445 ;
      RECT 38.78 1.065 38.825 1.385 ;
      RECT 38.705 1.065 38.78 1.333 ;
      RECT 38.7 1.065 38.705 1.298 ;
      RECT 38.695 1.065 38.7 1.288 ;
      RECT 38.69 1.065 38.695 1.268 ;
      RECT 38.955 0.285 39.125 0.755 ;
      RECT 38.9 0.278 39.095 0.739 ;
      RECT 38.9 0.292 39.13 0.738 ;
      RECT 38.885 0.293 39.13 0.719 ;
      RECT 38.88 0.311 39.13 0.705 ;
      RECT 38.885 0.294 39.135 0.703 ;
      RECT 38.87 0.325 39.135 0.688 ;
      RECT 38.885 0.3 39.14 0.673 ;
      RECT 38.865 0.34 39.14 0.67 ;
      RECT 38.88 0.312 39.145 0.655 ;
      RECT 38.88 0.324 39.15 0.635 ;
      RECT 38.865 0.34 39.155 0.618 ;
      RECT 38.865 0.35 39.16 0.473 ;
      RECT 38.86 0.35 39.16 0.43 ;
      RECT 38.86 0.365 39.165 0.408 ;
      RECT 38.955 0.275 39.095 0.755 ;
      RECT 38.955 0.273 39.065 0.755 ;
      RECT 39.041 0.27 39.065 0.755 ;
      RECT 38.7 1.937 38.705 1.983 ;
      RECT 38.69 1.785 38.7 2.007 ;
      RECT 38.685 1.63 38.69 2.032 ;
      RECT 38.67 1.592 38.685 2.043 ;
      RECT 38.665 1.575 38.67 2.05 ;
      RECT 38.655 1.563 38.665 2.057 ;
      RECT 38.65 1.554 38.655 2.059 ;
      RECT 38.645 1.552 38.65 2.063 ;
      RECT 38.6 1.543 38.645 2.078 ;
      RECT 38.595 1.535 38.6 2.092 ;
      RECT 38.59 1.532 38.595 2.096 ;
      RECT 38.575 1.527 38.59 2.104 ;
      RECT 38.52 1.517 38.575 2.115 ;
      RECT 38.485 1.505 38.52 2.116 ;
      RECT 38.476 1.5 38.485 2.11 ;
      RECT 38.39 1.5 38.476 2.1 ;
      RECT 38.36 1.5 38.39 2.078 ;
      RECT 38.35 1.5 38.355 2.058 ;
      RECT 38.345 1.5 38.35 2.02 ;
      RECT 38.34 1.5 38.345 1.978 ;
      RECT 38.335 1.5 38.34 1.938 ;
      RECT 38.33 1.5 38.335 1.868 ;
      RECT 38.32 1.5 38.33 1.79 ;
      RECT 38.315 1.5 38.32 1.69 ;
      RECT 38.355 1.5 38.36 2.06 ;
      RECT 37.85 1.582 37.94 2.06 ;
      RECT 37.835 1.585 37.955 2.058 ;
      RECT 37.85 1.584 37.955 2.058 ;
      RECT 37.815 1.591 37.98 2.048 ;
      RECT 37.835 1.585 37.98 2.048 ;
      RECT 37.8 1.597 37.98 2.036 ;
      RECT 37.835 1.588 38.03 2.029 ;
      RECT 37.786 1.605 38.03 2.027 ;
      RECT 37.815 1.595 38.04 2.015 ;
      RECT 37.786 1.616 38.07 2.006 ;
      RECT 37.7 1.64 38.07 2 ;
      RECT 37.7 1.653 38.11 1.983 ;
      RECT 37.695 1.675 38.11 1.976 ;
      RECT 37.665 1.69 38.11 1.966 ;
      RECT 37.66 1.701 38.11 1.956 ;
      RECT 37.63 1.714 38.11 1.947 ;
      RECT 37.615 1.732 38.11 1.936 ;
      RECT 37.59 1.745 38.11 1.926 ;
      RECT 37.85 1.581 37.86 2.06 ;
      RECT 37.896 1.005 37.935 1.25 ;
      RECT 37.81 1.005 37.945 1.248 ;
      RECT 37.695 1.03 37.945 1.245 ;
      RECT 37.695 1.03 37.95 1.243 ;
      RECT 37.695 1.03 37.965 1.238 ;
      RECT 37.801 1.005 37.98 1.218 ;
      RECT 37.715 1.013 37.98 1.218 ;
      RECT 37.385 0.365 37.555 0.8 ;
      RECT 37.375 0.399 37.555 0.783 ;
      RECT 37.455 0.335 37.625 0.77 ;
      RECT 37.36 0.41 37.625 0.748 ;
      RECT 37.455 0.345 37.63 0.738 ;
      RECT 37.385 0.397 37.66 0.723 ;
      RECT 37.345 0.423 37.66 0.708 ;
      RECT 37.345 0.465 37.67 0.688 ;
      RECT 37.34 0.49 37.675 0.67 ;
      RECT 37.34 0.5 37.68 0.655 ;
      RECT 37.335 0.437 37.66 0.653 ;
      RECT 37.335 0.51 37.685 0.638 ;
      RECT 37.33 0.447 37.66 0.635 ;
      RECT 37.325 0.531 37.69 0.618 ;
      RECT 37.325 0.563 37.695 0.598 ;
      RECT 37.32 0.477 37.67 0.59 ;
      RECT 37.325 0.462 37.66 0.618 ;
      RECT 37.34 0.432 37.66 0.67 ;
      RECT 37.185 1.019 37.41 1.275 ;
      RECT 37.185 1.052 37.43 1.265 ;
      RECT 37.15 1.052 37.43 1.263 ;
      RECT 37.15 1.065 37.435 1.253 ;
      RECT 37.15 1.085 37.445 1.245 ;
      RECT 37.15 1.182 37.45 1.238 ;
      RECT 37.13 0.93 37.26 1.228 ;
      RECT 37.085 1.085 37.445 1.17 ;
      RECT 37.075 0.93 37.26 1.115 ;
      RECT 37.075 0.962 37.346 1.115 ;
      RECT 37.04 1.492 37.06 1.67 ;
      RECT 37.005 1.445 37.04 1.67 ;
      RECT 36.99 1.385 37.005 1.67 ;
      RECT 36.965 1.332 36.99 1.67 ;
      RECT 36.95 1.285 36.965 1.67 ;
      RECT 36.93 1.262 36.95 1.67 ;
      RECT 36.905 1.227 36.93 1.67 ;
      RECT 36.895 1.073 36.905 1.67 ;
      RECT 36.865 1.068 36.895 1.661 ;
      RECT 36.86 1.065 36.865 1.651 ;
      RECT 36.845 1.065 36.86 1.625 ;
      RECT 36.84 1.065 36.845 1.588 ;
      RECT 36.815 1.065 36.84 1.54 ;
      RECT 36.795 1.065 36.815 1.465 ;
      RECT 36.785 1.065 36.795 1.425 ;
      RECT 36.78 1.065 36.785 1.4 ;
      RECT 36.775 1.065 36.78 1.383 ;
      RECT 36.77 1.065 36.775 1.365 ;
      RECT 36.765 1.066 36.77 1.355 ;
      RECT 36.755 1.068 36.765 1.323 ;
      RECT 36.745 1.07 36.755 1.29 ;
      RECT 36.735 1.073 36.745 1.263 ;
      RECT 37.06 1.5 37.285 1.67 ;
      RECT 36.39 0.312 36.56 0.765 ;
      RECT 36.39 0.312 36.65 0.731 ;
      RECT 36.39 0.312 36.68 0.715 ;
      RECT 36.39 0.312 36.71 0.688 ;
      RECT 36.646 0.29 36.725 0.67 ;
      RECT 36.425 0.297 36.73 0.655 ;
      RECT 36.425 0.305 36.74 0.618 ;
      RECT 36.385 0.332 36.74 0.59 ;
      RECT 36.37 0.345 36.74 0.555 ;
      RECT 36.39 0.32 36.76 0.545 ;
      RECT 36.365 0.385 36.76 0.515 ;
      RECT 36.365 0.415 36.765 0.498 ;
      RECT 36.36 0.445 36.765 0.485 ;
      RECT 36.425 0.294 36.725 0.67 ;
      RECT 36.56 0.291 36.646 0.749 ;
      RECT 36.511 0.292 36.725 0.67 ;
      RECT 36.655 1.952 36.7 2.145 ;
      RECT 36.645 1.922 36.655 2.145 ;
      RECT 36.64 1.907 36.645 2.145 ;
      RECT 36.6 1.817 36.64 2.145 ;
      RECT 36.595 1.73 36.6 2.145 ;
      RECT 36.585 1.7 36.595 2.145 ;
      RECT 36.58 1.66 36.585 2.145 ;
      RECT 36.57 1.622 36.58 2.145 ;
      RECT 36.565 1.587 36.57 2.145 ;
      RECT 36.545 1.54 36.565 2.145 ;
      RECT 36.53 1.465 36.545 2.145 ;
      RECT 36.525 1.42 36.53 2.14 ;
      RECT 36.52 1.4 36.525 2.113 ;
      RECT 36.515 1.38 36.52 2.098 ;
      RECT 36.51 1.355 36.515 2.078 ;
      RECT 36.505 1.333 36.51 2.063 ;
      RECT 36.5 1.311 36.505 2.045 ;
      RECT 36.495 1.29 36.5 2.035 ;
      RECT 36.485 1.262 36.495 2.005 ;
      RECT 36.475 1.225 36.485 1.973 ;
      RECT 36.465 1.185 36.475 1.94 ;
      RECT 36.455 1.163 36.465 1.91 ;
      RECT 36.425 1.115 36.455 1.842 ;
      RECT 36.41 1.075 36.425 1.769 ;
      RECT 36.4 1.075 36.41 1.735 ;
      RECT 36.395 1.075 36.4 1.71 ;
      RECT 36.39 1.075 36.395 1.695 ;
      RECT 36.385 1.075 36.39 1.673 ;
      RECT 36.38 1.075 36.385 1.66 ;
      RECT 36.365 1.075 36.38 1.625 ;
      RECT 36.345 1.075 36.365 1.565 ;
      RECT 36.335 1.075 36.345 1.515 ;
      RECT 36.315 1.075 36.335 1.463 ;
      RECT 36.295 1.075 36.315 1.42 ;
      RECT 36.285 1.075 36.295 1.408 ;
      RECT 36.255 1.075 36.285 1.395 ;
      RECT 36.225 1.096 36.255 1.375 ;
      RECT 36.215 1.124 36.225 1.355 ;
      RECT 36.2 1.141 36.215 1.323 ;
      RECT 36.195 1.155 36.2 1.29 ;
      RECT 36.19 1.163 36.195 1.263 ;
      RECT 36.185 1.171 36.19 1.225 ;
      RECT 36.19 1.695 36.195 2.03 ;
      RECT 36.155 1.682 36.19 2.029 ;
      RECT 36.085 1.622 36.155 2.028 ;
      RECT 36.005 1.565 36.085 2.027 ;
      RECT 35.87 1.525 36.005 2.026 ;
      RECT 35.87 1.712 36.205 2.015 ;
      RECT 35.83 1.712 36.205 2.005 ;
      RECT 35.83 1.73 36.21 2 ;
      RECT 35.83 1.82 36.215 1.99 ;
      RECT 35.825 1.515 35.99 1.97 ;
      RECT 35.82 1.515 35.99 1.713 ;
      RECT 35.82 1.672 36.185 1.713 ;
      RECT 35.82 1.66 36.18 1.713 ;
      RECT 35.085 1.875 35.6 2.285 ;
      RECT 35.26 0.895 35.6 2.285 ;
      RECT 34.37 0.895 35.6 1.065 ;
      RECT 35.08 0.29 35.325 1.065 ;
      RECT 32.48 2.295 34.51 2.465 ;
      RECT 34.34 1.44 34.51 2.465 ;
      RECT 32.48 0.995 32.65 2.465 ;
      RECT 34.34 1.44 35.09 1.63 ;
      RECT 32.455 0.995 32.65 1.325 ;
      RECT 33.16 1.615 34.17 1.785 ;
      RECT 33.98 0.255 34.17 1.785 ;
      RECT 33.16 0.815 33.33 1.785 ;
      RECT 32.82 1.955 33.945 2.125 ;
      RECT 32.82 0.255 32.99 2.125 ;
      RECT 31.975 0.995 32.23 1.325 ;
      RECT 32.06 0.655 32.23 1.325 ;
      RECT 32.06 0.655 32.99 0.825 ;
      RECT 32.815 0.255 32.99 0.825 ;
      RECT 32.815 0.255 33.345 0.62 ;
      RECT 31.635 1.495 31.97 2.465 ;
      RECT 31.635 0.255 31.805 2.465 ;
      RECT 31.635 0.255 31.89 0.825 ;
      RECT 30.885 1.485 31.215 2.465 ;
      RECT 30.985 0.255 31.215 2.465 ;
      RECT 30.885 1.855 31.345 2.015 ;
      RECT 30.885 0.255 31.215 0.885 ;
      RECT 29.505 1.485 29.835 2.465 ;
      RECT 29.605 0.255 29.835 2.465 ;
      RECT 29.605 1.075 30.815 1.315 ;
      RECT 29.505 0.255 29.835 0.885 ;
      RECT 28.125 1.485 28.455 2.465 ;
      RECT 28.225 0.255 28.455 2.465 ;
      RECT 28.125 1.515 28.59 1.69 ;
      RECT 28.125 0.255 28.455 0.885 ;
      RECT 26.745 1.485 27.075 2.465 ;
      RECT 26.845 0.255 27.075 2.465 ;
      RECT 26.845 1.075 28.055 1.315 ;
      RECT 26.745 0.255 27.075 0.885 ;
      RECT 25.425 1.875 25.94 2.285 ;
      RECT 25.6 0.895 25.94 2.285 ;
      RECT 24.71 0.895 25.94 1.065 ;
      RECT 25.42 0.29 25.665 1.065 ;
      RECT 22.82 2.295 24.85 2.465 ;
      RECT 24.68 1.44 24.85 2.465 ;
      RECT 22.82 0.995 22.99 2.465 ;
      RECT 24.68 1.44 25.43 1.63 ;
      RECT 22.795 0.995 22.99 1.325 ;
      RECT 23.5 1.615 24.51 1.785 ;
      RECT 24.32 0.255 24.51 1.785 ;
      RECT 23.5 0.815 23.67 1.785 ;
      RECT 23.16 1.955 24.285 2.125 ;
      RECT 23.16 0.255 23.33 2.125 ;
      RECT 22.315 0.995 22.57 1.325 ;
      RECT 22.4 0.655 22.57 1.325 ;
      RECT 22.4 0.655 23.33 0.825 ;
      RECT 23.155 0.255 23.33 0.825 ;
      RECT 23.155 0.255 23.685 0.62 ;
      RECT 21.975 1.495 22.31 2.465 ;
      RECT 21.975 0.255 22.145 2.465 ;
      RECT 21.975 0.255 22.23 0.825 ;
      RECT 21.29 1.875 21.805 2.285 ;
      RECT 21.465 0.895 21.805 2.285 ;
      RECT 20.575 0.895 21.805 1.065 ;
      RECT 21.285 0.29 21.53 1.065 ;
      RECT 18.685 2.295 20.715 2.465 ;
      RECT 20.545 1.44 20.715 2.465 ;
      RECT 18.685 0.995 18.855 2.465 ;
      RECT 20.545 1.44 21.295 1.63 ;
      RECT 18.66 0.995 18.855 1.325 ;
      RECT 19.365 1.615 20.375 1.785 ;
      RECT 20.185 0.255 20.375 1.785 ;
      RECT 19.365 0.815 19.535 1.785 ;
      RECT 19.025 1.955 20.15 2.125 ;
      RECT 19.025 0.255 19.195 2.125 ;
      RECT 18.18 0.995 18.435 1.325 ;
      RECT 18.265 0.655 18.435 1.325 ;
      RECT 18.265 0.655 19.195 0.825 ;
      RECT 19.02 0.255 19.195 0.825 ;
      RECT 19.02 0.255 19.55 0.62 ;
      RECT 17.84 1.495 18.175 2.465 ;
      RECT 17.84 0.255 18.01 2.465 ;
      RECT 17.84 0.255 18.095 0.825 ;
      RECT 16.745 0.475 17.475 0.715 ;
      RECT 17.287 0.27 17.475 0.715 ;
      RECT 17.115 0.282 17.49 0.709 ;
      RECT 17.03 0.297 17.51 0.694 ;
      RECT 17.03 0.312 17.515 0.684 ;
      RECT 16.985 0.332 17.53 0.676 ;
      RECT 16.962 0.367 17.545 0.63 ;
      RECT 16.876 0.39 17.55 0.59 ;
      RECT 16.876 0.408 17.56 0.56 ;
      RECT 16.745 0.477 17.565 0.523 ;
      RECT 16.79 0.42 17.56 0.56 ;
      RECT 16.876 0.372 17.545 0.63 ;
      RECT 16.962 0.341 17.53 0.676 ;
      RECT 16.985 0.322 17.515 0.684 ;
      RECT 17.03 0.295 17.49 0.709 ;
      RECT 17.115 0.277 17.475 0.715 ;
      RECT 17.201 0.271 17.475 0.715 ;
      RECT 17.287 0.266 17.42 0.715 ;
      RECT 17.373 0.261 17.42 0.715 ;
      RECT 17.065 1.159 17.235 1.545 ;
      RECT 17.06 1.159 17.235 1.54 ;
      RECT 17.035 1.159 17.235 1.505 ;
      RECT 17.035 1.187 17.245 1.495 ;
      RECT 17.015 1.187 17.245 1.455 ;
      RECT 17.01 1.187 17.245 1.428 ;
      RECT 17.01 1.205 17.25 1.42 ;
      RECT 16.955 1.205 17.25 1.355 ;
      RECT 16.955 1.222 17.26 1.338 ;
      RECT 16.945 1.222 17.26 1.278 ;
      RECT 16.945 1.239 17.265 1.275 ;
      RECT 16.94 1.075 17.11 1.253 ;
      RECT 16.94 1.109 17.196 1.253 ;
      RECT 16.935 1.875 16.94 1.888 ;
      RECT 16.93 1.77 16.935 1.893 ;
      RECT 16.905 1.63 16.93 1.908 ;
      RECT 16.87 1.581 16.905 1.94 ;
      RECT 16.865 1.549 16.87 1.96 ;
      RECT 16.86 1.54 16.865 1.96 ;
      RECT 16.78 1.505 16.86 1.96 ;
      RECT 16.717 1.475 16.78 1.96 ;
      RECT 16.631 1.463 16.717 1.96 ;
      RECT 16.545 1.449 16.631 1.96 ;
      RECT 16.465 1.436 16.545 1.946 ;
      RECT 16.43 1.428 16.465 1.926 ;
      RECT 16.42 1.425 16.43 1.917 ;
      RECT 16.39 1.42 16.42 1.904 ;
      RECT 16.34 1.395 16.39 1.88 ;
      RECT 16.326 1.369 16.34 1.862 ;
      RECT 16.24 1.329 16.326 1.838 ;
      RECT 16.195 1.277 16.24 1.807 ;
      RECT 16.185 1.252 16.195 1.794 ;
      RECT 16.18 1.033 16.185 1.055 ;
      RECT 16.175 1.235 16.185 1.79 ;
      RECT 16.175 1.031 16.18 1.145 ;
      RECT 16.165 1.027 16.175 1.786 ;
      RECT 16.121 1.025 16.165 1.774 ;
      RECT 16.035 1.025 16.121 1.745 ;
      RECT 16.005 1.025 16.035 1.718 ;
      RECT 15.99 1.025 16.005 1.706 ;
      RECT 15.95 1.037 15.99 1.691 ;
      RECT 15.93 1.056 15.95 1.67 ;
      RECT 15.92 1.066 15.93 1.654 ;
      RECT 15.91 1.072 15.92 1.643 ;
      RECT 15.89 1.082 15.91 1.626 ;
      RECT 15.885 1.091 15.89 1.613 ;
      RECT 15.88 1.095 15.885 1.563 ;
      RECT 15.87 1.101 15.88 1.48 ;
      RECT 15.865 1.105 15.87 1.394 ;
      RECT 15.86 1.125 15.865 1.331 ;
      RECT 15.855 1.148 15.86 1.278 ;
      RECT 15.85 1.166 15.855 1.223 ;
      RECT 16.46 0.985 16.63 1.245 ;
      RECT 16.63 0.95 16.675 1.231 ;
      RECT 16.591 0.952 16.68 1.214 ;
      RECT 16.48 0.969 16.766 1.185 ;
      RECT 16.48 0.984 16.77 1.157 ;
      RECT 16.48 0.965 16.68 1.214 ;
      RECT 16.505 0.953 16.63 1.245 ;
      RECT 16.591 0.951 16.675 1.231 ;
      RECT 15.645 0.34 15.815 0.83 ;
      RECT 15.645 0.34 15.85 0.81 ;
      RECT 15.78 0.26 15.89 0.77 ;
      RECT 15.761 0.264 15.91 0.74 ;
      RECT 15.675 0.272 15.93 0.723 ;
      RECT 15.675 0.278 15.935 0.713 ;
      RECT 15.675 0.287 15.955 0.701 ;
      RECT 15.65 0.312 15.985 0.679 ;
      RECT 15.65 0.332 15.99 0.659 ;
      RECT 15.645 0.345 16 0.639 ;
      RECT 15.645 0.412 16.005 0.62 ;
      RECT 15.645 0.545 16.01 0.607 ;
      RECT 15.64 0.35 16 0.44 ;
      RECT 15.65 0.307 15.955 0.701 ;
      RECT 15.761 0.262 15.89 0.77 ;
      RECT 15.635 2.015 15.935 2.27 ;
      RECT 15.72 1.981 15.935 2.27 ;
      RECT 15.72 1.984 15.94 2.13 ;
      RECT 15.655 2.005 15.94 2.13 ;
      RECT 15.69 1.995 15.935 2.27 ;
      RECT 15.685 2 15.94 2.13 ;
      RECT 15.72 1.979 15.921 2.27 ;
      RECT 15.806 1.97 15.921 2.27 ;
      RECT 15.806 1.964 15.835 2.27 ;
      RECT 15.295 1.605 15.305 2.095 ;
      RECT 14.955 1.54 14.965 1.84 ;
      RECT 15.47 1.712 15.475 1.931 ;
      RECT 15.46 1.692 15.47 1.948 ;
      RECT 15.45 1.672 15.46 1.978 ;
      RECT 15.445 1.662 15.45 1.993 ;
      RECT 15.44 1.658 15.445 1.998 ;
      RECT 15.425 1.65 15.44 2.005 ;
      RECT 15.385 1.63 15.425 2.03 ;
      RECT 15.36 1.612 15.385 2.063 ;
      RECT 15.355 1.61 15.36 2.076 ;
      RECT 15.335 1.607 15.355 2.08 ;
      RECT 15.305 1.605 15.335 2.09 ;
      RECT 15.235 1.607 15.295 2.091 ;
      RECT 15.215 1.607 15.235 2.085 ;
      RECT 15.19 1.605 15.215 2.082 ;
      RECT 15.155 1.6 15.19 2.078 ;
      RECT 15.135 1.594 15.155 2.065 ;
      RECT 15.125 1.591 15.135 2.053 ;
      RECT 15.105 1.588 15.125 2.038 ;
      RECT 15.085 1.584 15.105 2.02 ;
      RECT 15.08 1.581 15.085 2.01 ;
      RECT 15.075 1.58 15.08 2.008 ;
      RECT 15.065 1.577 15.075 2 ;
      RECT 15.055 1.571 15.065 1.983 ;
      RECT 15.045 1.565 15.055 1.965 ;
      RECT 15.035 1.559 15.045 1.953 ;
      RECT 15.025 1.553 15.035 1.933 ;
      RECT 15.02 1.549 15.025 1.918 ;
      RECT 15.015 1.547 15.02 1.91 ;
      RECT 15.01 1.545 15.015 1.903 ;
      RECT 15.005 1.543 15.01 1.893 ;
      RECT 15 1.541 15.005 1.887 ;
      RECT 14.99 1.54 15 1.877 ;
      RECT 14.98 1.54 14.99 1.868 ;
      RECT 14.965 1.54 14.98 1.853 ;
      RECT 14.925 1.54 14.955 1.837 ;
      RECT 14.905 1.542 14.925 1.832 ;
      RECT 14.9 1.547 14.905 1.83 ;
      RECT 14.87 1.555 14.9 1.828 ;
      RECT 14.84 1.57 14.87 1.827 ;
      RECT 14.795 1.592 14.84 1.832 ;
      RECT 14.79 1.607 14.795 1.836 ;
      RECT 14.775 1.612 14.79 1.838 ;
      RECT 14.77 1.616 14.775 1.84 ;
      RECT 14.71 1.639 14.77 1.849 ;
      RECT 14.69 1.665 14.71 1.862 ;
      RECT 14.68 1.672 14.69 1.866 ;
      RECT 14.665 1.679 14.68 1.869 ;
      RECT 14.645 1.689 14.665 1.872 ;
      RECT 14.64 1.697 14.645 1.875 ;
      RECT 14.595 1.702 14.64 1.882 ;
      RECT 14.585 1.705 14.595 1.889 ;
      RECT 14.575 1.705 14.585 1.893 ;
      RECT 14.54 1.707 14.575 1.905 ;
      RECT 14.52 1.71 14.54 1.918 ;
      RECT 14.48 1.713 14.52 1.929 ;
      RECT 14.465 1.715 14.48 1.942 ;
      RECT 14.455 1.715 14.465 1.947 ;
      RECT 14.43 1.716 14.455 1.955 ;
      RECT 14.42 1.718 14.43 1.96 ;
      RECT 14.415 1.719 14.42 1.963 ;
      RECT 14.39 1.717 14.415 1.966 ;
      RECT 14.375 1.715 14.39 1.967 ;
      RECT 14.355 1.712 14.375 1.969 ;
      RECT 14.335 1.707 14.355 1.969 ;
      RECT 14.275 1.702 14.335 1.966 ;
      RECT 14.24 1.677 14.275 1.962 ;
      RECT 14.23 1.654 14.24 1.96 ;
      RECT 14.2 1.631 14.23 1.96 ;
      RECT 14.19 1.61 14.2 1.96 ;
      RECT 14.165 1.592 14.19 1.958 ;
      RECT 14.15 1.57 14.165 1.955 ;
      RECT 14.135 1.552 14.15 1.953 ;
      RECT 14.115 1.542 14.135 1.951 ;
      RECT 14.1 1.537 14.115 1.95 ;
      RECT 14.085 1.535 14.1 1.949 ;
      RECT 14.055 1.536 14.085 1.947 ;
      RECT 14.035 1.539 14.055 1.945 ;
      RECT 13.978 1.543 14.035 1.945 ;
      RECT 13.892 1.552 13.978 1.945 ;
      RECT 13.806 1.563 13.892 1.945 ;
      RECT 13.72 1.574 13.806 1.945 ;
      RECT 13.7 1.581 13.72 1.953 ;
      RECT 13.69 1.584 13.7 1.96 ;
      RECT 13.625 1.589 13.69 1.978 ;
      RECT 13.595 1.596 13.625 2.003 ;
      RECT 13.585 1.599 13.595 2.01 ;
      RECT 13.54 1.603 13.585 2.015 ;
      RECT 13.51 1.608 13.54 2.02 ;
      RECT 13.509 1.61 13.51 2.02 ;
      RECT 13.423 1.616 13.509 2.02 ;
      RECT 13.337 1.627 13.423 2.02 ;
      RECT 13.251 1.639 13.337 2.02 ;
      RECT 13.165 1.65 13.251 2.02 ;
      RECT 13.15 1.657 13.165 2.015 ;
      RECT 13.145 1.659 13.15 2.009 ;
      RECT 13.125 1.67 13.145 2.004 ;
      RECT 13.115 1.688 13.125 1.998 ;
      RECT 13.11 1.7 13.115 1.798 ;
      RECT 15.405 0.453 15.425 0.54 ;
      RECT 15.4 0.388 15.405 0.572 ;
      RECT 15.39 0.355 15.4 0.577 ;
      RECT 15.385 0.335 15.39 0.583 ;
      RECT 15.355 0.335 15.385 0.6 ;
      RECT 15.306 0.335 15.355 0.636 ;
      RECT 15.22 0.335 15.306 0.694 ;
      RECT 15.191 0.345 15.22 0.743 ;
      RECT 15.105 0.387 15.191 0.796 ;
      RECT 15.085 0.425 15.105 0.843 ;
      RECT 15.06 0.442 15.085 0.863 ;
      RECT 15.05 0.456 15.06 0.883 ;
      RECT 15.045 0.462 15.05 0.893 ;
      RECT 15.04 0.466 15.045 0.9 ;
      RECT 14.99 0.486 15.04 0.905 ;
      RECT 14.925 0.53 14.99 0.905 ;
      RECT 14.9 0.58 14.925 0.905 ;
      RECT 14.89 0.61 14.9 0.905 ;
      RECT 14.885 0.637 14.89 0.905 ;
      RECT 14.88 0.655 14.885 0.905 ;
      RECT 14.87 0.697 14.88 0.905 ;
      RECT 15.22 1.255 15.39 1.43 ;
      RECT 15.16 1.083 15.22 1.418 ;
      RECT 15.15 1.076 15.16 1.401 ;
      RECT 15.105 1.255 15.39 1.381 ;
      RECT 15.086 1.255 15.39 1.359 ;
      RECT 15 1.255 15.39 1.324 ;
      RECT 14.98 1.075 15.15 1.28 ;
      RECT 14.98 1.222 15.385 1.28 ;
      RECT 14.98 1.17 15.36 1.28 ;
      RECT 14.98 1.125 15.325 1.28 ;
      RECT 14.98 1.107 15.29 1.28 ;
      RECT 14.98 1.097 15.285 1.28 ;
      RECT 14.7 2.055 14.89 2.28 ;
      RECT 14.69 2.056 14.895 2.275 ;
      RECT 14.69 2.058 14.905 2.255 ;
      RECT 14.69 2.062 14.91 2.24 ;
      RECT 14.69 2.049 14.86 2.275 ;
      RECT 14.69 2.052 14.885 2.275 ;
      RECT 14.7 2.048 14.86 2.28 ;
      RECT 14.786 2.046 14.86 2.28 ;
      RECT 14.41 1.297 14.58 1.535 ;
      RECT 14.41 1.297 14.666 1.449 ;
      RECT 14.41 1.297 14.67 1.359 ;
      RECT 14.46 1.07 14.68 1.338 ;
      RECT 14.455 1.087 14.685 1.311 ;
      RECT 14.42 1.245 14.685 1.311 ;
      RECT 14.44 1.095 14.58 1.535 ;
      RECT 14.43 1.177 14.69 1.294 ;
      RECT 14.425 1.225 14.69 1.294 ;
      RECT 14.43 1.135 14.685 1.311 ;
      RECT 14.455 1.072 14.68 1.338 ;
      RECT 14.02 1.047 14.19 1.245 ;
      RECT 14.02 1.047 14.235 1.22 ;
      RECT 14.09 0.99 14.26 1.178 ;
      RECT 14.065 1.005 14.26 1.178 ;
      RECT 13.68 1.051 13.71 1.245 ;
      RECT 13.675 1.023 13.68 1.245 ;
      RECT 13.645 0.997 13.675 1.247 ;
      RECT 13.62 0.955 13.645 1.25 ;
      RECT 13.61 0.927 13.62 1.252 ;
      RECT 13.575 0.907 13.61 1.254 ;
      RECT 13.51 0.892 13.575 1.26 ;
      RECT 13.46 0.89 13.51 1.266 ;
      RECT 13.437 0.892 13.46 1.271 ;
      RECT 13.351 0.903 13.437 1.277 ;
      RECT 13.265 0.921 13.351 1.287 ;
      RECT 13.25 0.932 13.265 1.293 ;
      RECT 13.18 0.955 13.25 1.299 ;
      RECT 13.125 0.987 13.18 1.307 ;
      RECT 13.085 1.01 13.125 1.313 ;
      RECT 13.071 1.023 13.085 1.316 ;
      RECT 12.985 1.045 13.071 1.322 ;
      RECT 12.97 1.07 12.985 1.328 ;
      RECT 12.93 1.085 12.97 1.332 ;
      RECT 12.88 1.1 12.93 1.337 ;
      RECT 12.855 1.107 12.88 1.341 ;
      RECT 12.795 1.102 12.855 1.345 ;
      RECT 12.78 1.093 12.795 1.349 ;
      RECT 12.71 1.083 12.78 1.345 ;
      RECT 12.685 1.075 12.705 1.335 ;
      RECT 12.626 1.075 12.685 1.313 ;
      RECT 12.54 1.075 12.626 1.27 ;
      RECT 12.705 1.075 12.71 1.34 ;
      RECT 13.4 0.306 13.57 0.64 ;
      RECT 13.37 0.306 13.57 0.635 ;
      RECT 13.31 0.273 13.37 0.623 ;
      RECT 13.31 0.329 13.58 0.618 ;
      RECT 13.285 0.329 13.58 0.612 ;
      RECT 13.28 0.27 13.31 0.609 ;
      RECT 13.265 0.276 13.4 0.607 ;
      RECT 13.26 0.284 13.485 0.595 ;
      RECT 13.26 0.336 13.595 0.548 ;
      RECT 13.245 0.292 13.485 0.543 ;
      RECT 13.245 0.362 13.605 0.484 ;
      RECT 13.215 0.312 13.57 0.445 ;
      RECT 13.215 0.402 13.615 0.441 ;
      RECT 13.265 0.281 13.485 0.607 ;
      RECT 12.605 0.611 12.66 0.875 ;
      RECT 12.605 0.611 12.725 0.874 ;
      RECT 12.605 0.611 12.75 0.873 ;
      RECT 12.605 0.611 12.815 0.872 ;
      RECT 12.75 0.577 12.83 0.871 ;
      RECT 12.565 0.621 12.975 0.87 ;
      RECT 12.605 0.618 12.975 0.87 ;
      RECT 12.565 0.626 12.98 0.863 ;
      RECT 12.55 0.628 12.98 0.862 ;
      RECT 12.55 0.635 12.985 0.858 ;
      RECT 12.53 0.634 12.98 0.854 ;
      RECT 12.53 0.642 12.99 0.853 ;
      RECT 12.525 0.639 12.985 0.849 ;
      RECT 12.525 0.652 13 0.848 ;
      RECT 12.51 0.642 12.99 0.847 ;
      RECT 12.475 0.655 13 0.84 ;
      RECT 12.66 0.61 12.97 0.87 ;
      RECT 12.66 0.595 12.92 0.87 ;
      RECT 12.725 0.582 12.855 0.87 ;
      RECT 12.27 1.671 12.285 2.064 ;
      RECT 12.235 1.676 12.285 2.063 ;
      RECT 12.27 1.675 12.33 2.062 ;
      RECT 12.215 1.686 12.33 2.061 ;
      RECT 12.23 1.682 12.33 2.061 ;
      RECT 12.195 1.692 12.405 2.058 ;
      RECT 12.195 1.711 12.45 2.056 ;
      RECT 12.195 1.718 12.455 2.053 ;
      RECT 12.18 1.695 12.405 2.05 ;
      RECT 12.16 1.7 12.405 2.043 ;
      RECT 12.155 1.704 12.405 2.039 ;
      RECT 12.155 1.721 12.465 2.038 ;
      RECT 12.135 1.715 12.45 2.034 ;
      RECT 12.135 1.724 12.47 2.028 ;
      RECT 12.13 1.73 12.47 1.8 ;
      RECT 12.195 1.69 12.33 2.058 ;
      RECT 12.07 1.053 12.27 1.365 ;
      RECT 12.145 1.031 12.27 1.365 ;
      RECT 12.085 1.05 12.275 1.35 ;
      RECT 12.055 1.061 12.275 1.348 ;
      RECT 12.07 1.056 12.28 1.314 ;
      RECT 12.055 1.16 12.285 1.281 ;
      RECT 12.085 1.032 12.27 1.365 ;
      RECT 12.145 1.01 12.245 1.365 ;
      RECT 12.17 1.007 12.245 1.365 ;
      RECT 12.17 1.002 12.19 1.365 ;
      RECT 11.575 1.07 11.75 1.245 ;
      RECT 11.57 1.07 11.75 1.243 ;
      RECT 11.545 1.07 11.75 1.238 ;
      RECT 11.49 1.05 11.66 1.228 ;
      RECT 11.49 1.057 11.725 1.228 ;
      RECT 11.575 1.737 11.59 1.92 ;
      RECT 11.565 1.715 11.575 1.92 ;
      RECT 11.55 1.695 11.565 1.92 ;
      RECT 11.54 1.67 11.55 1.92 ;
      RECT 11.51 1.635 11.54 1.92 ;
      RECT 11.475 1.575 11.51 1.92 ;
      RECT 11.47 1.537 11.475 1.92 ;
      RECT 11.42 1.488 11.47 1.92 ;
      RECT 11.41 1.438 11.42 1.908 ;
      RECT 11.395 1.417 11.41 1.868 ;
      RECT 11.375 1.385 11.395 1.818 ;
      RECT 11.35 1.341 11.375 1.758 ;
      RECT 11.345 1.313 11.35 1.713 ;
      RECT 11.34 1.304 11.345 1.699 ;
      RECT 11.335 1.297 11.34 1.686 ;
      RECT 11.33 1.292 11.335 1.675 ;
      RECT 11.325 1.277 11.33 1.665 ;
      RECT 11.32 1.255 11.325 1.652 ;
      RECT 11.31 1.215 11.32 1.627 ;
      RECT 11.285 1.145 11.31 1.583 ;
      RECT 11.28 1.085 11.285 1.548 ;
      RECT 11.265 1.065 11.28 1.515 ;
      RECT 11.26 1.065 11.265 1.49 ;
      RECT 11.23 1.065 11.26 1.445 ;
      RECT 11.185 1.065 11.23 1.385 ;
      RECT 11.11 1.065 11.185 1.333 ;
      RECT 11.105 1.065 11.11 1.298 ;
      RECT 11.1 1.065 11.105 1.288 ;
      RECT 11.095 1.065 11.1 1.268 ;
      RECT 11.36 0.285 11.53 0.755 ;
      RECT 11.305 0.278 11.5 0.739 ;
      RECT 11.305 0.292 11.535 0.738 ;
      RECT 11.29 0.293 11.535 0.719 ;
      RECT 11.285 0.311 11.535 0.705 ;
      RECT 11.29 0.294 11.54 0.703 ;
      RECT 11.275 0.325 11.54 0.688 ;
      RECT 11.29 0.3 11.545 0.673 ;
      RECT 11.27 0.34 11.545 0.67 ;
      RECT 11.285 0.312 11.55 0.655 ;
      RECT 11.285 0.324 11.555 0.635 ;
      RECT 11.27 0.34 11.56 0.618 ;
      RECT 11.27 0.35 11.565 0.473 ;
      RECT 11.265 0.35 11.565 0.43 ;
      RECT 11.265 0.365 11.57 0.408 ;
      RECT 11.36 0.275 11.5 0.755 ;
      RECT 11.36 0.273 11.47 0.755 ;
      RECT 11.446 0.27 11.47 0.755 ;
      RECT 11.105 1.937 11.11 1.983 ;
      RECT 11.095 1.785 11.105 2.007 ;
      RECT 11.09 1.63 11.095 2.032 ;
      RECT 11.075 1.592 11.09 2.043 ;
      RECT 11.07 1.575 11.075 2.05 ;
      RECT 11.06 1.563 11.07 2.057 ;
      RECT 11.055 1.554 11.06 2.059 ;
      RECT 11.05 1.552 11.055 2.063 ;
      RECT 11.005 1.543 11.05 2.078 ;
      RECT 11 1.535 11.005 2.092 ;
      RECT 10.995 1.532 11 2.096 ;
      RECT 10.98 1.527 10.995 2.104 ;
      RECT 10.925 1.517 10.98 2.115 ;
      RECT 10.89 1.505 10.925 2.116 ;
      RECT 10.881 1.5 10.89 2.11 ;
      RECT 10.795 1.5 10.881 2.1 ;
      RECT 10.765 1.5 10.795 2.078 ;
      RECT 10.755 1.5 10.76 2.058 ;
      RECT 10.75 1.5 10.755 2.02 ;
      RECT 10.745 1.5 10.75 1.978 ;
      RECT 10.74 1.5 10.745 1.938 ;
      RECT 10.735 1.5 10.74 1.868 ;
      RECT 10.725 1.5 10.735 1.79 ;
      RECT 10.72 1.5 10.725 1.69 ;
      RECT 10.76 1.5 10.765 2.06 ;
      RECT 10.255 1.582 10.345 2.06 ;
      RECT 10.24 1.585 10.36 2.058 ;
      RECT 10.255 1.584 10.36 2.058 ;
      RECT 10.22 1.591 10.385 2.048 ;
      RECT 10.24 1.585 10.385 2.048 ;
      RECT 10.205 1.597 10.385 2.036 ;
      RECT 10.24 1.588 10.435 2.029 ;
      RECT 10.191 1.605 10.435 2.027 ;
      RECT 10.22 1.595 10.445 2.015 ;
      RECT 10.191 1.616 10.475 2.006 ;
      RECT 10.105 1.64 10.475 2 ;
      RECT 10.105 1.653 10.515 1.983 ;
      RECT 10.1 1.675 10.515 1.976 ;
      RECT 10.07 1.69 10.515 1.966 ;
      RECT 10.065 1.701 10.515 1.956 ;
      RECT 10.035 1.714 10.515 1.947 ;
      RECT 10.02 1.732 10.515 1.936 ;
      RECT 9.995 1.745 10.515 1.926 ;
      RECT 10.255 1.581 10.265 2.06 ;
      RECT 10.301 1.005 10.34 1.25 ;
      RECT 10.215 1.005 10.35 1.248 ;
      RECT 10.1 1.03 10.35 1.245 ;
      RECT 10.1 1.03 10.355 1.243 ;
      RECT 10.1 1.03 10.37 1.238 ;
      RECT 10.206 1.005 10.385 1.218 ;
      RECT 10.12 1.013 10.385 1.218 ;
      RECT 9.79 0.365 9.96 0.8 ;
      RECT 9.78 0.399 9.96 0.783 ;
      RECT 9.86 0.335 10.03 0.77 ;
      RECT 9.765 0.41 10.03 0.748 ;
      RECT 9.86 0.345 10.035 0.738 ;
      RECT 9.79 0.397 10.065 0.723 ;
      RECT 9.75 0.423 10.065 0.708 ;
      RECT 9.75 0.465 10.075 0.688 ;
      RECT 9.745 0.49 10.08 0.67 ;
      RECT 9.745 0.5 10.085 0.655 ;
      RECT 9.74 0.437 10.065 0.653 ;
      RECT 9.74 0.51 10.09 0.638 ;
      RECT 9.735 0.447 10.065 0.635 ;
      RECT 9.73 0.531 10.095 0.618 ;
      RECT 9.73 0.563 10.1 0.598 ;
      RECT 9.725 0.477 10.075 0.59 ;
      RECT 9.73 0.462 10.065 0.618 ;
      RECT 9.745 0.432 10.065 0.67 ;
      RECT 9.59 1.019 9.815 1.275 ;
      RECT 9.59 1.052 9.835 1.265 ;
      RECT 9.555 1.052 9.835 1.263 ;
      RECT 9.555 1.065 9.84 1.253 ;
      RECT 9.555 1.085 9.85 1.245 ;
      RECT 9.555 1.182 9.855 1.238 ;
      RECT 9.535 0.93 9.665 1.228 ;
      RECT 9.49 1.085 9.85 1.17 ;
      RECT 9.48 0.93 9.665 1.115 ;
      RECT 9.48 0.962 9.751 1.115 ;
      RECT 9.445 1.492 9.465 1.67 ;
      RECT 9.41 1.445 9.445 1.67 ;
      RECT 9.395 1.385 9.41 1.67 ;
      RECT 9.37 1.332 9.395 1.67 ;
      RECT 9.355 1.285 9.37 1.67 ;
      RECT 9.335 1.262 9.355 1.67 ;
      RECT 9.31 1.227 9.335 1.67 ;
      RECT 9.3 1.073 9.31 1.67 ;
      RECT 9.27 1.068 9.3 1.661 ;
      RECT 9.265 1.065 9.27 1.651 ;
      RECT 9.25 1.065 9.265 1.625 ;
      RECT 9.245 1.065 9.25 1.588 ;
      RECT 9.22 1.065 9.245 1.54 ;
      RECT 9.2 1.065 9.22 1.465 ;
      RECT 9.19 1.065 9.2 1.425 ;
      RECT 9.185 1.065 9.19 1.4 ;
      RECT 9.18 1.065 9.185 1.383 ;
      RECT 9.175 1.065 9.18 1.365 ;
      RECT 9.17 1.066 9.175 1.355 ;
      RECT 9.16 1.068 9.17 1.323 ;
      RECT 9.15 1.07 9.16 1.29 ;
      RECT 9.14 1.073 9.15 1.263 ;
      RECT 9.465 1.5 9.69 1.67 ;
      RECT 8.795 0.312 8.965 0.765 ;
      RECT 8.795 0.312 9.055 0.731 ;
      RECT 8.795 0.312 9.085 0.715 ;
      RECT 8.795 0.312 9.115 0.688 ;
      RECT 9.051 0.29 9.13 0.67 ;
      RECT 8.83 0.297 9.135 0.655 ;
      RECT 8.83 0.305 9.145 0.618 ;
      RECT 8.79 0.332 9.145 0.59 ;
      RECT 8.775 0.345 9.145 0.555 ;
      RECT 8.795 0.32 9.165 0.545 ;
      RECT 8.77 0.385 9.165 0.515 ;
      RECT 8.77 0.415 9.17 0.498 ;
      RECT 8.765 0.445 9.17 0.485 ;
      RECT 8.83 0.294 9.13 0.67 ;
      RECT 8.965 0.291 9.051 0.749 ;
      RECT 8.916 0.292 9.13 0.67 ;
      RECT 9.06 1.952 9.105 2.145 ;
      RECT 9.05 1.922 9.06 2.145 ;
      RECT 9.045 1.907 9.05 2.145 ;
      RECT 9.005 1.817 9.045 2.145 ;
      RECT 9 1.73 9.005 2.145 ;
      RECT 8.99 1.7 9 2.145 ;
      RECT 8.985 1.66 8.99 2.145 ;
      RECT 8.975 1.622 8.985 2.145 ;
      RECT 8.97 1.587 8.975 2.145 ;
      RECT 8.95 1.54 8.97 2.145 ;
      RECT 8.935 1.465 8.95 2.145 ;
      RECT 8.93 1.42 8.935 2.14 ;
      RECT 8.925 1.4 8.93 2.113 ;
      RECT 8.92 1.38 8.925 2.098 ;
      RECT 8.915 1.355 8.92 2.078 ;
      RECT 8.91 1.333 8.915 2.063 ;
      RECT 8.905 1.311 8.91 2.045 ;
      RECT 8.9 1.29 8.905 2.035 ;
      RECT 8.89 1.262 8.9 2.005 ;
      RECT 8.88 1.225 8.89 1.973 ;
      RECT 8.87 1.185 8.88 1.94 ;
      RECT 8.86 1.163 8.87 1.91 ;
      RECT 8.83 1.115 8.86 1.842 ;
      RECT 8.815 1.075 8.83 1.769 ;
      RECT 8.805 1.075 8.815 1.735 ;
      RECT 8.8 1.075 8.805 1.71 ;
      RECT 8.795 1.075 8.8 1.695 ;
      RECT 8.79 1.075 8.795 1.673 ;
      RECT 8.785 1.075 8.79 1.66 ;
      RECT 8.77 1.075 8.785 1.625 ;
      RECT 8.75 1.075 8.77 1.565 ;
      RECT 8.74 1.075 8.75 1.515 ;
      RECT 8.72 1.075 8.74 1.463 ;
      RECT 8.7 1.075 8.72 1.42 ;
      RECT 8.69 1.075 8.7 1.408 ;
      RECT 8.66 1.075 8.69 1.395 ;
      RECT 8.63 1.096 8.66 1.375 ;
      RECT 8.62 1.124 8.63 1.355 ;
      RECT 8.605 1.141 8.62 1.323 ;
      RECT 8.6 1.155 8.605 1.29 ;
      RECT 8.595 1.163 8.6 1.263 ;
      RECT 8.59 1.171 8.595 1.225 ;
      RECT 8.595 1.695 8.6 2.03 ;
      RECT 8.56 1.682 8.595 2.029 ;
      RECT 8.49 1.622 8.56 2.028 ;
      RECT 8.41 1.565 8.49 2.027 ;
      RECT 8.275 1.525 8.41 2.026 ;
      RECT 8.275 1.712 8.61 2.015 ;
      RECT 8.235 1.712 8.61 2.005 ;
      RECT 8.235 1.73 8.615 2 ;
      RECT 8.235 1.82 8.62 1.99 ;
      RECT 8.23 1.515 8.395 1.97 ;
      RECT 8.225 1.515 8.395 1.713 ;
      RECT 8.225 1.672 8.59 1.713 ;
      RECT 8.225 1.66 8.585 1.713 ;
      RECT 7.49 1.875 8.005 2.285 ;
      RECT 7.665 0.895 8.005 2.285 ;
      RECT 6.775 0.895 8.005 1.065 ;
      RECT 7.485 0.29 7.73 1.065 ;
      RECT 4.885 2.295 6.915 2.465 ;
      RECT 6.745 1.44 6.915 2.465 ;
      RECT 4.885 0.995 5.055 2.465 ;
      RECT 6.745 1.44 7.495 1.63 ;
      RECT 4.86 0.995 5.055 1.325 ;
      RECT 5.565 1.615 6.575 1.785 ;
      RECT 6.385 0.255 6.575 1.785 ;
      RECT 5.565 0.815 5.735 1.785 ;
      RECT 5.225 1.955 6.35 2.125 ;
      RECT 5.225 0.255 5.395 2.125 ;
      RECT 4.38 0.995 4.635 1.325 ;
      RECT 4.465 0.655 4.635 1.325 ;
      RECT 4.465 0.655 5.395 0.825 ;
      RECT 5.22 0.255 5.395 0.825 ;
      RECT 5.22 0.255 5.75 0.62 ;
      RECT 4.04 1.495 4.375 2.465 ;
      RECT 3.54 1.875 4.375 2.285 ;
      RECT 3.715 0.895 4.21 2.285 ;
      RECT 2.825 0.895 4.21 1.065 ;
      RECT 3.535 0.29 3.78 1.065 ;
      RECT 4.04 0.255 4.21 2.465 ;
      RECT 4.04 0.255 4.295 0.825 ;
      RECT 0.935 2.295 2.965 2.465 ;
      RECT 2.795 1.44 2.965 2.465 ;
      RECT 0.935 0.995 1.105 2.465 ;
      RECT 2.795 1.44 3.545 1.63 ;
      RECT 0.91 0.995 1.105 1.325 ;
      RECT 2.455 0.255 2.625 1.87 ;
      RECT 1.615 1.615 2.625 1.785 ;
      RECT 2.435 0.255 2.625 1.785 ;
      RECT 1.615 0.815 1.785 1.785 ;
      RECT 1.275 1.955 2.4 2.125 ;
      RECT 1.275 0.255 1.445 2.125 ;
      RECT 0.43 0.995 0.685 1.325 ;
      RECT 0.515 0.655 0.685 1.325 ;
      RECT 0.515 0.655 1.445 0.825 ;
      RECT 1.27 0.255 1.445 0.825 ;
      RECT 1.27 0.255 1.8 0.62 ;
      RECT 0.09 1.495 0.425 2.465 ;
      RECT 0.09 0.255 0.26 2.465 ;
      RECT 0.09 0.255 0.345 0.825 ;
      RECT 139.485 1.075 139.815 1.315 ;
      RECT 136.725 1.075 137.055 1.315 ;
      RECT 134.255 0.255 134.53 1.415 ;
      RECT 130.12 0.255 130.395 1.415 ;
      RECT 117.815 1.7 117.985 1.87 ;
      RECT 111.89 1.075 112.22 1.315 ;
      RECT 109.13 1.075 109.46 1.315 ;
      RECT 106.66 0.255 106.935 1.415 ;
      RECT 102.525 0.255 102.8 1.415 ;
      RECT 90.22 1.7 90.39 1.87 ;
      RECT 84.295 1.075 84.625 1.315 ;
      RECT 81.535 1.075 81.865 1.315 ;
      RECT 79.065 0.255 79.34 1.415 ;
      RECT 74.93 0.255 75.205 1.415 ;
      RECT 62.625 1.7 62.795 1.87 ;
      RECT 56.7 1.075 57.03 1.315 ;
      RECT 53.94 1.075 54.27 1.315 ;
      RECT 51.47 0.255 51.745 1.415 ;
      RECT 47.335 0.255 47.61 1.415 ;
      RECT 35.03 1.7 35.2 1.87 ;
      RECT 29.105 1.075 29.435 1.315 ;
      RECT 26.345 1.075 26.675 1.315 ;
      RECT 23.875 0.255 24.15 1.415 ;
      RECT 19.74 0.255 20.015 1.415 ;
      RECT 7.435 1.7 7.605 1.87 ;
      RECT 3.115 1.68 3.24 1.87 ;
      RECT 1.99 0.255 2.265 1.415 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 4.14 1.65 ;
  SIZE 104.79 BY 7.63 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  OBS
    LAYER met4 ;
      RECT 84.755 -0.61 85.135 -0.23 ;
      RECT 95.51 -0.62 95.89 -0.24 ;
      RECT 84.755 -0.575 95.89 -0.27 ;
      RECT 89.245 4.855 89.67 5.28 ;
      RECT -0.01 4.85 0.415 5.275 ;
      RECT -0.01 4.91 89.67 5.23 ;
      RECT -0.015 4.905 0.415 5.225 ;
      RECT 66.815 -0.61 67.195 -0.23 ;
      RECT 77.57 -0.62 77.95 -0.24 ;
      RECT 66.815 -0.575 77.95 -0.27 ;
      RECT 48.88 -0.61 49.26 -0.23 ;
      RECT 59.635 -0.62 60.015 -0.24 ;
      RECT 48.88 -0.575 60.015 -0.27 ;
      RECT 30.94 -0.61 31.32 -0.23 ;
      RECT 41.695 -0.62 42.075 -0.24 ;
      RECT 30.94 -0.575 42.075 -0.27 ;
      RECT 13 -0.61 13.38 -0.23 ;
      RECT 23.755 -0.62 24.135 -0.24 ;
      RECT 13 -0.575 24.135 -0.27 ;
    LAYER via3 ;
      RECT 95.6 -0.53 95.8 -0.33 ;
      RECT 89.36 4.97 89.56 5.17 ;
      RECT 84.845 -0.52 85.045 -0.32 ;
      RECT 77.66 -0.53 77.86 -0.33 ;
      RECT 66.905 -0.52 67.105 -0.32 ;
      RECT 59.725 -0.53 59.925 -0.33 ;
      RECT 48.97 -0.52 49.17 -0.32 ;
      RECT 41.785 -0.53 41.985 -0.33 ;
      RECT 31.03 -0.52 31.23 -0.32 ;
      RECT 23.845 -0.53 24.045 -0.33 ;
      RECT 13.09 -0.52 13.29 -0.32 ;
      RECT 0.105 4.965 0.305 5.165 ;
    LAYER met3 ;
      RECT 95.51 -0.62 95.89 -0.24 ;
      RECT 95.25 -0.585 96.155 -0.275 ;
      RECT 83.1 2.31 83.47 2.68 ;
      RECT 83.1 2.345 83.775 2.645 ;
      RECT 83.43 -1.47 83.73 2.645 ;
      RECT 94.385 -0.43 94.755 -0.06 ;
      RECT 94.45 -1.435 94.75 -0.06 ;
      RECT 83.43 -1.435 94.76 -1.135 ;
      RECT 91.435 -0.385 91.765 -0.055 ;
      RECT 91.435 -0.37 92.235 -0.07 ;
      RECT 86.335 2.67 86.705 3.04 ;
      RECT 90.755 2.675 91.085 3.005 ;
      RECT 89.71 2.675 90.04 3.005 ;
      RECT 89.71 2.7 91.085 3 ;
      RECT 86.335 2.7 91.555 2.99 ;
      RECT 91.435 0.635 91.76 2.985 ;
      RECT 90.755 2.69 91.76 2.985 ;
      RECT 91.43 0.92 91.555 2.99 ;
      RECT 86.335 2.69 90.04 2.99 ;
      RECT 90.76 2.67 91.06 3.005 ;
      RECT 91.435 0.635 91.765 0.965 ;
      RECT 91.435 0.65 92.235 0.95 ;
      RECT 91.44 0.585 91.74 2.985 ;
      RECT 90.735 -0.045 91.065 0.285 ;
      RECT 90.265 -0.03 91.065 0.27 ;
      RECT 90.76 -0.06 91.06 0.285 ;
      RECT 90.075 1.655 90.405 1.985 ;
      RECT 90.075 1.67 90.875 1.97 ;
      RECT 89.245 4.855 89.665 5.28 ;
      RECT 88.93 4.9 89.96 5.245 ;
      RECT 89.395 -0.73 89.725 -0.4 ;
      RECT 88.925 -0.71 89.285 -0.41 ;
      RECT 89.285 -0.715 89.725 -0.415 ;
      RECT 89.005 3.37 89.305 3.785 ;
      RECT 89.035 3.355 89.365 3.685 ;
      RECT 88.565 3.37 89.365 3.67 ;
      RECT 84.805 2.165 85.175 2.535 ;
      RECT 84.785 -0.61 85.085 2.345 ;
      RECT 84.755 -0.61 85.135 -0.23 ;
      RECT 77.57 -0.62 77.95 -0.24 ;
      RECT 77.31 -0.585 78.215 -0.275 ;
      RECT 65.16 2.31 65.53 2.68 ;
      RECT 65.16 2.345 65.835 2.645 ;
      RECT 65.49 -1.47 65.79 2.645 ;
      RECT 76.445 -0.43 76.815 -0.06 ;
      RECT 76.51 -1.435 76.81 -0.06 ;
      RECT 65.49 -1.435 76.82 -1.135 ;
      RECT 73.495 -0.385 73.825 -0.055 ;
      RECT 73.495 -0.37 74.295 -0.07 ;
      RECT 68.395 2.67 68.765 3.04 ;
      RECT 72.815 2.675 73.145 3.005 ;
      RECT 71.77 2.675 72.1 3.005 ;
      RECT 71.77 2.7 73.145 3 ;
      RECT 68.395 2.7 73.615 2.99 ;
      RECT 73.495 0.635 73.82 2.985 ;
      RECT 72.815 2.69 73.82 2.985 ;
      RECT 73.49 0.92 73.615 2.99 ;
      RECT 68.395 2.69 72.1 2.99 ;
      RECT 72.82 2.67 73.12 3.005 ;
      RECT 73.495 0.635 73.825 0.965 ;
      RECT 73.495 0.65 74.295 0.95 ;
      RECT 73.5 0.585 73.8 2.985 ;
      RECT 72.795 -0.045 73.125 0.285 ;
      RECT 72.325 -0.03 73.125 0.27 ;
      RECT 72.82 -0.06 73.12 0.285 ;
      RECT 72.135 1.655 72.465 1.985 ;
      RECT 72.135 1.67 72.935 1.97 ;
      RECT 71.455 -0.73 71.785 -0.4 ;
      RECT 70.985 -0.71 71.345 -0.41 ;
      RECT 71.345 -0.715 71.785 -0.415 ;
      RECT 71.065 3.37 71.365 3.785 ;
      RECT 71.095 3.355 71.425 3.685 ;
      RECT 70.625 3.37 71.425 3.67 ;
      RECT 66.865 2.165 67.235 2.535 ;
      RECT 66.845 -0.61 67.145 2.345 ;
      RECT 66.815 -0.61 67.195 -0.23 ;
      RECT 59.635 -0.62 60.015 -0.24 ;
      RECT 59.375 -0.585 60.28 -0.275 ;
      RECT 47.225 2.31 47.595 2.68 ;
      RECT 47.225 2.345 47.9 2.645 ;
      RECT 47.555 -1.47 47.855 2.645 ;
      RECT 58.51 -0.43 58.88 -0.06 ;
      RECT 58.575 -1.435 58.875 -0.06 ;
      RECT 47.555 -1.435 58.885 -1.135 ;
      RECT 55.56 -0.385 55.89 -0.055 ;
      RECT 55.56 -0.37 56.36 -0.07 ;
      RECT 50.46 2.67 50.83 3.04 ;
      RECT 54.88 2.675 55.21 3.005 ;
      RECT 53.835 2.675 54.165 3.005 ;
      RECT 53.835 2.7 55.21 3 ;
      RECT 50.46 2.7 55.68 2.99 ;
      RECT 55.56 0.635 55.885 2.985 ;
      RECT 54.88 2.69 55.885 2.985 ;
      RECT 55.555 0.92 55.68 2.99 ;
      RECT 50.46 2.69 54.165 2.99 ;
      RECT 54.885 2.67 55.185 3.005 ;
      RECT 55.56 0.635 55.89 0.965 ;
      RECT 55.56 0.65 56.36 0.95 ;
      RECT 55.565 0.585 55.865 2.985 ;
      RECT 54.86 -0.045 55.19 0.285 ;
      RECT 54.39 -0.03 55.19 0.27 ;
      RECT 54.885 -0.06 55.185 0.285 ;
      RECT 54.2 1.655 54.53 1.985 ;
      RECT 54.2 1.67 55 1.97 ;
      RECT 53.52 -0.73 53.85 -0.4 ;
      RECT 53.05 -0.71 53.41 -0.41 ;
      RECT 53.41 -0.715 53.85 -0.415 ;
      RECT 53.13 3.37 53.43 3.785 ;
      RECT 53.16 3.355 53.49 3.685 ;
      RECT 52.69 3.37 53.49 3.67 ;
      RECT 48.93 2.165 49.3 2.535 ;
      RECT 48.91 -0.61 49.21 2.345 ;
      RECT 48.88 -0.61 49.26 -0.23 ;
      RECT 41.695 -0.62 42.075 -0.24 ;
      RECT 41.435 -0.585 42.34 -0.275 ;
      RECT 29.285 2.31 29.655 2.68 ;
      RECT 29.285 2.345 29.96 2.645 ;
      RECT 29.615 -1.47 29.915 2.645 ;
      RECT 40.57 -0.43 40.94 -0.06 ;
      RECT 40.635 -1.435 40.935 -0.06 ;
      RECT 29.615 -1.435 40.945 -1.135 ;
      RECT 37.62 -0.385 37.95 -0.055 ;
      RECT 37.62 -0.37 38.42 -0.07 ;
      RECT 32.52 2.67 32.89 3.04 ;
      RECT 36.94 2.675 37.27 3.005 ;
      RECT 35.895 2.675 36.225 3.005 ;
      RECT 35.895 2.7 37.27 3 ;
      RECT 32.52 2.7 37.74 2.99 ;
      RECT 37.62 0.635 37.945 2.985 ;
      RECT 36.94 2.69 37.945 2.985 ;
      RECT 37.615 0.92 37.74 2.99 ;
      RECT 32.52 2.69 36.225 2.99 ;
      RECT 36.945 2.67 37.245 3.005 ;
      RECT 37.62 0.635 37.95 0.965 ;
      RECT 37.62 0.65 38.42 0.95 ;
      RECT 37.625 0.585 37.925 2.985 ;
      RECT 36.92 -0.045 37.25 0.285 ;
      RECT 36.45 -0.03 37.25 0.27 ;
      RECT 36.945 -0.06 37.245 0.285 ;
      RECT 36.26 1.655 36.59 1.985 ;
      RECT 36.26 1.67 37.06 1.97 ;
      RECT 35.58 -0.73 35.91 -0.4 ;
      RECT 35.11 -0.71 35.47 -0.41 ;
      RECT 35.47 -0.715 35.91 -0.415 ;
      RECT 35.19 3.37 35.49 3.785 ;
      RECT 35.22 3.355 35.55 3.685 ;
      RECT 34.75 3.37 35.55 3.67 ;
      RECT 30.99 2.165 31.36 2.535 ;
      RECT 30.97 -0.61 31.27 2.345 ;
      RECT 30.94 -0.61 31.32 -0.23 ;
      RECT 23.755 -0.62 24.135 -0.24 ;
      RECT 23.495 -0.585 24.4 -0.275 ;
      RECT 11.345 2.31 11.715 2.68 ;
      RECT 11.345 2.345 12.02 2.645 ;
      RECT 11.675 -1.47 11.975 2.645 ;
      RECT 22.63 -0.43 23 -0.06 ;
      RECT 22.695 -1.435 22.995 -0.06 ;
      RECT 11.675 -1.435 23.005 -1.135 ;
      RECT 19.68 -0.385 20.01 -0.055 ;
      RECT 19.68 -0.37 20.48 -0.07 ;
      RECT 14.58 2.67 14.95 3.04 ;
      RECT 19 2.675 19.33 3.005 ;
      RECT 17.955 2.675 18.285 3.005 ;
      RECT 17.955 2.7 19.33 3 ;
      RECT 14.58 2.7 19.8 2.99 ;
      RECT 19.68 0.635 20.005 2.985 ;
      RECT 19 2.69 20.005 2.985 ;
      RECT 19.675 0.92 19.8 2.99 ;
      RECT 14.58 2.69 18.285 2.99 ;
      RECT 19.005 2.67 19.305 3.005 ;
      RECT 19.68 0.635 20.01 0.965 ;
      RECT 19.68 0.65 20.48 0.95 ;
      RECT 19.685 0.585 19.985 2.985 ;
      RECT 18.98 -0.045 19.31 0.285 ;
      RECT 18.51 -0.03 19.31 0.27 ;
      RECT 19.005 -0.06 19.305 0.285 ;
      RECT 18.32 1.655 18.65 1.985 ;
      RECT 18.32 1.67 19.12 1.97 ;
      RECT 17.64 -0.73 17.97 -0.4 ;
      RECT 17.17 -0.71 17.53 -0.41 ;
      RECT 17.53 -0.715 17.97 -0.415 ;
      RECT 17.25 3.37 17.55 3.785 ;
      RECT 17.28 3.355 17.61 3.685 ;
      RECT 16.81 3.37 17.61 3.67 ;
      RECT 13.05 2.165 13.42 2.535 ;
      RECT 13.03 -0.61 13.33 2.345 ;
      RECT 13 -0.61 13.38 -0.23 ;
      RECT -0.01 4.85 0.41 5.275 ;
      RECT -0.325 4.895 0.705 5.24 ;
    LAYER via2 ;
      RECT 95.605 -0.53 95.805 -0.33 ;
      RECT 94.47 -0.345 94.67 -0.145 ;
      RECT 91.5 -0.32 91.7 -0.12 ;
      RECT 91.5 0.7 91.7 0.9 ;
      RECT 90.82 2.74 91.02 2.94 ;
      RECT 90.8 0.02 91 0.22 ;
      RECT 90.14 1.72 90.34 1.92 ;
      RECT 89.775 2.74 89.975 2.94 ;
      RECT 89.46 -0.665 89.66 -0.465 ;
      RECT 89.36 4.97 89.56 5.17 ;
      RECT 89.1 3.42 89.3 3.62 ;
      RECT 86.42 2.755 86.62 2.955 ;
      RECT 84.89 2.25 85.09 2.45 ;
      RECT 83.185 2.395 83.385 2.595 ;
      RECT 77.665 -0.53 77.865 -0.33 ;
      RECT 76.53 -0.345 76.73 -0.145 ;
      RECT 73.56 -0.32 73.76 -0.12 ;
      RECT 73.56 0.7 73.76 0.9 ;
      RECT 72.88 2.74 73.08 2.94 ;
      RECT 72.86 0.02 73.06 0.22 ;
      RECT 72.2 1.72 72.4 1.92 ;
      RECT 71.835 2.74 72.035 2.94 ;
      RECT 71.52 -0.665 71.72 -0.465 ;
      RECT 71.16 3.42 71.36 3.62 ;
      RECT 68.48 2.755 68.68 2.955 ;
      RECT 66.95 2.25 67.15 2.45 ;
      RECT 65.245 2.395 65.445 2.595 ;
      RECT 59.73 -0.53 59.93 -0.33 ;
      RECT 58.595 -0.345 58.795 -0.145 ;
      RECT 55.625 -0.32 55.825 -0.12 ;
      RECT 55.625 0.7 55.825 0.9 ;
      RECT 54.945 2.74 55.145 2.94 ;
      RECT 54.925 0.02 55.125 0.22 ;
      RECT 54.265 1.72 54.465 1.92 ;
      RECT 53.9 2.74 54.1 2.94 ;
      RECT 53.585 -0.665 53.785 -0.465 ;
      RECT 53.225 3.42 53.425 3.62 ;
      RECT 50.545 2.755 50.745 2.955 ;
      RECT 49.015 2.25 49.215 2.45 ;
      RECT 47.31 2.395 47.51 2.595 ;
      RECT 41.79 -0.53 41.99 -0.33 ;
      RECT 40.655 -0.345 40.855 -0.145 ;
      RECT 37.685 -0.32 37.885 -0.12 ;
      RECT 37.685 0.7 37.885 0.9 ;
      RECT 37.005 2.74 37.205 2.94 ;
      RECT 36.985 0.02 37.185 0.22 ;
      RECT 36.325 1.72 36.525 1.92 ;
      RECT 35.96 2.74 36.16 2.94 ;
      RECT 35.645 -0.665 35.845 -0.465 ;
      RECT 35.285 3.42 35.485 3.62 ;
      RECT 32.605 2.755 32.805 2.955 ;
      RECT 31.075 2.25 31.275 2.45 ;
      RECT 29.37 2.395 29.57 2.595 ;
      RECT 23.85 -0.53 24.05 -0.33 ;
      RECT 22.715 -0.345 22.915 -0.145 ;
      RECT 19.745 -0.32 19.945 -0.12 ;
      RECT 19.745 0.7 19.945 0.9 ;
      RECT 19.065 2.74 19.265 2.94 ;
      RECT 19.045 0.02 19.245 0.22 ;
      RECT 18.385 1.72 18.585 1.92 ;
      RECT 18.02 2.74 18.22 2.94 ;
      RECT 17.705 -0.665 17.905 -0.465 ;
      RECT 17.345 3.42 17.545 3.62 ;
      RECT 14.665 2.755 14.865 2.955 ;
      RECT 13.135 2.25 13.335 2.45 ;
      RECT 11.43 2.395 11.63 2.595 ;
      RECT 0.105 4.965 0.305 5.165 ;
    LAYER met2 ;
      RECT 95.52 2.865 95.86 3.205 ;
      RECT 95.52 2.995 96.795 3.185 ;
      RECT 96.605 1.76 96.795 3.185 ;
      RECT 96.135 1.76 96.795 1.95 ;
      RECT 96.135 -0.01 96.325 1.95 ;
      RECT 95.985 -0.01 96.325 0.33 ;
      RECT 92.525 -0.01 92.865 0.33 ;
      RECT 92.815 -1.04 92.955 0.285 ;
      RECT 96.18 -1.04 96.32 1.95 ;
      RECT 92.815 -1.04 96.32 -0.9 ;
      RECT 95.94 2.26 96.28 2.6 ;
      RECT 95.165 2.26 96.28 2.43 ;
      RECT 95.165 -0.51 95.335 2.43 ;
      RECT 95.52 -0.615 95.89 -0.245 ;
      RECT 95.165 -0.51 95.89 -0.34 ;
      RECT 94.385 2.705 94.725 3.045 ;
      RECT 94.495 -0.43 94.665 3.045 ;
      RECT 94.385 -0.43 94.755 -0.06 ;
      RECT 93.16 1.66 93.42 1.98 ;
      RECT 93.22 -0.38 93.36 1.98 ;
      RECT 93.16 -0.38 93.42 -0.06 ;
      RECT 92.14 2.68 92.4 3 ;
      RECT 91.52 2.77 92.4 2.91 ;
      RECT 91.52 0.615 91.66 2.91 ;
      RECT 91.46 0.615 91.74 0.985 ;
      RECT 90.78 2.655 91.06 3.025 ;
      RECT 90.84 0.73 90.98 3.025 ;
      RECT 90.84 0.73 91.32 0.87 ;
      RECT 91.18 -1.06 91.32 0.87 ;
      RECT 91.12 -1.06 91.38 -0.74 ;
      RECT 90.1 1.635 90.38 2.005 ;
      RECT 90.16 -0.72 90.3 2.005 ;
      RECT 90.1 -0.72 90.36 -0.4 ;
      RECT 89.735 2.655 90.015 3.025 ;
      RECT 89.735 2.68 90.02 3 ;
      RECT 77.58 2.865 77.92 3.205 ;
      RECT 77.58 2.995 78.855 3.185 ;
      RECT 78.665 1.76 78.855 3.185 ;
      RECT 78.195 1.76 78.855 1.95 ;
      RECT 78.195 -0.01 78.385 1.95 ;
      RECT 78.045 -0.01 78.385 0.33 ;
      RECT 74.585 -0.01 74.925 0.33 ;
      RECT 74.875 -1.04 75.015 0.285 ;
      RECT 78.24 -1.04 78.38 1.95 ;
      RECT 74.875 -1.04 78.38 -0.9 ;
      RECT 78 2.26 78.34 2.6 ;
      RECT 77.225 2.26 78.34 2.43 ;
      RECT 77.225 -0.51 77.395 2.43 ;
      RECT 77.58 -0.615 77.95 -0.245 ;
      RECT 77.225 -0.51 77.95 -0.34 ;
      RECT 76.445 2.705 76.785 3.045 ;
      RECT 76.555 -0.43 76.725 3.045 ;
      RECT 76.445 -0.43 76.815 -0.06 ;
      RECT 75.22 1.66 75.48 1.98 ;
      RECT 75.28 -0.38 75.42 1.98 ;
      RECT 75.22 -0.38 75.48 -0.06 ;
      RECT 74.2 2.68 74.46 3 ;
      RECT 73.58 2.77 74.46 2.91 ;
      RECT 73.58 0.615 73.72 2.91 ;
      RECT 73.52 0.615 73.8 0.985 ;
      RECT 72.84 2.655 73.12 3.025 ;
      RECT 72.9 0.73 73.04 3.025 ;
      RECT 72.9 0.73 73.38 0.87 ;
      RECT 73.24 -1.06 73.38 0.87 ;
      RECT 73.18 -1.06 73.44 -0.74 ;
      RECT 72.16 1.635 72.44 2.005 ;
      RECT 72.22 -0.72 72.36 2.005 ;
      RECT 72.16 -0.72 72.42 -0.4 ;
      RECT 71.795 2.655 72.075 3.025 ;
      RECT 71.795 2.68 72.08 3 ;
      RECT 59.645 2.865 59.985 3.205 ;
      RECT 59.645 2.995 60.92 3.185 ;
      RECT 60.73 1.76 60.92 3.185 ;
      RECT 60.26 1.76 60.92 1.95 ;
      RECT 60.26 -0.01 60.45 1.95 ;
      RECT 60.11 -0.01 60.45 0.33 ;
      RECT 56.65 -0.01 56.99 0.33 ;
      RECT 56.94 -1.04 57.08 0.285 ;
      RECT 60.305 -1.04 60.445 1.95 ;
      RECT 56.94 -1.04 60.445 -0.9 ;
      RECT 60.065 2.26 60.405 2.6 ;
      RECT 59.29 2.26 60.405 2.43 ;
      RECT 59.29 -0.51 59.46 2.43 ;
      RECT 59.645 -0.615 60.015 -0.245 ;
      RECT 59.29 -0.51 60.015 -0.34 ;
      RECT 58.51 2.705 58.85 3.045 ;
      RECT 58.62 -0.43 58.79 3.045 ;
      RECT 58.51 -0.43 58.88 -0.06 ;
      RECT 57.285 1.66 57.545 1.98 ;
      RECT 57.345 -0.38 57.485 1.98 ;
      RECT 57.285 -0.38 57.545 -0.06 ;
      RECT 56.265 2.68 56.525 3 ;
      RECT 55.645 2.77 56.525 2.91 ;
      RECT 55.645 0.615 55.785 2.91 ;
      RECT 55.585 0.615 55.865 0.985 ;
      RECT 54.905 2.655 55.185 3.025 ;
      RECT 54.965 0.73 55.105 3.025 ;
      RECT 54.965 0.73 55.445 0.87 ;
      RECT 55.305 -1.06 55.445 0.87 ;
      RECT 55.245 -1.06 55.505 -0.74 ;
      RECT 54.225 1.635 54.505 2.005 ;
      RECT 54.285 -0.72 54.425 2.005 ;
      RECT 54.225 -0.72 54.485 -0.4 ;
      RECT 53.86 2.655 54.14 3.025 ;
      RECT 53.86 2.68 54.145 3 ;
      RECT 41.705 2.865 42.045 3.205 ;
      RECT 41.705 2.995 42.98 3.185 ;
      RECT 42.79 1.76 42.98 3.185 ;
      RECT 42.32 1.76 42.98 1.95 ;
      RECT 42.32 -0.01 42.51 1.95 ;
      RECT 42.17 -0.01 42.51 0.33 ;
      RECT 38.71 -0.01 39.05 0.33 ;
      RECT 39 -1.04 39.14 0.285 ;
      RECT 42.365 -1.04 42.505 1.95 ;
      RECT 39 -1.04 42.505 -0.9 ;
      RECT 42.125 2.26 42.465 2.6 ;
      RECT 41.35 2.26 42.465 2.43 ;
      RECT 41.35 -0.51 41.52 2.43 ;
      RECT 41.705 -0.615 42.075 -0.245 ;
      RECT 41.35 -0.51 42.075 -0.34 ;
      RECT 40.57 2.705 40.91 3.045 ;
      RECT 40.68 -0.43 40.85 3.045 ;
      RECT 40.57 -0.43 40.94 -0.06 ;
      RECT 39.345 1.66 39.605 1.98 ;
      RECT 39.405 -0.38 39.545 1.98 ;
      RECT 39.345 -0.38 39.605 -0.06 ;
      RECT 38.325 2.68 38.585 3 ;
      RECT 37.705 2.77 38.585 2.91 ;
      RECT 37.705 0.615 37.845 2.91 ;
      RECT 37.645 0.615 37.925 0.985 ;
      RECT 36.965 2.655 37.245 3.025 ;
      RECT 37.025 0.73 37.165 3.025 ;
      RECT 37.025 0.73 37.505 0.87 ;
      RECT 37.365 -1.06 37.505 0.87 ;
      RECT 37.305 -1.06 37.565 -0.74 ;
      RECT 36.285 1.635 36.565 2.005 ;
      RECT 36.345 -0.72 36.485 2.005 ;
      RECT 36.285 -0.72 36.545 -0.4 ;
      RECT 35.92 2.655 36.2 3.025 ;
      RECT 35.92 2.68 36.205 3 ;
      RECT 23.765 2.865 24.105 3.205 ;
      RECT 23.765 2.995 25.04 3.185 ;
      RECT 24.85 1.76 25.04 3.185 ;
      RECT 24.38 1.76 25.04 1.95 ;
      RECT 24.38 -0.01 24.57 1.95 ;
      RECT 24.23 -0.01 24.57 0.33 ;
      RECT 20.77 -0.01 21.11 0.33 ;
      RECT 21.06 -1.04 21.2 0.285 ;
      RECT 24.425 -1.04 24.565 1.95 ;
      RECT 21.06 -1.04 24.565 -0.9 ;
      RECT 24.185 2.26 24.525 2.6 ;
      RECT 23.41 2.26 24.525 2.43 ;
      RECT 23.41 -0.51 23.58 2.43 ;
      RECT 23.765 -0.615 24.135 -0.245 ;
      RECT 23.41 -0.51 24.135 -0.34 ;
      RECT 22.63 2.705 22.97 3.045 ;
      RECT 22.74 -0.43 22.91 3.045 ;
      RECT 22.63 -0.43 23 -0.06 ;
      RECT 21.405 1.66 21.665 1.98 ;
      RECT 21.465 -0.38 21.605 1.98 ;
      RECT 21.405 -0.38 21.665 -0.06 ;
      RECT 20.385 2.68 20.645 3 ;
      RECT 19.765 2.77 20.645 2.91 ;
      RECT 19.765 0.615 19.905 2.91 ;
      RECT 19.705 0.615 19.985 0.985 ;
      RECT 19.025 2.655 19.305 3.025 ;
      RECT 19.085 0.73 19.225 3.025 ;
      RECT 19.085 0.73 19.565 0.87 ;
      RECT 19.425 -1.06 19.565 0.87 ;
      RECT 19.365 -1.06 19.625 -0.74 ;
      RECT 18.345 1.635 18.625 2.005 ;
      RECT 18.405 -0.72 18.545 2.005 ;
      RECT 18.345 -0.72 18.605 -0.4 ;
      RECT 17.98 2.655 18.26 3.025 ;
      RECT 17.98 2.68 18.265 3 ;
      RECT 2.52 3.55 2.645 3.985 ;
      RECT 2.52 3.55 2.66 3.93 ;
      RECT -3.885 3.55 -3.505 3.93 ;
      RECT -3.885 3.55 2.66 3.69 ;
      RECT 91.46 -0.405 91.74 -0.035 ;
      RECT 90.76 -0.065 91.04 0.305 ;
      RECT 89.42 -0.75 89.7 -0.38 ;
      RECT 89.24 4.86 89.67 5.28 ;
      RECT 89.06 3.335 89.34 3.705 ;
      RECT 86.335 2.67 86.705 3.04 ;
      RECT 84.805 2.165 85.175 2.535 ;
      RECT 83.1 2.31 83.47 2.68 ;
      RECT 73.52 -0.405 73.8 -0.035 ;
      RECT 72.82 -0.065 73.1 0.305 ;
      RECT 71.48 -0.75 71.76 -0.38 ;
      RECT 71.12 3.335 71.4 3.705 ;
      RECT 68.395 2.67 68.765 3.04 ;
      RECT 66.865 2.165 67.235 2.535 ;
      RECT 65.16 2.31 65.53 2.68 ;
      RECT 55.585 -0.405 55.865 -0.035 ;
      RECT 54.885 -0.065 55.165 0.305 ;
      RECT 53.545 -0.75 53.825 -0.38 ;
      RECT 53.185 3.335 53.465 3.705 ;
      RECT 50.46 2.67 50.83 3.04 ;
      RECT 48.93 2.165 49.3 2.535 ;
      RECT 47.225 2.31 47.595 2.68 ;
      RECT 37.645 -0.405 37.925 -0.035 ;
      RECT 36.945 -0.065 37.225 0.305 ;
      RECT 35.605 -0.75 35.885 -0.38 ;
      RECT 35.245 3.335 35.525 3.705 ;
      RECT 32.52 2.67 32.89 3.04 ;
      RECT 30.99 2.165 31.36 2.535 ;
      RECT 29.285 2.31 29.655 2.68 ;
      RECT 19.705 -0.405 19.985 -0.035 ;
      RECT 19.005 -0.065 19.285 0.305 ;
      RECT 17.665 -0.75 17.945 -0.38 ;
      RECT 17.305 3.335 17.585 3.705 ;
      RECT 14.58 2.67 14.95 3.04 ;
      RECT 13.05 2.165 13.42 2.535 ;
      RECT 11.345 2.31 11.715 2.68 ;
      RECT -0.015 4.855 0.415 5.275 ;
    LAYER via1 ;
      RECT 96.08 0.085 96.23 0.235 ;
      RECT 96.035 2.355 96.185 2.505 ;
      RECT 95.63 -0.505 95.78 -0.355 ;
      RECT 95.615 2.96 95.765 3.11 ;
      RECT 94.485 -0.33 94.635 -0.18 ;
      RECT 94.48 2.8 94.63 2.95 ;
      RECT 93.215 -0.295 93.365 -0.145 ;
      RECT 93.215 1.745 93.365 1.895 ;
      RECT 92.62 0.085 92.77 0.235 ;
      RECT 92.195 2.765 92.345 2.915 ;
      RECT 91.515 -0.295 91.665 -0.145 ;
      RECT 91.515 0.725 91.665 0.875 ;
      RECT 91.175 -0.975 91.325 -0.825 ;
      RECT 90.835 0.045 90.985 0.195 ;
      RECT 90.835 2.765 90.985 2.915 ;
      RECT 90.155 -0.635 90.305 -0.485 ;
      RECT 90.155 1.745 90.305 1.895 ;
      RECT 89.815 2.765 89.965 2.915 ;
      RECT 89.475 -0.64 89.625 -0.49 ;
      RECT 89.385 4.995 89.535 5.145 ;
      RECT 89.135 3.445 89.285 3.595 ;
      RECT 86.445 2.78 86.595 2.93 ;
      RECT 84.915 2.275 85.065 2.425 ;
      RECT 83.21 2.42 83.36 2.57 ;
      RECT 78.14 0.085 78.29 0.235 ;
      RECT 78.095 2.355 78.245 2.505 ;
      RECT 77.69 -0.505 77.84 -0.355 ;
      RECT 77.675 2.96 77.825 3.11 ;
      RECT 76.545 -0.33 76.695 -0.18 ;
      RECT 76.54 2.8 76.69 2.95 ;
      RECT 75.275 -0.295 75.425 -0.145 ;
      RECT 75.275 1.745 75.425 1.895 ;
      RECT 74.68 0.085 74.83 0.235 ;
      RECT 74.255 2.765 74.405 2.915 ;
      RECT 73.575 -0.295 73.725 -0.145 ;
      RECT 73.575 0.725 73.725 0.875 ;
      RECT 73.235 -0.975 73.385 -0.825 ;
      RECT 72.895 0.045 73.045 0.195 ;
      RECT 72.895 2.765 73.045 2.915 ;
      RECT 72.215 -0.635 72.365 -0.485 ;
      RECT 72.215 1.745 72.365 1.895 ;
      RECT 71.875 2.765 72.025 2.915 ;
      RECT 71.535 -0.64 71.685 -0.49 ;
      RECT 71.195 3.445 71.345 3.595 ;
      RECT 68.505 2.78 68.655 2.93 ;
      RECT 66.975 2.275 67.125 2.425 ;
      RECT 65.27 2.42 65.42 2.57 ;
      RECT 60.205 0.085 60.355 0.235 ;
      RECT 60.16 2.355 60.31 2.505 ;
      RECT 59.755 -0.505 59.905 -0.355 ;
      RECT 59.74 2.96 59.89 3.11 ;
      RECT 58.61 -0.33 58.76 -0.18 ;
      RECT 58.605 2.8 58.755 2.95 ;
      RECT 57.34 -0.295 57.49 -0.145 ;
      RECT 57.34 1.745 57.49 1.895 ;
      RECT 56.745 0.085 56.895 0.235 ;
      RECT 56.32 2.765 56.47 2.915 ;
      RECT 55.64 -0.295 55.79 -0.145 ;
      RECT 55.64 0.725 55.79 0.875 ;
      RECT 55.3 -0.975 55.45 -0.825 ;
      RECT 54.96 0.045 55.11 0.195 ;
      RECT 54.96 2.765 55.11 2.915 ;
      RECT 54.28 -0.635 54.43 -0.485 ;
      RECT 54.28 1.745 54.43 1.895 ;
      RECT 53.94 2.765 54.09 2.915 ;
      RECT 53.6 -0.64 53.75 -0.49 ;
      RECT 53.26 3.445 53.41 3.595 ;
      RECT 50.57 2.78 50.72 2.93 ;
      RECT 49.04 2.275 49.19 2.425 ;
      RECT 47.335 2.42 47.485 2.57 ;
      RECT 42.265 0.085 42.415 0.235 ;
      RECT 42.22 2.355 42.37 2.505 ;
      RECT 41.815 -0.505 41.965 -0.355 ;
      RECT 41.8 2.96 41.95 3.11 ;
      RECT 40.67 -0.33 40.82 -0.18 ;
      RECT 40.665 2.8 40.815 2.95 ;
      RECT 39.4 -0.295 39.55 -0.145 ;
      RECT 39.4 1.745 39.55 1.895 ;
      RECT 38.805 0.085 38.955 0.235 ;
      RECT 38.38 2.765 38.53 2.915 ;
      RECT 37.7 -0.295 37.85 -0.145 ;
      RECT 37.7 0.725 37.85 0.875 ;
      RECT 37.36 -0.975 37.51 -0.825 ;
      RECT 37.02 0.045 37.17 0.195 ;
      RECT 37.02 2.765 37.17 2.915 ;
      RECT 36.34 -0.635 36.49 -0.485 ;
      RECT 36.34 1.745 36.49 1.895 ;
      RECT 36 2.765 36.15 2.915 ;
      RECT 35.66 -0.64 35.81 -0.49 ;
      RECT 35.32 3.445 35.47 3.595 ;
      RECT 32.63 2.78 32.78 2.93 ;
      RECT 31.1 2.275 31.25 2.425 ;
      RECT 29.395 2.42 29.545 2.57 ;
      RECT 24.325 0.085 24.475 0.235 ;
      RECT 24.28 2.355 24.43 2.505 ;
      RECT 23.875 -0.505 24.025 -0.355 ;
      RECT 23.86 2.96 24.01 3.11 ;
      RECT 22.73 -0.33 22.88 -0.18 ;
      RECT 22.725 2.8 22.875 2.95 ;
      RECT 21.46 -0.295 21.61 -0.145 ;
      RECT 21.46 1.745 21.61 1.895 ;
      RECT 20.865 0.085 21.015 0.235 ;
      RECT 20.44 2.765 20.59 2.915 ;
      RECT 19.76 -0.295 19.91 -0.145 ;
      RECT 19.76 0.725 19.91 0.875 ;
      RECT 19.42 -0.975 19.57 -0.825 ;
      RECT 19.08 0.045 19.23 0.195 ;
      RECT 19.08 2.765 19.23 2.915 ;
      RECT 18.4 -0.635 18.55 -0.485 ;
      RECT 18.4 1.745 18.55 1.895 ;
      RECT 18.06 2.765 18.21 2.915 ;
      RECT 17.72 -0.64 17.87 -0.49 ;
      RECT 17.38 3.445 17.53 3.595 ;
      RECT 14.69 2.78 14.84 2.93 ;
      RECT 13.16 2.275 13.31 2.425 ;
      RECT 11.455 2.42 11.605 2.57 ;
      RECT 0.13 4.99 0.28 5.14 ;
      RECT -3.77 3.665 -3.62 3.815 ;
    LAYER met1 ;
      RECT 10.765 3.79 100.46 4.27 ;
      RECT 89.09 3.39 89.335 4.27 ;
      RECT 71.15 3.655 74.4 4.27 ;
      RECT 53.215 3.655 56.5 4.27 ;
      RECT 35.275 3.655 38.52 4.27 ;
      RECT 17.335 3.655 20.685 4.27 ;
      RECT 71.15 3.625 71.565 4.27 ;
      RECT 53.215 3.625 53.63 4.27 ;
      RECT 35.275 3.625 35.69 4.27 ;
      RECT 17.335 3.61 17.765 4.27 ;
      RECT 89.05 3.39 89.37 3.65 ;
      RECT 71.11 3.39 71.43 3.65 ;
      RECT 53.175 3.39 53.495 3.65 ;
      RECT 35.235 3.39 35.555 3.65 ;
      RECT 17.295 3.39 17.615 3.65 ;
      RECT 88.12 3.45 90.47 3.59 ;
      RECT 90.33 2.725 90.47 3.59 ;
      RECT 70.18 3.45 72.53 3.59 ;
      RECT 72.39 2.725 72.53 3.59 ;
      RECT 52.245 3.45 54.595 3.59 ;
      RECT 54.455 2.725 54.595 3.59 ;
      RECT 34.305 3.45 36.655 3.59 ;
      RECT 36.515 2.725 36.655 3.59 ;
      RECT 16.365 3.45 18.715 3.59 ;
      RECT 18.575 2.725 18.715 3.59 ;
      RECT 88.12 2.725 88.26 3.59 ;
      RECT 70.18 2.725 70.32 3.59 ;
      RECT 52.245 2.725 52.385 3.59 ;
      RECT 34.305 2.725 34.445 3.59 ;
      RECT 16.365 2.725 16.505 3.59 ;
      RECT 90.255 2.725 90.545 2.955 ;
      RECT 88.045 2.725 88.335 2.955 ;
      RECT 72.315 2.725 72.605 2.955 ;
      RECT 70.105 2.725 70.395 2.955 ;
      RECT 54.38 2.725 54.67 2.955 ;
      RECT 52.17 2.725 52.46 2.955 ;
      RECT 36.44 2.725 36.73 2.955 ;
      RECT 34.23 2.725 34.52 2.955 ;
      RECT 18.5 2.725 18.79 2.955 ;
      RECT 16.29 2.725 16.58 2.955 ;
      RECT 93.815 3.475 98.265 3.64 ;
      RECT 98.1 2.725 98.265 3.64 ;
      RECT 93.735 3.26 93.905 3.525 ;
      RECT 93.675 3.28 93.955 3.525 ;
      RECT 98.1 2.725 98.27 3.015 ;
      RECT 98.065 2.755 98.315 2.99 ;
      RECT 98.08 -1.01 98.25 -0.105 ;
      RECT 98.05 -0.365 98.28 -0.13 ;
      RECT 93.64 -0.89 93.9 -0.66 ;
      RECT 93.64 -0.86 94.975 -0.69 ;
      RECT 94.805 -1.01 98.25 -0.84 ;
      RECT 93.13 -0.35 93.45 -0.09 ;
      RECT 92.855 -0.29 93.45 -0.15 ;
      RECT 92.525 -0.01 92.865 0.33 ;
      RECT 90.75 -0.01 91.07 0.25 ;
      RECT 92.525 0.005 93.015 0.235 ;
      RECT 90.75 0.05 93.015 0.19 ;
      RECT 92.11 2.71 92.43 2.97 ;
      RECT 92.11 2.77 92.705 2.91 ;
      RECT 91.43 -0.35 91.75 -0.09 ;
      RECT 86.69 -0.335 86.98 -0.105 ;
      RECT 86.69 -0.29 91.75 -0.15 ;
      RECT 91.52 -0.63 91.66 -0.09 ;
      RECT 91.52 -0.63 92 -0.49 ;
      RECT 91.86 -1.015 92 -0.49 ;
      RECT 91.785 -1.015 92.075 -0.785 ;
      RECT 91.43 0.67 91.75 0.93 ;
      RECT 90.765 0.685 91.055 0.915 ;
      RECT 88.555 0.685 88.845 0.915 ;
      RECT 88.555 0.73 91.75 0.87 ;
      RECT 89.73 2.71 90.05 2.97 ;
      RECT 91.445 2.725 91.735 2.955 ;
      RECT 89.065 2.725 89.355 2.955 ;
      RECT 89.065 2.77 90.05 2.91 ;
      RECT 91.52 2.43 91.66 2.955 ;
      RECT 89.82 2.43 89.96 2.97 ;
      RECT 89.82 2.43 91.66 2.57 ;
      RECT 88.725 -0.675 89.015 -0.445 ;
      RECT 88.8 -0.97 88.94 -0.445 ;
      RECT 91.09 -1.03 91.41 -0.77 ;
      RECT 90.99 -1.015 91.41 -0.785 ;
      RECT 88.8 -0.97 91.41 -0.83 ;
      RECT 90.07 -0.69 90.39 -0.43 ;
      RECT 90.07 -0.63 90.665 -0.49 ;
      RECT 90.07 1.69 90.39 1.95 ;
      RECT 87.365 1.705 87.655 1.935 ;
      RECT 87.365 1.75 90.39 1.89 ;
      RECT 89.395 -0.73 89.725 -0.4 ;
      RECT 89.39 -0.695 89.725 -0.435 ;
      RECT 89.74 -0.675 89.855 -0.445 ;
      RECT 89.39 -0.68 89.74 -0.45 ;
      RECT 89.39 -0.63 89.87 -0.49 ;
      RECT 89.275 -0.63 89.285 -0.49 ;
      RECT 89.285 -0.635 89.855 -0.495 ;
      RECT 75.875 3.475 80.325 3.64 ;
      RECT 80.16 2.725 80.325 3.64 ;
      RECT 75.795 3.26 75.965 3.525 ;
      RECT 75.735 3.28 76.015 3.525 ;
      RECT 80.16 2.725 80.33 3.015 ;
      RECT 80.125 2.755 80.375 2.99 ;
      RECT 80.14 -1.01 80.31 -0.105 ;
      RECT 80.11 -0.365 80.34 -0.13 ;
      RECT 75.7 -0.89 75.96 -0.66 ;
      RECT 75.7 -0.86 77.035 -0.69 ;
      RECT 76.865 -1.01 80.31 -0.84 ;
      RECT 75.19 -0.35 75.51 -0.09 ;
      RECT 74.915 -0.29 75.51 -0.15 ;
      RECT 74.585 -0.01 74.925 0.33 ;
      RECT 72.81 -0.01 73.13 0.25 ;
      RECT 74.585 0.005 75.075 0.235 ;
      RECT 72.81 0.05 75.075 0.19 ;
      RECT 74.17 2.71 74.49 2.97 ;
      RECT 74.17 2.77 74.765 2.91 ;
      RECT 73.49 -0.35 73.81 -0.09 ;
      RECT 68.75 -0.335 69.04 -0.105 ;
      RECT 68.75 -0.29 73.81 -0.15 ;
      RECT 73.58 -0.63 73.72 -0.09 ;
      RECT 73.58 -0.63 74.06 -0.49 ;
      RECT 73.92 -1.015 74.06 -0.49 ;
      RECT 73.845 -1.015 74.135 -0.785 ;
      RECT 73.49 0.67 73.81 0.93 ;
      RECT 72.825 0.685 73.115 0.915 ;
      RECT 70.615 0.685 70.905 0.915 ;
      RECT 70.615 0.73 73.81 0.87 ;
      RECT 71.79 2.71 72.11 2.97 ;
      RECT 73.505 2.725 73.795 2.955 ;
      RECT 71.125 2.725 71.415 2.955 ;
      RECT 71.125 2.77 72.11 2.91 ;
      RECT 73.58 2.43 73.72 2.955 ;
      RECT 71.88 2.43 72.02 2.97 ;
      RECT 71.88 2.43 73.72 2.57 ;
      RECT 70.785 -0.675 71.075 -0.445 ;
      RECT 70.86 -0.97 71 -0.445 ;
      RECT 73.15 -1.03 73.47 -0.77 ;
      RECT 73.05 -1.015 73.47 -0.785 ;
      RECT 70.86 -0.97 73.47 -0.83 ;
      RECT 72.13 -0.69 72.45 -0.43 ;
      RECT 72.13 -0.63 72.725 -0.49 ;
      RECT 72.13 1.69 72.45 1.95 ;
      RECT 69.425 1.705 69.715 1.935 ;
      RECT 69.425 1.75 72.45 1.89 ;
      RECT 71.455 -0.73 71.785 -0.4 ;
      RECT 71.45 -0.695 71.785 -0.435 ;
      RECT 71.8 -0.675 71.915 -0.445 ;
      RECT 71.45 -0.68 71.8 -0.45 ;
      RECT 71.45 -0.63 71.93 -0.49 ;
      RECT 71.335 -0.63 71.345 -0.49 ;
      RECT 71.345 -0.635 71.915 -0.495 ;
      RECT 57.94 3.475 62.39 3.64 ;
      RECT 62.225 2.725 62.39 3.64 ;
      RECT 57.86 3.26 58.03 3.525 ;
      RECT 57.8 3.28 58.08 3.525 ;
      RECT 62.225 2.725 62.395 3.015 ;
      RECT 62.19 2.755 62.44 2.99 ;
      RECT 62.205 -1.01 62.375 -0.105 ;
      RECT 62.175 -0.365 62.405 -0.13 ;
      RECT 57.765 -0.89 58.025 -0.66 ;
      RECT 57.765 -0.86 59.1 -0.69 ;
      RECT 58.93 -1.01 62.375 -0.84 ;
      RECT 57.255 -0.35 57.575 -0.09 ;
      RECT 56.98 -0.29 57.575 -0.15 ;
      RECT 56.65 -0.01 56.99 0.33 ;
      RECT 54.875 -0.01 55.195 0.25 ;
      RECT 56.65 0.005 57.14 0.235 ;
      RECT 54.875 0.05 57.14 0.19 ;
      RECT 56.235 2.71 56.555 2.97 ;
      RECT 56.235 2.77 56.83 2.91 ;
      RECT 55.555 -0.35 55.875 -0.09 ;
      RECT 50.815 -0.335 51.105 -0.105 ;
      RECT 50.815 -0.29 55.875 -0.15 ;
      RECT 55.645 -0.63 55.785 -0.09 ;
      RECT 55.645 -0.63 56.125 -0.49 ;
      RECT 55.985 -1.015 56.125 -0.49 ;
      RECT 55.91 -1.015 56.2 -0.785 ;
      RECT 55.555 0.67 55.875 0.93 ;
      RECT 54.89 0.685 55.18 0.915 ;
      RECT 52.68 0.685 52.97 0.915 ;
      RECT 52.68 0.73 55.875 0.87 ;
      RECT 53.855 2.71 54.175 2.97 ;
      RECT 55.57 2.725 55.86 2.955 ;
      RECT 53.19 2.725 53.48 2.955 ;
      RECT 53.19 2.77 54.175 2.91 ;
      RECT 55.645 2.43 55.785 2.955 ;
      RECT 53.945 2.43 54.085 2.97 ;
      RECT 53.945 2.43 55.785 2.57 ;
      RECT 52.85 -0.675 53.14 -0.445 ;
      RECT 52.925 -0.97 53.065 -0.445 ;
      RECT 55.215 -1.03 55.535 -0.77 ;
      RECT 55.115 -1.015 55.535 -0.785 ;
      RECT 52.925 -0.97 55.535 -0.83 ;
      RECT 54.195 -0.69 54.515 -0.43 ;
      RECT 54.195 -0.63 54.79 -0.49 ;
      RECT 54.195 1.69 54.515 1.95 ;
      RECT 51.49 1.705 51.78 1.935 ;
      RECT 51.49 1.75 54.515 1.89 ;
      RECT 53.52 -0.73 53.85 -0.4 ;
      RECT 53.515 -0.695 53.85 -0.435 ;
      RECT 53.865 -0.675 53.98 -0.445 ;
      RECT 53.515 -0.68 53.865 -0.45 ;
      RECT 53.515 -0.63 53.995 -0.49 ;
      RECT 53.4 -0.63 53.41 -0.49 ;
      RECT 53.41 -0.635 53.98 -0.495 ;
      RECT 40 3.475 44.45 3.64 ;
      RECT 44.285 2.725 44.45 3.64 ;
      RECT 39.92 3.26 40.09 3.525 ;
      RECT 39.86 3.28 40.14 3.525 ;
      RECT 44.285 2.725 44.455 3.015 ;
      RECT 44.25 2.755 44.5 2.99 ;
      RECT 44.265 -1.01 44.435 -0.105 ;
      RECT 44.235 -0.365 44.465 -0.13 ;
      RECT 39.825 -0.89 40.085 -0.66 ;
      RECT 39.825 -0.86 41.16 -0.69 ;
      RECT 40.99 -1.01 44.435 -0.84 ;
      RECT 39.315 -0.35 39.635 -0.09 ;
      RECT 39.04 -0.29 39.635 -0.15 ;
      RECT 38.71 -0.01 39.05 0.33 ;
      RECT 36.935 -0.01 37.255 0.25 ;
      RECT 38.71 0.005 39.2 0.235 ;
      RECT 36.935 0.05 39.2 0.19 ;
      RECT 38.295 2.71 38.615 2.97 ;
      RECT 38.295 2.77 38.89 2.91 ;
      RECT 37.615 -0.35 37.935 -0.09 ;
      RECT 32.875 -0.335 33.165 -0.105 ;
      RECT 32.875 -0.29 37.935 -0.15 ;
      RECT 37.705 -0.63 37.845 -0.09 ;
      RECT 37.705 -0.63 38.185 -0.49 ;
      RECT 38.045 -1.015 38.185 -0.49 ;
      RECT 37.97 -1.015 38.26 -0.785 ;
      RECT 37.615 0.67 37.935 0.93 ;
      RECT 36.95 0.685 37.24 0.915 ;
      RECT 34.74 0.685 35.03 0.915 ;
      RECT 34.74 0.73 37.935 0.87 ;
      RECT 35.915 2.71 36.235 2.97 ;
      RECT 37.63 2.725 37.92 2.955 ;
      RECT 35.25 2.725 35.54 2.955 ;
      RECT 35.25 2.77 36.235 2.91 ;
      RECT 37.705 2.43 37.845 2.955 ;
      RECT 36.005 2.43 36.145 2.97 ;
      RECT 36.005 2.43 37.845 2.57 ;
      RECT 34.91 -0.675 35.2 -0.445 ;
      RECT 34.985 -0.97 35.125 -0.445 ;
      RECT 37.275 -1.03 37.595 -0.77 ;
      RECT 37.175 -1.015 37.595 -0.785 ;
      RECT 34.985 -0.97 37.595 -0.83 ;
      RECT 36.255 -0.69 36.575 -0.43 ;
      RECT 36.255 -0.63 36.85 -0.49 ;
      RECT 36.255 1.69 36.575 1.95 ;
      RECT 33.55 1.705 33.84 1.935 ;
      RECT 33.55 1.75 36.575 1.89 ;
      RECT 35.58 -0.73 35.91 -0.4 ;
      RECT 35.575 -0.695 35.91 -0.435 ;
      RECT 35.925 -0.675 36.04 -0.445 ;
      RECT 35.575 -0.68 35.925 -0.45 ;
      RECT 35.575 -0.63 36.055 -0.49 ;
      RECT 35.46 -0.63 35.47 -0.49 ;
      RECT 35.47 -0.635 36.04 -0.495 ;
      RECT 22.06 3.475 26.51 3.64 ;
      RECT 26.345 2.725 26.51 3.64 ;
      RECT 21.98 3.26 22.15 3.525 ;
      RECT 21.92 3.28 22.2 3.525 ;
      RECT 26.345 2.725 26.515 3.015 ;
      RECT 26.31 2.755 26.56 2.99 ;
      RECT 26.325 -1.01 26.495 -0.105 ;
      RECT 26.295 -0.365 26.525 -0.13 ;
      RECT 21.885 -0.89 22.145 -0.66 ;
      RECT 21.885 -0.86 23.22 -0.69 ;
      RECT 23.05 -1.01 26.495 -0.84 ;
      RECT 21.375 -0.35 21.695 -0.09 ;
      RECT 21.1 -0.29 21.695 -0.15 ;
      RECT 20.77 -0.01 21.11 0.33 ;
      RECT 18.995 -0.01 19.315 0.25 ;
      RECT 20.77 0.005 21.26 0.235 ;
      RECT 18.995 0.05 21.26 0.19 ;
      RECT 20.355 2.71 20.675 2.97 ;
      RECT 20.355 2.77 20.95 2.91 ;
      RECT 19.675 -0.35 19.995 -0.09 ;
      RECT 14.935 -0.335 15.225 -0.105 ;
      RECT 14.935 -0.29 19.995 -0.15 ;
      RECT 19.765 -0.63 19.905 -0.09 ;
      RECT 19.765 -0.63 20.245 -0.49 ;
      RECT 20.105 -1.015 20.245 -0.49 ;
      RECT 20.03 -1.015 20.32 -0.785 ;
      RECT 19.675 0.67 19.995 0.93 ;
      RECT 19.01 0.685 19.3 0.915 ;
      RECT 16.8 0.685 17.09 0.915 ;
      RECT 16.8 0.73 19.995 0.87 ;
      RECT 17.975 2.71 18.295 2.97 ;
      RECT 19.69 2.725 19.98 2.955 ;
      RECT 17.31 2.725 17.6 2.955 ;
      RECT 17.31 2.77 18.295 2.91 ;
      RECT 19.765 2.43 19.905 2.955 ;
      RECT 18.065 2.43 18.205 2.97 ;
      RECT 18.065 2.43 19.905 2.57 ;
      RECT 16.97 -0.675 17.26 -0.445 ;
      RECT 17.045 -0.97 17.185 -0.445 ;
      RECT 19.335 -1.03 19.655 -0.77 ;
      RECT 19.235 -1.015 19.655 -0.785 ;
      RECT 17.045 -0.97 19.655 -0.83 ;
      RECT 18.315 -0.69 18.635 -0.43 ;
      RECT 18.315 -0.63 18.91 -0.49 ;
      RECT 18.315 1.69 18.635 1.95 ;
      RECT 15.61 1.705 15.9 1.935 ;
      RECT 15.61 1.75 18.635 1.89 ;
      RECT 17.64 -0.73 17.97 -0.4 ;
      RECT 17.635 -0.695 17.97 -0.435 ;
      RECT 17.985 -0.675 18.1 -0.445 ;
      RECT 17.635 -0.68 17.985 -0.45 ;
      RECT 17.635 -0.63 18.115 -0.49 ;
      RECT 17.52 -0.63 17.53 -0.49 ;
      RECT 17.53 -0.635 18.1 -0.495 ;
      RECT -0.015 4.855 0.415 5.275 ;
      RECT -1.855 4.925 0.415 5.115 ;
      RECT -1.855 4.645 -1.65 5.115 ;
      RECT -1.885 4.645 -1.65 4.875 ;
      RECT -1.855 4.615 -1.685 5.115 ;
      RECT -3.95 0.06 0.325 0.54 ;
      RECT -3.95 0.215 0.405 0.39 ;
      RECT -1.51 2.78 -1.32 4.365 ;
      RECT -1.53 4.07 -1.29 4.325 ;
      RECT -3.95 2.78 0.19 3.26 ;
      RECT -3.95 2.935 0.335 3.105 ;
      RECT 10.765 -1.65 100.46 -1.17 ;
      RECT 10.765 1.07 100.46 1.55 ;
      RECT 95.985 -0.01 96.325 0.33 ;
      RECT 95.94 2.26 96.28 2.6 ;
      RECT 95.535 -0.6 95.875 -0.26 ;
      RECT 95.52 2.865 95.86 3.205 ;
      RECT 94.385 2.705 94.725 3.045 ;
      RECT 94.4 -0.415 94.72 -0.095 ;
      RECT 92.805 1.69 93.45 1.95 ;
      RECT 90.75 2.71 91.07 2.97 ;
      RECT 89.24 4.86 89.67 5.28 ;
      RECT 86.335 2.67 86.705 3.04 ;
      RECT 84.805 2.165 85.175 2.535 ;
      RECT 83.1 2.31 83.47 2.68 ;
      RECT 78.045 -0.01 78.385 0.33 ;
      RECT 78 2.26 78.34 2.6 ;
      RECT 77.595 -0.6 77.935 -0.26 ;
      RECT 77.58 2.865 77.92 3.205 ;
      RECT 76.445 2.705 76.785 3.045 ;
      RECT 76.46 -0.415 76.78 -0.095 ;
      RECT 74.865 1.69 75.51 1.95 ;
      RECT 72.81 2.71 73.13 2.97 ;
      RECT 68.395 2.67 68.765 3.04 ;
      RECT 66.865 2.165 67.235 2.535 ;
      RECT 65.16 2.31 65.53 2.68 ;
      RECT 60.11 -0.01 60.45 0.33 ;
      RECT 60.065 2.26 60.405 2.6 ;
      RECT 59.66 -0.6 60 -0.26 ;
      RECT 59.645 2.865 59.985 3.205 ;
      RECT 58.51 2.705 58.85 3.045 ;
      RECT 58.525 -0.415 58.845 -0.095 ;
      RECT 56.93 1.69 57.575 1.95 ;
      RECT 54.875 2.71 55.195 2.97 ;
      RECT 50.46 2.67 50.83 3.04 ;
      RECT 48.93 2.165 49.3 2.535 ;
      RECT 47.225 2.31 47.595 2.68 ;
      RECT 42.17 -0.01 42.51 0.33 ;
      RECT 42.125 2.26 42.465 2.6 ;
      RECT 41.72 -0.6 42.06 -0.26 ;
      RECT 41.705 2.865 42.045 3.205 ;
      RECT 40.57 2.705 40.91 3.045 ;
      RECT 40.585 -0.415 40.905 -0.095 ;
      RECT 38.99 1.69 39.635 1.95 ;
      RECT 36.935 2.71 37.255 2.97 ;
      RECT 32.52 2.67 32.89 3.04 ;
      RECT 30.99 2.165 31.36 2.535 ;
      RECT 29.285 2.31 29.655 2.68 ;
      RECT 24.23 -0.01 24.57 0.33 ;
      RECT 24.185 2.26 24.525 2.6 ;
      RECT 23.78 -0.6 24.12 -0.26 ;
      RECT 23.765 2.865 24.105 3.205 ;
      RECT 22.63 2.705 22.97 3.045 ;
      RECT 22.645 -0.415 22.965 -0.095 ;
      RECT 21.05 1.69 21.695 1.95 ;
      RECT 18.995 2.71 19.315 2.97 ;
      RECT 14.58 2.67 14.95 3.04 ;
      RECT 13.05 2.165 13.42 2.535 ;
      RECT 11.345 2.31 11.715 2.68 ;
      RECT -3.95 5.5 0.19 5.98 ;
      RECT -3.885 3.55 -3.505 3.93 ;
    LAYER mcon ;
      RECT 100.145 -1.495 100.315 -1.325 ;
      RECT 100.145 1.225 100.315 1.395 ;
      RECT 100.145 3.945 100.315 4.115 ;
      RECT 99.685 -1.495 99.855 -1.325 ;
      RECT 99.685 1.225 99.855 1.395 ;
      RECT 99.685 3.945 99.855 4.115 ;
      RECT 99.225 -1.495 99.395 -1.325 ;
      RECT 99.225 1.225 99.395 1.395 ;
      RECT 99.225 3.945 99.395 4.115 ;
      RECT 98.765 -1.495 98.935 -1.325 ;
      RECT 98.765 1.225 98.935 1.395 ;
      RECT 98.765 3.945 98.935 4.115 ;
      RECT 98.305 -1.495 98.475 -1.325 ;
      RECT 98.305 1.225 98.475 1.395 ;
      RECT 98.305 3.945 98.475 4.115 ;
      RECT 98.1 2.785 98.27 2.955 ;
      RECT 98.08 -0.335 98.25 -0.165 ;
      RECT 97.845 -1.495 98.015 -1.325 ;
      RECT 97.845 1.225 98.015 1.395 ;
      RECT 97.845 3.945 98.015 4.115 ;
      RECT 97.385 -1.495 97.555 -1.325 ;
      RECT 97.385 1.225 97.555 1.395 ;
      RECT 97.385 3.945 97.555 4.115 ;
      RECT 96.925 -1.495 97.095 -1.325 ;
      RECT 96.925 1.225 97.095 1.395 ;
      RECT 96.925 3.945 97.095 4.115 ;
      RECT 96.465 -1.495 96.635 -1.325 ;
      RECT 96.465 1.225 96.635 1.395 ;
      RECT 96.465 3.945 96.635 4.115 ;
      RECT 96.015 0.05 96.185 0.22 ;
      RECT 96.015 2.4 96.185 2.57 ;
      RECT 96.005 -1.495 96.175 -1.325 ;
      RECT 96.005 1.225 96.175 1.395 ;
      RECT 96.005 3.945 96.175 4.115 ;
      RECT 95.655 -0.515 95.825 -0.345 ;
      RECT 95.655 2.965 95.825 3.135 ;
      RECT 95.545 -1.495 95.715 -1.325 ;
      RECT 95.545 1.225 95.715 1.395 ;
      RECT 95.545 3.945 95.715 4.115 ;
      RECT 95.085 -1.495 95.255 -1.325 ;
      RECT 95.085 1.225 95.255 1.395 ;
      RECT 95.085 3.945 95.255 4.115 ;
      RECT 94.625 -1.495 94.795 -1.325 ;
      RECT 94.625 1.225 94.795 1.395 ;
      RECT 94.625 3.945 94.795 4.115 ;
      RECT 94.47 -0.335 94.64 -0.165 ;
      RECT 94.47 2.785 94.64 2.955 ;
      RECT 94.165 -1.495 94.335 -1.325 ;
      RECT 94.165 1.225 94.335 1.395 ;
      RECT 94.165 3.945 94.335 4.115 ;
      RECT 93.735 3.32 93.905 3.49 ;
      RECT 93.705 -1.495 93.875 -1.325 ;
      RECT 93.705 1.225 93.875 1.395 ;
      RECT 93.705 3.945 93.875 4.115 ;
      RECT 93.7 -0.86 93.87 -0.69 ;
      RECT 93.245 -1.495 93.415 -1.325 ;
      RECT 93.245 1.225 93.415 1.395 ;
      RECT 93.245 3.945 93.415 4.115 ;
      RECT 93.205 -0.305 93.375 -0.135 ;
      RECT 92.865 1.735 93.035 1.905 ;
      RECT 92.785 -1.495 92.955 -1.325 ;
      RECT 92.785 0.035 92.955 0.205 ;
      RECT 92.785 1.225 92.955 1.395 ;
      RECT 92.785 3.945 92.955 4.115 ;
      RECT 92.325 -1.495 92.495 -1.325 ;
      RECT 92.325 1.225 92.495 1.395 ;
      RECT 92.325 3.945 92.495 4.115 ;
      RECT 92.185 2.755 92.355 2.925 ;
      RECT 91.865 -1.495 92.035 -1.325 ;
      RECT 91.865 1.225 92.035 1.395 ;
      RECT 91.865 3.945 92.035 4.115 ;
      RECT 91.845 -0.985 92.015 -0.815 ;
      RECT 91.505 2.755 91.675 2.925 ;
      RECT 91.405 -1.495 91.575 -1.325 ;
      RECT 91.405 1.225 91.575 1.395 ;
      RECT 91.405 3.945 91.575 4.115 ;
      RECT 91.05 -0.985 91.22 -0.815 ;
      RECT 90.945 -1.495 91.115 -1.325 ;
      RECT 90.945 1.225 91.115 1.395 ;
      RECT 90.945 3.945 91.115 4.115 ;
      RECT 90.825 0.715 90.995 0.885 ;
      RECT 90.825 2.755 90.995 2.925 ;
      RECT 90.485 -1.495 90.655 -1.325 ;
      RECT 90.485 1.225 90.655 1.395 ;
      RECT 90.485 3.945 90.655 4.115 ;
      RECT 90.315 2.755 90.485 2.925 ;
      RECT 90.145 -0.645 90.315 -0.475 ;
      RECT 90.025 -1.495 90.195 -1.325 ;
      RECT 90.025 1.225 90.195 1.395 ;
      RECT 90.025 3.945 90.195 4.115 ;
      RECT 89.565 -1.495 89.735 -1.325 ;
      RECT 89.565 1.225 89.735 1.395 ;
      RECT 89.565 3.945 89.735 4.115 ;
      RECT 89.305 4.915 89.475 5.085 ;
      RECT 89.125 2.755 89.295 2.925 ;
      RECT 89.105 -1.495 89.275 -1.325 ;
      RECT 89.105 1.225 89.275 1.395 ;
      RECT 89.105 3.945 89.275 4.115 ;
      RECT 88.785 -0.645 88.955 -0.475 ;
      RECT 88.645 -1.495 88.815 -1.325 ;
      RECT 88.645 1.225 88.815 1.395 ;
      RECT 88.645 3.945 88.815 4.115 ;
      RECT 88.615 0.715 88.785 0.885 ;
      RECT 88.185 -1.495 88.355 -1.325 ;
      RECT 88.185 1.225 88.355 1.395 ;
      RECT 88.185 3.945 88.355 4.115 ;
      RECT 88.105 2.755 88.275 2.925 ;
      RECT 87.725 -1.495 87.895 -1.325 ;
      RECT 87.725 1.225 87.895 1.395 ;
      RECT 87.725 3.945 87.895 4.115 ;
      RECT 87.425 1.735 87.595 1.905 ;
      RECT 87.265 -1.495 87.435 -1.325 ;
      RECT 87.265 1.225 87.435 1.395 ;
      RECT 87.265 3.945 87.435 4.115 ;
      RECT 86.805 -1.495 86.975 -1.325 ;
      RECT 86.805 1.225 86.975 1.395 ;
      RECT 86.805 3.945 86.975 4.115 ;
      RECT 86.75 -0.305 86.92 -0.135 ;
      RECT 86.405 2.775 86.575 2.945 ;
      RECT 86.345 1.225 86.515 1.395 ;
      RECT 86.345 3.945 86.515 4.115 ;
      RECT 85.885 1.225 86.055 1.395 ;
      RECT 85.885 3.945 86.055 4.115 ;
      RECT 85.425 1.225 85.595 1.395 ;
      RECT 85.425 3.945 85.595 4.115 ;
      RECT 84.965 1.225 85.135 1.395 ;
      RECT 84.965 3.945 85.135 4.115 ;
      RECT 84.875 2.27 85.045 2.44 ;
      RECT 84.505 1.225 84.675 1.395 ;
      RECT 84.505 3.945 84.675 4.115 ;
      RECT 84.045 1.225 84.215 1.395 ;
      RECT 84.045 3.945 84.215 4.115 ;
      RECT 83.585 1.225 83.755 1.395 ;
      RECT 83.585 3.945 83.755 4.115 ;
      RECT 83.195 2.4 83.365 2.57 ;
      RECT 83.125 1.225 83.295 1.395 ;
      RECT 83.125 3.945 83.295 4.115 ;
      RECT 82.665 1.225 82.835 1.395 ;
      RECT 82.665 3.945 82.835 4.115 ;
      RECT 82.205 -1.495 82.375 -1.325 ;
      RECT 82.205 1.225 82.375 1.395 ;
      RECT 82.205 3.945 82.375 4.115 ;
      RECT 81.745 -1.495 81.915 -1.325 ;
      RECT 81.745 1.225 81.915 1.395 ;
      RECT 81.745 3.945 81.915 4.115 ;
      RECT 81.285 -1.495 81.455 -1.325 ;
      RECT 81.285 1.225 81.455 1.395 ;
      RECT 81.285 3.945 81.455 4.115 ;
      RECT 80.825 -1.495 80.995 -1.325 ;
      RECT 80.825 1.225 80.995 1.395 ;
      RECT 80.825 3.945 80.995 4.115 ;
      RECT 80.365 -1.495 80.535 -1.325 ;
      RECT 80.365 1.225 80.535 1.395 ;
      RECT 80.365 3.945 80.535 4.115 ;
      RECT 80.16 2.785 80.33 2.955 ;
      RECT 80.14 -0.335 80.31 -0.165 ;
      RECT 79.905 -1.495 80.075 -1.325 ;
      RECT 79.905 1.225 80.075 1.395 ;
      RECT 79.905 3.945 80.075 4.115 ;
      RECT 79.445 -1.495 79.615 -1.325 ;
      RECT 79.445 1.225 79.615 1.395 ;
      RECT 79.445 3.945 79.615 4.115 ;
      RECT 78.985 -1.495 79.155 -1.325 ;
      RECT 78.985 1.225 79.155 1.395 ;
      RECT 78.985 3.945 79.155 4.115 ;
      RECT 78.525 -1.495 78.695 -1.325 ;
      RECT 78.525 1.225 78.695 1.395 ;
      RECT 78.525 3.945 78.695 4.115 ;
      RECT 78.075 0.05 78.245 0.22 ;
      RECT 78.075 2.4 78.245 2.57 ;
      RECT 78.065 -1.495 78.235 -1.325 ;
      RECT 78.065 1.225 78.235 1.395 ;
      RECT 78.065 3.945 78.235 4.115 ;
      RECT 77.715 -0.515 77.885 -0.345 ;
      RECT 77.715 2.965 77.885 3.135 ;
      RECT 77.605 -1.495 77.775 -1.325 ;
      RECT 77.605 1.225 77.775 1.395 ;
      RECT 77.605 3.945 77.775 4.115 ;
      RECT 77.145 -1.495 77.315 -1.325 ;
      RECT 77.145 1.225 77.315 1.395 ;
      RECT 77.145 3.945 77.315 4.115 ;
      RECT 76.685 -1.495 76.855 -1.325 ;
      RECT 76.685 1.225 76.855 1.395 ;
      RECT 76.685 3.945 76.855 4.115 ;
      RECT 76.53 -0.335 76.7 -0.165 ;
      RECT 76.53 2.785 76.7 2.955 ;
      RECT 76.225 -1.495 76.395 -1.325 ;
      RECT 76.225 1.225 76.395 1.395 ;
      RECT 76.225 3.945 76.395 4.115 ;
      RECT 75.795 3.32 75.965 3.49 ;
      RECT 75.765 -1.495 75.935 -1.325 ;
      RECT 75.765 1.225 75.935 1.395 ;
      RECT 75.765 3.945 75.935 4.115 ;
      RECT 75.76 -0.86 75.93 -0.69 ;
      RECT 75.305 -1.495 75.475 -1.325 ;
      RECT 75.305 1.225 75.475 1.395 ;
      RECT 75.305 3.945 75.475 4.115 ;
      RECT 75.265 -0.305 75.435 -0.135 ;
      RECT 74.925 1.735 75.095 1.905 ;
      RECT 74.845 -1.495 75.015 -1.325 ;
      RECT 74.845 0.035 75.015 0.205 ;
      RECT 74.845 1.225 75.015 1.395 ;
      RECT 74.845 3.945 75.015 4.115 ;
      RECT 74.385 -1.495 74.555 -1.325 ;
      RECT 74.385 1.225 74.555 1.395 ;
      RECT 74.385 3.945 74.555 4.115 ;
      RECT 74.245 2.755 74.415 2.925 ;
      RECT 73.925 -1.495 74.095 -1.325 ;
      RECT 73.925 1.225 74.095 1.395 ;
      RECT 73.925 3.945 74.095 4.115 ;
      RECT 73.905 -0.985 74.075 -0.815 ;
      RECT 73.565 2.755 73.735 2.925 ;
      RECT 73.465 -1.495 73.635 -1.325 ;
      RECT 73.465 1.225 73.635 1.395 ;
      RECT 73.465 3.945 73.635 4.115 ;
      RECT 73.11 -0.985 73.28 -0.815 ;
      RECT 73.005 -1.495 73.175 -1.325 ;
      RECT 73.005 1.225 73.175 1.395 ;
      RECT 73.005 3.945 73.175 4.115 ;
      RECT 72.885 0.715 73.055 0.885 ;
      RECT 72.885 2.755 73.055 2.925 ;
      RECT 72.545 -1.495 72.715 -1.325 ;
      RECT 72.545 1.225 72.715 1.395 ;
      RECT 72.545 3.945 72.715 4.115 ;
      RECT 72.375 2.755 72.545 2.925 ;
      RECT 72.205 -0.645 72.375 -0.475 ;
      RECT 72.085 -1.495 72.255 -1.325 ;
      RECT 72.085 1.225 72.255 1.395 ;
      RECT 72.085 3.945 72.255 4.115 ;
      RECT 71.625 -1.495 71.795 -1.325 ;
      RECT 71.625 1.225 71.795 1.395 ;
      RECT 71.625 3.945 71.795 4.115 ;
      RECT 71.365 3.655 71.535 3.825 ;
      RECT 71.185 2.755 71.355 2.925 ;
      RECT 71.165 -1.495 71.335 -1.325 ;
      RECT 71.165 1.225 71.335 1.395 ;
      RECT 71.165 3.945 71.335 4.115 ;
      RECT 70.845 -0.645 71.015 -0.475 ;
      RECT 70.705 -1.495 70.875 -1.325 ;
      RECT 70.705 1.225 70.875 1.395 ;
      RECT 70.705 3.945 70.875 4.115 ;
      RECT 70.675 0.715 70.845 0.885 ;
      RECT 70.245 -1.495 70.415 -1.325 ;
      RECT 70.245 1.225 70.415 1.395 ;
      RECT 70.245 3.945 70.415 4.115 ;
      RECT 70.165 2.755 70.335 2.925 ;
      RECT 69.785 -1.495 69.955 -1.325 ;
      RECT 69.785 1.225 69.955 1.395 ;
      RECT 69.785 3.945 69.955 4.115 ;
      RECT 69.485 1.735 69.655 1.905 ;
      RECT 69.325 -1.495 69.495 -1.325 ;
      RECT 69.325 1.225 69.495 1.395 ;
      RECT 69.325 3.945 69.495 4.115 ;
      RECT 68.865 -1.495 69.035 -1.325 ;
      RECT 68.865 1.225 69.035 1.395 ;
      RECT 68.865 3.945 69.035 4.115 ;
      RECT 68.81 -0.305 68.98 -0.135 ;
      RECT 68.465 2.775 68.635 2.945 ;
      RECT 68.405 1.225 68.575 1.395 ;
      RECT 68.405 3.945 68.575 4.115 ;
      RECT 67.945 1.225 68.115 1.395 ;
      RECT 67.945 3.945 68.115 4.115 ;
      RECT 67.485 1.225 67.655 1.395 ;
      RECT 67.485 3.945 67.655 4.115 ;
      RECT 67.025 1.225 67.195 1.395 ;
      RECT 67.025 3.945 67.195 4.115 ;
      RECT 66.935 2.27 67.105 2.44 ;
      RECT 66.565 1.225 66.735 1.395 ;
      RECT 66.565 3.945 66.735 4.115 ;
      RECT 66.105 1.225 66.275 1.395 ;
      RECT 66.105 3.945 66.275 4.115 ;
      RECT 65.645 1.225 65.815 1.395 ;
      RECT 65.645 3.945 65.815 4.115 ;
      RECT 65.255 2.4 65.425 2.57 ;
      RECT 65.185 1.225 65.355 1.395 ;
      RECT 65.185 3.945 65.355 4.115 ;
      RECT 64.725 1.225 64.895 1.395 ;
      RECT 64.725 3.945 64.895 4.115 ;
      RECT 64.27 -1.495 64.44 -1.325 ;
      RECT 64.27 1.225 64.44 1.395 ;
      RECT 64.27 3.945 64.44 4.115 ;
      RECT 63.81 -1.495 63.98 -1.325 ;
      RECT 63.81 1.225 63.98 1.395 ;
      RECT 63.81 3.945 63.98 4.115 ;
      RECT 63.35 -1.495 63.52 -1.325 ;
      RECT 63.35 1.225 63.52 1.395 ;
      RECT 63.35 3.945 63.52 4.115 ;
      RECT 62.89 -1.495 63.06 -1.325 ;
      RECT 62.89 1.225 63.06 1.395 ;
      RECT 62.89 3.945 63.06 4.115 ;
      RECT 62.43 -1.495 62.6 -1.325 ;
      RECT 62.43 1.225 62.6 1.395 ;
      RECT 62.43 3.945 62.6 4.115 ;
      RECT 62.225 2.785 62.395 2.955 ;
      RECT 62.205 -0.335 62.375 -0.165 ;
      RECT 61.97 -1.495 62.14 -1.325 ;
      RECT 61.97 1.225 62.14 1.395 ;
      RECT 61.97 3.945 62.14 4.115 ;
      RECT 61.51 -1.495 61.68 -1.325 ;
      RECT 61.51 1.225 61.68 1.395 ;
      RECT 61.51 3.945 61.68 4.115 ;
      RECT 61.05 -1.495 61.22 -1.325 ;
      RECT 61.05 1.225 61.22 1.395 ;
      RECT 61.05 3.945 61.22 4.115 ;
      RECT 60.59 -1.495 60.76 -1.325 ;
      RECT 60.59 1.225 60.76 1.395 ;
      RECT 60.59 3.945 60.76 4.115 ;
      RECT 60.14 0.05 60.31 0.22 ;
      RECT 60.14 2.4 60.31 2.57 ;
      RECT 60.13 -1.495 60.3 -1.325 ;
      RECT 60.13 1.225 60.3 1.395 ;
      RECT 60.13 3.945 60.3 4.115 ;
      RECT 59.78 -0.515 59.95 -0.345 ;
      RECT 59.78 2.965 59.95 3.135 ;
      RECT 59.67 -1.495 59.84 -1.325 ;
      RECT 59.67 1.225 59.84 1.395 ;
      RECT 59.67 3.945 59.84 4.115 ;
      RECT 59.21 -1.495 59.38 -1.325 ;
      RECT 59.21 1.225 59.38 1.395 ;
      RECT 59.21 3.945 59.38 4.115 ;
      RECT 58.75 -1.495 58.92 -1.325 ;
      RECT 58.75 1.225 58.92 1.395 ;
      RECT 58.75 3.945 58.92 4.115 ;
      RECT 58.595 -0.335 58.765 -0.165 ;
      RECT 58.595 2.785 58.765 2.955 ;
      RECT 58.29 -1.495 58.46 -1.325 ;
      RECT 58.29 1.225 58.46 1.395 ;
      RECT 58.29 3.945 58.46 4.115 ;
      RECT 57.86 3.32 58.03 3.49 ;
      RECT 57.83 -1.495 58 -1.325 ;
      RECT 57.83 1.225 58 1.395 ;
      RECT 57.83 3.945 58 4.115 ;
      RECT 57.825 -0.86 57.995 -0.69 ;
      RECT 57.37 -1.495 57.54 -1.325 ;
      RECT 57.37 1.225 57.54 1.395 ;
      RECT 57.37 3.945 57.54 4.115 ;
      RECT 57.33 -0.305 57.5 -0.135 ;
      RECT 56.99 1.735 57.16 1.905 ;
      RECT 56.91 -1.495 57.08 -1.325 ;
      RECT 56.91 0.035 57.08 0.205 ;
      RECT 56.91 1.225 57.08 1.395 ;
      RECT 56.91 3.945 57.08 4.115 ;
      RECT 56.45 -1.495 56.62 -1.325 ;
      RECT 56.45 1.225 56.62 1.395 ;
      RECT 56.45 3.945 56.62 4.115 ;
      RECT 56.31 2.755 56.48 2.925 ;
      RECT 55.99 -1.495 56.16 -1.325 ;
      RECT 55.99 1.225 56.16 1.395 ;
      RECT 55.99 3.945 56.16 4.115 ;
      RECT 55.97 -0.985 56.14 -0.815 ;
      RECT 55.63 2.755 55.8 2.925 ;
      RECT 55.53 -1.495 55.7 -1.325 ;
      RECT 55.53 1.225 55.7 1.395 ;
      RECT 55.53 3.945 55.7 4.115 ;
      RECT 55.175 -0.985 55.345 -0.815 ;
      RECT 55.07 -1.495 55.24 -1.325 ;
      RECT 55.07 1.225 55.24 1.395 ;
      RECT 55.07 3.945 55.24 4.115 ;
      RECT 54.95 0.715 55.12 0.885 ;
      RECT 54.95 2.755 55.12 2.925 ;
      RECT 54.61 -1.495 54.78 -1.325 ;
      RECT 54.61 1.225 54.78 1.395 ;
      RECT 54.61 3.945 54.78 4.115 ;
      RECT 54.44 2.755 54.61 2.925 ;
      RECT 54.27 -0.645 54.44 -0.475 ;
      RECT 54.15 -1.495 54.32 -1.325 ;
      RECT 54.15 1.225 54.32 1.395 ;
      RECT 54.15 3.945 54.32 4.115 ;
      RECT 53.69 -1.495 53.86 -1.325 ;
      RECT 53.69 1.225 53.86 1.395 ;
      RECT 53.69 3.945 53.86 4.115 ;
      RECT 53.43 3.655 53.6 3.825 ;
      RECT 53.25 2.755 53.42 2.925 ;
      RECT 53.23 -1.495 53.4 -1.325 ;
      RECT 53.23 1.225 53.4 1.395 ;
      RECT 53.23 3.945 53.4 4.115 ;
      RECT 52.91 -0.645 53.08 -0.475 ;
      RECT 52.77 -1.495 52.94 -1.325 ;
      RECT 52.77 1.225 52.94 1.395 ;
      RECT 52.77 3.945 52.94 4.115 ;
      RECT 52.74 0.715 52.91 0.885 ;
      RECT 52.31 -1.495 52.48 -1.325 ;
      RECT 52.31 1.225 52.48 1.395 ;
      RECT 52.31 3.945 52.48 4.115 ;
      RECT 52.23 2.755 52.4 2.925 ;
      RECT 51.85 -1.495 52.02 -1.325 ;
      RECT 51.85 1.225 52.02 1.395 ;
      RECT 51.85 3.945 52.02 4.115 ;
      RECT 51.55 1.735 51.72 1.905 ;
      RECT 51.39 -1.495 51.56 -1.325 ;
      RECT 51.39 1.225 51.56 1.395 ;
      RECT 51.39 3.945 51.56 4.115 ;
      RECT 50.93 -1.495 51.1 -1.325 ;
      RECT 50.93 1.225 51.1 1.395 ;
      RECT 50.93 3.945 51.1 4.115 ;
      RECT 50.875 -0.305 51.045 -0.135 ;
      RECT 50.53 2.775 50.7 2.945 ;
      RECT 50.47 1.225 50.64 1.395 ;
      RECT 50.47 3.945 50.64 4.115 ;
      RECT 50.01 1.225 50.18 1.395 ;
      RECT 50.01 3.945 50.18 4.115 ;
      RECT 49.55 1.225 49.72 1.395 ;
      RECT 49.55 3.945 49.72 4.115 ;
      RECT 49.09 1.225 49.26 1.395 ;
      RECT 49.09 3.945 49.26 4.115 ;
      RECT 49 2.27 49.17 2.44 ;
      RECT 48.63 1.225 48.8 1.395 ;
      RECT 48.63 3.945 48.8 4.115 ;
      RECT 48.17 1.225 48.34 1.395 ;
      RECT 48.17 3.945 48.34 4.115 ;
      RECT 47.71 1.225 47.88 1.395 ;
      RECT 47.71 3.945 47.88 4.115 ;
      RECT 47.32 2.4 47.49 2.57 ;
      RECT 47.25 1.225 47.42 1.395 ;
      RECT 47.25 3.945 47.42 4.115 ;
      RECT 46.79 1.225 46.96 1.395 ;
      RECT 46.79 3.945 46.96 4.115 ;
      RECT 46.33 -1.495 46.5 -1.325 ;
      RECT 46.33 1.225 46.5 1.395 ;
      RECT 46.33 3.945 46.5 4.115 ;
      RECT 45.87 -1.495 46.04 -1.325 ;
      RECT 45.87 1.225 46.04 1.395 ;
      RECT 45.87 3.945 46.04 4.115 ;
      RECT 45.41 -1.495 45.58 -1.325 ;
      RECT 45.41 1.225 45.58 1.395 ;
      RECT 45.41 3.945 45.58 4.115 ;
      RECT 44.95 -1.495 45.12 -1.325 ;
      RECT 44.95 1.225 45.12 1.395 ;
      RECT 44.95 3.945 45.12 4.115 ;
      RECT 44.49 -1.495 44.66 -1.325 ;
      RECT 44.49 1.225 44.66 1.395 ;
      RECT 44.49 3.945 44.66 4.115 ;
      RECT 44.285 2.785 44.455 2.955 ;
      RECT 44.265 -0.335 44.435 -0.165 ;
      RECT 44.03 -1.495 44.2 -1.325 ;
      RECT 44.03 1.225 44.2 1.395 ;
      RECT 44.03 3.945 44.2 4.115 ;
      RECT 43.57 -1.495 43.74 -1.325 ;
      RECT 43.57 1.225 43.74 1.395 ;
      RECT 43.57 3.945 43.74 4.115 ;
      RECT 43.11 -1.495 43.28 -1.325 ;
      RECT 43.11 1.225 43.28 1.395 ;
      RECT 43.11 3.945 43.28 4.115 ;
      RECT 42.65 -1.495 42.82 -1.325 ;
      RECT 42.65 1.225 42.82 1.395 ;
      RECT 42.65 3.945 42.82 4.115 ;
      RECT 42.2 0.05 42.37 0.22 ;
      RECT 42.2 2.4 42.37 2.57 ;
      RECT 42.19 -1.495 42.36 -1.325 ;
      RECT 42.19 1.225 42.36 1.395 ;
      RECT 42.19 3.945 42.36 4.115 ;
      RECT 41.84 -0.515 42.01 -0.345 ;
      RECT 41.84 2.965 42.01 3.135 ;
      RECT 41.73 -1.495 41.9 -1.325 ;
      RECT 41.73 1.225 41.9 1.395 ;
      RECT 41.73 3.945 41.9 4.115 ;
      RECT 41.27 -1.495 41.44 -1.325 ;
      RECT 41.27 1.225 41.44 1.395 ;
      RECT 41.27 3.945 41.44 4.115 ;
      RECT 40.81 -1.495 40.98 -1.325 ;
      RECT 40.81 1.225 40.98 1.395 ;
      RECT 40.81 3.945 40.98 4.115 ;
      RECT 40.655 -0.335 40.825 -0.165 ;
      RECT 40.655 2.785 40.825 2.955 ;
      RECT 40.35 -1.495 40.52 -1.325 ;
      RECT 40.35 1.225 40.52 1.395 ;
      RECT 40.35 3.945 40.52 4.115 ;
      RECT 39.92 3.32 40.09 3.49 ;
      RECT 39.89 -1.495 40.06 -1.325 ;
      RECT 39.89 1.225 40.06 1.395 ;
      RECT 39.89 3.945 40.06 4.115 ;
      RECT 39.885 -0.86 40.055 -0.69 ;
      RECT 39.43 -1.495 39.6 -1.325 ;
      RECT 39.43 1.225 39.6 1.395 ;
      RECT 39.43 3.945 39.6 4.115 ;
      RECT 39.39 -0.305 39.56 -0.135 ;
      RECT 39.05 1.735 39.22 1.905 ;
      RECT 38.97 -1.495 39.14 -1.325 ;
      RECT 38.97 0.035 39.14 0.205 ;
      RECT 38.97 1.225 39.14 1.395 ;
      RECT 38.97 3.945 39.14 4.115 ;
      RECT 38.51 -1.495 38.68 -1.325 ;
      RECT 38.51 1.225 38.68 1.395 ;
      RECT 38.51 3.945 38.68 4.115 ;
      RECT 38.37 2.755 38.54 2.925 ;
      RECT 38.05 -1.495 38.22 -1.325 ;
      RECT 38.05 1.225 38.22 1.395 ;
      RECT 38.05 3.945 38.22 4.115 ;
      RECT 38.03 -0.985 38.2 -0.815 ;
      RECT 37.69 2.755 37.86 2.925 ;
      RECT 37.59 -1.495 37.76 -1.325 ;
      RECT 37.59 1.225 37.76 1.395 ;
      RECT 37.59 3.945 37.76 4.115 ;
      RECT 37.235 -0.985 37.405 -0.815 ;
      RECT 37.13 -1.495 37.3 -1.325 ;
      RECT 37.13 1.225 37.3 1.395 ;
      RECT 37.13 3.945 37.3 4.115 ;
      RECT 37.01 0.715 37.18 0.885 ;
      RECT 37.01 2.755 37.18 2.925 ;
      RECT 36.67 -1.495 36.84 -1.325 ;
      RECT 36.67 1.225 36.84 1.395 ;
      RECT 36.67 3.945 36.84 4.115 ;
      RECT 36.5 2.755 36.67 2.925 ;
      RECT 36.33 -0.645 36.5 -0.475 ;
      RECT 36.21 -1.495 36.38 -1.325 ;
      RECT 36.21 1.225 36.38 1.395 ;
      RECT 36.21 3.945 36.38 4.115 ;
      RECT 35.75 -1.495 35.92 -1.325 ;
      RECT 35.75 1.225 35.92 1.395 ;
      RECT 35.75 3.945 35.92 4.115 ;
      RECT 35.49 3.655 35.66 3.825 ;
      RECT 35.31 2.755 35.48 2.925 ;
      RECT 35.29 -1.495 35.46 -1.325 ;
      RECT 35.29 1.225 35.46 1.395 ;
      RECT 35.29 3.945 35.46 4.115 ;
      RECT 34.97 -0.645 35.14 -0.475 ;
      RECT 34.83 -1.495 35 -1.325 ;
      RECT 34.83 1.225 35 1.395 ;
      RECT 34.83 3.945 35 4.115 ;
      RECT 34.8 0.715 34.97 0.885 ;
      RECT 34.37 -1.495 34.54 -1.325 ;
      RECT 34.37 1.225 34.54 1.395 ;
      RECT 34.37 3.945 34.54 4.115 ;
      RECT 34.29 2.755 34.46 2.925 ;
      RECT 33.91 -1.495 34.08 -1.325 ;
      RECT 33.91 1.225 34.08 1.395 ;
      RECT 33.91 3.945 34.08 4.115 ;
      RECT 33.61 1.735 33.78 1.905 ;
      RECT 33.45 -1.495 33.62 -1.325 ;
      RECT 33.45 1.225 33.62 1.395 ;
      RECT 33.45 3.945 33.62 4.115 ;
      RECT 32.99 -1.495 33.16 -1.325 ;
      RECT 32.99 1.225 33.16 1.395 ;
      RECT 32.99 3.945 33.16 4.115 ;
      RECT 32.935 -0.305 33.105 -0.135 ;
      RECT 32.59 2.775 32.76 2.945 ;
      RECT 32.53 1.225 32.7 1.395 ;
      RECT 32.53 3.945 32.7 4.115 ;
      RECT 32.07 1.225 32.24 1.395 ;
      RECT 32.07 3.945 32.24 4.115 ;
      RECT 31.61 1.225 31.78 1.395 ;
      RECT 31.61 3.945 31.78 4.115 ;
      RECT 31.15 1.225 31.32 1.395 ;
      RECT 31.15 3.945 31.32 4.115 ;
      RECT 31.06 2.27 31.23 2.44 ;
      RECT 30.69 1.225 30.86 1.395 ;
      RECT 30.69 3.945 30.86 4.115 ;
      RECT 30.23 1.225 30.4 1.395 ;
      RECT 30.23 3.945 30.4 4.115 ;
      RECT 29.77 1.225 29.94 1.395 ;
      RECT 29.77 3.945 29.94 4.115 ;
      RECT 29.38 2.4 29.55 2.57 ;
      RECT 29.31 1.225 29.48 1.395 ;
      RECT 29.31 3.945 29.48 4.115 ;
      RECT 28.85 1.225 29.02 1.395 ;
      RECT 28.85 3.945 29.02 4.115 ;
      RECT 28.39 -1.495 28.56 -1.325 ;
      RECT 28.39 1.225 28.56 1.395 ;
      RECT 28.39 3.945 28.56 4.115 ;
      RECT 27.93 -1.495 28.1 -1.325 ;
      RECT 27.93 1.225 28.1 1.395 ;
      RECT 27.93 3.945 28.1 4.115 ;
      RECT 27.47 -1.495 27.64 -1.325 ;
      RECT 27.47 1.225 27.64 1.395 ;
      RECT 27.47 3.945 27.64 4.115 ;
      RECT 27.01 -1.495 27.18 -1.325 ;
      RECT 27.01 1.225 27.18 1.395 ;
      RECT 27.01 3.945 27.18 4.115 ;
      RECT 26.55 -1.495 26.72 -1.325 ;
      RECT 26.55 1.225 26.72 1.395 ;
      RECT 26.55 3.945 26.72 4.115 ;
      RECT 26.345 2.785 26.515 2.955 ;
      RECT 26.325 -0.335 26.495 -0.165 ;
      RECT 26.09 -1.495 26.26 -1.325 ;
      RECT 26.09 1.225 26.26 1.395 ;
      RECT 26.09 3.945 26.26 4.115 ;
      RECT 25.63 -1.495 25.8 -1.325 ;
      RECT 25.63 1.225 25.8 1.395 ;
      RECT 25.63 3.945 25.8 4.115 ;
      RECT 25.17 -1.495 25.34 -1.325 ;
      RECT 25.17 1.225 25.34 1.395 ;
      RECT 25.17 3.945 25.34 4.115 ;
      RECT 24.71 -1.495 24.88 -1.325 ;
      RECT 24.71 1.225 24.88 1.395 ;
      RECT 24.71 3.945 24.88 4.115 ;
      RECT 24.26 0.05 24.43 0.22 ;
      RECT 24.26 2.4 24.43 2.57 ;
      RECT 24.25 -1.495 24.42 -1.325 ;
      RECT 24.25 1.225 24.42 1.395 ;
      RECT 24.25 3.945 24.42 4.115 ;
      RECT 23.9 -0.515 24.07 -0.345 ;
      RECT 23.9 2.965 24.07 3.135 ;
      RECT 23.79 -1.495 23.96 -1.325 ;
      RECT 23.79 1.225 23.96 1.395 ;
      RECT 23.79 3.945 23.96 4.115 ;
      RECT 23.33 -1.495 23.5 -1.325 ;
      RECT 23.33 1.225 23.5 1.395 ;
      RECT 23.33 3.945 23.5 4.115 ;
      RECT 22.87 -1.495 23.04 -1.325 ;
      RECT 22.87 1.225 23.04 1.395 ;
      RECT 22.87 3.945 23.04 4.115 ;
      RECT 22.715 -0.335 22.885 -0.165 ;
      RECT 22.715 2.785 22.885 2.955 ;
      RECT 22.41 -1.495 22.58 -1.325 ;
      RECT 22.41 1.225 22.58 1.395 ;
      RECT 22.41 3.945 22.58 4.115 ;
      RECT 21.98 3.32 22.15 3.49 ;
      RECT 21.95 -1.495 22.12 -1.325 ;
      RECT 21.95 1.225 22.12 1.395 ;
      RECT 21.95 3.945 22.12 4.115 ;
      RECT 21.945 -0.86 22.115 -0.69 ;
      RECT 21.49 -1.495 21.66 -1.325 ;
      RECT 21.49 1.225 21.66 1.395 ;
      RECT 21.49 3.945 21.66 4.115 ;
      RECT 21.45 -0.305 21.62 -0.135 ;
      RECT 21.11 1.735 21.28 1.905 ;
      RECT 21.03 -1.495 21.2 -1.325 ;
      RECT 21.03 0.035 21.2 0.205 ;
      RECT 21.03 1.225 21.2 1.395 ;
      RECT 21.03 3.945 21.2 4.115 ;
      RECT 20.57 -1.495 20.74 -1.325 ;
      RECT 20.57 1.225 20.74 1.395 ;
      RECT 20.57 3.945 20.74 4.115 ;
      RECT 20.43 2.755 20.6 2.925 ;
      RECT 20.11 -1.495 20.28 -1.325 ;
      RECT 20.11 1.225 20.28 1.395 ;
      RECT 20.11 3.945 20.28 4.115 ;
      RECT 20.09 -0.985 20.26 -0.815 ;
      RECT 19.75 2.755 19.92 2.925 ;
      RECT 19.65 -1.495 19.82 -1.325 ;
      RECT 19.65 1.225 19.82 1.395 ;
      RECT 19.65 3.945 19.82 4.115 ;
      RECT 19.295 -0.985 19.465 -0.815 ;
      RECT 19.19 -1.495 19.36 -1.325 ;
      RECT 19.19 1.225 19.36 1.395 ;
      RECT 19.19 3.945 19.36 4.115 ;
      RECT 19.07 0.715 19.24 0.885 ;
      RECT 19.07 2.755 19.24 2.925 ;
      RECT 18.73 -1.495 18.9 -1.325 ;
      RECT 18.73 1.225 18.9 1.395 ;
      RECT 18.73 3.945 18.9 4.115 ;
      RECT 18.56 2.755 18.73 2.925 ;
      RECT 18.39 -0.645 18.56 -0.475 ;
      RECT 18.27 -1.495 18.44 -1.325 ;
      RECT 18.27 1.225 18.44 1.395 ;
      RECT 18.27 3.945 18.44 4.115 ;
      RECT 17.81 -1.495 17.98 -1.325 ;
      RECT 17.81 1.225 17.98 1.395 ;
      RECT 17.81 3.945 17.98 4.115 ;
      RECT 17.55 3.655 17.72 3.825 ;
      RECT 17.37 2.755 17.54 2.925 ;
      RECT 17.35 -1.495 17.52 -1.325 ;
      RECT 17.35 1.225 17.52 1.395 ;
      RECT 17.35 3.945 17.52 4.115 ;
      RECT 17.03 -0.645 17.2 -0.475 ;
      RECT 16.89 -1.495 17.06 -1.325 ;
      RECT 16.89 1.225 17.06 1.395 ;
      RECT 16.89 3.945 17.06 4.115 ;
      RECT 16.86 0.715 17.03 0.885 ;
      RECT 16.43 -1.495 16.6 -1.325 ;
      RECT 16.43 1.225 16.6 1.395 ;
      RECT 16.43 3.945 16.6 4.115 ;
      RECT 16.35 2.755 16.52 2.925 ;
      RECT 15.97 -1.495 16.14 -1.325 ;
      RECT 15.97 1.225 16.14 1.395 ;
      RECT 15.97 3.945 16.14 4.115 ;
      RECT 15.67 1.735 15.84 1.905 ;
      RECT 15.51 -1.495 15.68 -1.325 ;
      RECT 15.51 1.225 15.68 1.395 ;
      RECT 15.51 3.945 15.68 4.115 ;
      RECT 15.05 -1.495 15.22 -1.325 ;
      RECT 15.05 1.225 15.22 1.395 ;
      RECT 15.05 3.945 15.22 4.115 ;
      RECT 14.995 -0.305 15.165 -0.135 ;
      RECT 14.65 2.775 14.82 2.945 ;
      RECT 14.59 1.225 14.76 1.395 ;
      RECT 14.59 3.945 14.76 4.115 ;
      RECT 14.13 1.225 14.3 1.395 ;
      RECT 14.13 3.945 14.3 4.115 ;
      RECT 13.67 1.225 13.84 1.395 ;
      RECT 13.67 3.945 13.84 4.115 ;
      RECT 13.21 1.225 13.38 1.395 ;
      RECT 13.21 3.945 13.38 4.115 ;
      RECT 13.12 2.27 13.29 2.44 ;
      RECT 12.75 1.225 12.92 1.395 ;
      RECT 12.75 3.945 12.92 4.115 ;
      RECT 12.29 1.225 12.46 1.395 ;
      RECT 12.29 3.945 12.46 4.115 ;
      RECT 11.83 1.225 12 1.395 ;
      RECT 11.83 3.945 12 4.115 ;
      RECT 11.44 2.4 11.61 2.57 ;
      RECT 11.37 1.225 11.54 1.395 ;
      RECT 11.37 3.945 11.54 4.115 ;
      RECT 10.91 1.225 11.08 1.395 ;
      RECT 10.91 3.945 11.08 4.115 ;
      RECT -0.125 2.935 0.045 3.105 ;
      RECT -0.125 5.655 0.045 5.825 ;
      RECT -0.585 2.935 -0.415 3.105 ;
      RECT -0.585 5.655 -0.415 5.825 ;
      RECT -1.045 2.935 -0.875 3.105 ;
      RECT -1.045 5.655 -0.875 5.825 ;
      RECT -1.495 4.11 -1.325 4.28 ;
      RECT -1.505 2.935 -1.335 3.105 ;
      RECT -1.505 5.655 -1.335 5.825 ;
      RECT -1.855 4.675 -1.685 4.845 ;
      RECT -1.965 2.935 -1.795 3.105 ;
      RECT -1.965 5.655 -1.795 5.825 ;
      RECT -2.425 2.935 -2.255 3.105 ;
      RECT -2.425 5.655 -2.255 5.825 ;
      RECT -2.885 2.935 -2.715 3.105 ;
      RECT -2.885 5.655 -2.715 5.825 ;
      RECT -3.345 2.935 -3.175 3.105 ;
      RECT -3.345 5.655 -3.175 5.825 ;
      RECT -3.775 3.655 -3.605 3.825 ;
      RECT -3.805 2.935 -3.635 3.105 ;
      RECT -3.805 5.655 -3.635 5.825 ;
    LAYER li ;
      RECT 99.4 -1.495 99.63 -0.505 ;
      RECT 98.02 -1.495 98.25 -0.505 ;
      RECT 86.745 -1.495 87.005 -0.505 ;
      RECT 81.46 -1.495 81.69 -0.505 ;
      RECT 80.08 -1.495 80.31 -0.505 ;
      RECT 68.805 -1.495 69.065 -0.505 ;
      RECT 63.525 -1.495 63.755 -0.505 ;
      RECT 62.145 -1.495 62.375 -0.505 ;
      RECT 50.87 -1.495 51.13 -0.505 ;
      RECT 45.585 -1.495 45.815 -0.505 ;
      RECT 44.205 -1.495 44.435 -0.505 ;
      RECT 32.93 -1.495 33.19 -0.505 ;
      RECT 27.645 -1.495 27.875 -0.505 ;
      RECT 26.265 -1.495 26.495 -0.505 ;
      RECT 14.99 -1.495 15.25 -0.505 ;
      RECT 93.195 -1.495 93.465 -0.515 ;
      RECT 92.285 -1.495 92.525 -0.515 ;
      RECT 75.255 -1.495 75.525 -0.515 ;
      RECT 74.345 -1.495 74.585 -0.515 ;
      RECT 57.32 -1.495 57.59 -0.515 ;
      RECT 56.41 -1.495 56.65 -0.515 ;
      RECT 39.38 -1.495 39.65 -0.515 ;
      RECT 38.47 -1.495 38.71 -0.515 ;
      RECT 21.44 -1.495 21.71 -0.515 ;
      RECT 20.53 -1.495 20.77 -0.515 ;
      RECT 91.415 -1.495 91.665 -0.785 ;
      RECT 73.475 -1.495 73.725 -0.785 ;
      RECT 55.54 -1.495 55.79 -0.785 ;
      RECT 37.6 -1.495 37.85 -0.785 ;
      RECT 19.66 -1.495 19.91 -0.785 ;
      RECT 96.365 -1.495 96.875 -0.79 ;
      RECT 78.425 -1.495 78.935 -0.79 ;
      RECT 60.49 -1.495 61 -0.79 ;
      RECT 42.55 -1.495 43.06 -0.79 ;
      RECT 24.61 -1.495 25.12 -0.79 ;
      RECT 89.035 -1.495 89.365 -0.865 ;
      RECT 71.095 -1.495 71.425 -0.865 ;
      RECT 53.16 -1.495 53.49 -0.865 ;
      RECT 35.22 -1.495 35.55 -0.865 ;
      RECT 17.28 -1.495 17.61 -0.865 ;
      RECT 94.075 -1.495 94.405 -0.925 ;
      RECT 76.135 -1.495 76.465 -0.925 ;
      RECT 58.2 -1.495 58.53 -0.925 ;
      RECT 40.26 -1.495 40.59 -0.925 ;
      RECT 22.32 -1.495 22.65 -0.925 ;
      RECT 10.765 -1.495 100.46 -1.325 ;
      RECT 99.42 0.085 99.63 2.535 ;
      RECT 98.04 0.085 98.25 2.535 ;
      RECT 94.155 0.085 94.325 2.535 ;
      RECT 85.895 1.225 86.065 2.535 ;
      RECT 81.48 0.085 81.69 2.535 ;
      RECT 80.1 0.085 80.31 2.535 ;
      RECT 76.215 0.085 76.385 2.535 ;
      RECT 67.955 1.225 68.125 2.535 ;
      RECT 63.545 0.085 63.755 2.535 ;
      RECT 62.165 0.085 62.375 2.535 ;
      RECT 58.28 0.085 58.45 2.535 ;
      RECT 50.02 1.225 50.19 2.535 ;
      RECT 45.605 0.085 45.815 2.535 ;
      RECT 44.225 0.085 44.435 2.535 ;
      RECT 40.34 0.085 40.51 2.535 ;
      RECT 32.08 1.225 32.25 2.535 ;
      RECT 27.665 0.085 27.875 2.535 ;
      RECT 26.285 0.085 26.495 2.535 ;
      RECT 22.4 0.085 22.57 2.535 ;
      RECT 14.14 1.225 14.31 2.535 ;
      RECT 90.015 0.57 90.28 2.175 ;
      RECT 72.075 0.57 72.34 2.175 ;
      RECT 54.14 0.57 54.405 2.175 ;
      RECT 36.2 0.57 36.465 2.175 ;
      RECT 18.26 0.57 18.525 2.175 ;
      RECT 96.695 0.465 96.865 2.155 ;
      RECT 83.355 1.225 83.525 2.155 ;
      RECT 78.755 0.465 78.925 2.155 ;
      RECT 65.415 1.225 65.585 2.155 ;
      RECT 60.82 0.465 60.99 2.155 ;
      RECT 47.48 1.225 47.65 2.155 ;
      RECT 42.88 0.465 43.05 2.155 ;
      RECT 29.54 1.225 29.71 2.155 ;
      RECT 24.94 0.465 25.11 2.155 ;
      RECT 11.6 1.225 11.77 2.155 ;
      RECT 87.855 0.72 88.185 2.115 ;
      RECT 69.915 0.72 70.245 2.115 ;
      RECT 51.98 0.72 52.31 2.115 ;
      RECT 34.04 0.72 34.37 2.115 ;
      RECT 16.1 0.72 16.43 2.115 ;
      RECT 88.855 1.225 89.135 2.065 ;
      RECT 70.915 1.225 71.195 2.065 ;
      RECT 52.98 1.225 53.26 2.065 ;
      RECT 35.04 1.225 35.32 2.065 ;
      RECT 17.1 1.225 17.38 2.065 ;
      RECT 89.325 1.125 89.555 1.875 ;
      RECT 71.385 1.125 71.615 1.875 ;
      RECT 53.45 1.125 53.68 1.875 ;
      RECT 35.51 1.125 35.74 1.875 ;
      RECT 17.57 1.125 17.8 1.875 ;
      RECT 90.83 1.225 91.205 1.775 ;
      RECT 72.89 1.225 73.265 1.775 ;
      RECT 54.955 1.225 55.33 1.775 ;
      RECT 37.015 1.225 37.39 1.775 ;
      RECT 19.075 1.225 19.45 1.775 ;
      RECT 10.765 1.225 100.46 1.395 ;
      RECT 93.135 0.085 93.465 1.395 ;
      RECT 91.395 0.68 91.65 1.395 ;
      RECT 89.965 0.57 90.57 1.395 ;
      RECT 89.095 0.68 89.31 1.395 ;
      RECT 87.665 0.72 88.28 1.395 ;
      RECT 88.085 0.355 88.28 1.395 ;
      RECT 86.745 0.715 87.005 1.395 ;
      RECT 75.195 0.085 75.525 1.395 ;
      RECT 73.455 0.68 73.71 1.395 ;
      RECT 72.025 0.57 72.63 1.395 ;
      RECT 71.155 0.68 71.37 1.395 ;
      RECT 69.725 0.72 70.34 1.395 ;
      RECT 70.145 0.355 70.34 1.395 ;
      RECT 68.805 0.715 69.065 1.395 ;
      RECT 57.26 0.085 57.59 1.395 ;
      RECT 55.52 0.68 55.775 1.395 ;
      RECT 54.09 0.57 54.695 1.395 ;
      RECT 53.22 0.68 53.435 1.395 ;
      RECT 51.79 0.72 52.405 1.395 ;
      RECT 52.21 0.355 52.405 1.395 ;
      RECT 50.87 0.715 51.13 1.395 ;
      RECT 39.32 0.085 39.65 1.395 ;
      RECT 37.58 0.68 37.835 1.395 ;
      RECT 36.15 0.57 36.755 1.395 ;
      RECT 35.28 0.68 35.495 1.395 ;
      RECT 33.85 0.72 34.465 1.395 ;
      RECT 34.27 0.355 34.465 1.395 ;
      RECT 32.93 0.715 33.19 1.395 ;
      RECT 21.38 0.085 21.71 1.395 ;
      RECT 19.64 0.68 19.895 1.395 ;
      RECT 18.21 0.57 18.815 1.395 ;
      RECT 17.34 0.68 17.555 1.395 ;
      RECT 15.91 0.72 16.525 1.395 ;
      RECT 16.33 0.355 16.525 1.395 ;
      RECT 14.99 0.715 15.25 1.395 ;
      RECT 90.395 0.3 90.58 0.67 ;
      RECT 72.455 0.3 72.64 0.67 ;
      RECT 54.52 0.3 54.705 0.67 ;
      RECT 36.58 0.3 36.765 0.67 ;
      RECT 18.64 0.3 18.825 0.67 ;
      RECT 90.395 0.3 90.725 0.545 ;
      RECT 88.085 0.355 88.415 0.545 ;
      RECT 72.455 0.3 72.785 0.545 ;
      RECT 70.145 0.355 70.475 0.545 ;
      RECT 54.52 0.3 54.85 0.545 ;
      RECT 52.21 0.355 52.54 0.545 ;
      RECT 36.58 0.3 36.91 0.545 ;
      RECT 34.27 0.355 34.6 0.545 ;
      RECT 18.64 0.3 18.97 0.545 ;
      RECT 16.33 0.355 16.66 0.545 ;
      RECT 72.62 3.945 72.79 4.28 ;
      RECT 54.68 3.945 54.85 4.28 ;
      RECT 36.745 3.945 36.915 4.28 ;
      RECT 18.805 3.945 18.975 4.28 ;
      RECT 10.765 3.945 100.46 4.115 ;
      RECT 99.4 3.125 99.63 4.115 ;
      RECT 98.02 3.125 98.25 4.115 ;
      RECT 96.365 3.41 96.875 4.115 ;
      RECT 94.075 3.545 94.405 4.115 ;
      RECT 92.095 3.435 92.545 4.115 ;
      RECT 90.005 3.545 90.335 4.115 ;
      RECT 87.935 3.485 88.185 4.115 ;
      RECT 85.815 3.545 86.145 4.115 ;
      RECT 84.395 2.615 84.67 4.115 ;
      RECT 83.345 3.41 83.855 4.115 ;
      RECT 81.46 3.125 81.69 4.115 ;
      RECT 80.08 3.125 80.31 4.115 ;
      RECT 78.425 3.41 78.935 4.115 ;
      RECT 76.135 3.545 76.465 4.115 ;
      RECT 74.155 3.435 74.605 4.115 ;
      RECT 72.065 3.545 72.395 4.115 ;
      RECT 69.995 3.485 70.245 4.115 ;
      RECT 67.875 3.545 68.205 4.115 ;
      RECT 66.455 2.615 66.73 4.115 ;
      RECT 65.405 3.41 65.915 4.115 ;
      RECT 63.525 3.125 63.755 4.115 ;
      RECT 62.145 3.125 62.375 4.115 ;
      RECT 60.49 3.41 61 4.115 ;
      RECT 58.2 3.545 58.53 4.115 ;
      RECT 56.22 3.435 56.67 4.115 ;
      RECT 54.13 3.545 54.46 4.115 ;
      RECT 52.06 3.485 52.31 4.115 ;
      RECT 49.94 3.545 50.27 4.115 ;
      RECT 48.52 2.615 48.795 4.115 ;
      RECT 47.47 3.41 47.98 4.115 ;
      RECT 45.585 3.125 45.815 4.115 ;
      RECT 44.205 3.125 44.435 4.115 ;
      RECT 42.55 3.41 43.06 4.115 ;
      RECT 40.26 3.545 40.59 4.115 ;
      RECT 38.28 3.435 38.73 4.115 ;
      RECT 36.19 3.545 36.52 4.115 ;
      RECT 34.12 3.485 34.37 4.115 ;
      RECT 32 3.545 32.33 4.115 ;
      RECT 30.58 2.615 30.855 4.115 ;
      RECT 29.53 3.41 30.04 4.115 ;
      RECT 27.645 3.125 27.875 4.115 ;
      RECT 26.265 3.125 26.495 4.115 ;
      RECT 24.61 3.41 25.12 4.115 ;
      RECT 22.32 3.545 22.65 4.115 ;
      RECT 20.34 3.435 20.79 4.115 ;
      RECT 18.25 3.545 18.58 4.115 ;
      RECT 16.18 3.485 16.43 4.115 ;
      RECT 14.06 3.545 14.39 4.115 ;
      RECT 12.64 2.615 12.915 4.115 ;
      RECT 11.59 3.41 12.1 4.115 ;
      RECT 99.8 0.075 100.13 1.055 ;
      RECT 99.9 -1.155 100.13 1.055 ;
      RECT 99.8 -1.155 100.13 -0.525 ;
      RECT 99.8 3.145 100.13 3.775 ;
      RECT 99.9 1.565 100.13 3.775 ;
      RECT 99.8 1.565 100.13 2.545 ;
      RECT 98.42 0.075 98.75 1.055 ;
      RECT 98.52 -1.155 98.75 1.055 ;
      RECT 99.4 -0.335 99.73 -0.095 ;
      RECT 98.52 -0.305 99.73 -0.135 ;
      RECT 98.42 -1.155 98.75 -0.525 ;
      RECT 98.42 3.145 98.75 3.775 ;
      RECT 98.52 1.565 98.75 3.775 ;
      RECT 99.4 2.715 99.73 2.955 ;
      RECT 98.52 2.72 99.73 2.89 ;
      RECT 98.42 1.565 98.75 2.545 ;
      RECT 97.1 0.465 97.615 0.875 ;
      RECT 97.275 -0.515 97.615 0.875 ;
      RECT 96.385 -0.515 97.615 -0.345 ;
      RECT 97.095 -1.12 97.34 -0.345 ;
      RECT 97.095 2.965 97.34 3.74 ;
      RECT 96.385 2.965 97.615 3.135 ;
      RECT 97.275 1.745 97.615 3.135 ;
      RECT 97.1 1.745 97.615 2.155 ;
      RECT 94.495 0.885 96.525 1.055 ;
      RECT 96.355 0.03 96.525 1.055 ;
      RECT 94.495 -0.415 94.665 1.055 ;
      RECT 96.355 0.03 97.105 0.22 ;
      RECT 94.47 -0.415 94.665 -0.085 ;
      RECT 94.47 2.705 94.665 3.035 ;
      RECT 94.495 1.565 94.665 3.035 ;
      RECT 96.355 2.4 97.105 2.59 ;
      RECT 96.355 1.565 96.525 2.59 ;
      RECT 94.495 1.565 96.525 1.735 ;
      RECT 95.175 0.205 96.185 0.375 ;
      RECT 95.995 -1.155 96.185 0.375 ;
      RECT 95.175 -0.595 95.345 0.375 ;
      RECT 95.995 2.245 96.185 3.775 ;
      RECT 95.175 2.245 95.345 3.215 ;
      RECT 95.175 2.245 96.185 2.415 ;
      RECT 94.835 0.545 95.96 0.715 ;
      RECT 94.835 -1.155 95.005 0.715 ;
      RECT 93.99 -0.415 94.245 -0.085 ;
      RECT 94.075 -0.755 94.245 -0.085 ;
      RECT 94.075 -0.755 95.005 -0.585 ;
      RECT 94.83 -1.155 95.005 -0.585 ;
      RECT 94.83 -1.155 95.36 -0.79 ;
      RECT 94.83 3.41 95.36 3.775 ;
      RECT 94.83 3.205 95.005 3.775 ;
      RECT 94.835 1.905 95.005 3.775 ;
      RECT 94.075 3.205 95.005 3.375 ;
      RECT 94.075 2.705 94.245 3.375 ;
      RECT 93.99 2.705 94.245 3.035 ;
      RECT 94.835 1.905 95.96 2.075 ;
      RECT 93.65 0.085 93.985 1.055 ;
      RECT 93.65 -1.155 93.82 1.055 ;
      RECT 93.65 -1.155 93.905 -0.585 ;
      RECT 93.65 3.205 93.905 3.775 ;
      RECT 93.65 1.565 93.82 3.775 ;
      RECT 93.65 1.565 93.985 2.535 ;
      RECT 90.515 3.525 91.82 3.775 ;
      RECT 90.515 3.205 90.695 3.775 ;
      RECT 89.965 3.205 90.695 3.375 ;
      RECT 89.965 2.365 90.135 3.375 ;
      RECT 90.8 2.405 92.545 2.585 ;
      RECT 92.215 1.565 92.545 2.585 ;
      RECT 89.965 2.365 91.025 2.535 ;
      RECT 92.215 1.735 93.035 1.905 ;
      RECT 91.375 1.565 91.705 1.775 ;
      RECT 91.375 1.565 92.545 1.735 ;
      RECT 92.275 0.085 92.605 1.04 ;
      RECT 92.275 0.085 92.955 0.255 ;
      RECT 92.785 -1.155 92.955 0.255 ;
      RECT 92.695 -1.155 93.025 -0.515 ;
      RECT 91.82 0.355 92.095 1.055 ;
      RECT 91.925 -1.155 92.095 1.055 ;
      RECT 92.265 -0.335 92.615 -0.085 ;
      RECT 91.925 -0.305 92.615 -0.135 ;
      RECT 91.835 -1.155 92.095 -0.675 ;
      RECT 91.165 1.995 92.045 2.235 ;
      RECT 91.815 1.905 92.045 2.235 ;
      RECT 90.515 1.995 92.045 2.195 ;
      RECT 91.43 1.945 92.045 2.235 ;
      RECT 90.515 1.865 90.685 2.195 ;
      RECT 91.4 2.755 91.65 3.355 ;
      RECT 91.4 2.755 91.875 2.955 ;
      RECT 90.895 -0.025 91.65 0.475 ;
      RECT 89.965 -0.22 90.225 0.4 ;
      RECT 90.88 -0.08 90.895 0.225 ;
      RECT 90.865 -0.095 90.885 0.19 ;
      RECT 91.525 -0.42 91.755 0.18 ;
      RECT 90.84 -0.15 90.86 0.165 ;
      RECT 90.82 -0.025 91.755 0.15 ;
      RECT 90.795 -0.025 91.755 0.14 ;
      RECT 90.725 -0.025 91.755 0.13 ;
      RECT 90.705 -0.025 91.755 0.1 ;
      RECT 90.685 -1.115 90.855 0.07 ;
      RECT 90.655 -0.025 91.755 0.04 ;
      RECT 90.62 -0.025 91.755 0.015 ;
      RECT 90.59 -0.03 90.98 -0.02 ;
      RECT 90.59 -0.04 90.955 -0.02 ;
      RECT 90.59 -0.045 90.94 -0.02 ;
      RECT 90.59 -0.055 90.925 -0.02 ;
      RECT 89.965 -0.22 90.855 -0.05 ;
      RECT 89.965 -0.065 90.915 -0.05 ;
      RECT 89.965 -0.07 90.905 -0.05 ;
      RECT 90.86 -0.125 90.87 0.18 ;
      RECT 89.965 -0.09 90.89 -0.05 ;
      RECT 89.965 -0.11 90.875 -0.05 ;
      RECT 89.965 -1.115 90.855 -0.945 ;
      RECT 91.025 -0.62 91.355 -0.195 ;
      RECT 91.025 -1.105 91.245 -0.195 ;
      RECT 90.94 2.755 91.15 3.355 ;
      RECT 90.8 2.755 91.15 2.955 ;
      RECT 89.52 0.355 89.795 1.055 ;
      RECT 89.74 -1.155 89.795 1.055 ;
      RECT 89.625 -0.35 89.795 1.055 ;
      RECT 89.625 -1.155 89.795 -0.355 ;
      RECT 89.535 -1.155 89.795 -0.68 ;
      RECT 87.665 0.015 87.915 0.55 ;
      RECT 88.635 0.015 89.35 0.48 ;
      RECT 87.665 0.015 89.455 0.185 ;
      RECT 89.225 -0.35 89.455 0.185 ;
      RECT 88.22 -1.105 88.475 0.185 ;
      RECT 89.225 -0.415 89.285 0.48 ;
      RECT 89.285 -0.42 89.455 -0.355 ;
      RECT 87.685 -1.105 88.475 -0.84 ;
      RECT 88.645 2.705 89.32 2.955 ;
      RECT 89.055 2.345 89.32 2.955 ;
      RECT 88.805 3.125 89.135 3.675 ;
      RECT 87.745 3.125 89.135 3.315 ;
      RECT 87.745 2.285 87.915 3.315 ;
      RECT 87.625 2.705 87.915 3.035 ;
      RECT 87.745 2.285 88.685 2.455 ;
      RECT 88.385 1.735 88.685 2.455 ;
      RECT 88.645 -0.685 89.055 -0.165 ;
      RECT 88.645 -1.105 88.845 -0.165 ;
      RECT 87.255 -0.925 87.425 1.055 ;
      RECT 87.255 -0.415 88.05 -0.165 ;
      RECT 87.255 -0.925 87.505 -0.165 ;
      RECT 87.175 -0.925 87.505 -0.505 ;
      RECT 87.205 3.485 87.765 3.775 ;
      RECT 87.205 1.565 87.455 3.775 ;
      RECT 87.205 1.565 87.665 2.115 ;
      RECT 86.315 3.205 86.57 3.775 ;
      RECT 86.4 1.565 86.57 3.775 ;
      RECT 86.4 2.775 86.575 2.945 ;
      RECT 86.235 1.565 86.57 2.535 ;
      RECT 84.86 3.41 85.39 3.775 ;
      RECT 85.215 3.205 85.39 3.775 ;
      RECT 85.215 3.205 86.145 3.375 ;
      RECT 85.975 2.705 86.145 3.375 ;
      RECT 85.215 1.905 85.385 3.775 ;
      RECT 85.975 2.705 86.23 3.035 ;
      RECT 84.26 1.905 85.385 2.075 ;
      RECT 85.555 2.705 85.75 3.035 ;
      RECT 85.555 1.565 85.725 3.035 ;
      RECT 83.115 2.4 83.865 2.59 ;
      RECT 83.695 1.565 83.865 2.59 ;
      RECT 83.695 1.565 85.725 1.735 ;
      RECT 84.035 2.245 84.225 3.775 ;
      RECT 84.875 2.245 85.045 3.215 ;
      RECT 84.87 2.245 85.045 2.5 ;
      RECT 84.035 2.245 85.045 2.415 ;
      RECT 82.88 2.965 83.125 3.74 ;
      RECT 82.605 2.965 83.835 3.135 ;
      RECT 82.605 1.745 82.945 3.135 ;
      RECT 82.605 1.745 83.12 2.155 ;
      RECT 81.86 0.075 82.19 1.055 ;
      RECT 81.96 -1.155 82.19 1.055 ;
      RECT 81.86 -1.155 82.19 -0.525 ;
      RECT 81.86 3.145 82.19 3.775 ;
      RECT 81.96 1.565 82.19 3.775 ;
      RECT 81.86 1.565 82.19 2.545 ;
      RECT 80.48 0.075 80.81 1.055 ;
      RECT 80.58 -1.155 80.81 1.055 ;
      RECT 81.46 -0.335 81.79 -0.095 ;
      RECT 80.58 -0.305 81.79 -0.135 ;
      RECT 80.48 -1.155 80.81 -0.525 ;
      RECT 80.48 3.145 80.81 3.775 ;
      RECT 80.58 1.565 80.81 3.775 ;
      RECT 81.46 2.715 81.79 2.955 ;
      RECT 80.58 2.72 81.79 2.89 ;
      RECT 80.48 1.565 80.81 2.545 ;
      RECT 79.16 0.465 79.675 0.875 ;
      RECT 79.335 -0.515 79.675 0.875 ;
      RECT 78.445 -0.515 79.675 -0.345 ;
      RECT 79.155 -1.12 79.4 -0.345 ;
      RECT 79.155 2.965 79.4 3.74 ;
      RECT 78.445 2.965 79.675 3.135 ;
      RECT 79.335 1.745 79.675 3.135 ;
      RECT 79.16 1.745 79.675 2.155 ;
      RECT 76.555 0.885 78.585 1.055 ;
      RECT 78.415 0.03 78.585 1.055 ;
      RECT 76.555 -0.415 76.725 1.055 ;
      RECT 78.415 0.03 79.165 0.22 ;
      RECT 76.53 -0.415 76.725 -0.085 ;
      RECT 76.53 2.705 76.725 3.035 ;
      RECT 76.555 1.565 76.725 3.035 ;
      RECT 78.415 2.4 79.165 2.59 ;
      RECT 78.415 1.565 78.585 2.59 ;
      RECT 76.555 1.565 78.585 1.735 ;
      RECT 77.235 0.205 78.245 0.375 ;
      RECT 78.055 -1.155 78.245 0.375 ;
      RECT 77.235 -0.595 77.405 0.375 ;
      RECT 78.055 2.245 78.245 3.775 ;
      RECT 77.235 2.245 77.405 3.215 ;
      RECT 77.235 2.245 78.245 2.415 ;
      RECT 76.895 0.545 78.02 0.715 ;
      RECT 76.895 -1.155 77.065 0.715 ;
      RECT 76.05 -0.415 76.305 -0.085 ;
      RECT 76.135 -0.755 76.305 -0.085 ;
      RECT 76.135 -0.755 77.065 -0.585 ;
      RECT 76.89 -1.155 77.065 -0.585 ;
      RECT 76.89 -1.155 77.42 -0.79 ;
      RECT 76.89 3.41 77.42 3.775 ;
      RECT 76.89 3.205 77.065 3.775 ;
      RECT 76.895 1.905 77.065 3.775 ;
      RECT 76.135 3.205 77.065 3.375 ;
      RECT 76.135 2.705 76.305 3.375 ;
      RECT 76.05 2.705 76.305 3.035 ;
      RECT 76.895 1.905 78.02 2.075 ;
      RECT 75.71 0.085 76.045 1.055 ;
      RECT 75.71 -1.155 75.88 1.055 ;
      RECT 75.71 -1.155 75.965 -0.585 ;
      RECT 75.71 3.205 75.965 3.775 ;
      RECT 75.71 1.565 75.88 3.775 ;
      RECT 75.71 1.565 76.045 2.535 ;
      RECT 72.575 3.525 73.88 3.775 ;
      RECT 72.575 3.205 72.755 3.775 ;
      RECT 72.025 3.205 72.755 3.375 ;
      RECT 72.025 2.365 72.195 3.375 ;
      RECT 72.86 2.405 74.605 2.585 ;
      RECT 74.275 1.565 74.605 2.585 ;
      RECT 72.025 2.365 73.085 2.535 ;
      RECT 74.275 1.735 75.095 1.905 ;
      RECT 73.435 1.565 73.765 1.775 ;
      RECT 73.435 1.565 74.605 1.735 ;
      RECT 74.335 0.085 74.665 1.04 ;
      RECT 74.335 0.085 75.015 0.255 ;
      RECT 74.845 -1.155 75.015 0.255 ;
      RECT 74.755 -1.155 75.085 -0.515 ;
      RECT 73.88 0.355 74.155 1.055 ;
      RECT 73.985 -1.155 74.155 1.055 ;
      RECT 74.325 -0.335 74.675 -0.085 ;
      RECT 73.985 -0.305 74.675 -0.135 ;
      RECT 73.895 -1.155 74.155 -0.675 ;
      RECT 73.225 1.995 74.105 2.235 ;
      RECT 73.875 1.905 74.105 2.235 ;
      RECT 72.575 1.995 74.105 2.195 ;
      RECT 73.49 1.945 74.105 2.235 ;
      RECT 72.575 1.865 72.745 2.195 ;
      RECT 73.46 2.755 73.71 3.355 ;
      RECT 73.46 2.755 73.935 2.955 ;
      RECT 72.955 -0.025 73.71 0.475 ;
      RECT 72.025 -0.22 72.285 0.4 ;
      RECT 72.94 -0.08 72.955 0.225 ;
      RECT 72.925 -0.095 72.945 0.19 ;
      RECT 73.585 -0.42 73.815 0.18 ;
      RECT 72.9 -0.15 72.92 0.165 ;
      RECT 72.88 -0.025 73.815 0.15 ;
      RECT 72.855 -0.025 73.815 0.14 ;
      RECT 72.785 -0.025 73.815 0.13 ;
      RECT 72.765 -0.025 73.815 0.1 ;
      RECT 72.745 -1.115 72.915 0.07 ;
      RECT 72.715 -0.025 73.815 0.04 ;
      RECT 72.68 -0.025 73.815 0.015 ;
      RECT 72.65 -0.03 73.04 -0.02 ;
      RECT 72.65 -0.04 73.015 -0.02 ;
      RECT 72.65 -0.045 73 -0.02 ;
      RECT 72.65 -0.055 72.985 -0.02 ;
      RECT 72.025 -0.22 72.915 -0.05 ;
      RECT 72.025 -0.065 72.975 -0.05 ;
      RECT 72.025 -0.07 72.965 -0.05 ;
      RECT 72.92 -0.125 72.93 0.18 ;
      RECT 72.025 -0.09 72.95 -0.05 ;
      RECT 72.025 -0.11 72.935 -0.05 ;
      RECT 72.025 -1.115 72.915 -0.945 ;
      RECT 73.085 -0.62 73.415 -0.195 ;
      RECT 73.085 -1.105 73.305 -0.195 ;
      RECT 73 2.755 73.21 3.355 ;
      RECT 72.86 2.755 73.21 2.955 ;
      RECT 71.58 0.355 71.855 1.055 ;
      RECT 71.8 -1.155 71.855 1.055 ;
      RECT 71.685 -0.35 71.855 1.055 ;
      RECT 71.685 -1.155 71.855 -0.355 ;
      RECT 71.595 -1.155 71.855 -0.68 ;
      RECT 69.725 0.015 69.975 0.55 ;
      RECT 70.695 0.015 71.41 0.48 ;
      RECT 69.725 0.015 71.515 0.185 ;
      RECT 71.285 -0.35 71.515 0.185 ;
      RECT 70.28 -1.105 70.535 0.185 ;
      RECT 71.285 -0.415 71.345 0.48 ;
      RECT 71.345 -0.42 71.515 -0.355 ;
      RECT 69.745 -1.105 70.535 -0.84 ;
      RECT 70.705 2.705 71.38 2.955 ;
      RECT 71.115 2.345 71.38 2.955 ;
      RECT 70.865 3.125 71.195 3.675 ;
      RECT 69.805 3.125 71.195 3.315 ;
      RECT 69.805 2.285 69.975 3.315 ;
      RECT 69.685 2.705 69.975 3.035 ;
      RECT 69.805 2.285 70.745 2.455 ;
      RECT 70.445 1.735 70.745 2.455 ;
      RECT 70.705 -0.685 71.115 -0.165 ;
      RECT 70.705 -1.105 70.905 -0.165 ;
      RECT 69.315 -0.925 69.485 1.055 ;
      RECT 69.315 -0.415 70.11 -0.165 ;
      RECT 69.315 -0.925 69.565 -0.165 ;
      RECT 69.235 -0.925 69.565 -0.505 ;
      RECT 69.265 3.485 69.825 3.775 ;
      RECT 69.265 1.565 69.515 3.775 ;
      RECT 69.265 1.565 69.725 2.115 ;
      RECT 68.375 3.205 68.63 3.775 ;
      RECT 68.46 1.565 68.63 3.775 ;
      RECT 68.46 2.775 68.635 2.945 ;
      RECT 68.295 1.565 68.63 2.535 ;
      RECT 66.92 3.41 67.45 3.775 ;
      RECT 67.275 3.205 67.45 3.775 ;
      RECT 67.275 3.205 68.205 3.375 ;
      RECT 68.035 2.705 68.205 3.375 ;
      RECT 67.275 1.905 67.445 3.775 ;
      RECT 68.035 2.705 68.29 3.035 ;
      RECT 66.32 1.905 67.445 2.075 ;
      RECT 67.615 2.705 67.81 3.035 ;
      RECT 67.615 1.565 67.785 3.035 ;
      RECT 65.175 2.4 65.925 2.59 ;
      RECT 65.755 1.565 65.925 2.59 ;
      RECT 65.755 1.565 67.785 1.735 ;
      RECT 66.095 2.245 66.285 3.775 ;
      RECT 66.935 2.245 67.105 3.215 ;
      RECT 66.93 2.245 67.105 2.5 ;
      RECT 66.095 2.245 67.105 2.415 ;
      RECT 64.94 2.965 65.185 3.74 ;
      RECT 64.665 2.965 65.895 3.135 ;
      RECT 64.665 1.745 65.005 3.135 ;
      RECT 64.665 1.745 65.18 2.155 ;
      RECT 63.925 0.075 64.255 1.055 ;
      RECT 64.025 -1.155 64.255 1.055 ;
      RECT 63.925 -1.155 64.255 -0.525 ;
      RECT 63.925 3.145 64.255 3.775 ;
      RECT 64.025 1.565 64.255 3.775 ;
      RECT 63.925 1.565 64.255 2.545 ;
      RECT 62.545 0.075 62.875 1.055 ;
      RECT 62.645 -1.155 62.875 1.055 ;
      RECT 63.525 -0.335 63.855 -0.095 ;
      RECT 62.645 -0.305 63.855 -0.135 ;
      RECT 62.545 -1.155 62.875 -0.525 ;
      RECT 62.545 3.145 62.875 3.775 ;
      RECT 62.645 1.565 62.875 3.775 ;
      RECT 63.525 2.715 63.855 2.955 ;
      RECT 62.645 2.72 63.855 2.89 ;
      RECT 62.545 1.565 62.875 2.545 ;
      RECT 61.225 0.465 61.74 0.875 ;
      RECT 61.4 -0.515 61.74 0.875 ;
      RECT 60.51 -0.515 61.74 -0.345 ;
      RECT 61.22 -1.12 61.465 -0.345 ;
      RECT 61.22 2.965 61.465 3.74 ;
      RECT 60.51 2.965 61.74 3.135 ;
      RECT 61.4 1.745 61.74 3.135 ;
      RECT 61.225 1.745 61.74 2.155 ;
      RECT 58.62 0.885 60.65 1.055 ;
      RECT 60.48 0.03 60.65 1.055 ;
      RECT 58.62 -0.415 58.79 1.055 ;
      RECT 60.48 0.03 61.23 0.22 ;
      RECT 58.595 -0.415 58.79 -0.085 ;
      RECT 58.595 2.705 58.79 3.035 ;
      RECT 58.62 1.565 58.79 3.035 ;
      RECT 60.48 2.4 61.23 2.59 ;
      RECT 60.48 1.565 60.65 2.59 ;
      RECT 58.62 1.565 60.65 1.735 ;
      RECT 59.3 0.205 60.31 0.375 ;
      RECT 60.12 -1.155 60.31 0.375 ;
      RECT 59.3 -0.595 59.47 0.375 ;
      RECT 60.12 2.245 60.31 3.775 ;
      RECT 59.3 2.245 59.47 3.215 ;
      RECT 59.3 2.245 60.31 2.415 ;
      RECT 58.96 0.545 60.085 0.715 ;
      RECT 58.96 -1.155 59.13 0.715 ;
      RECT 58.115 -0.415 58.37 -0.085 ;
      RECT 58.2 -0.755 58.37 -0.085 ;
      RECT 58.2 -0.755 59.13 -0.585 ;
      RECT 58.955 -1.155 59.13 -0.585 ;
      RECT 58.955 -1.155 59.485 -0.79 ;
      RECT 58.955 3.41 59.485 3.775 ;
      RECT 58.955 3.205 59.13 3.775 ;
      RECT 58.96 1.905 59.13 3.775 ;
      RECT 58.2 3.205 59.13 3.375 ;
      RECT 58.2 2.705 58.37 3.375 ;
      RECT 58.115 2.705 58.37 3.035 ;
      RECT 58.96 1.905 60.085 2.075 ;
      RECT 57.775 0.085 58.11 1.055 ;
      RECT 57.775 -1.155 57.945 1.055 ;
      RECT 57.775 -1.155 58.03 -0.585 ;
      RECT 57.775 3.205 58.03 3.775 ;
      RECT 57.775 1.565 57.945 3.775 ;
      RECT 57.775 1.565 58.11 2.535 ;
      RECT 54.64 3.525 55.945 3.775 ;
      RECT 54.64 3.205 54.82 3.775 ;
      RECT 54.09 3.205 54.82 3.375 ;
      RECT 54.09 2.365 54.26 3.375 ;
      RECT 54.925 2.405 56.67 2.585 ;
      RECT 56.34 1.565 56.67 2.585 ;
      RECT 54.09 2.365 55.15 2.535 ;
      RECT 56.34 1.735 57.16 1.905 ;
      RECT 55.5 1.565 55.83 1.775 ;
      RECT 55.5 1.565 56.67 1.735 ;
      RECT 56.4 0.085 56.73 1.04 ;
      RECT 56.4 0.085 57.08 0.255 ;
      RECT 56.91 -1.155 57.08 0.255 ;
      RECT 56.82 -1.155 57.15 -0.515 ;
      RECT 55.945 0.355 56.22 1.055 ;
      RECT 56.05 -1.155 56.22 1.055 ;
      RECT 56.39 -0.335 56.74 -0.085 ;
      RECT 56.05 -0.305 56.74 -0.135 ;
      RECT 55.96 -1.155 56.22 -0.675 ;
      RECT 55.29 1.995 56.17 2.235 ;
      RECT 55.94 1.905 56.17 2.235 ;
      RECT 54.64 1.995 56.17 2.195 ;
      RECT 55.555 1.945 56.17 2.235 ;
      RECT 54.64 1.865 54.81 2.195 ;
      RECT 55.525 2.755 55.775 3.355 ;
      RECT 55.525 2.755 56 2.955 ;
      RECT 55.02 -0.025 55.775 0.475 ;
      RECT 54.09 -0.22 54.35 0.4 ;
      RECT 55.005 -0.08 55.02 0.225 ;
      RECT 54.99 -0.095 55.01 0.19 ;
      RECT 55.65 -0.42 55.88 0.18 ;
      RECT 54.965 -0.15 54.985 0.165 ;
      RECT 54.945 -0.025 55.88 0.15 ;
      RECT 54.92 -0.025 55.88 0.14 ;
      RECT 54.85 -0.025 55.88 0.13 ;
      RECT 54.83 -0.025 55.88 0.1 ;
      RECT 54.81 -1.115 54.98 0.07 ;
      RECT 54.78 -0.025 55.88 0.04 ;
      RECT 54.745 -0.025 55.88 0.015 ;
      RECT 54.715 -0.03 55.105 -0.02 ;
      RECT 54.715 -0.04 55.08 -0.02 ;
      RECT 54.715 -0.045 55.065 -0.02 ;
      RECT 54.715 -0.055 55.05 -0.02 ;
      RECT 54.09 -0.22 54.98 -0.05 ;
      RECT 54.09 -0.065 55.04 -0.05 ;
      RECT 54.09 -0.07 55.03 -0.05 ;
      RECT 54.985 -0.125 54.995 0.18 ;
      RECT 54.09 -0.09 55.015 -0.05 ;
      RECT 54.09 -0.11 55 -0.05 ;
      RECT 54.09 -1.115 54.98 -0.945 ;
      RECT 55.15 -0.62 55.48 -0.195 ;
      RECT 55.15 -1.105 55.37 -0.195 ;
      RECT 55.065 2.755 55.275 3.355 ;
      RECT 54.925 2.755 55.275 2.955 ;
      RECT 53.645 0.355 53.92 1.055 ;
      RECT 53.865 -1.155 53.92 1.055 ;
      RECT 53.75 -0.35 53.92 1.055 ;
      RECT 53.75 -1.155 53.92 -0.355 ;
      RECT 53.66 -1.155 53.92 -0.68 ;
      RECT 51.79 0.015 52.04 0.55 ;
      RECT 52.76 0.015 53.475 0.48 ;
      RECT 51.79 0.015 53.58 0.185 ;
      RECT 53.35 -0.35 53.58 0.185 ;
      RECT 52.345 -1.105 52.6 0.185 ;
      RECT 53.35 -0.415 53.41 0.48 ;
      RECT 53.41 -0.42 53.58 -0.355 ;
      RECT 51.81 -1.105 52.6 -0.84 ;
      RECT 52.77 2.705 53.445 2.955 ;
      RECT 53.18 2.345 53.445 2.955 ;
      RECT 52.93 3.125 53.26 3.675 ;
      RECT 51.87 3.125 53.26 3.315 ;
      RECT 51.87 2.285 52.04 3.315 ;
      RECT 51.75 2.705 52.04 3.035 ;
      RECT 51.87 2.285 52.81 2.455 ;
      RECT 52.51 1.735 52.81 2.455 ;
      RECT 52.77 -0.685 53.18 -0.165 ;
      RECT 52.77 -1.105 52.97 -0.165 ;
      RECT 51.38 -0.925 51.55 1.055 ;
      RECT 51.38 -0.415 52.175 -0.165 ;
      RECT 51.38 -0.925 51.63 -0.165 ;
      RECT 51.3 -0.925 51.63 -0.505 ;
      RECT 51.33 3.485 51.89 3.775 ;
      RECT 51.33 1.565 51.58 3.775 ;
      RECT 51.33 1.565 51.79 2.115 ;
      RECT 50.44 3.205 50.695 3.775 ;
      RECT 50.525 1.565 50.695 3.775 ;
      RECT 50.525 2.775 50.7 2.945 ;
      RECT 50.36 1.565 50.695 2.535 ;
      RECT 48.985 3.41 49.515 3.775 ;
      RECT 49.34 3.205 49.515 3.775 ;
      RECT 49.34 3.205 50.27 3.375 ;
      RECT 50.1 2.705 50.27 3.375 ;
      RECT 49.34 1.905 49.51 3.775 ;
      RECT 50.1 2.705 50.355 3.035 ;
      RECT 48.385 1.905 49.51 2.075 ;
      RECT 49.68 2.705 49.875 3.035 ;
      RECT 49.68 1.565 49.85 3.035 ;
      RECT 47.24 2.4 47.99 2.59 ;
      RECT 47.82 1.565 47.99 2.59 ;
      RECT 47.82 1.565 49.85 1.735 ;
      RECT 48.16 2.245 48.35 3.775 ;
      RECT 49 2.245 49.17 3.215 ;
      RECT 48.995 2.245 49.17 2.5 ;
      RECT 48.16 2.245 49.17 2.415 ;
      RECT 47.005 2.965 47.25 3.74 ;
      RECT 46.73 2.965 47.96 3.135 ;
      RECT 46.73 1.745 47.07 3.135 ;
      RECT 46.73 1.745 47.245 2.155 ;
      RECT 45.985 0.075 46.315 1.055 ;
      RECT 46.085 -1.155 46.315 1.055 ;
      RECT 45.985 -1.155 46.315 -0.525 ;
      RECT 45.985 3.145 46.315 3.775 ;
      RECT 46.085 1.565 46.315 3.775 ;
      RECT 45.985 1.565 46.315 2.545 ;
      RECT 44.605 0.075 44.935 1.055 ;
      RECT 44.705 -1.155 44.935 1.055 ;
      RECT 45.585 -0.335 45.915 -0.095 ;
      RECT 44.705 -0.305 45.915 -0.135 ;
      RECT 44.605 -1.155 44.935 -0.525 ;
      RECT 44.605 3.145 44.935 3.775 ;
      RECT 44.705 1.565 44.935 3.775 ;
      RECT 45.585 2.715 45.915 2.955 ;
      RECT 44.705 2.72 45.915 2.89 ;
      RECT 44.605 1.565 44.935 2.545 ;
      RECT 43.285 0.465 43.8 0.875 ;
      RECT 43.46 -0.515 43.8 0.875 ;
      RECT 42.57 -0.515 43.8 -0.345 ;
      RECT 43.28 -1.12 43.525 -0.345 ;
      RECT 43.28 2.965 43.525 3.74 ;
      RECT 42.57 2.965 43.8 3.135 ;
      RECT 43.46 1.745 43.8 3.135 ;
      RECT 43.285 1.745 43.8 2.155 ;
      RECT 40.68 0.885 42.71 1.055 ;
      RECT 42.54 0.03 42.71 1.055 ;
      RECT 40.68 -0.415 40.85 1.055 ;
      RECT 42.54 0.03 43.29 0.22 ;
      RECT 40.655 -0.415 40.85 -0.085 ;
      RECT 40.655 2.705 40.85 3.035 ;
      RECT 40.68 1.565 40.85 3.035 ;
      RECT 42.54 2.4 43.29 2.59 ;
      RECT 42.54 1.565 42.71 2.59 ;
      RECT 40.68 1.565 42.71 1.735 ;
      RECT 41.36 0.205 42.37 0.375 ;
      RECT 42.18 -1.155 42.37 0.375 ;
      RECT 41.36 -0.595 41.53 0.375 ;
      RECT 42.18 2.245 42.37 3.775 ;
      RECT 41.36 2.245 41.53 3.215 ;
      RECT 41.36 2.245 42.37 2.415 ;
      RECT 41.02 0.545 42.145 0.715 ;
      RECT 41.02 -1.155 41.19 0.715 ;
      RECT 40.175 -0.415 40.43 -0.085 ;
      RECT 40.26 -0.755 40.43 -0.085 ;
      RECT 40.26 -0.755 41.19 -0.585 ;
      RECT 41.015 -1.155 41.19 -0.585 ;
      RECT 41.015 -1.155 41.545 -0.79 ;
      RECT 41.015 3.41 41.545 3.775 ;
      RECT 41.015 3.205 41.19 3.775 ;
      RECT 41.02 1.905 41.19 3.775 ;
      RECT 40.26 3.205 41.19 3.375 ;
      RECT 40.26 2.705 40.43 3.375 ;
      RECT 40.175 2.705 40.43 3.035 ;
      RECT 41.02 1.905 42.145 2.075 ;
      RECT 39.835 0.085 40.17 1.055 ;
      RECT 39.835 -1.155 40.005 1.055 ;
      RECT 39.835 -1.155 40.09 -0.585 ;
      RECT 39.835 3.205 40.09 3.775 ;
      RECT 39.835 1.565 40.005 3.775 ;
      RECT 39.835 1.565 40.17 2.535 ;
      RECT 36.7 3.525 38.005 3.775 ;
      RECT 36.7 3.205 36.88 3.775 ;
      RECT 36.15 3.205 36.88 3.375 ;
      RECT 36.15 2.365 36.32 3.375 ;
      RECT 36.985 2.405 38.73 2.585 ;
      RECT 38.4 1.565 38.73 2.585 ;
      RECT 36.15 2.365 37.21 2.535 ;
      RECT 38.4 1.735 39.22 1.905 ;
      RECT 37.56 1.565 37.89 1.775 ;
      RECT 37.56 1.565 38.73 1.735 ;
      RECT 38.46 0.085 38.79 1.04 ;
      RECT 38.46 0.085 39.14 0.255 ;
      RECT 38.97 -1.155 39.14 0.255 ;
      RECT 38.88 -1.155 39.21 -0.515 ;
      RECT 38.005 0.355 38.28 1.055 ;
      RECT 38.11 -1.155 38.28 1.055 ;
      RECT 38.45 -0.335 38.8 -0.085 ;
      RECT 38.11 -0.305 38.8 -0.135 ;
      RECT 38.02 -1.155 38.28 -0.675 ;
      RECT 37.35 1.995 38.23 2.235 ;
      RECT 38 1.905 38.23 2.235 ;
      RECT 36.7 1.995 38.23 2.195 ;
      RECT 37.615 1.945 38.23 2.235 ;
      RECT 36.7 1.865 36.87 2.195 ;
      RECT 37.585 2.755 37.835 3.355 ;
      RECT 37.585 2.755 38.06 2.955 ;
      RECT 37.08 -0.025 37.835 0.475 ;
      RECT 36.15 -0.22 36.41 0.4 ;
      RECT 37.065 -0.08 37.08 0.225 ;
      RECT 37.05 -0.095 37.07 0.19 ;
      RECT 37.71 -0.42 37.94 0.18 ;
      RECT 37.025 -0.15 37.045 0.165 ;
      RECT 37.005 -0.025 37.94 0.15 ;
      RECT 36.98 -0.025 37.94 0.14 ;
      RECT 36.91 -0.025 37.94 0.13 ;
      RECT 36.89 -0.025 37.94 0.1 ;
      RECT 36.87 -1.115 37.04 0.07 ;
      RECT 36.84 -0.025 37.94 0.04 ;
      RECT 36.805 -0.025 37.94 0.015 ;
      RECT 36.775 -0.03 37.165 -0.02 ;
      RECT 36.775 -0.04 37.14 -0.02 ;
      RECT 36.775 -0.045 37.125 -0.02 ;
      RECT 36.775 -0.055 37.11 -0.02 ;
      RECT 36.15 -0.22 37.04 -0.05 ;
      RECT 36.15 -0.065 37.1 -0.05 ;
      RECT 36.15 -0.07 37.09 -0.05 ;
      RECT 37.045 -0.125 37.055 0.18 ;
      RECT 36.15 -0.09 37.075 -0.05 ;
      RECT 36.15 -0.11 37.06 -0.05 ;
      RECT 36.15 -1.115 37.04 -0.945 ;
      RECT 37.21 -0.62 37.54 -0.195 ;
      RECT 37.21 -1.105 37.43 -0.195 ;
      RECT 37.125 2.755 37.335 3.355 ;
      RECT 36.985 2.755 37.335 2.955 ;
      RECT 35.705 0.355 35.98 1.055 ;
      RECT 35.925 -1.155 35.98 1.055 ;
      RECT 35.81 -0.35 35.98 1.055 ;
      RECT 35.81 -1.155 35.98 -0.355 ;
      RECT 35.72 -1.155 35.98 -0.68 ;
      RECT 33.85 0.015 34.1 0.55 ;
      RECT 34.82 0.015 35.535 0.48 ;
      RECT 33.85 0.015 35.64 0.185 ;
      RECT 35.41 -0.35 35.64 0.185 ;
      RECT 34.405 -1.105 34.66 0.185 ;
      RECT 35.41 -0.415 35.47 0.48 ;
      RECT 35.47 -0.42 35.64 -0.355 ;
      RECT 33.87 -1.105 34.66 -0.84 ;
      RECT 34.83 2.705 35.505 2.955 ;
      RECT 35.24 2.345 35.505 2.955 ;
      RECT 34.99 3.125 35.32 3.675 ;
      RECT 33.93 3.125 35.32 3.315 ;
      RECT 33.93 2.285 34.1 3.315 ;
      RECT 33.81 2.705 34.1 3.035 ;
      RECT 33.93 2.285 34.87 2.455 ;
      RECT 34.57 1.735 34.87 2.455 ;
      RECT 34.83 -0.685 35.24 -0.165 ;
      RECT 34.83 -1.105 35.03 -0.165 ;
      RECT 33.44 -0.925 33.61 1.055 ;
      RECT 33.44 -0.415 34.235 -0.165 ;
      RECT 33.44 -0.925 33.69 -0.165 ;
      RECT 33.36 -0.925 33.69 -0.505 ;
      RECT 33.39 3.485 33.95 3.775 ;
      RECT 33.39 1.565 33.64 3.775 ;
      RECT 33.39 1.565 33.85 2.115 ;
      RECT 32.5 3.205 32.755 3.775 ;
      RECT 32.585 1.565 32.755 3.775 ;
      RECT 32.585 2.775 32.76 2.945 ;
      RECT 32.42 1.565 32.755 2.535 ;
      RECT 31.045 3.41 31.575 3.775 ;
      RECT 31.4 3.205 31.575 3.775 ;
      RECT 31.4 3.205 32.33 3.375 ;
      RECT 32.16 2.705 32.33 3.375 ;
      RECT 31.4 1.905 31.57 3.775 ;
      RECT 32.16 2.705 32.415 3.035 ;
      RECT 30.445 1.905 31.57 2.075 ;
      RECT 31.74 2.705 31.935 3.035 ;
      RECT 31.74 1.565 31.91 3.035 ;
      RECT 29.3 2.4 30.05 2.59 ;
      RECT 29.88 1.565 30.05 2.59 ;
      RECT 29.88 1.565 31.91 1.735 ;
      RECT 30.22 2.245 30.41 3.775 ;
      RECT 31.06 2.245 31.23 3.215 ;
      RECT 31.055 2.245 31.23 2.5 ;
      RECT 30.22 2.245 31.23 2.415 ;
      RECT 29.065 2.965 29.31 3.74 ;
      RECT 28.79 2.965 30.02 3.135 ;
      RECT 28.79 1.745 29.13 3.135 ;
      RECT 28.79 1.745 29.305 2.155 ;
      RECT 28.045 0.075 28.375 1.055 ;
      RECT 28.145 -1.155 28.375 1.055 ;
      RECT 28.045 -1.155 28.375 -0.525 ;
      RECT 28.045 3.145 28.375 3.775 ;
      RECT 28.145 1.565 28.375 3.775 ;
      RECT 28.045 1.565 28.375 2.545 ;
      RECT 26.665 0.075 26.995 1.055 ;
      RECT 26.765 -1.155 26.995 1.055 ;
      RECT 27.645 -0.335 27.975 -0.095 ;
      RECT 26.765 -0.305 27.975 -0.135 ;
      RECT 26.665 -1.155 26.995 -0.525 ;
      RECT 26.665 3.145 26.995 3.775 ;
      RECT 26.765 1.565 26.995 3.775 ;
      RECT 27.645 2.715 27.975 2.955 ;
      RECT 26.765 2.72 27.975 2.89 ;
      RECT 26.665 1.565 26.995 2.545 ;
      RECT 25.345 0.465 25.86 0.875 ;
      RECT 25.52 -0.515 25.86 0.875 ;
      RECT 24.63 -0.515 25.86 -0.345 ;
      RECT 25.34 -1.12 25.585 -0.345 ;
      RECT 25.34 2.965 25.585 3.74 ;
      RECT 24.63 2.965 25.86 3.135 ;
      RECT 25.52 1.745 25.86 3.135 ;
      RECT 25.345 1.745 25.86 2.155 ;
      RECT 22.74 0.885 24.77 1.055 ;
      RECT 24.6 0.03 24.77 1.055 ;
      RECT 22.74 -0.415 22.91 1.055 ;
      RECT 24.6 0.03 25.35 0.22 ;
      RECT 22.715 -0.415 22.91 -0.085 ;
      RECT 22.715 2.705 22.91 3.035 ;
      RECT 22.74 1.565 22.91 3.035 ;
      RECT 24.6 2.4 25.35 2.59 ;
      RECT 24.6 1.565 24.77 2.59 ;
      RECT 22.74 1.565 24.77 1.735 ;
      RECT 23.42 0.205 24.43 0.375 ;
      RECT 24.24 -1.155 24.43 0.375 ;
      RECT 23.42 -0.595 23.59 0.375 ;
      RECT 24.24 2.245 24.43 3.775 ;
      RECT 23.42 2.245 23.59 3.215 ;
      RECT 23.42 2.245 24.43 2.415 ;
      RECT 23.08 0.545 24.205 0.715 ;
      RECT 23.08 -1.155 23.25 0.715 ;
      RECT 22.235 -0.415 22.49 -0.085 ;
      RECT 22.32 -0.755 22.49 -0.085 ;
      RECT 22.32 -0.755 23.25 -0.585 ;
      RECT 23.075 -1.155 23.25 -0.585 ;
      RECT 23.075 -1.155 23.605 -0.79 ;
      RECT 23.075 3.41 23.605 3.775 ;
      RECT 23.075 3.205 23.25 3.775 ;
      RECT 23.08 1.905 23.25 3.775 ;
      RECT 22.32 3.205 23.25 3.375 ;
      RECT 22.32 2.705 22.49 3.375 ;
      RECT 22.235 2.705 22.49 3.035 ;
      RECT 23.08 1.905 24.205 2.075 ;
      RECT 21.895 0.085 22.23 1.055 ;
      RECT 21.895 -1.155 22.065 1.055 ;
      RECT 21.895 -1.155 22.15 -0.585 ;
      RECT 21.895 3.205 22.15 3.775 ;
      RECT 21.895 1.565 22.065 3.775 ;
      RECT 21.895 1.565 22.23 2.535 ;
      RECT 18.76 3.525 20.065 3.775 ;
      RECT 18.76 3.205 18.94 3.775 ;
      RECT 18.21 3.205 18.94 3.375 ;
      RECT 18.21 2.365 18.38 3.375 ;
      RECT 19.045 2.405 20.79 2.585 ;
      RECT 20.46 1.565 20.79 2.585 ;
      RECT 18.21 2.365 19.27 2.535 ;
      RECT 20.46 1.735 21.28 1.905 ;
      RECT 19.62 1.565 19.95 1.775 ;
      RECT 19.62 1.565 20.79 1.735 ;
      RECT 20.52 0.085 20.85 1.04 ;
      RECT 20.52 0.085 21.2 0.255 ;
      RECT 21.03 -1.155 21.2 0.255 ;
      RECT 20.94 -1.155 21.27 -0.515 ;
      RECT 20.065 0.355 20.34 1.055 ;
      RECT 20.17 -1.155 20.34 1.055 ;
      RECT 20.51 -0.335 20.86 -0.085 ;
      RECT 20.17 -0.305 20.86 -0.135 ;
      RECT 20.08 -1.155 20.34 -0.675 ;
      RECT 19.41 1.995 20.29 2.235 ;
      RECT 20.06 1.905 20.29 2.235 ;
      RECT 18.76 1.995 20.29 2.195 ;
      RECT 19.675 1.945 20.29 2.235 ;
      RECT 18.76 1.865 18.93 2.195 ;
      RECT 19.645 2.755 19.895 3.355 ;
      RECT 19.645 2.755 20.12 2.955 ;
      RECT 19.14 -0.025 19.895 0.475 ;
      RECT 18.21 -0.22 18.47 0.4 ;
      RECT 19.125 -0.08 19.14 0.225 ;
      RECT 19.11 -0.095 19.13 0.19 ;
      RECT 19.77 -0.42 20 0.18 ;
      RECT 19.085 -0.15 19.105 0.165 ;
      RECT 19.065 -0.025 20 0.15 ;
      RECT 19.04 -0.025 20 0.14 ;
      RECT 18.97 -0.025 20 0.13 ;
      RECT 18.95 -0.025 20 0.1 ;
      RECT 18.93 -1.115 19.1 0.07 ;
      RECT 18.9 -0.025 20 0.04 ;
      RECT 18.865 -0.025 20 0.015 ;
      RECT 18.835 -0.03 19.225 -0.02 ;
      RECT 18.835 -0.04 19.2 -0.02 ;
      RECT 18.835 -0.045 19.185 -0.02 ;
      RECT 18.835 -0.055 19.17 -0.02 ;
      RECT 18.21 -0.22 19.1 -0.05 ;
      RECT 18.21 -0.065 19.16 -0.05 ;
      RECT 18.21 -0.07 19.15 -0.05 ;
      RECT 19.105 -0.125 19.115 0.18 ;
      RECT 18.21 -0.09 19.135 -0.05 ;
      RECT 18.21 -0.11 19.12 -0.05 ;
      RECT 18.21 -1.115 19.1 -0.945 ;
      RECT 19.27 -0.62 19.6 -0.195 ;
      RECT 19.27 -1.105 19.49 -0.195 ;
      RECT 19.185 2.755 19.395 3.355 ;
      RECT 19.045 2.755 19.395 2.955 ;
      RECT 17.765 0.355 18.04 1.055 ;
      RECT 17.985 -1.155 18.04 1.055 ;
      RECT 17.87 -0.35 18.04 1.055 ;
      RECT 17.87 -1.155 18.04 -0.355 ;
      RECT 17.78 -1.155 18.04 -0.68 ;
      RECT 15.91 0.015 16.16 0.55 ;
      RECT 16.88 0.015 17.595 0.48 ;
      RECT 15.91 0.015 17.7 0.185 ;
      RECT 17.47 -0.35 17.7 0.185 ;
      RECT 16.465 -1.105 16.72 0.185 ;
      RECT 17.47 -0.415 17.53 0.48 ;
      RECT 17.53 -0.42 17.7 -0.355 ;
      RECT 15.93 -1.105 16.72 -0.84 ;
      RECT 16.89 2.705 17.565 2.955 ;
      RECT 17.3 2.345 17.565 2.955 ;
      RECT 17.05 3.125 17.38 3.675 ;
      RECT 15.99 3.125 17.38 3.315 ;
      RECT 15.99 2.285 16.16 3.315 ;
      RECT 15.87 2.705 16.16 3.035 ;
      RECT 15.99 2.285 16.93 2.455 ;
      RECT 16.63 1.735 16.93 2.455 ;
      RECT 16.89 -0.685 17.3 -0.165 ;
      RECT 16.89 -1.105 17.09 -0.165 ;
      RECT 15.5 -0.925 15.67 1.055 ;
      RECT 15.5 -0.415 16.295 -0.165 ;
      RECT 15.5 -0.925 15.75 -0.165 ;
      RECT 15.42 -0.925 15.75 -0.505 ;
      RECT 15.45 3.485 16.01 3.775 ;
      RECT 15.45 1.565 15.7 3.775 ;
      RECT 15.45 1.565 15.91 2.115 ;
      RECT 14.56 3.205 14.815 3.775 ;
      RECT 14.645 1.565 14.815 3.775 ;
      RECT 14.645 2.775 14.82 2.945 ;
      RECT 14.48 1.565 14.815 2.535 ;
      RECT 13.105 3.41 13.635 3.775 ;
      RECT 13.46 3.205 13.635 3.775 ;
      RECT 13.46 3.205 14.39 3.375 ;
      RECT 14.22 2.705 14.39 3.375 ;
      RECT 13.46 1.905 13.63 3.775 ;
      RECT 14.22 2.705 14.475 3.035 ;
      RECT 12.505 1.905 13.63 2.075 ;
      RECT 13.8 2.705 13.995 3.035 ;
      RECT 13.8 1.565 13.97 3.035 ;
      RECT 11.36 2.4 12.11 2.59 ;
      RECT 11.94 1.565 12.11 2.59 ;
      RECT 11.94 1.565 13.97 1.735 ;
      RECT 12.28 2.245 12.47 3.775 ;
      RECT 13.12 2.245 13.29 3.215 ;
      RECT 13.115 2.245 13.29 2.5 ;
      RECT 12.28 2.245 13.29 2.415 ;
      RECT 11.125 2.965 11.37 3.74 ;
      RECT 10.85 2.965 12.08 3.135 ;
      RECT 10.85 1.745 11.19 3.135 ;
      RECT 10.85 1.745 11.365 2.155 ;
      RECT -3.355 2.935 -3.185 4.245 ;
      RECT -0.815 2.935 -0.645 3.865 ;
      RECT -3.95 2.935 0.335 3.105 ;
      RECT -3.95 5.655 0.19 5.825 ;
      RECT -1.145 5.12 -0.635 5.825 ;
      RECT -3.435 5.255 -3.105 5.825 ;
      RECT -0.415 4.675 -0.17 5.45 ;
      RECT -1.125 4.675 0.105 4.845 ;
      RECT -0.235 3.455 0.105 4.845 ;
      RECT -0.41 3.455 0.105 3.865 ;
      RECT -3.04 4.415 -2.845 4.745 ;
      RECT -3.015 3.275 -2.845 4.745 ;
      RECT -1.155 4.11 -0.405 4.3 ;
      RECT -1.155 3.275 -0.985 4.3 ;
      RECT -3.015 3.275 -0.985 3.445 ;
      RECT -1.515 3.955 -1.325 5.485 ;
      RECT -2.335 3.955 -2.165 4.925 ;
      RECT -2.335 3.955 -1.325 4.125 ;
      RECT -2.68 5.12 -2.15 5.485 ;
      RECT -2.68 4.915 -2.505 5.485 ;
      RECT -2.675 3.615 -2.505 5.485 ;
      RECT -3.435 4.915 -2.505 5.085 ;
      RECT -3.435 4.415 -3.265 5.085 ;
      RECT -3.52 4.415 -3.265 4.745 ;
      RECT -2.675 3.615 -1.55 3.785 ;
      RECT -3.86 4.915 -3.605 5.485 ;
      RECT -3.86 3.275 -3.69 5.485 ;
      RECT -3.86 3.275 -3.525 4.245 ;
      RECT 98.02 -0.335 98.35 -0.095 ;
      RECT 98.02 2.715 98.35 2.955 ;
      RECT 95.55 -1.155 95.825 0.005 ;
      RECT 95.55 2.615 95.825 3.775 ;
      RECT 93.125 -0.335 93.475 -0.085 ;
      RECT 92.065 2.755 92.515 3.265 ;
      RECT 90.745 0.715 91.225 1.055 ;
      RECT 90.305 2.705 90.63 3.035 ;
      RECT 89.965 -0.775 90.515 -0.39 ;
      RECT 89.305 4.915 89.475 5.085 ;
      RECT 88.45 0.715 88.925 1.055 ;
      RECT 88.085 2.705 88.425 2.955 ;
      RECT 86.745 -0.335 87.085 0.545 ;
      RECT 80.08 -0.335 80.41 -0.095 ;
      RECT 80.08 2.715 80.41 2.955 ;
      RECT 77.61 -1.155 77.885 0.005 ;
      RECT 77.61 2.615 77.885 3.775 ;
      RECT 75.185 -0.335 75.535 -0.085 ;
      RECT 74.125 2.755 74.575 3.265 ;
      RECT 72.805 0.715 73.285 1.055 ;
      RECT 72.365 2.705 72.69 3.035 ;
      RECT 72.025 -0.775 72.575 -0.39 ;
      RECT 71.365 3.655 71.535 3.825 ;
      RECT 70.51 0.715 70.985 1.055 ;
      RECT 70.145 2.705 70.485 2.955 ;
      RECT 68.805 -0.335 69.145 0.545 ;
      RECT 62.145 -0.335 62.475 -0.095 ;
      RECT 62.145 2.715 62.475 2.955 ;
      RECT 59.675 -1.155 59.95 0.005 ;
      RECT 59.675 2.615 59.95 3.775 ;
      RECT 57.25 -0.335 57.6 -0.085 ;
      RECT 56.19 2.755 56.64 3.265 ;
      RECT 54.87 0.715 55.35 1.055 ;
      RECT 54.43 2.705 54.755 3.035 ;
      RECT 54.09 -0.775 54.64 -0.39 ;
      RECT 53.43 3.655 53.6 3.825 ;
      RECT 52.575 0.715 53.05 1.055 ;
      RECT 52.21 2.705 52.55 2.955 ;
      RECT 50.87 -0.335 51.21 0.545 ;
      RECT 44.205 -0.335 44.535 -0.095 ;
      RECT 44.205 2.715 44.535 2.955 ;
      RECT 41.735 -1.155 42.01 0.005 ;
      RECT 41.735 2.615 42.01 3.775 ;
      RECT 39.31 -0.335 39.66 -0.085 ;
      RECT 38.25 2.755 38.7 3.265 ;
      RECT 36.93 0.715 37.41 1.055 ;
      RECT 36.49 2.705 36.815 3.035 ;
      RECT 36.15 -0.775 36.7 -0.39 ;
      RECT 35.46 3.625 35.69 3.855 ;
      RECT 34.635 0.715 35.11 1.055 ;
      RECT 34.27 2.705 34.61 2.955 ;
      RECT 32.93 -0.335 33.27 0.545 ;
      RECT 26.265 -0.335 26.595 -0.095 ;
      RECT 26.265 2.715 26.595 2.955 ;
      RECT 23.795 -1.155 24.07 0.005 ;
      RECT 23.795 2.615 24.07 3.775 ;
      RECT 21.37 -0.335 21.72 -0.085 ;
      RECT 20.31 2.755 20.76 3.265 ;
      RECT 18.99 0.715 19.47 1.055 ;
      RECT 18.55 2.705 18.875 3.035 ;
      RECT 18.21 -0.775 18.76 -0.39 ;
      RECT 17.55 3.655 17.72 3.825 ;
      RECT 16.695 0.715 17.17 1.055 ;
      RECT 16.33 2.705 16.67 2.955 ;
      RECT 14.99 -0.335 15.33 0.545 ;
      RECT 0.865 4.11 1.035 4.28 ;
      RECT -3.95 0.215 0.405 0.39 ;
      RECT 0.31 5.71 0.335 5.76 ;
      RECT 0.31 5.82 0.335 5.825 ;
      RECT -1.96 4.325 -1.685 5.485 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r1

END LIBRARY
