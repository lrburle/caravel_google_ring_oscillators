magic
tech sky130A
magscale 1 2
timestamp 1703004377
<< obsli1 >>
rect 292000 197600 526832 451376
<< obsm1 >>
rect 289722 195848 580230 451376
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
<< obsm2 >>
rect 289728 6559 580318 452849
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 291009 444988 583520 452845
rect 291009 444588 583440 444988
rect 291009 431796 583520 444588
rect 291009 431396 583440 431796
rect 291009 418468 583520 431396
rect 291009 418068 583440 418468
rect 291009 405140 583520 418068
rect 291009 404740 583440 405140
rect 291009 391948 583520 404740
rect 291009 391548 583440 391948
rect 291009 378620 583520 391548
rect 291009 378220 583440 378620
rect 291009 365292 583520 378220
rect 291009 364892 583440 365292
rect 291009 352100 583520 364892
rect 291009 351700 583440 352100
rect 291009 338772 583520 351700
rect 291009 338372 583440 338772
rect 291009 325444 583520 338372
rect 291009 325044 583440 325444
rect 291009 312252 583520 325044
rect 291009 311852 583440 312252
rect 291009 298924 583520 311852
rect 291009 298524 583440 298924
rect 291009 285596 583520 298524
rect 291009 285196 583440 285596
rect 291009 272404 583520 285196
rect 291009 272004 583440 272404
rect 291009 259076 583520 272004
rect 291009 258676 583440 259076
rect 291009 245748 583520 258676
rect 291009 245348 583440 245748
rect 291009 232556 583520 245348
rect 291009 232156 583440 232556
rect 291009 219228 583520 232156
rect 291009 218828 583440 219228
rect 291009 205900 583520 218828
rect 291009 205500 583440 205900
rect 291009 192708 583520 205500
rect 291009 192308 583440 192708
rect 291009 179380 583520 192308
rect 291009 178980 583440 179380
rect 291009 166052 583520 178980
rect 291009 165652 583440 166052
rect 291009 152860 583520 165652
rect 291009 152460 583440 152860
rect 291009 139532 583520 152460
rect 291009 139132 583440 139532
rect 291009 126204 583520 139132
rect 291009 125804 583440 126204
rect 291009 113012 583520 125804
rect 291009 112612 583440 113012
rect 291009 99684 583520 112612
rect 291009 99284 583440 99684
rect 291009 86356 583520 99284
rect 291009 85956 583440 86356
rect 291009 73164 583520 85956
rect 291009 72764 583440 73164
rect 291009 59836 583520 72764
rect 291009 59436 583440 59836
rect 291009 46508 583520 59436
rect 291009 46108 583440 46508
rect 291009 33316 583520 46108
rect 291009 32916 583440 33316
rect 291009 19988 583520 32916
rect 291009 19588 583440 19988
rect 291009 6796 583520 19588
rect 291009 6563 583440 6796
<< metal4 >>
rect -4950 -3878 -3538 707814
rect -3198 -2126 -1786 706062
rect 1144 -2294 1464 706230
rect 2876 -2294 3196 706230
rect 8144 -2294 8464 706230
rect 9876 -2294 10196 706230
rect 15144 -2294 15464 706230
rect 16876 -2294 17196 706230
rect 22144 -2294 22464 706230
rect 23876 -2294 24196 706230
rect 29144 -2294 29464 706230
rect 30876 -2294 31196 706230
rect 36144 -2294 36464 706230
rect 37876 -2294 38196 706230
rect 43144 -2294 43464 706230
rect 44876 -2294 45196 706230
rect 50144 -2294 50464 706230
rect 51876 -2294 52196 706230
rect 57144 -2294 57464 706230
rect 58876 -2294 59196 706230
rect 64144 -2294 64464 706230
rect 65876 -2294 66196 706230
rect 71144 -2294 71464 706230
rect 72876 -2294 73196 706230
rect 78144 -2294 78464 706230
rect 79876 -2294 80196 706230
rect 85144 -2294 85464 706230
rect 86876 -2294 87196 706230
rect 92144 -2294 92464 706230
rect 93876 -2294 94196 706230
rect 99144 -2294 99464 706230
rect 100876 -2294 101196 706230
rect 106144 -2294 106464 706230
rect 107876 -2294 108196 706230
rect 113144 -2294 113464 706230
rect 114876 -2294 115196 706230
rect 120144 -2294 120464 706230
rect 121876 -2294 122196 706230
rect 127144 -2294 127464 706230
rect 128876 -2294 129196 706230
rect 134144 -2294 134464 706230
rect 135876 -2294 136196 706230
rect 141144 -2294 141464 706230
rect 142876 -2294 143196 706230
rect 148144 -2294 148464 706230
rect 149876 -2294 150196 706230
rect 155144 -2294 155464 706230
rect 156876 -2294 157196 706230
rect 162144 -2294 162464 706230
rect 163876 -2294 164196 706230
rect 169144 -2294 169464 706230
rect 170876 -2294 171196 706230
rect 176144 -2294 176464 706230
rect 177876 -2294 178196 706230
rect 183144 -2294 183464 706230
rect 184876 -2294 185196 706230
rect 190144 -2294 190464 706230
rect 191876 -2294 192196 706230
rect 197144 -2294 197464 706230
rect 198876 -2294 199196 706230
rect 204144 -2294 204464 706230
rect 205876 -2294 206196 706230
rect 211144 -2294 211464 706230
rect 212876 -2294 213196 706230
rect 218144 -2294 218464 706230
rect 219876 -2294 220196 706230
rect 225144 -2294 225464 706230
rect 226876 -2294 227196 706230
rect 232144 -2294 232464 706230
rect 233876 -2294 234196 706230
rect 239144 -2294 239464 706230
rect 240876 -2294 241196 706230
rect 246144 -2294 246464 706230
rect 247876 -2294 248196 706230
rect 253144 -2294 253464 706230
rect 254876 -2294 255196 706230
rect 260144 -2294 260464 706230
rect 261876 -2294 262196 706230
rect 267144 -2294 267464 706230
rect 268876 -2294 269196 706230
rect 274144 -2294 274464 706230
rect 275876 -2294 276196 706230
rect 281144 -2294 281464 706230
rect 282876 -2294 283196 706230
rect 288144 -2294 288464 706230
rect 289876 -2294 290196 706230
rect 295144 368380 295464 706230
rect 296876 368380 297196 706230
rect 302144 368380 302464 706230
rect 303876 368380 304196 706230
rect 295144 200380 295464 363976
rect 296876 200380 297196 363976
rect 302144 200380 302464 363976
rect 303876 200380 304196 363976
rect 295144 -2294 295464 195976
rect 296876 -2294 297196 195976
rect 302144 -2294 302464 195976
rect 303876 -2294 304196 195976
rect 309144 -2294 309464 706230
rect 310876 -2294 311196 706230
rect 316144 -2294 316464 706230
rect 317876 -2294 318196 706230
rect 323144 -2294 323464 706230
rect 324876 -2294 325196 706230
rect 330144 -2294 330464 706230
rect 331876 -2294 332196 706230
rect 337144 -2294 337464 706230
rect 338876 -2294 339196 706230
rect 344144 -2294 344464 706230
rect 345876 -2294 346196 706230
rect 351144 -2294 351464 706230
rect 352876 -2294 353196 706230
rect 358144 -2294 358464 706230
rect 359876 -2294 360196 706230
rect 365144 -2294 365464 706230
rect 366876 -2294 367196 706230
rect 372144 -2294 372464 706230
rect 373876 -2294 374196 706230
rect 379144 -2294 379464 706230
rect 380876 -2294 381196 706230
rect 386144 -2294 386464 706230
rect 387876 -2294 388196 706230
rect 393144 -2294 393464 706230
rect 394876 -2294 395196 706230
rect 400144 -2294 400464 706230
rect 401876 -2294 402196 706230
rect 407144 -2294 407464 706230
rect 408876 -2294 409196 706230
rect 414144 -2294 414464 706230
rect 415876 -2294 416196 706230
rect 421144 -2294 421464 706230
rect 422876 -2294 423196 706230
rect 428144 -2294 428464 706230
rect 429876 -2294 430196 706230
rect 435144 -2294 435464 706230
rect 436876 -2294 437196 706230
rect 442144 -2294 442464 706230
rect 443876 -2294 444196 706230
rect 449144 -2294 449464 706230
rect 450876 -2294 451196 706230
rect 456144 -2294 456464 706230
rect 457876 -2294 458196 706230
rect 463144 -2294 463464 706230
rect 464876 -2294 465196 706230
rect 470144 -2294 470464 706230
rect 471876 -2294 472196 706230
rect 477144 -2294 477464 706230
rect 478876 -2294 479196 706230
rect 484144 -2294 484464 706230
rect 485876 -2294 486196 706230
rect 491144 -2294 491464 706230
rect 492876 -2294 493196 706230
rect 498144 -2294 498464 706230
rect 499876 -2294 500196 706230
rect 505144 -2294 505464 706230
rect 506876 -2294 507196 706230
rect 512144 -2294 512464 706230
rect 513876 -2294 514196 706230
rect 519144 -2294 519464 706230
rect 520876 421752 521196 706230
rect 526144 421752 526464 706230
rect 520876 381752 521196 400008
rect 526144 381752 526464 400008
rect 520876 341752 521196 360008
rect 526144 341752 526464 360008
rect 520876 301752 521196 320008
rect 526144 301752 526464 320008
rect 520876 261752 521196 280008
rect 526144 261752 526464 280008
rect 520876 -2294 521196 240008
rect 526144 -2294 526464 240008
rect 527876 -2294 528196 706230
rect 533144 -2294 533464 706230
rect 534876 -2294 535196 706230
rect 540144 -2294 540464 706230
rect 541876 -2294 542196 706230
rect 547144 -2294 547464 706230
rect 548876 -2294 549196 706230
rect 554144 -2294 554464 706230
rect 555876 -2294 556196 706230
rect 561144 -2294 561464 706230
rect 562876 -2294 563196 706230
rect 568144 -2294 568464 706230
rect 569876 -2294 570196 706230
rect 575144 -2294 575464 706230
rect 576876 -2294 577196 706230
rect 582144 -2294 582464 706230
rect 585710 -2126 587122 706062
rect 587462 -3878 588874 707814
<< obsm4 >>
rect 293139 368300 295064 419632
rect 295544 368300 296796 419632
rect 297276 368300 302064 419632
rect 302544 368300 303796 419632
rect 304276 368300 309064 419632
rect 293139 364056 309064 368300
rect 293139 200300 295064 364056
rect 295544 200300 296796 364056
rect 297276 200300 302064 364056
rect 302544 200300 303796 364056
rect 304276 200300 309064 364056
rect 293139 198096 309064 200300
rect 309544 198096 310796 419632
rect 311276 198096 316064 419632
rect 316544 198096 317796 419632
rect 318276 198096 323064 419632
rect 323544 198096 324796 419632
rect 325276 198096 330064 419632
rect 330544 198096 331796 419632
rect 332276 198096 337064 419632
rect 337544 198096 338796 419632
rect 339276 198096 344064 419632
rect 344544 198096 345796 419632
rect 346276 198096 351064 419632
rect 351544 198096 352796 419632
rect 353276 198096 358064 419632
rect 358544 198096 359796 419632
rect 360276 198096 365064 419632
rect 365544 198096 366796 419632
rect 367276 198096 372064 419632
rect 372544 198096 373796 419632
rect 374276 198096 379064 419632
rect 379544 198096 380796 419632
rect 381276 198096 386064 419632
rect 386544 198096 387796 419632
rect 388276 198096 393064 419632
rect 393544 198096 394796 419632
rect 395276 198096 400064 419632
rect 400544 198096 401796 419632
rect 402276 198096 407064 419632
rect 407544 198096 408796 419632
rect 409276 198096 414064 419632
rect 414544 198096 415796 419632
rect 416276 198096 421064 419632
rect 421544 198096 422796 419632
rect 423276 198096 428064 419632
rect 428544 198096 429796 419632
rect 430276 198096 435064 419632
rect 435544 198096 436796 419632
rect 437276 198096 442064 419632
rect 442544 198096 443796 419632
rect 444276 198096 449064 419632
rect 449544 198096 450796 419632
rect 451276 198096 456064 419632
rect 456544 198096 457796 419632
rect 458276 198096 463064 419632
rect 463544 198096 464796 419632
rect 465276 198096 470064 419632
rect 470544 198096 471796 419632
rect 472276 198096 477064 419632
rect 477544 198096 478796 419632
rect 479276 198096 484064 419632
rect 484544 198096 485796 419632
rect 486276 198096 491064 419632
rect 491544 198096 492796 419632
rect 493276 198096 498064 419632
rect 498544 198096 499796 419632
rect 500276 198096 505064 419632
rect 505544 198096 506796 419632
rect 507276 198096 512064 419632
rect 512544 198096 513796 419632
rect 514276 198096 519064 419632
rect 519544 400088 526992 419632
rect 519544 381672 520796 400088
rect 521276 381672 526064 400088
rect 526544 381672 526992 400088
rect 519544 360088 526992 381672
rect 519544 341672 520796 360088
rect 521276 341672 526064 360088
rect 526544 341672 526992 360088
rect 519544 320088 526992 341672
rect 519544 301672 520796 320088
rect 521276 301672 526064 320088
rect 526544 301672 526992 320088
rect 519544 280088 526992 301672
rect 519544 261672 520796 280088
rect 521276 261672 526064 280088
rect 526544 261672 526992 280088
rect 519544 240088 526992 261672
rect 519544 198096 520796 240088
rect 521276 198096 526064 240088
rect 526544 198096 526992 240088
<< metal5 >>
rect -3366 705610 587290 706230
rect -2406 704650 587122 705270
rect -4950 696156 588874 696476
rect -4950 695216 588874 695536
rect -4950 689156 588874 689476
rect -4950 688216 588874 688536
rect -4950 682156 588874 682476
rect -4950 681216 588874 681536
rect -4950 675156 588874 675476
rect -4950 674216 588874 674536
rect -4950 668156 588874 668476
rect -4950 667216 588874 667536
rect -4950 661156 588874 661476
rect -4950 660216 588874 660536
rect -4950 654156 588874 654476
rect -4950 653216 588874 653536
rect -4950 647156 588874 647476
rect -4950 646216 588874 646536
rect -4950 640156 588874 640476
rect -4950 639216 588874 639536
rect -4950 633156 588874 633476
rect -4950 632216 588874 632536
rect -4950 626156 588874 626476
rect -4950 625216 588874 625536
rect -4950 619156 588874 619476
rect -4950 618216 588874 618536
rect -4950 612156 588874 612476
rect -4950 611216 588874 611536
rect -4950 605156 588874 605476
rect -4950 604216 588874 604536
rect -4950 598156 588874 598476
rect -4950 597216 588874 597536
rect -4950 591156 588874 591476
rect -4950 590216 588874 590536
rect -4950 584156 588874 584476
rect -4950 583216 588874 583536
rect -4950 577156 588874 577476
rect -4950 576216 588874 576536
rect -4950 570156 588874 570476
rect -4950 569216 588874 569536
rect -4950 563156 588874 563476
rect -4950 562216 588874 562536
rect -4950 556156 588874 556476
rect -4950 555216 588874 555536
rect -4950 549156 588874 549476
rect -4950 548216 588874 548536
rect -4950 542156 588874 542476
rect -4950 541216 588874 541536
rect -4950 535156 588874 535476
rect -4950 534216 588874 534536
rect -4950 528156 588874 528476
rect -4950 527216 588874 527536
rect -4950 521156 588874 521476
rect -4950 520216 588874 520536
rect -4950 514156 588874 514476
rect -4950 513216 588874 513536
rect -4950 507156 588874 507476
rect -4950 506216 588874 506536
rect -4950 500156 588874 500476
rect -4950 499216 588874 499536
rect -4950 493156 588874 493476
rect -4950 492216 588874 492536
rect -4950 486156 588874 486476
rect -4950 485216 588874 485536
rect -4950 479156 588874 479476
rect -4950 478216 588874 478536
rect -4950 472156 588874 472476
rect -4950 471216 588874 471536
rect -4950 465156 588874 465476
rect -4950 464216 588874 464536
rect -4950 458156 588874 458476
rect -4950 457216 588874 457536
rect -4950 451156 588874 451476
rect -4950 450216 588874 450536
rect -4950 444156 588874 444476
rect -4950 443216 588874 443536
rect -4950 437156 588874 437476
rect -4950 436216 588874 436536
rect -4950 430156 588874 430476
rect -4950 429216 588874 429536
rect -4950 423156 588874 423476
rect -4950 422216 588874 422536
rect -4950 416156 588874 416476
rect -4950 415216 588874 415536
rect -4950 409156 588874 409476
rect -4950 408216 588874 408536
rect -4950 402156 588874 402476
rect -4950 401216 588874 401536
rect -4950 395156 588874 395476
rect -4950 394216 588874 394536
rect -4950 388156 588874 388476
rect -4950 387216 588874 387536
rect -4950 381156 588874 381476
rect -4950 380216 588874 380536
rect -4950 374156 588874 374476
rect -4950 373216 588874 373536
rect -4950 367156 588874 367476
rect -4950 366216 588874 366536
rect -4950 360156 588874 360476
rect -4950 359216 588874 359536
rect -4950 353156 588874 353476
rect -4950 352216 588874 352536
rect -4950 346156 588874 346476
rect -4950 345216 588874 345536
rect -4950 339156 588874 339476
rect -4950 338216 588874 338536
rect -4950 332156 588874 332476
rect -4950 331216 588874 331536
rect -4950 325156 588874 325476
rect -4950 324216 588874 324536
rect -4950 318156 588874 318476
rect -4950 317216 588874 317536
rect -4950 311156 588874 311476
rect -4950 310216 588874 310536
rect -4950 304156 588874 304476
rect -4950 303216 588874 303536
rect -4950 297156 588874 297476
rect -4950 296216 588874 296536
rect -4950 290156 588874 290476
rect -4950 289216 588874 289536
rect -4950 283156 588874 283476
rect -4950 282216 588874 282536
rect -4950 276156 588874 276476
rect -4950 275216 588874 275536
rect -4950 269156 588874 269476
rect -4950 268216 588874 268536
rect -4950 262156 588874 262476
rect -4950 261216 588874 261536
rect -4950 255156 588874 255476
rect -4950 254216 588874 254536
rect -4950 248156 588874 248476
rect -4950 247216 588874 247536
rect -4950 241156 588874 241476
rect -4950 240216 588874 240536
rect -4950 234156 588874 234476
rect -4950 233216 588874 233536
rect -4950 227156 588874 227476
rect -4950 226216 588874 226536
rect -4950 220156 588874 220476
rect -4950 219216 588874 219536
rect -4950 213156 588874 213476
rect -4950 212216 588874 212536
rect -4950 206156 588874 206476
rect -4950 205216 588874 205536
rect -4950 199156 588874 199476
rect -4950 198216 588874 198536
rect -4950 192156 588874 192476
rect -4950 191216 588874 191536
rect -4950 185156 588874 185476
rect -4950 184216 588874 184536
rect -4950 178156 588874 178476
rect -4950 177216 588874 177536
rect -4950 171156 588874 171476
rect -4950 170216 588874 170536
rect -4950 164156 588874 164476
rect -4950 163216 588874 163536
rect -4950 157156 588874 157476
rect -4950 156216 588874 156536
rect -4950 150156 588874 150476
rect -4950 149216 588874 149536
rect -4950 143156 588874 143476
rect -4950 142216 588874 142536
rect -4950 136156 588874 136476
rect -4950 135216 588874 135536
rect -4950 129156 588874 129476
rect -4950 128216 588874 128536
rect -4950 122156 588874 122476
rect -4950 121216 588874 121536
rect -4950 115156 588874 115476
rect -4950 114216 588874 114536
rect -4950 108156 588874 108476
rect -4950 107216 588874 107536
rect -4950 101156 588874 101476
rect -4950 100216 588874 100536
rect -4950 94156 588874 94476
rect -4950 93216 588874 93536
rect -4950 87156 588874 87476
rect -4950 86216 588874 86536
rect -4950 80156 588874 80476
rect -4950 79216 588874 79536
rect -4950 73156 588874 73476
rect -4950 72216 588874 72536
rect -4950 66156 588874 66476
rect -4950 65216 588874 65536
rect -4950 59156 588874 59476
rect -4950 58216 588874 58536
rect -4950 52156 588874 52476
rect -4950 51216 588874 51536
rect -4950 45156 588874 45476
rect -4950 44216 588874 44536
rect -4950 38156 588874 38476
rect -4950 37216 588874 37536
rect -4950 31156 588874 31476
rect -4950 30216 588874 30536
rect -4950 24156 588874 24476
rect -4950 23216 588874 23536
rect -4950 17156 588874 17476
rect -4950 16216 588874 16536
rect -4950 10156 588874 10476
rect -4950 9216 588874 9536
rect -4950 3156 588874 3476
rect -4950 2216 588874 2536
rect -2406 -1334 587122 -714
rect -3366 -2294 587290 -1674
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal4 s -3198 -2126 -1786 706062 4 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -2406 -1334 587122 -714 8 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -2406 704650 587122 705270 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 585710 -2126 587122 706062 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 1144 -2294 1464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 8144 -2294 8464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 15144 -2294 15464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 22144 -2294 22464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 29144 -2294 29464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 36144 -2294 36464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 43144 -2294 43464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 50144 -2294 50464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 57144 -2294 57464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 64144 -2294 64464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 71144 -2294 71464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 78144 -2294 78464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 85144 -2294 85464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 92144 -2294 92464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 99144 -2294 99464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 106144 -2294 106464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 113144 -2294 113464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 120144 -2294 120464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 127144 -2294 127464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 134144 -2294 134464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 141144 -2294 141464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 148144 -2294 148464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 155144 -2294 155464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 162144 -2294 162464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 169144 -2294 169464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 176144 -2294 176464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 183144 -2294 183464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 190144 -2294 190464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 197144 -2294 197464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 204144 -2294 204464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 211144 -2294 211464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 218144 -2294 218464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 225144 -2294 225464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 232144 -2294 232464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 239144 -2294 239464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 246144 -2294 246464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 253144 -2294 253464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 260144 -2294 260464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 267144 -2294 267464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 274144 -2294 274464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 281144 -2294 281464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 288144 -2294 288464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 295144 -2294 295464 195976 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 295144 200380 295464 363976 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 295144 368380 295464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 302144 -2294 302464 195976 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 302144 200380 302464 363976 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 302144 368380 302464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 309144 -2294 309464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 316144 -2294 316464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 323144 -2294 323464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 330144 -2294 330464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 337144 -2294 337464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 344144 -2294 344464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 351144 -2294 351464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 358144 -2294 358464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 365144 -2294 365464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 372144 -2294 372464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 379144 -2294 379464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 386144 -2294 386464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 393144 -2294 393464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 400144 -2294 400464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 407144 -2294 407464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 414144 -2294 414464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 421144 -2294 421464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 428144 -2294 428464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 435144 -2294 435464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 442144 -2294 442464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 449144 -2294 449464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 456144 -2294 456464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 463144 -2294 463464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 470144 -2294 470464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 477144 -2294 477464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 484144 -2294 484464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 491144 -2294 491464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 498144 -2294 498464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 505144 -2294 505464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 512144 -2294 512464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 519144 -2294 519464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 526144 -2294 526464 240008 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 526144 261752 526464 280008 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 526144 301752 526464 320008 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 526144 341752 526464 360008 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 526144 381752 526464 400008 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 526144 421752 526464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 533144 -2294 533464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 540144 -2294 540464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 547144 -2294 547464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 554144 -2294 554464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 561144 -2294 561464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 568144 -2294 568464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 575144 -2294 575464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 582144 -2294 582464 706230 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 2216 588874 2536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 9216 588874 9536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 16216 588874 16536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 23216 588874 23536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 30216 588874 30536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 37216 588874 37536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 44216 588874 44536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 51216 588874 51536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 58216 588874 58536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 65216 588874 65536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 72216 588874 72536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 79216 588874 79536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 86216 588874 86536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 93216 588874 93536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 100216 588874 100536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 107216 588874 107536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 114216 588874 114536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 121216 588874 121536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 128216 588874 128536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 135216 588874 135536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 142216 588874 142536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 149216 588874 149536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 156216 588874 156536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 163216 588874 163536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 170216 588874 170536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 177216 588874 177536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 184216 588874 184536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 191216 588874 191536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 198216 588874 198536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 205216 588874 205536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 212216 588874 212536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 219216 588874 219536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 226216 588874 226536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 233216 588874 233536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 240216 588874 240536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 247216 588874 247536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 254216 588874 254536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 261216 588874 261536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 268216 588874 268536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 275216 588874 275536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 282216 588874 282536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 289216 588874 289536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 296216 588874 296536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 303216 588874 303536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 310216 588874 310536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 317216 588874 317536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 324216 588874 324536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 331216 588874 331536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 338216 588874 338536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 345216 588874 345536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 352216 588874 352536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 359216 588874 359536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 366216 588874 366536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 373216 588874 373536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 380216 588874 380536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 387216 588874 387536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 394216 588874 394536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 401216 588874 401536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 408216 588874 408536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 415216 588874 415536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 422216 588874 422536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 429216 588874 429536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 436216 588874 436536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 443216 588874 443536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 450216 588874 450536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 457216 588874 457536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 464216 588874 464536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 471216 588874 471536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 478216 588874 478536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 485216 588874 485536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 492216 588874 492536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 499216 588874 499536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 506216 588874 506536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 513216 588874 513536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 520216 588874 520536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 527216 588874 527536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 534216 588874 534536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 541216 588874 541536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 548216 588874 548536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 555216 588874 555536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 562216 588874 562536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 569216 588874 569536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 576216 588874 576536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 583216 588874 583536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 590216 588874 590536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 597216 588874 597536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 604216 588874 604536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 611216 588874 611536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 618216 588874 618536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 625216 588874 625536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 632216 588874 632536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 639216 588874 639536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 646216 588874 646536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 653216 588874 653536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 660216 588874 660536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 667216 588874 667536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 674216 588874 674536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 681216 588874 681536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 688216 588874 688536 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -4950 695216 588874 695536 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s -4950 -3878 -3538 707814 4 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3366 -2294 587290 -1674 8 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3366 705610 587290 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 587462 -3878 588874 707814 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 2876 -2294 3196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 9876 -2294 10196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 16876 -2294 17196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 23876 -2294 24196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 30876 -2294 31196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 37876 -2294 38196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 44876 -2294 45196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 51876 -2294 52196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 58876 -2294 59196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 65876 -2294 66196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 72876 -2294 73196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 79876 -2294 80196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 86876 -2294 87196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 93876 -2294 94196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 100876 -2294 101196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 107876 -2294 108196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 114876 -2294 115196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 121876 -2294 122196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 128876 -2294 129196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 135876 -2294 136196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 142876 -2294 143196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 149876 -2294 150196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 156876 -2294 157196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 163876 -2294 164196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 170876 -2294 171196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 177876 -2294 178196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 184876 -2294 185196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 191876 -2294 192196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 198876 -2294 199196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 205876 -2294 206196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 212876 -2294 213196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 219876 -2294 220196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 226876 -2294 227196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 233876 -2294 234196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 240876 -2294 241196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 247876 -2294 248196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 254876 -2294 255196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 261876 -2294 262196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 268876 -2294 269196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 275876 -2294 276196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 282876 -2294 283196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 289876 -2294 290196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 296876 -2294 297196 195976 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 296876 200380 297196 363976 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 296876 368380 297196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 303876 -2294 304196 195976 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 303876 200380 304196 363976 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 303876 368380 304196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 310876 -2294 311196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 317876 -2294 318196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 324876 -2294 325196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 331876 -2294 332196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 338876 -2294 339196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 345876 -2294 346196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 352876 -2294 353196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 359876 -2294 360196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 366876 -2294 367196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 373876 -2294 374196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 380876 -2294 381196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 387876 -2294 388196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 394876 -2294 395196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 401876 -2294 402196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 408876 -2294 409196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 415876 -2294 416196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 422876 -2294 423196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 429876 -2294 430196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 436876 -2294 437196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 443876 -2294 444196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 450876 -2294 451196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 457876 -2294 458196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 464876 -2294 465196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 471876 -2294 472196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 478876 -2294 479196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 485876 -2294 486196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 492876 -2294 493196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 499876 -2294 500196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 506876 -2294 507196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 513876 -2294 514196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 520876 -2294 521196 240008 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 520876 261752 521196 280008 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 520876 301752 521196 320008 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 520876 341752 521196 360008 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 520876 381752 521196 400008 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 520876 421752 521196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 527876 -2294 528196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 534876 -2294 535196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 541876 -2294 542196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 548876 -2294 549196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 555876 -2294 556196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 562876 -2294 563196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 569876 -2294 570196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 576876 -2294 577196 706230 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 3156 588874 3476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 10156 588874 10476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 17156 588874 17476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 24156 588874 24476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 31156 588874 31476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 38156 588874 38476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 45156 588874 45476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 52156 588874 52476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 59156 588874 59476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 66156 588874 66476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 73156 588874 73476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 80156 588874 80476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 87156 588874 87476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 94156 588874 94476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 101156 588874 101476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 108156 588874 108476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 115156 588874 115476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 122156 588874 122476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 129156 588874 129476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 136156 588874 136476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 143156 588874 143476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 150156 588874 150476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 157156 588874 157476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 164156 588874 164476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 171156 588874 171476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 178156 588874 178476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 185156 588874 185476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 192156 588874 192476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 199156 588874 199476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 206156 588874 206476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 213156 588874 213476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 220156 588874 220476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 227156 588874 227476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 234156 588874 234476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 241156 588874 241476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 248156 588874 248476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 255156 588874 255476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 262156 588874 262476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 269156 588874 269476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 276156 588874 276476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 283156 588874 283476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 290156 588874 290476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 297156 588874 297476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 304156 588874 304476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 311156 588874 311476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 318156 588874 318476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 325156 588874 325476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 332156 588874 332476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 339156 588874 339476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 346156 588874 346476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 353156 588874 353476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 360156 588874 360476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 367156 588874 367476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 374156 588874 374476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 381156 588874 381476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 388156 588874 388476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 395156 588874 395476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 402156 588874 402476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 409156 588874 409476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 416156 588874 416476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 423156 588874 423476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 430156 588874 430476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 437156 588874 437476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 444156 588874 444476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 451156 588874 451476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 458156 588874 458476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 465156 588874 465476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 472156 588874 472476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 479156 588874 479476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 486156 588874 486476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 493156 588874 493476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 500156 588874 500476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 507156 588874 507476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 514156 588874 514476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 521156 588874 521476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 528156 588874 528476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 535156 588874 535476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 542156 588874 542476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 549156 588874 549476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 556156 588874 556476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 563156 588874 563476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 570156 588874 570476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 577156 588874 577476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 584156 588874 584476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 591156 588874 591476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 598156 588874 598476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 605156 588874 605476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 612156 588874 612476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 619156 588874 619476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 626156 588874 626476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 633156 588874 633476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 640156 588874 640476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 647156 588874 647476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 654156 588874 654476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 661156 588874 661476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 668156 588874 668476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 675156 588874 675476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 682156 588874 682476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 689156 588874 689476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -4950 696156 588874 696476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 146 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 147 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 148 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 149 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 150 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 151 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 152 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 153 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 154 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 155 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 156 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 157 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 158 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 159 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 160 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 161 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 162 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 163 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 164 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 165 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 166 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 167 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 168 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 169 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 170 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 171 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 172 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 173 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 174 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 175 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 176 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 177 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 178 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 179 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 180 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 181 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 182 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 183 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 184 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 185 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 186 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 187 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 188 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 189 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 190 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 191 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 192 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 193 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 194 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 195 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 196 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 197 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 198 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 199 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 200 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 201 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 202 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 203 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 204 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 205 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 206 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 207 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 208 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 209 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 210 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 211 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 212 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 213 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 214 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 215 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 216 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 217 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 218 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 219 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 220 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 221 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 222 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 223 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 224 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 225 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 226 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 227 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 228 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 229 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 230 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 231 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 232 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 233 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 234 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 235 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 236 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 237 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 238 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 239 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 240 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 241 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 242 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 243 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 244 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 245 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 246 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 247 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 248 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 249 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 250 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 251 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2644206
string GDS_FILE /import/yukari1/lrburle/google_ring_oscillator/caravel/openlane/user_project_wrapper/runs/23_12_19_10_44/results/signoff/user_project_wrapper.magic.gds
string GDS_START 1096046
<< end >>

