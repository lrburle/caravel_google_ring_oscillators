magic
tech sky130A
magscale 1 2
timestamp 1604095905
<< checkpaint >>
rect -1269 2461 1439 2601
rect -1760 -1129 6260 2461
rect -1269 -1260 1439 -1129
<< nwell >>
rect -9 485 179 897
<< locali >>
rect 0 827 176 888
rect 0 0 176 61
<< metal1 >>
rect 0 827 176 888
rect 0 0 176 61
<< labels >>
rlabel metal1 111 859 111 859 1 vccd1
rlabel metal1 112 28 112 28 1 vssd1
<< end >>
