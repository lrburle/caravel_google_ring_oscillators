magic
tech sky130A
magscale 1 2
timestamp 1716047795
<< nwell >>
rect 3000 1019 5943 1749
rect 6909 1730 7316 1751
rect 10618 1729 11025 1750
rect 14463 1741 14720 1750
rect 18132 1730 18444 1750
rect 8908 1635 8966 1693
rect 12620 1635 12678 1693
rect 16332 1635 16390 1693
rect 20044 1635 20102 1693
rect 7251 1407 7288 1408
rect 10955 1406 10986 1408
rect 14675 1407 14708 1408
rect 18387 1407 18410 1408
rect 3000 820 4966 1019
rect 7151 986 7209 1044
rect 10863 986 10921 1044
rect 14575 986 14633 1044
rect 18287 986 18345 1044
rect 21999 986 22057 1044
rect 7271 819 7424 820
rect 10983 819 11136 820
rect 14695 819 14848 820
rect 18407 819 18560 820
<< ndiff >>
rect 7162 442 7197 476
rect 10874 442 10909 476
rect 14586 442 14621 476
rect 18298 442 18333 476
rect 22010 442 22045 476
rect 7162 441 7196 442
rect 10874 441 10908 442
rect 14586 441 14620 442
rect 18298 441 18332 442
rect 22010 441 22044 442
<< pdiff >>
rect 3045 1648 3079 1682
rect 5209 1647 5243 1681
rect 8908 1635 8966 1693
rect 12620 1635 12678 1693
rect 16332 1635 16390 1693
rect 20044 1635 20102 1693
<< locali >>
rect 0 2173 22120 2493
rect 9055 1756 9079 1758
rect 3406 1408 3440 1479
rect 0 1088 22099 1408
rect 0 0 22119 320
<< viali >>
rect 3045 1648 3079 1682
rect 7163 442 7197 476
rect 10875 442 10909 476
rect 14587 442 14621 476
rect 18299 442 18333 476
rect 22011 442 22045 476
<< metal1 >>
rect 0 2173 22120 2493
rect 22040 2010 22046 2013
rect 22005 2000 22058 2010
rect 22005 1983 22070 2000
rect 22005 1977 22075 1983
rect 3302 1864 3308 1922
rect 3366 1864 3372 1922
rect 22005 1919 22011 1977
rect 22069 1919 22075 1977
rect 22005 1913 22075 1919
rect 7161 1853 7231 1859
rect 5598 1843 5668 1849
rect 5598 1785 5604 1843
rect 5662 1785 5668 1843
rect 5598 1779 5668 1785
rect 7161 1795 7167 1853
rect 7225 1795 7231 1853
rect 10872 1854 10943 1861
rect 7161 1789 7231 1795
rect 9310 1844 9380 1850
rect 3227 1715 3233 1773
rect 3291 1715 3297 1773
rect 7161 1771 7221 1789
rect 9310 1786 9316 1844
rect 9374 1786 9380 1844
rect 9310 1780 9380 1786
rect 10872 1796 10879 1854
rect 10937 1796 10943 1854
rect 14576 1853 14646 1859
rect 10872 1790 10943 1796
rect 13021 1845 13091 1851
rect 10872 1770 10933 1790
rect 13021 1787 13027 1845
rect 13085 1787 13091 1845
rect 13021 1781 13091 1787
rect 14576 1795 14582 1853
rect 14640 1795 14646 1853
rect 18288 1853 18358 1859
rect 14576 1789 14646 1795
rect 16733 1844 16803 1850
rect 14576 1771 14645 1789
rect 16733 1786 16739 1844
rect 16797 1786 16803 1844
rect 16733 1780 16803 1786
rect 18288 1795 18294 1853
rect 18352 1795 18358 1853
rect 18288 1789 18358 1795
rect 20445 1844 20515 1850
rect 18288 1771 18357 1789
rect 20445 1786 20451 1844
rect 20509 1786 20515 1844
rect 20445 1780 20515 1786
rect 5343 1756 5377 1758
rect 9055 1756 9079 1758
rect 12767 1756 12796 1758
rect 16479 1756 16511 1758
rect 20191 1756 20227 1758
rect 3028 1682 3096 1691
rect 3028 1648 3045 1682
rect 3079 1648 3096 1682
rect 3028 1639 3096 1648
rect 5196 1635 5254 1693
rect 8908 1635 8966 1693
rect 12620 1635 12678 1693
rect 16332 1635 16390 1693
rect 20044 1635 20102 1693
rect 0 1088 22099 1408
rect 7162 441 7196 442
rect 10874 441 10908 442
rect 14586 441 14620 442
rect 18298 441 18332 442
rect 22010 441 22044 442
rect 0 0 22119 320
<< via1 >>
rect 3308 1864 3366 1922
rect 22011 1919 22069 1977
rect 5604 1785 5662 1843
rect 7167 1795 7225 1853
rect 3233 1715 3291 1773
rect 9316 1786 9374 1844
rect 10879 1796 10937 1854
rect 13027 1787 13085 1845
rect 14582 1795 14640 1853
rect 16739 1786 16797 1844
rect 18294 1795 18352 1853
rect 20451 1786 20509 1844
<< metal2 >>
rect 3245 2138 22045 2172
rect 3245 1779 3279 2138
rect 22011 1983 22045 2138
rect 22005 1977 22075 1983
rect 3308 1922 3366 1928
rect 22005 1919 22011 1977
rect 22069 1919 22075 1977
rect 22005 1913 22075 1919
rect 3366 1903 3372 1904
rect 3366 1869 3546 1903
rect 3308 1858 3366 1864
rect 3512 1829 3546 1869
rect 7161 1853 7231 1859
rect 5598 1843 5668 1849
rect 5598 1829 5604 1843
rect 3512 1795 5604 1829
rect 5598 1785 5604 1795
rect 5662 1785 5668 1843
rect 7161 1795 7167 1853
rect 7225 1835 7231 1853
rect 10873 1854 10943 1860
rect 9310 1844 9380 1850
rect 9310 1835 9316 1844
rect 7225 1795 9316 1835
rect 7161 1789 7231 1795
rect 5598 1779 5668 1785
rect 9310 1786 9316 1795
rect 9374 1786 9380 1844
rect 10873 1796 10879 1854
rect 10937 1836 10943 1854
rect 14576 1853 14646 1859
rect 13021 1845 13091 1851
rect 13021 1836 13027 1845
rect 10937 1796 13027 1836
rect 10873 1790 10943 1796
rect 9310 1780 9380 1786
rect 13021 1787 13027 1796
rect 13085 1787 13091 1845
rect 14576 1795 14582 1853
rect 14640 1835 14646 1853
rect 18288 1853 18358 1859
rect 16733 1844 16803 1850
rect 16733 1835 16739 1844
rect 14640 1795 16739 1835
rect 14576 1789 14646 1795
rect 13021 1781 13091 1787
rect 16733 1786 16739 1795
rect 16797 1786 16803 1844
rect 18288 1795 18294 1853
rect 18352 1835 18358 1853
rect 20445 1844 20515 1850
rect 20445 1835 20451 1844
rect 18352 1795 20451 1835
rect 18288 1789 18358 1795
rect 16733 1780 16803 1786
rect 20445 1786 20451 1795
rect 20509 1786 20515 1844
rect 20445 1780 20515 1786
rect 3233 1773 3291 1779
rect 3233 1709 3291 1715
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1714057206
transform 1 0 3009 0 -1 2234
box -10 0 552 902
use sky130_osu_single_mpr2et_8_b0r2  sky130_osu_single_mpr2et_8_b0r2_0
timestamp 1716047795
transform 1 0 18406 0 1 0
box 0 0 3714 2493
use sky130_osu_single_mpr2et_8_b0r2  sky130_osu_single_mpr2et_8_b0r2_1
timestamp 1716047795
transform 1 0 3558 0 1 0
box 0 0 3714 2493
use sky130_osu_single_mpr2et_8_b0r2  sky130_osu_single_mpr2et_8_b0r2_2
timestamp 1716047795
transform 1 0 7270 0 1 0
box 0 0 3714 2493
use sky130_osu_single_mpr2et_8_b0r2  sky130_osu_single_mpr2et_8_b0r2_3
timestamp 1716047795
transform 1 0 10982 0 1 0
box 0 0 3714 2493
use sky130_osu_single_mpr2et_8_b0r2  sky130_osu_single_mpr2et_8_b0r2_4
timestamp 1716047795
transform 1 0 14694 0 1 0
box 0 0 3714 2493
<< labels >>
flabel metal1 s 3032 1641 3092 1687 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel metal1 s 0 2173 22120 2493 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal1 s 0 1088 22099 1408 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 0 0 22119 320 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel viali s 5208 1648 5242 1682 0 FreeSans 100 0 0 0 s1
port 1 nw signal input
flabel viali s 8920 1648 8954 1682 0 FreeSans 100 0 0 0 s2
port 2 nw signal input
flabel viali s 12632 1648 12666 1682 0 FreeSans 100 0 0 0 s3
port 3 nw signal input
flabel viali s 16344 1648 16378 1682 0 FreeSans 100 0 0 0 s4
port 4 nw signal input
flabel viali s 20056 1648 20090 1682 0 FreeSans 100 0 0 0 s5
port 5 nw signal input
flabel viali s 22011 442 22045 476 0 FreeSans 100 0 0 0 X5_Y1
port 10 se signal output
flabel viali s 18299 442 18333 476 0 FreeSans 100 0 0 0 X4_Y1
port 9 se signal output
flabel viali s 14587 442 14621 476 0 FreeSans 100 0 0 0 X3_Y1
port 8 se signal output
flabel viali s 10875 442 10909 476 0 FreeSans 100 0 0 0 X2_Y1
port 7 se signal output
flabel viali s 7163 442 7197 476 0 FreeSans 100 0 0 0 X1_Y1
port 6 se signal output
<< end >>
