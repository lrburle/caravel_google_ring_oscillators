magic
tech sky130A
magscale 1 2
timestamp 1710268143
<< checkpaint >>
rect -12658 -11586 596582 715522
<< viali >>
rect 481557 432429 481591 432463
rect 473362 411417 473396 411451
rect 478581 410057 478615 410091
rect 485111 410057 485145 410091
rect 473809 390473 473843 390507
rect 479474 389045 479508 389079
rect 475138 369461 475172 369495
rect 477091 367965 477125 367999
rect 475441 347021 475475 347055
rect 478758 347021 478792 347055
rect 482075 347021 482109 347055
rect 478938 326009 478972 326043
rect 473361 306425 473395 306459
rect 478580 305473 478614 305507
rect 485110 305473 485144 305507
rect 479474 284053 479508 284087
rect 477101 263041 477135 263075
rect 544117 212789 544151 212823
<< metal1 >>
rect 470234 451485 470854 451491
rect 470234 451177 470262 451485
rect 470826 451177 470854 451485
rect 470234 451171 470854 451177
rect 471330 450644 471336 450696
rect 471388 450684 471394 450696
rect 471388 450656 471652 450684
rect 471388 450644 471394 450656
rect 468994 450399 469614 450405
rect 468994 450091 469022 450399
rect 469586 450091 469614 450399
rect 468994 450085 469614 450091
rect 488258 450004 488264 450016
rect 484504 449936 484532 449990
rect 487830 449976 488264 450004
rect 488258 449964 488264 449976
rect 488316 449964 488322 450016
rect 484504 449908 485774 449936
rect 485746 449868 485774 449908
rect 488994 449868 489000 449880
rect 485746 449840 487752 449868
rect 487724 449732 487752 449840
rect 488276 449840 489000 449868
rect 488276 449732 488304 449840
rect 488994 449828 489000 449840
rect 489052 449828 489058 449880
rect 487724 449704 488304 449732
rect 475384 449485 475436 449491
rect 475384 449427 475436 449433
rect 478696 449485 478748 449491
rect 478696 449427 478748 449433
rect 482008 449485 482060 449491
rect 482008 449427 482060 449433
rect 485320 449485 485372 449491
rect 488810 449473 488816 449485
rect 488658 449445 488816 449473
rect 488810 449433 488816 449445
rect 488868 449433 488874 449485
rect 485320 449427 485372 449433
rect 470234 449314 470854 449320
rect 470234 449006 470262 449314
rect 470826 449006 470854 449314
rect 470234 449000 470854 449006
rect 544562 445136 544568 445188
rect 544620 445176 544626 445188
rect 547874 445176 547880 445188
rect 544620 445148 547880 445176
rect 544620 445136 544626 445148
rect 547874 445136 547880 445148
rect 547932 445136 547938 445188
rect 493502 434732 493508 434784
rect 493560 434772 493566 434784
rect 535454 434772 535460 434784
rect 493560 434744 535460 434772
rect 493560 434732 493566 434744
rect 535454 434732 535460 434744
rect 535512 434732 535518 434784
rect 470234 433086 470854 433092
rect 470234 432778 470262 433086
rect 470826 432778 470854 433086
rect 470234 432772 470854 432778
rect 481542 432692 481548 432744
rect 481600 432692 481606 432744
rect 483106 432692 483112 432744
rect 483164 432692 483170 432744
rect 481560 432469 481588 432692
rect 481545 432463 481603 432469
rect 481545 432429 481557 432463
rect 481591 432429 481603 432463
rect 481545 432423 481603 432429
rect 483124 432392 483152 432692
rect 482940 432364 483152 432392
rect 471612 432290 471664 432296
rect 482940 432278 482968 432364
rect 471612 432232 471664 432238
rect 471790 432216 471796 432268
rect 471848 432256 471854 432268
rect 472084 432256 472374 432278
rect 471848 432250 472374 432256
rect 482678 432250 482968 432278
rect 483124 432278 483152 432364
rect 483124 432250 483157 432278
rect 471848 432228 472112 432250
rect 471848 432216 471854 432228
rect 483129 432188 483157 432250
rect 483124 432160 483157 432188
rect 483124 432132 483152 432160
rect 483106 432080 483112 432132
rect 483164 432080 483170 432132
rect 468994 431999 469614 432005
rect 468994 431691 469022 431999
rect 469586 431691 469614 431999
rect 468994 431685 469614 431691
rect 489638 431440 489644 431452
rect 477954 431128 477960 431180
rect 478012 431168 478018 431180
rect 478156 431168 478184 431428
rect 488460 431412 489644 431440
rect 489638 431400 489644 431412
rect 489696 431400 489702 431452
rect 478012 431140 478184 431168
rect 478012 431128 478018 431140
rect 470234 430914 470854 430920
rect 470234 430606 470262 430914
rect 470826 430606 470854 430914
rect 470234 430600 470854 430606
rect 470234 412086 470854 412092
rect 470234 411778 470262 412086
rect 470826 411778 470854 412086
rect 470234 411772 470854 411778
rect 471606 411544 471612 411596
rect 471664 411584 471670 411596
rect 471664 411556 473400 411584
rect 471664 411544 471670 411556
rect 473372 411457 473400 411556
rect 473350 411451 473408 411457
rect 473350 411417 473362 411451
rect 473396 411417 473408 411451
rect 473350 411411 473408 411417
rect 471238 411272 471244 411324
rect 471296 411277 471302 411324
rect 471296 411272 471638 411277
rect 471256 411249 471638 411272
rect 468994 411000 469614 411006
rect 468994 410692 469022 411000
rect 469586 410692 469614 411000
rect 468994 410686 469614 410692
rect 488534 410496 488540 410508
rect 487724 410468 488540 410496
rect 487724 410428 487752 410468
rect 488534 410456 488540 410468
rect 488592 410496 488598 410508
rect 489086 410496 489092 410508
rect 488592 410468 489092 410496
rect 488592 410456 488598 410468
rect 489086 410456 489092 410468
rect 489144 410456 489150 410508
rect 487554 410400 487752 410428
rect 478569 410091 478627 410097
rect 475292 410085 475344 410091
rect 478569 410057 478581 410091
rect 478615 410088 478627 410091
rect 478690 410088 478696 410100
rect 478615 410060 478696 410088
rect 478615 410057 478627 410060
rect 478569 410051 478627 410057
rect 478690 410048 478696 410060
rect 478748 410048 478754 410100
rect 485099 410091 485157 410097
rect 481824 410085 481876 410091
rect 475292 410027 475344 410033
rect 485099 410057 485111 410091
rect 485145 410088 485157 410091
rect 485222 410088 485228 410100
rect 485145 410060 485228 410088
rect 485145 410057 485157 410060
rect 485099 410051 485157 410057
rect 485222 410048 485228 410060
rect 485280 410048 485286 410100
rect 488534 410073 488540 410085
rect 488382 410045 488540 410073
rect 488534 410033 488540 410045
rect 488592 410033 488598 410085
rect 481824 410027 481876 410033
rect 470234 409914 470854 409920
rect 470234 409606 470262 409914
rect 470826 409606 470854 409914
rect 470234 409600 470854 409606
rect 544654 409164 544660 409216
rect 544712 409204 544718 409216
rect 547874 409204 547880 409216
rect 544712 409176 547880 409204
rect 544712 409164 544718 409176
rect 547874 409164 547880 409176
rect 547932 409164 547938 409216
rect 488534 407736 488540 407788
rect 488592 407776 488598 407788
rect 489454 407776 489460 407788
rect 488592 407748 489460 407776
rect 488592 407736 488598 407748
rect 489454 407736 489460 407748
rect 489512 407736 489518 407788
rect 470234 391087 470854 391093
rect 470234 390779 470262 391087
rect 470826 390779 470854 391087
rect 470234 390773 470854 390779
rect 471698 390464 471704 390516
rect 471756 390504 471762 390516
rect 473797 390507 473855 390513
rect 473797 390504 473809 390507
rect 471756 390476 473809 390504
rect 471756 390464 471762 390476
rect 473797 390473 473809 390476
rect 473843 390473 473855 390507
rect 473797 390467 473855 390473
rect 471514 390238 471520 390290
rect 471572 390278 471578 390290
rect 471572 390264 471638 390278
rect 471572 390250 471652 390264
rect 471572 390238 471578 390250
rect 471624 390096 471652 390250
rect 478046 390238 478052 390290
rect 478104 390238 478110 390290
rect 471698 390096 471704 390108
rect 471624 390068 471704 390096
rect 471698 390056 471704 390068
rect 471756 390056 471762 390108
rect 468994 390004 469614 390010
rect 468994 389696 469022 390004
rect 469586 389696 469614 390004
rect 468994 389690 469614 389696
rect 487172 389592 489914 389620
rect 487172 389552 487200 389592
rect 486068 389524 487200 389552
rect 489886 389552 489914 389592
rect 490834 389552 490840 389564
rect 489886 389524 490840 389552
rect 486068 389470 486096 389524
rect 490834 389512 490840 389524
rect 490892 389512 490898 389564
rect 475752 389085 475804 389091
rect 479462 389079 479520 389085
rect 479462 389045 479474 389079
rect 479508 389076 479520 389079
rect 479610 389076 479616 389088
rect 479508 389048 479616 389076
rect 479508 389045 479520 389048
rect 479462 389039 479520 389045
rect 479610 389036 479616 389048
rect 479668 389036 479674 389088
rect 483204 389085 483256 389091
rect 475752 389027 475804 389033
rect 483204 389027 483256 389033
rect 486884 389085 486936 389091
rect 486884 389027 486936 389033
rect 470234 388914 470854 388920
rect 470234 388606 470262 388914
rect 470826 388606 470854 388914
rect 470234 388600 470854 388606
rect 545022 373192 545028 373244
rect 545080 373232 545086 373244
rect 548518 373232 548524 373244
rect 545080 373204 548524 373232
rect 545080 373192 545086 373204
rect 548518 373192 548524 373204
rect 548576 373192 548582 373244
rect 470234 370087 470854 370093
rect 470234 369779 470262 370087
rect 470826 369779 470854 370087
rect 470234 369773 470854 369779
rect 473722 369452 473728 369504
rect 473780 369492 473786 369504
rect 475126 369495 475184 369501
rect 475126 369492 475138 369495
rect 473780 369464 475138 369492
rect 473780 369452 473786 369464
rect 475126 369461 475138 369464
rect 475172 369461 475184 369495
rect 475126 369455 475184 369461
rect 471698 369316 471704 369368
rect 471756 369356 471762 369368
rect 471756 369328 473676 369356
rect 471756 369316 471762 369328
rect 473648 369265 473676 369328
rect 481272 369290 481324 369296
rect 478874 369238 478880 369290
rect 478932 369238 478938 369290
rect 488902 369288 488908 369300
rect 488474 369260 488908 369288
rect 488902 369248 488908 369260
rect 488960 369288 488966 369300
rect 489822 369288 489828 369300
rect 488960 369260 489828 369288
rect 488960 369248 488966 369260
rect 489822 369248 489828 369260
rect 489880 369248 489886 369300
rect 481272 369232 481324 369238
rect 473906 369112 473912 369164
rect 473964 369152 473970 369164
rect 481266 369152 481272 369164
rect 473964 369124 481272 369152
rect 473964 369112 473970 369124
rect 481266 369112 481272 369124
rect 481324 369152 481330 369164
rect 481818 369152 481824 369164
rect 481324 369124 481824 369152
rect 481324 369112 481330 369124
rect 481818 369112 481824 369124
rect 481876 369112 481882 369164
rect 468994 369001 469614 369007
rect 468994 368693 469022 369001
rect 469586 368693 469614 369001
rect 468994 368687 469614 368693
rect 485314 368568 485320 368620
rect 485372 368608 485378 368620
rect 485372 368580 485452 368608
rect 485372 368568 485378 368580
rect 485424 368540 485452 368580
rect 489638 368540 489644 368552
rect 485424 368512 489644 368540
rect 485424 368458 485452 368512
rect 489638 368500 489644 368512
rect 489696 368500 489702 368552
rect 489454 368072 489460 368084
rect 489302 368044 489460 368072
rect 489454 368032 489460 368044
rect 489512 368032 489518 368084
rect 477079 367999 477137 368005
rect 477079 367965 477091 367999
rect 477125 367996 477137 367999
rect 477218 367996 477224 368008
rect 477125 367968 477224 367996
rect 477125 367965 477137 367968
rect 477079 367959 477137 367965
rect 477218 367956 477224 367968
rect 477276 367956 477282 368008
rect 470234 367914 470854 367920
rect 470234 367606 470262 367914
rect 470826 367606 470854 367914
rect 470234 367600 470854 367606
rect 490558 363604 490564 363656
rect 490616 363644 490622 363656
rect 536190 363644 536196 363656
rect 490616 363616 536196 363644
rect 490616 363604 490622 363616
rect 536190 363604 536196 363616
rect 536248 363604 536254 363656
rect 470234 349086 470854 349092
rect 470234 348778 470262 349086
rect 470826 348778 470854 349086
rect 470234 348772 470854 348778
rect 475654 348508 475660 348560
rect 475712 348508 475718 348560
rect 471606 348440 471612 348492
rect 471664 348480 471670 348492
rect 471664 348452 471744 348480
rect 471664 348440 471670 348452
rect 471716 348263 471744 348452
rect 475672 348344 475700 348508
rect 475580 348316 475700 348344
rect 475580 348276 475608 348316
rect 487922 348276 488028 348279
rect 489086 348276 489092 348288
rect 475396 348248 475686 348276
rect 487922 348251 489092 348276
rect 488000 348248 489092 348251
rect 471790 348100 471796 348152
rect 471848 348140 471854 348152
rect 475396 348140 475424 348248
rect 489086 348236 489092 348248
rect 489144 348236 489150 348288
rect 471848 348112 473216 348140
rect 471848 348100 471854 348112
rect 468994 347999 469614 348005
rect 468994 347691 469022 347999
rect 469586 347691 469614 347999
rect 473188 347936 473216 348112
rect 473832 348112 475424 348140
rect 473832 347936 473860 348112
rect 473188 347908 473860 347936
rect 468994 347685 469614 347691
rect 484780 347445 487752 347460
rect 484610 347432 487752 347445
rect 484610 347417 484808 347432
rect 487724 347324 487752 347432
rect 488534 347324 488540 347336
rect 487724 347296 488540 347324
rect 488534 347284 488540 347296
rect 488592 347284 488598 347336
rect 485412 347087 485464 347093
rect 475429 347055 475487 347061
rect 475429 347021 475441 347055
rect 475475 347052 475487 347055
rect 475562 347052 475568 347064
rect 475475 347024 475568 347052
rect 475475 347021 475487 347024
rect 475429 347015 475487 347021
rect 475562 347012 475568 347024
rect 475620 347012 475626 347064
rect 478598 347012 478604 347064
rect 478656 347052 478662 347064
rect 478746 347055 478804 347061
rect 478746 347052 478758 347055
rect 478656 347024 478758 347052
rect 478656 347012 478662 347024
rect 478746 347021 478758 347024
rect 478792 347021 478804 347055
rect 478746 347015 478804 347021
rect 482063 347055 482121 347061
rect 482063 347021 482075 347055
rect 482109 347052 482121 347055
rect 482186 347052 482192 347064
rect 482109 347024 482192 347052
rect 482109 347021 482121 347024
rect 482063 347015 482121 347021
rect 482186 347012 482192 347024
rect 482244 347012 482250 347064
rect 488750 347052 488948 347075
rect 488994 347052 489000 347064
rect 488750 347047 489000 347052
rect 485412 347029 485464 347035
rect 488920 347024 489000 347047
rect 488994 347012 489000 347024
rect 489052 347012 489058 347064
rect 470234 346914 470854 346920
rect 470234 346606 470262 346914
rect 470826 346606 470854 346914
rect 470234 346600 470854 346606
rect 485406 328176 485412 328228
rect 485464 328216 485470 328228
rect 488810 328216 488816 328228
rect 485464 328188 488816 328216
rect 485464 328176 485470 328188
rect 488810 328176 488816 328188
rect 488868 328216 488874 328228
rect 489730 328216 489736 328228
rect 488868 328188 489736 328216
rect 488868 328176 488874 328188
rect 489730 328176 489736 328188
rect 489788 328176 489794 328228
rect 470234 328086 470854 328092
rect 470234 327778 470262 328086
rect 470826 327778 470854 328086
rect 470234 327772 470854 327778
rect 471238 327292 471244 327344
rect 471296 327332 471302 327344
rect 471296 327304 471652 327332
rect 471296 327292 471302 327304
rect 471624 327264 471652 327304
rect 468994 326999 469614 327005
rect 468994 326691 469022 326999
rect 469586 326691 469614 326999
rect 468994 326685 469614 326691
rect 489546 326448 489552 326460
rect 488552 326442 489552 326448
rect 488474 326420 489552 326442
rect 488474 326414 488580 326420
rect 489546 326408 489552 326420
rect 489604 326408 489610 326460
rect 536282 326448 536288 326460
rect 495406 326420 536288 326448
rect 489362 326340 489368 326392
rect 489420 326380 489426 326392
rect 495406 326380 495434 326420
rect 536282 326408 536288 326420
rect 536340 326408 536346 326460
rect 489420 326352 495434 326380
rect 489420 326340 489426 326352
rect 478926 326043 478984 326049
rect 478926 326009 478938 326043
rect 478972 326040 478984 326043
rect 479058 326040 479064 326052
rect 478972 326012 479064 326040
rect 478972 326009 478984 326012
rect 478926 326003 478984 326009
rect 479058 326000 479064 326012
rect 479116 326000 479122 326052
rect 489288 326040 489316 326058
rect 492030 326040 492036 326052
rect 489288 326012 492036 326040
rect 492030 326000 492036 326012
rect 492088 326000 492094 326052
rect 470234 325914 470854 325920
rect 470234 325606 470262 325914
rect 470826 325606 470854 325914
rect 470234 325600 470854 325606
rect 470234 307086 470854 307092
rect 470234 306778 470262 307086
rect 470826 306778 470854 307086
rect 470234 306772 470854 306778
rect 471698 306484 471704 306536
rect 471756 306524 471762 306536
rect 471756 306496 473400 306524
rect 471756 306484 471762 306496
rect 473372 306465 473400 306496
rect 473349 306459 473407 306465
rect 473349 306425 473361 306459
rect 473395 306425 473407 306459
rect 473349 306419 473407 306425
rect 471238 306280 471244 306332
rect 471296 306320 471302 306332
rect 471296 306292 471652 306320
rect 471296 306280 471302 306292
rect 471624 306264 471652 306292
rect 468994 306001 469614 306007
rect 468994 305693 469022 306001
rect 469586 305693 469614 306001
rect 468994 305687 469614 305693
rect 478598 305513 478604 305516
rect 478568 305507 478604 305513
rect 478568 305473 478580 305507
rect 478568 305467 478604 305473
rect 478598 305464 478604 305467
rect 478656 305464 478662 305516
rect 485130 305513 485136 305516
rect 485098 305507 485136 305513
rect 485098 305473 485110 305507
rect 485098 305467 485136 305473
rect 485130 305464 485136 305467
rect 485188 305464 485194 305516
rect 489270 305436 489276 305448
rect 487554 305408 489276 305436
rect 489270 305396 489276 305408
rect 489328 305396 489334 305448
rect 475292 305085 475344 305091
rect 475292 305027 475344 305033
rect 481824 305085 481876 305091
rect 488382 305045 488672 305073
rect 481824 305027 481876 305033
rect 488644 305028 488672 305045
rect 490650 305028 490656 305040
rect 488644 305000 490656 305028
rect 490650 304988 490656 305000
rect 490708 304988 490714 305040
rect 470234 304914 470854 304920
rect 470234 304606 470262 304914
rect 470826 304606 470854 304914
rect 470234 304600 470854 304606
rect 478524 303640 478736 303668
rect 475286 303560 475292 303612
rect 475344 303600 475350 303612
rect 478524 303600 478552 303640
rect 475344 303572 478552 303600
rect 475344 303560 475350 303572
rect 478598 303560 478604 303612
rect 478656 303560 478662 303612
rect 478616 303464 478644 303560
rect 478708 303532 478736 303640
rect 485130 303560 485136 303612
rect 485188 303600 485194 303612
rect 536374 303600 536380 303612
rect 485188 303572 536380 303600
rect 485188 303560 485194 303572
rect 536374 303560 536380 303572
rect 536432 303560 536438 303612
rect 493502 303532 493508 303544
rect 478708 303504 493508 303532
rect 493502 303492 493508 303504
rect 493560 303492 493566 303544
rect 490558 303464 490564 303476
rect 478616 303436 490564 303464
rect 490558 303424 490564 303436
rect 490616 303424 490622 303476
rect 481818 303356 481824 303408
rect 481876 303396 481882 303408
rect 489178 303396 489184 303408
rect 481876 303368 489184 303396
rect 481876 303356 481882 303368
rect 489178 303356 489184 303368
rect 489236 303356 489242 303408
rect 490650 292476 490656 292528
rect 490708 292516 490714 292528
rect 535454 292516 535460 292528
rect 490708 292488 535460 292516
rect 490708 292476 490714 292488
rect 535454 292476 535460 292488
rect 535512 292476 535518 292528
rect 470234 286087 470854 286093
rect 470234 285779 470262 286087
rect 470826 285779 470854 286087
rect 470234 285773 470854 285779
rect 471422 285239 471428 285291
rect 471480 285279 471486 285291
rect 471480 285265 471638 285279
rect 471480 285251 471652 285265
rect 471480 285239 471486 285251
rect 471624 285104 471652 285251
rect 478046 285238 478052 285290
rect 478104 285238 478110 285290
rect 486071 285240 486099 285278
rect 486068 285212 486099 285240
rect 489270 285238 489276 285290
rect 489328 285238 489334 285290
rect 486068 285172 486096 285212
rect 491386 285172 491392 285184
rect 486068 285144 491392 285172
rect 491386 285132 491392 285144
rect 491444 285132 491450 285184
rect 471698 285104 471704 285116
rect 471624 285076 471704 285104
rect 471698 285064 471704 285076
rect 471756 285064 471762 285116
rect 468994 285002 469614 285008
rect 468994 284694 469022 285002
rect 469586 284694 469614 285002
rect 468994 284688 469614 284694
rect 475752 284085 475804 284091
rect 479462 284087 479520 284093
rect 479462 284053 479474 284087
rect 479508 284084 479520 284087
rect 479610 284084 479616 284096
rect 479508 284056 479616 284084
rect 479508 284053 479520 284056
rect 479462 284047 479520 284053
rect 479610 284044 479616 284056
rect 479668 284044 479674 284096
rect 483204 284085 483256 284091
rect 475752 284027 475804 284033
rect 483204 284027 483256 284033
rect 486884 284085 486936 284091
rect 486884 284027 486936 284033
rect 470234 283914 470854 283920
rect 470234 283606 470262 283914
rect 470826 283606 470854 283914
rect 470234 283600 470854 283606
rect 471698 266364 471704 266416
rect 471756 266404 471762 266416
rect 473722 266404 473728 266416
rect 471756 266376 473728 266404
rect 471756 266364 471762 266376
rect 473722 266364 473728 266376
rect 473780 266364 473786 266416
rect 470234 265087 470854 265093
rect 470234 264779 470262 265087
rect 470826 264779 470854 265087
rect 470234 264773 470854 264779
rect 473648 264092 473676 264264
rect 473722 264092 473728 264104
rect 473648 264064 473728 264092
rect 473722 264052 473728 264064
rect 473780 264052 473786 264104
rect 468994 264001 469614 264007
rect 468994 263693 469022 264001
rect 469586 263693 469614 264001
rect 468994 263687 469614 263693
rect 477089 263075 477147 263081
rect 477089 263041 477101 263075
rect 477135 263072 477147 263075
rect 477218 263072 477224 263084
rect 477135 263044 477224 263072
rect 477135 263041 477147 263044
rect 477089 263035 477147 263041
rect 477218 263032 477224 263044
rect 477276 263032 477282 263084
rect 470234 262914 470854 262920
rect 470234 262606 470262 262914
rect 470826 262606 470854 262914
rect 470234 262600 470854 262606
rect 536742 212780 536748 212832
rect 536800 212820 536806 212832
rect 544105 212823 544163 212829
rect 544105 212820 544117 212823
rect 536800 212792 544117 212820
rect 536800 212780 536806 212792
rect 544105 212789 544117 212792
rect 544151 212789 544163 212823
rect 544105 212783 544163 212789
rect 473722 206932 473728 206984
rect 473780 206972 473786 206984
rect 580166 206972 580172 206984
rect 473780 206944 580172 206972
rect 473780 206932 473786 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
<< via1 >>
rect 470262 451177 470826 451485
rect 471336 450644 471388 450696
rect 469022 450091 469586 450399
rect 488264 449964 488316 450016
rect 489000 449828 489052 449880
rect 475384 449433 475436 449485
rect 478696 449433 478748 449485
rect 482008 449433 482060 449485
rect 485320 449433 485372 449485
rect 488816 449433 488868 449485
rect 470262 449006 470826 449314
rect 544568 445136 544620 445188
rect 547880 445136 547932 445188
rect 493508 434732 493560 434784
rect 535460 434732 535512 434784
rect 470262 432778 470826 433086
rect 481548 432692 481600 432744
rect 483112 432692 483164 432744
rect 471612 432238 471664 432290
rect 471796 432216 471848 432268
rect 483112 432080 483164 432132
rect 469022 431691 469586 431999
rect 477960 431128 478012 431180
rect 489644 431400 489696 431452
rect 470262 430606 470826 430914
rect 470262 411778 470826 412086
rect 471612 411544 471664 411596
rect 471244 411272 471296 411324
rect 469022 410692 469586 411000
rect 488540 410456 488592 410508
rect 489092 410456 489144 410508
rect 475292 410033 475344 410085
rect 478696 410048 478748 410100
rect 481824 410033 481876 410085
rect 485228 410048 485280 410100
rect 488540 410033 488592 410085
rect 470262 409606 470826 409914
rect 544660 409164 544712 409216
rect 547880 409164 547932 409216
rect 488540 407736 488592 407788
rect 489460 407736 489512 407788
rect 470262 390779 470826 391087
rect 471704 390464 471756 390516
rect 471520 390238 471572 390290
rect 478052 390238 478104 390290
rect 471704 390056 471756 390108
rect 469022 389696 469586 390004
rect 490840 389512 490892 389564
rect 475752 389033 475804 389085
rect 479616 389036 479668 389088
rect 483204 389033 483256 389085
rect 486884 389033 486936 389085
rect 470262 388606 470826 388914
rect 545028 373192 545080 373244
rect 548524 373192 548576 373244
rect 470262 369779 470826 370087
rect 473728 369452 473780 369504
rect 471704 369316 471756 369368
rect 478880 369238 478932 369290
rect 481272 369238 481324 369290
rect 488908 369248 488960 369300
rect 489828 369248 489880 369300
rect 473912 369112 473964 369164
rect 481272 369112 481324 369164
rect 481824 369112 481876 369164
rect 469022 368693 469586 369001
rect 485320 368568 485372 368620
rect 489644 368500 489696 368552
rect 489460 368032 489512 368084
rect 477224 367956 477276 368008
rect 470262 367606 470826 367914
rect 490564 363604 490616 363656
rect 536196 363604 536248 363656
rect 470262 348778 470826 349086
rect 475660 348508 475712 348560
rect 471612 348440 471664 348492
rect 471796 348100 471848 348152
rect 489092 348236 489144 348288
rect 469022 347691 469586 347999
rect 488540 347284 488592 347336
rect 475568 347012 475620 347064
rect 478604 347012 478656 347064
rect 482192 347012 482244 347064
rect 485412 347035 485464 347087
rect 489000 347012 489052 347064
rect 470262 346606 470826 346914
rect 485412 328176 485464 328228
rect 488816 328176 488868 328228
rect 489736 328176 489788 328228
rect 470262 327778 470826 328086
rect 471244 327292 471296 327344
rect 469022 326691 469586 326999
rect 489552 326408 489604 326460
rect 489368 326340 489420 326392
rect 536288 326408 536340 326460
rect 479064 326000 479116 326052
rect 492036 326000 492088 326052
rect 470262 325606 470826 325914
rect 470262 306778 470826 307086
rect 471704 306484 471756 306536
rect 471244 306280 471296 306332
rect 469022 305693 469586 306001
rect 478604 305507 478656 305516
rect 478604 305473 478614 305507
rect 478614 305473 478656 305507
rect 478604 305464 478656 305473
rect 485136 305507 485188 305516
rect 485136 305473 485144 305507
rect 485144 305473 485188 305507
rect 485136 305464 485188 305473
rect 489276 305396 489328 305448
rect 475292 305033 475344 305085
rect 481824 305033 481876 305085
rect 490656 304988 490708 305040
rect 470262 304606 470826 304914
rect 475292 303560 475344 303612
rect 478604 303560 478656 303612
rect 485136 303560 485188 303612
rect 536380 303560 536432 303612
rect 493508 303492 493560 303544
rect 490564 303424 490616 303476
rect 481824 303356 481876 303408
rect 489184 303356 489236 303408
rect 490656 292476 490708 292528
rect 535460 292476 535512 292528
rect 470262 285779 470826 286087
rect 471428 285239 471480 285291
rect 478052 285238 478104 285290
rect 489276 285238 489328 285290
rect 491392 285132 491444 285184
rect 471704 285064 471756 285116
rect 469022 284694 469586 285002
rect 475752 284033 475804 284085
rect 479616 284044 479668 284096
rect 483204 284033 483256 284085
rect 486884 284033 486936 284085
rect 470262 283606 470826 283914
rect 471704 266364 471756 266416
rect 473728 266364 473780 266416
rect 470262 264779 470826 265087
rect 473728 264052 473780 264104
rect 469022 263693 469586 264001
rect 477224 263032 477276 263084
rect 470262 262606 470826 262914
rect 536748 212780 536800 212832
rect 473728 206932 473780 206984
rect 580172 206932 580224 206984
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 470138 451616 470194 451625
rect 470138 451551 470194 451560
rect 488906 451616 488962 451625
rect 488906 451551 488962 451560
rect 469022 450399 469586 450405
rect 469022 450085 469586 450091
rect 469022 431999 469586 432005
rect 469022 431685 469586 431691
rect 470152 429865 470180 451551
rect 470262 451485 470826 451491
rect 470262 451171 470826 451177
rect 481160 450800 481216 450809
rect 471256 450758 471376 450786
rect 470262 449314 470826 449320
rect 470262 449000 470826 449006
rect 470262 433086 470826 433092
rect 470262 432772 470826 432778
rect 471256 432290 471284 450758
rect 471348 450702 471376 450758
rect 481160 450735 481216 450744
rect 471336 450696 471388 450702
rect 471336 450638 471388 450644
rect 472772 450622 473308 450650
rect 473280 450514 473308 450622
rect 476052 450608 476061 450664
rect 476117 450608 476126 450664
rect 473280 450486 473400 450514
rect 473372 434625 473400 450486
rect 488264 450016 488316 450022
rect 488316 449964 488580 449970
rect 488264 449958 488580 449964
rect 488276 449942 488580 449958
rect 475384 449485 475436 449491
rect 475384 449427 475436 449433
rect 478696 449485 478748 449491
rect 478696 449427 478748 449433
rect 482008 449485 482060 449491
rect 482008 449427 482060 449433
rect 485320 449485 485372 449491
rect 485320 449427 485372 449433
rect 475396 444961 475424 449427
rect 478708 447953 478736 449427
rect 478694 447944 478750 447953
rect 478694 447879 478750 447888
rect 482020 447817 482048 449427
rect 482006 447808 482062 447817
rect 482006 447743 482062 447752
rect 475382 444952 475438 444961
rect 475382 444887 475438 444896
rect 483202 435160 483258 435169
rect 483124 435118 483202 435146
rect 481546 435024 481602 435033
rect 481546 434959 481602 434968
rect 471886 434616 471942 434625
rect 471716 434574 471886 434602
rect 471612 432290 471664 432296
rect 471256 432262 471612 432290
rect 470262 430914 470826 430920
rect 470262 430600 470826 430606
rect 470138 429856 470194 429865
rect 470138 429791 470194 429800
rect 470262 412086 470826 412092
rect 470262 411772 470826 411778
rect 471256 411330 471284 432262
rect 471612 432232 471664 432238
rect 471716 432154 471744 434574
rect 471886 434551 471942 434560
rect 473358 434616 473414 434625
rect 473358 434551 473414 434560
rect 481560 432750 481588 434959
rect 483124 432750 483152 435118
rect 483202 435095 483258 435104
rect 485332 433945 485360 449427
rect 488552 445890 488580 449942
rect 488816 449485 488868 449491
rect 488814 449440 488816 449449
rect 488868 449440 488870 449449
rect 488814 449375 488870 449384
rect 488920 446434 488948 451551
rect 489000 449880 489052 449886
rect 489000 449822 489052 449828
rect 488460 445862 488580 445890
rect 488828 446406 488948 446434
rect 488460 434625 488488 445862
rect 488828 441614 488856 446406
rect 488828 441586 488948 441614
rect 488920 435033 488948 441586
rect 489012 435169 489040 449822
rect 497462 449440 497518 449449
rect 497462 449375 497518 449384
rect 490562 447944 490618 447953
rect 490562 447879 490618 447888
rect 488998 435160 489054 435169
rect 488998 435095 489054 435104
rect 488906 435024 488962 435033
rect 488962 434982 489500 435010
rect 488906 434959 488962 434968
rect 488446 434616 488502 434625
rect 488446 434551 488502 434560
rect 485318 433936 485374 433945
rect 485318 433871 485374 433880
rect 481548 432744 481600 432750
rect 481548 432686 481600 432692
rect 483112 432744 483164 432750
rect 483112 432686 483164 432692
rect 471796 432268 471848 432274
rect 471796 432210 471848 432216
rect 471808 432154 471836 432210
rect 471716 432126 471836 432154
rect 483112 432132 483164 432138
rect 471716 422294 471744 432126
rect 483112 432074 483164 432080
rect 483124 431954 483152 432074
rect 483124 431926 483244 431954
rect 475488 429185 475516 431596
rect 478998 431582 479288 431610
rect 477960 431180 478012 431186
rect 477960 431122 478012 431128
rect 477972 429865 478000 431122
rect 477958 429856 478014 429865
rect 477958 429791 478014 429800
rect 475474 429176 475530 429185
rect 475474 429111 475530 429120
rect 471624 422266 471744 422294
rect 471518 412312 471574 412321
rect 471518 412247 471574 412256
rect 471244 411324 471296 411330
rect 471244 411266 471296 411272
rect 469022 411000 469586 411006
rect 469022 410686 469586 410692
rect 470262 409914 470826 409920
rect 470262 409600 470826 409606
rect 470138 392592 470194 392601
rect 470138 392527 470194 392536
rect 469022 390004 469586 390010
rect 469022 389690 469586 389696
rect 470152 370297 470180 392527
rect 470262 391087 470826 391093
rect 470262 390773 470826 390779
rect 471256 390402 471284 411266
rect 471532 392601 471560 412247
rect 471624 411602 471652 422266
rect 477972 412634 478000 429791
rect 479260 428505 479288 431582
rect 479246 428496 479302 428505
rect 479246 428431 479302 428440
rect 482388 413409 482416 431596
rect 483216 430681 483244 431926
rect 489090 431624 489146 431633
rect 489146 431582 489302 431610
rect 489090 431559 489146 431568
rect 483202 430672 483258 430681
rect 483202 430607 483258 430616
rect 484306 430672 484362 430681
rect 484306 430607 484362 430616
rect 482374 413400 482430 413409
rect 482374 413335 482430 413344
rect 481086 412720 481142 412729
rect 481086 412655 481142 412664
rect 477788 412606 478000 412634
rect 477788 412321 477816 412606
rect 477774 412312 477830 412321
rect 477774 412247 477830 412256
rect 477788 411913 477816 412247
rect 481100 411913 481128 412655
rect 484320 412321 484348 430607
rect 485870 430400 485926 430409
rect 485870 430335 485926 430344
rect 485884 413273 485912 430335
rect 489274 428496 489330 428505
rect 489274 428431 489330 428440
rect 488538 413944 488594 413953
rect 488538 413879 488594 413888
rect 485870 413264 485926 413273
rect 485870 413199 485926 413208
rect 484306 412312 484362 412321
rect 484306 412247 484362 412256
rect 484320 411913 484348 412247
rect 477774 411904 477830 411913
rect 477774 411839 477830 411848
rect 481086 411904 481142 411913
rect 481086 411839 481142 411848
rect 484306 411904 484362 411913
rect 484306 411839 484362 411848
rect 477682 411632 477738 411641
rect 471612 411596 471664 411602
rect 471612 411538 471664 411544
rect 477604 411590 477682 411618
rect 471518 392592 471574 392601
rect 471518 392527 471574 392536
rect 471532 392057 471560 392527
rect 471518 392048 471574 392057
rect 471518 391983 471574 391992
rect 471256 390374 471560 390402
rect 471532 390296 471560 390374
rect 471520 390290 471572 390296
rect 471520 390232 471572 390238
rect 471624 390266 471652 411538
rect 477604 410938 477632 411590
rect 481086 411632 481142 411641
rect 477682 411567 477738 411576
rect 481008 411590 481086 411618
rect 481008 411482 481036 411590
rect 481086 411567 481142 411576
rect 484306 411632 484362 411641
rect 484306 411567 484362 411576
rect 484320 411482 484348 411567
rect 481008 411454 481047 411482
rect 481019 411196 481047 411454
rect 484284 411454 484348 411482
rect 484284 411196 484312 411454
rect 477604 410910 477768 410938
rect 488552 410514 488580 413879
rect 488722 412312 488778 412321
rect 488722 412247 488778 412256
rect 488540 410508 488592 410514
rect 488540 410450 488592 410456
rect 488538 410136 488594 410145
rect 478696 410100 478748 410106
rect 475292 410085 475344 410091
rect 485228 410100 485280 410106
rect 478696 410042 478748 410048
rect 481824 410085 481876 410091
rect 475292 410027 475344 410033
rect 475304 408513 475332 410027
rect 475290 408504 475346 408513
rect 475290 408439 475346 408448
rect 478708 406201 478736 410042
rect 488538 410071 488540 410080
rect 485228 410042 485280 410048
rect 481824 410027 481876 410033
rect 478694 406192 478750 406201
rect 478694 406127 478750 406136
rect 481836 392601 481864 410027
rect 485240 393961 485268 410042
rect 488592 410071 488594 410080
rect 488540 410027 488592 410033
rect 488540 407788 488592 407794
rect 488540 407730 488592 407736
rect 485226 393952 485282 393961
rect 485226 393887 485282 393896
rect 481822 392592 481878 392601
rect 481822 392527 481878 392536
rect 488552 392193 488580 407730
rect 488736 393314 488764 412247
rect 489092 410508 489144 410514
rect 489092 410450 489144 410456
rect 489104 402974 489132 410450
rect 489288 407561 489316 428431
rect 489472 412729 489500 434982
rect 489642 434616 489698 434625
rect 489642 434551 489698 434560
rect 489656 431458 489684 434551
rect 489644 431452 489696 431458
rect 489644 431394 489696 431400
rect 489656 413953 489684 431394
rect 489642 413944 489698 413953
rect 489642 413879 489698 413888
rect 489458 412720 489514 412729
rect 489458 412655 489514 412664
rect 489472 407794 489500 412655
rect 490576 408921 490604 447879
rect 490746 443592 490802 443601
rect 490746 443527 490802 443536
rect 490654 442232 490710 442241
rect 490654 442167 490710 442176
rect 490562 408912 490618 408921
rect 490562 408847 490618 408856
rect 490668 408513 490696 442167
rect 490760 429185 490788 443527
rect 492126 440872 492182 440881
rect 492126 440807 492182 440816
rect 492034 438152 492090 438161
rect 492034 438087 492090 438096
rect 491942 431624 491998 431633
rect 491942 431559 491998 431568
rect 490746 429176 490802 429185
rect 490746 429111 490802 429120
rect 490654 408504 490710 408513
rect 490654 408439 490710 408448
rect 489460 407788 489512 407794
rect 489460 407730 489512 407736
rect 489274 407552 489330 407561
rect 489274 407487 489330 407496
rect 489104 402946 489224 402974
rect 488644 393286 488764 393314
rect 482558 392184 482614 392193
rect 482558 392119 482614 392128
rect 488538 392184 488594 392193
rect 488538 392119 488594 392128
rect 477866 392048 477922 392057
rect 477866 391983 477922 391992
rect 477880 390969 477908 391983
rect 482572 390969 482600 392119
rect 488644 392057 488672 393286
rect 488630 392048 488686 392057
rect 488630 391983 488686 391992
rect 489196 390969 489224 402946
rect 490746 392184 490802 392193
rect 490746 392119 490802 392128
rect 477866 390960 477922 390969
rect 477866 390895 477922 390904
rect 482558 390960 482614 390969
rect 482558 390895 482614 390904
rect 489182 390960 489238 390969
rect 489182 390895 489238 390904
rect 478050 390688 478106 390697
rect 478050 390623 478106 390632
rect 482374 390688 482430 390697
rect 482374 390623 482430 390632
rect 489458 390688 489514 390697
rect 489458 390623 489514 390632
rect 471704 390516 471756 390522
rect 471704 390458 471756 390464
rect 471716 390266 471744 390458
rect 478064 390296 478092 390623
rect 471624 390238 471744 390266
rect 478052 390290 478104 390296
rect 482388 390252 482416 390623
rect 489472 390266 489500 390623
rect 489472 390252 489798 390266
rect 489472 390238 489812 390252
rect 470262 388914 470826 388920
rect 470262 388600 470826 388606
rect 471624 371385 471652 390238
rect 478052 390232 478104 390238
rect 471704 390108 471756 390114
rect 471704 390050 471756 390056
rect 471610 371376 471666 371385
rect 471610 371311 471666 371320
rect 470138 370288 470194 370297
rect 470138 370223 470194 370232
rect 470262 370087 470826 370093
rect 470262 369773 470826 369779
rect 471716 369374 471744 390050
rect 489784 389178 489812 390238
rect 489784 389150 489960 389178
rect 475752 389085 475804 389091
rect 475752 389027 475804 389033
rect 479616 389088 479668 389094
rect 479616 389030 479668 389036
rect 483204 389085 483256 389091
rect 475764 387705 475792 389027
rect 475750 387696 475806 387705
rect 475750 387631 475806 387640
rect 479628 387569 479656 389030
rect 483204 389027 483256 389033
rect 486884 389085 486936 389091
rect 486884 389027 486936 389033
rect 479614 387560 479670 387569
rect 479614 387495 479670 387504
rect 483216 386481 483244 389027
rect 483202 386472 483258 386481
rect 483202 386407 483258 386416
rect 485686 382392 485742 382401
rect 485686 382327 485742 382336
rect 482374 371920 482430 371929
rect 482374 371855 482430 371864
rect 473726 371376 473782 371385
rect 473726 371311 473782 371320
rect 473266 370288 473322 370297
rect 473266 370223 473322 370232
rect 471704 369368 471756 369374
rect 471704 369310 471756 369316
rect 469022 369001 469586 369007
rect 469022 368687 469586 368693
rect 470262 367914 470826 367920
rect 470262 367600 470826 367606
rect 471716 354674 471744 369310
rect 473280 359553 473308 370223
rect 473740 369510 473768 371311
rect 482388 369889 482416 371855
rect 485700 369889 485728 382327
rect 486896 372065 486924 389027
rect 489550 386472 489606 386481
rect 489550 386407 489606 386416
rect 486882 372056 486938 372065
rect 486882 371991 486938 372000
rect 482374 369880 482430 369889
rect 482374 369815 482430 369824
rect 485686 369880 485742 369889
rect 485686 369815 485742 369824
rect 478878 369608 478934 369617
rect 478878 369543 478934 369552
rect 481822 369608 481878 369617
rect 481822 369543 481878 369552
rect 485318 369608 485374 369617
rect 485318 369543 485374 369552
rect 473728 369504 473780 369510
rect 473728 369446 473780 369452
rect 473740 368914 473768 369446
rect 478892 369296 478920 369543
rect 478880 369290 478932 369296
rect 478880 369232 478932 369238
rect 481272 369290 481324 369296
rect 481272 369232 481324 369238
rect 481284 369170 481312 369232
rect 481836 369170 481864 369543
rect 473912 369164 473964 369170
rect 473912 369106 473964 369112
rect 481272 369164 481324 369170
rect 481272 369106 481324 369112
rect 481824 369164 481876 369170
rect 481824 369106 481876 369112
rect 473372 368886 473768 368914
rect 473266 359544 473322 359553
rect 473266 359479 473322 359488
rect 471624 354646 471744 354674
rect 470262 349086 470826 349092
rect 470262 348772 470826 348778
rect 471624 348498 471652 354646
rect 473372 349217 473400 368886
rect 473924 354674 473952 369106
rect 477224 368008 477276 368014
rect 477224 367950 477276 367956
rect 477236 367033 477264 367950
rect 477222 367024 477278 367033
rect 477222 366959 477278 366968
rect 480180 366897 480208 368628
rect 480166 366888 480222 366897
rect 480166 366823 480222 366832
rect 483216 366761 483244 368628
rect 485332 368626 485360 369543
rect 488908 369300 488960 369306
rect 488908 369242 488960 369248
rect 485320 368620 485372 368626
rect 486266 368614 486464 368642
rect 485320 368562 485372 368568
rect 483202 366752 483258 366761
rect 483202 366687 483258 366696
rect 476118 359544 476174 359553
rect 476118 359479 476174 359488
rect 473740 354646 473952 354674
rect 473740 350577 473768 354646
rect 473726 350568 473782 350577
rect 473726 350503 473782 350512
rect 471702 349208 471758 349217
rect 471702 349143 471758 349152
rect 473358 349208 473414 349217
rect 473358 349143 473414 349152
rect 471612 348492 471664 348498
rect 471612 348434 471664 348440
rect 469022 347999 469586 348005
rect 469022 347685 469586 347691
rect 470262 346914 470826 346920
rect 470262 346600 470826 346606
rect 471624 345014 471652 348434
rect 471256 344986 471652 345014
rect 470262 328086 470826 328092
rect 470262 327772 470826 327778
rect 471256 327350 471284 344986
rect 471716 342281 471744 349143
rect 476132 348809 476160 359479
rect 481270 350568 481326 350577
rect 481270 350503 481326 350512
rect 481284 348809 481312 350503
rect 486436 349761 486464 368614
rect 488920 364334 488948 369242
rect 489564 368801 489592 386407
rect 489932 371362 489960 389150
rect 490654 372056 490710 372065
rect 490654 371991 490710 372000
rect 489840 371334 489960 371362
rect 489840 369306 489868 371334
rect 489828 369300 489880 369306
rect 489828 369242 489880 369248
rect 489550 368792 489606 368801
rect 489550 368727 489606 368736
rect 489644 368552 489696 368558
rect 489644 368494 489696 368500
rect 489458 368112 489514 368121
rect 489458 368047 489460 368056
rect 489512 368047 489514 368056
rect 489460 368026 489512 368032
rect 489366 367296 489422 367305
rect 489366 367231 489422 367240
rect 488920 364306 489132 364334
rect 488814 350704 488870 350713
rect 488814 350639 488870 350648
rect 486422 349752 486478 349761
rect 486422 349687 486478 349696
rect 476118 348800 476174 348809
rect 476118 348735 476174 348744
rect 481270 348800 481326 348809
rect 481270 348735 481326 348744
rect 475660 348560 475712 348566
rect 475658 348528 475660 348537
rect 475712 348528 475714 348537
rect 475658 348463 475714 348472
rect 474186 348392 474242 348401
rect 481232 348392 481288 348401
rect 474242 348350 474626 348378
rect 474186 348327 474242 348336
rect 481232 348327 481288 348336
rect 471796 348152 471848 348158
rect 471796 348094 471848 348100
rect 471702 342272 471758 342281
rect 471702 342207 471758 342216
rect 471808 335354 471836 348094
rect 488540 347336 488592 347342
rect 488828 347290 488856 350639
rect 488906 350568 488962 350577
rect 488906 350503 488962 350512
rect 488592 347284 488856 347290
rect 488540 347278 488856 347284
rect 488552 347262 488856 347278
rect 485412 347087 485464 347093
rect 475568 347064 475620 347070
rect 475568 347006 475620 347012
rect 478604 347064 478656 347070
rect 478604 347006 478656 347012
rect 482192 347064 482244 347070
rect 485412 347029 485464 347035
rect 482192 347006 482244 347012
rect 475580 346361 475608 347006
rect 475566 346352 475622 346361
rect 475566 346287 475622 346296
rect 478616 345001 478644 347006
rect 478602 344992 478658 345001
rect 478602 344927 478658 344936
rect 482204 344865 482232 347006
rect 482190 344856 482246 344865
rect 482190 344791 482246 344800
rect 474646 342272 474702 342281
rect 474646 342207 474702 342216
rect 471532 335326 471836 335354
rect 471244 327344 471296 327350
rect 471244 327286 471296 327292
rect 469022 326999 469586 327005
rect 469022 326685 469586 326691
rect 470262 325914 470826 325920
rect 470262 325600 470826 325606
rect 470262 307086 470826 307092
rect 470262 306772 470826 306778
rect 471256 306338 471284 327286
rect 471532 326913 471560 335326
rect 471610 329896 471666 329905
rect 471610 329831 471666 329840
rect 471518 326904 471574 326913
rect 471518 326839 471574 326848
rect 471532 307873 471560 326839
rect 471624 308417 471652 329831
rect 474660 327865 474688 342207
rect 485424 330041 485452 347029
rect 488828 335354 488856 347262
rect 488736 335326 488856 335354
rect 488736 331214 488764 335326
rect 488736 331186 488856 331214
rect 485410 330032 485466 330041
rect 485410 329967 485466 329976
rect 481546 329896 481602 329905
rect 481546 329831 481602 329840
rect 481560 327865 481588 329831
rect 488828 328234 488856 331186
rect 488920 329905 488948 350503
rect 489104 348294 489132 364306
rect 489092 348288 489144 348294
rect 489092 348230 489144 348236
rect 489000 347064 489052 347070
rect 488998 347032 489000 347041
rect 489052 347032 489054 347041
rect 488998 346967 489054 346976
rect 489104 345014 489132 348230
rect 489104 344986 489224 345014
rect 489196 330970 489224 344986
rect 489380 331214 489408 367231
rect 489656 350713 489684 368494
rect 490564 363656 490616 363662
rect 490564 363598 490616 363604
rect 489642 350704 489698 350713
rect 489642 350639 489698 350648
rect 489380 331186 489684 331214
rect 489196 330942 489592 330970
rect 488906 329896 488962 329905
rect 488906 329831 488962 329840
rect 485412 328228 485464 328234
rect 485412 328170 485464 328176
rect 488816 328228 488868 328234
rect 488816 328170 488868 328176
rect 485424 327865 485452 328170
rect 474646 327856 474702 327865
rect 474646 327791 474702 327800
rect 481546 327856 481602 327865
rect 481546 327791 481602 327800
rect 485410 327856 485466 327865
rect 485410 327791 485466 327800
rect 471702 327720 471758 327729
rect 471702 327655 471758 327664
rect 471610 308408 471666 308417
rect 471610 308343 471666 308352
rect 471518 307864 471574 307873
rect 471518 307799 471574 307808
rect 471244 306332 471296 306338
rect 471244 306274 471296 306280
rect 469022 306001 469586 306007
rect 469022 305687 469586 305693
rect 470262 304914 470826 304920
rect 470262 304600 470826 304606
rect 471256 302234 471284 306274
rect 471256 302206 471376 302234
rect 471348 287054 471376 302206
rect 471532 287337 471560 307799
rect 471716 306542 471744 327655
rect 481542 327448 481598 327457
rect 474644 327392 474653 327448
rect 474709 327392 474718 327448
rect 484977 327392 484986 327448
rect 485042 327392 485051 327448
rect 481542 327383 481598 327392
rect 476224 326913 476252 327298
rect 476210 326904 476266 326913
rect 476210 326839 476266 326848
rect 475488 325417 475516 326604
rect 479064 326052 479116 326058
rect 479064 325994 479116 326000
rect 475474 325408 475530 325417
rect 475474 325343 475530 325352
rect 479076 324193 479104 325994
rect 479062 324184 479118 324193
rect 479062 324119 479118 324128
rect 482388 324057 482416 326604
rect 489564 326466 489592 330942
rect 489552 326460 489604 326466
rect 489552 326402 489604 326408
rect 489368 326392 489420 326398
rect 489368 326334 489420 326340
rect 482374 324048 482430 324057
rect 482374 323983 482430 323992
rect 489380 316034 489408 326334
rect 489564 316034 489592 326402
rect 489656 324193 489684 331186
rect 489918 328672 489974 328681
rect 489918 328607 489974 328616
rect 489736 328228 489788 328234
rect 489736 328170 489788 328176
rect 489642 324184 489698 324193
rect 489642 324119 489698 324128
rect 489748 318794 489776 328170
rect 489932 326913 489960 328607
rect 489918 326904 489974 326913
rect 489918 326839 489974 326848
rect 489196 316006 489408 316034
rect 489472 316006 489592 316034
rect 489656 318766 489776 318794
rect 488630 313304 488686 313313
rect 488630 313239 488686 313248
rect 480902 308408 480958 308417
rect 480902 308343 480958 308352
rect 488538 308408 488594 308417
rect 488538 308343 488594 308352
rect 477498 307864 477554 307873
rect 477498 307799 477554 307808
rect 477512 306921 477540 307799
rect 480916 306921 480944 308343
rect 477498 306912 477554 306921
rect 477498 306847 477554 306856
rect 480902 306912 480958 306921
rect 480902 306847 480958 306856
rect 477590 306640 477646 306649
rect 477590 306575 477646 306584
rect 480902 306640 480958 306649
rect 480902 306575 480958 306584
rect 484306 306640 484362 306649
rect 484306 306575 484362 306584
rect 471704 306536 471756 306542
rect 471704 306478 471756 306484
rect 471716 296714 471744 306478
rect 477604 306082 477632 306575
rect 480916 306082 480944 306575
rect 484320 306374 484348 306575
rect 484283 306346 484348 306374
rect 484283 306204 484311 306346
rect 477604 306054 477767 306082
rect 480916 306054 481032 306082
rect 478604 305516 478656 305522
rect 478604 305458 478656 305464
rect 485136 305516 485188 305522
rect 485136 305458 485188 305464
rect 475292 305085 475344 305091
rect 475292 305027 475344 305033
rect 475304 303618 475332 305027
rect 478616 303618 478644 305458
rect 481824 305085 481876 305091
rect 481824 305027 481876 305033
rect 475292 303612 475344 303618
rect 475292 303554 475344 303560
rect 478604 303612 478656 303618
rect 478604 303554 478656 303560
rect 481836 303414 481864 305027
rect 485148 303618 485176 305458
rect 485136 303612 485188 303618
rect 485136 303554 485188 303560
rect 481824 303408 481876 303414
rect 481824 303350 481876 303356
rect 471624 296686 471744 296714
rect 471518 287328 471574 287337
rect 471518 287263 471574 287272
rect 471348 287026 471468 287054
rect 470262 286087 470826 286093
rect 470262 285773 470826 285779
rect 471440 285297 471468 287026
rect 471428 285291 471480 285297
rect 471428 285233 471480 285239
rect 469022 285002 469586 285008
rect 469022 284688 469586 284694
rect 470262 283914 470826 283920
rect 470262 283600 470826 283606
rect 471532 266801 471560 287263
rect 471624 287201 471652 296686
rect 488552 287473 488580 308343
rect 488644 306785 488672 313239
rect 488630 306776 488686 306785
rect 488630 306711 488686 306720
rect 482558 287464 482614 287473
rect 482558 287399 482614 287408
rect 488538 287464 488594 287473
rect 488538 287399 488594 287408
rect 477866 287328 477922 287337
rect 477866 287263 477922 287272
rect 471610 287192 471666 287201
rect 471610 287127 471666 287136
rect 474738 287192 474794 287201
rect 474738 287127 474794 287136
rect 471518 266792 471574 266801
rect 471518 266727 471574 266736
rect 471624 266393 471652 287127
rect 474752 285977 474780 287127
rect 477880 285977 477908 287263
rect 482572 285977 482600 287399
rect 488644 287337 488672 306711
rect 489196 303414 489224 316006
rect 489472 306374 489500 316006
rect 489656 313313 489684 318766
rect 489642 313304 489698 313313
rect 489642 313239 489698 313248
rect 489288 306346 489500 306374
rect 489288 305454 489316 306346
rect 489276 305448 489328 305454
rect 489276 305390 489328 305396
rect 489184 303408 489236 303414
rect 489184 303350 489236 303356
rect 488630 287328 488686 287337
rect 488630 287263 488686 287272
rect 489288 287201 489316 305390
rect 490576 303482 490604 363598
rect 490668 332761 490696 371991
rect 490760 371929 490788 392119
rect 490838 392048 490894 392057
rect 490838 391983 490894 391992
rect 490852 389570 490880 391983
rect 490840 389564 490892 389570
rect 490840 389506 490892 389512
rect 490852 382401 490880 389506
rect 490838 382392 490894 382401
rect 490838 382327 490894 382336
rect 490746 371920 490802 371929
rect 490746 371855 490802 371864
rect 490746 364984 490802 364993
rect 490746 364919 490802 364928
rect 490760 344865 490788 364919
rect 490746 344856 490802 344865
rect 490746 344791 490802 344800
rect 490654 332752 490710 332761
rect 490654 332687 490710 332696
rect 490746 325000 490802 325009
rect 490746 324935 490802 324944
rect 490656 305040 490708 305046
rect 490656 304982 490708 304988
rect 490564 303476 490616 303482
rect 490564 303418 490616 303424
rect 490668 292534 490696 304982
rect 490656 292528 490708 292534
rect 490656 292470 490708 292476
rect 489274 287192 489330 287201
rect 489274 287127 489330 287136
rect 489288 285977 489316 287127
rect 474738 285968 474794 285977
rect 474738 285903 474794 285912
rect 477866 285968 477922 285977
rect 477866 285903 477922 285912
rect 482558 285968 482614 285977
rect 482558 285903 482614 285912
rect 489274 285968 489330 285977
rect 489274 285903 489330 285912
rect 474738 285696 474794 285705
rect 474738 285631 474794 285640
rect 478050 285696 478106 285705
rect 478050 285631 478106 285640
rect 482374 285696 482430 285705
rect 482374 285631 482430 285640
rect 489274 285696 489330 285705
rect 489274 285631 489330 285640
rect 474752 285274 474780 285631
rect 478064 285296 478092 285631
rect 478052 285290 478104 285296
rect 474752 285246 474949 285274
rect 482388 285260 482416 285631
rect 489288 285296 489316 285631
rect 489276 285290 489328 285296
rect 478052 285232 478104 285238
rect 489276 285232 489328 285238
rect 471704 285116 471756 285122
rect 471704 285058 471756 285064
rect 471716 266422 471744 285058
rect 479616 284096 479668 284102
rect 475752 284085 475804 284091
rect 479616 284038 479668 284044
rect 483204 284085 483256 284091
rect 475752 284027 475804 284033
rect 475764 282713 475792 284027
rect 475750 282704 475806 282713
rect 475750 282639 475806 282648
rect 479628 282441 479656 284038
rect 483204 284027 483256 284033
rect 486884 284085 486936 284091
rect 486884 284027 486936 284033
rect 483216 282577 483244 284027
rect 486896 282849 486924 284027
rect 486882 282840 486938 282849
rect 486882 282775 486938 282784
rect 483202 282568 483258 282577
rect 483202 282503 483258 282512
rect 479614 282432 479670 282441
rect 479614 282367 479670 282376
rect 476118 266928 476174 266937
rect 476118 266863 476174 266872
rect 490562 266928 490618 266937
rect 490562 266863 490618 266872
rect 471704 266416 471756 266422
rect 471610 266384 471666 266393
rect 471704 266358 471756 266364
rect 473728 266416 473780 266422
rect 476132 266393 476160 266863
rect 479062 266792 479118 266801
rect 479062 266727 479118 266736
rect 473728 266358 473780 266364
rect 476118 266384 476174 266393
rect 471610 266319 471666 266328
rect 470262 265087 470826 265093
rect 470262 264773 470826 264779
rect 473740 264110 473768 266358
rect 476118 266319 476174 266328
rect 476132 264897 476160 266319
rect 479076 264897 479104 266727
rect 482558 266656 482614 266665
rect 482558 266591 482614 266600
rect 489826 266656 489882 266665
rect 489826 266591 489882 266600
rect 482572 264897 482600 266591
rect 488446 266520 488502 266529
rect 488446 266455 488502 266464
rect 485318 266384 485374 266393
rect 485318 266319 485374 266328
rect 485332 264897 485360 266319
rect 488460 264897 488488 266455
rect 476118 264888 476174 264897
rect 476118 264823 476174 264832
rect 479062 264888 479118 264897
rect 479062 264823 479118 264832
rect 482558 264888 482614 264897
rect 482558 264823 482614 264832
rect 485318 264888 485374 264897
rect 485318 264823 485374 264832
rect 488446 264888 488502 264897
rect 488446 264823 488502 264832
rect 476118 264616 476174 264625
rect 476118 264551 476174 264560
rect 479062 264616 479118 264625
rect 479062 264551 479118 264560
rect 482374 264616 482430 264625
rect 482374 264551 482430 264560
rect 485410 264616 485466 264625
rect 485410 264551 485466 264560
rect 488446 264616 488502 264625
rect 488446 264551 488502 264560
rect 476132 264194 476160 264551
rect 479076 264194 479104 264551
rect 482388 264466 482416 264551
rect 482379 264438 482416 264466
rect 476132 264166 476289 264194
rect 479076 264166 479341 264194
rect 482379 264180 482407 264438
rect 485424 264166 485452 264551
rect 488460 264194 488488 264551
rect 488460 264166 488497 264194
rect 473728 264104 473780 264110
rect 473728 264046 473780 264052
rect 469022 264001 469586 264007
rect 469022 263687 469586 263693
rect 470262 262914 470826 262920
rect 470262 262600 470826 262606
rect 473740 206990 473768 264046
rect 477224 263084 477276 263090
rect 477224 263026 477276 263032
rect 477236 261769 477264 263026
rect 480180 261905 480208 263636
rect 483216 262041 483244 263636
rect 486252 262177 486280 263636
rect 489302 263622 489500 263650
rect 489472 263537 489500 263622
rect 489458 263528 489514 263537
rect 489458 263463 489514 263472
rect 486238 262168 486294 262177
rect 486238 262103 486294 262112
rect 483202 262032 483258 262041
rect 483202 261967 483258 261976
rect 480166 261896 480222 261905
rect 480166 261831 480222 261840
rect 477222 261760 477278 261769
rect 477222 261695 477278 261704
rect 473728 206984 473780 206990
rect 473728 206926 473780 206932
rect 489840 86193 489868 266591
rect 489826 86184 489882 86193
rect 489826 86119 489882 86128
rect 490576 6633 490604 266863
rect 490760 261905 490788 324935
rect 491956 299441 491984 431559
rect 492048 346361 492076 438087
rect 492140 387433 492168 440807
rect 493598 436792 493654 436801
rect 493598 436727 493654 436736
rect 493508 434784 493560 434790
rect 493508 434726 493560 434732
rect 493322 434072 493378 434081
rect 493322 434007 493378 434016
rect 492218 432576 492274 432585
rect 492218 432511 492274 432520
rect 492126 387424 492182 387433
rect 492126 387359 492182 387368
rect 492126 368112 492182 368121
rect 492126 368047 492182 368056
rect 492034 346352 492090 346361
rect 492034 346287 492090 346296
rect 492036 326052 492088 326058
rect 492036 325994 492088 326000
rect 491942 299432 491998 299441
rect 491942 299367 491998 299376
rect 492048 292777 492076 325994
rect 492140 295497 492168 368047
rect 492232 367033 492260 432511
rect 492218 367024 492274 367033
rect 492218 366959 492274 366968
rect 492218 347032 492274 347041
rect 492218 346967 492274 346976
rect 492126 295488 492182 295497
rect 492126 295423 492182 295432
rect 492232 294137 492260 346967
rect 492218 294128 492274 294137
rect 492218 294063 492274 294072
rect 492034 292768 492090 292777
rect 492034 292703 492090 292712
rect 491298 287736 491354 287745
rect 491298 287671 491354 287680
rect 490838 287464 490894 287473
rect 490838 287399 490894 287408
rect 490852 266665 490880 287399
rect 491312 282849 491340 287671
rect 491390 287328 491446 287337
rect 491390 287263 491446 287272
rect 491404 285190 491432 287263
rect 491392 285184 491444 285190
rect 491392 285126 491444 285132
rect 491298 282840 491354 282849
rect 491298 282775 491354 282784
rect 491404 277394 491432 285126
rect 493336 282713 493364 434007
rect 493414 396808 493470 396817
rect 493414 396743 493470 396752
rect 493322 282704 493378 282713
rect 493322 282639 493378 282648
rect 491312 277366 491432 277394
rect 491312 267734 491340 277366
rect 491312 267706 491984 267734
rect 490838 266656 490894 266665
rect 490838 266591 490894 266600
rect 491956 266393 491984 267706
rect 491942 266384 491998 266393
rect 491942 266319 491998 266328
rect 491206 265568 491262 265577
rect 491206 265503 491262 265512
rect 491220 262177 491248 265503
rect 491206 262168 491262 262177
rect 491206 262103 491262 262112
rect 490746 261896 490802 261905
rect 490746 261831 490802 261840
rect 491956 126041 491984 266319
rect 493428 261769 493456 396743
rect 493520 303550 493548 434726
rect 493612 325417 493640 436727
rect 496266 413400 496322 413409
rect 496266 413335 496322 413344
rect 494794 404832 494850 404841
rect 494794 404767 494850 404776
rect 494702 392592 494758 392601
rect 494702 392527 494758 392536
rect 493690 388104 493746 388113
rect 493690 388039 493746 388048
rect 493598 325408 493654 325417
rect 493598 325343 493654 325352
rect 493508 303544 493560 303550
rect 493508 303486 493560 303492
rect 493704 301481 493732 388039
rect 494716 370161 494744 392527
rect 494808 387569 494836 404767
rect 496174 402112 496230 402121
rect 496174 402047 496230 402056
rect 496082 393952 496138 393961
rect 496082 393887 496138 393896
rect 494794 387560 494850 387569
rect 494794 387495 494850 387504
rect 494702 370152 494758 370161
rect 494702 370087 494758 370096
rect 494702 361992 494758 362001
rect 494702 361927 494758 361936
rect 493690 301472 493746 301481
rect 493690 301407 493746 301416
rect 493506 290048 493562 290057
rect 493506 289983 493562 289992
rect 493520 284209 493548 289983
rect 494058 287192 494114 287201
rect 494058 287127 494114 287136
rect 493506 284200 493562 284209
rect 493506 284135 493562 284144
rect 494072 266529 494100 287127
rect 494716 282577 494744 361927
rect 494794 349752 494850 349761
rect 494794 349687 494850 349696
rect 494808 331401 494836 349687
rect 496096 334121 496124 393887
rect 496188 345001 496216 402047
rect 496280 371521 496308 413335
rect 496266 371512 496322 371521
rect 496266 371447 496322 371456
rect 496174 344992 496230 345001
rect 496174 344927 496230 344936
rect 496082 334112 496138 334121
rect 496082 334047 496138 334056
rect 494794 331392 494850 331401
rect 494794 331327 494850 331336
rect 497476 300801 497504 449375
rect 501602 447808 501658 447817
rect 501602 447743 501658 447752
rect 499026 433936 499082 433945
rect 499026 433871 499082 433880
rect 498934 410136 498990 410145
rect 498934 410071 498990 410080
rect 497554 403472 497610 403481
rect 497554 403407 497610 403416
rect 497568 366897 497596 403407
rect 498842 398032 498898 398041
rect 498842 397967 498898 397976
rect 497554 366888 497610 366897
rect 497554 366823 497610 366832
rect 497554 360632 497610 360641
rect 497554 360567 497610 360576
rect 497462 300792 497518 300801
rect 497462 300727 497518 300736
rect 494702 282568 494758 282577
rect 494702 282503 494758 282512
rect 494058 266520 494114 266529
rect 494058 266455 494114 266464
rect 494072 264217 494100 266455
rect 494058 264208 494114 264217
rect 494058 264143 494114 264152
rect 497568 262041 497596 360567
rect 498856 282441 498884 397967
rect 498948 298081 498976 410071
rect 499040 336841 499068 433871
rect 500222 413264 500278 413273
rect 500222 413199 500278 413208
rect 499118 344312 499174 344321
rect 499118 344247 499174 344256
rect 499026 336832 499082 336841
rect 499026 336767 499082 336776
rect 499132 324057 499160 344247
rect 500236 335481 500264 413199
rect 501616 372881 501644 447743
rect 538126 447264 538182 447273
rect 538126 447199 538182 447208
rect 541714 447264 541770 447273
rect 541714 447199 541770 447208
rect 535550 439376 535606 439385
rect 535550 439311 535606 439320
rect 535458 435296 535514 435305
rect 535458 435231 535514 435240
rect 535472 434790 535500 435231
rect 535460 434784 535512 434790
rect 535460 434726 535512 434732
rect 535564 432585 535592 439311
rect 535550 432576 535606 432585
rect 535550 432511 535606 432520
rect 536286 432576 536342 432585
rect 536286 432511 536342 432520
rect 536194 398848 536250 398857
rect 536194 398783 536250 398792
rect 536102 396128 536158 396137
rect 536102 396063 536158 396072
rect 501602 372872 501658 372881
rect 501602 372807 501658 372816
rect 535458 366072 535514 366081
rect 535458 366007 535514 366016
rect 535472 364993 535500 366007
rect 535458 364984 535514 364993
rect 535458 364919 535514 364928
rect 500222 335472 500278 335481
rect 500222 335407 500278 335416
rect 536116 325009 536144 396063
rect 536208 363662 536236 398783
rect 536300 396817 536328 432511
rect 536746 424416 536802 424425
rect 536746 424351 536802 424360
rect 536378 400344 536434 400353
rect 536378 400279 536434 400288
rect 536286 396808 536342 396817
rect 536286 396743 536342 396752
rect 536392 367305 536420 400279
rect 536760 396001 536788 424351
rect 538140 422929 538168 447199
rect 541728 445740 541756 447199
rect 538692 445182 539258 445210
rect 544226 445194 544608 445210
rect 544226 445188 544620 445194
rect 544226 445182 544568 445188
rect 538126 422920 538182 422929
rect 538126 422855 538182 422864
rect 538692 422294 538720 445182
rect 546710 445182 547368 445210
rect 544568 445130 544620 445136
rect 540978 422920 541034 422929
rect 540978 422855 541034 422864
rect 538692 422266 538904 422294
rect 538126 411360 538182 411369
rect 538126 411295 538182 411304
rect 536746 395992 536802 396001
rect 536746 395927 536802 395936
rect 536746 388376 536802 388385
rect 536746 388311 536802 388320
rect 536378 367296 536434 367305
rect 536378 367231 536434 367240
rect 536378 364712 536434 364721
rect 536378 364647 536434 364656
rect 536196 363656 536248 363662
rect 536196 363598 536248 363604
rect 536286 363352 536342 363361
rect 536286 363287 536342 363296
rect 536300 326466 536328 363287
rect 536392 344321 536420 364647
rect 536760 359281 536788 388311
rect 538140 387025 538168 411295
rect 538876 409170 538904 422266
rect 540992 411369 541020 422855
rect 545026 422376 545082 422385
rect 545026 422311 545082 422320
rect 545040 412634 545068 422311
rect 547340 412634 547368 445182
rect 547880 445188 547932 445194
rect 547880 445130 547932 445136
rect 547892 422385 547920 445130
rect 549258 434752 549314 434761
rect 549258 434687 549314 434696
rect 547878 422376 547934 422385
rect 547878 422311 547934 422320
rect 544672 412606 545068 412634
rect 547064 412606 547368 412634
rect 540978 411360 541034 411369
rect 540978 411295 541034 411304
rect 540992 409714 541020 411295
rect 540992 409686 541742 409714
rect 544672 409222 544700 412606
rect 547064 409714 547092 412606
rect 546710 409686 547368 409714
rect 544660 409216 544712 409222
rect 538876 409142 539258 409170
rect 544226 409164 544660 409170
rect 544226 409158 544712 409164
rect 544226 409142 544700 409158
rect 538876 409034 538904 409142
rect 538784 409006 538904 409034
rect 538784 393314 538812 409006
rect 547340 404977 547368 409686
rect 547880 409216 547932 409222
rect 547880 409158 547932 409164
rect 547326 404968 547382 404977
rect 547326 404903 547382 404912
rect 538692 393286 538812 393314
rect 538126 387016 538182 387025
rect 538126 386951 538182 386960
rect 538692 383654 538720 393286
rect 545026 387696 545082 387705
rect 545026 387631 545082 387640
rect 540978 387016 541034 387025
rect 540978 386951 541034 386960
rect 538692 383626 538812 383654
rect 538126 375456 538182 375465
rect 538126 375391 538182 375400
rect 536746 359272 536802 359281
rect 536746 359207 536802 359216
rect 536746 352472 536802 352481
rect 536746 352407 536802 352416
rect 536378 344312 536434 344321
rect 536378 344247 536434 344256
rect 536378 327312 536434 327321
rect 536378 327247 536434 327256
rect 536288 326460 536340 326466
rect 536288 326402 536340 326408
rect 536194 325952 536250 325961
rect 536194 325887 536250 325896
rect 536102 325000 536158 325009
rect 536102 324935 536158 324944
rect 499118 324048 499174 324057
rect 499118 323983 499174 323992
rect 536102 301472 536158 301481
rect 536102 301407 536158 301416
rect 498934 298072 498990 298081
rect 498934 298007 498990 298016
rect 536116 296721 536144 301407
rect 536102 296712 536158 296721
rect 536102 296647 536158 296656
rect 535460 292528 535512 292534
rect 535460 292470 535512 292476
rect 535472 291281 535500 292470
rect 535458 291272 535514 291281
rect 535458 291207 535514 291216
rect 536102 288552 536158 288561
rect 536102 288487 536158 288496
rect 498842 282432 498898 282441
rect 498842 282367 498898 282376
rect 504362 266792 504418 266801
rect 504362 266727 504418 266736
rect 497554 262032 497610 262041
rect 497554 261967 497610 261976
rect 493414 261760 493470 261769
rect 493414 261695 493470 261704
rect 491942 126032 491998 126041
rect 491942 125967 491998 125976
rect 504376 46345 504404 266727
rect 536116 263537 536144 288487
rect 536208 287745 536236 325887
rect 536286 324592 536342 324601
rect 536286 324527 536342 324536
rect 536194 287736 536250 287745
rect 536194 287671 536250 287680
rect 536300 265577 536328 324527
rect 536392 303618 536420 327247
rect 536760 323241 536788 352407
rect 538140 351121 538168 375391
rect 538784 373266 538812 383626
rect 540992 375465 541020 386951
rect 540978 375456 541034 375465
rect 540978 375391 541034 375400
rect 540992 373994 541020 375391
rect 540992 373966 541756 373994
rect 541728 373660 541756 373966
rect 545040 373402 545068 387631
rect 547340 373994 547368 404903
rect 547892 387705 547920 409158
rect 549272 398313 549300 434687
rect 549258 398304 549314 398313
rect 549258 398239 549314 398248
rect 547878 387696 547934 387705
rect 547878 387631 547934 387640
rect 544226 373374 545068 373402
rect 538784 373238 539258 373266
rect 545040 373250 545068 373374
rect 547064 373966 547368 373994
rect 547064 373266 547092 373966
rect 545028 373244 545080 373250
rect 538784 354674 538812 373238
rect 546710 373238 547092 373266
rect 545028 373186 545080 373192
rect 547064 364334 547092 373238
rect 548524 373244 548576 373250
rect 548524 373186 548576 373192
rect 547064 364306 547368 364334
rect 538692 354646 538812 354674
rect 538126 351112 538182 351121
rect 538126 351047 538182 351056
rect 538692 345014 538720 354646
rect 540978 351112 541034 351121
rect 540978 351047 541034 351056
rect 540992 345014 541020 351047
rect 547340 345014 547368 364306
rect 548536 351937 548564 373186
rect 549272 362817 549300 398239
rect 549258 362808 549314 362817
rect 549258 362743 549314 362752
rect 548522 351928 548578 351937
rect 548522 351863 548578 351872
rect 538692 344986 538904 345014
rect 540992 344986 541296 345014
rect 538126 339552 538182 339561
rect 538126 339487 538182 339496
rect 536746 323232 536802 323241
rect 536746 323167 536802 323176
rect 536746 316432 536802 316441
rect 536746 316367 536802 316376
rect 536380 303612 536432 303618
rect 536380 303554 536432 303560
rect 536760 287201 536788 316367
rect 538140 315353 538168 339487
rect 538876 337770 538904 344986
rect 541268 339561 541296 344986
rect 547064 344986 547368 345014
rect 541254 339552 541310 339561
rect 541254 339487 541310 339496
rect 544198 339552 544254 339561
rect 544198 339487 544254 339496
rect 541268 337770 541296 339487
rect 538784 337742 539258 337770
rect 541268 337742 541742 337770
rect 544212 337756 544240 339487
rect 547064 337770 547092 344986
rect 548536 339561 548564 351863
rect 547878 339552 547934 339561
rect 547878 339487 547934 339496
rect 548522 339552 548578 339561
rect 548522 339487 548578 339496
rect 546710 337742 547092 337770
rect 538784 316034 538812 337742
rect 547064 335354 547092 337742
rect 547064 335326 547368 335354
rect 538784 316006 538904 316034
rect 538126 315344 538182 315353
rect 538126 315279 538182 315288
rect 538876 306374 538904 316006
rect 541714 315344 541770 315353
rect 541714 315279 541770 315288
rect 538876 306346 539272 306374
rect 539244 303657 539272 306346
rect 541728 303793 541756 315279
rect 547340 306374 547368 335326
rect 547064 306346 547368 306374
rect 544198 305008 544254 305017
rect 544198 304943 544254 304952
rect 541714 303784 541770 303793
rect 541714 303719 541770 303728
rect 539230 303648 539286 303657
rect 539230 303583 539286 303592
rect 539244 301716 539272 303583
rect 541728 301716 541756 303719
rect 544212 301716 544240 304943
rect 547064 301730 547092 306346
rect 547892 305017 547920 339487
rect 549272 326777 549300 362743
rect 549258 326768 549314 326777
rect 549258 326703 549314 326712
rect 547878 305008 547934 305017
rect 547878 304943 547934 304952
rect 549166 303784 549222 303793
rect 549166 303719 549222 303728
rect 548522 303648 548578 303657
rect 548522 303583 548578 303592
rect 546710 301702 547092 301730
rect 536746 287192 536802 287201
rect 536746 287127 536802 287136
rect 548536 282169 548564 303583
rect 549180 298761 549208 303719
rect 549166 298752 549222 298761
rect 549166 298687 549222 298696
rect 549272 290737 549300 326703
rect 549258 290728 549314 290737
rect 549258 290663 549314 290672
rect 549902 290728 549958 290737
rect 549902 290663 549958 290672
rect 548522 282160 548578 282169
rect 548522 282095 548578 282104
rect 536746 280392 536802 280401
rect 536746 280327 536802 280336
rect 536286 265568 536342 265577
rect 536286 265503 536342 265512
rect 536102 263528 536158 263537
rect 536102 263463 536158 263472
rect 536760 212838 536788 280327
rect 536748 212832 536800 212838
rect 536748 212774 536800 212780
rect 504362 46336 504418 46345
rect 504362 46271 504418 46280
rect 549916 19825 549944 290663
rect 580354 282160 580410 282169
rect 580354 282095 580410 282104
rect 580262 264208 580318 264217
rect 580262 264143 580318 264152
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580276 165889 580304 264143
rect 580368 245585 580396 282095
rect 580354 245576 580410 245585
rect 580354 245511 580410 245520
rect 580262 165880 580318 165889
rect 580262 165815 580318 165824
rect 549902 19816 549958 19825
rect 549902 19751 549958 19760
rect 490562 6624 490618 6633
rect 490562 6559 490618 6568
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 470138 451560 470194 451616
rect 488906 451560 488962 451616
rect 469036 450097 469572 450393
rect 469036 431697 469572 431993
rect 470276 451183 470812 451479
rect 470276 449012 470812 449308
rect 470276 432784 470812 433080
rect 481160 450744 481216 450800
rect 476061 450608 476117 450664
rect 478694 447888 478750 447944
rect 482006 447752 482062 447808
rect 475382 444896 475438 444952
rect 481546 434968 481602 435024
rect 470276 430612 470812 430908
rect 470138 429800 470194 429856
rect 470276 411784 470812 412080
rect 471886 434560 471942 434616
rect 473358 434560 473414 434616
rect 483202 435104 483258 435160
rect 488814 449433 488816 449440
rect 488816 449433 488868 449440
rect 488868 449433 488870 449440
rect 488814 449384 488870 449433
rect 497462 449384 497518 449440
rect 490562 447888 490618 447944
rect 488998 435104 489054 435160
rect 488906 434968 488962 435024
rect 488446 434560 488502 434616
rect 485318 433880 485374 433936
rect 477958 429800 478014 429856
rect 475474 429120 475530 429176
rect 471518 412256 471574 412312
rect 469036 410698 469572 410994
rect 470276 409612 470812 409908
rect 470138 392536 470194 392592
rect 469036 389702 469572 389998
rect 470276 390785 470812 391081
rect 479246 428440 479302 428496
rect 489090 431568 489146 431624
rect 483202 430616 483258 430672
rect 484306 430616 484362 430672
rect 482374 413344 482430 413400
rect 481086 412664 481142 412720
rect 477774 412256 477830 412312
rect 485870 430344 485926 430400
rect 489274 428440 489330 428496
rect 488538 413888 488594 413944
rect 485870 413208 485926 413264
rect 484306 412256 484362 412312
rect 477774 411848 477830 411904
rect 481086 411848 481142 411904
rect 484306 411848 484362 411904
rect 471518 392536 471574 392592
rect 471518 391992 471574 392048
rect 477682 411576 477738 411632
rect 481086 411576 481142 411632
rect 484306 411576 484362 411632
rect 488722 412256 488778 412312
rect 475290 408448 475346 408504
rect 488538 410085 488594 410136
rect 488538 410080 488540 410085
rect 488540 410080 488592 410085
rect 488592 410080 488594 410085
rect 478694 406136 478750 406192
rect 485226 393896 485282 393952
rect 481822 392536 481878 392592
rect 489642 434560 489698 434616
rect 489642 413888 489698 413944
rect 489458 412664 489514 412720
rect 490746 443536 490802 443592
rect 490654 442176 490710 442232
rect 490562 408856 490618 408912
rect 492126 440816 492182 440872
rect 492034 438096 492090 438152
rect 491942 431568 491998 431624
rect 490746 429120 490802 429176
rect 490654 408448 490710 408504
rect 489274 407496 489330 407552
rect 482558 392128 482614 392184
rect 488538 392128 488594 392184
rect 477866 391992 477922 392048
rect 488630 391992 488686 392048
rect 490746 392128 490802 392184
rect 477866 390904 477922 390960
rect 482558 390904 482614 390960
rect 489182 390904 489238 390960
rect 478050 390632 478106 390688
rect 482374 390632 482430 390688
rect 489458 390632 489514 390688
rect 470276 388612 470812 388908
rect 471610 371320 471666 371376
rect 470138 370232 470194 370288
rect 470276 369785 470812 370081
rect 475750 387640 475806 387696
rect 479614 387504 479670 387560
rect 483202 386416 483258 386472
rect 485686 382336 485742 382392
rect 482374 371864 482430 371920
rect 473726 371320 473782 371376
rect 473266 370232 473322 370288
rect 469036 368699 469572 368995
rect 470276 367612 470812 367908
rect 489550 386416 489606 386472
rect 486882 372000 486938 372056
rect 482374 369824 482430 369880
rect 485686 369824 485742 369880
rect 478878 369552 478934 369608
rect 481822 369552 481878 369608
rect 485318 369552 485374 369608
rect 473266 359488 473322 359544
rect 470276 348784 470812 349080
rect 477222 366968 477278 367024
rect 480166 366832 480222 366888
rect 483202 366696 483258 366752
rect 476118 359488 476174 359544
rect 473726 350512 473782 350568
rect 471702 349152 471758 349208
rect 473358 349152 473414 349208
rect 469036 347697 469572 347993
rect 470276 346612 470812 346908
rect 470276 327784 470812 328080
rect 481270 350512 481326 350568
rect 490654 372000 490710 372056
rect 489550 368736 489606 368792
rect 489458 368084 489514 368112
rect 489458 368056 489460 368084
rect 489460 368056 489512 368084
rect 489512 368056 489514 368084
rect 489366 367240 489422 367296
rect 488814 350648 488870 350704
rect 486422 349696 486478 349752
rect 476118 348744 476174 348800
rect 481270 348744 481326 348800
rect 475658 348508 475660 348528
rect 475660 348508 475712 348528
rect 475712 348508 475714 348528
rect 475658 348472 475714 348508
rect 474186 348336 474242 348392
rect 481232 348336 481288 348392
rect 471702 342216 471758 342272
rect 488906 350512 488962 350568
rect 475566 346296 475622 346352
rect 478602 344936 478658 344992
rect 482190 344800 482246 344856
rect 474646 342216 474702 342272
rect 469036 326697 469572 326993
rect 470276 325612 470812 325908
rect 470276 306784 470812 307080
rect 471610 329840 471666 329896
rect 471518 326848 471574 326904
rect 485410 329976 485466 330032
rect 481546 329840 481602 329896
rect 488998 347012 489000 347032
rect 489000 347012 489052 347032
rect 489052 347012 489054 347032
rect 488998 346976 489054 347012
rect 489642 350648 489698 350704
rect 488906 329840 488962 329896
rect 474646 327800 474702 327856
rect 481546 327800 481602 327856
rect 485410 327800 485466 327856
rect 471702 327664 471758 327720
rect 471610 308352 471666 308408
rect 471518 307808 471574 307864
rect 469036 305699 469572 305995
rect 470276 304612 470812 304908
rect 474653 327392 474709 327448
rect 481542 327392 481598 327448
rect 484986 327392 485042 327448
rect 476210 326848 476266 326904
rect 475474 325352 475530 325408
rect 479062 324128 479118 324184
rect 482374 323992 482430 324048
rect 489918 328616 489974 328672
rect 489642 324128 489698 324184
rect 489918 326848 489974 326904
rect 488630 313248 488686 313304
rect 480902 308352 480958 308408
rect 488538 308352 488594 308408
rect 477498 307808 477554 307864
rect 477498 306856 477554 306912
rect 480902 306856 480958 306912
rect 477590 306584 477646 306640
rect 480902 306584 480958 306640
rect 484306 306584 484362 306640
rect 471518 287272 471574 287328
rect 470276 285785 470812 286081
rect 469036 284700 469572 284996
rect 470276 283612 470812 283908
rect 488630 306720 488686 306776
rect 482558 287408 482614 287464
rect 488538 287408 488594 287464
rect 477866 287272 477922 287328
rect 471610 287136 471666 287192
rect 474738 287136 474794 287192
rect 471518 266736 471574 266792
rect 489642 313248 489698 313304
rect 488630 287272 488686 287328
rect 490838 391992 490894 392048
rect 490838 382336 490894 382392
rect 490746 371864 490802 371920
rect 490746 364928 490802 364984
rect 490746 344800 490802 344856
rect 490654 332696 490710 332752
rect 490746 324944 490802 325000
rect 489274 287136 489330 287192
rect 474738 285912 474794 285968
rect 477866 285912 477922 285968
rect 482558 285912 482614 285968
rect 489274 285912 489330 285968
rect 474738 285640 474794 285696
rect 478050 285640 478106 285696
rect 482374 285640 482430 285696
rect 489274 285640 489330 285696
rect 475750 282648 475806 282704
rect 486882 282784 486938 282840
rect 483202 282512 483258 282568
rect 479614 282376 479670 282432
rect 476118 266872 476174 266928
rect 490562 266872 490618 266928
rect 471610 266328 471666 266384
rect 479062 266736 479118 266792
rect 470276 264785 470812 265081
rect 476118 266328 476174 266384
rect 482558 266600 482614 266656
rect 489826 266600 489882 266656
rect 488446 266464 488502 266520
rect 485318 266328 485374 266384
rect 476118 264832 476174 264888
rect 479062 264832 479118 264888
rect 482558 264832 482614 264888
rect 485318 264832 485374 264888
rect 488446 264832 488502 264888
rect 476118 264560 476174 264616
rect 479062 264560 479118 264616
rect 482374 264560 482430 264616
rect 485410 264560 485466 264616
rect 488446 264560 488502 264616
rect 469036 263699 469572 263995
rect 470276 262612 470812 262908
rect 489458 263472 489514 263528
rect 486238 262112 486294 262168
rect 483202 261976 483258 262032
rect 480166 261840 480222 261896
rect 477222 261704 477278 261760
rect 489826 86128 489882 86184
rect 493598 436736 493654 436792
rect 493322 434016 493378 434072
rect 492218 432520 492274 432576
rect 492126 387368 492182 387424
rect 492126 368056 492182 368112
rect 492034 346296 492090 346352
rect 491942 299376 491998 299432
rect 492218 366968 492274 367024
rect 492218 346976 492274 347032
rect 492126 295432 492182 295488
rect 492218 294072 492274 294128
rect 492034 292712 492090 292768
rect 491298 287680 491354 287736
rect 490838 287408 490894 287464
rect 491390 287272 491446 287328
rect 491298 282784 491354 282840
rect 493414 396752 493470 396808
rect 493322 282648 493378 282704
rect 490838 266600 490894 266656
rect 491942 266328 491998 266384
rect 491206 265512 491262 265568
rect 491206 262112 491262 262168
rect 490746 261840 490802 261896
rect 496266 413344 496322 413400
rect 494794 404776 494850 404832
rect 494702 392536 494758 392592
rect 493690 388048 493746 388104
rect 493598 325352 493654 325408
rect 496174 402056 496230 402112
rect 496082 393896 496138 393952
rect 494794 387504 494850 387560
rect 494702 370096 494758 370152
rect 494702 361936 494758 361992
rect 493690 301416 493746 301472
rect 493506 289992 493562 290048
rect 494058 287136 494114 287192
rect 493506 284144 493562 284200
rect 494794 349696 494850 349752
rect 496266 371456 496322 371512
rect 496174 344936 496230 344992
rect 496082 334056 496138 334112
rect 494794 331336 494850 331392
rect 501602 447752 501658 447808
rect 499026 433880 499082 433936
rect 498934 410080 498990 410136
rect 497554 403416 497610 403472
rect 498842 397976 498898 398032
rect 497554 366832 497610 366888
rect 497554 360576 497610 360632
rect 497462 300736 497518 300792
rect 494702 282512 494758 282568
rect 494058 266464 494114 266520
rect 494058 264152 494114 264208
rect 500222 413208 500278 413264
rect 499118 344256 499174 344312
rect 499026 336776 499082 336832
rect 538126 447208 538182 447264
rect 541714 447208 541770 447264
rect 535550 439320 535606 439376
rect 535458 435240 535514 435296
rect 535550 432520 535606 432576
rect 536286 432520 536342 432576
rect 536194 398792 536250 398848
rect 536102 396072 536158 396128
rect 501602 372816 501658 372872
rect 535458 366016 535514 366072
rect 535458 364928 535514 364984
rect 500222 335416 500278 335472
rect 536746 424360 536802 424416
rect 536378 400288 536434 400344
rect 536286 396752 536342 396808
rect 538126 422864 538182 422920
rect 540978 422864 541034 422920
rect 538126 411304 538182 411360
rect 536746 395936 536802 395992
rect 536746 388320 536802 388376
rect 536378 367240 536434 367296
rect 536378 364656 536434 364712
rect 536286 363296 536342 363352
rect 545026 422320 545082 422376
rect 549258 434696 549314 434752
rect 547878 422320 547934 422376
rect 540978 411304 541034 411360
rect 547326 404912 547382 404968
rect 538126 386960 538182 387016
rect 545026 387640 545082 387696
rect 540978 386960 541034 387016
rect 538126 375400 538182 375456
rect 536746 359216 536802 359272
rect 536746 352416 536802 352472
rect 536378 344256 536434 344312
rect 536378 327256 536434 327312
rect 536194 325896 536250 325952
rect 536102 324944 536158 325000
rect 499118 323992 499174 324048
rect 536102 301416 536158 301472
rect 498934 298016 498990 298072
rect 536102 296656 536158 296712
rect 535458 291216 535514 291272
rect 536102 288496 536158 288552
rect 498842 282376 498898 282432
rect 504362 266736 504418 266792
rect 497554 261976 497610 262032
rect 493414 261704 493470 261760
rect 491942 125976 491998 126032
rect 536286 324536 536342 324592
rect 536194 287680 536250 287736
rect 540978 375400 541034 375456
rect 549258 398248 549314 398304
rect 547878 387640 547934 387696
rect 538126 351056 538182 351112
rect 540978 351056 541034 351112
rect 549258 362752 549314 362808
rect 548522 351872 548578 351928
rect 538126 339496 538182 339552
rect 536746 323176 536802 323232
rect 536746 316376 536802 316432
rect 541254 339496 541310 339552
rect 544198 339496 544254 339552
rect 547878 339496 547934 339552
rect 548522 339496 548578 339552
rect 538126 315288 538182 315344
rect 541714 315288 541770 315344
rect 544198 304952 544254 305008
rect 541714 303728 541770 303784
rect 539230 303592 539286 303648
rect 549258 326712 549314 326768
rect 547878 304952 547934 305008
rect 549166 303728 549222 303784
rect 548522 303592 548578 303648
rect 536746 287136 536802 287192
rect 549166 298696 549222 298752
rect 549258 290672 549314 290728
rect 549902 290672 549958 290728
rect 548522 282104 548578 282160
rect 536746 280336 536802 280392
rect 536286 265512 536342 265568
rect 536102 263472 536158 263528
rect 504362 46280 504418 46336
rect 580354 282104 580410 282160
rect 580262 264152 580318 264208
rect 580170 205672 580226 205728
rect 580354 245520 580410 245576
rect 580262 165824 580318 165880
rect 549902 19760 549958 19816
rect 490562 6568 490618 6624
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect 470133 451618 470199 451621
rect 488901 451618 488967 451621
rect 470133 451616 475762 451618
rect 470133 451560 470138 451616
rect 470194 451560 475762 451616
rect 470133 451558 475762 451560
rect 470133 451555 470199 451558
rect 470266 451483 470822 451484
rect 470266 451179 470272 451483
rect 470816 451179 470822 451483
rect 470266 451178 470822 451179
rect 475702 450666 475762 451558
rect 481406 451616 488967 451618
rect 481406 451560 488906 451616
rect 488962 451560 488967 451616
rect 481406 451558 488967 451560
rect 481155 450802 481221 450805
rect 481406 450802 481466 451558
rect 488901 451555 488967 451558
rect 481155 450800 481466 450802
rect 481155 450744 481160 450800
rect 481216 450744 481466 450800
rect 481155 450742 481466 450744
rect 481155 450739 481221 450742
rect 476056 450666 476122 450669
rect 475702 450664 476122 450666
rect 475702 450608 476061 450664
rect 476117 450608 476122 450664
rect 475702 450606 476122 450608
rect 476056 450603 476122 450606
rect 469026 450397 469582 450398
rect 469026 450093 469032 450397
rect 469576 450093 469582 450397
rect 469026 450092 469582 450093
rect -960 449428 480 449668
rect 488809 449442 488875 449445
rect 497457 449442 497523 449445
rect 488809 449440 497523 449442
rect 488809 449384 488814 449440
rect 488870 449384 497462 449440
rect 497518 449384 497523 449440
rect 488809 449382 497523 449384
rect 488809 449379 488875 449382
rect 497457 449379 497523 449382
rect 470266 449312 470822 449313
rect 470266 449008 470272 449312
rect 470816 449008 470822 449312
rect 470266 449007 470822 449008
rect 478689 447946 478755 447949
rect 490557 447946 490623 447949
rect 478689 447944 490623 447946
rect 478689 447888 478694 447944
rect 478750 447888 490562 447944
rect 490618 447888 490623 447944
rect 478689 447886 490623 447888
rect 478689 447883 478755 447886
rect 490557 447883 490623 447886
rect 482001 447810 482067 447813
rect 501597 447810 501663 447813
rect 482001 447808 501663 447810
rect 482001 447752 482006 447808
rect 482062 447752 501602 447808
rect 501658 447752 501663 447808
rect 482001 447750 501663 447752
rect 482001 447747 482067 447750
rect 501597 447747 501663 447750
rect 538121 447266 538187 447269
rect 541709 447266 541775 447269
rect 538121 447264 541775 447266
rect 538121 447208 538126 447264
rect 538182 447208 541714 447264
rect 541770 447208 541775 447264
rect 538121 447206 541775 447208
rect 538121 447203 538187 447206
rect 541709 447203 541775 447206
rect 475377 444954 475443 444957
rect 475377 444952 528570 444954
rect 475377 444896 475382 444952
rect 475438 444896 528570 444952
rect 475377 444894 528570 444896
rect 475377 444891 475443 444894
rect 528510 444818 528570 444894
rect 528510 444758 538108 444818
rect 583520 444668 584960 444908
rect 490741 443594 490807 443597
rect 490741 443592 528570 443594
rect 490741 443536 490746 443592
rect 490802 443536 528570 443592
rect 490741 443534 528570 443536
rect 490741 443531 490807 443534
rect 528510 443458 528570 443534
rect 528510 443398 538108 443458
rect 490649 442234 490715 442237
rect 490649 442232 528570 442234
rect 490649 442176 490654 442232
rect 490710 442176 528570 442232
rect 490649 442174 528570 442176
rect 490649 442171 490715 442174
rect 528510 442098 528570 442174
rect 528510 442038 538108 442098
rect 492121 440874 492187 440877
rect 492121 440872 528570 440874
rect 492121 440816 492126 440872
rect 492182 440816 528570 440872
rect 492121 440814 528570 440816
rect 492121 440811 492187 440814
rect 528510 440738 528570 440814
rect 528510 440678 538108 440738
rect 535545 439378 535611 439381
rect 535545 439376 538108 439378
rect 535545 439320 535550 439376
rect 535606 439320 538108 439376
rect 535545 439318 538108 439320
rect 535545 439315 535611 439318
rect 492029 438154 492095 438157
rect 492029 438152 528570 438154
rect 492029 438096 492034 438152
rect 492090 438096 528570 438152
rect 492029 438094 528570 438096
rect 492029 438091 492095 438094
rect 528510 438018 528570 438094
rect 528510 437958 538108 438018
rect 493593 436794 493659 436797
rect 493593 436792 528570 436794
rect -960 436508 480 436748
rect 493593 436736 493598 436792
rect 493654 436736 528570 436792
rect 493593 436734 528570 436736
rect 493593 436731 493659 436734
rect 528510 436658 528570 436734
rect 528510 436598 538108 436658
rect 535453 435298 535519 435301
rect 535453 435296 538108 435298
rect 535453 435240 535458 435296
rect 535514 435240 538108 435296
rect 535453 435238 538108 435240
rect 535453 435235 535519 435238
rect 483197 435162 483263 435165
rect 488993 435162 489059 435165
rect 483197 435160 489059 435162
rect 483197 435104 483202 435160
rect 483258 435104 488998 435160
rect 489054 435104 489059 435160
rect 483197 435102 489059 435104
rect 483197 435099 483263 435102
rect 488993 435099 489059 435102
rect 481541 435026 481607 435029
rect 488901 435026 488967 435029
rect 481541 435024 488967 435026
rect 481541 434968 481546 435024
rect 481602 434968 488906 435024
rect 488962 434968 488967 435024
rect 481541 434966 488967 434968
rect 481541 434963 481607 434966
rect 488901 434963 488967 434966
rect 549253 434754 549319 434757
rect 547860 434752 549319 434754
rect 547860 434696 549258 434752
rect 549314 434696 549319 434752
rect 547860 434694 549319 434696
rect 549253 434691 549319 434694
rect 471881 434618 471947 434621
rect 473353 434618 473419 434621
rect 471881 434616 473419 434618
rect 471881 434560 471886 434616
rect 471942 434560 473358 434616
rect 473414 434560 473419 434616
rect 471881 434558 473419 434560
rect 471881 434555 471947 434558
rect 473353 434555 473419 434558
rect 488441 434618 488507 434621
rect 489637 434618 489703 434621
rect 488441 434616 489703 434618
rect 488441 434560 488446 434616
rect 488502 434560 489642 434616
rect 489698 434560 489703 434616
rect 488441 434558 489703 434560
rect 488441 434555 488507 434558
rect 489637 434555 489703 434558
rect 493317 434074 493383 434077
rect 493317 434072 528570 434074
rect 493317 434016 493322 434072
rect 493378 434016 528570 434072
rect 493317 434014 528570 434016
rect 493317 434011 493383 434014
rect 485313 433938 485379 433941
rect 499021 433938 499087 433941
rect 485313 433936 499087 433938
rect 485313 433880 485318 433936
rect 485374 433880 499026 433936
rect 499082 433880 499087 433936
rect 485313 433878 499087 433880
rect 528510 433938 528570 434014
rect 528510 433878 538108 433938
rect 485313 433875 485379 433878
rect 499021 433875 499087 433878
rect 470266 433084 470822 433085
rect 470266 432780 470272 433084
rect 470816 432780 470822 433084
rect 470266 432779 470822 432780
rect 492213 432578 492279 432581
rect 535545 432578 535611 432581
rect 492213 432576 535611 432578
rect 492213 432520 492218 432576
rect 492274 432520 535550 432576
rect 535606 432520 535611 432576
rect 492213 432518 535611 432520
rect 492213 432515 492279 432518
rect 535545 432515 535611 432518
rect 536281 432578 536347 432581
rect 536281 432576 538108 432578
rect 536281 432520 536286 432576
rect 536342 432520 538108 432576
rect 536281 432518 538108 432520
rect 536281 432515 536347 432518
rect 469026 431997 469582 431998
rect 469026 431693 469032 431997
rect 469576 431693 469582 431997
rect 469026 431692 469582 431693
rect 489085 431626 489151 431629
rect 491937 431626 492003 431629
rect 489085 431624 492003 431626
rect 489085 431568 489090 431624
rect 489146 431568 491942 431624
rect 491998 431568 492003 431624
rect 489085 431566 492003 431568
rect 489085 431563 489151 431566
rect 491937 431563 492003 431566
rect 583520 431476 584960 431716
rect 470266 430912 470822 430913
rect 470266 430608 470272 430912
rect 470816 430608 470822 430912
rect 483197 430674 483263 430677
rect 484301 430674 484367 430677
rect 483197 430672 484367 430674
rect 483197 430616 483202 430672
rect 483258 430616 484306 430672
rect 484362 430616 484367 430672
rect 483197 430614 484367 430616
rect 483197 430611 483263 430614
rect 484301 430611 484367 430614
rect 470266 430607 470822 430608
rect 485822 430405 485882 430644
rect 485822 430400 485931 430405
rect 485822 430344 485870 430400
rect 485926 430344 485931 430400
rect 485822 430342 485931 430344
rect 485865 430339 485931 430342
rect 470133 429858 470199 429861
rect 477953 429858 478019 429861
rect 470133 429856 478019 429858
rect 470133 429800 470138 429856
rect 470194 429800 477958 429856
rect 478014 429800 478019 429856
rect 470133 429798 478019 429800
rect 470133 429795 470199 429798
rect 477953 429795 478019 429798
rect 475469 429178 475535 429181
rect 490741 429178 490807 429181
rect 475469 429176 490807 429178
rect 475469 429120 475474 429176
rect 475530 429120 490746 429176
rect 490802 429120 490807 429176
rect 475469 429118 490807 429120
rect 475469 429115 475535 429118
rect 490741 429115 490807 429118
rect 479241 428498 479307 428501
rect 489269 428498 489335 428501
rect 479241 428496 489335 428498
rect 479241 428440 479246 428496
rect 479302 428440 489274 428496
rect 489330 428440 489335 428496
rect 479241 428438 489335 428440
rect 479241 428435 479307 428438
rect 489269 428435 489335 428438
rect 536741 424418 536807 424421
rect 538078 424418 538138 431188
rect 536741 424416 538138 424418
rect 536741 424360 536746 424416
rect 536802 424388 538138 424416
rect 536802 424360 538108 424388
rect 536741 424358 538108 424360
rect 536741 424355 536807 424358
rect -960 423452 480 423692
rect 538121 422922 538187 422925
rect 540973 422922 541039 422925
rect 538121 422920 541039 422922
rect 538121 422864 538126 422920
rect 538182 422864 540978 422920
rect 541034 422864 541039 422920
rect 538121 422862 541039 422864
rect 538121 422859 538187 422862
rect 540973 422859 541039 422862
rect 545021 422378 545087 422381
rect 547873 422378 547939 422381
rect 545021 422376 547939 422378
rect 545021 422320 545026 422376
rect 545082 422320 547878 422376
rect 547934 422320 547939 422376
rect 545021 422318 547939 422320
rect 545021 422315 545087 422318
rect 547873 422315 547939 422318
rect 583520 418148 584960 418388
rect 488533 413946 488599 413949
rect 489637 413946 489703 413949
rect 488533 413944 489703 413946
rect 488533 413888 488538 413944
rect 488594 413888 489642 413944
rect 489698 413888 489703 413944
rect 488533 413886 489703 413888
rect 488533 413883 488599 413886
rect 489637 413883 489703 413886
rect 482369 413402 482435 413405
rect 496261 413402 496327 413405
rect 482369 413400 496327 413402
rect 482369 413344 482374 413400
rect 482430 413344 496266 413400
rect 496322 413344 496327 413400
rect 482369 413342 496327 413344
rect 482369 413339 482435 413342
rect 496261 413339 496327 413342
rect 485865 413266 485931 413269
rect 500217 413266 500283 413269
rect 485865 413264 500283 413266
rect 485865 413208 485870 413264
rect 485926 413208 500222 413264
rect 500278 413208 500283 413264
rect 485865 413206 500283 413208
rect 485865 413203 485931 413206
rect 500217 413203 500283 413206
rect 481081 412722 481147 412725
rect 489453 412722 489519 412725
rect 481081 412720 489519 412722
rect 481081 412664 481086 412720
rect 481142 412664 489458 412720
rect 489514 412664 489519 412720
rect 481081 412662 489519 412664
rect 481081 412659 481147 412662
rect 489453 412659 489519 412662
rect 471513 412314 471579 412317
rect 477769 412314 477835 412317
rect 471513 412312 477835 412314
rect 471513 412256 471518 412312
rect 471574 412256 477774 412312
rect 477830 412256 477835 412312
rect 471513 412254 477835 412256
rect 471513 412251 471579 412254
rect 477769 412251 477835 412254
rect 484301 412314 484367 412317
rect 488717 412314 488783 412317
rect 484301 412312 488783 412314
rect 484301 412256 484306 412312
rect 484362 412256 488722 412312
rect 488778 412256 488783 412312
rect 484301 412254 488783 412256
rect 484301 412251 484367 412254
rect 488717 412251 488783 412254
rect 470266 412084 470822 412085
rect 470266 411780 470272 412084
rect 470816 411780 470822 412084
rect 477769 411906 477835 411909
rect 470266 411779 470822 411780
rect 477726 411904 477835 411906
rect 477726 411848 477774 411904
rect 477830 411848 477835 411904
rect 477726 411843 477835 411848
rect 481081 411904 481147 411909
rect 481081 411848 481086 411904
rect 481142 411848 481147 411904
rect 481081 411843 481147 411848
rect 484301 411906 484367 411909
rect 484301 411904 484410 411906
rect 484301 411848 484306 411904
rect 484362 411848 484410 411904
rect 484301 411843 484410 411848
rect 477726 411637 477786 411843
rect 481084 411637 481144 411843
rect 484350 411637 484410 411843
rect 477677 411632 477786 411637
rect 477677 411576 477682 411632
rect 477738 411576 477786 411632
rect 477677 411574 477786 411576
rect 481081 411632 481147 411637
rect 481081 411576 481086 411632
rect 481142 411576 481147 411632
rect 477677 411571 477743 411574
rect 481081 411571 481147 411576
rect 484301 411632 484410 411637
rect 484301 411576 484306 411632
rect 484362 411576 484410 411632
rect 484301 411574 484410 411576
rect 484301 411571 484367 411574
rect 538121 411362 538187 411365
rect 540973 411362 541039 411365
rect 538121 411360 541039 411362
rect 538121 411304 538126 411360
rect 538182 411304 540978 411360
rect 541034 411304 541039 411360
rect 538121 411302 541039 411304
rect 538121 411299 538187 411302
rect 540973 411299 541039 411302
rect 469026 410998 469582 410999
rect 469026 410694 469032 410998
rect 469576 410694 469582 410998
rect 469026 410693 469582 410694
rect -960 410396 480 410636
rect 488533 410138 488599 410141
rect 498929 410138 498995 410141
rect 488533 410136 498995 410138
rect 488533 410080 488538 410136
rect 488594 410080 498934 410136
rect 498990 410080 498995 410136
rect 488533 410078 498995 410080
rect 488533 410075 488599 410078
rect 498929 410075 498995 410078
rect 470266 409912 470822 409913
rect 470266 409608 470272 409912
rect 470816 409608 470822 409912
rect 470266 409607 470822 409608
rect 490557 408914 490623 408917
rect 490557 408912 538138 408914
rect 490557 408856 490562 408912
rect 490618 408856 538138 408912
rect 490557 408854 538138 408856
rect 490557 408851 490623 408854
rect 538078 408816 538138 408854
rect 475285 408506 475351 408509
rect 490649 408506 490715 408509
rect 475285 408504 490715 408506
rect 475285 408448 475290 408504
rect 475346 408448 490654 408504
rect 490710 408448 490715 408504
rect 475285 408446 490715 408448
rect 475285 408443 475351 408446
rect 490649 408443 490715 408446
rect 489269 407554 489335 407557
rect 489269 407552 538138 407554
rect 489269 407496 489274 407552
rect 489330 407496 538138 407552
rect 489269 407494 538138 407496
rect 489269 407491 489335 407494
rect 538078 407456 538138 407494
rect 478689 406194 478755 406197
rect 478689 406192 538138 406194
rect 478689 406136 478694 406192
rect 478750 406136 538138 406192
rect 478689 406134 538138 406136
rect 478689 406131 478755 406134
rect 538078 406096 538138 406134
rect 547321 404970 547387 404973
rect 583520 404970 584960 405060
rect 547321 404968 584960 404970
rect 547321 404912 547326 404968
rect 547382 404912 584960 404968
rect 547321 404910 584960 404912
rect 547321 404907 547387 404910
rect 494789 404834 494855 404837
rect 494789 404832 538138 404834
rect 494789 404776 494794 404832
rect 494850 404776 538138 404832
rect 583520 404820 584960 404910
rect 494789 404774 538138 404776
rect 494789 404771 494855 404774
rect 538078 404736 538138 404774
rect 497549 403474 497615 403477
rect 497549 403472 538138 403474
rect 497549 403416 497554 403472
rect 497610 403416 538138 403472
rect 497549 403414 538138 403416
rect 497549 403411 497615 403414
rect 538078 403376 538138 403414
rect 496169 402114 496235 402117
rect 496169 402112 538138 402114
rect 496169 402056 496174 402112
rect 496230 402056 538138 402112
rect 496169 402054 538138 402056
rect 496169 402051 496235 402054
rect 538078 402016 538138 402054
rect 536373 400346 536439 400349
rect 538078 400346 538138 400656
rect 536373 400344 538138 400346
rect 536373 400288 536378 400344
rect 536434 400288 538138 400344
rect 536373 400286 538138 400288
rect 536373 400283 536439 400286
rect 536189 398850 536255 398853
rect 538078 398850 538138 399296
rect 536189 398848 538138 398850
rect 536189 398792 536194 398848
rect 536250 398792 538138 398848
rect 536189 398790 538138 398792
rect 536189 398787 536255 398790
rect 547830 398306 547890 398752
rect 549253 398306 549319 398309
rect 547830 398304 549319 398306
rect 547830 398248 549258 398304
rect 549314 398248 549319 398304
rect 547830 398246 549319 398248
rect 549253 398243 549319 398246
rect 498837 398034 498903 398037
rect 498837 398032 538138 398034
rect 498837 397976 498842 398032
rect 498898 397976 538138 398032
rect 498837 397974 538138 397976
rect 498837 397971 498903 397974
rect 538078 397936 538138 397974
rect -960 397340 480 397580
rect 493409 396810 493475 396813
rect 536281 396810 536347 396813
rect 493409 396808 536347 396810
rect 493409 396752 493414 396808
rect 493470 396752 536286 396808
rect 536342 396752 536347 396808
rect 493409 396750 536347 396752
rect 493409 396747 493475 396750
rect 536281 396747 536347 396750
rect 536097 396130 536163 396133
rect 538078 396130 538138 396576
rect 536097 396128 538138 396130
rect 536097 396072 536102 396128
rect 536158 396072 538138 396128
rect 536097 396070 538138 396072
rect 536097 396067 536163 396070
rect 536741 395994 536807 395997
rect 536741 395992 538138 395994
rect 536741 395936 536746 395992
rect 536802 395936 538138 395992
rect 536741 395934 538138 395936
rect 536741 395931 536807 395934
rect 485221 393954 485287 393957
rect 496077 393954 496143 393957
rect 485221 393952 496143 393954
rect 485221 393896 485226 393952
rect 485282 393896 496082 393952
rect 496138 393896 496143 393952
rect 485221 393894 496143 393896
rect 485221 393891 485287 393894
rect 496077 393891 496143 393894
rect 470133 392594 470199 392597
rect 471513 392594 471579 392597
rect 470133 392592 471579 392594
rect 470133 392536 470138 392592
rect 470194 392536 471518 392592
rect 471574 392536 471579 392592
rect 470133 392534 471579 392536
rect 470133 392531 470199 392534
rect 471513 392531 471579 392534
rect 481817 392594 481883 392597
rect 494697 392594 494763 392597
rect 481817 392592 494763 392594
rect 481817 392536 481822 392592
rect 481878 392536 494702 392592
rect 494758 392536 494763 392592
rect 481817 392534 494763 392536
rect 481817 392531 481883 392534
rect 494697 392531 494763 392534
rect 482553 392186 482619 392189
rect 488533 392186 488599 392189
rect 490741 392186 490807 392189
rect 482553 392184 490807 392186
rect 482553 392128 482558 392184
rect 482614 392128 488538 392184
rect 488594 392128 490746 392184
rect 490802 392128 490807 392184
rect 482553 392126 490807 392128
rect 482553 392123 482619 392126
rect 488533 392123 488599 392126
rect 490741 392123 490807 392126
rect 471513 392050 471579 392053
rect 477861 392050 477927 392053
rect 471513 392048 477927 392050
rect 471513 391992 471518 392048
rect 471574 391992 477866 392048
rect 477922 391992 477927 392048
rect 471513 391990 477927 391992
rect 471513 391987 471579 391990
rect 477861 391987 477927 391990
rect 488625 392050 488691 392053
rect 490833 392050 490899 392053
rect 488625 392048 490899 392050
rect 488625 391992 488630 392048
rect 488686 391992 490838 392048
rect 490894 391992 490899 392048
rect 488625 391990 490899 391992
rect 488625 391987 488691 391990
rect 490833 391987 490899 391990
rect 470266 391085 470822 391086
rect 470266 390781 470272 391085
rect 470816 390781 470822 391085
rect 477861 390962 477927 390965
rect 482553 390962 482619 390965
rect 477861 390960 477970 390962
rect 477861 390904 477866 390960
rect 477922 390904 477970 390960
rect 477861 390899 477970 390904
rect 470266 390780 470822 390781
rect 477910 390690 477970 390899
rect 482510 390960 482619 390962
rect 482510 390904 482558 390960
rect 482614 390904 482619 390960
rect 482510 390899 482619 390904
rect 489177 390962 489243 390965
rect 489177 390960 489378 390962
rect 489177 390904 489182 390960
rect 489238 390904 489378 390960
rect 489177 390902 489378 390904
rect 489177 390899 489243 390902
rect 478045 390690 478111 390693
rect 477910 390688 478111 390690
rect 477910 390632 478050 390688
rect 478106 390632 478111 390688
rect 477910 390630 478111 390632
rect 478045 390627 478111 390630
rect 482369 390690 482435 390693
rect 482510 390690 482570 390899
rect 482369 390688 482570 390690
rect 482369 390632 482374 390688
rect 482430 390632 482570 390688
rect 482369 390630 482570 390632
rect 489318 390690 489378 390902
rect 489453 390690 489519 390693
rect 489318 390688 489519 390690
rect 489318 390632 489458 390688
rect 489514 390632 489519 390688
rect 489318 390630 489519 390632
rect 482369 390627 482435 390630
rect 489453 390627 489519 390630
rect 469026 390002 469582 390003
rect 469026 389698 469032 390002
rect 469576 389698 469582 390002
rect 469026 389697 469582 389698
rect 470266 388912 470822 388913
rect 470266 388608 470272 388912
rect 470816 388608 470822 388912
rect 470266 388607 470822 388608
rect 490606 388106 490666 388620
rect 536741 388378 536807 388381
rect 538078 388378 538138 395934
rect 583520 391628 584960 391868
rect 536741 388376 538138 388378
rect 536741 388320 536746 388376
rect 536802 388320 538138 388376
rect 536741 388318 538138 388320
rect 536741 388315 536807 388318
rect 493685 388106 493751 388109
rect 490606 388104 493751 388106
rect 490606 388048 493690 388104
rect 493746 388048 493751 388104
rect 490606 388046 493751 388048
rect 493685 388043 493751 388046
rect 475745 387698 475811 387701
rect 545021 387698 545087 387701
rect 547873 387698 547939 387701
rect 475745 387696 476130 387698
rect 475745 387640 475750 387696
rect 475806 387640 476130 387696
rect 475745 387638 476130 387640
rect 475745 387635 475811 387638
rect 476070 387426 476130 387638
rect 545021 387696 547939 387698
rect 545021 387640 545026 387696
rect 545082 387640 547878 387696
rect 547934 387640 547939 387696
rect 545021 387638 547939 387640
rect 545021 387635 545087 387638
rect 547873 387635 547939 387638
rect 479609 387562 479675 387565
rect 494789 387562 494855 387565
rect 479609 387560 494855 387562
rect 479609 387504 479614 387560
rect 479670 387504 494794 387560
rect 494850 387504 494855 387560
rect 479609 387502 494855 387504
rect 479609 387499 479675 387502
rect 494789 387499 494855 387502
rect 492121 387426 492187 387429
rect 476070 387424 492187 387426
rect 476070 387368 492126 387424
rect 492182 387368 492187 387424
rect 476070 387366 492187 387368
rect 492121 387363 492187 387366
rect 538121 387018 538187 387021
rect 540973 387018 541039 387021
rect 538121 387016 541039 387018
rect 538121 386960 538126 387016
rect 538182 386960 540978 387016
rect 541034 386960 541039 387016
rect 538121 386958 541039 386960
rect 538121 386955 538187 386958
rect 540973 386955 541039 386958
rect 483197 386474 483263 386477
rect 489545 386474 489611 386477
rect 483197 386472 489611 386474
rect 483197 386416 483202 386472
rect 483258 386416 489550 386472
rect 489606 386416 489611 386472
rect 483197 386414 489611 386416
rect 483197 386411 483263 386414
rect 489545 386411 489611 386414
rect -960 384284 480 384524
rect 485681 382394 485747 382397
rect 490833 382394 490899 382397
rect 485681 382392 490899 382394
rect 485681 382336 485686 382392
rect 485742 382336 490838 382392
rect 490894 382336 490899 382392
rect 485681 382334 490899 382336
rect 485681 382331 485747 382334
rect 490833 382331 490899 382334
rect 583520 378300 584960 378540
rect 538121 375458 538187 375461
rect 540973 375458 541039 375461
rect 538121 375456 541039 375458
rect 538121 375400 538126 375456
rect 538182 375400 540978 375456
rect 541034 375400 541039 375456
rect 538121 375398 541039 375400
rect 538121 375395 538187 375398
rect 540973 375395 541039 375398
rect 501597 372874 501663 372877
rect 501597 372872 538108 372874
rect 501597 372816 501602 372872
rect 501658 372816 538108 372872
rect 501597 372814 538108 372816
rect 501597 372811 501663 372814
rect 486877 372058 486943 372061
rect 490649 372058 490715 372061
rect 486877 372056 490715 372058
rect 486877 372000 486882 372056
rect 486938 372000 490654 372056
rect 490710 372000 490715 372056
rect 486877 371998 490715 372000
rect 486877 371995 486943 371998
rect 490649 371995 490715 371998
rect 482369 371922 482435 371925
rect 490741 371922 490807 371925
rect 482369 371920 490807 371922
rect 482369 371864 482374 371920
rect 482430 371864 490746 371920
rect 490802 371864 490807 371920
rect 482369 371862 490807 371864
rect 482369 371859 482435 371862
rect 490741 371859 490807 371862
rect 496261 371514 496327 371517
rect 496261 371512 538108 371514
rect -960 371228 480 371468
rect 496261 371456 496266 371512
rect 496322 371456 538108 371512
rect 496261 371454 538108 371456
rect 496261 371451 496327 371454
rect 471605 371378 471671 371381
rect 473721 371378 473787 371381
rect 471605 371376 473787 371378
rect 471605 371320 471610 371376
rect 471666 371320 473726 371376
rect 473782 371320 473787 371376
rect 471605 371318 473787 371320
rect 471605 371315 471671 371318
rect 473721 371315 473787 371318
rect 470133 370290 470199 370293
rect 473261 370290 473327 370293
rect 470133 370288 478890 370290
rect 470133 370232 470138 370288
rect 470194 370232 473266 370288
rect 473322 370232 478890 370288
rect 470133 370230 478890 370232
rect 470133 370227 470199 370230
rect 473261 370227 473327 370230
rect 470266 370085 470822 370086
rect 470266 369781 470272 370085
rect 470816 369781 470822 370085
rect 470266 369780 470822 369781
rect 478830 369613 478890 370230
rect 494697 370154 494763 370157
rect 494697 370152 538108 370154
rect 494697 370096 494702 370152
rect 494758 370096 538108 370152
rect 494697 370094 538108 370096
rect 494697 370091 494763 370094
rect 482369 369882 482435 369885
rect 485681 369882 485747 369885
rect 482326 369880 482435 369882
rect 482326 369824 482374 369880
rect 482430 369824 482435 369880
rect 482326 369819 482435 369824
rect 485454 369880 485747 369882
rect 485454 369824 485686 369880
rect 485742 369824 485747 369880
rect 485454 369822 485747 369824
rect 482326 369746 482386 369819
rect 481958 369686 482386 369746
rect 478830 369608 478939 369613
rect 478830 369552 478878 369608
rect 478934 369552 478939 369608
rect 478830 369550 478939 369552
rect 478873 369547 478939 369550
rect 481817 369610 481883 369613
rect 481958 369610 482018 369686
rect 481817 369608 482018 369610
rect 481817 369552 481822 369608
rect 481878 369552 482018 369608
rect 481817 369550 482018 369552
rect 485313 369610 485379 369613
rect 485454 369610 485514 369822
rect 485681 369819 485747 369822
rect 485313 369608 485514 369610
rect 485313 369552 485318 369608
rect 485374 369552 485514 369608
rect 485313 369550 485514 369552
rect 481817 369547 481883 369550
rect 485313 369547 485379 369550
rect 469026 368999 469582 369000
rect 469026 368695 469032 368999
rect 469576 368695 469582 368999
rect 489545 368794 489611 368797
rect 489545 368792 538108 368794
rect 489545 368736 489550 368792
rect 489606 368736 538108 368792
rect 489545 368734 538108 368736
rect 489545 368731 489611 368734
rect 469026 368694 469582 368695
rect 489453 368114 489519 368117
rect 492121 368114 492187 368117
rect 489453 368112 492187 368114
rect 489453 368056 489458 368112
rect 489514 368056 492126 368112
rect 492182 368056 492187 368112
rect 489453 368054 492187 368056
rect 489453 368051 489519 368054
rect 492121 368051 492187 368054
rect 470266 367912 470822 367913
rect 470266 367608 470272 367912
rect 470816 367608 470822 367912
rect 470266 367607 470822 367608
rect 489361 367298 489427 367301
rect 536373 367298 536439 367301
rect 489361 367296 536439 367298
rect 489361 367240 489366 367296
rect 489422 367240 536378 367296
rect 536434 367240 536439 367296
rect 489361 367238 536439 367240
rect 489361 367235 489427 367238
rect 536373 367235 536439 367238
rect 538078 367162 538138 367404
rect 536790 367102 538138 367162
rect 477217 367026 477283 367029
rect 492213 367026 492279 367029
rect 536790 367026 536850 367102
rect 477217 367024 492279 367026
rect 477217 366968 477222 367024
rect 477278 366968 492218 367024
rect 492274 366968 492279 367024
rect 477217 366966 492279 366968
rect 477217 366963 477283 366966
rect 492213 366963 492279 366966
rect 528510 366966 536850 367026
rect 480161 366890 480227 366893
rect 497549 366890 497615 366893
rect 480161 366888 497615 366890
rect 480161 366832 480166 366888
rect 480222 366832 497554 366888
rect 497610 366832 497615 366888
rect 480161 366830 497615 366832
rect 480161 366827 480227 366830
rect 497549 366827 497615 366830
rect 483197 366754 483263 366757
rect 528510 366754 528570 366966
rect 483197 366752 528570 366754
rect 483197 366696 483202 366752
rect 483258 366696 528570 366752
rect 483197 366694 528570 366696
rect 483197 366691 483263 366694
rect 535453 366074 535519 366077
rect 535453 366072 538108 366074
rect 535453 366016 535458 366072
rect 535514 366016 538108 366072
rect 535453 366014 538108 366016
rect 535453 366011 535519 366014
rect 490741 364986 490807 364989
rect 535453 364986 535519 364989
rect 490741 364984 535519 364986
rect 490741 364928 490746 364984
rect 490802 364928 535458 364984
rect 535514 364928 535519 364984
rect 583520 364972 584960 365212
rect 490741 364926 535519 364928
rect 490741 364923 490807 364926
rect 535453 364923 535519 364926
rect 536373 364714 536439 364717
rect 536373 364712 538108 364714
rect 536373 364656 536378 364712
rect 536434 364656 538108 364712
rect 536373 364654 538108 364656
rect 536373 364651 536439 364654
rect 536281 363354 536347 363357
rect 536281 363352 538108 363354
rect 536281 363296 536286 363352
rect 536342 363296 538108 363352
rect 536281 363294 538108 363296
rect 536281 363291 536347 363294
rect 549253 362810 549319 362813
rect 547860 362808 549319 362810
rect 547860 362752 549258 362808
rect 549314 362752 549319 362808
rect 547860 362750 549319 362752
rect 549253 362747 549319 362750
rect 494697 361994 494763 361997
rect 494697 361992 538108 361994
rect 494697 361936 494702 361992
rect 494758 361936 538108 361992
rect 494697 361934 538108 361936
rect 494697 361931 494763 361934
rect 497549 360634 497615 360637
rect 497549 360632 538108 360634
rect 497549 360576 497554 360632
rect 497610 360576 538108 360632
rect 497549 360574 538108 360576
rect 497549 360571 497615 360574
rect 473261 359546 473327 359549
rect 476113 359546 476179 359549
rect 473261 359544 476179 359546
rect 473261 359488 473266 359544
rect 473322 359488 476118 359544
rect 476174 359488 476179 359544
rect 473261 359486 476179 359488
rect 473261 359483 473327 359486
rect 476113 359483 476179 359486
rect 536741 359274 536807 359277
rect 536741 359272 538108 359274
rect 536741 359216 536746 359272
rect 536802 359244 538108 359272
rect 536802 359216 538138 359244
rect 536741 359214 538138 359216
rect 536741 359211 536807 359214
rect -960 358308 480 358548
rect 536741 352474 536807 352477
rect 538078 352474 538138 359214
rect 536741 352472 538138 352474
rect 536741 352416 536746 352472
rect 536802 352444 538138 352472
rect 536802 352416 538108 352444
rect 536741 352414 538108 352416
rect 536741 352411 536807 352414
rect 548517 351930 548583 351933
rect 583520 351930 584960 352020
rect 548517 351928 584960 351930
rect 548517 351872 548522 351928
rect 548578 351872 584960 351928
rect 548517 351870 584960 351872
rect 548517 351867 548583 351870
rect 583520 351780 584960 351870
rect 538121 351114 538187 351117
rect 540973 351114 541039 351117
rect 538121 351112 541039 351114
rect 538121 351056 538126 351112
rect 538182 351056 540978 351112
rect 541034 351056 541039 351112
rect 538121 351054 541039 351056
rect 538121 351051 538187 351054
rect 540973 351051 541039 351054
rect 488809 350706 488875 350709
rect 489637 350706 489703 350709
rect 488809 350704 489703 350706
rect 488809 350648 488814 350704
rect 488870 350648 489642 350704
rect 489698 350648 489703 350704
rect 488809 350646 489703 350648
rect 488809 350643 488875 350646
rect 489637 350643 489703 350646
rect 473721 350570 473787 350573
rect 481265 350570 481331 350573
rect 488901 350570 488967 350573
rect 473721 350568 488967 350570
rect 473721 350512 473726 350568
rect 473782 350512 481270 350568
rect 481326 350512 488906 350568
rect 488962 350512 488967 350568
rect 473721 350510 488967 350512
rect 473721 350507 473787 350510
rect 481265 350507 481331 350510
rect 488901 350507 488967 350510
rect 486417 349754 486483 349757
rect 494789 349754 494855 349757
rect 486417 349752 494855 349754
rect 486417 349696 486422 349752
rect 486478 349696 494794 349752
rect 494850 349696 494855 349752
rect 486417 349694 494855 349696
rect 486417 349691 486483 349694
rect 494789 349691 494855 349694
rect 471697 349210 471763 349213
rect 473353 349210 473419 349213
rect 471697 349208 474290 349210
rect 471697 349152 471702 349208
rect 471758 349152 473358 349208
rect 473414 349152 474290 349208
rect 471697 349150 474290 349152
rect 471697 349147 471763 349150
rect 473353 349147 473419 349150
rect 470266 349084 470822 349085
rect 470266 348780 470272 349084
rect 470816 348780 470822 349084
rect 470266 348779 470822 348780
rect 474230 348397 474290 349150
rect 476113 348802 476179 348805
rect 481265 348802 481331 348805
rect 475702 348800 476179 348802
rect 475702 348744 476118 348800
rect 476174 348744 476179 348800
rect 475702 348742 476179 348744
rect 475702 348533 475762 348742
rect 476113 348739 476179 348742
rect 481222 348800 481331 348802
rect 481222 348744 481270 348800
rect 481326 348744 481331 348800
rect 481222 348739 481331 348744
rect 475653 348528 475762 348533
rect 475653 348472 475658 348528
rect 475714 348472 475762 348528
rect 475653 348470 475762 348472
rect 475653 348467 475719 348470
rect 474181 348392 474290 348397
rect 474181 348336 474186 348392
rect 474242 348336 474290 348392
rect 474181 348334 474290 348336
rect 481222 348397 481282 348739
rect 481222 348392 481293 348397
rect 481222 348336 481232 348392
rect 481288 348336 481293 348392
rect 481222 348334 481293 348336
rect 474181 348331 474247 348334
rect 481227 348331 481293 348334
rect 469026 347997 469582 347998
rect 469026 347693 469032 347997
rect 469576 347693 469582 347997
rect 469026 347692 469582 347693
rect 488993 347034 489059 347037
rect 492213 347034 492279 347037
rect 488993 347032 492279 347034
rect 488993 346976 488998 347032
rect 489054 346976 492218 347032
rect 492274 346976 492279 347032
rect 488993 346974 492279 346976
rect 488993 346971 489059 346974
rect 492213 346971 492279 346974
rect 470266 346912 470822 346913
rect 470266 346608 470272 346912
rect 470816 346608 470822 346912
rect 470266 346607 470822 346608
rect 475561 346354 475627 346357
rect 492029 346354 492095 346357
rect 475561 346352 492095 346354
rect 475561 346296 475566 346352
rect 475622 346296 492034 346352
rect 492090 346296 492095 346352
rect 475561 346294 492095 346296
rect 475561 346291 475627 346294
rect 492029 346291 492095 346294
rect -960 345252 480 345492
rect 478597 344994 478663 344997
rect 496169 344994 496235 344997
rect 478597 344992 496235 344994
rect 478597 344936 478602 344992
rect 478658 344936 496174 344992
rect 496230 344936 496235 344992
rect 478597 344934 496235 344936
rect 478597 344931 478663 344934
rect 496169 344931 496235 344934
rect 482185 344858 482251 344861
rect 490741 344858 490807 344861
rect 482185 344856 490807 344858
rect 482185 344800 482190 344856
rect 482246 344800 490746 344856
rect 490802 344800 490807 344856
rect 482185 344798 490807 344800
rect 482185 344795 482251 344798
rect 490741 344795 490807 344798
rect 499113 344314 499179 344317
rect 536373 344314 536439 344317
rect 499113 344312 536439 344314
rect 499113 344256 499118 344312
rect 499174 344256 536378 344312
rect 536434 344256 536439 344312
rect 499113 344254 536439 344256
rect 499113 344251 499179 344254
rect 536373 344251 536439 344254
rect 471697 342274 471763 342277
rect 474641 342274 474707 342277
rect 471697 342272 474707 342274
rect 471697 342216 471702 342272
rect 471758 342216 474646 342272
rect 474702 342216 474707 342272
rect 471697 342214 474707 342216
rect 471697 342211 471763 342214
rect 474641 342211 474707 342214
rect 538121 339554 538187 339557
rect 541249 339554 541315 339557
rect 538121 339552 541315 339554
rect 538121 339496 538126 339552
rect 538182 339496 541254 339552
rect 541310 339496 541315 339552
rect 538121 339494 541315 339496
rect 538121 339491 538187 339494
rect 541249 339491 541315 339494
rect 544193 339554 544259 339557
rect 547873 339554 547939 339557
rect 548517 339554 548583 339557
rect 544193 339552 548583 339554
rect 544193 339496 544198 339552
rect 544254 339496 547878 339552
rect 547934 339496 548522 339552
rect 548578 339496 548583 339552
rect 544193 339494 548583 339496
rect 544193 339491 544259 339494
rect 547873 339491 547939 339494
rect 548517 339491 548583 339494
rect 583520 338452 584960 338692
rect 499021 336834 499087 336837
rect 499021 336832 538108 336834
rect 499021 336776 499026 336832
rect 499082 336776 538108 336832
rect 499021 336774 538108 336776
rect 499021 336771 499087 336774
rect 500217 335474 500283 335477
rect 500217 335472 538108 335474
rect 500217 335416 500222 335472
rect 500278 335416 538108 335472
rect 500217 335414 538108 335416
rect 500217 335411 500283 335414
rect 496077 334114 496143 334117
rect 496077 334112 538108 334114
rect 496077 334056 496082 334112
rect 496138 334056 538108 334112
rect 496077 334054 538108 334056
rect 496077 334051 496143 334054
rect 490649 332754 490715 332757
rect 490649 332752 538108 332754
rect 490649 332696 490654 332752
rect 490710 332696 538108 332752
rect 490649 332694 538108 332696
rect 490649 332691 490715 332694
rect -960 332196 480 332436
rect 494789 331394 494855 331397
rect 494789 331392 538108 331394
rect 494789 331336 494794 331392
rect 494850 331336 538108 331392
rect 494789 331334 538108 331336
rect 494789 331331 494855 331334
rect 485405 330034 485471 330037
rect 485405 330032 538108 330034
rect 485405 329976 485410 330032
rect 485466 329976 538108 330032
rect 485405 329974 538108 329976
rect 485405 329971 485471 329974
rect 471605 329898 471671 329901
rect 481541 329898 481607 329901
rect 488901 329898 488967 329901
rect 471605 329896 488967 329898
rect 471605 329840 471610 329896
rect 471666 329840 481546 329896
rect 481602 329840 488906 329896
rect 488962 329840 488967 329896
rect 471605 329838 488967 329840
rect 471605 329835 471671 329838
rect 481541 329835 481607 329838
rect 488901 329835 488967 329838
rect 489913 328674 489979 328677
rect 489913 328672 538108 328674
rect 489913 328616 489918 328672
rect 489974 328616 538108 328672
rect 489913 328614 538108 328616
rect 489913 328611 489979 328614
rect 470266 328084 470822 328085
rect 470266 327780 470272 328084
rect 470816 327780 470822 328084
rect 474641 327858 474707 327861
rect 470266 327779 470822 327780
rect 474598 327856 474707 327858
rect 474598 327800 474646 327856
rect 474702 327800 474707 327856
rect 474598 327795 474707 327800
rect 481541 327858 481607 327861
rect 485405 327858 485471 327861
rect 481541 327856 481650 327858
rect 481541 327800 481546 327856
rect 481602 327800 481650 327856
rect 481541 327795 481650 327800
rect 471697 327722 471763 327725
rect 474598 327722 474658 327795
rect 471697 327720 474658 327722
rect 471697 327664 471702 327720
rect 471758 327664 474658 327720
rect 471697 327662 474658 327664
rect 471697 327659 471763 327662
rect 474598 327453 474658 327662
rect 481590 327453 481650 327795
rect 485270 327856 485471 327858
rect 485270 327800 485410 327856
rect 485466 327800 485471 327856
rect 485270 327798 485471 327800
rect 474598 327448 474714 327453
rect 474598 327392 474653 327448
rect 474709 327392 474714 327448
rect 474598 327390 474714 327392
rect 474648 327387 474714 327390
rect 481537 327448 481650 327453
rect 481537 327392 481542 327448
rect 481598 327392 481650 327448
rect 481537 327390 481650 327392
rect 484981 327450 485047 327453
rect 485270 327450 485330 327798
rect 485405 327795 485471 327798
rect 484981 327448 485330 327450
rect 484981 327392 484986 327448
rect 485042 327392 485330 327448
rect 484981 327390 485330 327392
rect 481537 327387 481603 327390
rect 484981 327387 485047 327390
rect 536373 327314 536439 327317
rect 536373 327312 538108 327314
rect 536373 327256 536378 327312
rect 536434 327256 538108 327312
rect 536373 327254 538108 327256
rect 536373 327251 536439 327254
rect 469026 326997 469582 326998
rect 469026 326693 469032 326997
rect 469576 326693 469582 326997
rect 471513 326906 471579 326909
rect 476205 326906 476271 326909
rect 489913 326906 489979 326909
rect 471513 326904 476271 326906
rect 471513 326848 471518 326904
rect 471574 326848 476210 326904
rect 476266 326848 476271 326904
rect 471513 326846 476271 326848
rect 471513 326843 471579 326846
rect 476205 326843 476271 326846
rect 485822 326904 489979 326906
rect 485822 326848 489918 326904
rect 489974 326848 489979 326904
rect 485822 326846 489979 326848
rect 469026 326692 469582 326693
rect 485822 326604 485882 326846
rect 489913 326843 489979 326846
rect 549253 326770 549319 326773
rect 547860 326768 549319 326770
rect 547860 326712 549258 326768
rect 549314 326712 549319 326768
rect 547860 326710 549319 326712
rect 549253 326707 549319 326710
rect 536189 325954 536255 325957
rect 536189 325952 538108 325954
rect 470266 325912 470822 325913
rect 470266 325608 470272 325912
rect 470816 325608 470822 325912
rect 536189 325896 536194 325952
rect 536250 325896 538108 325952
rect 536189 325894 538108 325896
rect 536189 325891 536255 325894
rect 470266 325607 470822 325608
rect 475469 325410 475535 325413
rect 493593 325410 493659 325413
rect 475469 325408 493659 325410
rect 475469 325352 475474 325408
rect 475530 325352 493598 325408
rect 493654 325352 493659 325408
rect 475469 325350 493659 325352
rect 475469 325347 475535 325350
rect 493593 325347 493659 325350
rect 583520 325124 584960 325364
rect 490741 325002 490807 325005
rect 536097 325002 536163 325005
rect 490741 325000 536163 325002
rect 490741 324944 490746 325000
rect 490802 324944 536102 325000
rect 536158 324944 536163 325000
rect 490741 324942 536163 324944
rect 490741 324939 490807 324942
rect 536097 324939 536163 324942
rect 536281 324594 536347 324597
rect 536281 324592 538108 324594
rect 536281 324536 536286 324592
rect 536342 324536 538108 324592
rect 536281 324534 538108 324536
rect 536281 324531 536347 324534
rect 479057 324186 479123 324189
rect 489637 324186 489703 324189
rect 479057 324184 489703 324186
rect 479057 324128 479062 324184
rect 479118 324128 489642 324184
rect 489698 324128 489703 324184
rect 479057 324126 489703 324128
rect 479057 324123 479123 324126
rect 489637 324123 489703 324126
rect 482369 324050 482435 324053
rect 499113 324050 499179 324053
rect 482369 324048 499179 324050
rect 482369 323992 482374 324048
rect 482430 323992 499118 324048
rect 499174 323992 499179 324048
rect 482369 323990 499179 323992
rect 482369 323987 482435 323990
rect 499113 323987 499179 323990
rect 536741 323234 536807 323237
rect 536741 323232 538108 323234
rect 536741 323176 536746 323232
rect 536802 323204 538108 323232
rect 536802 323176 538138 323204
rect 536741 323174 538138 323176
rect 536741 323171 536807 323174
rect -960 319140 480 319380
rect 536741 316434 536807 316437
rect 538078 316434 538138 323174
rect 536741 316432 538138 316434
rect 536741 316376 536746 316432
rect 536802 316404 538138 316432
rect 536802 316376 538108 316404
rect 536741 316374 538108 316376
rect 536741 316371 536807 316374
rect 538121 315346 538187 315349
rect 541709 315346 541775 315349
rect 538121 315344 541775 315346
rect 538121 315288 538126 315344
rect 538182 315288 541714 315344
rect 541770 315288 541775 315344
rect 538121 315286 541775 315288
rect 538121 315283 538187 315286
rect 541709 315283 541775 315286
rect 488625 313306 488691 313309
rect 489637 313306 489703 313309
rect 488625 313304 489703 313306
rect 488625 313248 488630 313304
rect 488686 313248 489642 313304
rect 489698 313248 489703 313304
rect 488625 313246 489703 313248
rect 488625 313243 488691 313246
rect 489637 313243 489703 313246
rect 583520 311932 584960 312172
rect 471605 308410 471671 308413
rect 480897 308410 480963 308413
rect 488533 308410 488599 308413
rect 471605 308408 488599 308410
rect 471605 308352 471610 308408
rect 471666 308352 480902 308408
rect 480958 308352 488538 308408
rect 488594 308352 488599 308408
rect 471605 308350 488599 308352
rect 471605 308347 471671 308350
rect 480897 308347 480963 308350
rect 488533 308347 488599 308350
rect 471513 307866 471579 307869
rect 477493 307866 477559 307869
rect 471513 307864 477559 307866
rect 471513 307808 471518 307864
rect 471574 307808 477498 307864
rect 477554 307808 477559 307864
rect 471513 307806 477559 307808
rect 471513 307803 471579 307806
rect 477493 307803 477559 307806
rect 470266 307084 470822 307085
rect 470266 306780 470272 307084
rect 470816 306780 470822 307084
rect 477493 306914 477559 306917
rect 480897 306914 480963 306917
rect 477493 306912 477602 306914
rect 477493 306856 477498 306912
rect 477554 306856 477602 306912
rect 477493 306851 477602 306856
rect 470266 306779 470822 306780
rect 477542 306645 477602 306851
rect 480854 306912 480963 306914
rect 480854 306856 480902 306912
rect 480958 306856 480963 306912
rect 480854 306851 480963 306856
rect 480854 306645 480914 306851
rect 488625 306778 488691 306781
rect 484350 306776 488691 306778
rect 484350 306720 488630 306776
rect 488686 306720 488691 306776
rect 484350 306718 488691 306720
rect 484350 306645 484410 306718
rect 488625 306715 488691 306718
rect 477542 306640 477651 306645
rect 477542 306584 477590 306640
rect 477646 306584 477651 306640
rect 477542 306582 477651 306584
rect 480854 306640 480963 306645
rect 480854 306584 480902 306640
rect 480958 306584 480963 306640
rect 480854 306582 480963 306584
rect 477585 306579 477651 306582
rect 480897 306579 480963 306582
rect 484301 306640 484410 306645
rect 484301 306584 484306 306640
rect 484362 306584 484410 306640
rect 484301 306582 484410 306584
rect 484301 306579 484367 306582
rect -960 306084 480 306324
rect 469026 305999 469582 306000
rect 469026 305695 469032 305999
rect 469576 305695 469582 305999
rect 469026 305694 469582 305695
rect 544193 305010 544259 305013
rect 547873 305010 547939 305013
rect 544193 305008 547939 305010
rect 544193 304952 544198 305008
rect 544254 304952 547878 305008
rect 547934 304952 547939 305008
rect 544193 304950 547939 304952
rect 544193 304947 544259 304950
rect 547873 304947 547939 304950
rect 470266 304912 470822 304913
rect 470266 304608 470272 304912
rect 470816 304608 470822 304912
rect 470266 304607 470822 304608
rect 541709 303786 541775 303789
rect 549161 303786 549227 303789
rect 541709 303784 549227 303786
rect 541709 303728 541714 303784
rect 541770 303728 549166 303784
rect 549222 303728 549227 303784
rect 541709 303726 549227 303728
rect 541709 303723 541775 303726
rect 549161 303723 549227 303726
rect 539225 303650 539291 303653
rect 548517 303650 548583 303653
rect 539225 303648 548583 303650
rect 539225 303592 539230 303648
rect 539286 303592 548522 303648
rect 548578 303592 548583 303648
rect 539225 303590 548583 303592
rect 539225 303587 539291 303590
rect 548517 303587 548583 303590
rect 493685 301474 493751 301477
rect 536097 301474 536163 301477
rect 493685 301472 536163 301474
rect 493685 301416 493690 301472
rect 493746 301416 536102 301472
rect 536158 301416 536163 301472
rect 493685 301414 536163 301416
rect 493685 301411 493751 301414
rect 536097 301411 536163 301414
rect 497457 300794 497523 300797
rect 497457 300792 538108 300794
rect 497457 300736 497462 300792
rect 497518 300736 538108 300792
rect 497457 300734 538108 300736
rect 497457 300731 497523 300734
rect 491937 299434 492003 299437
rect 491937 299432 538108 299434
rect 491937 299376 491942 299432
rect 491998 299376 538108 299432
rect 491937 299374 538108 299376
rect 491937 299371 492003 299374
rect 549161 298754 549227 298757
rect 583520 298754 584960 298844
rect 549161 298752 584960 298754
rect 549161 298696 549166 298752
rect 549222 298696 584960 298752
rect 549161 298694 584960 298696
rect 549161 298691 549227 298694
rect 583520 298604 584960 298694
rect 498929 298074 498995 298077
rect 498929 298072 538108 298074
rect 498929 298016 498934 298072
rect 498990 298016 538108 298072
rect 498929 298014 538108 298016
rect 498929 298011 498995 298014
rect 536097 296714 536163 296717
rect 536097 296712 538108 296714
rect 536097 296656 536102 296712
rect 536158 296656 538108 296712
rect 536097 296654 538108 296656
rect 536097 296651 536163 296654
rect 492121 295490 492187 295493
rect 492121 295488 538138 295490
rect 492121 295432 492126 295488
rect 492182 295432 538138 295488
rect 492121 295430 538138 295432
rect 492121 295427 492187 295430
rect 538078 295324 538138 295430
rect 492213 294130 492279 294133
rect 492213 294128 538138 294130
rect 492213 294072 492218 294128
rect 492274 294072 538138 294128
rect 492213 294070 538138 294072
rect 492213 294067 492279 294070
rect 538078 293964 538138 294070
rect -960 293028 480 293268
rect 492029 292770 492095 292773
rect 492029 292768 538138 292770
rect 492029 292712 492034 292768
rect 492090 292712 538138 292768
rect 492029 292710 538138 292712
rect 492029 292707 492095 292710
rect 538078 292604 538138 292710
rect 535453 291274 535519 291277
rect 535453 291272 538108 291274
rect 535453 291216 535458 291272
rect 535514 291216 538108 291272
rect 535453 291214 538108 291216
rect 535453 291211 535519 291214
rect 549253 290730 549319 290733
rect 549897 290730 549963 290733
rect 547860 290728 549963 290730
rect 547860 290672 549258 290728
rect 549314 290672 549902 290728
rect 549958 290672 549963 290728
rect 547860 290670 549963 290672
rect 549253 290667 549319 290670
rect 549897 290667 549963 290670
rect 493501 290050 493567 290053
rect 493501 290048 538138 290050
rect 493501 289992 493506 290048
rect 493562 289992 538138 290048
rect 493501 289990 538138 289992
rect 493501 289987 493567 289990
rect 538078 289884 538138 289990
rect 536097 288554 536163 288557
rect 536097 288552 538108 288554
rect 536097 288496 536102 288552
rect 536158 288496 538108 288552
rect 536097 288494 538108 288496
rect 536097 288491 536163 288494
rect 491293 287738 491359 287741
rect 536189 287738 536255 287741
rect 491293 287736 536255 287738
rect 491293 287680 491298 287736
rect 491354 287680 536194 287736
rect 536250 287680 536255 287736
rect 491293 287678 536255 287680
rect 491293 287675 491359 287678
rect 536189 287675 536255 287678
rect 482553 287466 482619 287469
rect 488533 287466 488599 287469
rect 490833 287466 490899 287469
rect 482553 287464 490899 287466
rect 482553 287408 482558 287464
rect 482614 287408 488538 287464
rect 488594 287408 490838 287464
rect 490894 287408 490899 287464
rect 482553 287406 490899 287408
rect 482553 287403 482619 287406
rect 488533 287403 488599 287406
rect 490833 287403 490899 287406
rect 471513 287330 471579 287333
rect 477861 287330 477927 287333
rect 471513 287328 477927 287330
rect 471513 287272 471518 287328
rect 471574 287272 477866 287328
rect 477922 287272 477927 287328
rect 471513 287270 477927 287272
rect 471513 287267 471579 287270
rect 477861 287267 477927 287270
rect 488625 287330 488691 287333
rect 491385 287330 491451 287333
rect 488625 287328 491451 287330
rect 488625 287272 488630 287328
rect 488686 287272 491390 287328
rect 491446 287272 491451 287328
rect 488625 287270 491451 287272
rect 488625 287267 488691 287270
rect 491385 287267 491451 287270
rect 471605 287194 471671 287197
rect 474733 287194 474799 287197
rect 471605 287192 474799 287194
rect 471605 287136 471610 287192
rect 471666 287136 474738 287192
rect 474794 287136 474799 287192
rect 471605 287134 474799 287136
rect 471605 287131 471671 287134
rect 474733 287131 474799 287134
rect 489269 287194 489335 287197
rect 494053 287194 494119 287197
rect 489269 287192 494119 287194
rect 489269 287136 489274 287192
rect 489330 287136 494058 287192
rect 494114 287136 494119 287192
rect 489269 287134 494119 287136
rect 489269 287131 489335 287134
rect 494053 287131 494119 287134
rect 536741 287194 536807 287197
rect 536741 287192 538108 287194
rect 536741 287136 536746 287192
rect 536802 287164 538108 287192
rect 536802 287136 538138 287164
rect 536741 287134 538138 287136
rect 536741 287131 536807 287134
rect 470266 286085 470822 286086
rect 470266 285781 470272 286085
rect 470816 285781 470822 286085
rect 474733 285968 474799 285973
rect 474733 285912 474738 285968
rect 474794 285912 474799 285968
rect 474733 285907 474799 285912
rect 477861 285968 477927 285973
rect 477861 285912 477866 285968
rect 477922 285912 477927 285968
rect 477861 285907 477927 285912
rect 482553 285968 482619 285973
rect 482553 285912 482558 285968
rect 482614 285912 482619 285968
rect 482553 285907 482619 285912
rect 489269 285968 489335 285973
rect 489269 285912 489274 285968
rect 489330 285912 489335 285968
rect 489269 285907 489335 285912
rect 470266 285780 470822 285781
rect 474736 285701 474796 285907
rect 474733 285696 474799 285701
rect 474733 285640 474738 285696
rect 474794 285640 474799 285696
rect 474733 285635 474799 285640
rect 477864 285698 477924 285907
rect 478045 285698 478111 285701
rect 477864 285696 478111 285698
rect 477864 285640 478050 285696
rect 478106 285640 478111 285696
rect 477864 285638 478111 285640
rect 478045 285635 478111 285638
rect 482369 285698 482435 285701
rect 482556 285698 482616 285907
rect 489272 285701 489332 285907
rect 482369 285696 482616 285698
rect 482369 285640 482374 285696
rect 482430 285640 482616 285696
rect 482369 285638 482616 285640
rect 489269 285696 489335 285701
rect 489269 285640 489274 285696
rect 489330 285640 489335 285696
rect 482369 285635 482435 285638
rect 489269 285635 489335 285640
rect 469026 285000 469582 285001
rect 469026 284696 469032 285000
rect 469576 284696 469582 285000
rect 469026 284695 469582 284696
rect 493501 284202 493567 284205
rect 490636 284200 493567 284202
rect 490636 284144 493506 284200
rect 493562 284144 493567 284200
rect 490636 284142 493567 284144
rect 493501 284139 493567 284142
rect 470266 283912 470822 283913
rect 470266 283608 470272 283912
rect 470816 283608 470822 283912
rect 470266 283607 470822 283608
rect 486877 282842 486943 282845
rect 491293 282842 491359 282845
rect 486877 282840 491359 282842
rect 486877 282784 486882 282840
rect 486938 282784 491298 282840
rect 491354 282784 491359 282840
rect 486877 282782 491359 282784
rect 486877 282779 486943 282782
rect 491293 282779 491359 282782
rect 475745 282706 475811 282709
rect 493317 282706 493383 282709
rect 475745 282704 493383 282706
rect 475745 282648 475750 282704
rect 475806 282648 493322 282704
rect 493378 282648 493383 282704
rect 475745 282646 493383 282648
rect 475745 282643 475811 282646
rect 493317 282643 493383 282646
rect 483197 282570 483263 282573
rect 494697 282570 494763 282573
rect 483197 282568 494763 282570
rect 483197 282512 483202 282568
rect 483258 282512 494702 282568
rect 494758 282512 494763 282568
rect 483197 282510 494763 282512
rect 483197 282507 483263 282510
rect 494697 282507 494763 282510
rect 479609 282434 479675 282437
rect 498837 282434 498903 282437
rect 479609 282432 498903 282434
rect 479609 282376 479614 282432
rect 479670 282376 498842 282432
rect 498898 282376 498903 282432
rect 479609 282374 498903 282376
rect 479609 282371 479675 282374
rect 498837 282371 498903 282374
rect 536741 280394 536807 280397
rect 538078 280394 538138 287134
rect 583520 285276 584960 285516
rect 548517 282162 548583 282165
rect 580349 282162 580415 282165
rect 548517 282160 580415 282162
rect 548517 282104 548522 282160
rect 548578 282104 580354 282160
rect 580410 282104 580415 282160
rect 548517 282102 580415 282104
rect 548517 282099 548583 282102
rect 580349 282099 580415 282102
rect 536741 280392 538138 280394
rect 536741 280336 536746 280392
rect 536802 280364 538138 280392
rect 536802 280336 538108 280364
rect 536741 280334 538108 280336
rect 536741 280331 536807 280334
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 476113 266930 476179 266933
rect 490557 266930 490623 266933
rect 476113 266928 490623 266930
rect 476113 266872 476118 266928
rect 476174 266872 490562 266928
rect 490618 266872 490623 266928
rect 476113 266870 490623 266872
rect 476113 266867 476179 266870
rect 490557 266867 490623 266870
rect 471513 266794 471579 266797
rect 479057 266794 479123 266797
rect 504357 266794 504423 266797
rect 471513 266792 504423 266794
rect 471513 266736 471518 266792
rect 471574 266736 479062 266792
rect 479118 266736 504362 266792
rect 504418 266736 504423 266792
rect 471513 266734 504423 266736
rect 471513 266731 471579 266734
rect 479057 266731 479123 266734
rect 504357 266731 504423 266734
rect 482553 266658 482619 266661
rect 489821 266658 489887 266661
rect 490833 266658 490899 266661
rect 482553 266656 490899 266658
rect 482553 266600 482558 266656
rect 482614 266600 489826 266656
rect 489882 266600 490838 266656
rect 490894 266600 490899 266656
rect 482553 266598 490899 266600
rect 482553 266595 482619 266598
rect 489821 266595 489887 266598
rect 490833 266595 490899 266598
rect 488441 266522 488507 266525
rect 494053 266522 494119 266525
rect 488441 266520 494119 266522
rect 488441 266464 488446 266520
rect 488502 266464 494058 266520
rect 494114 266464 494119 266520
rect 488441 266462 494119 266464
rect 488441 266459 488507 266462
rect 494053 266459 494119 266462
rect 471605 266386 471671 266389
rect 476113 266386 476179 266389
rect 471605 266384 476179 266386
rect 471605 266328 471610 266384
rect 471666 266328 476118 266384
rect 476174 266328 476179 266384
rect 471605 266326 476179 266328
rect 471605 266323 471671 266326
rect 476113 266323 476179 266326
rect 485313 266386 485379 266389
rect 491937 266386 492003 266389
rect 485313 266384 492003 266386
rect 485313 266328 485318 266384
rect 485374 266328 491942 266384
rect 491998 266328 492003 266384
rect 485313 266326 492003 266328
rect 485313 266323 485379 266326
rect 491937 266323 492003 266326
rect 491201 265570 491267 265573
rect 536281 265570 536347 265573
rect 491201 265568 536347 265570
rect 491201 265512 491206 265568
rect 491262 265512 536286 265568
rect 536342 265512 536347 265568
rect 491201 265510 536347 265512
rect 491201 265507 491267 265510
rect 536281 265507 536347 265510
rect 470266 265085 470822 265086
rect 470266 264781 470272 265085
rect 470816 264781 470822 265085
rect 476113 264890 476179 264893
rect 479057 264890 479123 264893
rect 482553 264890 482619 264893
rect 485313 264890 485379 264893
rect 488441 264890 488507 264893
rect 470266 264780 470822 264781
rect 476070 264888 476179 264890
rect 476070 264832 476118 264888
rect 476174 264832 476179 264888
rect 476070 264827 476179 264832
rect 479014 264888 479123 264890
rect 479014 264832 479062 264888
rect 479118 264832 479123 264888
rect 479014 264827 479123 264832
rect 482510 264888 482619 264890
rect 482510 264832 482558 264888
rect 482614 264832 482619 264888
rect 482510 264827 482619 264832
rect 485270 264888 485379 264890
rect 485270 264832 485318 264888
rect 485374 264832 485379 264888
rect 485270 264827 485379 264832
rect 488398 264888 488507 264890
rect 488398 264832 488446 264888
rect 488502 264832 488507 264888
rect 488398 264827 488507 264832
rect 476070 264621 476130 264827
rect 479014 264621 479074 264827
rect 476070 264616 476179 264621
rect 476070 264560 476118 264616
rect 476174 264560 476179 264616
rect 476070 264558 476179 264560
rect 479014 264616 479123 264621
rect 479014 264560 479062 264616
rect 479118 264560 479123 264616
rect 479014 264558 479123 264560
rect 476113 264555 476179 264558
rect 479057 264555 479123 264558
rect 482369 264618 482435 264621
rect 482510 264618 482570 264827
rect 482369 264616 482570 264618
rect 482369 264560 482374 264616
rect 482430 264560 482570 264616
rect 482369 264558 482570 264560
rect 485270 264618 485330 264827
rect 488398 264621 488458 264827
rect 485405 264618 485471 264621
rect 485270 264616 485471 264618
rect 485270 264560 485410 264616
rect 485466 264560 485471 264616
rect 485270 264558 485471 264560
rect 488398 264616 488507 264621
rect 488398 264560 488446 264616
rect 488502 264560 488507 264616
rect 488398 264558 488507 264560
rect 482369 264555 482435 264558
rect 485405 264555 485471 264558
rect 488441 264555 488507 264558
rect 494053 264210 494119 264213
rect 580257 264210 580323 264213
rect 494053 264208 580323 264210
rect 494053 264152 494058 264208
rect 494114 264152 580262 264208
rect 580318 264152 580323 264208
rect 494053 264150 580323 264152
rect 494053 264147 494119 264150
rect 580257 264147 580323 264150
rect 469026 263999 469582 264000
rect 469026 263695 469032 263999
rect 469576 263695 469582 263999
rect 469026 263694 469582 263695
rect 489453 263530 489519 263533
rect 536097 263530 536163 263533
rect 489453 263528 536163 263530
rect 489453 263472 489458 263528
rect 489514 263472 536102 263528
rect 536158 263472 536163 263528
rect 489453 263470 536163 263472
rect 489453 263467 489519 263470
rect 536097 263467 536163 263470
rect 470266 262912 470822 262913
rect 470266 262608 470272 262912
rect 470816 262608 470822 262912
rect 470266 262607 470822 262608
rect 486233 262170 486299 262173
rect 491201 262170 491267 262173
rect 486233 262168 491267 262170
rect 486233 262112 486238 262168
rect 486294 262112 491206 262168
rect 491262 262112 491267 262168
rect 486233 262110 491267 262112
rect 486233 262107 486299 262110
rect 491201 262107 491267 262110
rect 483197 262034 483263 262037
rect 497549 262034 497615 262037
rect 483197 262032 497615 262034
rect 483197 261976 483202 262032
rect 483258 261976 497554 262032
rect 497610 261976 497615 262032
rect 483197 261974 497615 261976
rect 483197 261971 483263 261974
rect 497549 261971 497615 261974
rect 480161 261898 480227 261901
rect 490741 261898 490807 261901
rect 480161 261896 490807 261898
rect 480161 261840 480166 261896
rect 480222 261840 490746 261896
rect 490802 261840 490807 261896
rect 480161 261838 490807 261840
rect 480161 261835 480227 261838
rect 490741 261835 490807 261838
rect 477217 261762 477283 261765
rect 493409 261762 493475 261765
rect 477217 261760 493475 261762
rect 477217 261704 477222 261760
rect 477278 261704 493414 261760
rect 493470 261704 493475 261760
rect 477217 261702 493475 261704
rect 477217 261699 477283 261702
rect 493409 261699 493475 261702
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 580349 245578 580415 245581
rect 583520 245578 584960 245668
rect 580349 245576 584960 245578
rect 580349 245520 580354 245576
rect 580410 245520 584960 245576
rect 580349 245518 584960 245520
rect 580349 245515 580415 245518
rect 583520 245428 584960 245518
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 580257 165882 580323 165885
rect 583520 165882 584960 165972
rect 580257 165880 584960 165882
rect 580257 165824 580262 165880
rect 580318 165824 584960 165880
rect 580257 165822 584960 165824
rect 580257 165819 580323 165822
rect 583520 165732 584960 165822
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 491937 126034 492003 126037
rect 583520 126034 584960 126124
rect 491937 126032 584960 126034
rect 491937 125976 491942 126032
rect 491998 125976 584960 126032
rect 491937 125974 584960 125976
rect 491937 125971 492003 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 489821 86186 489887 86189
rect 583520 86186 584960 86276
rect 489821 86184 584960 86186
rect 489821 86128 489826 86184
rect 489882 86128 584960 86184
rect 489821 86126 584960 86128
rect 489821 86123 489887 86126
rect 583520 86036 584960 86126
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 504357 46338 504423 46341
rect 583520 46338 584960 46428
rect 504357 46336 584960 46338
rect 504357 46280 504362 46336
rect 504418 46280 584960 46336
rect 504357 46278 584960 46280
rect 504357 46275 504423 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 549897 19818 549963 19821
rect 583520 19818 584960 19908
rect 549897 19816 584960 19818
rect 549897 19760 549902 19816
rect 549958 19760 584960 19816
rect 549897 19758 584960 19760
rect 549897 19755 549963 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect 490557 6626 490623 6629
rect 583520 6626 584960 6716
rect 490557 6624 584960 6626
rect -960 6340 480 6580
rect 490557 6568 490562 6624
rect 490618 6568 584960 6624
rect 490557 6566 584960 6568
rect 490557 6563 490623 6566
rect 583520 6476 584960 6566
<< via3 >>
rect 470272 451479 470816 451483
rect 470272 451183 470276 451479
rect 470276 451183 470812 451479
rect 470812 451183 470816 451479
rect 470272 451179 470816 451183
rect 469032 450393 469576 450397
rect 469032 450097 469036 450393
rect 469036 450097 469572 450393
rect 469572 450097 469576 450393
rect 469032 450093 469576 450097
rect 470272 449308 470816 449312
rect 470272 449012 470276 449308
rect 470276 449012 470812 449308
rect 470812 449012 470816 449308
rect 470272 449008 470816 449012
rect 470272 433080 470816 433084
rect 470272 432784 470276 433080
rect 470276 432784 470812 433080
rect 470812 432784 470816 433080
rect 470272 432780 470816 432784
rect 469032 431993 469576 431997
rect 469032 431697 469036 431993
rect 469036 431697 469572 431993
rect 469572 431697 469576 431993
rect 469032 431693 469576 431697
rect 470272 430908 470816 430912
rect 470272 430612 470276 430908
rect 470276 430612 470812 430908
rect 470812 430612 470816 430908
rect 470272 430608 470816 430612
rect 470272 412080 470816 412084
rect 470272 411784 470276 412080
rect 470276 411784 470812 412080
rect 470812 411784 470816 412080
rect 470272 411780 470816 411784
rect 469032 410994 469576 410998
rect 469032 410698 469036 410994
rect 469036 410698 469572 410994
rect 469572 410698 469576 410994
rect 469032 410694 469576 410698
rect 470272 409908 470816 409912
rect 470272 409612 470276 409908
rect 470276 409612 470812 409908
rect 470812 409612 470816 409908
rect 470272 409608 470816 409612
rect 470272 391081 470816 391085
rect 470272 390785 470276 391081
rect 470276 390785 470812 391081
rect 470812 390785 470816 391081
rect 470272 390781 470816 390785
rect 469032 389998 469576 390002
rect 469032 389702 469036 389998
rect 469036 389702 469572 389998
rect 469572 389702 469576 389998
rect 469032 389698 469576 389702
rect 470272 388908 470816 388912
rect 470272 388612 470276 388908
rect 470276 388612 470812 388908
rect 470812 388612 470816 388908
rect 470272 388608 470816 388612
rect 470272 370081 470816 370085
rect 470272 369785 470276 370081
rect 470276 369785 470812 370081
rect 470812 369785 470816 370081
rect 470272 369781 470816 369785
rect 469032 368995 469576 368999
rect 469032 368699 469036 368995
rect 469036 368699 469572 368995
rect 469572 368699 469576 368995
rect 469032 368695 469576 368699
rect 470272 367908 470816 367912
rect 470272 367612 470276 367908
rect 470276 367612 470812 367908
rect 470812 367612 470816 367908
rect 470272 367608 470816 367612
rect 470272 349080 470816 349084
rect 470272 348784 470276 349080
rect 470276 348784 470812 349080
rect 470812 348784 470816 349080
rect 470272 348780 470816 348784
rect 469032 347993 469576 347997
rect 469032 347697 469036 347993
rect 469036 347697 469572 347993
rect 469572 347697 469576 347993
rect 469032 347693 469576 347697
rect 470272 346908 470816 346912
rect 470272 346612 470276 346908
rect 470276 346612 470812 346908
rect 470812 346612 470816 346908
rect 470272 346608 470816 346612
rect 470272 328080 470816 328084
rect 470272 327784 470276 328080
rect 470276 327784 470812 328080
rect 470812 327784 470816 328080
rect 470272 327780 470816 327784
rect 469032 326993 469576 326997
rect 469032 326697 469036 326993
rect 469036 326697 469572 326993
rect 469572 326697 469576 326993
rect 469032 326693 469576 326697
rect 470272 325908 470816 325912
rect 470272 325612 470276 325908
rect 470276 325612 470812 325908
rect 470812 325612 470816 325908
rect 470272 325608 470816 325612
rect 470272 307080 470816 307084
rect 470272 306784 470276 307080
rect 470276 306784 470812 307080
rect 470812 306784 470816 307080
rect 470272 306780 470816 306784
rect 469032 305995 469576 305999
rect 469032 305699 469036 305995
rect 469036 305699 469572 305995
rect 469572 305699 469576 305995
rect 469032 305695 469576 305699
rect 470272 304908 470816 304912
rect 470272 304612 470276 304908
rect 470276 304612 470812 304908
rect 470812 304612 470816 304908
rect 470272 304608 470816 304612
rect 470272 286081 470816 286085
rect 470272 285785 470276 286081
rect 470276 285785 470812 286081
rect 470812 285785 470816 286081
rect 470272 285781 470816 285785
rect 469032 284996 469576 285000
rect 469032 284700 469036 284996
rect 469036 284700 469572 284996
rect 469572 284700 469576 284996
rect 469032 284696 469576 284700
rect 470272 283908 470816 283912
rect 470272 283612 470276 283908
rect 470276 283612 470812 283908
rect 470812 283612 470816 283908
rect 470272 283608 470816 283612
rect 470272 265081 470816 265085
rect 470272 264785 470276 265081
rect 470276 264785 470812 265081
rect 470812 264785 470816 265081
rect 470272 264781 470816 264785
rect 469032 263995 469576 263999
rect 469032 263699 469036 263995
rect 469036 263699 469572 263995
rect 469572 263699 469576 263995
rect 469032 263695 469576 263699
rect 470272 262908 470816 262912
rect 470272 262612 470276 262908
rect 470276 262612 470812 262908
rect 470812 262612 470816 262908
rect 470272 262608 470816 262612
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711002 -8694 711558
rect -8138 711002 -8106 711558
rect -8726 695334 -8106 711002
rect -8726 694778 -8694 695334
rect -8138 694778 -8106 695334
rect -8726 659334 -8106 694778
rect -8726 658778 -8694 659334
rect -8138 658778 -8106 659334
rect -8726 623334 -8106 658778
rect -8726 622778 -8694 623334
rect -8138 622778 -8106 623334
rect -8726 587334 -8106 622778
rect -8726 586778 -8694 587334
rect -8138 586778 -8106 587334
rect -8726 551334 -8106 586778
rect -8726 550778 -8694 551334
rect -8138 550778 -8106 551334
rect -8726 515334 -8106 550778
rect -8726 514778 -8694 515334
rect -8138 514778 -8106 515334
rect -8726 479334 -8106 514778
rect -8726 478778 -8694 479334
rect -8138 478778 -8106 479334
rect -8726 443334 -8106 478778
rect -8726 442778 -8694 443334
rect -8138 442778 -8106 443334
rect -8726 407334 -8106 442778
rect -8726 406778 -8694 407334
rect -8138 406778 -8106 407334
rect -8726 371334 -8106 406778
rect -8726 370778 -8694 371334
rect -8138 370778 -8106 371334
rect -8726 335334 -8106 370778
rect -8726 334778 -8694 335334
rect -8138 334778 -8106 335334
rect -8726 299334 -8106 334778
rect -8726 298778 -8694 299334
rect -8138 298778 -8106 299334
rect -8726 263334 -8106 298778
rect -8726 262778 -8694 263334
rect -8138 262778 -8106 263334
rect -8726 227334 -8106 262778
rect -8726 226778 -8694 227334
rect -8138 226778 -8106 227334
rect -8726 191334 -8106 226778
rect -8726 190778 -8694 191334
rect -8138 190778 -8106 191334
rect -8726 155334 -8106 190778
rect -8726 154778 -8694 155334
rect -8138 154778 -8106 155334
rect -8726 119334 -8106 154778
rect -8726 118778 -8694 119334
rect -8138 118778 -8106 119334
rect -8726 83334 -8106 118778
rect -8726 82778 -8694 83334
rect -8138 82778 -8106 83334
rect -8726 47334 -8106 82778
rect -8726 46778 -8694 47334
rect -8138 46778 -8106 47334
rect -8726 11334 -8106 46778
rect -8726 10778 -8694 11334
rect -8138 10778 -8106 11334
rect -8726 -7066 -8106 10778
rect -7766 710598 -7146 710630
rect -7766 710042 -7734 710598
rect -7178 710042 -7146 710598
rect -7766 694094 -7146 710042
rect -7766 693538 -7734 694094
rect -7178 693538 -7146 694094
rect -7766 658094 -7146 693538
rect -7766 657538 -7734 658094
rect -7178 657538 -7146 658094
rect -7766 622094 -7146 657538
rect -7766 621538 -7734 622094
rect -7178 621538 -7146 622094
rect -7766 586094 -7146 621538
rect -7766 585538 -7734 586094
rect -7178 585538 -7146 586094
rect -7766 550094 -7146 585538
rect -7766 549538 -7734 550094
rect -7178 549538 -7146 550094
rect -7766 514094 -7146 549538
rect -7766 513538 -7734 514094
rect -7178 513538 -7146 514094
rect -7766 478094 -7146 513538
rect -7766 477538 -7734 478094
rect -7178 477538 -7146 478094
rect -7766 442094 -7146 477538
rect -7766 441538 -7734 442094
rect -7178 441538 -7146 442094
rect -7766 406094 -7146 441538
rect -7766 405538 -7734 406094
rect -7178 405538 -7146 406094
rect -7766 370094 -7146 405538
rect -7766 369538 -7734 370094
rect -7178 369538 -7146 370094
rect -7766 334094 -7146 369538
rect -7766 333538 -7734 334094
rect -7178 333538 -7146 334094
rect -7766 298094 -7146 333538
rect -7766 297538 -7734 298094
rect -7178 297538 -7146 298094
rect -7766 262094 -7146 297538
rect -7766 261538 -7734 262094
rect -7178 261538 -7146 262094
rect -7766 226094 -7146 261538
rect -7766 225538 -7734 226094
rect -7178 225538 -7146 226094
rect -7766 190094 -7146 225538
rect -7766 189538 -7734 190094
rect -7178 189538 -7146 190094
rect -7766 154094 -7146 189538
rect -7766 153538 -7734 154094
rect -7178 153538 -7146 154094
rect -7766 118094 -7146 153538
rect -7766 117538 -7734 118094
rect -7178 117538 -7146 118094
rect -7766 82094 -7146 117538
rect -7766 81538 -7734 82094
rect -7178 81538 -7146 82094
rect -7766 46094 -7146 81538
rect -7766 45538 -7734 46094
rect -7178 45538 -7146 46094
rect -7766 10094 -7146 45538
rect -7766 9538 -7734 10094
rect -7178 9538 -7146 10094
rect -7766 -6106 -7146 9538
rect -6806 709638 -6186 709670
rect -6806 709082 -6774 709638
rect -6218 709082 -6186 709638
rect -6806 692854 -6186 709082
rect -6806 692298 -6774 692854
rect -6218 692298 -6186 692854
rect -6806 656854 -6186 692298
rect -6806 656298 -6774 656854
rect -6218 656298 -6186 656854
rect -6806 620854 -6186 656298
rect -6806 620298 -6774 620854
rect -6218 620298 -6186 620854
rect -6806 584854 -6186 620298
rect -6806 584298 -6774 584854
rect -6218 584298 -6186 584854
rect -6806 548854 -6186 584298
rect -6806 548298 -6774 548854
rect -6218 548298 -6186 548854
rect -6806 512854 -6186 548298
rect -6806 512298 -6774 512854
rect -6218 512298 -6186 512854
rect -6806 476854 -6186 512298
rect -6806 476298 -6774 476854
rect -6218 476298 -6186 476854
rect -6806 440854 -6186 476298
rect -6806 440298 -6774 440854
rect -6218 440298 -6186 440854
rect -6806 404854 -6186 440298
rect -6806 404298 -6774 404854
rect -6218 404298 -6186 404854
rect -6806 368854 -6186 404298
rect -6806 368298 -6774 368854
rect -6218 368298 -6186 368854
rect -6806 332854 -6186 368298
rect -6806 332298 -6774 332854
rect -6218 332298 -6186 332854
rect -6806 296854 -6186 332298
rect -6806 296298 -6774 296854
rect -6218 296298 -6186 296854
rect -6806 260854 -6186 296298
rect -6806 260298 -6774 260854
rect -6218 260298 -6186 260854
rect -6806 224854 -6186 260298
rect -6806 224298 -6774 224854
rect -6218 224298 -6186 224854
rect -6806 188854 -6186 224298
rect -6806 188298 -6774 188854
rect -6218 188298 -6186 188854
rect -6806 152854 -6186 188298
rect -6806 152298 -6774 152854
rect -6218 152298 -6186 152854
rect -6806 116854 -6186 152298
rect -6806 116298 -6774 116854
rect -6218 116298 -6186 116854
rect -6806 80854 -6186 116298
rect -6806 80298 -6774 80854
rect -6218 80298 -6186 80854
rect -6806 44854 -6186 80298
rect -6806 44298 -6774 44854
rect -6218 44298 -6186 44854
rect -6806 8854 -6186 44298
rect -6806 8298 -6774 8854
rect -6218 8298 -6186 8854
rect -6806 -5146 -6186 8298
rect -5846 708678 -5226 708710
rect -5846 708122 -5814 708678
rect -5258 708122 -5226 708678
rect -5846 691614 -5226 708122
rect -5846 691058 -5814 691614
rect -5258 691058 -5226 691614
rect -5846 655614 -5226 691058
rect -5846 655058 -5814 655614
rect -5258 655058 -5226 655614
rect -5846 619614 -5226 655058
rect -5846 619058 -5814 619614
rect -5258 619058 -5226 619614
rect -5846 583614 -5226 619058
rect -5846 583058 -5814 583614
rect -5258 583058 -5226 583614
rect -5846 547614 -5226 583058
rect -5846 547058 -5814 547614
rect -5258 547058 -5226 547614
rect -5846 511614 -5226 547058
rect -5846 511058 -5814 511614
rect -5258 511058 -5226 511614
rect -5846 475614 -5226 511058
rect -5846 475058 -5814 475614
rect -5258 475058 -5226 475614
rect -5846 439614 -5226 475058
rect -5846 439058 -5814 439614
rect -5258 439058 -5226 439614
rect -5846 403614 -5226 439058
rect -5846 403058 -5814 403614
rect -5258 403058 -5226 403614
rect -5846 367614 -5226 403058
rect -5846 367058 -5814 367614
rect -5258 367058 -5226 367614
rect -5846 331614 -5226 367058
rect -5846 331058 -5814 331614
rect -5258 331058 -5226 331614
rect -5846 295614 -5226 331058
rect -5846 295058 -5814 295614
rect -5258 295058 -5226 295614
rect -5846 259614 -5226 295058
rect -5846 259058 -5814 259614
rect -5258 259058 -5226 259614
rect -5846 223614 -5226 259058
rect -5846 223058 -5814 223614
rect -5258 223058 -5226 223614
rect -5846 187614 -5226 223058
rect -5846 187058 -5814 187614
rect -5258 187058 -5226 187614
rect -5846 151614 -5226 187058
rect -5846 151058 -5814 151614
rect -5258 151058 -5226 151614
rect -5846 115614 -5226 151058
rect -5846 115058 -5814 115614
rect -5258 115058 -5226 115614
rect -5846 79614 -5226 115058
rect -5846 79058 -5814 79614
rect -5258 79058 -5226 79614
rect -5846 43614 -5226 79058
rect -5846 43058 -5814 43614
rect -5258 43058 -5226 43614
rect -5846 7614 -5226 43058
rect -5846 7058 -5814 7614
rect -5258 7058 -5226 7614
rect -5846 -4186 -5226 7058
rect -4886 707718 -4266 707750
rect -4886 707162 -4854 707718
rect -4298 707162 -4266 707718
rect -4886 690374 -4266 707162
rect -4886 689818 -4854 690374
rect -4298 689818 -4266 690374
rect -4886 654374 -4266 689818
rect -4886 653818 -4854 654374
rect -4298 653818 -4266 654374
rect -4886 618374 -4266 653818
rect -4886 617818 -4854 618374
rect -4298 617818 -4266 618374
rect -4886 582374 -4266 617818
rect -4886 581818 -4854 582374
rect -4298 581818 -4266 582374
rect -4886 546374 -4266 581818
rect -4886 545818 -4854 546374
rect -4298 545818 -4266 546374
rect -4886 510374 -4266 545818
rect -4886 509818 -4854 510374
rect -4298 509818 -4266 510374
rect -4886 474374 -4266 509818
rect -4886 473818 -4854 474374
rect -4298 473818 -4266 474374
rect -4886 438374 -4266 473818
rect -4886 437818 -4854 438374
rect -4298 437818 -4266 438374
rect -4886 402374 -4266 437818
rect -4886 401818 -4854 402374
rect -4298 401818 -4266 402374
rect -4886 366374 -4266 401818
rect -4886 365818 -4854 366374
rect -4298 365818 -4266 366374
rect -4886 330374 -4266 365818
rect -4886 329818 -4854 330374
rect -4298 329818 -4266 330374
rect -4886 294374 -4266 329818
rect -4886 293818 -4854 294374
rect -4298 293818 -4266 294374
rect -4886 258374 -4266 293818
rect -4886 257818 -4854 258374
rect -4298 257818 -4266 258374
rect -4886 222374 -4266 257818
rect -4886 221818 -4854 222374
rect -4298 221818 -4266 222374
rect -4886 186374 -4266 221818
rect -4886 185818 -4854 186374
rect -4298 185818 -4266 186374
rect -4886 150374 -4266 185818
rect -4886 149818 -4854 150374
rect -4298 149818 -4266 150374
rect -4886 114374 -4266 149818
rect -4886 113818 -4854 114374
rect -4298 113818 -4266 114374
rect -4886 78374 -4266 113818
rect -4886 77818 -4854 78374
rect -4298 77818 -4266 78374
rect -4886 42374 -4266 77818
rect -4886 41818 -4854 42374
rect -4298 41818 -4266 42374
rect -4886 6374 -4266 41818
rect -4886 5818 -4854 6374
rect -4298 5818 -4266 6374
rect -4886 -3226 -4266 5818
rect -3926 706758 -3306 706790
rect -3926 706202 -3894 706758
rect -3338 706202 -3306 706758
rect -3926 689134 -3306 706202
rect -3926 688578 -3894 689134
rect -3338 688578 -3306 689134
rect -3926 653134 -3306 688578
rect -3926 652578 -3894 653134
rect -3338 652578 -3306 653134
rect -3926 617134 -3306 652578
rect -3926 616578 -3894 617134
rect -3338 616578 -3306 617134
rect -3926 581134 -3306 616578
rect -3926 580578 -3894 581134
rect -3338 580578 -3306 581134
rect -3926 545134 -3306 580578
rect -3926 544578 -3894 545134
rect -3338 544578 -3306 545134
rect -3926 509134 -3306 544578
rect -3926 508578 -3894 509134
rect -3338 508578 -3306 509134
rect -3926 473134 -3306 508578
rect -3926 472578 -3894 473134
rect -3338 472578 -3306 473134
rect -3926 437134 -3306 472578
rect -3926 436578 -3894 437134
rect -3338 436578 -3306 437134
rect -3926 401134 -3306 436578
rect -3926 400578 -3894 401134
rect -3338 400578 -3306 401134
rect -3926 365134 -3306 400578
rect -3926 364578 -3894 365134
rect -3338 364578 -3306 365134
rect -3926 329134 -3306 364578
rect -3926 328578 -3894 329134
rect -3338 328578 -3306 329134
rect -3926 293134 -3306 328578
rect -3926 292578 -3894 293134
rect -3338 292578 -3306 293134
rect -3926 257134 -3306 292578
rect -3926 256578 -3894 257134
rect -3338 256578 -3306 257134
rect -3926 221134 -3306 256578
rect -3926 220578 -3894 221134
rect -3338 220578 -3306 221134
rect -3926 185134 -3306 220578
rect -3926 184578 -3894 185134
rect -3338 184578 -3306 185134
rect -3926 149134 -3306 184578
rect -3926 148578 -3894 149134
rect -3338 148578 -3306 149134
rect -3926 113134 -3306 148578
rect -3926 112578 -3894 113134
rect -3338 112578 -3306 113134
rect -3926 77134 -3306 112578
rect -3926 76578 -3894 77134
rect -3338 76578 -3306 77134
rect -3926 41134 -3306 76578
rect -3926 40578 -3894 41134
rect -3338 40578 -3306 41134
rect -3926 5134 -3306 40578
rect -3926 4578 -3894 5134
rect -3338 4578 -3306 5134
rect -3926 -2266 -3306 4578
rect -2966 705798 -2346 705830
rect -2966 705242 -2934 705798
rect -2378 705242 -2346 705798
rect -2966 687894 -2346 705242
rect -2966 687338 -2934 687894
rect -2378 687338 -2346 687894
rect -2966 651894 -2346 687338
rect -2966 651338 -2934 651894
rect -2378 651338 -2346 651894
rect -2966 615894 -2346 651338
rect -2966 615338 -2934 615894
rect -2378 615338 -2346 615894
rect -2966 579894 -2346 615338
rect -2966 579338 -2934 579894
rect -2378 579338 -2346 579894
rect -2966 543894 -2346 579338
rect -2966 543338 -2934 543894
rect -2378 543338 -2346 543894
rect -2966 507894 -2346 543338
rect -2966 507338 -2934 507894
rect -2378 507338 -2346 507894
rect -2966 471894 -2346 507338
rect -2966 471338 -2934 471894
rect -2378 471338 -2346 471894
rect -2966 435894 -2346 471338
rect -2966 435338 -2934 435894
rect -2378 435338 -2346 435894
rect -2966 399894 -2346 435338
rect -2966 399338 -2934 399894
rect -2378 399338 -2346 399894
rect -2966 363894 -2346 399338
rect -2966 363338 -2934 363894
rect -2378 363338 -2346 363894
rect -2966 327894 -2346 363338
rect -2966 327338 -2934 327894
rect -2378 327338 -2346 327894
rect -2966 291894 -2346 327338
rect -2966 291338 -2934 291894
rect -2378 291338 -2346 291894
rect -2966 255894 -2346 291338
rect -2966 255338 -2934 255894
rect -2378 255338 -2346 255894
rect -2966 219894 -2346 255338
rect -2966 219338 -2934 219894
rect -2378 219338 -2346 219894
rect -2966 183894 -2346 219338
rect -2966 183338 -2934 183894
rect -2378 183338 -2346 183894
rect -2966 147894 -2346 183338
rect -2966 147338 -2934 147894
rect -2378 147338 -2346 147894
rect -2966 111894 -2346 147338
rect -2966 111338 -2934 111894
rect -2378 111338 -2346 111894
rect -2966 75894 -2346 111338
rect -2966 75338 -2934 75894
rect -2378 75338 -2346 75894
rect -2966 39894 -2346 75338
rect -2966 39338 -2934 39894
rect -2378 39338 -2346 39894
rect -2966 3894 -2346 39338
rect -2966 3338 -2934 3894
rect -2378 3338 -2346 3894
rect -2966 -1306 -2346 3338
rect -2006 704838 -1386 704870
rect -2006 704282 -1974 704838
rect -1418 704282 -1386 704838
rect -2006 686654 -1386 704282
rect -2006 686098 -1974 686654
rect -1418 686098 -1386 686654
rect -2006 650654 -1386 686098
rect -2006 650098 -1974 650654
rect -1418 650098 -1386 650654
rect -2006 614654 -1386 650098
rect -2006 614098 -1974 614654
rect -1418 614098 -1386 614654
rect -2006 578654 -1386 614098
rect -2006 578098 -1974 578654
rect -1418 578098 -1386 578654
rect -2006 542654 -1386 578098
rect -2006 542098 -1974 542654
rect -1418 542098 -1386 542654
rect -2006 506654 -1386 542098
rect -2006 506098 -1974 506654
rect -1418 506098 -1386 506654
rect -2006 470654 -1386 506098
rect -2006 470098 -1974 470654
rect -1418 470098 -1386 470654
rect -2006 434654 -1386 470098
rect -2006 434098 -1974 434654
rect -1418 434098 -1386 434654
rect -2006 398654 -1386 434098
rect -2006 398098 -1974 398654
rect -1418 398098 -1386 398654
rect -2006 362654 -1386 398098
rect -2006 362098 -1974 362654
rect -1418 362098 -1386 362654
rect -2006 326654 -1386 362098
rect -2006 326098 -1974 326654
rect -1418 326098 -1386 326654
rect -2006 290654 -1386 326098
rect -2006 290098 -1974 290654
rect -1418 290098 -1386 290654
rect -2006 254654 -1386 290098
rect -2006 254098 -1974 254654
rect -1418 254098 -1386 254654
rect -2006 218654 -1386 254098
rect -2006 218098 -1974 218654
rect -1418 218098 -1386 218654
rect -2006 182654 -1386 218098
rect -2006 182098 -1974 182654
rect -1418 182098 -1386 182654
rect -2006 146654 -1386 182098
rect -2006 146098 -1974 146654
rect -1418 146098 -1386 146654
rect -2006 110654 -1386 146098
rect -2006 110098 -1974 110654
rect -1418 110098 -1386 110654
rect -2006 74654 -1386 110098
rect -2006 74098 -1974 74654
rect -1418 74098 -1386 74654
rect -2006 38654 -1386 74098
rect -2006 38098 -1974 38654
rect -1418 38098 -1386 38654
rect -2006 2654 -1386 38098
rect -2006 2098 -1974 2654
rect -1418 2098 -1386 2654
rect -2006 -346 -1386 2098
rect -2006 -902 -1974 -346
rect -1418 -902 -1386 -346
rect -2006 -934 -1386 -902
rect 994 704838 1614 711590
rect 994 704282 1026 704838
rect 1582 704282 1614 704838
rect 994 686654 1614 704282
rect 994 686098 1026 686654
rect 1582 686098 1614 686654
rect 994 650654 1614 686098
rect 994 650098 1026 650654
rect 1582 650098 1614 650654
rect 994 614654 1614 650098
rect 994 614098 1026 614654
rect 1582 614098 1614 614654
rect 994 578654 1614 614098
rect 994 578098 1026 578654
rect 1582 578098 1614 578654
rect 994 542654 1614 578098
rect 994 542098 1026 542654
rect 1582 542098 1614 542654
rect 994 506654 1614 542098
rect 994 506098 1026 506654
rect 1582 506098 1614 506654
rect 994 470654 1614 506098
rect 994 470098 1026 470654
rect 1582 470098 1614 470654
rect 994 434654 1614 470098
rect 994 434098 1026 434654
rect 1582 434098 1614 434654
rect 994 398654 1614 434098
rect 994 398098 1026 398654
rect 1582 398098 1614 398654
rect 994 362654 1614 398098
rect 994 362098 1026 362654
rect 1582 362098 1614 362654
rect 994 326654 1614 362098
rect 994 326098 1026 326654
rect 1582 326098 1614 326654
rect 994 290654 1614 326098
rect 994 290098 1026 290654
rect 1582 290098 1614 290654
rect 994 254654 1614 290098
rect 994 254098 1026 254654
rect 1582 254098 1614 254654
rect 994 218654 1614 254098
rect 994 218098 1026 218654
rect 1582 218098 1614 218654
rect 994 182654 1614 218098
rect 994 182098 1026 182654
rect 1582 182098 1614 182654
rect 994 146654 1614 182098
rect 994 146098 1026 146654
rect 1582 146098 1614 146654
rect 994 110654 1614 146098
rect 994 110098 1026 110654
rect 1582 110098 1614 110654
rect 994 74654 1614 110098
rect 994 74098 1026 74654
rect 1582 74098 1614 74654
rect 994 38654 1614 74098
rect 994 38098 1026 38654
rect 1582 38098 1614 38654
rect 994 2654 1614 38098
rect 994 2098 1026 2654
rect 1582 2098 1614 2654
rect 994 -346 1614 2098
rect 994 -902 1026 -346
rect 1582 -902 1614 -346
rect -2966 -1862 -2934 -1306
rect -2378 -1862 -2346 -1306
rect -2966 -1894 -2346 -1862
rect -3926 -2822 -3894 -2266
rect -3338 -2822 -3306 -2266
rect -3926 -2854 -3306 -2822
rect -4886 -3782 -4854 -3226
rect -4298 -3782 -4266 -3226
rect -4886 -3814 -4266 -3782
rect -5846 -4742 -5814 -4186
rect -5258 -4742 -5226 -4186
rect -5846 -4774 -5226 -4742
rect -6806 -5702 -6774 -5146
rect -6218 -5702 -6186 -5146
rect -6806 -5734 -6186 -5702
rect -7766 -6662 -7734 -6106
rect -7178 -6662 -7146 -6106
rect -7766 -6694 -7146 -6662
rect -8726 -7622 -8694 -7066
rect -8138 -7622 -8106 -7066
rect -8726 -7654 -8106 -7622
rect 994 -7654 1614 -902
rect 2234 705798 2854 711590
rect 2234 705242 2266 705798
rect 2822 705242 2854 705798
rect 2234 687894 2854 705242
rect 2234 687338 2266 687894
rect 2822 687338 2854 687894
rect 2234 651894 2854 687338
rect 2234 651338 2266 651894
rect 2822 651338 2854 651894
rect 2234 615894 2854 651338
rect 2234 615338 2266 615894
rect 2822 615338 2854 615894
rect 2234 579894 2854 615338
rect 2234 579338 2266 579894
rect 2822 579338 2854 579894
rect 2234 543894 2854 579338
rect 2234 543338 2266 543894
rect 2822 543338 2854 543894
rect 2234 507894 2854 543338
rect 2234 507338 2266 507894
rect 2822 507338 2854 507894
rect 2234 471894 2854 507338
rect 2234 471338 2266 471894
rect 2822 471338 2854 471894
rect 2234 435894 2854 471338
rect 2234 435338 2266 435894
rect 2822 435338 2854 435894
rect 2234 399894 2854 435338
rect 2234 399338 2266 399894
rect 2822 399338 2854 399894
rect 2234 363894 2854 399338
rect 2234 363338 2266 363894
rect 2822 363338 2854 363894
rect 2234 327894 2854 363338
rect 2234 327338 2266 327894
rect 2822 327338 2854 327894
rect 2234 291894 2854 327338
rect 2234 291338 2266 291894
rect 2822 291338 2854 291894
rect 2234 255894 2854 291338
rect 2234 255338 2266 255894
rect 2822 255338 2854 255894
rect 2234 219894 2854 255338
rect 2234 219338 2266 219894
rect 2822 219338 2854 219894
rect 2234 183894 2854 219338
rect 2234 183338 2266 183894
rect 2822 183338 2854 183894
rect 2234 147894 2854 183338
rect 2234 147338 2266 147894
rect 2822 147338 2854 147894
rect 2234 111894 2854 147338
rect 2234 111338 2266 111894
rect 2822 111338 2854 111894
rect 2234 75894 2854 111338
rect 2234 75338 2266 75894
rect 2822 75338 2854 75894
rect 2234 39894 2854 75338
rect 2234 39338 2266 39894
rect 2822 39338 2854 39894
rect 2234 3894 2854 39338
rect 2234 3338 2266 3894
rect 2822 3338 2854 3894
rect 2234 -1306 2854 3338
rect 2234 -1862 2266 -1306
rect 2822 -1862 2854 -1306
rect 2234 -7654 2854 -1862
rect 3474 706758 4094 711590
rect 3474 706202 3506 706758
rect 4062 706202 4094 706758
rect 3474 689134 4094 706202
rect 3474 688578 3506 689134
rect 4062 688578 4094 689134
rect 3474 653134 4094 688578
rect 3474 652578 3506 653134
rect 4062 652578 4094 653134
rect 3474 617134 4094 652578
rect 3474 616578 3506 617134
rect 4062 616578 4094 617134
rect 3474 581134 4094 616578
rect 3474 580578 3506 581134
rect 4062 580578 4094 581134
rect 3474 545134 4094 580578
rect 3474 544578 3506 545134
rect 4062 544578 4094 545134
rect 3474 509134 4094 544578
rect 3474 508578 3506 509134
rect 4062 508578 4094 509134
rect 3474 473134 4094 508578
rect 3474 472578 3506 473134
rect 4062 472578 4094 473134
rect 3474 437134 4094 472578
rect 3474 436578 3506 437134
rect 4062 436578 4094 437134
rect 3474 401134 4094 436578
rect 3474 400578 3506 401134
rect 4062 400578 4094 401134
rect 3474 365134 4094 400578
rect 3474 364578 3506 365134
rect 4062 364578 4094 365134
rect 3474 329134 4094 364578
rect 3474 328578 3506 329134
rect 4062 328578 4094 329134
rect 3474 293134 4094 328578
rect 3474 292578 3506 293134
rect 4062 292578 4094 293134
rect 3474 257134 4094 292578
rect 3474 256578 3506 257134
rect 4062 256578 4094 257134
rect 3474 221134 4094 256578
rect 3474 220578 3506 221134
rect 4062 220578 4094 221134
rect 3474 185134 4094 220578
rect 3474 184578 3506 185134
rect 4062 184578 4094 185134
rect 3474 149134 4094 184578
rect 3474 148578 3506 149134
rect 4062 148578 4094 149134
rect 3474 113134 4094 148578
rect 3474 112578 3506 113134
rect 4062 112578 4094 113134
rect 3474 77134 4094 112578
rect 3474 76578 3506 77134
rect 4062 76578 4094 77134
rect 3474 41134 4094 76578
rect 3474 40578 3506 41134
rect 4062 40578 4094 41134
rect 3474 5134 4094 40578
rect 3474 4578 3506 5134
rect 4062 4578 4094 5134
rect 3474 -2266 4094 4578
rect 3474 -2822 3506 -2266
rect 4062 -2822 4094 -2266
rect 3474 -7654 4094 -2822
rect 4714 707718 5334 711590
rect 4714 707162 4746 707718
rect 5302 707162 5334 707718
rect 4714 690374 5334 707162
rect 4714 689818 4746 690374
rect 5302 689818 5334 690374
rect 4714 654374 5334 689818
rect 4714 653818 4746 654374
rect 5302 653818 5334 654374
rect 4714 618374 5334 653818
rect 4714 617818 4746 618374
rect 5302 617818 5334 618374
rect 4714 582374 5334 617818
rect 4714 581818 4746 582374
rect 5302 581818 5334 582374
rect 4714 546374 5334 581818
rect 4714 545818 4746 546374
rect 5302 545818 5334 546374
rect 4714 510374 5334 545818
rect 4714 509818 4746 510374
rect 5302 509818 5334 510374
rect 4714 474374 5334 509818
rect 4714 473818 4746 474374
rect 5302 473818 5334 474374
rect 4714 438374 5334 473818
rect 4714 437818 4746 438374
rect 5302 437818 5334 438374
rect 4714 402374 5334 437818
rect 4714 401818 4746 402374
rect 5302 401818 5334 402374
rect 4714 366374 5334 401818
rect 4714 365818 4746 366374
rect 5302 365818 5334 366374
rect 4714 330374 5334 365818
rect 4714 329818 4746 330374
rect 5302 329818 5334 330374
rect 4714 294374 5334 329818
rect 4714 293818 4746 294374
rect 5302 293818 5334 294374
rect 4714 258374 5334 293818
rect 4714 257818 4746 258374
rect 5302 257818 5334 258374
rect 4714 222374 5334 257818
rect 4714 221818 4746 222374
rect 5302 221818 5334 222374
rect 4714 186374 5334 221818
rect 4714 185818 4746 186374
rect 5302 185818 5334 186374
rect 4714 150374 5334 185818
rect 4714 149818 4746 150374
rect 5302 149818 5334 150374
rect 4714 114374 5334 149818
rect 4714 113818 4746 114374
rect 5302 113818 5334 114374
rect 4714 78374 5334 113818
rect 4714 77818 4746 78374
rect 5302 77818 5334 78374
rect 4714 42374 5334 77818
rect 4714 41818 4746 42374
rect 5302 41818 5334 42374
rect 4714 6374 5334 41818
rect 4714 5818 4746 6374
rect 5302 5818 5334 6374
rect 4714 -3226 5334 5818
rect 4714 -3782 4746 -3226
rect 5302 -3782 5334 -3226
rect 4714 -7654 5334 -3782
rect 5954 708678 6574 711590
rect 5954 708122 5986 708678
rect 6542 708122 6574 708678
rect 5954 691614 6574 708122
rect 5954 691058 5986 691614
rect 6542 691058 6574 691614
rect 5954 655614 6574 691058
rect 5954 655058 5986 655614
rect 6542 655058 6574 655614
rect 5954 619614 6574 655058
rect 5954 619058 5986 619614
rect 6542 619058 6574 619614
rect 5954 583614 6574 619058
rect 5954 583058 5986 583614
rect 6542 583058 6574 583614
rect 5954 547614 6574 583058
rect 5954 547058 5986 547614
rect 6542 547058 6574 547614
rect 5954 511614 6574 547058
rect 5954 511058 5986 511614
rect 6542 511058 6574 511614
rect 5954 475614 6574 511058
rect 5954 475058 5986 475614
rect 6542 475058 6574 475614
rect 5954 439614 6574 475058
rect 5954 439058 5986 439614
rect 6542 439058 6574 439614
rect 5954 403614 6574 439058
rect 5954 403058 5986 403614
rect 6542 403058 6574 403614
rect 5954 367614 6574 403058
rect 5954 367058 5986 367614
rect 6542 367058 6574 367614
rect 5954 331614 6574 367058
rect 5954 331058 5986 331614
rect 6542 331058 6574 331614
rect 5954 295614 6574 331058
rect 5954 295058 5986 295614
rect 6542 295058 6574 295614
rect 5954 259614 6574 295058
rect 5954 259058 5986 259614
rect 6542 259058 6574 259614
rect 5954 223614 6574 259058
rect 5954 223058 5986 223614
rect 6542 223058 6574 223614
rect 5954 187614 6574 223058
rect 5954 187058 5986 187614
rect 6542 187058 6574 187614
rect 5954 151614 6574 187058
rect 5954 151058 5986 151614
rect 6542 151058 6574 151614
rect 5954 115614 6574 151058
rect 5954 115058 5986 115614
rect 6542 115058 6574 115614
rect 5954 79614 6574 115058
rect 5954 79058 5986 79614
rect 6542 79058 6574 79614
rect 5954 43614 6574 79058
rect 5954 43058 5986 43614
rect 6542 43058 6574 43614
rect 5954 7614 6574 43058
rect 5954 7058 5986 7614
rect 6542 7058 6574 7614
rect 5954 -4186 6574 7058
rect 5954 -4742 5986 -4186
rect 6542 -4742 6574 -4186
rect 5954 -7654 6574 -4742
rect 7194 709638 7814 711590
rect 7194 709082 7226 709638
rect 7782 709082 7814 709638
rect 7194 692854 7814 709082
rect 7194 692298 7226 692854
rect 7782 692298 7814 692854
rect 7194 656854 7814 692298
rect 7194 656298 7226 656854
rect 7782 656298 7814 656854
rect 7194 620854 7814 656298
rect 7194 620298 7226 620854
rect 7782 620298 7814 620854
rect 7194 584854 7814 620298
rect 7194 584298 7226 584854
rect 7782 584298 7814 584854
rect 7194 548854 7814 584298
rect 7194 548298 7226 548854
rect 7782 548298 7814 548854
rect 7194 512854 7814 548298
rect 7194 512298 7226 512854
rect 7782 512298 7814 512854
rect 7194 476854 7814 512298
rect 7194 476298 7226 476854
rect 7782 476298 7814 476854
rect 7194 440854 7814 476298
rect 7194 440298 7226 440854
rect 7782 440298 7814 440854
rect 7194 404854 7814 440298
rect 7194 404298 7226 404854
rect 7782 404298 7814 404854
rect 7194 368854 7814 404298
rect 7194 368298 7226 368854
rect 7782 368298 7814 368854
rect 7194 332854 7814 368298
rect 7194 332298 7226 332854
rect 7782 332298 7814 332854
rect 7194 296854 7814 332298
rect 7194 296298 7226 296854
rect 7782 296298 7814 296854
rect 7194 260854 7814 296298
rect 7194 260298 7226 260854
rect 7782 260298 7814 260854
rect 7194 224854 7814 260298
rect 7194 224298 7226 224854
rect 7782 224298 7814 224854
rect 7194 188854 7814 224298
rect 7194 188298 7226 188854
rect 7782 188298 7814 188854
rect 7194 152854 7814 188298
rect 7194 152298 7226 152854
rect 7782 152298 7814 152854
rect 7194 116854 7814 152298
rect 7194 116298 7226 116854
rect 7782 116298 7814 116854
rect 7194 80854 7814 116298
rect 7194 80298 7226 80854
rect 7782 80298 7814 80854
rect 7194 44854 7814 80298
rect 7194 44298 7226 44854
rect 7782 44298 7814 44854
rect 7194 8854 7814 44298
rect 7194 8298 7226 8854
rect 7782 8298 7814 8854
rect 7194 -5146 7814 8298
rect 7194 -5702 7226 -5146
rect 7782 -5702 7814 -5146
rect 7194 -7654 7814 -5702
rect 8434 710598 9054 711590
rect 8434 710042 8466 710598
rect 9022 710042 9054 710598
rect 8434 694094 9054 710042
rect 8434 693538 8466 694094
rect 9022 693538 9054 694094
rect 8434 658094 9054 693538
rect 8434 657538 8466 658094
rect 9022 657538 9054 658094
rect 8434 622094 9054 657538
rect 8434 621538 8466 622094
rect 9022 621538 9054 622094
rect 8434 586094 9054 621538
rect 8434 585538 8466 586094
rect 9022 585538 9054 586094
rect 8434 550094 9054 585538
rect 8434 549538 8466 550094
rect 9022 549538 9054 550094
rect 8434 514094 9054 549538
rect 8434 513538 8466 514094
rect 9022 513538 9054 514094
rect 8434 478094 9054 513538
rect 8434 477538 8466 478094
rect 9022 477538 9054 478094
rect 8434 442094 9054 477538
rect 8434 441538 8466 442094
rect 9022 441538 9054 442094
rect 8434 406094 9054 441538
rect 8434 405538 8466 406094
rect 9022 405538 9054 406094
rect 8434 370094 9054 405538
rect 8434 369538 8466 370094
rect 9022 369538 9054 370094
rect 8434 334094 9054 369538
rect 8434 333538 8466 334094
rect 9022 333538 9054 334094
rect 8434 298094 9054 333538
rect 8434 297538 8466 298094
rect 9022 297538 9054 298094
rect 8434 262094 9054 297538
rect 8434 261538 8466 262094
rect 9022 261538 9054 262094
rect 8434 226094 9054 261538
rect 8434 225538 8466 226094
rect 9022 225538 9054 226094
rect 8434 190094 9054 225538
rect 8434 189538 8466 190094
rect 9022 189538 9054 190094
rect 8434 154094 9054 189538
rect 8434 153538 8466 154094
rect 9022 153538 9054 154094
rect 8434 118094 9054 153538
rect 8434 117538 8466 118094
rect 9022 117538 9054 118094
rect 8434 82094 9054 117538
rect 8434 81538 8466 82094
rect 9022 81538 9054 82094
rect 8434 46094 9054 81538
rect 8434 45538 8466 46094
rect 9022 45538 9054 46094
rect 8434 10094 9054 45538
rect 8434 9538 8466 10094
rect 9022 9538 9054 10094
rect 8434 -6106 9054 9538
rect 8434 -6662 8466 -6106
rect 9022 -6662 9054 -6106
rect 8434 -7654 9054 -6662
rect 9674 711558 10294 711590
rect 9674 711002 9706 711558
rect 10262 711002 10294 711558
rect 9674 695334 10294 711002
rect 9674 694778 9706 695334
rect 10262 694778 10294 695334
rect 9674 659334 10294 694778
rect 9674 658778 9706 659334
rect 10262 658778 10294 659334
rect 9674 623334 10294 658778
rect 9674 622778 9706 623334
rect 10262 622778 10294 623334
rect 9674 587334 10294 622778
rect 9674 586778 9706 587334
rect 10262 586778 10294 587334
rect 9674 551334 10294 586778
rect 9674 550778 9706 551334
rect 10262 550778 10294 551334
rect 9674 515334 10294 550778
rect 9674 514778 9706 515334
rect 10262 514778 10294 515334
rect 9674 479334 10294 514778
rect 9674 478778 9706 479334
rect 10262 478778 10294 479334
rect 9674 443334 10294 478778
rect 9674 442778 9706 443334
rect 10262 442778 10294 443334
rect 9674 407334 10294 442778
rect 9674 406778 9706 407334
rect 10262 406778 10294 407334
rect 9674 371334 10294 406778
rect 9674 370778 9706 371334
rect 10262 370778 10294 371334
rect 9674 335334 10294 370778
rect 9674 334778 9706 335334
rect 10262 334778 10294 335334
rect 9674 299334 10294 334778
rect 9674 298778 9706 299334
rect 10262 298778 10294 299334
rect 9674 263334 10294 298778
rect 9674 262778 9706 263334
rect 10262 262778 10294 263334
rect 9674 227334 10294 262778
rect 9674 226778 9706 227334
rect 10262 226778 10294 227334
rect 9674 191334 10294 226778
rect 9674 190778 9706 191334
rect 10262 190778 10294 191334
rect 9674 155334 10294 190778
rect 9674 154778 9706 155334
rect 10262 154778 10294 155334
rect 9674 119334 10294 154778
rect 9674 118778 9706 119334
rect 10262 118778 10294 119334
rect 9674 83334 10294 118778
rect 9674 82778 9706 83334
rect 10262 82778 10294 83334
rect 9674 47334 10294 82778
rect 9674 46778 9706 47334
rect 10262 46778 10294 47334
rect 9674 11334 10294 46778
rect 9674 10778 9706 11334
rect 10262 10778 10294 11334
rect 9674 -7066 10294 10778
rect 9674 -7622 9706 -7066
rect 10262 -7622 10294 -7066
rect 9674 -7654 10294 -7622
rect 36994 704838 37614 711590
rect 36994 704282 37026 704838
rect 37582 704282 37614 704838
rect 36994 686654 37614 704282
rect 36994 686098 37026 686654
rect 37582 686098 37614 686654
rect 36994 650654 37614 686098
rect 36994 650098 37026 650654
rect 37582 650098 37614 650654
rect 36994 614654 37614 650098
rect 36994 614098 37026 614654
rect 37582 614098 37614 614654
rect 36994 578654 37614 614098
rect 36994 578098 37026 578654
rect 37582 578098 37614 578654
rect 36994 542654 37614 578098
rect 36994 542098 37026 542654
rect 37582 542098 37614 542654
rect 36994 506654 37614 542098
rect 36994 506098 37026 506654
rect 37582 506098 37614 506654
rect 36994 470654 37614 506098
rect 36994 470098 37026 470654
rect 37582 470098 37614 470654
rect 36994 434654 37614 470098
rect 36994 434098 37026 434654
rect 37582 434098 37614 434654
rect 36994 398654 37614 434098
rect 36994 398098 37026 398654
rect 37582 398098 37614 398654
rect 36994 362654 37614 398098
rect 36994 362098 37026 362654
rect 37582 362098 37614 362654
rect 36994 326654 37614 362098
rect 36994 326098 37026 326654
rect 37582 326098 37614 326654
rect 36994 290654 37614 326098
rect 36994 290098 37026 290654
rect 37582 290098 37614 290654
rect 36994 254654 37614 290098
rect 36994 254098 37026 254654
rect 37582 254098 37614 254654
rect 36994 218654 37614 254098
rect 36994 218098 37026 218654
rect 37582 218098 37614 218654
rect 36994 182654 37614 218098
rect 36994 182098 37026 182654
rect 37582 182098 37614 182654
rect 36994 146654 37614 182098
rect 36994 146098 37026 146654
rect 37582 146098 37614 146654
rect 36994 110654 37614 146098
rect 36994 110098 37026 110654
rect 37582 110098 37614 110654
rect 36994 74654 37614 110098
rect 36994 74098 37026 74654
rect 37582 74098 37614 74654
rect 36994 38654 37614 74098
rect 36994 38098 37026 38654
rect 37582 38098 37614 38654
rect 36994 2654 37614 38098
rect 36994 2098 37026 2654
rect 37582 2098 37614 2654
rect 36994 -346 37614 2098
rect 36994 -902 37026 -346
rect 37582 -902 37614 -346
rect 36994 -7654 37614 -902
rect 38234 705798 38854 711590
rect 38234 705242 38266 705798
rect 38822 705242 38854 705798
rect 38234 687894 38854 705242
rect 38234 687338 38266 687894
rect 38822 687338 38854 687894
rect 38234 651894 38854 687338
rect 38234 651338 38266 651894
rect 38822 651338 38854 651894
rect 38234 615894 38854 651338
rect 38234 615338 38266 615894
rect 38822 615338 38854 615894
rect 38234 579894 38854 615338
rect 38234 579338 38266 579894
rect 38822 579338 38854 579894
rect 38234 543894 38854 579338
rect 38234 543338 38266 543894
rect 38822 543338 38854 543894
rect 38234 507894 38854 543338
rect 38234 507338 38266 507894
rect 38822 507338 38854 507894
rect 38234 471894 38854 507338
rect 38234 471338 38266 471894
rect 38822 471338 38854 471894
rect 38234 435894 38854 471338
rect 38234 435338 38266 435894
rect 38822 435338 38854 435894
rect 38234 399894 38854 435338
rect 38234 399338 38266 399894
rect 38822 399338 38854 399894
rect 38234 363894 38854 399338
rect 38234 363338 38266 363894
rect 38822 363338 38854 363894
rect 38234 327894 38854 363338
rect 38234 327338 38266 327894
rect 38822 327338 38854 327894
rect 38234 291894 38854 327338
rect 38234 291338 38266 291894
rect 38822 291338 38854 291894
rect 38234 255894 38854 291338
rect 38234 255338 38266 255894
rect 38822 255338 38854 255894
rect 38234 219894 38854 255338
rect 38234 219338 38266 219894
rect 38822 219338 38854 219894
rect 38234 183894 38854 219338
rect 38234 183338 38266 183894
rect 38822 183338 38854 183894
rect 38234 147894 38854 183338
rect 38234 147338 38266 147894
rect 38822 147338 38854 147894
rect 38234 111894 38854 147338
rect 38234 111338 38266 111894
rect 38822 111338 38854 111894
rect 38234 75894 38854 111338
rect 38234 75338 38266 75894
rect 38822 75338 38854 75894
rect 38234 39894 38854 75338
rect 38234 39338 38266 39894
rect 38822 39338 38854 39894
rect 38234 3894 38854 39338
rect 38234 3338 38266 3894
rect 38822 3338 38854 3894
rect 38234 -1306 38854 3338
rect 38234 -1862 38266 -1306
rect 38822 -1862 38854 -1306
rect 38234 -7654 38854 -1862
rect 39474 706758 40094 711590
rect 39474 706202 39506 706758
rect 40062 706202 40094 706758
rect 39474 689134 40094 706202
rect 39474 688578 39506 689134
rect 40062 688578 40094 689134
rect 39474 653134 40094 688578
rect 39474 652578 39506 653134
rect 40062 652578 40094 653134
rect 39474 617134 40094 652578
rect 39474 616578 39506 617134
rect 40062 616578 40094 617134
rect 39474 581134 40094 616578
rect 39474 580578 39506 581134
rect 40062 580578 40094 581134
rect 39474 545134 40094 580578
rect 39474 544578 39506 545134
rect 40062 544578 40094 545134
rect 39474 509134 40094 544578
rect 39474 508578 39506 509134
rect 40062 508578 40094 509134
rect 39474 473134 40094 508578
rect 39474 472578 39506 473134
rect 40062 472578 40094 473134
rect 39474 437134 40094 472578
rect 39474 436578 39506 437134
rect 40062 436578 40094 437134
rect 39474 401134 40094 436578
rect 39474 400578 39506 401134
rect 40062 400578 40094 401134
rect 39474 365134 40094 400578
rect 39474 364578 39506 365134
rect 40062 364578 40094 365134
rect 39474 329134 40094 364578
rect 39474 328578 39506 329134
rect 40062 328578 40094 329134
rect 39474 293134 40094 328578
rect 39474 292578 39506 293134
rect 40062 292578 40094 293134
rect 39474 257134 40094 292578
rect 39474 256578 39506 257134
rect 40062 256578 40094 257134
rect 39474 221134 40094 256578
rect 39474 220578 39506 221134
rect 40062 220578 40094 221134
rect 39474 185134 40094 220578
rect 39474 184578 39506 185134
rect 40062 184578 40094 185134
rect 39474 149134 40094 184578
rect 39474 148578 39506 149134
rect 40062 148578 40094 149134
rect 39474 113134 40094 148578
rect 39474 112578 39506 113134
rect 40062 112578 40094 113134
rect 39474 77134 40094 112578
rect 39474 76578 39506 77134
rect 40062 76578 40094 77134
rect 39474 41134 40094 76578
rect 39474 40578 39506 41134
rect 40062 40578 40094 41134
rect 39474 5134 40094 40578
rect 39474 4578 39506 5134
rect 40062 4578 40094 5134
rect 39474 -2266 40094 4578
rect 39474 -2822 39506 -2266
rect 40062 -2822 40094 -2266
rect 39474 -7654 40094 -2822
rect 40714 707718 41334 711590
rect 40714 707162 40746 707718
rect 41302 707162 41334 707718
rect 40714 690374 41334 707162
rect 40714 689818 40746 690374
rect 41302 689818 41334 690374
rect 40714 654374 41334 689818
rect 40714 653818 40746 654374
rect 41302 653818 41334 654374
rect 40714 618374 41334 653818
rect 40714 617818 40746 618374
rect 41302 617818 41334 618374
rect 40714 582374 41334 617818
rect 40714 581818 40746 582374
rect 41302 581818 41334 582374
rect 40714 546374 41334 581818
rect 40714 545818 40746 546374
rect 41302 545818 41334 546374
rect 40714 510374 41334 545818
rect 40714 509818 40746 510374
rect 41302 509818 41334 510374
rect 40714 474374 41334 509818
rect 40714 473818 40746 474374
rect 41302 473818 41334 474374
rect 40714 438374 41334 473818
rect 40714 437818 40746 438374
rect 41302 437818 41334 438374
rect 40714 402374 41334 437818
rect 40714 401818 40746 402374
rect 41302 401818 41334 402374
rect 40714 366374 41334 401818
rect 40714 365818 40746 366374
rect 41302 365818 41334 366374
rect 40714 330374 41334 365818
rect 40714 329818 40746 330374
rect 41302 329818 41334 330374
rect 40714 294374 41334 329818
rect 40714 293818 40746 294374
rect 41302 293818 41334 294374
rect 40714 258374 41334 293818
rect 40714 257818 40746 258374
rect 41302 257818 41334 258374
rect 40714 222374 41334 257818
rect 40714 221818 40746 222374
rect 41302 221818 41334 222374
rect 40714 186374 41334 221818
rect 40714 185818 40746 186374
rect 41302 185818 41334 186374
rect 40714 150374 41334 185818
rect 40714 149818 40746 150374
rect 41302 149818 41334 150374
rect 40714 114374 41334 149818
rect 40714 113818 40746 114374
rect 41302 113818 41334 114374
rect 40714 78374 41334 113818
rect 40714 77818 40746 78374
rect 41302 77818 41334 78374
rect 40714 42374 41334 77818
rect 40714 41818 40746 42374
rect 41302 41818 41334 42374
rect 40714 6374 41334 41818
rect 40714 5818 40746 6374
rect 41302 5818 41334 6374
rect 40714 -3226 41334 5818
rect 40714 -3782 40746 -3226
rect 41302 -3782 41334 -3226
rect 40714 -7654 41334 -3782
rect 41954 708678 42574 711590
rect 41954 708122 41986 708678
rect 42542 708122 42574 708678
rect 41954 691614 42574 708122
rect 41954 691058 41986 691614
rect 42542 691058 42574 691614
rect 41954 655614 42574 691058
rect 41954 655058 41986 655614
rect 42542 655058 42574 655614
rect 41954 619614 42574 655058
rect 41954 619058 41986 619614
rect 42542 619058 42574 619614
rect 41954 583614 42574 619058
rect 41954 583058 41986 583614
rect 42542 583058 42574 583614
rect 41954 547614 42574 583058
rect 41954 547058 41986 547614
rect 42542 547058 42574 547614
rect 41954 511614 42574 547058
rect 41954 511058 41986 511614
rect 42542 511058 42574 511614
rect 41954 475614 42574 511058
rect 41954 475058 41986 475614
rect 42542 475058 42574 475614
rect 41954 439614 42574 475058
rect 41954 439058 41986 439614
rect 42542 439058 42574 439614
rect 41954 403614 42574 439058
rect 41954 403058 41986 403614
rect 42542 403058 42574 403614
rect 41954 367614 42574 403058
rect 41954 367058 41986 367614
rect 42542 367058 42574 367614
rect 41954 331614 42574 367058
rect 41954 331058 41986 331614
rect 42542 331058 42574 331614
rect 41954 295614 42574 331058
rect 41954 295058 41986 295614
rect 42542 295058 42574 295614
rect 41954 259614 42574 295058
rect 41954 259058 41986 259614
rect 42542 259058 42574 259614
rect 41954 223614 42574 259058
rect 41954 223058 41986 223614
rect 42542 223058 42574 223614
rect 41954 187614 42574 223058
rect 41954 187058 41986 187614
rect 42542 187058 42574 187614
rect 41954 151614 42574 187058
rect 41954 151058 41986 151614
rect 42542 151058 42574 151614
rect 41954 115614 42574 151058
rect 41954 115058 41986 115614
rect 42542 115058 42574 115614
rect 41954 79614 42574 115058
rect 41954 79058 41986 79614
rect 42542 79058 42574 79614
rect 41954 43614 42574 79058
rect 41954 43058 41986 43614
rect 42542 43058 42574 43614
rect 41954 7614 42574 43058
rect 41954 7058 41986 7614
rect 42542 7058 42574 7614
rect 41954 -4186 42574 7058
rect 41954 -4742 41986 -4186
rect 42542 -4742 42574 -4186
rect 41954 -7654 42574 -4742
rect 43194 709638 43814 711590
rect 43194 709082 43226 709638
rect 43782 709082 43814 709638
rect 43194 692854 43814 709082
rect 43194 692298 43226 692854
rect 43782 692298 43814 692854
rect 43194 656854 43814 692298
rect 43194 656298 43226 656854
rect 43782 656298 43814 656854
rect 43194 620854 43814 656298
rect 43194 620298 43226 620854
rect 43782 620298 43814 620854
rect 43194 584854 43814 620298
rect 43194 584298 43226 584854
rect 43782 584298 43814 584854
rect 43194 548854 43814 584298
rect 43194 548298 43226 548854
rect 43782 548298 43814 548854
rect 43194 512854 43814 548298
rect 43194 512298 43226 512854
rect 43782 512298 43814 512854
rect 43194 476854 43814 512298
rect 43194 476298 43226 476854
rect 43782 476298 43814 476854
rect 43194 440854 43814 476298
rect 43194 440298 43226 440854
rect 43782 440298 43814 440854
rect 43194 404854 43814 440298
rect 43194 404298 43226 404854
rect 43782 404298 43814 404854
rect 43194 368854 43814 404298
rect 43194 368298 43226 368854
rect 43782 368298 43814 368854
rect 43194 332854 43814 368298
rect 43194 332298 43226 332854
rect 43782 332298 43814 332854
rect 43194 296854 43814 332298
rect 43194 296298 43226 296854
rect 43782 296298 43814 296854
rect 43194 260854 43814 296298
rect 43194 260298 43226 260854
rect 43782 260298 43814 260854
rect 43194 224854 43814 260298
rect 43194 224298 43226 224854
rect 43782 224298 43814 224854
rect 43194 188854 43814 224298
rect 43194 188298 43226 188854
rect 43782 188298 43814 188854
rect 43194 152854 43814 188298
rect 43194 152298 43226 152854
rect 43782 152298 43814 152854
rect 43194 116854 43814 152298
rect 43194 116298 43226 116854
rect 43782 116298 43814 116854
rect 43194 80854 43814 116298
rect 43194 80298 43226 80854
rect 43782 80298 43814 80854
rect 43194 44854 43814 80298
rect 43194 44298 43226 44854
rect 43782 44298 43814 44854
rect 43194 8854 43814 44298
rect 43194 8298 43226 8854
rect 43782 8298 43814 8854
rect 43194 -5146 43814 8298
rect 43194 -5702 43226 -5146
rect 43782 -5702 43814 -5146
rect 43194 -7654 43814 -5702
rect 44434 710598 45054 711590
rect 44434 710042 44466 710598
rect 45022 710042 45054 710598
rect 44434 694094 45054 710042
rect 44434 693538 44466 694094
rect 45022 693538 45054 694094
rect 44434 658094 45054 693538
rect 44434 657538 44466 658094
rect 45022 657538 45054 658094
rect 44434 622094 45054 657538
rect 44434 621538 44466 622094
rect 45022 621538 45054 622094
rect 44434 586094 45054 621538
rect 44434 585538 44466 586094
rect 45022 585538 45054 586094
rect 44434 550094 45054 585538
rect 44434 549538 44466 550094
rect 45022 549538 45054 550094
rect 44434 514094 45054 549538
rect 44434 513538 44466 514094
rect 45022 513538 45054 514094
rect 44434 478094 45054 513538
rect 44434 477538 44466 478094
rect 45022 477538 45054 478094
rect 44434 442094 45054 477538
rect 44434 441538 44466 442094
rect 45022 441538 45054 442094
rect 44434 406094 45054 441538
rect 44434 405538 44466 406094
rect 45022 405538 45054 406094
rect 44434 370094 45054 405538
rect 44434 369538 44466 370094
rect 45022 369538 45054 370094
rect 44434 334094 45054 369538
rect 44434 333538 44466 334094
rect 45022 333538 45054 334094
rect 44434 298094 45054 333538
rect 44434 297538 44466 298094
rect 45022 297538 45054 298094
rect 44434 262094 45054 297538
rect 44434 261538 44466 262094
rect 45022 261538 45054 262094
rect 44434 226094 45054 261538
rect 44434 225538 44466 226094
rect 45022 225538 45054 226094
rect 44434 190094 45054 225538
rect 44434 189538 44466 190094
rect 45022 189538 45054 190094
rect 44434 154094 45054 189538
rect 44434 153538 44466 154094
rect 45022 153538 45054 154094
rect 44434 118094 45054 153538
rect 44434 117538 44466 118094
rect 45022 117538 45054 118094
rect 44434 82094 45054 117538
rect 44434 81538 44466 82094
rect 45022 81538 45054 82094
rect 44434 46094 45054 81538
rect 44434 45538 44466 46094
rect 45022 45538 45054 46094
rect 44434 10094 45054 45538
rect 44434 9538 44466 10094
rect 45022 9538 45054 10094
rect 44434 -6106 45054 9538
rect 44434 -6662 44466 -6106
rect 45022 -6662 45054 -6106
rect 44434 -7654 45054 -6662
rect 45674 711558 46294 711590
rect 45674 711002 45706 711558
rect 46262 711002 46294 711558
rect 45674 695334 46294 711002
rect 45674 694778 45706 695334
rect 46262 694778 46294 695334
rect 45674 659334 46294 694778
rect 45674 658778 45706 659334
rect 46262 658778 46294 659334
rect 45674 623334 46294 658778
rect 45674 622778 45706 623334
rect 46262 622778 46294 623334
rect 45674 587334 46294 622778
rect 45674 586778 45706 587334
rect 46262 586778 46294 587334
rect 45674 551334 46294 586778
rect 45674 550778 45706 551334
rect 46262 550778 46294 551334
rect 45674 515334 46294 550778
rect 45674 514778 45706 515334
rect 46262 514778 46294 515334
rect 45674 479334 46294 514778
rect 45674 478778 45706 479334
rect 46262 478778 46294 479334
rect 45674 443334 46294 478778
rect 45674 442778 45706 443334
rect 46262 442778 46294 443334
rect 45674 407334 46294 442778
rect 45674 406778 45706 407334
rect 46262 406778 46294 407334
rect 45674 371334 46294 406778
rect 45674 370778 45706 371334
rect 46262 370778 46294 371334
rect 45674 335334 46294 370778
rect 45674 334778 45706 335334
rect 46262 334778 46294 335334
rect 45674 299334 46294 334778
rect 45674 298778 45706 299334
rect 46262 298778 46294 299334
rect 45674 263334 46294 298778
rect 45674 262778 45706 263334
rect 46262 262778 46294 263334
rect 45674 227334 46294 262778
rect 45674 226778 45706 227334
rect 46262 226778 46294 227334
rect 45674 191334 46294 226778
rect 45674 190778 45706 191334
rect 46262 190778 46294 191334
rect 45674 155334 46294 190778
rect 45674 154778 45706 155334
rect 46262 154778 46294 155334
rect 45674 119334 46294 154778
rect 45674 118778 45706 119334
rect 46262 118778 46294 119334
rect 45674 83334 46294 118778
rect 45674 82778 45706 83334
rect 46262 82778 46294 83334
rect 45674 47334 46294 82778
rect 45674 46778 45706 47334
rect 46262 46778 46294 47334
rect 45674 11334 46294 46778
rect 45674 10778 45706 11334
rect 46262 10778 46294 11334
rect 45674 -7066 46294 10778
rect 45674 -7622 45706 -7066
rect 46262 -7622 46294 -7066
rect 45674 -7654 46294 -7622
rect 72994 704838 73614 711590
rect 72994 704282 73026 704838
rect 73582 704282 73614 704838
rect 72994 686654 73614 704282
rect 72994 686098 73026 686654
rect 73582 686098 73614 686654
rect 72994 650654 73614 686098
rect 72994 650098 73026 650654
rect 73582 650098 73614 650654
rect 72994 614654 73614 650098
rect 72994 614098 73026 614654
rect 73582 614098 73614 614654
rect 72994 578654 73614 614098
rect 72994 578098 73026 578654
rect 73582 578098 73614 578654
rect 72994 542654 73614 578098
rect 72994 542098 73026 542654
rect 73582 542098 73614 542654
rect 72994 506654 73614 542098
rect 72994 506098 73026 506654
rect 73582 506098 73614 506654
rect 72994 470654 73614 506098
rect 72994 470098 73026 470654
rect 73582 470098 73614 470654
rect 72994 434654 73614 470098
rect 72994 434098 73026 434654
rect 73582 434098 73614 434654
rect 72994 398654 73614 434098
rect 72994 398098 73026 398654
rect 73582 398098 73614 398654
rect 72994 362654 73614 398098
rect 72994 362098 73026 362654
rect 73582 362098 73614 362654
rect 72994 326654 73614 362098
rect 72994 326098 73026 326654
rect 73582 326098 73614 326654
rect 72994 290654 73614 326098
rect 72994 290098 73026 290654
rect 73582 290098 73614 290654
rect 72994 254654 73614 290098
rect 72994 254098 73026 254654
rect 73582 254098 73614 254654
rect 72994 218654 73614 254098
rect 72994 218098 73026 218654
rect 73582 218098 73614 218654
rect 72994 182654 73614 218098
rect 72994 182098 73026 182654
rect 73582 182098 73614 182654
rect 72994 146654 73614 182098
rect 72994 146098 73026 146654
rect 73582 146098 73614 146654
rect 72994 110654 73614 146098
rect 72994 110098 73026 110654
rect 73582 110098 73614 110654
rect 72994 74654 73614 110098
rect 72994 74098 73026 74654
rect 73582 74098 73614 74654
rect 72994 38654 73614 74098
rect 72994 38098 73026 38654
rect 73582 38098 73614 38654
rect 72994 2654 73614 38098
rect 72994 2098 73026 2654
rect 73582 2098 73614 2654
rect 72994 -346 73614 2098
rect 72994 -902 73026 -346
rect 73582 -902 73614 -346
rect 72994 -7654 73614 -902
rect 74234 705798 74854 711590
rect 74234 705242 74266 705798
rect 74822 705242 74854 705798
rect 74234 687894 74854 705242
rect 74234 687338 74266 687894
rect 74822 687338 74854 687894
rect 74234 651894 74854 687338
rect 74234 651338 74266 651894
rect 74822 651338 74854 651894
rect 74234 615894 74854 651338
rect 74234 615338 74266 615894
rect 74822 615338 74854 615894
rect 74234 579894 74854 615338
rect 74234 579338 74266 579894
rect 74822 579338 74854 579894
rect 74234 543894 74854 579338
rect 74234 543338 74266 543894
rect 74822 543338 74854 543894
rect 74234 507894 74854 543338
rect 74234 507338 74266 507894
rect 74822 507338 74854 507894
rect 74234 471894 74854 507338
rect 74234 471338 74266 471894
rect 74822 471338 74854 471894
rect 74234 435894 74854 471338
rect 74234 435338 74266 435894
rect 74822 435338 74854 435894
rect 74234 399894 74854 435338
rect 74234 399338 74266 399894
rect 74822 399338 74854 399894
rect 74234 363894 74854 399338
rect 74234 363338 74266 363894
rect 74822 363338 74854 363894
rect 74234 327894 74854 363338
rect 74234 327338 74266 327894
rect 74822 327338 74854 327894
rect 74234 291894 74854 327338
rect 74234 291338 74266 291894
rect 74822 291338 74854 291894
rect 74234 255894 74854 291338
rect 74234 255338 74266 255894
rect 74822 255338 74854 255894
rect 74234 219894 74854 255338
rect 74234 219338 74266 219894
rect 74822 219338 74854 219894
rect 74234 183894 74854 219338
rect 74234 183338 74266 183894
rect 74822 183338 74854 183894
rect 74234 147894 74854 183338
rect 74234 147338 74266 147894
rect 74822 147338 74854 147894
rect 74234 111894 74854 147338
rect 74234 111338 74266 111894
rect 74822 111338 74854 111894
rect 74234 75894 74854 111338
rect 74234 75338 74266 75894
rect 74822 75338 74854 75894
rect 74234 39894 74854 75338
rect 74234 39338 74266 39894
rect 74822 39338 74854 39894
rect 74234 3894 74854 39338
rect 74234 3338 74266 3894
rect 74822 3338 74854 3894
rect 74234 -1306 74854 3338
rect 74234 -1862 74266 -1306
rect 74822 -1862 74854 -1306
rect 74234 -7654 74854 -1862
rect 75474 706758 76094 711590
rect 75474 706202 75506 706758
rect 76062 706202 76094 706758
rect 75474 689134 76094 706202
rect 75474 688578 75506 689134
rect 76062 688578 76094 689134
rect 75474 653134 76094 688578
rect 75474 652578 75506 653134
rect 76062 652578 76094 653134
rect 75474 617134 76094 652578
rect 75474 616578 75506 617134
rect 76062 616578 76094 617134
rect 75474 581134 76094 616578
rect 75474 580578 75506 581134
rect 76062 580578 76094 581134
rect 75474 545134 76094 580578
rect 75474 544578 75506 545134
rect 76062 544578 76094 545134
rect 75474 509134 76094 544578
rect 75474 508578 75506 509134
rect 76062 508578 76094 509134
rect 75474 473134 76094 508578
rect 75474 472578 75506 473134
rect 76062 472578 76094 473134
rect 75474 437134 76094 472578
rect 75474 436578 75506 437134
rect 76062 436578 76094 437134
rect 75474 401134 76094 436578
rect 75474 400578 75506 401134
rect 76062 400578 76094 401134
rect 75474 365134 76094 400578
rect 75474 364578 75506 365134
rect 76062 364578 76094 365134
rect 75474 329134 76094 364578
rect 75474 328578 75506 329134
rect 76062 328578 76094 329134
rect 75474 293134 76094 328578
rect 75474 292578 75506 293134
rect 76062 292578 76094 293134
rect 75474 257134 76094 292578
rect 75474 256578 75506 257134
rect 76062 256578 76094 257134
rect 75474 221134 76094 256578
rect 75474 220578 75506 221134
rect 76062 220578 76094 221134
rect 75474 185134 76094 220578
rect 75474 184578 75506 185134
rect 76062 184578 76094 185134
rect 75474 149134 76094 184578
rect 75474 148578 75506 149134
rect 76062 148578 76094 149134
rect 75474 113134 76094 148578
rect 75474 112578 75506 113134
rect 76062 112578 76094 113134
rect 75474 77134 76094 112578
rect 75474 76578 75506 77134
rect 76062 76578 76094 77134
rect 75474 41134 76094 76578
rect 75474 40578 75506 41134
rect 76062 40578 76094 41134
rect 75474 5134 76094 40578
rect 75474 4578 75506 5134
rect 76062 4578 76094 5134
rect 75474 -2266 76094 4578
rect 75474 -2822 75506 -2266
rect 76062 -2822 76094 -2266
rect 75474 -7654 76094 -2822
rect 76714 707718 77334 711590
rect 76714 707162 76746 707718
rect 77302 707162 77334 707718
rect 76714 690374 77334 707162
rect 76714 689818 76746 690374
rect 77302 689818 77334 690374
rect 76714 654374 77334 689818
rect 76714 653818 76746 654374
rect 77302 653818 77334 654374
rect 76714 618374 77334 653818
rect 76714 617818 76746 618374
rect 77302 617818 77334 618374
rect 76714 582374 77334 617818
rect 76714 581818 76746 582374
rect 77302 581818 77334 582374
rect 76714 546374 77334 581818
rect 76714 545818 76746 546374
rect 77302 545818 77334 546374
rect 76714 510374 77334 545818
rect 76714 509818 76746 510374
rect 77302 509818 77334 510374
rect 76714 474374 77334 509818
rect 76714 473818 76746 474374
rect 77302 473818 77334 474374
rect 76714 438374 77334 473818
rect 76714 437818 76746 438374
rect 77302 437818 77334 438374
rect 76714 402374 77334 437818
rect 76714 401818 76746 402374
rect 77302 401818 77334 402374
rect 76714 366374 77334 401818
rect 76714 365818 76746 366374
rect 77302 365818 77334 366374
rect 76714 330374 77334 365818
rect 76714 329818 76746 330374
rect 77302 329818 77334 330374
rect 76714 294374 77334 329818
rect 76714 293818 76746 294374
rect 77302 293818 77334 294374
rect 76714 258374 77334 293818
rect 76714 257818 76746 258374
rect 77302 257818 77334 258374
rect 76714 222374 77334 257818
rect 76714 221818 76746 222374
rect 77302 221818 77334 222374
rect 76714 186374 77334 221818
rect 76714 185818 76746 186374
rect 77302 185818 77334 186374
rect 76714 150374 77334 185818
rect 76714 149818 76746 150374
rect 77302 149818 77334 150374
rect 76714 114374 77334 149818
rect 76714 113818 76746 114374
rect 77302 113818 77334 114374
rect 76714 78374 77334 113818
rect 76714 77818 76746 78374
rect 77302 77818 77334 78374
rect 76714 42374 77334 77818
rect 76714 41818 76746 42374
rect 77302 41818 77334 42374
rect 76714 6374 77334 41818
rect 76714 5818 76746 6374
rect 77302 5818 77334 6374
rect 76714 -3226 77334 5818
rect 76714 -3782 76746 -3226
rect 77302 -3782 77334 -3226
rect 76714 -7654 77334 -3782
rect 77954 708678 78574 711590
rect 77954 708122 77986 708678
rect 78542 708122 78574 708678
rect 77954 691614 78574 708122
rect 77954 691058 77986 691614
rect 78542 691058 78574 691614
rect 77954 655614 78574 691058
rect 77954 655058 77986 655614
rect 78542 655058 78574 655614
rect 77954 619614 78574 655058
rect 77954 619058 77986 619614
rect 78542 619058 78574 619614
rect 77954 583614 78574 619058
rect 77954 583058 77986 583614
rect 78542 583058 78574 583614
rect 77954 547614 78574 583058
rect 77954 547058 77986 547614
rect 78542 547058 78574 547614
rect 77954 511614 78574 547058
rect 77954 511058 77986 511614
rect 78542 511058 78574 511614
rect 77954 475614 78574 511058
rect 77954 475058 77986 475614
rect 78542 475058 78574 475614
rect 77954 439614 78574 475058
rect 77954 439058 77986 439614
rect 78542 439058 78574 439614
rect 77954 403614 78574 439058
rect 77954 403058 77986 403614
rect 78542 403058 78574 403614
rect 77954 367614 78574 403058
rect 77954 367058 77986 367614
rect 78542 367058 78574 367614
rect 77954 331614 78574 367058
rect 77954 331058 77986 331614
rect 78542 331058 78574 331614
rect 77954 295614 78574 331058
rect 77954 295058 77986 295614
rect 78542 295058 78574 295614
rect 77954 259614 78574 295058
rect 77954 259058 77986 259614
rect 78542 259058 78574 259614
rect 77954 223614 78574 259058
rect 77954 223058 77986 223614
rect 78542 223058 78574 223614
rect 77954 187614 78574 223058
rect 77954 187058 77986 187614
rect 78542 187058 78574 187614
rect 77954 151614 78574 187058
rect 77954 151058 77986 151614
rect 78542 151058 78574 151614
rect 77954 115614 78574 151058
rect 77954 115058 77986 115614
rect 78542 115058 78574 115614
rect 77954 79614 78574 115058
rect 77954 79058 77986 79614
rect 78542 79058 78574 79614
rect 77954 43614 78574 79058
rect 77954 43058 77986 43614
rect 78542 43058 78574 43614
rect 77954 7614 78574 43058
rect 77954 7058 77986 7614
rect 78542 7058 78574 7614
rect 77954 -4186 78574 7058
rect 77954 -4742 77986 -4186
rect 78542 -4742 78574 -4186
rect 77954 -7654 78574 -4742
rect 79194 709638 79814 711590
rect 79194 709082 79226 709638
rect 79782 709082 79814 709638
rect 79194 692854 79814 709082
rect 79194 692298 79226 692854
rect 79782 692298 79814 692854
rect 79194 656854 79814 692298
rect 79194 656298 79226 656854
rect 79782 656298 79814 656854
rect 79194 620854 79814 656298
rect 79194 620298 79226 620854
rect 79782 620298 79814 620854
rect 79194 584854 79814 620298
rect 79194 584298 79226 584854
rect 79782 584298 79814 584854
rect 79194 548854 79814 584298
rect 79194 548298 79226 548854
rect 79782 548298 79814 548854
rect 79194 512854 79814 548298
rect 79194 512298 79226 512854
rect 79782 512298 79814 512854
rect 79194 476854 79814 512298
rect 79194 476298 79226 476854
rect 79782 476298 79814 476854
rect 79194 440854 79814 476298
rect 79194 440298 79226 440854
rect 79782 440298 79814 440854
rect 79194 404854 79814 440298
rect 79194 404298 79226 404854
rect 79782 404298 79814 404854
rect 79194 368854 79814 404298
rect 79194 368298 79226 368854
rect 79782 368298 79814 368854
rect 79194 332854 79814 368298
rect 79194 332298 79226 332854
rect 79782 332298 79814 332854
rect 79194 296854 79814 332298
rect 79194 296298 79226 296854
rect 79782 296298 79814 296854
rect 79194 260854 79814 296298
rect 79194 260298 79226 260854
rect 79782 260298 79814 260854
rect 79194 224854 79814 260298
rect 79194 224298 79226 224854
rect 79782 224298 79814 224854
rect 79194 188854 79814 224298
rect 79194 188298 79226 188854
rect 79782 188298 79814 188854
rect 79194 152854 79814 188298
rect 79194 152298 79226 152854
rect 79782 152298 79814 152854
rect 79194 116854 79814 152298
rect 79194 116298 79226 116854
rect 79782 116298 79814 116854
rect 79194 80854 79814 116298
rect 79194 80298 79226 80854
rect 79782 80298 79814 80854
rect 79194 44854 79814 80298
rect 79194 44298 79226 44854
rect 79782 44298 79814 44854
rect 79194 8854 79814 44298
rect 79194 8298 79226 8854
rect 79782 8298 79814 8854
rect 79194 -5146 79814 8298
rect 79194 -5702 79226 -5146
rect 79782 -5702 79814 -5146
rect 79194 -7654 79814 -5702
rect 80434 710598 81054 711590
rect 80434 710042 80466 710598
rect 81022 710042 81054 710598
rect 80434 694094 81054 710042
rect 80434 693538 80466 694094
rect 81022 693538 81054 694094
rect 80434 658094 81054 693538
rect 80434 657538 80466 658094
rect 81022 657538 81054 658094
rect 80434 622094 81054 657538
rect 80434 621538 80466 622094
rect 81022 621538 81054 622094
rect 80434 586094 81054 621538
rect 80434 585538 80466 586094
rect 81022 585538 81054 586094
rect 80434 550094 81054 585538
rect 80434 549538 80466 550094
rect 81022 549538 81054 550094
rect 80434 514094 81054 549538
rect 80434 513538 80466 514094
rect 81022 513538 81054 514094
rect 80434 478094 81054 513538
rect 80434 477538 80466 478094
rect 81022 477538 81054 478094
rect 80434 442094 81054 477538
rect 80434 441538 80466 442094
rect 81022 441538 81054 442094
rect 80434 406094 81054 441538
rect 80434 405538 80466 406094
rect 81022 405538 81054 406094
rect 80434 370094 81054 405538
rect 80434 369538 80466 370094
rect 81022 369538 81054 370094
rect 80434 334094 81054 369538
rect 80434 333538 80466 334094
rect 81022 333538 81054 334094
rect 80434 298094 81054 333538
rect 80434 297538 80466 298094
rect 81022 297538 81054 298094
rect 80434 262094 81054 297538
rect 80434 261538 80466 262094
rect 81022 261538 81054 262094
rect 80434 226094 81054 261538
rect 80434 225538 80466 226094
rect 81022 225538 81054 226094
rect 80434 190094 81054 225538
rect 80434 189538 80466 190094
rect 81022 189538 81054 190094
rect 80434 154094 81054 189538
rect 80434 153538 80466 154094
rect 81022 153538 81054 154094
rect 80434 118094 81054 153538
rect 80434 117538 80466 118094
rect 81022 117538 81054 118094
rect 80434 82094 81054 117538
rect 80434 81538 80466 82094
rect 81022 81538 81054 82094
rect 80434 46094 81054 81538
rect 80434 45538 80466 46094
rect 81022 45538 81054 46094
rect 80434 10094 81054 45538
rect 80434 9538 80466 10094
rect 81022 9538 81054 10094
rect 80434 -6106 81054 9538
rect 80434 -6662 80466 -6106
rect 81022 -6662 81054 -6106
rect 80434 -7654 81054 -6662
rect 81674 711558 82294 711590
rect 81674 711002 81706 711558
rect 82262 711002 82294 711558
rect 81674 695334 82294 711002
rect 81674 694778 81706 695334
rect 82262 694778 82294 695334
rect 81674 659334 82294 694778
rect 81674 658778 81706 659334
rect 82262 658778 82294 659334
rect 81674 623334 82294 658778
rect 81674 622778 81706 623334
rect 82262 622778 82294 623334
rect 81674 587334 82294 622778
rect 81674 586778 81706 587334
rect 82262 586778 82294 587334
rect 81674 551334 82294 586778
rect 81674 550778 81706 551334
rect 82262 550778 82294 551334
rect 81674 515334 82294 550778
rect 81674 514778 81706 515334
rect 82262 514778 82294 515334
rect 81674 479334 82294 514778
rect 81674 478778 81706 479334
rect 82262 478778 82294 479334
rect 81674 443334 82294 478778
rect 81674 442778 81706 443334
rect 82262 442778 82294 443334
rect 81674 407334 82294 442778
rect 81674 406778 81706 407334
rect 82262 406778 82294 407334
rect 81674 371334 82294 406778
rect 81674 370778 81706 371334
rect 82262 370778 82294 371334
rect 81674 335334 82294 370778
rect 81674 334778 81706 335334
rect 82262 334778 82294 335334
rect 81674 299334 82294 334778
rect 81674 298778 81706 299334
rect 82262 298778 82294 299334
rect 81674 263334 82294 298778
rect 81674 262778 81706 263334
rect 82262 262778 82294 263334
rect 81674 227334 82294 262778
rect 81674 226778 81706 227334
rect 82262 226778 82294 227334
rect 81674 191334 82294 226778
rect 81674 190778 81706 191334
rect 82262 190778 82294 191334
rect 81674 155334 82294 190778
rect 81674 154778 81706 155334
rect 82262 154778 82294 155334
rect 81674 119334 82294 154778
rect 81674 118778 81706 119334
rect 82262 118778 82294 119334
rect 81674 83334 82294 118778
rect 81674 82778 81706 83334
rect 82262 82778 82294 83334
rect 81674 47334 82294 82778
rect 81674 46778 81706 47334
rect 82262 46778 82294 47334
rect 81674 11334 82294 46778
rect 81674 10778 81706 11334
rect 82262 10778 82294 11334
rect 81674 -7066 82294 10778
rect 81674 -7622 81706 -7066
rect 82262 -7622 82294 -7066
rect 81674 -7654 82294 -7622
rect 108994 704838 109614 711590
rect 108994 704282 109026 704838
rect 109582 704282 109614 704838
rect 108994 686654 109614 704282
rect 108994 686098 109026 686654
rect 109582 686098 109614 686654
rect 108994 650654 109614 686098
rect 108994 650098 109026 650654
rect 109582 650098 109614 650654
rect 108994 614654 109614 650098
rect 108994 614098 109026 614654
rect 109582 614098 109614 614654
rect 108994 578654 109614 614098
rect 108994 578098 109026 578654
rect 109582 578098 109614 578654
rect 108994 542654 109614 578098
rect 108994 542098 109026 542654
rect 109582 542098 109614 542654
rect 108994 506654 109614 542098
rect 108994 506098 109026 506654
rect 109582 506098 109614 506654
rect 108994 470654 109614 506098
rect 108994 470098 109026 470654
rect 109582 470098 109614 470654
rect 108994 434654 109614 470098
rect 108994 434098 109026 434654
rect 109582 434098 109614 434654
rect 108994 398654 109614 434098
rect 108994 398098 109026 398654
rect 109582 398098 109614 398654
rect 108994 362654 109614 398098
rect 108994 362098 109026 362654
rect 109582 362098 109614 362654
rect 108994 326654 109614 362098
rect 108994 326098 109026 326654
rect 109582 326098 109614 326654
rect 108994 290654 109614 326098
rect 108994 290098 109026 290654
rect 109582 290098 109614 290654
rect 108994 254654 109614 290098
rect 108994 254098 109026 254654
rect 109582 254098 109614 254654
rect 108994 218654 109614 254098
rect 108994 218098 109026 218654
rect 109582 218098 109614 218654
rect 108994 182654 109614 218098
rect 108994 182098 109026 182654
rect 109582 182098 109614 182654
rect 108994 146654 109614 182098
rect 108994 146098 109026 146654
rect 109582 146098 109614 146654
rect 108994 110654 109614 146098
rect 108994 110098 109026 110654
rect 109582 110098 109614 110654
rect 108994 74654 109614 110098
rect 108994 74098 109026 74654
rect 109582 74098 109614 74654
rect 108994 38654 109614 74098
rect 108994 38098 109026 38654
rect 109582 38098 109614 38654
rect 108994 2654 109614 38098
rect 108994 2098 109026 2654
rect 109582 2098 109614 2654
rect 108994 -346 109614 2098
rect 108994 -902 109026 -346
rect 109582 -902 109614 -346
rect 108994 -7654 109614 -902
rect 110234 705798 110854 711590
rect 110234 705242 110266 705798
rect 110822 705242 110854 705798
rect 110234 687894 110854 705242
rect 110234 687338 110266 687894
rect 110822 687338 110854 687894
rect 110234 651894 110854 687338
rect 110234 651338 110266 651894
rect 110822 651338 110854 651894
rect 110234 615894 110854 651338
rect 110234 615338 110266 615894
rect 110822 615338 110854 615894
rect 110234 579894 110854 615338
rect 110234 579338 110266 579894
rect 110822 579338 110854 579894
rect 110234 543894 110854 579338
rect 110234 543338 110266 543894
rect 110822 543338 110854 543894
rect 110234 507894 110854 543338
rect 110234 507338 110266 507894
rect 110822 507338 110854 507894
rect 110234 471894 110854 507338
rect 110234 471338 110266 471894
rect 110822 471338 110854 471894
rect 110234 435894 110854 471338
rect 110234 435338 110266 435894
rect 110822 435338 110854 435894
rect 110234 399894 110854 435338
rect 110234 399338 110266 399894
rect 110822 399338 110854 399894
rect 110234 363894 110854 399338
rect 110234 363338 110266 363894
rect 110822 363338 110854 363894
rect 110234 327894 110854 363338
rect 110234 327338 110266 327894
rect 110822 327338 110854 327894
rect 110234 291894 110854 327338
rect 110234 291338 110266 291894
rect 110822 291338 110854 291894
rect 110234 255894 110854 291338
rect 110234 255338 110266 255894
rect 110822 255338 110854 255894
rect 110234 219894 110854 255338
rect 110234 219338 110266 219894
rect 110822 219338 110854 219894
rect 110234 183894 110854 219338
rect 110234 183338 110266 183894
rect 110822 183338 110854 183894
rect 110234 147894 110854 183338
rect 110234 147338 110266 147894
rect 110822 147338 110854 147894
rect 110234 111894 110854 147338
rect 110234 111338 110266 111894
rect 110822 111338 110854 111894
rect 110234 75894 110854 111338
rect 110234 75338 110266 75894
rect 110822 75338 110854 75894
rect 110234 39894 110854 75338
rect 110234 39338 110266 39894
rect 110822 39338 110854 39894
rect 110234 3894 110854 39338
rect 110234 3338 110266 3894
rect 110822 3338 110854 3894
rect 110234 -1306 110854 3338
rect 110234 -1862 110266 -1306
rect 110822 -1862 110854 -1306
rect 110234 -7654 110854 -1862
rect 111474 706758 112094 711590
rect 111474 706202 111506 706758
rect 112062 706202 112094 706758
rect 111474 689134 112094 706202
rect 111474 688578 111506 689134
rect 112062 688578 112094 689134
rect 111474 653134 112094 688578
rect 111474 652578 111506 653134
rect 112062 652578 112094 653134
rect 111474 617134 112094 652578
rect 111474 616578 111506 617134
rect 112062 616578 112094 617134
rect 111474 581134 112094 616578
rect 111474 580578 111506 581134
rect 112062 580578 112094 581134
rect 111474 545134 112094 580578
rect 111474 544578 111506 545134
rect 112062 544578 112094 545134
rect 111474 509134 112094 544578
rect 111474 508578 111506 509134
rect 112062 508578 112094 509134
rect 111474 473134 112094 508578
rect 111474 472578 111506 473134
rect 112062 472578 112094 473134
rect 111474 437134 112094 472578
rect 111474 436578 111506 437134
rect 112062 436578 112094 437134
rect 111474 401134 112094 436578
rect 111474 400578 111506 401134
rect 112062 400578 112094 401134
rect 111474 365134 112094 400578
rect 111474 364578 111506 365134
rect 112062 364578 112094 365134
rect 111474 329134 112094 364578
rect 111474 328578 111506 329134
rect 112062 328578 112094 329134
rect 111474 293134 112094 328578
rect 111474 292578 111506 293134
rect 112062 292578 112094 293134
rect 111474 257134 112094 292578
rect 111474 256578 111506 257134
rect 112062 256578 112094 257134
rect 111474 221134 112094 256578
rect 111474 220578 111506 221134
rect 112062 220578 112094 221134
rect 111474 185134 112094 220578
rect 111474 184578 111506 185134
rect 112062 184578 112094 185134
rect 111474 149134 112094 184578
rect 111474 148578 111506 149134
rect 112062 148578 112094 149134
rect 111474 113134 112094 148578
rect 111474 112578 111506 113134
rect 112062 112578 112094 113134
rect 111474 77134 112094 112578
rect 111474 76578 111506 77134
rect 112062 76578 112094 77134
rect 111474 41134 112094 76578
rect 111474 40578 111506 41134
rect 112062 40578 112094 41134
rect 111474 5134 112094 40578
rect 111474 4578 111506 5134
rect 112062 4578 112094 5134
rect 111474 -2266 112094 4578
rect 111474 -2822 111506 -2266
rect 112062 -2822 112094 -2266
rect 111474 -7654 112094 -2822
rect 112714 707718 113334 711590
rect 112714 707162 112746 707718
rect 113302 707162 113334 707718
rect 112714 690374 113334 707162
rect 112714 689818 112746 690374
rect 113302 689818 113334 690374
rect 112714 654374 113334 689818
rect 112714 653818 112746 654374
rect 113302 653818 113334 654374
rect 112714 618374 113334 653818
rect 112714 617818 112746 618374
rect 113302 617818 113334 618374
rect 112714 582374 113334 617818
rect 112714 581818 112746 582374
rect 113302 581818 113334 582374
rect 112714 546374 113334 581818
rect 112714 545818 112746 546374
rect 113302 545818 113334 546374
rect 112714 510374 113334 545818
rect 112714 509818 112746 510374
rect 113302 509818 113334 510374
rect 112714 474374 113334 509818
rect 112714 473818 112746 474374
rect 113302 473818 113334 474374
rect 112714 438374 113334 473818
rect 112714 437818 112746 438374
rect 113302 437818 113334 438374
rect 112714 402374 113334 437818
rect 112714 401818 112746 402374
rect 113302 401818 113334 402374
rect 112714 366374 113334 401818
rect 112714 365818 112746 366374
rect 113302 365818 113334 366374
rect 112714 330374 113334 365818
rect 112714 329818 112746 330374
rect 113302 329818 113334 330374
rect 112714 294374 113334 329818
rect 112714 293818 112746 294374
rect 113302 293818 113334 294374
rect 112714 258374 113334 293818
rect 112714 257818 112746 258374
rect 113302 257818 113334 258374
rect 112714 222374 113334 257818
rect 112714 221818 112746 222374
rect 113302 221818 113334 222374
rect 112714 186374 113334 221818
rect 112714 185818 112746 186374
rect 113302 185818 113334 186374
rect 112714 150374 113334 185818
rect 112714 149818 112746 150374
rect 113302 149818 113334 150374
rect 112714 114374 113334 149818
rect 112714 113818 112746 114374
rect 113302 113818 113334 114374
rect 112714 78374 113334 113818
rect 112714 77818 112746 78374
rect 113302 77818 113334 78374
rect 112714 42374 113334 77818
rect 112714 41818 112746 42374
rect 113302 41818 113334 42374
rect 112714 6374 113334 41818
rect 112714 5818 112746 6374
rect 113302 5818 113334 6374
rect 112714 -3226 113334 5818
rect 112714 -3782 112746 -3226
rect 113302 -3782 113334 -3226
rect 112714 -7654 113334 -3782
rect 113954 708678 114574 711590
rect 113954 708122 113986 708678
rect 114542 708122 114574 708678
rect 113954 691614 114574 708122
rect 113954 691058 113986 691614
rect 114542 691058 114574 691614
rect 113954 655614 114574 691058
rect 113954 655058 113986 655614
rect 114542 655058 114574 655614
rect 113954 619614 114574 655058
rect 113954 619058 113986 619614
rect 114542 619058 114574 619614
rect 113954 583614 114574 619058
rect 113954 583058 113986 583614
rect 114542 583058 114574 583614
rect 113954 547614 114574 583058
rect 113954 547058 113986 547614
rect 114542 547058 114574 547614
rect 113954 511614 114574 547058
rect 113954 511058 113986 511614
rect 114542 511058 114574 511614
rect 113954 475614 114574 511058
rect 113954 475058 113986 475614
rect 114542 475058 114574 475614
rect 113954 439614 114574 475058
rect 113954 439058 113986 439614
rect 114542 439058 114574 439614
rect 113954 403614 114574 439058
rect 113954 403058 113986 403614
rect 114542 403058 114574 403614
rect 113954 367614 114574 403058
rect 113954 367058 113986 367614
rect 114542 367058 114574 367614
rect 113954 331614 114574 367058
rect 113954 331058 113986 331614
rect 114542 331058 114574 331614
rect 113954 295614 114574 331058
rect 113954 295058 113986 295614
rect 114542 295058 114574 295614
rect 113954 259614 114574 295058
rect 113954 259058 113986 259614
rect 114542 259058 114574 259614
rect 113954 223614 114574 259058
rect 113954 223058 113986 223614
rect 114542 223058 114574 223614
rect 113954 187614 114574 223058
rect 113954 187058 113986 187614
rect 114542 187058 114574 187614
rect 113954 151614 114574 187058
rect 113954 151058 113986 151614
rect 114542 151058 114574 151614
rect 113954 115614 114574 151058
rect 113954 115058 113986 115614
rect 114542 115058 114574 115614
rect 113954 79614 114574 115058
rect 113954 79058 113986 79614
rect 114542 79058 114574 79614
rect 113954 43614 114574 79058
rect 113954 43058 113986 43614
rect 114542 43058 114574 43614
rect 113954 7614 114574 43058
rect 113954 7058 113986 7614
rect 114542 7058 114574 7614
rect 113954 -4186 114574 7058
rect 113954 -4742 113986 -4186
rect 114542 -4742 114574 -4186
rect 113954 -7654 114574 -4742
rect 115194 709638 115814 711590
rect 115194 709082 115226 709638
rect 115782 709082 115814 709638
rect 115194 692854 115814 709082
rect 115194 692298 115226 692854
rect 115782 692298 115814 692854
rect 115194 656854 115814 692298
rect 115194 656298 115226 656854
rect 115782 656298 115814 656854
rect 115194 620854 115814 656298
rect 115194 620298 115226 620854
rect 115782 620298 115814 620854
rect 115194 584854 115814 620298
rect 115194 584298 115226 584854
rect 115782 584298 115814 584854
rect 115194 548854 115814 584298
rect 115194 548298 115226 548854
rect 115782 548298 115814 548854
rect 115194 512854 115814 548298
rect 115194 512298 115226 512854
rect 115782 512298 115814 512854
rect 115194 476854 115814 512298
rect 115194 476298 115226 476854
rect 115782 476298 115814 476854
rect 115194 440854 115814 476298
rect 115194 440298 115226 440854
rect 115782 440298 115814 440854
rect 115194 404854 115814 440298
rect 115194 404298 115226 404854
rect 115782 404298 115814 404854
rect 115194 368854 115814 404298
rect 115194 368298 115226 368854
rect 115782 368298 115814 368854
rect 115194 332854 115814 368298
rect 115194 332298 115226 332854
rect 115782 332298 115814 332854
rect 115194 296854 115814 332298
rect 115194 296298 115226 296854
rect 115782 296298 115814 296854
rect 115194 260854 115814 296298
rect 115194 260298 115226 260854
rect 115782 260298 115814 260854
rect 115194 224854 115814 260298
rect 115194 224298 115226 224854
rect 115782 224298 115814 224854
rect 115194 188854 115814 224298
rect 115194 188298 115226 188854
rect 115782 188298 115814 188854
rect 115194 152854 115814 188298
rect 115194 152298 115226 152854
rect 115782 152298 115814 152854
rect 115194 116854 115814 152298
rect 115194 116298 115226 116854
rect 115782 116298 115814 116854
rect 115194 80854 115814 116298
rect 115194 80298 115226 80854
rect 115782 80298 115814 80854
rect 115194 44854 115814 80298
rect 115194 44298 115226 44854
rect 115782 44298 115814 44854
rect 115194 8854 115814 44298
rect 115194 8298 115226 8854
rect 115782 8298 115814 8854
rect 115194 -5146 115814 8298
rect 115194 -5702 115226 -5146
rect 115782 -5702 115814 -5146
rect 115194 -7654 115814 -5702
rect 116434 710598 117054 711590
rect 116434 710042 116466 710598
rect 117022 710042 117054 710598
rect 116434 694094 117054 710042
rect 116434 693538 116466 694094
rect 117022 693538 117054 694094
rect 116434 658094 117054 693538
rect 116434 657538 116466 658094
rect 117022 657538 117054 658094
rect 116434 622094 117054 657538
rect 116434 621538 116466 622094
rect 117022 621538 117054 622094
rect 116434 586094 117054 621538
rect 116434 585538 116466 586094
rect 117022 585538 117054 586094
rect 116434 550094 117054 585538
rect 116434 549538 116466 550094
rect 117022 549538 117054 550094
rect 116434 514094 117054 549538
rect 116434 513538 116466 514094
rect 117022 513538 117054 514094
rect 116434 478094 117054 513538
rect 116434 477538 116466 478094
rect 117022 477538 117054 478094
rect 116434 442094 117054 477538
rect 116434 441538 116466 442094
rect 117022 441538 117054 442094
rect 116434 406094 117054 441538
rect 116434 405538 116466 406094
rect 117022 405538 117054 406094
rect 116434 370094 117054 405538
rect 116434 369538 116466 370094
rect 117022 369538 117054 370094
rect 116434 334094 117054 369538
rect 116434 333538 116466 334094
rect 117022 333538 117054 334094
rect 116434 298094 117054 333538
rect 116434 297538 116466 298094
rect 117022 297538 117054 298094
rect 116434 262094 117054 297538
rect 116434 261538 116466 262094
rect 117022 261538 117054 262094
rect 116434 226094 117054 261538
rect 116434 225538 116466 226094
rect 117022 225538 117054 226094
rect 116434 190094 117054 225538
rect 116434 189538 116466 190094
rect 117022 189538 117054 190094
rect 116434 154094 117054 189538
rect 116434 153538 116466 154094
rect 117022 153538 117054 154094
rect 116434 118094 117054 153538
rect 116434 117538 116466 118094
rect 117022 117538 117054 118094
rect 116434 82094 117054 117538
rect 116434 81538 116466 82094
rect 117022 81538 117054 82094
rect 116434 46094 117054 81538
rect 116434 45538 116466 46094
rect 117022 45538 117054 46094
rect 116434 10094 117054 45538
rect 116434 9538 116466 10094
rect 117022 9538 117054 10094
rect 116434 -6106 117054 9538
rect 116434 -6662 116466 -6106
rect 117022 -6662 117054 -6106
rect 116434 -7654 117054 -6662
rect 117674 711558 118294 711590
rect 117674 711002 117706 711558
rect 118262 711002 118294 711558
rect 117674 695334 118294 711002
rect 117674 694778 117706 695334
rect 118262 694778 118294 695334
rect 117674 659334 118294 694778
rect 117674 658778 117706 659334
rect 118262 658778 118294 659334
rect 117674 623334 118294 658778
rect 117674 622778 117706 623334
rect 118262 622778 118294 623334
rect 117674 587334 118294 622778
rect 117674 586778 117706 587334
rect 118262 586778 118294 587334
rect 117674 551334 118294 586778
rect 117674 550778 117706 551334
rect 118262 550778 118294 551334
rect 117674 515334 118294 550778
rect 117674 514778 117706 515334
rect 118262 514778 118294 515334
rect 117674 479334 118294 514778
rect 117674 478778 117706 479334
rect 118262 478778 118294 479334
rect 117674 443334 118294 478778
rect 117674 442778 117706 443334
rect 118262 442778 118294 443334
rect 117674 407334 118294 442778
rect 117674 406778 117706 407334
rect 118262 406778 118294 407334
rect 117674 371334 118294 406778
rect 117674 370778 117706 371334
rect 118262 370778 118294 371334
rect 117674 335334 118294 370778
rect 117674 334778 117706 335334
rect 118262 334778 118294 335334
rect 117674 299334 118294 334778
rect 117674 298778 117706 299334
rect 118262 298778 118294 299334
rect 117674 263334 118294 298778
rect 117674 262778 117706 263334
rect 118262 262778 118294 263334
rect 117674 227334 118294 262778
rect 117674 226778 117706 227334
rect 118262 226778 118294 227334
rect 117674 191334 118294 226778
rect 117674 190778 117706 191334
rect 118262 190778 118294 191334
rect 117674 155334 118294 190778
rect 117674 154778 117706 155334
rect 118262 154778 118294 155334
rect 117674 119334 118294 154778
rect 117674 118778 117706 119334
rect 118262 118778 118294 119334
rect 117674 83334 118294 118778
rect 117674 82778 117706 83334
rect 118262 82778 118294 83334
rect 117674 47334 118294 82778
rect 117674 46778 117706 47334
rect 118262 46778 118294 47334
rect 117674 11334 118294 46778
rect 117674 10778 117706 11334
rect 118262 10778 118294 11334
rect 117674 -7066 118294 10778
rect 117674 -7622 117706 -7066
rect 118262 -7622 118294 -7066
rect 117674 -7654 118294 -7622
rect 144994 704838 145614 711590
rect 144994 704282 145026 704838
rect 145582 704282 145614 704838
rect 144994 686654 145614 704282
rect 144994 686098 145026 686654
rect 145582 686098 145614 686654
rect 144994 650654 145614 686098
rect 144994 650098 145026 650654
rect 145582 650098 145614 650654
rect 144994 614654 145614 650098
rect 144994 614098 145026 614654
rect 145582 614098 145614 614654
rect 144994 578654 145614 614098
rect 144994 578098 145026 578654
rect 145582 578098 145614 578654
rect 144994 542654 145614 578098
rect 144994 542098 145026 542654
rect 145582 542098 145614 542654
rect 144994 506654 145614 542098
rect 144994 506098 145026 506654
rect 145582 506098 145614 506654
rect 144994 470654 145614 506098
rect 144994 470098 145026 470654
rect 145582 470098 145614 470654
rect 144994 434654 145614 470098
rect 144994 434098 145026 434654
rect 145582 434098 145614 434654
rect 144994 398654 145614 434098
rect 144994 398098 145026 398654
rect 145582 398098 145614 398654
rect 144994 362654 145614 398098
rect 144994 362098 145026 362654
rect 145582 362098 145614 362654
rect 144994 326654 145614 362098
rect 144994 326098 145026 326654
rect 145582 326098 145614 326654
rect 144994 290654 145614 326098
rect 144994 290098 145026 290654
rect 145582 290098 145614 290654
rect 144994 254654 145614 290098
rect 144994 254098 145026 254654
rect 145582 254098 145614 254654
rect 144994 218654 145614 254098
rect 144994 218098 145026 218654
rect 145582 218098 145614 218654
rect 144994 182654 145614 218098
rect 144994 182098 145026 182654
rect 145582 182098 145614 182654
rect 144994 146654 145614 182098
rect 144994 146098 145026 146654
rect 145582 146098 145614 146654
rect 144994 110654 145614 146098
rect 144994 110098 145026 110654
rect 145582 110098 145614 110654
rect 144994 74654 145614 110098
rect 144994 74098 145026 74654
rect 145582 74098 145614 74654
rect 144994 38654 145614 74098
rect 144994 38098 145026 38654
rect 145582 38098 145614 38654
rect 144994 2654 145614 38098
rect 144994 2098 145026 2654
rect 145582 2098 145614 2654
rect 144994 -346 145614 2098
rect 144994 -902 145026 -346
rect 145582 -902 145614 -346
rect 144994 -7654 145614 -902
rect 146234 705798 146854 711590
rect 146234 705242 146266 705798
rect 146822 705242 146854 705798
rect 146234 687894 146854 705242
rect 146234 687338 146266 687894
rect 146822 687338 146854 687894
rect 146234 651894 146854 687338
rect 146234 651338 146266 651894
rect 146822 651338 146854 651894
rect 146234 615894 146854 651338
rect 146234 615338 146266 615894
rect 146822 615338 146854 615894
rect 146234 579894 146854 615338
rect 146234 579338 146266 579894
rect 146822 579338 146854 579894
rect 146234 543894 146854 579338
rect 146234 543338 146266 543894
rect 146822 543338 146854 543894
rect 146234 507894 146854 543338
rect 146234 507338 146266 507894
rect 146822 507338 146854 507894
rect 146234 471894 146854 507338
rect 146234 471338 146266 471894
rect 146822 471338 146854 471894
rect 146234 435894 146854 471338
rect 146234 435338 146266 435894
rect 146822 435338 146854 435894
rect 146234 399894 146854 435338
rect 146234 399338 146266 399894
rect 146822 399338 146854 399894
rect 146234 363894 146854 399338
rect 146234 363338 146266 363894
rect 146822 363338 146854 363894
rect 146234 327894 146854 363338
rect 146234 327338 146266 327894
rect 146822 327338 146854 327894
rect 146234 291894 146854 327338
rect 146234 291338 146266 291894
rect 146822 291338 146854 291894
rect 146234 255894 146854 291338
rect 146234 255338 146266 255894
rect 146822 255338 146854 255894
rect 146234 219894 146854 255338
rect 146234 219338 146266 219894
rect 146822 219338 146854 219894
rect 146234 183894 146854 219338
rect 146234 183338 146266 183894
rect 146822 183338 146854 183894
rect 146234 147894 146854 183338
rect 146234 147338 146266 147894
rect 146822 147338 146854 147894
rect 146234 111894 146854 147338
rect 146234 111338 146266 111894
rect 146822 111338 146854 111894
rect 146234 75894 146854 111338
rect 146234 75338 146266 75894
rect 146822 75338 146854 75894
rect 146234 39894 146854 75338
rect 146234 39338 146266 39894
rect 146822 39338 146854 39894
rect 146234 3894 146854 39338
rect 146234 3338 146266 3894
rect 146822 3338 146854 3894
rect 146234 -1306 146854 3338
rect 146234 -1862 146266 -1306
rect 146822 -1862 146854 -1306
rect 146234 -7654 146854 -1862
rect 147474 706758 148094 711590
rect 147474 706202 147506 706758
rect 148062 706202 148094 706758
rect 147474 689134 148094 706202
rect 147474 688578 147506 689134
rect 148062 688578 148094 689134
rect 147474 653134 148094 688578
rect 147474 652578 147506 653134
rect 148062 652578 148094 653134
rect 147474 617134 148094 652578
rect 147474 616578 147506 617134
rect 148062 616578 148094 617134
rect 147474 581134 148094 616578
rect 147474 580578 147506 581134
rect 148062 580578 148094 581134
rect 147474 545134 148094 580578
rect 147474 544578 147506 545134
rect 148062 544578 148094 545134
rect 147474 509134 148094 544578
rect 147474 508578 147506 509134
rect 148062 508578 148094 509134
rect 147474 473134 148094 508578
rect 147474 472578 147506 473134
rect 148062 472578 148094 473134
rect 147474 437134 148094 472578
rect 147474 436578 147506 437134
rect 148062 436578 148094 437134
rect 147474 401134 148094 436578
rect 147474 400578 147506 401134
rect 148062 400578 148094 401134
rect 147474 365134 148094 400578
rect 147474 364578 147506 365134
rect 148062 364578 148094 365134
rect 147474 329134 148094 364578
rect 147474 328578 147506 329134
rect 148062 328578 148094 329134
rect 147474 293134 148094 328578
rect 147474 292578 147506 293134
rect 148062 292578 148094 293134
rect 147474 257134 148094 292578
rect 147474 256578 147506 257134
rect 148062 256578 148094 257134
rect 147474 221134 148094 256578
rect 147474 220578 147506 221134
rect 148062 220578 148094 221134
rect 147474 185134 148094 220578
rect 147474 184578 147506 185134
rect 148062 184578 148094 185134
rect 147474 149134 148094 184578
rect 147474 148578 147506 149134
rect 148062 148578 148094 149134
rect 147474 113134 148094 148578
rect 147474 112578 147506 113134
rect 148062 112578 148094 113134
rect 147474 77134 148094 112578
rect 147474 76578 147506 77134
rect 148062 76578 148094 77134
rect 147474 41134 148094 76578
rect 147474 40578 147506 41134
rect 148062 40578 148094 41134
rect 147474 5134 148094 40578
rect 147474 4578 147506 5134
rect 148062 4578 148094 5134
rect 147474 -2266 148094 4578
rect 147474 -2822 147506 -2266
rect 148062 -2822 148094 -2266
rect 147474 -7654 148094 -2822
rect 148714 707718 149334 711590
rect 148714 707162 148746 707718
rect 149302 707162 149334 707718
rect 148714 690374 149334 707162
rect 148714 689818 148746 690374
rect 149302 689818 149334 690374
rect 148714 654374 149334 689818
rect 148714 653818 148746 654374
rect 149302 653818 149334 654374
rect 148714 618374 149334 653818
rect 148714 617818 148746 618374
rect 149302 617818 149334 618374
rect 148714 582374 149334 617818
rect 148714 581818 148746 582374
rect 149302 581818 149334 582374
rect 148714 546374 149334 581818
rect 148714 545818 148746 546374
rect 149302 545818 149334 546374
rect 148714 510374 149334 545818
rect 148714 509818 148746 510374
rect 149302 509818 149334 510374
rect 148714 474374 149334 509818
rect 148714 473818 148746 474374
rect 149302 473818 149334 474374
rect 148714 438374 149334 473818
rect 148714 437818 148746 438374
rect 149302 437818 149334 438374
rect 148714 402374 149334 437818
rect 148714 401818 148746 402374
rect 149302 401818 149334 402374
rect 148714 366374 149334 401818
rect 148714 365818 148746 366374
rect 149302 365818 149334 366374
rect 148714 330374 149334 365818
rect 148714 329818 148746 330374
rect 149302 329818 149334 330374
rect 148714 294374 149334 329818
rect 148714 293818 148746 294374
rect 149302 293818 149334 294374
rect 148714 258374 149334 293818
rect 148714 257818 148746 258374
rect 149302 257818 149334 258374
rect 148714 222374 149334 257818
rect 148714 221818 148746 222374
rect 149302 221818 149334 222374
rect 148714 186374 149334 221818
rect 148714 185818 148746 186374
rect 149302 185818 149334 186374
rect 148714 150374 149334 185818
rect 148714 149818 148746 150374
rect 149302 149818 149334 150374
rect 148714 114374 149334 149818
rect 148714 113818 148746 114374
rect 149302 113818 149334 114374
rect 148714 78374 149334 113818
rect 148714 77818 148746 78374
rect 149302 77818 149334 78374
rect 148714 42374 149334 77818
rect 148714 41818 148746 42374
rect 149302 41818 149334 42374
rect 148714 6374 149334 41818
rect 148714 5818 148746 6374
rect 149302 5818 149334 6374
rect 148714 -3226 149334 5818
rect 148714 -3782 148746 -3226
rect 149302 -3782 149334 -3226
rect 148714 -7654 149334 -3782
rect 149954 708678 150574 711590
rect 149954 708122 149986 708678
rect 150542 708122 150574 708678
rect 149954 691614 150574 708122
rect 149954 691058 149986 691614
rect 150542 691058 150574 691614
rect 149954 655614 150574 691058
rect 149954 655058 149986 655614
rect 150542 655058 150574 655614
rect 149954 619614 150574 655058
rect 149954 619058 149986 619614
rect 150542 619058 150574 619614
rect 149954 583614 150574 619058
rect 149954 583058 149986 583614
rect 150542 583058 150574 583614
rect 149954 547614 150574 583058
rect 149954 547058 149986 547614
rect 150542 547058 150574 547614
rect 149954 511614 150574 547058
rect 149954 511058 149986 511614
rect 150542 511058 150574 511614
rect 149954 475614 150574 511058
rect 149954 475058 149986 475614
rect 150542 475058 150574 475614
rect 149954 439614 150574 475058
rect 149954 439058 149986 439614
rect 150542 439058 150574 439614
rect 149954 403614 150574 439058
rect 149954 403058 149986 403614
rect 150542 403058 150574 403614
rect 149954 367614 150574 403058
rect 149954 367058 149986 367614
rect 150542 367058 150574 367614
rect 149954 331614 150574 367058
rect 149954 331058 149986 331614
rect 150542 331058 150574 331614
rect 149954 295614 150574 331058
rect 149954 295058 149986 295614
rect 150542 295058 150574 295614
rect 149954 259614 150574 295058
rect 149954 259058 149986 259614
rect 150542 259058 150574 259614
rect 149954 223614 150574 259058
rect 149954 223058 149986 223614
rect 150542 223058 150574 223614
rect 149954 187614 150574 223058
rect 149954 187058 149986 187614
rect 150542 187058 150574 187614
rect 149954 151614 150574 187058
rect 149954 151058 149986 151614
rect 150542 151058 150574 151614
rect 149954 115614 150574 151058
rect 149954 115058 149986 115614
rect 150542 115058 150574 115614
rect 149954 79614 150574 115058
rect 149954 79058 149986 79614
rect 150542 79058 150574 79614
rect 149954 43614 150574 79058
rect 149954 43058 149986 43614
rect 150542 43058 150574 43614
rect 149954 7614 150574 43058
rect 149954 7058 149986 7614
rect 150542 7058 150574 7614
rect 149954 -4186 150574 7058
rect 149954 -4742 149986 -4186
rect 150542 -4742 150574 -4186
rect 149954 -7654 150574 -4742
rect 151194 709638 151814 711590
rect 151194 709082 151226 709638
rect 151782 709082 151814 709638
rect 151194 692854 151814 709082
rect 151194 692298 151226 692854
rect 151782 692298 151814 692854
rect 151194 656854 151814 692298
rect 151194 656298 151226 656854
rect 151782 656298 151814 656854
rect 151194 620854 151814 656298
rect 151194 620298 151226 620854
rect 151782 620298 151814 620854
rect 151194 584854 151814 620298
rect 151194 584298 151226 584854
rect 151782 584298 151814 584854
rect 151194 548854 151814 584298
rect 151194 548298 151226 548854
rect 151782 548298 151814 548854
rect 151194 512854 151814 548298
rect 151194 512298 151226 512854
rect 151782 512298 151814 512854
rect 151194 476854 151814 512298
rect 151194 476298 151226 476854
rect 151782 476298 151814 476854
rect 151194 440854 151814 476298
rect 151194 440298 151226 440854
rect 151782 440298 151814 440854
rect 151194 404854 151814 440298
rect 151194 404298 151226 404854
rect 151782 404298 151814 404854
rect 151194 368854 151814 404298
rect 151194 368298 151226 368854
rect 151782 368298 151814 368854
rect 151194 332854 151814 368298
rect 151194 332298 151226 332854
rect 151782 332298 151814 332854
rect 151194 296854 151814 332298
rect 151194 296298 151226 296854
rect 151782 296298 151814 296854
rect 151194 260854 151814 296298
rect 151194 260298 151226 260854
rect 151782 260298 151814 260854
rect 151194 224854 151814 260298
rect 151194 224298 151226 224854
rect 151782 224298 151814 224854
rect 151194 188854 151814 224298
rect 151194 188298 151226 188854
rect 151782 188298 151814 188854
rect 151194 152854 151814 188298
rect 151194 152298 151226 152854
rect 151782 152298 151814 152854
rect 151194 116854 151814 152298
rect 151194 116298 151226 116854
rect 151782 116298 151814 116854
rect 151194 80854 151814 116298
rect 151194 80298 151226 80854
rect 151782 80298 151814 80854
rect 151194 44854 151814 80298
rect 151194 44298 151226 44854
rect 151782 44298 151814 44854
rect 151194 8854 151814 44298
rect 151194 8298 151226 8854
rect 151782 8298 151814 8854
rect 151194 -5146 151814 8298
rect 151194 -5702 151226 -5146
rect 151782 -5702 151814 -5146
rect 151194 -7654 151814 -5702
rect 152434 710598 153054 711590
rect 152434 710042 152466 710598
rect 153022 710042 153054 710598
rect 152434 694094 153054 710042
rect 152434 693538 152466 694094
rect 153022 693538 153054 694094
rect 152434 658094 153054 693538
rect 152434 657538 152466 658094
rect 153022 657538 153054 658094
rect 152434 622094 153054 657538
rect 152434 621538 152466 622094
rect 153022 621538 153054 622094
rect 152434 586094 153054 621538
rect 152434 585538 152466 586094
rect 153022 585538 153054 586094
rect 152434 550094 153054 585538
rect 152434 549538 152466 550094
rect 153022 549538 153054 550094
rect 152434 514094 153054 549538
rect 152434 513538 152466 514094
rect 153022 513538 153054 514094
rect 152434 478094 153054 513538
rect 152434 477538 152466 478094
rect 153022 477538 153054 478094
rect 152434 442094 153054 477538
rect 152434 441538 152466 442094
rect 153022 441538 153054 442094
rect 152434 406094 153054 441538
rect 152434 405538 152466 406094
rect 153022 405538 153054 406094
rect 152434 370094 153054 405538
rect 152434 369538 152466 370094
rect 153022 369538 153054 370094
rect 152434 334094 153054 369538
rect 152434 333538 152466 334094
rect 153022 333538 153054 334094
rect 152434 298094 153054 333538
rect 152434 297538 152466 298094
rect 153022 297538 153054 298094
rect 152434 262094 153054 297538
rect 152434 261538 152466 262094
rect 153022 261538 153054 262094
rect 152434 226094 153054 261538
rect 152434 225538 152466 226094
rect 153022 225538 153054 226094
rect 152434 190094 153054 225538
rect 152434 189538 152466 190094
rect 153022 189538 153054 190094
rect 152434 154094 153054 189538
rect 152434 153538 152466 154094
rect 153022 153538 153054 154094
rect 152434 118094 153054 153538
rect 152434 117538 152466 118094
rect 153022 117538 153054 118094
rect 152434 82094 153054 117538
rect 152434 81538 152466 82094
rect 153022 81538 153054 82094
rect 152434 46094 153054 81538
rect 152434 45538 152466 46094
rect 153022 45538 153054 46094
rect 152434 10094 153054 45538
rect 152434 9538 152466 10094
rect 153022 9538 153054 10094
rect 152434 -6106 153054 9538
rect 152434 -6662 152466 -6106
rect 153022 -6662 153054 -6106
rect 152434 -7654 153054 -6662
rect 153674 711558 154294 711590
rect 153674 711002 153706 711558
rect 154262 711002 154294 711558
rect 153674 695334 154294 711002
rect 153674 694778 153706 695334
rect 154262 694778 154294 695334
rect 153674 659334 154294 694778
rect 153674 658778 153706 659334
rect 154262 658778 154294 659334
rect 153674 623334 154294 658778
rect 153674 622778 153706 623334
rect 154262 622778 154294 623334
rect 153674 587334 154294 622778
rect 153674 586778 153706 587334
rect 154262 586778 154294 587334
rect 153674 551334 154294 586778
rect 153674 550778 153706 551334
rect 154262 550778 154294 551334
rect 153674 515334 154294 550778
rect 153674 514778 153706 515334
rect 154262 514778 154294 515334
rect 153674 479334 154294 514778
rect 153674 478778 153706 479334
rect 154262 478778 154294 479334
rect 153674 443334 154294 478778
rect 153674 442778 153706 443334
rect 154262 442778 154294 443334
rect 153674 407334 154294 442778
rect 153674 406778 153706 407334
rect 154262 406778 154294 407334
rect 153674 371334 154294 406778
rect 153674 370778 153706 371334
rect 154262 370778 154294 371334
rect 153674 335334 154294 370778
rect 153674 334778 153706 335334
rect 154262 334778 154294 335334
rect 153674 299334 154294 334778
rect 153674 298778 153706 299334
rect 154262 298778 154294 299334
rect 153674 263334 154294 298778
rect 153674 262778 153706 263334
rect 154262 262778 154294 263334
rect 153674 227334 154294 262778
rect 153674 226778 153706 227334
rect 154262 226778 154294 227334
rect 153674 191334 154294 226778
rect 153674 190778 153706 191334
rect 154262 190778 154294 191334
rect 153674 155334 154294 190778
rect 153674 154778 153706 155334
rect 154262 154778 154294 155334
rect 153674 119334 154294 154778
rect 153674 118778 153706 119334
rect 154262 118778 154294 119334
rect 153674 83334 154294 118778
rect 153674 82778 153706 83334
rect 154262 82778 154294 83334
rect 153674 47334 154294 82778
rect 153674 46778 153706 47334
rect 154262 46778 154294 47334
rect 153674 11334 154294 46778
rect 153674 10778 153706 11334
rect 154262 10778 154294 11334
rect 153674 -7066 154294 10778
rect 153674 -7622 153706 -7066
rect 154262 -7622 154294 -7066
rect 153674 -7654 154294 -7622
rect 180994 704838 181614 711590
rect 180994 704282 181026 704838
rect 181582 704282 181614 704838
rect 180994 686654 181614 704282
rect 180994 686098 181026 686654
rect 181582 686098 181614 686654
rect 180994 650654 181614 686098
rect 180994 650098 181026 650654
rect 181582 650098 181614 650654
rect 180994 614654 181614 650098
rect 180994 614098 181026 614654
rect 181582 614098 181614 614654
rect 180994 578654 181614 614098
rect 180994 578098 181026 578654
rect 181582 578098 181614 578654
rect 180994 542654 181614 578098
rect 180994 542098 181026 542654
rect 181582 542098 181614 542654
rect 180994 506654 181614 542098
rect 180994 506098 181026 506654
rect 181582 506098 181614 506654
rect 180994 470654 181614 506098
rect 180994 470098 181026 470654
rect 181582 470098 181614 470654
rect 180994 434654 181614 470098
rect 180994 434098 181026 434654
rect 181582 434098 181614 434654
rect 180994 398654 181614 434098
rect 180994 398098 181026 398654
rect 181582 398098 181614 398654
rect 180994 362654 181614 398098
rect 180994 362098 181026 362654
rect 181582 362098 181614 362654
rect 180994 326654 181614 362098
rect 180994 326098 181026 326654
rect 181582 326098 181614 326654
rect 180994 290654 181614 326098
rect 180994 290098 181026 290654
rect 181582 290098 181614 290654
rect 180994 254654 181614 290098
rect 180994 254098 181026 254654
rect 181582 254098 181614 254654
rect 180994 218654 181614 254098
rect 180994 218098 181026 218654
rect 181582 218098 181614 218654
rect 180994 182654 181614 218098
rect 180994 182098 181026 182654
rect 181582 182098 181614 182654
rect 180994 146654 181614 182098
rect 180994 146098 181026 146654
rect 181582 146098 181614 146654
rect 180994 110654 181614 146098
rect 180994 110098 181026 110654
rect 181582 110098 181614 110654
rect 180994 74654 181614 110098
rect 180994 74098 181026 74654
rect 181582 74098 181614 74654
rect 180994 38654 181614 74098
rect 180994 38098 181026 38654
rect 181582 38098 181614 38654
rect 180994 2654 181614 38098
rect 180994 2098 181026 2654
rect 181582 2098 181614 2654
rect 180994 -346 181614 2098
rect 180994 -902 181026 -346
rect 181582 -902 181614 -346
rect 180994 -7654 181614 -902
rect 182234 705798 182854 711590
rect 182234 705242 182266 705798
rect 182822 705242 182854 705798
rect 182234 687894 182854 705242
rect 182234 687338 182266 687894
rect 182822 687338 182854 687894
rect 182234 651894 182854 687338
rect 182234 651338 182266 651894
rect 182822 651338 182854 651894
rect 182234 615894 182854 651338
rect 182234 615338 182266 615894
rect 182822 615338 182854 615894
rect 182234 579894 182854 615338
rect 182234 579338 182266 579894
rect 182822 579338 182854 579894
rect 182234 543894 182854 579338
rect 182234 543338 182266 543894
rect 182822 543338 182854 543894
rect 182234 507894 182854 543338
rect 182234 507338 182266 507894
rect 182822 507338 182854 507894
rect 182234 471894 182854 507338
rect 182234 471338 182266 471894
rect 182822 471338 182854 471894
rect 182234 435894 182854 471338
rect 182234 435338 182266 435894
rect 182822 435338 182854 435894
rect 182234 399894 182854 435338
rect 182234 399338 182266 399894
rect 182822 399338 182854 399894
rect 182234 363894 182854 399338
rect 182234 363338 182266 363894
rect 182822 363338 182854 363894
rect 182234 327894 182854 363338
rect 182234 327338 182266 327894
rect 182822 327338 182854 327894
rect 182234 291894 182854 327338
rect 182234 291338 182266 291894
rect 182822 291338 182854 291894
rect 182234 255894 182854 291338
rect 182234 255338 182266 255894
rect 182822 255338 182854 255894
rect 182234 219894 182854 255338
rect 182234 219338 182266 219894
rect 182822 219338 182854 219894
rect 182234 183894 182854 219338
rect 182234 183338 182266 183894
rect 182822 183338 182854 183894
rect 182234 147894 182854 183338
rect 182234 147338 182266 147894
rect 182822 147338 182854 147894
rect 182234 111894 182854 147338
rect 182234 111338 182266 111894
rect 182822 111338 182854 111894
rect 182234 75894 182854 111338
rect 182234 75338 182266 75894
rect 182822 75338 182854 75894
rect 182234 39894 182854 75338
rect 182234 39338 182266 39894
rect 182822 39338 182854 39894
rect 182234 3894 182854 39338
rect 182234 3338 182266 3894
rect 182822 3338 182854 3894
rect 182234 -1306 182854 3338
rect 182234 -1862 182266 -1306
rect 182822 -1862 182854 -1306
rect 182234 -7654 182854 -1862
rect 183474 706758 184094 711590
rect 183474 706202 183506 706758
rect 184062 706202 184094 706758
rect 183474 689134 184094 706202
rect 183474 688578 183506 689134
rect 184062 688578 184094 689134
rect 183474 653134 184094 688578
rect 183474 652578 183506 653134
rect 184062 652578 184094 653134
rect 183474 617134 184094 652578
rect 183474 616578 183506 617134
rect 184062 616578 184094 617134
rect 183474 581134 184094 616578
rect 183474 580578 183506 581134
rect 184062 580578 184094 581134
rect 183474 545134 184094 580578
rect 183474 544578 183506 545134
rect 184062 544578 184094 545134
rect 183474 509134 184094 544578
rect 183474 508578 183506 509134
rect 184062 508578 184094 509134
rect 183474 473134 184094 508578
rect 183474 472578 183506 473134
rect 184062 472578 184094 473134
rect 183474 437134 184094 472578
rect 183474 436578 183506 437134
rect 184062 436578 184094 437134
rect 183474 401134 184094 436578
rect 183474 400578 183506 401134
rect 184062 400578 184094 401134
rect 183474 365134 184094 400578
rect 183474 364578 183506 365134
rect 184062 364578 184094 365134
rect 183474 329134 184094 364578
rect 183474 328578 183506 329134
rect 184062 328578 184094 329134
rect 183474 293134 184094 328578
rect 183474 292578 183506 293134
rect 184062 292578 184094 293134
rect 183474 257134 184094 292578
rect 183474 256578 183506 257134
rect 184062 256578 184094 257134
rect 183474 221134 184094 256578
rect 183474 220578 183506 221134
rect 184062 220578 184094 221134
rect 183474 185134 184094 220578
rect 183474 184578 183506 185134
rect 184062 184578 184094 185134
rect 183474 149134 184094 184578
rect 183474 148578 183506 149134
rect 184062 148578 184094 149134
rect 183474 113134 184094 148578
rect 183474 112578 183506 113134
rect 184062 112578 184094 113134
rect 183474 77134 184094 112578
rect 183474 76578 183506 77134
rect 184062 76578 184094 77134
rect 183474 41134 184094 76578
rect 183474 40578 183506 41134
rect 184062 40578 184094 41134
rect 183474 5134 184094 40578
rect 183474 4578 183506 5134
rect 184062 4578 184094 5134
rect 183474 -2266 184094 4578
rect 183474 -2822 183506 -2266
rect 184062 -2822 184094 -2266
rect 183474 -7654 184094 -2822
rect 184714 707718 185334 711590
rect 184714 707162 184746 707718
rect 185302 707162 185334 707718
rect 184714 690374 185334 707162
rect 184714 689818 184746 690374
rect 185302 689818 185334 690374
rect 184714 654374 185334 689818
rect 184714 653818 184746 654374
rect 185302 653818 185334 654374
rect 184714 618374 185334 653818
rect 184714 617818 184746 618374
rect 185302 617818 185334 618374
rect 184714 582374 185334 617818
rect 184714 581818 184746 582374
rect 185302 581818 185334 582374
rect 184714 546374 185334 581818
rect 184714 545818 184746 546374
rect 185302 545818 185334 546374
rect 184714 510374 185334 545818
rect 184714 509818 184746 510374
rect 185302 509818 185334 510374
rect 184714 474374 185334 509818
rect 184714 473818 184746 474374
rect 185302 473818 185334 474374
rect 184714 438374 185334 473818
rect 184714 437818 184746 438374
rect 185302 437818 185334 438374
rect 184714 402374 185334 437818
rect 184714 401818 184746 402374
rect 185302 401818 185334 402374
rect 184714 366374 185334 401818
rect 184714 365818 184746 366374
rect 185302 365818 185334 366374
rect 184714 330374 185334 365818
rect 184714 329818 184746 330374
rect 185302 329818 185334 330374
rect 184714 294374 185334 329818
rect 184714 293818 184746 294374
rect 185302 293818 185334 294374
rect 184714 258374 185334 293818
rect 184714 257818 184746 258374
rect 185302 257818 185334 258374
rect 184714 222374 185334 257818
rect 184714 221818 184746 222374
rect 185302 221818 185334 222374
rect 184714 186374 185334 221818
rect 184714 185818 184746 186374
rect 185302 185818 185334 186374
rect 184714 150374 185334 185818
rect 184714 149818 184746 150374
rect 185302 149818 185334 150374
rect 184714 114374 185334 149818
rect 184714 113818 184746 114374
rect 185302 113818 185334 114374
rect 184714 78374 185334 113818
rect 184714 77818 184746 78374
rect 185302 77818 185334 78374
rect 184714 42374 185334 77818
rect 184714 41818 184746 42374
rect 185302 41818 185334 42374
rect 184714 6374 185334 41818
rect 184714 5818 184746 6374
rect 185302 5818 185334 6374
rect 184714 -3226 185334 5818
rect 184714 -3782 184746 -3226
rect 185302 -3782 185334 -3226
rect 184714 -7654 185334 -3782
rect 185954 708678 186574 711590
rect 185954 708122 185986 708678
rect 186542 708122 186574 708678
rect 185954 691614 186574 708122
rect 185954 691058 185986 691614
rect 186542 691058 186574 691614
rect 185954 655614 186574 691058
rect 185954 655058 185986 655614
rect 186542 655058 186574 655614
rect 185954 619614 186574 655058
rect 185954 619058 185986 619614
rect 186542 619058 186574 619614
rect 185954 583614 186574 619058
rect 185954 583058 185986 583614
rect 186542 583058 186574 583614
rect 185954 547614 186574 583058
rect 185954 547058 185986 547614
rect 186542 547058 186574 547614
rect 185954 511614 186574 547058
rect 185954 511058 185986 511614
rect 186542 511058 186574 511614
rect 185954 475614 186574 511058
rect 185954 475058 185986 475614
rect 186542 475058 186574 475614
rect 185954 439614 186574 475058
rect 185954 439058 185986 439614
rect 186542 439058 186574 439614
rect 185954 403614 186574 439058
rect 185954 403058 185986 403614
rect 186542 403058 186574 403614
rect 185954 367614 186574 403058
rect 185954 367058 185986 367614
rect 186542 367058 186574 367614
rect 185954 331614 186574 367058
rect 185954 331058 185986 331614
rect 186542 331058 186574 331614
rect 185954 295614 186574 331058
rect 185954 295058 185986 295614
rect 186542 295058 186574 295614
rect 185954 259614 186574 295058
rect 185954 259058 185986 259614
rect 186542 259058 186574 259614
rect 185954 223614 186574 259058
rect 185954 223058 185986 223614
rect 186542 223058 186574 223614
rect 185954 187614 186574 223058
rect 185954 187058 185986 187614
rect 186542 187058 186574 187614
rect 185954 151614 186574 187058
rect 185954 151058 185986 151614
rect 186542 151058 186574 151614
rect 185954 115614 186574 151058
rect 185954 115058 185986 115614
rect 186542 115058 186574 115614
rect 185954 79614 186574 115058
rect 185954 79058 185986 79614
rect 186542 79058 186574 79614
rect 185954 43614 186574 79058
rect 185954 43058 185986 43614
rect 186542 43058 186574 43614
rect 185954 7614 186574 43058
rect 185954 7058 185986 7614
rect 186542 7058 186574 7614
rect 185954 -4186 186574 7058
rect 185954 -4742 185986 -4186
rect 186542 -4742 186574 -4186
rect 185954 -7654 186574 -4742
rect 187194 709638 187814 711590
rect 187194 709082 187226 709638
rect 187782 709082 187814 709638
rect 187194 692854 187814 709082
rect 187194 692298 187226 692854
rect 187782 692298 187814 692854
rect 187194 656854 187814 692298
rect 187194 656298 187226 656854
rect 187782 656298 187814 656854
rect 187194 620854 187814 656298
rect 187194 620298 187226 620854
rect 187782 620298 187814 620854
rect 187194 584854 187814 620298
rect 187194 584298 187226 584854
rect 187782 584298 187814 584854
rect 187194 548854 187814 584298
rect 187194 548298 187226 548854
rect 187782 548298 187814 548854
rect 187194 512854 187814 548298
rect 187194 512298 187226 512854
rect 187782 512298 187814 512854
rect 187194 476854 187814 512298
rect 187194 476298 187226 476854
rect 187782 476298 187814 476854
rect 187194 440854 187814 476298
rect 187194 440298 187226 440854
rect 187782 440298 187814 440854
rect 187194 404854 187814 440298
rect 187194 404298 187226 404854
rect 187782 404298 187814 404854
rect 187194 368854 187814 404298
rect 187194 368298 187226 368854
rect 187782 368298 187814 368854
rect 187194 332854 187814 368298
rect 187194 332298 187226 332854
rect 187782 332298 187814 332854
rect 187194 296854 187814 332298
rect 187194 296298 187226 296854
rect 187782 296298 187814 296854
rect 187194 260854 187814 296298
rect 187194 260298 187226 260854
rect 187782 260298 187814 260854
rect 187194 224854 187814 260298
rect 187194 224298 187226 224854
rect 187782 224298 187814 224854
rect 187194 188854 187814 224298
rect 187194 188298 187226 188854
rect 187782 188298 187814 188854
rect 187194 152854 187814 188298
rect 187194 152298 187226 152854
rect 187782 152298 187814 152854
rect 187194 116854 187814 152298
rect 187194 116298 187226 116854
rect 187782 116298 187814 116854
rect 187194 80854 187814 116298
rect 187194 80298 187226 80854
rect 187782 80298 187814 80854
rect 187194 44854 187814 80298
rect 187194 44298 187226 44854
rect 187782 44298 187814 44854
rect 187194 8854 187814 44298
rect 187194 8298 187226 8854
rect 187782 8298 187814 8854
rect 187194 -5146 187814 8298
rect 187194 -5702 187226 -5146
rect 187782 -5702 187814 -5146
rect 187194 -7654 187814 -5702
rect 188434 710598 189054 711590
rect 188434 710042 188466 710598
rect 189022 710042 189054 710598
rect 188434 694094 189054 710042
rect 188434 693538 188466 694094
rect 189022 693538 189054 694094
rect 188434 658094 189054 693538
rect 188434 657538 188466 658094
rect 189022 657538 189054 658094
rect 188434 622094 189054 657538
rect 188434 621538 188466 622094
rect 189022 621538 189054 622094
rect 188434 586094 189054 621538
rect 188434 585538 188466 586094
rect 189022 585538 189054 586094
rect 188434 550094 189054 585538
rect 188434 549538 188466 550094
rect 189022 549538 189054 550094
rect 188434 514094 189054 549538
rect 188434 513538 188466 514094
rect 189022 513538 189054 514094
rect 188434 478094 189054 513538
rect 188434 477538 188466 478094
rect 189022 477538 189054 478094
rect 188434 442094 189054 477538
rect 188434 441538 188466 442094
rect 189022 441538 189054 442094
rect 188434 406094 189054 441538
rect 188434 405538 188466 406094
rect 189022 405538 189054 406094
rect 188434 370094 189054 405538
rect 188434 369538 188466 370094
rect 189022 369538 189054 370094
rect 188434 334094 189054 369538
rect 188434 333538 188466 334094
rect 189022 333538 189054 334094
rect 188434 298094 189054 333538
rect 188434 297538 188466 298094
rect 189022 297538 189054 298094
rect 188434 262094 189054 297538
rect 188434 261538 188466 262094
rect 189022 261538 189054 262094
rect 188434 226094 189054 261538
rect 188434 225538 188466 226094
rect 189022 225538 189054 226094
rect 188434 190094 189054 225538
rect 188434 189538 188466 190094
rect 189022 189538 189054 190094
rect 188434 154094 189054 189538
rect 188434 153538 188466 154094
rect 189022 153538 189054 154094
rect 188434 118094 189054 153538
rect 188434 117538 188466 118094
rect 189022 117538 189054 118094
rect 188434 82094 189054 117538
rect 188434 81538 188466 82094
rect 189022 81538 189054 82094
rect 188434 46094 189054 81538
rect 188434 45538 188466 46094
rect 189022 45538 189054 46094
rect 188434 10094 189054 45538
rect 188434 9538 188466 10094
rect 189022 9538 189054 10094
rect 188434 -6106 189054 9538
rect 188434 -6662 188466 -6106
rect 189022 -6662 189054 -6106
rect 188434 -7654 189054 -6662
rect 189674 711558 190294 711590
rect 189674 711002 189706 711558
rect 190262 711002 190294 711558
rect 189674 695334 190294 711002
rect 189674 694778 189706 695334
rect 190262 694778 190294 695334
rect 189674 659334 190294 694778
rect 189674 658778 189706 659334
rect 190262 658778 190294 659334
rect 189674 623334 190294 658778
rect 189674 622778 189706 623334
rect 190262 622778 190294 623334
rect 189674 587334 190294 622778
rect 189674 586778 189706 587334
rect 190262 586778 190294 587334
rect 189674 551334 190294 586778
rect 189674 550778 189706 551334
rect 190262 550778 190294 551334
rect 189674 515334 190294 550778
rect 189674 514778 189706 515334
rect 190262 514778 190294 515334
rect 189674 479334 190294 514778
rect 189674 478778 189706 479334
rect 190262 478778 190294 479334
rect 189674 443334 190294 478778
rect 189674 442778 189706 443334
rect 190262 442778 190294 443334
rect 189674 407334 190294 442778
rect 189674 406778 189706 407334
rect 190262 406778 190294 407334
rect 189674 371334 190294 406778
rect 189674 370778 189706 371334
rect 190262 370778 190294 371334
rect 189674 335334 190294 370778
rect 189674 334778 189706 335334
rect 190262 334778 190294 335334
rect 189674 299334 190294 334778
rect 189674 298778 189706 299334
rect 190262 298778 190294 299334
rect 189674 263334 190294 298778
rect 189674 262778 189706 263334
rect 190262 262778 190294 263334
rect 189674 227334 190294 262778
rect 189674 226778 189706 227334
rect 190262 226778 190294 227334
rect 189674 191334 190294 226778
rect 189674 190778 189706 191334
rect 190262 190778 190294 191334
rect 189674 155334 190294 190778
rect 189674 154778 189706 155334
rect 190262 154778 190294 155334
rect 189674 119334 190294 154778
rect 189674 118778 189706 119334
rect 190262 118778 190294 119334
rect 189674 83334 190294 118778
rect 189674 82778 189706 83334
rect 190262 82778 190294 83334
rect 189674 47334 190294 82778
rect 189674 46778 189706 47334
rect 190262 46778 190294 47334
rect 189674 11334 190294 46778
rect 189674 10778 189706 11334
rect 190262 10778 190294 11334
rect 189674 -7066 190294 10778
rect 189674 -7622 189706 -7066
rect 190262 -7622 190294 -7066
rect 189674 -7654 190294 -7622
rect 216994 704838 217614 711590
rect 216994 704282 217026 704838
rect 217582 704282 217614 704838
rect 216994 686654 217614 704282
rect 216994 686098 217026 686654
rect 217582 686098 217614 686654
rect 216994 650654 217614 686098
rect 216994 650098 217026 650654
rect 217582 650098 217614 650654
rect 216994 614654 217614 650098
rect 216994 614098 217026 614654
rect 217582 614098 217614 614654
rect 216994 578654 217614 614098
rect 216994 578098 217026 578654
rect 217582 578098 217614 578654
rect 216994 542654 217614 578098
rect 216994 542098 217026 542654
rect 217582 542098 217614 542654
rect 216994 506654 217614 542098
rect 216994 506098 217026 506654
rect 217582 506098 217614 506654
rect 216994 470654 217614 506098
rect 216994 470098 217026 470654
rect 217582 470098 217614 470654
rect 216994 434654 217614 470098
rect 216994 434098 217026 434654
rect 217582 434098 217614 434654
rect 216994 398654 217614 434098
rect 216994 398098 217026 398654
rect 217582 398098 217614 398654
rect 216994 362654 217614 398098
rect 216994 362098 217026 362654
rect 217582 362098 217614 362654
rect 216994 326654 217614 362098
rect 216994 326098 217026 326654
rect 217582 326098 217614 326654
rect 216994 290654 217614 326098
rect 216994 290098 217026 290654
rect 217582 290098 217614 290654
rect 216994 254654 217614 290098
rect 216994 254098 217026 254654
rect 217582 254098 217614 254654
rect 216994 218654 217614 254098
rect 216994 218098 217026 218654
rect 217582 218098 217614 218654
rect 216994 182654 217614 218098
rect 216994 182098 217026 182654
rect 217582 182098 217614 182654
rect 216994 146654 217614 182098
rect 216994 146098 217026 146654
rect 217582 146098 217614 146654
rect 216994 110654 217614 146098
rect 216994 110098 217026 110654
rect 217582 110098 217614 110654
rect 216994 74654 217614 110098
rect 216994 74098 217026 74654
rect 217582 74098 217614 74654
rect 216994 38654 217614 74098
rect 216994 38098 217026 38654
rect 217582 38098 217614 38654
rect 216994 2654 217614 38098
rect 216994 2098 217026 2654
rect 217582 2098 217614 2654
rect 216994 -346 217614 2098
rect 216994 -902 217026 -346
rect 217582 -902 217614 -346
rect 216994 -7654 217614 -902
rect 218234 705798 218854 711590
rect 218234 705242 218266 705798
rect 218822 705242 218854 705798
rect 218234 687894 218854 705242
rect 218234 687338 218266 687894
rect 218822 687338 218854 687894
rect 218234 651894 218854 687338
rect 218234 651338 218266 651894
rect 218822 651338 218854 651894
rect 218234 615894 218854 651338
rect 218234 615338 218266 615894
rect 218822 615338 218854 615894
rect 218234 579894 218854 615338
rect 218234 579338 218266 579894
rect 218822 579338 218854 579894
rect 218234 543894 218854 579338
rect 218234 543338 218266 543894
rect 218822 543338 218854 543894
rect 218234 507894 218854 543338
rect 218234 507338 218266 507894
rect 218822 507338 218854 507894
rect 218234 471894 218854 507338
rect 218234 471338 218266 471894
rect 218822 471338 218854 471894
rect 218234 435894 218854 471338
rect 218234 435338 218266 435894
rect 218822 435338 218854 435894
rect 218234 399894 218854 435338
rect 218234 399338 218266 399894
rect 218822 399338 218854 399894
rect 218234 363894 218854 399338
rect 218234 363338 218266 363894
rect 218822 363338 218854 363894
rect 218234 327894 218854 363338
rect 218234 327338 218266 327894
rect 218822 327338 218854 327894
rect 218234 291894 218854 327338
rect 218234 291338 218266 291894
rect 218822 291338 218854 291894
rect 218234 255894 218854 291338
rect 218234 255338 218266 255894
rect 218822 255338 218854 255894
rect 218234 219894 218854 255338
rect 218234 219338 218266 219894
rect 218822 219338 218854 219894
rect 218234 183894 218854 219338
rect 218234 183338 218266 183894
rect 218822 183338 218854 183894
rect 218234 147894 218854 183338
rect 218234 147338 218266 147894
rect 218822 147338 218854 147894
rect 218234 111894 218854 147338
rect 218234 111338 218266 111894
rect 218822 111338 218854 111894
rect 218234 75894 218854 111338
rect 218234 75338 218266 75894
rect 218822 75338 218854 75894
rect 218234 39894 218854 75338
rect 218234 39338 218266 39894
rect 218822 39338 218854 39894
rect 218234 3894 218854 39338
rect 218234 3338 218266 3894
rect 218822 3338 218854 3894
rect 218234 -1306 218854 3338
rect 218234 -1862 218266 -1306
rect 218822 -1862 218854 -1306
rect 218234 -7654 218854 -1862
rect 219474 706758 220094 711590
rect 219474 706202 219506 706758
rect 220062 706202 220094 706758
rect 219474 689134 220094 706202
rect 219474 688578 219506 689134
rect 220062 688578 220094 689134
rect 219474 653134 220094 688578
rect 219474 652578 219506 653134
rect 220062 652578 220094 653134
rect 219474 617134 220094 652578
rect 219474 616578 219506 617134
rect 220062 616578 220094 617134
rect 219474 581134 220094 616578
rect 219474 580578 219506 581134
rect 220062 580578 220094 581134
rect 219474 545134 220094 580578
rect 219474 544578 219506 545134
rect 220062 544578 220094 545134
rect 219474 509134 220094 544578
rect 219474 508578 219506 509134
rect 220062 508578 220094 509134
rect 219474 473134 220094 508578
rect 219474 472578 219506 473134
rect 220062 472578 220094 473134
rect 219474 437134 220094 472578
rect 219474 436578 219506 437134
rect 220062 436578 220094 437134
rect 219474 401134 220094 436578
rect 219474 400578 219506 401134
rect 220062 400578 220094 401134
rect 219474 365134 220094 400578
rect 219474 364578 219506 365134
rect 220062 364578 220094 365134
rect 219474 329134 220094 364578
rect 219474 328578 219506 329134
rect 220062 328578 220094 329134
rect 219474 293134 220094 328578
rect 219474 292578 219506 293134
rect 220062 292578 220094 293134
rect 219474 257134 220094 292578
rect 219474 256578 219506 257134
rect 220062 256578 220094 257134
rect 219474 221134 220094 256578
rect 219474 220578 219506 221134
rect 220062 220578 220094 221134
rect 219474 185134 220094 220578
rect 219474 184578 219506 185134
rect 220062 184578 220094 185134
rect 219474 149134 220094 184578
rect 219474 148578 219506 149134
rect 220062 148578 220094 149134
rect 219474 113134 220094 148578
rect 219474 112578 219506 113134
rect 220062 112578 220094 113134
rect 219474 77134 220094 112578
rect 219474 76578 219506 77134
rect 220062 76578 220094 77134
rect 219474 41134 220094 76578
rect 219474 40578 219506 41134
rect 220062 40578 220094 41134
rect 219474 5134 220094 40578
rect 219474 4578 219506 5134
rect 220062 4578 220094 5134
rect 219474 -2266 220094 4578
rect 219474 -2822 219506 -2266
rect 220062 -2822 220094 -2266
rect 219474 -7654 220094 -2822
rect 220714 707718 221334 711590
rect 220714 707162 220746 707718
rect 221302 707162 221334 707718
rect 220714 690374 221334 707162
rect 220714 689818 220746 690374
rect 221302 689818 221334 690374
rect 220714 654374 221334 689818
rect 220714 653818 220746 654374
rect 221302 653818 221334 654374
rect 220714 618374 221334 653818
rect 220714 617818 220746 618374
rect 221302 617818 221334 618374
rect 220714 582374 221334 617818
rect 220714 581818 220746 582374
rect 221302 581818 221334 582374
rect 220714 546374 221334 581818
rect 220714 545818 220746 546374
rect 221302 545818 221334 546374
rect 220714 510374 221334 545818
rect 220714 509818 220746 510374
rect 221302 509818 221334 510374
rect 220714 474374 221334 509818
rect 220714 473818 220746 474374
rect 221302 473818 221334 474374
rect 220714 438374 221334 473818
rect 220714 437818 220746 438374
rect 221302 437818 221334 438374
rect 220714 402374 221334 437818
rect 220714 401818 220746 402374
rect 221302 401818 221334 402374
rect 220714 366374 221334 401818
rect 220714 365818 220746 366374
rect 221302 365818 221334 366374
rect 220714 330374 221334 365818
rect 220714 329818 220746 330374
rect 221302 329818 221334 330374
rect 220714 294374 221334 329818
rect 220714 293818 220746 294374
rect 221302 293818 221334 294374
rect 220714 258374 221334 293818
rect 220714 257818 220746 258374
rect 221302 257818 221334 258374
rect 220714 222374 221334 257818
rect 220714 221818 220746 222374
rect 221302 221818 221334 222374
rect 220714 186374 221334 221818
rect 220714 185818 220746 186374
rect 221302 185818 221334 186374
rect 220714 150374 221334 185818
rect 220714 149818 220746 150374
rect 221302 149818 221334 150374
rect 220714 114374 221334 149818
rect 220714 113818 220746 114374
rect 221302 113818 221334 114374
rect 220714 78374 221334 113818
rect 220714 77818 220746 78374
rect 221302 77818 221334 78374
rect 220714 42374 221334 77818
rect 220714 41818 220746 42374
rect 221302 41818 221334 42374
rect 220714 6374 221334 41818
rect 220714 5818 220746 6374
rect 221302 5818 221334 6374
rect 220714 -3226 221334 5818
rect 220714 -3782 220746 -3226
rect 221302 -3782 221334 -3226
rect 220714 -7654 221334 -3782
rect 221954 708678 222574 711590
rect 221954 708122 221986 708678
rect 222542 708122 222574 708678
rect 221954 691614 222574 708122
rect 221954 691058 221986 691614
rect 222542 691058 222574 691614
rect 221954 655614 222574 691058
rect 221954 655058 221986 655614
rect 222542 655058 222574 655614
rect 221954 619614 222574 655058
rect 221954 619058 221986 619614
rect 222542 619058 222574 619614
rect 221954 583614 222574 619058
rect 221954 583058 221986 583614
rect 222542 583058 222574 583614
rect 221954 547614 222574 583058
rect 221954 547058 221986 547614
rect 222542 547058 222574 547614
rect 221954 511614 222574 547058
rect 221954 511058 221986 511614
rect 222542 511058 222574 511614
rect 221954 475614 222574 511058
rect 221954 475058 221986 475614
rect 222542 475058 222574 475614
rect 221954 439614 222574 475058
rect 221954 439058 221986 439614
rect 222542 439058 222574 439614
rect 221954 403614 222574 439058
rect 221954 403058 221986 403614
rect 222542 403058 222574 403614
rect 221954 367614 222574 403058
rect 221954 367058 221986 367614
rect 222542 367058 222574 367614
rect 221954 331614 222574 367058
rect 221954 331058 221986 331614
rect 222542 331058 222574 331614
rect 221954 295614 222574 331058
rect 221954 295058 221986 295614
rect 222542 295058 222574 295614
rect 221954 259614 222574 295058
rect 221954 259058 221986 259614
rect 222542 259058 222574 259614
rect 221954 223614 222574 259058
rect 221954 223058 221986 223614
rect 222542 223058 222574 223614
rect 221954 187614 222574 223058
rect 221954 187058 221986 187614
rect 222542 187058 222574 187614
rect 221954 151614 222574 187058
rect 221954 151058 221986 151614
rect 222542 151058 222574 151614
rect 221954 115614 222574 151058
rect 221954 115058 221986 115614
rect 222542 115058 222574 115614
rect 221954 79614 222574 115058
rect 221954 79058 221986 79614
rect 222542 79058 222574 79614
rect 221954 43614 222574 79058
rect 221954 43058 221986 43614
rect 222542 43058 222574 43614
rect 221954 7614 222574 43058
rect 221954 7058 221986 7614
rect 222542 7058 222574 7614
rect 221954 -4186 222574 7058
rect 221954 -4742 221986 -4186
rect 222542 -4742 222574 -4186
rect 221954 -7654 222574 -4742
rect 223194 709638 223814 711590
rect 223194 709082 223226 709638
rect 223782 709082 223814 709638
rect 223194 692854 223814 709082
rect 223194 692298 223226 692854
rect 223782 692298 223814 692854
rect 223194 656854 223814 692298
rect 223194 656298 223226 656854
rect 223782 656298 223814 656854
rect 223194 620854 223814 656298
rect 223194 620298 223226 620854
rect 223782 620298 223814 620854
rect 223194 584854 223814 620298
rect 223194 584298 223226 584854
rect 223782 584298 223814 584854
rect 223194 548854 223814 584298
rect 223194 548298 223226 548854
rect 223782 548298 223814 548854
rect 223194 512854 223814 548298
rect 223194 512298 223226 512854
rect 223782 512298 223814 512854
rect 223194 476854 223814 512298
rect 223194 476298 223226 476854
rect 223782 476298 223814 476854
rect 223194 440854 223814 476298
rect 223194 440298 223226 440854
rect 223782 440298 223814 440854
rect 223194 404854 223814 440298
rect 223194 404298 223226 404854
rect 223782 404298 223814 404854
rect 223194 368854 223814 404298
rect 223194 368298 223226 368854
rect 223782 368298 223814 368854
rect 223194 332854 223814 368298
rect 223194 332298 223226 332854
rect 223782 332298 223814 332854
rect 223194 296854 223814 332298
rect 223194 296298 223226 296854
rect 223782 296298 223814 296854
rect 223194 260854 223814 296298
rect 223194 260298 223226 260854
rect 223782 260298 223814 260854
rect 223194 224854 223814 260298
rect 223194 224298 223226 224854
rect 223782 224298 223814 224854
rect 223194 188854 223814 224298
rect 223194 188298 223226 188854
rect 223782 188298 223814 188854
rect 223194 152854 223814 188298
rect 223194 152298 223226 152854
rect 223782 152298 223814 152854
rect 223194 116854 223814 152298
rect 223194 116298 223226 116854
rect 223782 116298 223814 116854
rect 223194 80854 223814 116298
rect 223194 80298 223226 80854
rect 223782 80298 223814 80854
rect 223194 44854 223814 80298
rect 223194 44298 223226 44854
rect 223782 44298 223814 44854
rect 223194 8854 223814 44298
rect 223194 8298 223226 8854
rect 223782 8298 223814 8854
rect 223194 -5146 223814 8298
rect 223194 -5702 223226 -5146
rect 223782 -5702 223814 -5146
rect 223194 -7654 223814 -5702
rect 224434 710598 225054 711590
rect 224434 710042 224466 710598
rect 225022 710042 225054 710598
rect 224434 694094 225054 710042
rect 224434 693538 224466 694094
rect 225022 693538 225054 694094
rect 224434 658094 225054 693538
rect 224434 657538 224466 658094
rect 225022 657538 225054 658094
rect 224434 622094 225054 657538
rect 224434 621538 224466 622094
rect 225022 621538 225054 622094
rect 224434 586094 225054 621538
rect 224434 585538 224466 586094
rect 225022 585538 225054 586094
rect 224434 550094 225054 585538
rect 224434 549538 224466 550094
rect 225022 549538 225054 550094
rect 224434 514094 225054 549538
rect 224434 513538 224466 514094
rect 225022 513538 225054 514094
rect 224434 478094 225054 513538
rect 224434 477538 224466 478094
rect 225022 477538 225054 478094
rect 224434 442094 225054 477538
rect 224434 441538 224466 442094
rect 225022 441538 225054 442094
rect 224434 406094 225054 441538
rect 224434 405538 224466 406094
rect 225022 405538 225054 406094
rect 224434 370094 225054 405538
rect 224434 369538 224466 370094
rect 225022 369538 225054 370094
rect 224434 334094 225054 369538
rect 224434 333538 224466 334094
rect 225022 333538 225054 334094
rect 224434 298094 225054 333538
rect 224434 297538 224466 298094
rect 225022 297538 225054 298094
rect 224434 262094 225054 297538
rect 224434 261538 224466 262094
rect 225022 261538 225054 262094
rect 224434 226094 225054 261538
rect 224434 225538 224466 226094
rect 225022 225538 225054 226094
rect 224434 190094 225054 225538
rect 224434 189538 224466 190094
rect 225022 189538 225054 190094
rect 224434 154094 225054 189538
rect 224434 153538 224466 154094
rect 225022 153538 225054 154094
rect 224434 118094 225054 153538
rect 224434 117538 224466 118094
rect 225022 117538 225054 118094
rect 224434 82094 225054 117538
rect 224434 81538 224466 82094
rect 225022 81538 225054 82094
rect 224434 46094 225054 81538
rect 224434 45538 224466 46094
rect 225022 45538 225054 46094
rect 224434 10094 225054 45538
rect 224434 9538 224466 10094
rect 225022 9538 225054 10094
rect 224434 -6106 225054 9538
rect 224434 -6662 224466 -6106
rect 225022 -6662 225054 -6106
rect 224434 -7654 225054 -6662
rect 225674 711558 226294 711590
rect 225674 711002 225706 711558
rect 226262 711002 226294 711558
rect 225674 695334 226294 711002
rect 225674 694778 225706 695334
rect 226262 694778 226294 695334
rect 225674 659334 226294 694778
rect 225674 658778 225706 659334
rect 226262 658778 226294 659334
rect 225674 623334 226294 658778
rect 225674 622778 225706 623334
rect 226262 622778 226294 623334
rect 225674 587334 226294 622778
rect 225674 586778 225706 587334
rect 226262 586778 226294 587334
rect 225674 551334 226294 586778
rect 225674 550778 225706 551334
rect 226262 550778 226294 551334
rect 225674 515334 226294 550778
rect 225674 514778 225706 515334
rect 226262 514778 226294 515334
rect 225674 479334 226294 514778
rect 225674 478778 225706 479334
rect 226262 478778 226294 479334
rect 225674 443334 226294 478778
rect 225674 442778 225706 443334
rect 226262 442778 226294 443334
rect 225674 407334 226294 442778
rect 225674 406778 225706 407334
rect 226262 406778 226294 407334
rect 225674 371334 226294 406778
rect 225674 370778 225706 371334
rect 226262 370778 226294 371334
rect 225674 335334 226294 370778
rect 225674 334778 225706 335334
rect 226262 334778 226294 335334
rect 225674 299334 226294 334778
rect 225674 298778 225706 299334
rect 226262 298778 226294 299334
rect 225674 263334 226294 298778
rect 225674 262778 225706 263334
rect 226262 262778 226294 263334
rect 225674 227334 226294 262778
rect 225674 226778 225706 227334
rect 226262 226778 226294 227334
rect 225674 191334 226294 226778
rect 225674 190778 225706 191334
rect 226262 190778 226294 191334
rect 225674 155334 226294 190778
rect 225674 154778 225706 155334
rect 226262 154778 226294 155334
rect 225674 119334 226294 154778
rect 225674 118778 225706 119334
rect 226262 118778 226294 119334
rect 225674 83334 226294 118778
rect 225674 82778 225706 83334
rect 226262 82778 226294 83334
rect 225674 47334 226294 82778
rect 225674 46778 225706 47334
rect 226262 46778 226294 47334
rect 225674 11334 226294 46778
rect 225674 10778 225706 11334
rect 226262 10778 226294 11334
rect 225674 -7066 226294 10778
rect 225674 -7622 225706 -7066
rect 226262 -7622 226294 -7066
rect 225674 -7654 226294 -7622
rect 252994 704838 253614 711590
rect 252994 704282 253026 704838
rect 253582 704282 253614 704838
rect 252994 686654 253614 704282
rect 252994 686098 253026 686654
rect 253582 686098 253614 686654
rect 252994 650654 253614 686098
rect 252994 650098 253026 650654
rect 253582 650098 253614 650654
rect 252994 614654 253614 650098
rect 252994 614098 253026 614654
rect 253582 614098 253614 614654
rect 252994 578654 253614 614098
rect 252994 578098 253026 578654
rect 253582 578098 253614 578654
rect 252994 542654 253614 578098
rect 252994 542098 253026 542654
rect 253582 542098 253614 542654
rect 252994 506654 253614 542098
rect 252994 506098 253026 506654
rect 253582 506098 253614 506654
rect 252994 470654 253614 506098
rect 252994 470098 253026 470654
rect 253582 470098 253614 470654
rect 252994 434654 253614 470098
rect 252994 434098 253026 434654
rect 253582 434098 253614 434654
rect 252994 398654 253614 434098
rect 252994 398098 253026 398654
rect 253582 398098 253614 398654
rect 252994 362654 253614 398098
rect 252994 362098 253026 362654
rect 253582 362098 253614 362654
rect 252994 326654 253614 362098
rect 252994 326098 253026 326654
rect 253582 326098 253614 326654
rect 252994 290654 253614 326098
rect 252994 290098 253026 290654
rect 253582 290098 253614 290654
rect 252994 254654 253614 290098
rect 252994 254098 253026 254654
rect 253582 254098 253614 254654
rect 252994 218654 253614 254098
rect 252994 218098 253026 218654
rect 253582 218098 253614 218654
rect 252994 182654 253614 218098
rect 252994 182098 253026 182654
rect 253582 182098 253614 182654
rect 252994 146654 253614 182098
rect 252994 146098 253026 146654
rect 253582 146098 253614 146654
rect 252994 110654 253614 146098
rect 252994 110098 253026 110654
rect 253582 110098 253614 110654
rect 252994 74654 253614 110098
rect 252994 74098 253026 74654
rect 253582 74098 253614 74654
rect 252994 38654 253614 74098
rect 252994 38098 253026 38654
rect 253582 38098 253614 38654
rect 252994 2654 253614 38098
rect 252994 2098 253026 2654
rect 253582 2098 253614 2654
rect 252994 -346 253614 2098
rect 252994 -902 253026 -346
rect 253582 -902 253614 -346
rect 252994 -7654 253614 -902
rect 254234 705798 254854 711590
rect 254234 705242 254266 705798
rect 254822 705242 254854 705798
rect 254234 687894 254854 705242
rect 254234 687338 254266 687894
rect 254822 687338 254854 687894
rect 254234 651894 254854 687338
rect 254234 651338 254266 651894
rect 254822 651338 254854 651894
rect 254234 615894 254854 651338
rect 254234 615338 254266 615894
rect 254822 615338 254854 615894
rect 254234 579894 254854 615338
rect 254234 579338 254266 579894
rect 254822 579338 254854 579894
rect 254234 543894 254854 579338
rect 254234 543338 254266 543894
rect 254822 543338 254854 543894
rect 254234 507894 254854 543338
rect 254234 507338 254266 507894
rect 254822 507338 254854 507894
rect 254234 471894 254854 507338
rect 254234 471338 254266 471894
rect 254822 471338 254854 471894
rect 254234 435894 254854 471338
rect 254234 435338 254266 435894
rect 254822 435338 254854 435894
rect 254234 399894 254854 435338
rect 254234 399338 254266 399894
rect 254822 399338 254854 399894
rect 254234 363894 254854 399338
rect 254234 363338 254266 363894
rect 254822 363338 254854 363894
rect 254234 327894 254854 363338
rect 254234 327338 254266 327894
rect 254822 327338 254854 327894
rect 254234 291894 254854 327338
rect 254234 291338 254266 291894
rect 254822 291338 254854 291894
rect 254234 255894 254854 291338
rect 254234 255338 254266 255894
rect 254822 255338 254854 255894
rect 254234 219894 254854 255338
rect 254234 219338 254266 219894
rect 254822 219338 254854 219894
rect 254234 183894 254854 219338
rect 254234 183338 254266 183894
rect 254822 183338 254854 183894
rect 254234 147894 254854 183338
rect 254234 147338 254266 147894
rect 254822 147338 254854 147894
rect 254234 111894 254854 147338
rect 254234 111338 254266 111894
rect 254822 111338 254854 111894
rect 254234 75894 254854 111338
rect 254234 75338 254266 75894
rect 254822 75338 254854 75894
rect 254234 39894 254854 75338
rect 254234 39338 254266 39894
rect 254822 39338 254854 39894
rect 254234 3894 254854 39338
rect 254234 3338 254266 3894
rect 254822 3338 254854 3894
rect 254234 -1306 254854 3338
rect 254234 -1862 254266 -1306
rect 254822 -1862 254854 -1306
rect 254234 -7654 254854 -1862
rect 255474 706758 256094 711590
rect 255474 706202 255506 706758
rect 256062 706202 256094 706758
rect 255474 689134 256094 706202
rect 255474 688578 255506 689134
rect 256062 688578 256094 689134
rect 255474 653134 256094 688578
rect 255474 652578 255506 653134
rect 256062 652578 256094 653134
rect 255474 617134 256094 652578
rect 255474 616578 255506 617134
rect 256062 616578 256094 617134
rect 255474 581134 256094 616578
rect 255474 580578 255506 581134
rect 256062 580578 256094 581134
rect 255474 545134 256094 580578
rect 255474 544578 255506 545134
rect 256062 544578 256094 545134
rect 255474 509134 256094 544578
rect 255474 508578 255506 509134
rect 256062 508578 256094 509134
rect 255474 473134 256094 508578
rect 255474 472578 255506 473134
rect 256062 472578 256094 473134
rect 255474 437134 256094 472578
rect 255474 436578 255506 437134
rect 256062 436578 256094 437134
rect 255474 401134 256094 436578
rect 255474 400578 255506 401134
rect 256062 400578 256094 401134
rect 255474 365134 256094 400578
rect 255474 364578 255506 365134
rect 256062 364578 256094 365134
rect 255474 329134 256094 364578
rect 255474 328578 255506 329134
rect 256062 328578 256094 329134
rect 255474 293134 256094 328578
rect 255474 292578 255506 293134
rect 256062 292578 256094 293134
rect 255474 257134 256094 292578
rect 255474 256578 255506 257134
rect 256062 256578 256094 257134
rect 255474 221134 256094 256578
rect 255474 220578 255506 221134
rect 256062 220578 256094 221134
rect 255474 185134 256094 220578
rect 255474 184578 255506 185134
rect 256062 184578 256094 185134
rect 255474 149134 256094 184578
rect 255474 148578 255506 149134
rect 256062 148578 256094 149134
rect 255474 113134 256094 148578
rect 255474 112578 255506 113134
rect 256062 112578 256094 113134
rect 255474 77134 256094 112578
rect 255474 76578 255506 77134
rect 256062 76578 256094 77134
rect 255474 41134 256094 76578
rect 255474 40578 255506 41134
rect 256062 40578 256094 41134
rect 255474 5134 256094 40578
rect 255474 4578 255506 5134
rect 256062 4578 256094 5134
rect 255474 -2266 256094 4578
rect 255474 -2822 255506 -2266
rect 256062 -2822 256094 -2266
rect 255474 -7654 256094 -2822
rect 256714 707718 257334 711590
rect 256714 707162 256746 707718
rect 257302 707162 257334 707718
rect 256714 690374 257334 707162
rect 256714 689818 256746 690374
rect 257302 689818 257334 690374
rect 256714 654374 257334 689818
rect 256714 653818 256746 654374
rect 257302 653818 257334 654374
rect 256714 618374 257334 653818
rect 256714 617818 256746 618374
rect 257302 617818 257334 618374
rect 256714 582374 257334 617818
rect 256714 581818 256746 582374
rect 257302 581818 257334 582374
rect 256714 546374 257334 581818
rect 256714 545818 256746 546374
rect 257302 545818 257334 546374
rect 256714 510374 257334 545818
rect 256714 509818 256746 510374
rect 257302 509818 257334 510374
rect 256714 474374 257334 509818
rect 256714 473818 256746 474374
rect 257302 473818 257334 474374
rect 256714 438374 257334 473818
rect 256714 437818 256746 438374
rect 257302 437818 257334 438374
rect 256714 402374 257334 437818
rect 256714 401818 256746 402374
rect 257302 401818 257334 402374
rect 256714 366374 257334 401818
rect 256714 365818 256746 366374
rect 257302 365818 257334 366374
rect 256714 330374 257334 365818
rect 256714 329818 256746 330374
rect 257302 329818 257334 330374
rect 256714 294374 257334 329818
rect 256714 293818 256746 294374
rect 257302 293818 257334 294374
rect 256714 258374 257334 293818
rect 256714 257818 256746 258374
rect 257302 257818 257334 258374
rect 256714 222374 257334 257818
rect 256714 221818 256746 222374
rect 257302 221818 257334 222374
rect 256714 186374 257334 221818
rect 256714 185818 256746 186374
rect 257302 185818 257334 186374
rect 256714 150374 257334 185818
rect 256714 149818 256746 150374
rect 257302 149818 257334 150374
rect 256714 114374 257334 149818
rect 256714 113818 256746 114374
rect 257302 113818 257334 114374
rect 256714 78374 257334 113818
rect 256714 77818 256746 78374
rect 257302 77818 257334 78374
rect 256714 42374 257334 77818
rect 256714 41818 256746 42374
rect 257302 41818 257334 42374
rect 256714 6374 257334 41818
rect 256714 5818 256746 6374
rect 257302 5818 257334 6374
rect 256714 -3226 257334 5818
rect 256714 -3782 256746 -3226
rect 257302 -3782 257334 -3226
rect 256714 -7654 257334 -3782
rect 257954 708678 258574 711590
rect 257954 708122 257986 708678
rect 258542 708122 258574 708678
rect 257954 691614 258574 708122
rect 257954 691058 257986 691614
rect 258542 691058 258574 691614
rect 257954 655614 258574 691058
rect 257954 655058 257986 655614
rect 258542 655058 258574 655614
rect 257954 619614 258574 655058
rect 257954 619058 257986 619614
rect 258542 619058 258574 619614
rect 257954 583614 258574 619058
rect 257954 583058 257986 583614
rect 258542 583058 258574 583614
rect 257954 547614 258574 583058
rect 257954 547058 257986 547614
rect 258542 547058 258574 547614
rect 257954 511614 258574 547058
rect 257954 511058 257986 511614
rect 258542 511058 258574 511614
rect 257954 475614 258574 511058
rect 257954 475058 257986 475614
rect 258542 475058 258574 475614
rect 257954 439614 258574 475058
rect 257954 439058 257986 439614
rect 258542 439058 258574 439614
rect 257954 403614 258574 439058
rect 257954 403058 257986 403614
rect 258542 403058 258574 403614
rect 257954 367614 258574 403058
rect 257954 367058 257986 367614
rect 258542 367058 258574 367614
rect 257954 331614 258574 367058
rect 257954 331058 257986 331614
rect 258542 331058 258574 331614
rect 257954 295614 258574 331058
rect 257954 295058 257986 295614
rect 258542 295058 258574 295614
rect 257954 259614 258574 295058
rect 257954 259058 257986 259614
rect 258542 259058 258574 259614
rect 257954 223614 258574 259058
rect 257954 223058 257986 223614
rect 258542 223058 258574 223614
rect 257954 187614 258574 223058
rect 257954 187058 257986 187614
rect 258542 187058 258574 187614
rect 257954 151614 258574 187058
rect 257954 151058 257986 151614
rect 258542 151058 258574 151614
rect 257954 115614 258574 151058
rect 257954 115058 257986 115614
rect 258542 115058 258574 115614
rect 257954 79614 258574 115058
rect 257954 79058 257986 79614
rect 258542 79058 258574 79614
rect 257954 43614 258574 79058
rect 257954 43058 257986 43614
rect 258542 43058 258574 43614
rect 257954 7614 258574 43058
rect 257954 7058 257986 7614
rect 258542 7058 258574 7614
rect 257954 -4186 258574 7058
rect 257954 -4742 257986 -4186
rect 258542 -4742 258574 -4186
rect 257954 -7654 258574 -4742
rect 259194 709638 259814 711590
rect 259194 709082 259226 709638
rect 259782 709082 259814 709638
rect 259194 692854 259814 709082
rect 259194 692298 259226 692854
rect 259782 692298 259814 692854
rect 259194 656854 259814 692298
rect 259194 656298 259226 656854
rect 259782 656298 259814 656854
rect 259194 620854 259814 656298
rect 259194 620298 259226 620854
rect 259782 620298 259814 620854
rect 259194 584854 259814 620298
rect 259194 584298 259226 584854
rect 259782 584298 259814 584854
rect 259194 548854 259814 584298
rect 259194 548298 259226 548854
rect 259782 548298 259814 548854
rect 259194 512854 259814 548298
rect 259194 512298 259226 512854
rect 259782 512298 259814 512854
rect 259194 476854 259814 512298
rect 259194 476298 259226 476854
rect 259782 476298 259814 476854
rect 259194 440854 259814 476298
rect 259194 440298 259226 440854
rect 259782 440298 259814 440854
rect 259194 404854 259814 440298
rect 259194 404298 259226 404854
rect 259782 404298 259814 404854
rect 259194 368854 259814 404298
rect 259194 368298 259226 368854
rect 259782 368298 259814 368854
rect 259194 332854 259814 368298
rect 259194 332298 259226 332854
rect 259782 332298 259814 332854
rect 259194 296854 259814 332298
rect 259194 296298 259226 296854
rect 259782 296298 259814 296854
rect 259194 260854 259814 296298
rect 259194 260298 259226 260854
rect 259782 260298 259814 260854
rect 259194 224854 259814 260298
rect 259194 224298 259226 224854
rect 259782 224298 259814 224854
rect 259194 188854 259814 224298
rect 259194 188298 259226 188854
rect 259782 188298 259814 188854
rect 259194 152854 259814 188298
rect 259194 152298 259226 152854
rect 259782 152298 259814 152854
rect 259194 116854 259814 152298
rect 259194 116298 259226 116854
rect 259782 116298 259814 116854
rect 259194 80854 259814 116298
rect 259194 80298 259226 80854
rect 259782 80298 259814 80854
rect 259194 44854 259814 80298
rect 259194 44298 259226 44854
rect 259782 44298 259814 44854
rect 259194 8854 259814 44298
rect 259194 8298 259226 8854
rect 259782 8298 259814 8854
rect 259194 -5146 259814 8298
rect 259194 -5702 259226 -5146
rect 259782 -5702 259814 -5146
rect 259194 -7654 259814 -5702
rect 260434 710598 261054 711590
rect 260434 710042 260466 710598
rect 261022 710042 261054 710598
rect 260434 694094 261054 710042
rect 260434 693538 260466 694094
rect 261022 693538 261054 694094
rect 260434 658094 261054 693538
rect 260434 657538 260466 658094
rect 261022 657538 261054 658094
rect 260434 622094 261054 657538
rect 260434 621538 260466 622094
rect 261022 621538 261054 622094
rect 260434 586094 261054 621538
rect 260434 585538 260466 586094
rect 261022 585538 261054 586094
rect 260434 550094 261054 585538
rect 260434 549538 260466 550094
rect 261022 549538 261054 550094
rect 260434 514094 261054 549538
rect 260434 513538 260466 514094
rect 261022 513538 261054 514094
rect 260434 478094 261054 513538
rect 260434 477538 260466 478094
rect 261022 477538 261054 478094
rect 260434 442094 261054 477538
rect 260434 441538 260466 442094
rect 261022 441538 261054 442094
rect 260434 406094 261054 441538
rect 260434 405538 260466 406094
rect 261022 405538 261054 406094
rect 260434 370094 261054 405538
rect 260434 369538 260466 370094
rect 261022 369538 261054 370094
rect 260434 334094 261054 369538
rect 260434 333538 260466 334094
rect 261022 333538 261054 334094
rect 260434 298094 261054 333538
rect 260434 297538 260466 298094
rect 261022 297538 261054 298094
rect 260434 262094 261054 297538
rect 260434 261538 260466 262094
rect 261022 261538 261054 262094
rect 260434 226094 261054 261538
rect 260434 225538 260466 226094
rect 261022 225538 261054 226094
rect 260434 190094 261054 225538
rect 260434 189538 260466 190094
rect 261022 189538 261054 190094
rect 260434 154094 261054 189538
rect 260434 153538 260466 154094
rect 261022 153538 261054 154094
rect 260434 118094 261054 153538
rect 260434 117538 260466 118094
rect 261022 117538 261054 118094
rect 260434 82094 261054 117538
rect 260434 81538 260466 82094
rect 261022 81538 261054 82094
rect 260434 46094 261054 81538
rect 260434 45538 260466 46094
rect 261022 45538 261054 46094
rect 260434 10094 261054 45538
rect 260434 9538 260466 10094
rect 261022 9538 261054 10094
rect 260434 -6106 261054 9538
rect 260434 -6662 260466 -6106
rect 261022 -6662 261054 -6106
rect 260434 -7654 261054 -6662
rect 261674 711558 262294 711590
rect 261674 711002 261706 711558
rect 262262 711002 262294 711558
rect 261674 695334 262294 711002
rect 261674 694778 261706 695334
rect 262262 694778 262294 695334
rect 261674 659334 262294 694778
rect 261674 658778 261706 659334
rect 262262 658778 262294 659334
rect 261674 623334 262294 658778
rect 261674 622778 261706 623334
rect 262262 622778 262294 623334
rect 261674 587334 262294 622778
rect 261674 586778 261706 587334
rect 262262 586778 262294 587334
rect 261674 551334 262294 586778
rect 261674 550778 261706 551334
rect 262262 550778 262294 551334
rect 261674 515334 262294 550778
rect 261674 514778 261706 515334
rect 262262 514778 262294 515334
rect 261674 479334 262294 514778
rect 261674 478778 261706 479334
rect 262262 478778 262294 479334
rect 261674 443334 262294 478778
rect 261674 442778 261706 443334
rect 262262 442778 262294 443334
rect 261674 407334 262294 442778
rect 261674 406778 261706 407334
rect 262262 406778 262294 407334
rect 261674 371334 262294 406778
rect 261674 370778 261706 371334
rect 262262 370778 262294 371334
rect 261674 335334 262294 370778
rect 261674 334778 261706 335334
rect 262262 334778 262294 335334
rect 261674 299334 262294 334778
rect 261674 298778 261706 299334
rect 262262 298778 262294 299334
rect 261674 263334 262294 298778
rect 261674 262778 261706 263334
rect 262262 262778 262294 263334
rect 261674 227334 262294 262778
rect 261674 226778 261706 227334
rect 262262 226778 262294 227334
rect 261674 191334 262294 226778
rect 261674 190778 261706 191334
rect 262262 190778 262294 191334
rect 261674 155334 262294 190778
rect 261674 154778 261706 155334
rect 262262 154778 262294 155334
rect 261674 119334 262294 154778
rect 261674 118778 261706 119334
rect 262262 118778 262294 119334
rect 261674 83334 262294 118778
rect 261674 82778 261706 83334
rect 262262 82778 262294 83334
rect 261674 47334 262294 82778
rect 261674 46778 261706 47334
rect 262262 46778 262294 47334
rect 261674 11334 262294 46778
rect 261674 10778 261706 11334
rect 262262 10778 262294 11334
rect 261674 -7066 262294 10778
rect 261674 -7622 261706 -7066
rect 262262 -7622 262294 -7066
rect 261674 -7654 262294 -7622
rect 288994 704838 289614 711590
rect 288994 704282 289026 704838
rect 289582 704282 289614 704838
rect 288994 686654 289614 704282
rect 288994 686098 289026 686654
rect 289582 686098 289614 686654
rect 288994 650654 289614 686098
rect 288994 650098 289026 650654
rect 289582 650098 289614 650654
rect 288994 614654 289614 650098
rect 288994 614098 289026 614654
rect 289582 614098 289614 614654
rect 288994 578654 289614 614098
rect 288994 578098 289026 578654
rect 289582 578098 289614 578654
rect 288994 542654 289614 578098
rect 288994 542098 289026 542654
rect 289582 542098 289614 542654
rect 288994 506654 289614 542098
rect 288994 506098 289026 506654
rect 289582 506098 289614 506654
rect 288994 470654 289614 506098
rect 288994 470098 289026 470654
rect 289582 470098 289614 470654
rect 288994 434654 289614 470098
rect 288994 434098 289026 434654
rect 289582 434098 289614 434654
rect 288994 398654 289614 434098
rect 288994 398098 289026 398654
rect 289582 398098 289614 398654
rect 288994 362654 289614 398098
rect 288994 362098 289026 362654
rect 289582 362098 289614 362654
rect 288994 326654 289614 362098
rect 288994 326098 289026 326654
rect 289582 326098 289614 326654
rect 288994 290654 289614 326098
rect 288994 290098 289026 290654
rect 289582 290098 289614 290654
rect 288994 254654 289614 290098
rect 288994 254098 289026 254654
rect 289582 254098 289614 254654
rect 288994 218654 289614 254098
rect 288994 218098 289026 218654
rect 289582 218098 289614 218654
rect 288994 182654 289614 218098
rect 288994 182098 289026 182654
rect 289582 182098 289614 182654
rect 288994 146654 289614 182098
rect 288994 146098 289026 146654
rect 289582 146098 289614 146654
rect 288994 110654 289614 146098
rect 288994 110098 289026 110654
rect 289582 110098 289614 110654
rect 288994 74654 289614 110098
rect 288994 74098 289026 74654
rect 289582 74098 289614 74654
rect 288994 38654 289614 74098
rect 288994 38098 289026 38654
rect 289582 38098 289614 38654
rect 288994 2654 289614 38098
rect 288994 2098 289026 2654
rect 289582 2098 289614 2654
rect 288994 -346 289614 2098
rect 288994 -902 289026 -346
rect 289582 -902 289614 -346
rect 288994 -7654 289614 -902
rect 290234 705798 290854 711590
rect 290234 705242 290266 705798
rect 290822 705242 290854 705798
rect 290234 687894 290854 705242
rect 290234 687338 290266 687894
rect 290822 687338 290854 687894
rect 290234 651894 290854 687338
rect 290234 651338 290266 651894
rect 290822 651338 290854 651894
rect 290234 615894 290854 651338
rect 290234 615338 290266 615894
rect 290822 615338 290854 615894
rect 290234 579894 290854 615338
rect 290234 579338 290266 579894
rect 290822 579338 290854 579894
rect 290234 543894 290854 579338
rect 290234 543338 290266 543894
rect 290822 543338 290854 543894
rect 290234 507894 290854 543338
rect 290234 507338 290266 507894
rect 290822 507338 290854 507894
rect 290234 471894 290854 507338
rect 290234 471338 290266 471894
rect 290822 471338 290854 471894
rect 290234 435894 290854 471338
rect 290234 435338 290266 435894
rect 290822 435338 290854 435894
rect 290234 399894 290854 435338
rect 290234 399338 290266 399894
rect 290822 399338 290854 399894
rect 290234 363894 290854 399338
rect 290234 363338 290266 363894
rect 290822 363338 290854 363894
rect 290234 327894 290854 363338
rect 290234 327338 290266 327894
rect 290822 327338 290854 327894
rect 290234 291894 290854 327338
rect 290234 291338 290266 291894
rect 290822 291338 290854 291894
rect 290234 255894 290854 291338
rect 290234 255338 290266 255894
rect 290822 255338 290854 255894
rect 290234 219894 290854 255338
rect 290234 219338 290266 219894
rect 290822 219338 290854 219894
rect 290234 183894 290854 219338
rect 290234 183338 290266 183894
rect 290822 183338 290854 183894
rect 290234 147894 290854 183338
rect 290234 147338 290266 147894
rect 290822 147338 290854 147894
rect 290234 111894 290854 147338
rect 290234 111338 290266 111894
rect 290822 111338 290854 111894
rect 290234 75894 290854 111338
rect 290234 75338 290266 75894
rect 290822 75338 290854 75894
rect 290234 39894 290854 75338
rect 290234 39338 290266 39894
rect 290822 39338 290854 39894
rect 290234 3894 290854 39338
rect 290234 3338 290266 3894
rect 290822 3338 290854 3894
rect 290234 -1306 290854 3338
rect 290234 -1862 290266 -1306
rect 290822 -1862 290854 -1306
rect 290234 -7654 290854 -1862
rect 291474 706758 292094 711590
rect 291474 706202 291506 706758
rect 292062 706202 292094 706758
rect 291474 689134 292094 706202
rect 291474 688578 291506 689134
rect 292062 688578 292094 689134
rect 291474 653134 292094 688578
rect 291474 652578 291506 653134
rect 292062 652578 292094 653134
rect 291474 617134 292094 652578
rect 291474 616578 291506 617134
rect 292062 616578 292094 617134
rect 291474 581134 292094 616578
rect 291474 580578 291506 581134
rect 292062 580578 292094 581134
rect 291474 545134 292094 580578
rect 291474 544578 291506 545134
rect 292062 544578 292094 545134
rect 291474 509134 292094 544578
rect 291474 508578 291506 509134
rect 292062 508578 292094 509134
rect 291474 473134 292094 508578
rect 291474 472578 291506 473134
rect 292062 472578 292094 473134
rect 291474 437134 292094 472578
rect 291474 436578 291506 437134
rect 292062 436578 292094 437134
rect 291474 401134 292094 436578
rect 291474 400578 291506 401134
rect 292062 400578 292094 401134
rect 291474 365134 292094 400578
rect 291474 364578 291506 365134
rect 292062 364578 292094 365134
rect 291474 329134 292094 364578
rect 291474 328578 291506 329134
rect 292062 328578 292094 329134
rect 291474 293134 292094 328578
rect 291474 292578 291506 293134
rect 292062 292578 292094 293134
rect 291474 257134 292094 292578
rect 291474 256578 291506 257134
rect 292062 256578 292094 257134
rect 291474 221134 292094 256578
rect 291474 220578 291506 221134
rect 292062 220578 292094 221134
rect 291474 185134 292094 220578
rect 291474 184578 291506 185134
rect 292062 184578 292094 185134
rect 291474 149134 292094 184578
rect 291474 148578 291506 149134
rect 292062 148578 292094 149134
rect 291474 113134 292094 148578
rect 291474 112578 291506 113134
rect 292062 112578 292094 113134
rect 291474 77134 292094 112578
rect 291474 76578 291506 77134
rect 292062 76578 292094 77134
rect 291474 41134 292094 76578
rect 291474 40578 291506 41134
rect 292062 40578 292094 41134
rect 291474 5134 292094 40578
rect 291474 4578 291506 5134
rect 292062 4578 292094 5134
rect 291474 -2266 292094 4578
rect 291474 -2822 291506 -2266
rect 292062 -2822 292094 -2266
rect 291474 -7654 292094 -2822
rect 292714 707718 293334 711590
rect 292714 707162 292746 707718
rect 293302 707162 293334 707718
rect 292714 690374 293334 707162
rect 292714 689818 292746 690374
rect 293302 689818 293334 690374
rect 292714 654374 293334 689818
rect 292714 653818 292746 654374
rect 293302 653818 293334 654374
rect 292714 618374 293334 653818
rect 292714 617818 292746 618374
rect 293302 617818 293334 618374
rect 292714 582374 293334 617818
rect 292714 581818 292746 582374
rect 293302 581818 293334 582374
rect 292714 546374 293334 581818
rect 292714 545818 292746 546374
rect 293302 545818 293334 546374
rect 292714 510374 293334 545818
rect 292714 509818 292746 510374
rect 293302 509818 293334 510374
rect 292714 474374 293334 509818
rect 292714 473818 292746 474374
rect 293302 473818 293334 474374
rect 292714 438374 293334 473818
rect 292714 437818 292746 438374
rect 293302 437818 293334 438374
rect 292714 402374 293334 437818
rect 292714 401818 292746 402374
rect 293302 401818 293334 402374
rect 292714 366374 293334 401818
rect 292714 365818 292746 366374
rect 293302 365818 293334 366374
rect 292714 330374 293334 365818
rect 292714 329818 292746 330374
rect 293302 329818 293334 330374
rect 292714 294374 293334 329818
rect 292714 293818 292746 294374
rect 293302 293818 293334 294374
rect 292714 258374 293334 293818
rect 292714 257818 292746 258374
rect 293302 257818 293334 258374
rect 292714 222374 293334 257818
rect 292714 221818 292746 222374
rect 293302 221818 293334 222374
rect 292714 186374 293334 221818
rect 292714 185818 292746 186374
rect 293302 185818 293334 186374
rect 292714 150374 293334 185818
rect 292714 149818 292746 150374
rect 293302 149818 293334 150374
rect 292714 114374 293334 149818
rect 292714 113818 292746 114374
rect 293302 113818 293334 114374
rect 292714 78374 293334 113818
rect 292714 77818 292746 78374
rect 293302 77818 293334 78374
rect 292714 42374 293334 77818
rect 292714 41818 292746 42374
rect 293302 41818 293334 42374
rect 292714 6374 293334 41818
rect 292714 5818 292746 6374
rect 293302 5818 293334 6374
rect 292714 -3226 293334 5818
rect 292714 -3782 292746 -3226
rect 293302 -3782 293334 -3226
rect 292714 -7654 293334 -3782
rect 293954 708678 294574 711590
rect 293954 708122 293986 708678
rect 294542 708122 294574 708678
rect 293954 691614 294574 708122
rect 293954 691058 293986 691614
rect 294542 691058 294574 691614
rect 293954 655614 294574 691058
rect 293954 655058 293986 655614
rect 294542 655058 294574 655614
rect 293954 619614 294574 655058
rect 293954 619058 293986 619614
rect 294542 619058 294574 619614
rect 293954 583614 294574 619058
rect 293954 583058 293986 583614
rect 294542 583058 294574 583614
rect 293954 547614 294574 583058
rect 293954 547058 293986 547614
rect 294542 547058 294574 547614
rect 293954 511614 294574 547058
rect 293954 511058 293986 511614
rect 294542 511058 294574 511614
rect 293954 475614 294574 511058
rect 293954 475058 293986 475614
rect 294542 475058 294574 475614
rect 293954 439614 294574 475058
rect 293954 439058 293986 439614
rect 294542 439058 294574 439614
rect 293954 403614 294574 439058
rect 293954 403058 293986 403614
rect 294542 403058 294574 403614
rect 293954 367614 294574 403058
rect 293954 367058 293986 367614
rect 294542 367058 294574 367614
rect 293954 331614 294574 367058
rect 293954 331058 293986 331614
rect 294542 331058 294574 331614
rect 293954 295614 294574 331058
rect 293954 295058 293986 295614
rect 294542 295058 294574 295614
rect 293954 259614 294574 295058
rect 293954 259058 293986 259614
rect 294542 259058 294574 259614
rect 293954 223614 294574 259058
rect 293954 223058 293986 223614
rect 294542 223058 294574 223614
rect 293954 187614 294574 223058
rect 293954 187058 293986 187614
rect 294542 187058 294574 187614
rect 293954 151614 294574 187058
rect 293954 151058 293986 151614
rect 294542 151058 294574 151614
rect 293954 115614 294574 151058
rect 293954 115058 293986 115614
rect 294542 115058 294574 115614
rect 293954 79614 294574 115058
rect 293954 79058 293986 79614
rect 294542 79058 294574 79614
rect 293954 43614 294574 79058
rect 293954 43058 293986 43614
rect 294542 43058 294574 43614
rect 293954 7614 294574 43058
rect 293954 7058 293986 7614
rect 294542 7058 294574 7614
rect 293954 -4186 294574 7058
rect 293954 -4742 293986 -4186
rect 294542 -4742 294574 -4186
rect 293954 -7654 294574 -4742
rect 295194 709638 295814 711590
rect 295194 709082 295226 709638
rect 295782 709082 295814 709638
rect 295194 692854 295814 709082
rect 295194 692298 295226 692854
rect 295782 692298 295814 692854
rect 295194 656854 295814 692298
rect 295194 656298 295226 656854
rect 295782 656298 295814 656854
rect 295194 620854 295814 656298
rect 295194 620298 295226 620854
rect 295782 620298 295814 620854
rect 295194 584854 295814 620298
rect 295194 584298 295226 584854
rect 295782 584298 295814 584854
rect 295194 548854 295814 584298
rect 295194 548298 295226 548854
rect 295782 548298 295814 548854
rect 295194 512854 295814 548298
rect 295194 512298 295226 512854
rect 295782 512298 295814 512854
rect 295194 476854 295814 512298
rect 295194 476298 295226 476854
rect 295782 476298 295814 476854
rect 295194 440854 295814 476298
rect 295194 440298 295226 440854
rect 295782 440298 295814 440854
rect 295194 404854 295814 440298
rect 295194 404298 295226 404854
rect 295782 404298 295814 404854
rect 295194 368854 295814 404298
rect 295194 368298 295226 368854
rect 295782 368298 295814 368854
rect 295194 332854 295814 368298
rect 295194 332298 295226 332854
rect 295782 332298 295814 332854
rect 295194 296854 295814 332298
rect 295194 296298 295226 296854
rect 295782 296298 295814 296854
rect 295194 260854 295814 296298
rect 295194 260298 295226 260854
rect 295782 260298 295814 260854
rect 295194 224854 295814 260298
rect 295194 224298 295226 224854
rect 295782 224298 295814 224854
rect 295194 188854 295814 224298
rect 295194 188298 295226 188854
rect 295782 188298 295814 188854
rect 295194 152854 295814 188298
rect 295194 152298 295226 152854
rect 295782 152298 295814 152854
rect 295194 116854 295814 152298
rect 295194 116298 295226 116854
rect 295782 116298 295814 116854
rect 295194 80854 295814 116298
rect 295194 80298 295226 80854
rect 295782 80298 295814 80854
rect 295194 44854 295814 80298
rect 295194 44298 295226 44854
rect 295782 44298 295814 44854
rect 295194 8854 295814 44298
rect 295194 8298 295226 8854
rect 295782 8298 295814 8854
rect 295194 -5146 295814 8298
rect 295194 -5702 295226 -5146
rect 295782 -5702 295814 -5146
rect 295194 -7654 295814 -5702
rect 296434 710598 297054 711590
rect 296434 710042 296466 710598
rect 297022 710042 297054 710598
rect 296434 694094 297054 710042
rect 296434 693538 296466 694094
rect 297022 693538 297054 694094
rect 296434 658094 297054 693538
rect 296434 657538 296466 658094
rect 297022 657538 297054 658094
rect 296434 622094 297054 657538
rect 296434 621538 296466 622094
rect 297022 621538 297054 622094
rect 296434 586094 297054 621538
rect 296434 585538 296466 586094
rect 297022 585538 297054 586094
rect 296434 550094 297054 585538
rect 296434 549538 296466 550094
rect 297022 549538 297054 550094
rect 296434 514094 297054 549538
rect 296434 513538 296466 514094
rect 297022 513538 297054 514094
rect 296434 478094 297054 513538
rect 296434 477538 296466 478094
rect 297022 477538 297054 478094
rect 296434 442094 297054 477538
rect 296434 441538 296466 442094
rect 297022 441538 297054 442094
rect 296434 406094 297054 441538
rect 296434 405538 296466 406094
rect 297022 405538 297054 406094
rect 296434 370094 297054 405538
rect 296434 369538 296466 370094
rect 297022 369538 297054 370094
rect 296434 334094 297054 369538
rect 296434 333538 296466 334094
rect 297022 333538 297054 334094
rect 296434 298094 297054 333538
rect 296434 297538 296466 298094
rect 297022 297538 297054 298094
rect 296434 262094 297054 297538
rect 296434 261538 296466 262094
rect 297022 261538 297054 262094
rect 296434 226094 297054 261538
rect 296434 225538 296466 226094
rect 297022 225538 297054 226094
rect 296434 190094 297054 225538
rect 296434 189538 296466 190094
rect 297022 189538 297054 190094
rect 296434 154094 297054 189538
rect 296434 153538 296466 154094
rect 297022 153538 297054 154094
rect 296434 118094 297054 153538
rect 296434 117538 296466 118094
rect 297022 117538 297054 118094
rect 296434 82094 297054 117538
rect 296434 81538 296466 82094
rect 297022 81538 297054 82094
rect 296434 46094 297054 81538
rect 296434 45538 296466 46094
rect 297022 45538 297054 46094
rect 296434 10094 297054 45538
rect 296434 9538 296466 10094
rect 297022 9538 297054 10094
rect 296434 -6106 297054 9538
rect 296434 -6662 296466 -6106
rect 297022 -6662 297054 -6106
rect 296434 -7654 297054 -6662
rect 297674 711558 298294 711590
rect 297674 711002 297706 711558
rect 298262 711002 298294 711558
rect 297674 695334 298294 711002
rect 297674 694778 297706 695334
rect 298262 694778 298294 695334
rect 297674 659334 298294 694778
rect 297674 658778 297706 659334
rect 298262 658778 298294 659334
rect 297674 623334 298294 658778
rect 297674 622778 297706 623334
rect 298262 622778 298294 623334
rect 297674 587334 298294 622778
rect 297674 586778 297706 587334
rect 298262 586778 298294 587334
rect 297674 551334 298294 586778
rect 297674 550778 297706 551334
rect 298262 550778 298294 551334
rect 297674 515334 298294 550778
rect 297674 514778 297706 515334
rect 298262 514778 298294 515334
rect 297674 479334 298294 514778
rect 297674 478778 297706 479334
rect 298262 478778 298294 479334
rect 297674 443334 298294 478778
rect 297674 442778 297706 443334
rect 298262 442778 298294 443334
rect 297674 407334 298294 442778
rect 297674 406778 297706 407334
rect 298262 406778 298294 407334
rect 297674 371334 298294 406778
rect 297674 370778 297706 371334
rect 298262 370778 298294 371334
rect 297674 335334 298294 370778
rect 297674 334778 297706 335334
rect 298262 334778 298294 335334
rect 297674 299334 298294 334778
rect 297674 298778 297706 299334
rect 298262 298778 298294 299334
rect 297674 263334 298294 298778
rect 297674 262778 297706 263334
rect 298262 262778 298294 263334
rect 297674 227334 298294 262778
rect 297674 226778 297706 227334
rect 298262 226778 298294 227334
rect 297674 191334 298294 226778
rect 297674 190778 297706 191334
rect 298262 190778 298294 191334
rect 297674 155334 298294 190778
rect 297674 154778 297706 155334
rect 298262 154778 298294 155334
rect 297674 119334 298294 154778
rect 297674 118778 297706 119334
rect 298262 118778 298294 119334
rect 297674 83334 298294 118778
rect 297674 82778 297706 83334
rect 298262 82778 298294 83334
rect 297674 47334 298294 82778
rect 297674 46778 297706 47334
rect 298262 46778 298294 47334
rect 297674 11334 298294 46778
rect 297674 10778 297706 11334
rect 298262 10778 298294 11334
rect 297674 -7066 298294 10778
rect 297674 -7622 297706 -7066
rect 298262 -7622 298294 -7066
rect 297674 -7654 298294 -7622
rect 324994 704838 325614 711590
rect 324994 704282 325026 704838
rect 325582 704282 325614 704838
rect 324994 686654 325614 704282
rect 324994 686098 325026 686654
rect 325582 686098 325614 686654
rect 324994 650654 325614 686098
rect 324994 650098 325026 650654
rect 325582 650098 325614 650654
rect 324994 614654 325614 650098
rect 324994 614098 325026 614654
rect 325582 614098 325614 614654
rect 324994 578654 325614 614098
rect 324994 578098 325026 578654
rect 325582 578098 325614 578654
rect 324994 542654 325614 578098
rect 324994 542098 325026 542654
rect 325582 542098 325614 542654
rect 324994 506654 325614 542098
rect 324994 506098 325026 506654
rect 325582 506098 325614 506654
rect 324994 470654 325614 506098
rect 324994 470098 325026 470654
rect 325582 470098 325614 470654
rect 324994 434654 325614 470098
rect 324994 434098 325026 434654
rect 325582 434098 325614 434654
rect 324994 398654 325614 434098
rect 324994 398098 325026 398654
rect 325582 398098 325614 398654
rect 324994 362654 325614 398098
rect 324994 362098 325026 362654
rect 325582 362098 325614 362654
rect 324994 326654 325614 362098
rect 324994 326098 325026 326654
rect 325582 326098 325614 326654
rect 324994 290654 325614 326098
rect 324994 290098 325026 290654
rect 325582 290098 325614 290654
rect 324994 254654 325614 290098
rect 324994 254098 325026 254654
rect 325582 254098 325614 254654
rect 324994 218654 325614 254098
rect 324994 218098 325026 218654
rect 325582 218098 325614 218654
rect 324994 182654 325614 218098
rect 324994 182098 325026 182654
rect 325582 182098 325614 182654
rect 324994 146654 325614 182098
rect 324994 146098 325026 146654
rect 325582 146098 325614 146654
rect 324994 110654 325614 146098
rect 324994 110098 325026 110654
rect 325582 110098 325614 110654
rect 324994 74654 325614 110098
rect 324994 74098 325026 74654
rect 325582 74098 325614 74654
rect 324994 38654 325614 74098
rect 324994 38098 325026 38654
rect 325582 38098 325614 38654
rect 324994 2654 325614 38098
rect 324994 2098 325026 2654
rect 325582 2098 325614 2654
rect 324994 -346 325614 2098
rect 324994 -902 325026 -346
rect 325582 -902 325614 -346
rect 324994 -7654 325614 -902
rect 326234 705798 326854 711590
rect 326234 705242 326266 705798
rect 326822 705242 326854 705798
rect 326234 687894 326854 705242
rect 326234 687338 326266 687894
rect 326822 687338 326854 687894
rect 326234 651894 326854 687338
rect 326234 651338 326266 651894
rect 326822 651338 326854 651894
rect 326234 615894 326854 651338
rect 326234 615338 326266 615894
rect 326822 615338 326854 615894
rect 326234 579894 326854 615338
rect 326234 579338 326266 579894
rect 326822 579338 326854 579894
rect 326234 543894 326854 579338
rect 326234 543338 326266 543894
rect 326822 543338 326854 543894
rect 326234 507894 326854 543338
rect 326234 507338 326266 507894
rect 326822 507338 326854 507894
rect 326234 471894 326854 507338
rect 326234 471338 326266 471894
rect 326822 471338 326854 471894
rect 326234 435894 326854 471338
rect 326234 435338 326266 435894
rect 326822 435338 326854 435894
rect 326234 399894 326854 435338
rect 326234 399338 326266 399894
rect 326822 399338 326854 399894
rect 326234 363894 326854 399338
rect 326234 363338 326266 363894
rect 326822 363338 326854 363894
rect 326234 327894 326854 363338
rect 326234 327338 326266 327894
rect 326822 327338 326854 327894
rect 326234 291894 326854 327338
rect 326234 291338 326266 291894
rect 326822 291338 326854 291894
rect 326234 255894 326854 291338
rect 326234 255338 326266 255894
rect 326822 255338 326854 255894
rect 326234 219894 326854 255338
rect 326234 219338 326266 219894
rect 326822 219338 326854 219894
rect 326234 183894 326854 219338
rect 326234 183338 326266 183894
rect 326822 183338 326854 183894
rect 326234 147894 326854 183338
rect 326234 147338 326266 147894
rect 326822 147338 326854 147894
rect 326234 111894 326854 147338
rect 326234 111338 326266 111894
rect 326822 111338 326854 111894
rect 326234 75894 326854 111338
rect 326234 75338 326266 75894
rect 326822 75338 326854 75894
rect 326234 39894 326854 75338
rect 326234 39338 326266 39894
rect 326822 39338 326854 39894
rect 326234 3894 326854 39338
rect 326234 3338 326266 3894
rect 326822 3338 326854 3894
rect 326234 -1306 326854 3338
rect 326234 -1862 326266 -1306
rect 326822 -1862 326854 -1306
rect 326234 -7654 326854 -1862
rect 327474 706758 328094 711590
rect 327474 706202 327506 706758
rect 328062 706202 328094 706758
rect 327474 689134 328094 706202
rect 327474 688578 327506 689134
rect 328062 688578 328094 689134
rect 327474 653134 328094 688578
rect 327474 652578 327506 653134
rect 328062 652578 328094 653134
rect 327474 617134 328094 652578
rect 327474 616578 327506 617134
rect 328062 616578 328094 617134
rect 327474 581134 328094 616578
rect 327474 580578 327506 581134
rect 328062 580578 328094 581134
rect 327474 545134 328094 580578
rect 327474 544578 327506 545134
rect 328062 544578 328094 545134
rect 327474 509134 328094 544578
rect 327474 508578 327506 509134
rect 328062 508578 328094 509134
rect 327474 473134 328094 508578
rect 327474 472578 327506 473134
rect 328062 472578 328094 473134
rect 327474 437134 328094 472578
rect 327474 436578 327506 437134
rect 328062 436578 328094 437134
rect 327474 401134 328094 436578
rect 327474 400578 327506 401134
rect 328062 400578 328094 401134
rect 327474 365134 328094 400578
rect 327474 364578 327506 365134
rect 328062 364578 328094 365134
rect 327474 329134 328094 364578
rect 327474 328578 327506 329134
rect 328062 328578 328094 329134
rect 327474 293134 328094 328578
rect 327474 292578 327506 293134
rect 328062 292578 328094 293134
rect 327474 257134 328094 292578
rect 327474 256578 327506 257134
rect 328062 256578 328094 257134
rect 327474 221134 328094 256578
rect 327474 220578 327506 221134
rect 328062 220578 328094 221134
rect 327474 185134 328094 220578
rect 327474 184578 327506 185134
rect 328062 184578 328094 185134
rect 327474 149134 328094 184578
rect 327474 148578 327506 149134
rect 328062 148578 328094 149134
rect 327474 113134 328094 148578
rect 327474 112578 327506 113134
rect 328062 112578 328094 113134
rect 327474 77134 328094 112578
rect 327474 76578 327506 77134
rect 328062 76578 328094 77134
rect 327474 41134 328094 76578
rect 327474 40578 327506 41134
rect 328062 40578 328094 41134
rect 327474 5134 328094 40578
rect 327474 4578 327506 5134
rect 328062 4578 328094 5134
rect 327474 -2266 328094 4578
rect 327474 -2822 327506 -2266
rect 328062 -2822 328094 -2266
rect 327474 -7654 328094 -2822
rect 328714 707718 329334 711590
rect 328714 707162 328746 707718
rect 329302 707162 329334 707718
rect 328714 690374 329334 707162
rect 328714 689818 328746 690374
rect 329302 689818 329334 690374
rect 328714 654374 329334 689818
rect 328714 653818 328746 654374
rect 329302 653818 329334 654374
rect 328714 618374 329334 653818
rect 328714 617818 328746 618374
rect 329302 617818 329334 618374
rect 328714 582374 329334 617818
rect 328714 581818 328746 582374
rect 329302 581818 329334 582374
rect 328714 546374 329334 581818
rect 328714 545818 328746 546374
rect 329302 545818 329334 546374
rect 328714 510374 329334 545818
rect 328714 509818 328746 510374
rect 329302 509818 329334 510374
rect 328714 474374 329334 509818
rect 328714 473818 328746 474374
rect 329302 473818 329334 474374
rect 328714 438374 329334 473818
rect 328714 437818 328746 438374
rect 329302 437818 329334 438374
rect 328714 402374 329334 437818
rect 328714 401818 328746 402374
rect 329302 401818 329334 402374
rect 328714 366374 329334 401818
rect 328714 365818 328746 366374
rect 329302 365818 329334 366374
rect 328714 330374 329334 365818
rect 328714 329818 328746 330374
rect 329302 329818 329334 330374
rect 328714 294374 329334 329818
rect 328714 293818 328746 294374
rect 329302 293818 329334 294374
rect 328714 258374 329334 293818
rect 328714 257818 328746 258374
rect 329302 257818 329334 258374
rect 328714 222374 329334 257818
rect 328714 221818 328746 222374
rect 329302 221818 329334 222374
rect 328714 186374 329334 221818
rect 328714 185818 328746 186374
rect 329302 185818 329334 186374
rect 328714 150374 329334 185818
rect 328714 149818 328746 150374
rect 329302 149818 329334 150374
rect 328714 114374 329334 149818
rect 328714 113818 328746 114374
rect 329302 113818 329334 114374
rect 328714 78374 329334 113818
rect 328714 77818 328746 78374
rect 329302 77818 329334 78374
rect 328714 42374 329334 77818
rect 328714 41818 328746 42374
rect 329302 41818 329334 42374
rect 328714 6374 329334 41818
rect 328714 5818 328746 6374
rect 329302 5818 329334 6374
rect 328714 -3226 329334 5818
rect 328714 -3782 328746 -3226
rect 329302 -3782 329334 -3226
rect 328714 -7654 329334 -3782
rect 329954 708678 330574 711590
rect 329954 708122 329986 708678
rect 330542 708122 330574 708678
rect 329954 691614 330574 708122
rect 329954 691058 329986 691614
rect 330542 691058 330574 691614
rect 329954 655614 330574 691058
rect 329954 655058 329986 655614
rect 330542 655058 330574 655614
rect 329954 619614 330574 655058
rect 329954 619058 329986 619614
rect 330542 619058 330574 619614
rect 329954 583614 330574 619058
rect 329954 583058 329986 583614
rect 330542 583058 330574 583614
rect 329954 547614 330574 583058
rect 329954 547058 329986 547614
rect 330542 547058 330574 547614
rect 329954 511614 330574 547058
rect 329954 511058 329986 511614
rect 330542 511058 330574 511614
rect 329954 475614 330574 511058
rect 329954 475058 329986 475614
rect 330542 475058 330574 475614
rect 329954 439614 330574 475058
rect 329954 439058 329986 439614
rect 330542 439058 330574 439614
rect 329954 403614 330574 439058
rect 329954 403058 329986 403614
rect 330542 403058 330574 403614
rect 329954 367614 330574 403058
rect 329954 367058 329986 367614
rect 330542 367058 330574 367614
rect 329954 331614 330574 367058
rect 329954 331058 329986 331614
rect 330542 331058 330574 331614
rect 329954 295614 330574 331058
rect 329954 295058 329986 295614
rect 330542 295058 330574 295614
rect 329954 259614 330574 295058
rect 329954 259058 329986 259614
rect 330542 259058 330574 259614
rect 329954 223614 330574 259058
rect 329954 223058 329986 223614
rect 330542 223058 330574 223614
rect 329954 187614 330574 223058
rect 329954 187058 329986 187614
rect 330542 187058 330574 187614
rect 329954 151614 330574 187058
rect 329954 151058 329986 151614
rect 330542 151058 330574 151614
rect 329954 115614 330574 151058
rect 329954 115058 329986 115614
rect 330542 115058 330574 115614
rect 329954 79614 330574 115058
rect 329954 79058 329986 79614
rect 330542 79058 330574 79614
rect 329954 43614 330574 79058
rect 329954 43058 329986 43614
rect 330542 43058 330574 43614
rect 329954 7614 330574 43058
rect 329954 7058 329986 7614
rect 330542 7058 330574 7614
rect 329954 -4186 330574 7058
rect 329954 -4742 329986 -4186
rect 330542 -4742 330574 -4186
rect 329954 -7654 330574 -4742
rect 331194 709638 331814 711590
rect 331194 709082 331226 709638
rect 331782 709082 331814 709638
rect 331194 692854 331814 709082
rect 331194 692298 331226 692854
rect 331782 692298 331814 692854
rect 331194 656854 331814 692298
rect 331194 656298 331226 656854
rect 331782 656298 331814 656854
rect 331194 620854 331814 656298
rect 331194 620298 331226 620854
rect 331782 620298 331814 620854
rect 331194 584854 331814 620298
rect 331194 584298 331226 584854
rect 331782 584298 331814 584854
rect 331194 548854 331814 584298
rect 331194 548298 331226 548854
rect 331782 548298 331814 548854
rect 331194 512854 331814 548298
rect 331194 512298 331226 512854
rect 331782 512298 331814 512854
rect 331194 476854 331814 512298
rect 331194 476298 331226 476854
rect 331782 476298 331814 476854
rect 331194 440854 331814 476298
rect 331194 440298 331226 440854
rect 331782 440298 331814 440854
rect 331194 404854 331814 440298
rect 331194 404298 331226 404854
rect 331782 404298 331814 404854
rect 331194 368854 331814 404298
rect 331194 368298 331226 368854
rect 331782 368298 331814 368854
rect 331194 332854 331814 368298
rect 331194 332298 331226 332854
rect 331782 332298 331814 332854
rect 331194 296854 331814 332298
rect 331194 296298 331226 296854
rect 331782 296298 331814 296854
rect 331194 260854 331814 296298
rect 331194 260298 331226 260854
rect 331782 260298 331814 260854
rect 331194 224854 331814 260298
rect 331194 224298 331226 224854
rect 331782 224298 331814 224854
rect 331194 188854 331814 224298
rect 331194 188298 331226 188854
rect 331782 188298 331814 188854
rect 331194 152854 331814 188298
rect 331194 152298 331226 152854
rect 331782 152298 331814 152854
rect 331194 116854 331814 152298
rect 331194 116298 331226 116854
rect 331782 116298 331814 116854
rect 331194 80854 331814 116298
rect 331194 80298 331226 80854
rect 331782 80298 331814 80854
rect 331194 44854 331814 80298
rect 331194 44298 331226 44854
rect 331782 44298 331814 44854
rect 331194 8854 331814 44298
rect 331194 8298 331226 8854
rect 331782 8298 331814 8854
rect 331194 -5146 331814 8298
rect 331194 -5702 331226 -5146
rect 331782 -5702 331814 -5146
rect 331194 -7654 331814 -5702
rect 332434 710598 333054 711590
rect 332434 710042 332466 710598
rect 333022 710042 333054 710598
rect 332434 694094 333054 710042
rect 332434 693538 332466 694094
rect 333022 693538 333054 694094
rect 332434 658094 333054 693538
rect 332434 657538 332466 658094
rect 333022 657538 333054 658094
rect 332434 622094 333054 657538
rect 332434 621538 332466 622094
rect 333022 621538 333054 622094
rect 332434 586094 333054 621538
rect 332434 585538 332466 586094
rect 333022 585538 333054 586094
rect 332434 550094 333054 585538
rect 332434 549538 332466 550094
rect 333022 549538 333054 550094
rect 332434 514094 333054 549538
rect 332434 513538 332466 514094
rect 333022 513538 333054 514094
rect 332434 478094 333054 513538
rect 332434 477538 332466 478094
rect 333022 477538 333054 478094
rect 332434 442094 333054 477538
rect 332434 441538 332466 442094
rect 333022 441538 333054 442094
rect 332434 406094 333054 441538
rect 332434 405538 332466 406094
rect 333022 405538 333054 406094
rect 332434 370094 333054 405538
rect 332434 369538 332466 370094
rect 333022 369538 333054 370094
rect 332434 334094 333054 369538
rect 332434 333538 332466 334094
rect 333022 333538 333054 334094
rect 332434 298094 333054 333538
rect 332434 297538 332466 298094
rect 333022 297538 333054 298094
rect 332434 262094 333054 297538
rect 332434 261538 332466 262094
rect 333022 261538 333054 262094
rect 332434 226094 333054 261538
rect 332434 225538 332466 226094
rect 333022 225538 333054 226094
rect 332434 190094 333054 225538
rect 332434 189538 332466 190094
rect 333022 189538 333054 190094
rect 332434 154094 333054 189538
rect 332434 153538 332466 154094
rect 333022 153538 333054 154094
rect 332434 118094 333054 153538
rect 332434 117538 332466 118094
rect 333022 117538 333054 118094
rect 332434 82094 333054 117538
rect 332434 81538 332466 82094
rect 333022 81538 333054 82094
rect 332434 46094 333054 81538
rect 332434 45538 332466 46094
rect 333022 45538 333054 46094
rect 332434 10094 333054 45538
rect 332434 9538 332466 10094
rect 333022 9538 333054 10094
rect 332434 -6106 333054 9538
rect 332434 -6662 332466 -6106
rect 333022 -6662 333054 -6106
rect 332434 -7654 333054 -6662
rect 333674 711558 334294 711590
rect 333674 711002 333706 711558
rect 334262 711002 334294 711558
rect 333674 695334 334294 711002
rect 333674 694778 333706 695334
rect 334262 694778 334294 695334
rect 333674 659334 334294 694778
rect 333674 658778 333706 659334
rect 334262 658778 334294 659334
rect 333674 623334 334294 658778
rect 333674 622778 333706 623334
rect 334262 622778 334294 623334
rect 333674 587334 334294 622778
rect 333674 586778 333706 587334
rect 334262 586778 334294 587334
rect 333674 551334 334294 586778
rect 333674 550778 333706 551334
rect 334262 550778 334294 551334
rect 333674 515334 334294 550778
rect 333674 514778 333706 515334
rect 334262 514778 334294 515334
rect 333674 479334 334294 514778
rect 333674 478778 333706 479334
rect 334262 478778 334294 479334
rect 333674 443334 334294 478778
rect 333674 442778 333706 443334
rect 334262 442778 334294 443334
rect 333674 407334 334294 442778
rect 333674 406778 333706 407334
rect 334262 406778 334294 407334
rect 333674 371334 334294 406778
rect 333674 370778 333706 371334
rect 334262 370778 334294 371334
rect 333674 335334 334294 370778
rect 333674 334778 333706 335334
rect 334262 334778 334294 335334
rect 333674 299334 334294 334778
rect 333674 298778 333706 299334
rect 334262 298778 334294 299334
rect 333674 263334 334294 298778
rect 333674 262778 333706 263334
rect 334262 262778 334294 263334
rect 333674 227334 334294 262778
rect 333674 226778 333706 227334
rect 334262 226778 334294 227334
rect 333674 191334 334294 226778
rect 333674 190778 333706 191334
rect 334262 190778 334294 191334
rect 333674 155334 334294 190778
rect 333674 154778 333706 155334
rect 334262 154778 334294 155334
rect 333674 119334 334294 154778
rect 333674 118778 333706 119334
rect 334262 118778 334294 119334
rect 333674 83334 334294 118778
rect 333674 82778 333706 83334
rect 334262 82778 334294 83334
rect 333674 47334 334294 82778
rect 333674 46778 333706 47334
rect 334262 46778 334294 47334
rect 333674 11334 334294 46778
rect 333674 10778 333706 11334
rect 334262 10778 334294 11334
rect 333674 -7066 334294 10778
rect 333674 -7622 333706 -7066
rect 334262 -7622 334294 -7066
rect 333674 -7654 334294 -7622
rect 360994 704838 361614 711590
rect 360994 704282 361026 704838
rect 361582 704282 361614 704838
rect 360994 686654 361614 704282
rect 360994 686098 361026 686654
rect 361582 686098 361614 686654
rect 360994 650654 361614 686098
rect 360994 650098 361026 650654
rect 361582 650098 361614 650654
rect 360994 614654 361614 650098
rect 360994 614098 361026 614654
rect 361582 614098 361614 614654
rect 360994 578654 361614 614098
rect 360994 578098 361026 578654
rect 361582 578098 361614 578654
rect 360994 542654 361614 578098
rect 360994 542098 361026 542654
rect 361582 542098 361614 542654
rect 360994 506654 361614 542098
rect 360994 506098 361026 506654
rect 361582 506098 361614 506654
rect 360994 470654 361614 506098
rect 360994 470098 361026 470654
rect 361582 470098 361614 470654
rect 360994 434654 361614 470098
rect 360994 434098 361026 434654
rect 361582 434098 361614 434654
rect 360994 398654 361614 434098
rect 360994 398098 361026 398654
rect 361582 398098 361614 398654
rect 360994 362654 361614 398098
rect 360994 362098 361026 362654
rect 361582 362098 361614 362654
rect 360994 326654 361614 362098
rect 360994 326098 361026 326654
rect 361582 326098 361614 326654
rect 360994 290654 361614 326098
rect 360994 290098 361026 290654
rect 361582 290098 361614 290654
rect 360994 254654 361614 290098
rect 360994 254098 361026 254654
rect 361582 254098 361614 254654
rect 360994 218654 361614 254098
rect 360994 218098 361026 218654
rect 361582 218098 361614 218654
rect 360994 182654 361614 218098
rect 360994 182098 361026 182654
rect 361582 182098 361614 182654
rect 360994 146654 361614 182098
rect 360994 146098 361026 146654
rect 361582 146098 361614 146654
rect 360994 110654 361614 146098
rect 360994 110098 361026 110654
rect 361582 110098 361614 110654
rect 360994 74654 361614 110098
rect 360994 74098 361026 74654
rect 361582 74098 361614 74654
rect 360994 38654 361614 74098
rect 360994 38098 361026 38654
rect 361582 38098 361614 38654
rect 360994 2654 361614 38098
rect 360994 2098 361026 2654
rect 361582 2098 361614 2654
rect 360994 -346 361614 2098
rect 360994 -902 361026 -346
rect 361582 -902 361614 -346
rect 360994 -7654 361614 -902
rect 362234 705798 362854 711590
rect 362234 705242 362266 705798
rect 362822 705242 362854 705798
rect 362234 687894 362854 705242
rect 362234 687338 362266 687894
rect 362822 687338 362854 687894
rect 362234 651894 362854 687338
rect 362234 651338 362266 651894
rect 362822 651338 362854 651894
rect 362234 615894 362854 651338
rect 362234 615338 362266 615894
rect 362822 615338 362854 615894
rect 362234 579894 362854 615338
rect 362234 579338 362266 579894
rect 362822 579338 362854 579894
rect 362234 543894 362854 579338
rect 362234 543338 362266 543894
rect 362822 543338 362854 543894
rect 362234 507894 362854 543338
rect 362234 507338 362266 507894
rect 362822 507338 362854 507894
rect 362234 471894 362854 507338
rect 362234 471338 362266 471894
rect 362822 471338 362854 471894
rect 362234 435894 362854 471338
rect 362234 435338 362266 435894
rect 362822 435338 362854 435894
rect 362234 399894 362854 435338
rect 362234 399338 362266 399894
rect 362822 399338 362854 399894
rect 362234 363894 362854 399338
rect 362234 363338 362266 363894
rect 362822 363338 362854 363894
rect 362234 327894 362854 363338
rect 362234 327338 362266 327894
rect 362822 327338 362854 327894
rect 362234 291894 362854 327338
rect 362234 291338 362266 291894
rect 362822 291338 362854 291894
rect 362234 255894 362854 291338
rect 362234 255338 362266 255894
rect 362822 255338 362854 255894
rect 362234 219894 362854 255338
rect 362234 219338 362266 219894
rect 362822 219338 362854 219894
rect 362234 183894 362854 219338
rect 362234 183338 362266 183894
rect 362822 183338 362854 183894
rect 362234 147894 362854 183338
rect 362234 147338 362266 147894
rect 362822 147338 362854 147894
rect 362234 111894 362854 147338
rect 362234 111338 362266 111894
rect 362822 111338 362854 111894
rect 362234 75894 362854 111338
rect 362234 75338 362266 75894
rect 362822 75338 362854 75894
rect 362234 39894 362854 75338
rect 362234 39338 362266 39894
rect 362822 39338 362854 39894
rect 362234 3894 362854 39338
rect 362234 3338 362266 3894
rect 362822 3338 362854 3894
rect 362234 -1306 362854 3338
rect 362234 -1862 362266 -1306
rect 362822 -1862 362854 -1306
rect 362234 -7654 362854 -1862
rect 363474 706758 364094 711590
rect 363474 706202 363506 706758
rect 364062 706202 364094 706758
rect 363474 689134 364094 706202
rect 363474 688578 363506 689134
rect 364062 688578 364094 689134
rect 363474 653134 364094 688578
rect 363474 652578 363506 653134
rect 364062 652578 364094 653134
rect 363474 617134 364094 652578
rect 363474 616578 363506 617134
rect 364062 616578 364094 617134
rect 363474 581134 364094 616578
rect 363474 580578 363506 581134
rect 364062 580578 364094 581134
rect 363474 545134 364094 580578
rect 363474 544578 363506 545134
rect 364062 544578 364094 545134
rect 363474 509134 364094 544578
rect 363474 508578 363506 509134
rect 364062 508578 364094 509134
rect 363474 473134 364094 508578
rect 363474 472578 363506 473134
rect 364062 472578 364094 473134
rect 363474 437134 364094 472578
rect 363474 436578 363506 437134
rect 364062 436578 364094 437134
rect 363474 401134 364094 436578
rect 363474 400578 363506 401134
rect 364062 400578 364094 401134
rect 363474 365134 364094 400578
rect 363474 364578 363506 365134
rect 364062 364578 364094 365134
rect 363474 329134 364094 364578
rect 363474 328578 363506 329134
rect 364062 328578 364094 329134
rect 363474 293134 364094 328578
rect 363474 292578 363506 293134
rect 364062 292578 364094 293134
rect 363474 257134 364094 292578
rect 363474 256578 363506 257134
rect 364062 256578 364094 257134
rect 363474 221134 364094 256578
rect 363474 220578 363506 221134
rect 364062 220578 364094 221134
rect 363474 185134 364094 220578
rect 363474 184578 363506 185134
rect 364062 184578 364094 185134
rect 363474 149134 364094 184578
rect 363474 148578 363506 149134
rect 364062 148578 364094 149134
rect 363474 113134 364094 148578
rect 363474 112578 363506 113134
rect 364062 112578 364094 113134
rect 363474 77134 364094 112578
rect 363474 76578 363506 77134
rect 364062 76578 364094 77134
rect 363474 41134 364094 76578
rect 363474 40578 363506 41134
rect 364062 40578 364094 41134
rect 363474 5134 364094 40578
rect 363474 4578 363506 5134
rect 364062 4578 364094 5134
rect 363474 -2266 364094 4578
rect 363474 -2822 363506 -2266
rect 364062 -2822 364094 -2266
rect 363474 -7654 364094 -2822
rect 364714 707718 365334 711590
rect 364714 707162 364746 707718
rect 365302 707162 365334 707718
rect 364714 690374 365334 707162
rect 364714 689818 364746 690374
rect 365302 689818 365334 690374
rect 364714 654374 365334 689818
rect 364714 653818 364746 654374
rect 365302 653818 365334 654374
rect 364714 618374 365334 653818
rect 364714 617818 364746 618374
rect 365302 617818 365334 618374
rect 364714 582374 365334 617818
rect 364714 581818 364746 582374
rect 365302 581818 365334 582374
rect 364714 546374 365334 581818
rect 364714 545818 364746 546374
rect 365302 545818 365334 546374
rect 364714 510374 365334 545818
rect 364714 509818 364746 510374
rect 365302 509818 365334 510374
rect 364714 474374 365334 509818
rect 364714 473818 364746 474374
rect 365302 473818 365334 474374
rect 364714 438374 365334 473818
rect 364714 437818 364746 438374
rect 365302 437818 365334 438374
rect 364714 402374 365334 437818
rect 364714 401818 364746 402374
rect 365302 401818 365334 402374
rect 364714 366374 365334 401818
rect 364714 365818 364746 366374
rect 365302 365818 365334 366374
rect 364714 330374 365334 365818
rect 364714 329818 364746 330374
rect 365302 329818 365334 330374
rect 364714 294374 365334 329818
rect 364714 293818 364746 294374
rect 365302 293818 365334 294374
rect 364714 258374 365334 293818
rect 364714 257818 364746 258374
rect 365302 257818 365334 258374
rect 364714 222374 365334 257818
rect 364714 221818 364746 222374
rect 365302 221818 365334 222374
rect 364714 186374 365334 221818
rect 364714 185818 364746 186374
rect 365302 185818 365334 186374
rect 364714 150374 365334 185818
rect 364714 149818 364746 150374
rect 365302 149818 365334 150374
rect 364714 114374 365334 149818
rect 364714 113818 364746 114374
rect 365302 113818 365334 114374
rect 364714 78374 365334 113818
rect 364714 77818 364746 78374
rect 365302 77818 365334 78374
rect 364714 42374 365334 77818
rect 364714 41818 364746 42374
rect 365302 41818 365334 42374
rect 364714 6374 365334 41818
rect 364714 5818 364746 6374
rect 365302 5818 365334 6374
rect 364714 -3226 365334 5818
rect 364714 -3782 364746 -3226
rect 365302 -3782 365334 -3226
rect 364714 -7654 365334 -3782
rect 365954 708678 366574 711590
rect 365954 708122 365986 708678
rect 366542 708122 366574 708678
rect 365954 691614 366574 708122
rect 365954 691058 365986 691614
rect 366542 691058 366574 691614
rect 365954 655614 366574 691058
rect 365954 655058 365986 655614
rect 366542 655058 366574 655614
rect 365954 619614 366574 655058
rect 365954 619058 365986 619614
rect 366542 619058 366574 619614
rect 365954 583614 366574 619058
rect 365954 583058 365986 583614
rect 366542 583058 366574 583614
rect 365954 547614 366574 583058
rect 365954 547058 365986 547614
rect 366542 547058 366574 547614
rect 365954 511614 366574 547058
rect 365954 511058 365986 511614
rect 366542 511058 366574 511614
rect 365954 475614 366574 511058
rect 365954 475058 365986 475614
rect 366542 475058 366574 475614
rect 365954 439614 366574 475058
rect 365954 439058 365986 439614
rect 366542 439058 366574 439614
rect 365954 403614 366574 439058
rect 365954 403058 365986 403614
rect 366542 403058 366574 403614
rect 365954 367614 366574 403058
rect 365954 367058 365986 367614
rect 366542 367058 366574 367614
rect 365954 331614 366574 367058
rect 365954 331058 365986 331614
rect 366542 331058 366574 331614
rect 365954 295614 366574 331058
rect 365954 295058 365986 295614
rect 366542 295058 366574 295614
rect 365954 259614 366574 295058
rect 365954 259058 365986 259614
rect 366542 259058 366574 259614
rect 365954 223614 366574 259058
rect 365954 223058 365986 223614
rect 366542 223058 366574 223614
rect 365954 187614 366574 223058
rect 365954 187058 365986 187614
rect 366542 187058 366574 187614
rect 365954 151614 366574 187058
rect 365954 151058 365986 151614
rect 366542 151058 366574 151614
rect 365954 115614 366574 151058
rect 365954 115058 365986 115614
rect 366542 115058 366574 115614
rect 365954 79614 366574 115058
rect 365954 79058 365986 79614
rect 366542 79058 366574 79614
rect 365954 43614 366574 79058
rect 365954 43058 365986 43614
rect 366542 43058 366574 43614
rect 365954 7614 366574 43058
rect 365954 7058 365986 7614
rect 366542 7058 366574 7614
rect 365954 -4186 366574 7058
rect 365954 -4742 365986 -4186
rect 366542 -4742 366574 -4186
rect 365954 -7654 366574 -4742
rect 367194 709638 367814 711590
rect 367194 709082 367226 709638
rect 367782 709082 367814 709638
rect 367194 692854 367814 709082
rect 367194 692298 367226 692854
rect 367782 692298 367814 692854
rect 367194 656854 367814 692298
rect 367194 656298 367226 656854
rect 367782 656298 367814 656854
rect 367194 620854 367814 656298
rect 367194 620298 367226 620854
rect 367782 620298 367814 620854
rect 367194 584854 367814 620298
rect 367194 584298 367226 584854
rect 367782 584298 367814 584854
rect 367194 548854 367814 584298
rect 367194 548298 367226 548854
rect 367782 548298 367814 548854
rect 367194 512854 367814 548298
rect 367194 512298 367226 512854
rect 367782 512298 367814 512854
rect 367194 476854 367814 512298
rect 367194 476298 367226 476854
rect 367782 476298 367814 476854
rect 367194 440854 367814 476298
rect 367194 440298 367226 440854
rect 367782 440298 367814 440854
rect 367194 404854 367814 440298
rect 367194 404298 367226 404854
rect 367782 404298 367814 404854
rect 367194 368854 367814 404298
rect 367194 368298 367226 368854
rect 367782 368298 367814 368854
rect 367194 332854 367814 368298
rect 367194 332298 367226 332854
rect 367782 332298 367814 332854
rect 367194 296854 367814 332298
rect 367194 296298 367226 296854
rect 367782 296298 367814 296854
rect 367194 260854 367814 296298
rect 367194 260298 367226 260854
rect 367782 260298 367814 260854
rect 367194 224854 367814 260298
rect 367194 224298 367226 224854
rect 367782 224298 367814 224854
rect 367194 188854 367814 224298
rect 367194 188298 367226 188854
rect 367782 188298 367814 188854
rect 367194 152854 367814 188298
rect 367194 152298 367226 152854
rect 367782 152298 367814 152854
rect 367194 116854 367814 152298
rect 367194 116298 367226 116854
rect 367782 116298 367814 116854
rect 367194 80854 367814 116298
rect 367194 80298 367226 80854
rect 367782 80298 367814 80854
rect 367194 44854 367814 80298
rect 367194 44298 367226 44854
rect 367782 44298 367814 44854
rect 367194 8854 367814 44298
rect 367194 8298 367226 8854
rect 367782 8298 367814 8854
rect 367194 -5146 367814 8298
rect 367194 -5702 367226 -5146
rect 367782 -5702 367814 -5146
rect 367194 -7654 367814 -5702
rect 368434 710598 369054 711590
rect 368434 710042 368466 710598
rect 369022 710042 369054 710598
rect 368434 694094 369054 710042
rect 368434 693538 368466 694094
rect 369022 693538 369054 694094
rect 368434 658094 369054 693538
rect 368434 657538 368466 658094
rect 369022 657538 369054 658094
rect 368434 622094 369054 657538
rect 368434 621538 368466 622094
rect 369022 621538 369054 622094
rect 368434 586094 369054 621538
rect 368434 585538 368466 586094
rect 369022 585538 369054 586094
rect 368434 550094 369054 585538
rect 368434 549538 368466 550094
rect 369022 549538 369054 550094
rect 368434 514094 369054 549538
rect 368434 513538 368466 514094
rect 369022 513538 369054 514094
rect 368434 478094 369054 513538
rect 368434 477538 368466 478094
rect 369022 477538 369054 478094
rect 368434 442094 369054 477538
rect 368434 441538 368466 442094
rect 369022 441538 369054 442094
rect 368434 406094 369054 441538
rect 368434 405538 368466 406094
rect 369022 405538 369054 406094
rect 368434 370094 369054 405538
rect 368434 369538 368466 370094
rect 369022 369538 369054 370094
rect 368434 334094 369054 369538
rect 368434 333538 368466 334094
rect 369022 333538 369054 334094
rect 368434 298094 369054 333538
rect 368434 297538 368466 298094
rect 369022 297538 369054 298094
rect 368434 262094 369054 297538
rect 368434 261538 368466 262094
rect 369022 261538 369054 262094
rect 368434 226094 369054 261538
rect 368434 225538 368466 226094
rect 369022 225538 369054 226094
rect 368434 190094 369054 225538
rect 368434 189538 368466 190094
rect 369022 189538 369054 190094
rect 368434 154094 369054 189538
rect 368434 153538 368466 154094
rect 369022 153538 369054 154094
rect 368434 118094 369054 153538
rect 368434 117538 368466 118094
rect 369022 117538 369054 118094
rect 368434 82094 369054 117538
rect 368434 81538 368466 82094
rect 369022 81538 369054 82094
rect 368434 46094 369054 81538
rect 368434 45538 368466 46094
rect 369022 45538 369054 46094
rect 368434 10094 369054 45538
rect 368434 9538 368466 10094
rect 369022 9538 369054 10094
rect 368434 -6106 369054 9538
rect 368434 -6662 368466 -6106
rect 369022 -6662 369054 -6106
rect 368434 -7654 369054 -6662
rect 369674 711558 370294 711590
rect 369674 711002 369706 711558
rect 370262 711002 370294 711558
rect 369674 695334 370294 711002
rect 369674 694778 369706 695334
rect 370262 694778 370294 695334
rect 369674 659334 370294 694778
rect 369674 658778 369706 659334
rect 370262 658778 370294 659334
rect 369674 623334 370294 658778
rect 369674 622778 369706 623334
rect 370262 622778 370294 623334
rect 369674 587334 370294 622778
rect 369674 586778 369706 587334
rect 370262 586778 370294 587334
rect 369674 551334 370294 586778
rect 369674 550778 369706 551334
rect 370262 550778 370294 551334
rect 369674 515334 370294 550778
rect 369674 514778 369706 515334
rect 370262 514778 370294 515334
rect 369674 479334 370294 514778
rect 369674 478778 369706 479334
rect 370262 478778 370294 479334
rect 369674 443334 370294 478778
rect 369674 442778 369706 443334
rect 370262 442778 370294 443334
rect 369674 407334 370294 442778
rect 369674 406778 369706 407334
rect 370262 406778 370294 407334
rect 369674 371334 370294 406778
rect 369674 370778 369706 371334
rect 370262 370778 370294 371334
rect 369674 335334 370294 370778
rect 369674 334778 369706 335334
rect 370262 334778 370294 335334
rect 369674 299334 370294 334778
rect 369674 298778 369706 299334
rect 370262 298778 370294 299334
rect 369674 263334 370294 298778
rect 369674 262778 369706 263334
rect 370262 262778 370294 263334
rect 369674 227334 370294 262778
rect 369674 226778 369706 227334
rect 370262 226778 370294 227334
rect 369674 191334 370294 226778
rect 369674 190778 369706 191334
rect 370262 190778 370294 191334
rect 369674 155334 370294 190778
rect 369674 154778 369706 155334
rect 370262 154778 370294 155334
rect 369674 119334 370294 154778
rect 369674 118778 369706 119334
rect 370262 118778 370294 119334
rect 369674 83334 370294 118778
rect 369674 82778 369706 83334
rect 370262 82778 370294 83334
rect 369674 47334 370294 82778
rect 369674 46778 369706 47334
rect 370262 46778 370294 47334
rect 369674 11334 370294 46778
rect 369674 10778 369706 11334
rect 370262 10778 370294 11334
rect 369674 -7066 370294 10778
rect 369674 -7622 369706 -7066
rect 370262 -7622 370294 -7066
rect 369674 -7654 370294 -7622
rect 396994 704838 397614 711590
rect 396994 704282 397026 704838
rect 397582 704282 397614 704838
rect 396994 686654 397614 704282
rect 396994 686098 397026 686654
rect 397582 686098 397614 686654
rect 396994 650654 397614 686098
rect 396994 650098 397026 650654
rect 397582 650098 397614 650654
rect 396994 614654 397614 650098
rect 396994 614098 397026 614654
rect 397582 614098 397614 614654
rect 396994 578654 397614 614098
rect 396994 578098 397026 578654
rect 397582 578098 397614 578654
rect 396994 542654 397614 578098
rect 396994 542098 397026 542654
rect 397582 542098 397614 542654
rect 396994 506654 397614 542098
rect 396994 506098 397026 506654
rect 397582 506098 397614 506654
rect 396994 470654 397614 506098
rect 396994 470098 397026 470654
rect 397582 470098 397614 470654
rect 396994 434654 397614 470098
rect 396994 434098 397026 434654
rect 397582 434098 397614 434654
rect 396994 398654 397614 434098
rect 396994 398098 397026 398654
rect 397582 398098 397614 398654
rect 396994 362654 397614 398098
rect 396994 362098 397026 362654
rect 397582 362098 397614 362654
rect 396994 326654 397614 362098
rect 396994 326098 397026 326654
rect 397582 326098 397614 326654
rect 396994 290654 397614 326098
rect 396994 290098 397026 290654
rect 397582 290098 397614 290654
rect 396994 254654 397614 290098
rect 396994 254098 397026 254654
rect 397582 254098 397614 254654
rect 396994 218654 397614 254098
rect 396994 218098 397026 218654
rect 397582 218098 397614 218654
rect 396994 182654 397614 218098
rect 396994 182098 397026 182654
rect 397582 182098 397614 182654
rect 396994 146654 397614 182098
rect 396994 146098 397026 146654
rect 397582 146098 397614 146654
rect 396994 110654 397614 146098
rect 396994 110098 397026 110654
rect 397582 110098 397614 110654
rect 396994 74654 397614 110098
rect 396994 74098 397026 74654
rect 397582 74098 397614 74654
rect 396994 38654 397614 74098
rect 396994 38098 397026 38654
rect 397582 38098 397614 38654
rect 396994 2654 397614 38098
rect 396994 2098 397026 2654
rect 397582 2098 397614 2654
rect 396994 -346 397614 2098
rect 396994 -902 397026 -346
rect 397582 -902 397614 -346
rect 396994 -7654 397614 -902
rect 398234 705798 398854 711590
rect 398234 705242 398266 705798
rect 398822 705242 398854 705798
rect 398234 687894 398854 705242
rect 398234 687338 398266 687894
rect 398822 687338 398854 687894
rect 398234 651894 398854 687338
rect 398234 651338 398266 651894
rect 398822 651338 398854 651894
rect 398234 615894 398854 651338
rect 398234 615338 398266 615894
rect 398822 615338 398854 615894
rect 398234 579894 398854 615338
rect 398234 579338 398266 579894
rect 398822 579338 398854 579894
rect 398234 543894 398854 579338
rect 398234 543338 398266 543894
rect 398822 543338 398854 543894
rect 398234 507894 398854 543338
rect 398234 507338 398266 507894
rect 398822 507338 398854 507894
rect 398234 471894 398854 507338
rect 398234 471338 398266 471894
rect 398822 471338 398854 471894
rect 398234 435894 398854 471338
rect 398234 435338 398266 435894
rect 398822 435338 398854 435894
rect 398234 399894 398854 435338
rect 398234 399338 398266 399894
rect 398822 399338 398854 399894
rect 398234 363894 398854 399338
rect 398234 363338 398266 363894
rect 398822 363338 398854 363894
rect 398234 327894 398854 363338
rect 398234 327338 398266 327894
rect 398822 327338 398854 327894
rect 398234 291894 398854 327338
rect 398234 291338 398266 291894
rect 398822 291338 398854 291894
rect 398234 255894 398854 291338
rect 398234 255338 398266 255894
rect 398822 255338 398854 255894
rect 398234 219894 398854 255338
rect 398234 219338 398266 219894
rect 398822 219338 398854 219894
rect 398234 183894 398854 219338
rect 398234 183338 398266 183894
rect 398822 183338 398854 183894
rect 398234 147894 398854 183338
rect 398234 147338 398266 147894
rect 398822 147338 398854 147894
rect 398234 111894 398854 147338
rect 398234 111338 398266 111894
rect 398822 111338 398854 111894
rect 398234 75894 398854 111338
rect 398234 75338 398266 75894
rect 398822 75338 398854 75894
rect 398234 39894 398854 75338
rect 398234 39338 398266 39894
rect 398822 39338 398854 39894
rect 398234 3894 398854 39338
rect 398234 3338 398266 3894
rect 398822 3338 398854 3894
rect 398234 -1306 398854 3338
rect 398234 -1862 398266 -1306
rect 398822 -1862 398854 -1306
rect 398234 -7654 398854 -1862
rect 399474 706758 400094 711590
rect 399474 706202 399506 706758
rect 400062 706202 400094 706758
rect 399474 689134 400094 706202
rect 399474 688578 399506 689134
rect 400062 688578 400094 689134
rect 399474 653134 400094 688578
rect 399474 652578 399506 653134
rect 400062 652578 400094 653134
rect 399474 617134 400094 652578
rect 399474 616578 399506 617134
rect 400062 616578 400094 617134
rect 399474 581134 400094 616578
rect 399474 580578 399506 581134
rect 400062 580578 400094 581134
rect 399474 545134 400094 580578
rect 399474 544578 399506 545134
rect 400062 544578 400094 545134
rect 399474 509134 400094 544578
rect 399474 508578 399506 509134
rect 400062 508578 400094 509134
rect 399474 473134 400094 508578
rect 399474 472578 399506 473134
rect 400062 472578 400094 473134
rect 399474 437134 400094 472578
rect 399474 436578 399506 437134
rect 400062 436578 400094 437134
rect 399474 401134 400094 436578
rect 399474 400578 399506 401134
rect 400062 400578 400094 401134
rect 399474 365134 400094 400578
rect 399474 364578 399506 365134
rect 400062 364578 400094 365134
rect 399474 329134 400094 364578
rect 399474 328578 399506 329134
rect 400062 328578 400094 329134
rect 399474 293134 400094 328578
rect 399474 292578 399506 293134
rect 400062 292578 400094 293134
rect 399474 257134 400094 292578
rect 399474 256578 399506 257134
rect 400062 256578 400094 257134
rect 399474 221134 400094 256578
rect 399474 220578 399506 221134
rect 400062 220578 400094 221134
rect 399474 185134 400094 220578
rect 399474 184578 399506 185134
rect 400062 184578 400094 185134
rect 399474 149134 400094 184578
rect 399474 148578 399506 149134
rect 400062 148578 400094 149134
rect 399474 113134 400094 148578
rect 399474 112578 399506 113134
rect 400062 112578 400094 113134
rect 399474 77134 400094 112578
rect 399474 76578 399506 77134
rect 400062 76578 400094 77134
rect 399474 41134 400094 76578
rect 399474 40578 399506 41134
rect 400062 40578 400094 41134
rect 399474 5134 400094 40578
rect 399474 4578 399506 5134
rect 400062 4578 400094 5134
rect 399474 -2266 400094 4578
rect 399474 -2822 399506 -2266
rect 400062 -2822 400094 -2266
rect 399474 -7654 400094 -2822
rect 400714 707718 401334 711590
rect 400714 707162 400746 707718
rect 401302 707162 401334 707718
rect 400714 690374 401334 707162
rect 400714 689818 400746 690374
rect 401302 689818 401334 690374
rect 400714 654374 401334 689818
rect 400714 653818 400746 654374
rect 401302 653818 401334 654374
rect 400714 618374 401334 653818
rect 400714 617818 400746 618374
rect 401302 617818 401334 618374
rect 400714 582374 401334 617818
rect 400714 581818 400746 582374
rect 401302 581818 401334 582374
rect 400714 546374 401334 581818
rect 400714 545818 400746 546374
rect 401302 545818 401334 546374
rect 400714 510374 401334 545818
rect 400714 509818 400746 510374
rect 401302 509818 401334 510374
rect 400714 474374 401334 509818
rect 400714 473818 400746 474374
rect 401302 473818 401334 474374
rect 400714 438374 401334 473818
rect 400714 437818 400746 438374
rect 401302 437818 401334 438374
rect 400714 402374 401334 437818
rect 400714 401818 400746 402374
rect 401302 401818 401334 402374
rect 400714 366374 401334 401818
rect 400714 365818 400746 366374
rect 401302 365818 401334 366374
rect 400714 330374 401334 365818
rect 400714 329818 400746 330374
rect 401302 329818 401334 330374
rect 400714 294374 401334 329818
rect 400714 293818 400746 294374
rect 401302 293818 401334 294374
rect 400714 258374 401334 293818
rect 400714 257818 400746 258374
rect 401302 257818 401334 258374
rect 400714 222374 401334 257818
rect 400714 221818 400746 222374
rect 401302 221818 401334 222374
rect 400714 186374 401334 221818
rect 400714 185818 400746 186374
rect 401302 185818 401334 186374
rect 400714 150374 401334 185818
rect 400714 149818 400746 150374
rect 401302 149818 401334 150374
rect 400714 114374 401334 149818
rect 400714 113818 400746 114374
rect 401302 113818 401334 114374
rect 400714 78374 401334 113818
rect 400714 77818 400746 78374
rect 401302 77818 401334 78374
rect 400714 42374 401334 77818
rect 400714 41818 400746 42374
rect 401302 41818 401334 42374
rect 400714 6374 401334 41818
rect 400714 5818 400746 6374
rect 401302 5818 401334 6374
rect 400714 -3226 401334 5818
rect 400714 -3782 400746 -3226
rect 401302 -3782 401334 -3226
rect 400714 -7654 401334 -3782
rect 401954 708678 402574 711590
rect 401954 708122 401986 708678
rect 402542 708122 402574 708678
rect 401954 691614 402574 708122
rect 401954 691058 401986 691614
rect 402542 691058 402574 691614
rect 401954 655614 402574 691058
rect 401954 655058 401986 655614
rect 402542 655058 402574 655614
rect 401954 619614 402574 655058
rect 401954 619058 401986 619614
rect 402542 619058 402574 619614
rect 401954 583614 402574 619058
rect 401954 583058 401986 583614
rect 402542 583058 402574 583614
rect 401954 547614 402574 583058
rect 401954 547058 401986 547614
rect 402542 547058 402574 547614
rect 401954 511614 402574 547058
rect 401954 511058 401986 511614
rect 402542 511058 402574 511614
rect 401954 475614 402574 511058
rect 401954 475058 401986 475614
rect 402542 475058 402574 475614
rect 401954 439614 402574 475058
rect 401954 439058 401986 439614
rect 402542 439058 402574 439614
rect 401954 403614 402574 439058
rect 401954 403058 401986 403614
rect 402542 403058 402574 403614
rect 401954 367614 402574 403058
rect 401954 367058 401986 367614
rect 402542 367058 402574 367614
rect 401954 331614 402574 367058
rect 401954 331058 401986 331614
rect 402542 331058 402574 331614
rect 401954 295614 402574 331058
rect 401954 295058 401986 295614
rect 402542 295058 402574 295614
rect 401954 259614 402574 295058
rect 401954 259058 401986 259614
rect 402542 259058 402574 259614
rect 401954 223614 402574 259058
rect 401954 223058 401986 223614
rect 402542 223058 402574 223614
rect 401954 187614 402574 223058
rect 401954 187058 401986 187614
rect 402542 187058 402574 187614
rect 401954 151614 402574 187058
rect 401954 151058 401986 151614
rect 402542 151058 402574 151614
rect 401954 115614 402574 151058
rect 401954 115058 401986 115614
rect 402542 115058 402574 115614
rect 401954 79614 402574 115058
rect 401954 79058 401986 79614
rect 402542 79058 402574 79614
rect 401954 43614 402574 79058
rect 401954 43058 401986 43614
rect 402542 43058 402574 43614
rect 401954 7614 402574 43058
rect 401954 7058 401986 7614
rect 402542 7058 402574 7614
rect 401954 -4186 402574 7058
rect 401954 -4742 401986 -4186
rect 402542 -4742 402574 -4186
rect 401954 -7654 402574 -4742
rect 403194 709638 403814 711590
rect 403194 709082 403226 709638
rect 403782 709082 403814 709638
rect 403194 692854 403814 709082
rect 403194 692298 403226 692854
rect 403782 692298 403814 692854
rect 403194 656854 403814 692298
rect 403194 656298 403226 656854
rect 403782 656298 403814 656854
rect 403194 620854 403814 656298
rect 403194 620298 403226 620854
rect 403782 620298 403814 620854
rect 403194 584854 403814 620298
rect 403194 584298 403226 584854
rect 403782 584298 403814 584854
rect 403194 548854 403814 584298
rect 403194 548298 403226 548854
rect 403782 548298 403814 548854
rect 403194 512854 403814 548298
rect 403194 512298 403226 512854
rect 403782 512298 403814 512854
rect 403194 476854 403814 512298
rect 403194 476298 403226 476854
rect 403782 476298 403814 476854
rect 403194 440854 403814 476298
rect 403194 440298 403226 440854
rect 403782 440298 403814 440854
rect 403194 404854 403814 440298
rect 403194 404298 403226 404854
rect 403782 404298 403814 404854
rect 403194 368854 403814 404298
rect 403194 368298 403226 368854
rect 403782 368298 403814 368854
rect 403194 332854 403814 368298
rect 403194 332298 403226 332854
rect 403782 332298 403814 332854
rect 403194 296854 403814 332298
rect 403194 296298 403226 296854
rect 403782 296298 403814 296854
rect 403194 260854 403814 296298
rect 403194 260298 403226 260854
rect 403782 260298 403814 260854
rect 403194 224854 403814 260298
rect 403194 224298 403226 224854
rect 403782 224298 403814 224854
rect 403194 188854 403814 224298
rect 403194 188298 403226 188854
rect 403782 188298 403814 188854
rect 403194 152854 403814 188298
rect 403194 152298 403226 152854
rect 403782 152298 403814 152854
rect 403194 116854 403814 152298
rect 403194 116298 403226 116854
rect 403782 116298 403814 116854
rect 403194 80854 403814 116298
rect 403194 80298 403226 80854
rect 403782 80298 403814 80854
rect 403194 44854 403814 80298
rect 403194 44298 403226 44854
rect 403782 44298 403814 44854
rect 403194 8854 403814 44298
rect 403194 8298 403226 8854
rect 403782 8298 403814 8854
rect 403194 -5146 403814 8298
rect 403194 -5702 403226 -5146
rect 403782 -5702 403814 -5146
rect 403194 -7654 403814 -5702
rect 404434 710598 405054 711590
rect 404434 710042 404466 710598
rect 405022 710042 405054 710598
rect 404434 694094 405054 710042
rect 404434 693538 404466 694094
rect 405022 693538 405054 694094
rect 404434 658094 405054 693538
rect 404434 657538 404466 658094
rect 405022 657538 405054 658094
rect 404434 622094 405054 657538
rect 404434 621538 404466 622094
rect 405022 621538 405054 622094
rect 404434 586094 405054 621538
rect 404434 585538 404466 586094
rect 405022 585538 405054 586094
rect 404434 550094 405054 585538
rect 404434 549538 404466 550094
rect 405022 549538 405054 550094
rect 404434 514094 405054 549538
rect 404434 513538 404466 514094
rect 405022 513538 405054 514094
rect 404434 478094 405054 513538
rect 404434 477538 404466 478094
rect 405022 477538 405054 478094
rect 404434 442094 405054 477538
rect 404434 441538 404466 442094
rect 405022 441538 405054 442094
rect 404434 406094 405054 441538
rect 404434 405538 404466 406094
rect 405022 405538 405054 406094
rect 404434 370094 405054 405538
rect 404434 369538 404466 370094
rect 405022 369538 405054 370094
rect 404434 334094 405054 369538
rect 404434 333538 404466 334094
rect 405022 333538 405054 334094
rect 404434 298094 405054 333538
rect 404434 297538 404466 298094
rect 405022 297538 405054 298094
rect 404434 262094 405054 297538
rect 404434 261538 404466 262094
rect 405022 261538 405054 262094
rect 404434 226094 405054 261538
rect 404434 225538 404466 226094
rect 405022 225538 405054 226094
rect 404434 190094 405054 225538
rect 404434 189538 404466 190094
rect 405022 189538 405054 190094
rect 404434 154094 405054 189538
rect 404434 153538 404466 154094
rect 405022 153538 405054 154094
rect 404434 118094 405054 153538
rect 404434 117538 404466 118094
rect 405022 117538 405054 118094
rect 404434 82094 405054 117538
rect 404434 81538 404466 82094
rect 405022 81538 405054 82094
rect 404434 46094 405054 81538
rect 404434 45538 404466 46094
rect 405022 45538 405054 46094
rect 404434 10094 405054 45538
rect 404434 9538 404466 10094
rect 405022 9538 405054 10094
rect 404434 -6106 405054 9538
rect 404434 -6662 404466 -6106
rect 405022 -6662 405054 -6106
rect 404434 -7654 405054 -6662
rect 405674 711558 406294 711590
rect 405674 711002 405706 711558
rect 406262 711002 406294 711558
rect 405674 695334 406294 711002
rect 405674 694778 405706 695334
rect 406262 694778 406294 695334
rect 405674 659334 406294 694778
rect 405674 658778 405706 659334
rect 406262 658778 406294 659334
rect 405674 623334 406294 658778
rect 405674 622778 405706 623334
rect 406262 622778 406294 623334
rect 405674 587334 406294 622778
rect 405674 586778 405706 587334
rect 406262 586778 406294 587334
rect 405674 551334 406294 586778
rect 405674 550778 405706 551334
rect 406262 550778 406294 551334
rect 405674 515334 406294 550778
rect 405674 514778 405706 515334
rect 406262 514778 406294 515334
rect 405674 479334 406294 514778
rect 405674 478778 405706 479334
rect 406262 478778 406294 479334
rect 405674 443334 406294 478778
rect 405674 442778 405706 443334
rect 406262 442778 406294 443334
rect 405674 407334 406294 442778
rect 405674 406778 405706 407334
rect 406262 406778 406294 407334
rect 405674 371334 406294 406778
rect 405674 370778 405706 371334
rect 406262 370778 406294 371334
rect 405674 335334 406294 370778
rect 405674 334778 405706 335334
rect 406262 334778 406294 335334
rect 405674 299334 406294 334778
rect 405674 298778 405706 299334
rect 406262 298778 406294 299334
rect 405674 263334 406294 298778
rect 405674 262778 405706 263334
rect 406262 262778 406294 263334
rect 405674 227334 406294 262778
rect 405674 226778 405706 227334
rect 406262 226778 406294 227334
rect 405674 191334 406294 226778
rect 405674 190778 405706 191334
rect 406262 190778 406294 191334
rect 405674 155334 406294 190778
rect 405674 154778 405706 155334
rect 406262 154778 406294 155334
rect 405674 119334 406294 154778
rect 405674 118778 405706 119334
rect 406262 118778 406294 119334
rect 405674 83334 406294 118778
rect 405674 82778 405706 83334
rect 406262 82778 406294 83334
rect 405674 47334 406294 82778
rect 405674 46778 405706 47334
rect 406262 46778 406294 47334
rect 405674 11334 406294 46778
rect 405674 10778 405706 11334
rect 406262 10778 406294 11334
rect 405674 -7066 406294 10778
rect 405674 -7622 405706 -7066
rect 406262 -7622 406294 -7066
rect 405674 -7654 406294 -7622
rect 432994 704838 433614 711590
rect 432994 704282 433026 704838
rect 433582 704282 433614 704838
rect 432994 686654 433614 704282
rect 432994 686098 433026 686654
rect 433582 686098 433614 686654
rect 432994 650654 433614 686098
rect 432994 650098 433026 650654
rect 433582 650098 433614 650654
rect 432994 614654 433614 650098
rect 432994 614098 433026 614654
rect 433582 614098 433614 614654
rect 432994 578654 433614 614098
rect 432994 578098 433026 578654
rect 433582 578098 433614 578654
rect 432994 542654 433614 578098
rect 432994 542098 433026 542654
rect 433582 542098 433614 542654
rect 432994 506654 433614 542098
rect 432994 506098 433026 506654
rect 433582 506098 433614 506654
rect 432994 470654 433614 506098
rect 432994 470098 433026 470654
rect 433582 470098 433614 470654
rect 432994 434654 433614 470098
rect 432994 434098 433026 434654
rect 433582 434098 433614 434654
rect 432994 398654 433614 434098
rect 432994 398098 433026 398654
rect 433582 398098 433614 398654
rect 432994 362654 433614 398098
rect 432994 362098 433026 362654
rect 433582 362098 433614 362654
rect 432994 326654 433614 362098
rect 432994 326098 433026 326654
rect 433582 326098 433614 326654
rect 432994 290654 433614 326098
rect 432994 290098 433026 290654
rect 433582 290098 433614 290654
rect 432994 254654 433614 290098
rect 432994 254098 433026 254654
rect 433582 254098 433614 254654
rect 432994 218654 433614 254098
rect 432994 218098 433026 218654
rect 433582 218098 433614 218654
rect 432994 182654 433614 218098
rect 432994 182098 433026 182654
rect 433582 182098 433614 182654
rect 432994 146654 433614 182098
rect 432994 146098 433026 146654
rect 433582 146098 433614 146654
rect 432994 110654 433614 146098
rect 432994 110098 433026 110654
rect 433582 110098 433614 110654
rect 432994 74654 433614 110098
rect 432994 74098 433026 74654
rect 433582 74098 433614 74654
rect 432994 38654 433614 74098
rect 432994 38098 433026 38654
rect 433582 38098 433614 38654
rect 432994 2654 433614 38098
rect 432994 2098 433026 2654
rect 433582 2098 433614 2654
rect 432994 -346 433614 2098
rect 432994 -902 433026 -346
rect 433582 -902 433614 -346
rect 432994 -7654 433614 -902
rect 434234 705798 434854 711590
rect 434234 705242 434266 705798
rect 434822 705242 434854 705798
rect 434234 687894 434854 705242
rect 434234 687338 434266 687894
rect 434822 687338 434854 687894
rect 434234 651894 434854 687338
rect 434234 651338 434266 651894
rect 434822 651338 434854 651894
rect 434234 615894 434854 651338
rect 434234 615338 434266 615894
rect 434822 615338 434854 615894
rect 434234 579894 434854 615338
rect 434234 579338 434266 579894
rect 434822 579338 434854 579894
rect 434234 543894 434854 579338
rect 434234 543338 434266 543894
rect 434822 543338 434854 543894
rect 434234 507894 434854 543338
rect 434234 507338 434266 507894
rect 434822 507338 434854 507894
rect 434234 471894 434854 507338
rect 434234 471338 434266 471894
rect 434822 471338 434854 471894
rect 434234 435894 434854 471338
rect 434234 435338 434266 435894
rect 434822 435338 434854 435894
rect 434234 399894 434854 435338
rect 434234 399338 434266 399894
rect 434822 399338 434854 399894
rect 434234 363894 434854 399338
rect 434234 363338 434266 363894
rect 434822 363338 434854 363894
rect 434234 327894 434854 363338
rect 434234 327338 434266 327894
rect 434822 327338 434854 327894
rect 434234 291894 434854 327338
rect 434234 291338 434266 291894
rect 434822 291338 434854 291894
rect 434234 255894 434854 291338
rect 434234 255338 434266 255894
rect 434822 255338 434854 255894
rect 434234 219894 434854 255338
rect 434234 219338 434266 219894
rect 434822 219338 434854 219894
rect 434234 183894 434854 219338
rect 434234 183338 434266 183894
rect 434822 183338 434854 183894
rect 434234 147894 434854 183338
rect 434234 147338 434266 147894
rect 434822 147338 434854 147894
rect 434234 111894 434854 147338
rect 434234 111338 434266 111894
rect 434822 111338 434854 111894
rect 434234 75894 434854 111338
rect 434234 75338 434266 75894
rect 434822 75338 434854 75894
rect 434234 39894 434854 75338
rect 434234 39338 434266 39894
rect 434822 39338 434854 39894
rect 434234 3894 434854 39338
rect 434234 3338 434266 3894
rect 434822 3338 434854 3894
rect 434234 -1306 434854 3338
rect 434234 -1862 434266 -1306
rect 434822 -1862 434854 -1306
rect 434234 -7654 434854 -1862
rect 435474 706758 436094 711590
rect 435474 706202 435506 706758
rect 436062 706202 436094 706758
rect 435474 689134 436094 706202
rect 435474 688578 435506 689134
rect 436062 688578 436094 689134
rect 435474 653134 436094 688578
rect 435474 652578 435506 653134
rect 436062 652578 436094 653134
rect 435474 617134 436094 652578
rect 435474 616578 435506 617134
rect 436062 616578 436094 617134
rect 435474 581134 436094 616578
rect 435474 580578 435506 581134
rect 436062 580578 436094 581134
rect 435474 545134 436094 580578
rect 435474 544578 435506 545134
rect 436062 544578 436094 545134
rect 435474 509134 436094 544578
rect 435474 508578 435506 509134
rect 436062 508578 436094 509134
rect 435474 473134 436094 508578
rect 435474 472578 435506 473134
rect 436062 472578 436094 473134
rect 435474 437134 436094 472578
rect 435474 436578 435506 437134
rect 436062 436578 436094 437134
rect 435474 401134 436094 436578
rect 435474 400578 435506 401134
rect 436062 400578 436094 401134
rect 435474 365134 436094 400578
rect 435474 364578 435506 365134
rect 436062 364578 436094 365134
rect 435474 329134 436094 364578
rect 435474 328578 435506 329134
rect 436062 328578 436094 329134
rect 435474 293134 436094 328578
rect 435474 292578 435506 293134
rect 436062 292578 436094 293134
rect 435474 257134 436094 292578
rect 435474 256578 435506 257134
rect 436062 256578 436094 257134
rect 435474 221134 436094 256578
rect 435474 220578 435506 221134
rect 436062 220578 436094 221134
rect 435474 185134 436094 220578
rect 435474 184578 435506 185134
rect 436062 184578 436094 185134
rect 435474 149134 436094 184578
rect 435474 148578 435506 149134
rect 436062 148578 436094 149134
rect 435474 113134 436094 148578
rect 435474 112578 435506 113134
rect 436062 112578 436094 113134
rect 435474 77134 436094 112578
rect 435474 76578 435506 77134
rect 436062 76578 436094 77134
rect 435474 41134 436094 76578
rect 435474 40578 435506 41134
rect 436062 40578 436094 41134
rect 435474 5134 436094 40578
rect 435474 4578 435506 5134
rect 436062 4578 436094 5134
rect 435474 -2266 436094 4578
rect 435474 -2822 435506 -2266
rect 436062 -2822 436094 -2266
rect 435474 -7654 436094 -2822
rect 436714 707718 437334 711590
rect 436714 707162 436746 707718
rect 437302 707162 437334 707718
rect 436714 690374 437334 707162
rect 436714 689818 436746 690374
rect 437302 689818 437334 690374
rect 436714 654374 437334 689818
rect 436714 653818 436746 654374
rect 437302 653818 437334 654374
rect 436714 618374 437334 653818
rect 436714 617818 436746 618374
rect 437302 617818 437334 618374
rect 436714 582374 437334 617818
rect 436714 581818 436746 582374
rect 437302 581818 437334 582374
rect 436714 546374 437334 581818
rect 436714 545818 436746 546374
rect 437302 545818 437334 546374
rect 436714 510374 437334 545818
rect 436714 509818 436746 510374
rect 437302 509818 437334 510374
rect 436714 474374 437334 509818
rect 436714 473818 436746 474374
rect 437302 473818 437334 474374
rect 436714 438374 437334 473818
rect 436714 437818 436746 438374
rect 437302 437818 437334 438374
rect 436714 402374 437334 437818
rect 436714 401818 436746 402374
rect 437302 401818 437334 402374
rect 436714 366374 437334 401818
rect 436714 365818 436746 366374
rect 437302 365818 437334 366374
rect 436714 330374 437334 365818
rect 436714 329818 436746 330374
rect 437302 329818 437334 330374
rect 436714 294374 437334 329818
rect 436714 293818 436746 294374
rect 437302 293818 437334 294374
rect 436714 258374 437334 293818
rect 436714 257818 436746 258374
rect 437302 257818 437334 258374
rect 436714 222374 437334 257818
rect 436714 221818 436746 222374
rect 437302 221818 437334 222374
rect 436714 186374 437334 221818
rect 436714 185818 436746 186374
rect 437302 185818 437334 186374
rect 436714 150374 437334 185818
rect 436714 149818 436746 150374
rect 437302 149818 437334 150374
rect 436714 114374 437334 149818
rect 436714 113818 436746 114374
rect 437302 113818 437334 114374
rect 436714 78374 437334 113818
rect 436714 77818 436746 78374
rect 437302 77818 437334 78374
rect 436714 42374 437334 77818
rect 436714 41818 436746 42374
rect 437302 41818 437334 42374
rect 436714 6374 437334 41818
rect 436714 5818 436746 6374
rect 437302 5818 437334 6374
rect 436714 -3226 437334 5818
rect 436714 -3782 436746 -3226
rect 437302 -3782 437334 -3226
rect 436714 -7654 437334 -3782
rect 437954 708678 438574 711590
rect 437954 708122 437986 708678
rect 438542 708122 438574 708678
rect 437954 691614 438574 708122
rect 437954 691058 437986 691614
rect 438542 691058 438574 691614
rect 437954 655614 438574 691058
rect 437954 655058 437986 655614
rect 438542 655058 438574 655614
rect 437954 619614 438574 655058
rect 437954 619058 437986 619614
rect 438542 619058 438574 619614
rect 437954 583614 438574 619058
rect 437954 583058 437986 583614
rect 438542 583058 438574 583614
rect 437954 547614 438574 583058
rect 437954 547058 437986 547614
rect 438542 547058 438574 547614
rect 437954 511614 438574 547058
rect 437954 511058 437986 511614
rect 438542 511058 438574 511614
rect 437954 475614 438574 511058
rect 437954 475058 437986 475614
rect 438542 475058 438574 475614
rect 437954 439614 438574 475058
rect 437954 439058 437986 439614
rect 438542 439058 438574 439614
rect 437954 403614 438574 439058
rect 437954 403058 437986 403614
rect 438542 403058 438574 403614
rect 437954 367614 438574 403058
rect 437954 367058 437986 367614
rect 438542 367058 438574 367614
rect 437954 331614 438574 367058
rect 437954 331058 437986 331614
rect 438542 331058 438574 331614
rect 437954 295614 438574 331058
rect 437954 295058 437986 295614
rect 438542 295058 438574 295614
rect 437954 259614 438574 295058
rect 437954 259058 437986 259614
rect 438542 259058 438574 259614
rect 437954 223614 438574 259058
rect 437954 223058 437986 223614
rect 438542 223058 438574 223614
rect 437954 187614 438574 223058
rect 437954 187058 437986 187614
rect 438542 187058 438574 187614
rect 437954 151614 438574 187058
rect 437954 151058 437986 151614
rect 438542 151058 438574 151614
rect 437954 115614 438574 151058
rect 437954 115058 437986 115614
rect 438542 115058 438574 115614
rect 437954 79614 438574 115058
rect 437954 79058 437986 79614
rect 438542 79058 438574 79614
rect 437954 43614 438574 79058
rect 437954 43058 437986 43614
rect 438542 43058 438574 43614
rect 437954 7614 438574 43058
rect 437954 7058 437986 7614
rect 438542 7058 438574 7614
rect 437954 -4186 438574 7058
rect 437954 -4742 437986 -4186
rect 438542 -4742 438574 -4186
rect 437954 -7654 438574 -4742
rect 439194 709638 439814 711590
rect 439194 709082 439226 709638
rect 439782 709082 439814 709638
rect 439194 692854 439814 709082
rect 439194 692298 439226 692854
rect 439782 692298 439814 692854
rect 439194 656854 439814 692298
rect 439194 656298 439226 656854
rect 439782 656298 439814 656854
rect 439194 620854 439814 656298
rect 439194 620298 439226 620854
rect 439782 620298 439814 620854
rect 439194 584854 439814 620298
rect 439194 584298 439226 584854
rect 439782 584298 439814 584854
rect 439194 548854 439814 584298
rect 439194 548298 439226 548854
rect 439782 548298 439814 548854
rect 439194 512854 439814 548298
rect 439194 512298 439226 512854
rect 439782 512298 439814 512854
rect 439194 476854 439814 512298
rect 439194 476298 439226 476854
rect 439782 476298 439814 476854
rect 439194 440854 439814 476298
rect 439194 440298 439226 440854
rect 439782 440298 439814 440854
rect 439194 404854 439814 440298
rect 439194 404298 439226 404854
rect 439782 404298 439814 404854
rect 439194 368854 439814 404298
rect 439194 368298 439226 368854
rect 439782 368298 439814 368854
rect 439194 332854 439814 368298
rect 439194 332298 439226 332854
rect 439782 332298 439814 332854
rect 439194 296854 439814 332298
rect 439194 296298 439226 296854
rect 439782 296298 439814 296854
rect 439194 260854 439814 296298
rect 439194 260298 439226 260854
rect 439782 260298 439814 260854
rect 439194 224854 439814 260298
rect 439194 224298 439226 224854
rect 439782 224298 439814 224854
rect 439194 188854 439814 224298
rect 439194 188298 439226 188854
rect 439782 188298 439814 188854
rect 439194 152854 439814 188298
rect 439194 152298 439226 152854
rect 439782 152298 439814 152854
rect 439194 116854 439814 152298
rect 439194 116298 439226 116854
rect 439782 116298 439814 116854
rect 439194 80854 439814 116298
rect 439194 80298 439226 80854
rect 439782 80298 439814 80854
rect 439194 44854 439814 80298
rect 439194 44298 439226 44854
rect 439782 44298 439814 44854
rect 439194 8854 439814 44298
rect 439194 8298 439226 8854
rect 439782 8298 439814 8854
rect 439194 -5146 439814 8298
rect 439194 -5702 439226 -5146
rect 439782 -5702 439814 -5146
rect 439194 -7654 439814 -5702
rect 440434 710598 441054 711590
rect 440434 710042 440466 710598
rect 441022 710042 441054 710598
rect 440434 694094 441054 710042
rect 440434 693538 440466 694094
rect 441022 693538 441054 694094
rect 440434 658094 441054 693538
rect 440434 657538 440466 658094
rect 441022 657538 441054 658094
rect 440434 622094 441054 657538
rect 440434 621538 440466 622094
rect 441022 621538 441054 622094
rect 440434 586094 441054 621538
rect 440434 585538 440466 586094
rect 441022 585538 441054 586094
rect 440434 550094 441054 585538
rect 440434 549538 440466 550094
rect 441022 549538 441054 550094
rect 440434 514094 441054 549538
rect 440434 513538 440466 514094
rect 441022 513538 441054 514094
rect 440434 478094 441054 513538
rect 440434 477538 440466 478094
rect 441022 477538 441054 478094
rect 440434 442094 441054 477538
rect 440434 441538 440466 442094
rect 441022 441538 441054 442094
rect 440434 406094 441054 441538
rect 440434 405538 440466 406094
rect 441022 405538 441054 406094
rect 440434 370094 441054 405538
rect 440434 369538 440466 370094
rect 441022 369538 441054 370094
rect 440434 334094 441054 369538
rect 440434 333538 440466 334094
rect 441022 333538 441054 334094
rect 440434 298094 441054 333538
rect 440434 297538 440466 298094
rect 441022 297538 441054 298094
rect 440434 262094 441054 297538
rect 440434 261538 440466 262094
rect 441022 261538 441054 262094
rect 440434 226094 441054 261538
rect 440434 225538 440466 226094
rect 441022 225538 441054 226094
rect 440434 190094 441054 225538
rect 440434 189538 440466 190094
rect 441022 189538 441054 190094
rect 440434 154094 441054 189538
rect 440434 153538 440466 154094
rect 441022 153538 441054 154094
rect 440434 118094 441054 153538
rect 440434 117538 440466 118094
rect 441022 117538 441054 118094
rect 440434 82094 441054 117538
rect 440434 81538 440466 82094
rect 441022 81538 441054 82094
rect 440434 46094 441054 81538
rect 440434 45538 440466 46094
rect 441022 45538 441054 46094
rect 440434 10094 441054 45538
rect 440434 9538 440466 10094
rect 441022 9538 441054 10094
rect 440434 -6106 441054 9538
rect 440434 -6662 440466 -6106
rect 441022 -6662 441054 -6106
rect 440434 -7654 441054 -6662
rect 441674 711558 442294 711590
rect 441674 711002 441706 711558
rect 442262 711002 442294 711558
rect 441674 695334 442294 711002
rect 441674 694778 441706 695334
rect 442262 694778 442294 695334
rect 441674 659334 442294 694778
rect 441674 658778 441706 659334
rect 442262 658778 442294 659334
rect 441674 623334 442294 658778
rect 441674 622778 441706 623334
rect 442262 622778 442294 623334
rect 441674 587334 442294 622778
rect 441674 586778 441706 587334
rect 442262 586778 442294 587334
rect 441674 551334 442294 586778
rect 441674 550778 441706 551334
rect 442262 550778 442294 551334
rect 441674 515334 442294 550778
rect 441674 514778 441706 515334
rect 442262 514778 442294 515334
rect 441674 479334 442294 514778
rect 441674 478778 441706 479334
rect 442262 478778 442294 479334
rect 441674 443334 442294 478778
rect 441674 442778 441706 443334
rect 442262 442778 442294 443334
rect 441674 407334 442294 442778
rect 441674 406778 441706 407334
rect 442262 406778 442294 407334
rect 441674 371334 442294 406778
rect 441674 370778 441706 371334
rect 442262 370778 442294 371334
rect 441674 335334 442294 370778
rect 441674 334778 441706 335334
rect 442262 334778 442294 335334
rect 441674 299334 442294 334778
rect 441674 298778 441706 299334
rect 442262 298778 442294 299334
rect 441674 263334 442294 298778
rect 441674 262778 441706 263334
rect 442262 262778 442294 263334
rect 441674 227334 442294 262778
rect 441674 226778 441706 227334
rect 442262 226778 442294 227334
rect 441674 191334 442294 226778
rect 441674 190778 441706 191334
rect 442262 190778 442294 191334
rect 441674 155334 442294 190778
rect 441674 154778 441706 155334
rect 442262 154778 442294 155334
rect 441674 119334 442294 154778
rect 441674 118778 441706 119334
rect 442262 118778 442294 119334
rect 441674 83334 442294 118778
rect 441674 82778 441706 83334
rect 442262 82778 442294 83334
rect 441674 47334 442294 82778
rect 441674 46778 441706 47334
rect 442262 46778 442294 47334
rect 441674 11334 442294 46778
rect 441674 10778 441706 11334
rect 442262 10778 442294 11334
rect 441674 -7066 442294 10778
rect 441674 -7622 441706 -7066
rect 442262 -7622 442294 -7066
rect 441674 -7654 442294 -7622
rect 468994 704838 469614 711590
rect 468994 704282 469026 704838
rect 469582 704282 469614 704838
rect 468994 686654 469614 704282
rect 468994 686098 469026 686654
rect 469582 686098 469614 686654
rect 468994 650654 469614 686098
rect 468994 650098 469026 650654
rect 469582 650098 469614 650654
rect 468994 614654 469614 650098
rect 468994 614098 469026 614654
rect 469582 614098 469614 614654
rect 468994 578654 469614 614098
rect 468994 578098 469026 578654
rect 469582 578098 469614 578654
rect 468994 542654 469614 578098
rect 468994 542098 469026 542654
rect 469582 542098 469614 542654
rect 468994 506654 469614 542098
rect 468994 506098 469026 506654
rect 469582 506098 469614 506654
rect 468994 470654 469614 506098
rect 468994 470098 469026 470654
rect 469582 470098 469614 470654
rect 468994 450397 469614 470098
rect 468994 450093 469032 450397
rect 469576 450093 469614 450397
rect 468994 434654 469614 450093
rect 468994 434098 469026 434654
rect 469582 434098 469614 434654
rect 468994 431997 469614 434098
rect 468994 431693 469032 431997
rect 469576 431693 469614 431997
rect 468994 410998 469614 431693
rect 468994 410694 469032 410998
rect 469576 410694 469614 410998
rect 468994 398654 469614 410694
rect 468994 398098 469026 398654
rect 469582 398098 469614 398654
rect 468994 390002 469614 398098
rect 468994 389698 469032 390002
rect 469576 389698 469614 390002
rect 468994 368999 469614 389698
rect 468994 368695 469032 368999
rect 469576 368695 469614 368999
rect 468994 362654 469614 368695
rect 468994 362098 469026 362654
rect 469582 362098 469614 362654
rect 468994 347997 469614 362098
rect 468994 347693 469032 347997
rect 469576 347693 469614 347997
rect 468994 326997 469614 347693
rect 468994 326693 469032 326997
rect 469576 326693 469614 326997
rect 468994 326654 469614 326693
rect 468994 326098 469026 326654
rect 469582 326098 469614 326654
rect 468994 305999 469614 326098
rect 468994 305695 469032 305999
rect 469576 305695 469614 305999
rect 468994 290654 469614 305695
rect 468994 290098 469026 290654
rect 469582 290098 469614 290654
rect 468994 285000 469614 290098
rect 468994 284696 469032 285000
rect 469576 284696 469614 285000
rect 468994 263999 469614 284696
rect 468994 263695 469032 263999
rect 469576 263695 469614 263999
rect 468994 254654 469614 263695
rect 468994 254098 469026 254654
rect 469582 254098 469614 254654
rect 468994 218654 469614 254098
rect 468994 218098 469026 218654
rect 469582 218098 469614 218654
rect 468994 182654 469614 218098
rect 468994 182098 469026 182654
rect 469582 182098 469614 182654
rect 468994 146654 469614 182098
rect 468994 146098 469026 146654
rect 469582 146098 469614 146654
rect 468994 110654 469614 146098
rect 468994 110098 469026 110654
rect 469582 110098 469614 110654
rect 468994 74654 469614 110098
rect 468994 74098 469026 74654
rect 469582 74098 469614 74654
rect 468994 38654 469614 74098
rect 468994 38098 469026 38654
rect 469582 38098 469614 38654
rect 468994 2654 469614 38098
rect 468994 2098 469026 2654
rect 469582 2098 469614 2654
rect 468994 -346 469614 2098
rect 468994 -902 469026 -346
rect 469582 -902 469614 -346
rect 468994 -7654 469614 -902
rect 470234 705798 470854 711590
rect 470234 705242 470266 705798
rect 470822 705242 470854 705798
rect 470234 687894 470854 705242
rect 470234 687338 470266 687894
rect 470822 687338 470854 687894
rect 470234 651894 470854 687338
rect 470234 651338 470266 651894
rect 470822 651338 470854 651894
rect 470234 615894 470854 651338
rect 470234 615338 470266 615894
rect 470822 615338 470854 615894
rect 470234 579894 470854 615338
rect 470234 579338 470266 579894
rect 470822 579338 470854 579894
rect 470234 543894 470854 579338
rect 470234 543338 470266 543894
rect 470822 543338 470854 543894
rect 470234 507894 470854 543338
rect 470234 507338 470266 507894
rect 470822 507338 470854 507894
rect 470234 471894 470854 507338
rect 470234 471338 470266 471894
rect 470822 471338 470854 471894
rect 470234 451483 470854 471338
rect 470234 451179 470272 451483
rect 470816 451179 470854 451483
rect 470234 449312 470854 451179
rect 470234 449008 470272 449312
rect 470816 449008 470854 449312
rect 470234 435894 470854 449008
rect 470234 435338 470266 435894
rect 470822 435338 470854 435894
rect 470234 433084 470854 435338
rect 470234 432780 470272 433084
rect 470816 432780 470854 433084
rect 470234 430912 470854 432780
rect 470234 430608 470272 430912
rect 470816 430608 470854 430912
rect 470234 412084 470854 430608
rect 470234 411780 470272 412084
rect 470816 411780 470854 412084
rect 470234 409912 470854 411780
rect 470234 409608 470272 409912
rect 470816 409608 470854 409912
rect 470234 399894 470854 409608
rect 470234 399338 470266 399894
rect 470822 399338 470854 399894
rect 470234 391085 470854 399338
rect 470234 390781 470272 391085
rect 470816 390781 470854 391085
rect 470234 388912 470854 390781
rect 470234 388608 470272 388912
rect 470816 388608 470854 388912
rect 470234 370085 470854 388608
rect 470234 369781 470272 370085
rect 470816 369781 470854 370085
rect 470234 367912 470854 369781
rect 470234 367608 470272 367912
rect 470816 367608 470854 367912
rect 470234 363894 470854 367608
rect 470234 363338 470266 363894
rect 470822 363338 470854 363894
rect 470234 349084 470854 363338
rect 470234 348780 470272 349084
rect 470816 348780 470854 349084
rect 470234 346912 470854 348780
rect 470234 346608 470272 346912
rect 470816 346608 470854 346912
rect 470234 328084 470854 346608
rect 470234 327894 470272 328084
rect 470816 327894 470854 328084
rect 470234 327338 470266 327894
rect 470822 327338 470854 327894
rect 470234 325912 470854 327338
rect 470234 325608 470272 325912
rect 470816 325608 470854 325912
rect 470234 307084 470854 325608
rect 470234 306780 470272 307084
rect 470816 306780 470854 307084
rect 470234 304912 470854 306780
rect 470234 304608 470272 304912
rect 470816 304608 470854 304912
rect 470234 291894 470854 304608
rect 470234 291338 470266 291894
rect 470822 291338 470854 291894
rect 470234 286085 470854 291338
rect 470234 285781 470272 286085
rect 470816 285781 470854 286085
rect 470234 283912 470854 285781
rect 470234 283608 470272 283912
rect 470816 283608 470854 283912
rect 470234 265085 470854 283608
rect 470234 264781 470272 265085
rect 470816 264781 470854 265085
rect 470234 262912 470854 264781
rect 470234 262608 470272 262912
rect 470816 262608 470854 262912
rect 470234 255894 470854 262608
rect 470234 255338 470266 255894
rect 470822 255338 470854 255894
rect 470234 219894 470854 255338
rect 470234 219338 470266 219894
rect 470822 219338 470854 219894
rect 470234 183894 470854 219338
rect 470234 183338 470266 183894
rect 470822 183338 470854 183894
rect 470234 147894 470854 183338
rect 470234 147338 470266 147894
rect 470822 147338 470854 147894
rect 470234 111894 470854 147338
rect 470234 111338 470266 111894
rect 470822 111338 470854 111894
rect 470234 75894 470854 111338
rect 470234 75338 470266 75894
rect 470822 75338 470854 75894
rect 470234 39894 470854 75338
rect 470234 39338 470266 39894
rect 470822 39338 470854 39894
rect 470234 3894 470854 39338
rect 470234 3338 470266 3894
rect 470822 3338 470854 3894
rect 470234 -1306 470854 3338
rect 470234 -1862 470266 -1306
rect 470822 -1862 470854 -1306
rect 470234 -7654 470854 -1862
rect 471474 706758 472094 711590
rect 471474 706202 471506 706758
rect 472062 706202 472094 706758
rect 471474 689134 472094 706202
rect 471474 688578 471506 689134
rect 472062 688578 472094 689134
rect 471474 653134 472094 688578
rect 471474 652578 471506 653134
rect 472062 652578 472094 653134
rect 471474 617134 472094 652578
rect 471474 616578 471506 617134
rect 472062 616578 472094 617134
rect 471474 581134 472094 616578
rect 471474 580578 471506 581134
rect 472062 580578 472094 581134
rect 471474 545134 472094 580578
rect 471474 544578 471506 545134
rect 472062 544578 472094 545134
rect 471474 509134 472094 544578
rect 471474 508578 471506 509134
rect 472062 508578 472094 509134
rect 471474 473134 472094 508578
rect 471474 472578 471506 473134
rect 472062 472578 472094 473134
rect 471474 437134 472094 472578
rect 471474 436578 471506 437134
rect 472062 436578 472094 437134
rect 471474 401134 472094 436578
rect 471474 400578 471506 401134
rect 472062 400578 472094 401134
rect 471474 365134 472094 400578
rect 472714 707718 473334 711590
rect 472714 707162 472746 707718
rect 473302 707162 473334 707718
rect 472714 690374 473334 707162
rect 472714 689818 472746 690374
rect 473302 689818 473334 690374
rect 472714 654374 473334 689818
rect 472714 653818 472746 654374
rect 473302 653818 473334 654374
rect 472714 618374 473334 653818
rect 472714 617818 472746 618374
rect 473302 617818 473334 618374
rect 472714 582374 473334 617818
rect 472714 581818 472746 582374
rect 473302 581818 473334 582374
rect 472714 546374 473334 581818
rect 472714 545818 472746 546374
rect 473302 545818 473334 546374
rect 472714 510374 473334 545818
rect 472714 509818 472746 510374
rect 473302 509818 473334 510374
rect 472714 474374 473334 509818
rect 472714 473818 472746 474374
rect 473302 473818 473334 474374
rect 472714 438374 473334 473818
rect 472714 437818 472746 438374
rect 473302 437818 473334 438374
rect 472714 402374 473334 437818
rect 472714 401818 472746 402374
rect 473302 401818 473334 402374
rect 472714 370660 473334 401818
rect 473954 708678 474574 711590
rect 473954 708122 473986 708678
rect 474542 708122 474574 708678
rect 473954 691614 474574 708122
rect 473954 691058 473986 691614
rect 474542 691058 474574 691614
rect 473954 655614 474574 691058
rect 473954 655058 473986 655614
rect 474542 655058 474574 655614
rect 473954 619614 474574 655058
rect 473954 619058 473986 619614
rect 474542 619058 474574 619614
rect 473954 583614 474574 619058
rect 473954 583058 473986 583614
rect 474542 583058 474574 583614
rect 473954 547614 474574 583058
rect 473954 547058 473986 547614
rect 474542 547058 474574 547614
rect 473954 511614 474574 547058
rect 473954 511058 473986 511614
rect 474542 511058 474574 511614
rect 473954 475614 474574 511058
rect 473954 475058 473986 475614
rect 474542 475058 474574 475614
rect 473954 439614 474574 475058
rect 473954 439058 473986 439614
rect 474542 439058 474574 439614
rect 473954 403614 474574 439058
rect 473954 403058 473986 403614
rect 474542 403058 474574 403614
rect 473954 370660 474574 403058
rect 475194 709638 475814 711590
rect 475194 709082 475226 709638
rect 475782 709082 475814 709638
rect 475194 692854 475814 709082
rect 475194 692298 475226 692854
rect 475782 692298 475814 692854
rect 475194 656854 475814 692298
rect 475194 656298 475226 656854
rect 475782 656298 475814 656854
rect 475194 620854 475814 656298
rect 475194 620298 475226 620854
rect 475782 620298 475814 620854
rect 475194 584854 475814 620298
rect 475194 584298 475226 584854
rect 475782 584298 475814 584854
rect 475194 548854 475814 584298
rect 475194 548298 475226 548854
rect 475782 548298 475814 548854
rect 475194 512854 475814 548298
rect 475194 512298 475226 512854
rect 475782 512298 475814 512854
rect 475194 476854 475814 512298
rect 475194 476298 475226 476854
rect 475782 476298 475814 476854
rect 475194 440854 475814 476298
rect 475194 440298 475226 440854
rect 475782 440298 475814 440854
rect 475194 404854 475814 440298
rect 475194 404298 475226 404854
rect 475782 404298 475814 404854
rect 475194 370660 475814 404298
rect 476434 710598 477054 711590
rect 476434 710042 476466 710598
rect 477022 710042 477054 710598
rect 476434 694094 477054 710042
rect 476434 693538 476466 694094
rect 477022 693538 477054 694094
rect 476434 658094 477054 693538
rect 476434 657538 476466 658094
rect 477022 657538 477054 658094
rect 476434 622094 477054 657538
rect 476434 621538 476466 622094
rect 477022 621538 477054 622094
rect 476434 586094 477054 621538
rect 476434 585538 476466 586094
rect 477022 585538 477054 586094
rect 476434 550094 477054 585538
rect 476434 549538 476466 550094
rect 477022 549538 477054 550094
rect 476434 514094 477054 549538
rect 476434 513538 476466 514094
rect 477022 513538 477054 514094
rect 476434 478094 477054 513538
rect 476434 477538 476466 478094
rect 477022 477538 477054 478094
rect 476434 442094 477054 477538
rect 476434 441538 476466 442094
rect 477022 441538 477054 442094
rect 476434 406094 477054 441538
rect 476434 405538 476466 406094
rect 477022 405538 477054 406094
rect 476434 370660 477054 405538
rect 477674 711558 478294 711590
rect 477674 711002 477706 711558
rect 478262 711002 478294 711558
rect 477674 695334 478294 711002
rect 477674 694778 477706 695334
rect 478262 694778 478294 695334
rect 477674 659334 478294 694778
rect 477674 658778 477706 659334
rect 478262 658778 478294 659334
rect 477674 623334 478294 658778
rect 477674 622778 477706 623334
rect 478262 622778 478294 623334
rect 477674 587334 478294 622778
rect 477674 586778 477706 587334
rect 478262 586778 478294 587334
rect 477674 551334 478294 586778
rect 477674 550778 477706 551334
rect 478262 550778 478294 551334
rect 477674 515334 478294 550778
rect 477674 514778 477706 515334
rect 478262 514778 478294 515334
rect 477674 479334 478294 514778
rect 477674 478778 477706 479334
rect 478262 478778 478294 479334
rect 477674 443334 478294 478778
rect 477674 442778 477706 443334
rect 478262 442778 478294 443334
rect 477674 407334 478294 442778
rect 477674 406778 477706 407334
rect 478262 406778 478294 407334
rect 477674 371334 478294 406778
rect 477674 370778 477706 371334
rect 478262 370778 478294 371334
rect 477674 370660 478294 370778
rect 504994 704838 505614 711590
rect 504994 704282 505026 704838
rect 505582 704282 505614 704838
rect 504994 686654 505614 704282
rect 504994 686098 505026 686654
rect 505582 686098 505614 686654
rect 504994 650654 505614 686098
rect 504994 650098 505026 650654
rect 505582 650098 505614 650654
rect 504994 614654 505614 650098
rect 504994 614098 505026 614654
rect 505582 614098 505614 614654
rect 504994 578654 505614 614098
rect 504994 578098 505026 578654
rect 505582 578098 505614 578654
rect 504994 542654 505614 578098
rect 504994 542098 505026 542654
rect 505582 542098 505614 542654
rect 504994 506654 505614 542098
rect 504994 506098 505026 506654
rect 505582 506098 505614 506654
rect 504994 470654 505614 506098
rect 504994 470098 505026 470654
rect 505582 470098 505614 470654
rect 504994 434654 505614 470098
rect 504994 434098 505026 434654
rect 505582 434098 505614 434654
rect 504994 398654 505614 434098
rect 504994 398098 505026 398654
rect 505582 398098 505614 398654
rect 471474 364578 471506 365134
rect 472062 364578 472094 365134
rect 471474 329134 472094 364578
rect 471474 328578 471506 329134
rect 472062 328578 472094 329134
rect 471474 293134 472094 328578
rect 471474 292578 471506 293134
rect 472062 292578 472094 293134
rect 471474 257134 472094 292578
rect 472714 366119 473334 366216
rect 472714 365883 472746 366119
rect 472982 365883 473066 366119
rect 473302 365883 473334 366119
rect 472714 330374 473334 365883
rect 472714 329818 472746 330374
rect 473302 329818 473334 330374
rect 472714 294374 473334 329818
rect 472714 293818 472746 294374
rect 473302 293818 473334 294374
rect 472714 265660 473334 293818
rect 473954 331614 474574 366216
rect 473954 331058 473986 331614
rect 474542 331058 474574 331614
rect 473954 295614 474574 331058
rect 473954 295058 473986 295614
rect 474542 295058 474574 295614
rect 473954 265660 474574 295058
rect 475194 332854 475814 366216
rect 475194 332298 475226 332854
rect 475782 332298 475814 332854
rect 475194 296854 475814 332298
rect 475194 296298 475226 296854
rect 475782 296298 475814 296854
rect 475194 265660 475814 296298
rect 476434 334094 477054 366216
rect 476434 333538 476466 334094
rect 477022 333538 477054 334094
rect 476434 298094 477054 333538
rect 476434 297538 476466 298094
rect 477022 297538 477054 298094
rect 476434 265660 477054 297538
rect 477674 335334 478294 366216
rect 477674 334778 477706 335334
rect 478262 334778 478294 335334
rect 477674 299334 478294 334778
rect 477674 298778 477706 299334
rect 478262 298778 478294 299334
rect 477674 265660 478294 298778
rect 504994 362654 505614 398098
rect 504994 362098 505026 362654
rect 505582 362098 505614 362654
rect 504994 326654 505614 362098
rect 504994 326098 505026 326654
rect 505582 326098 505614 326654
rect 504994 290654 505614 326098
rect 504994 290098 505026 290654
rect 505582 290098 505614 290654
rect 471474 256578 471506 257134
rect 472062 256578 472094 257134
rect 471474 221134 472094 256578
rect 471474 220578 471506 221134
rect 472062 220578 472094 221134
rect 471474 185134 472094 220578
rect 471474 184578 471506 185134
rect 472062 184578 472094 185134
rect 471474 149134 472094 184578
rect 471474 148578 471506 149134
rect 472062 148578 472094 149134
rect 471474 113134 472094 148578
rect 471474 112578 471506 113134
rect 472062 112578 472094 113134
rect 471474 77134 472094 112578
rect 471474 76578 471506 77134
rect 472062 76578 472094 77134
rect 471474 41134 472094 76578
rect 471474 40578 471506 41134
rect 472062 40578 472094 41134
rect 471474 5134 472094 40578
rect 471474 4578 471506 5134
rect 472062 4578 472094 5134
rect 471474 -2266 472094 4578
rect 471474 -2822 471506 -2266
rect 472062 -2822 472094 -2266
rect 471474 -7654 472094 -2822
rect 472714 258374 473334 261216
rect 472714 257818 472746 258374
rect 473302 257818 473334 258374
rect 472714 222374 473334 257818
rect 472714 221818 472746 222374
rect 473302 221818 473334 222374
rect 472714 186374 473334 221818
rect 472714 185818 472746 186374
rect 473302 185818 473334 186374
rect 472714 150374 473334 185818
rect 472714 149818 472746 150374
rect 473302 149818 473334 150374
rect 472714 114374 473334 149818
rect 472714 113818 472746 114374
rect 473302 113818 473334 114374
rect 472714 78374 473334 113818
rect 472714 77818 472746 78374
rect 473302 77818 473334 78374
rect 472714 42374 473334 77818
rect 472714 41818 472746 42374
rect 473302 41818 473334 42374
rect 472714 6374 473334 41818
rect 472714 5818 472746 6374
rect 473302 5818 473334 6374
rect 472714 -3226 473334 5818
rect 472714 -3782 472746 -3226
rect 473302 -3782 473334 -3226
rect 472714 -7654 473334 -3782
rect 473954 259614 474574 261216
rect 473954 259058 473986 259614
rect 474542 259058 474574 259614
rect 473954 223614 474574 259058
rect 473954 223058 473986 223614
rect 474542 223058 474574 223614
rect 473954 187614 474574 223058
rect 473954 187058 473986 187614
rect 474542 187058 474574 187614
rect 473954 151614 474574 187058
rect 473954 151058 473986 151614
rect 474542 151058 474574 151614
rect 473954 115614 474574 151058
rect 473954 115058 473986 115614
rect 474542 115058 474574 115614
rect 473954 79614 474574 115058
rect 473954 79058 473986 79614
rect 474542 79058 474574 79614
rect 473954 43614 474574 79058
rect 473954 43058 473986 43614
rect 474542 43058 474574 43614
rect 473954 7614 474574 43058
rect 473954 7058 473986 7614
rect 474542 7058 474574 7614
rect 473954 -4186 474574 7058
rect 473954 -4742 473986 -4186
rect 474542 -4742 474574 -4186
rect 473954 -7654 474574 -4742
rect 475194 260854 475814 261216
rect 475194 260298 475226 260854
rect 475782 260298 475814 260854
rect 475194 224854 475814 260298
rect 475194 224298 475226 224854
rect 475782 224298 475814 224854
rect 475194 188854 475814 224298
rect 475194 188298 475226 188854
rect 475782 188298 475814 188854
rect 475194 152854 475814 188298
rect 475194 152298 475226 152854
rect 475782 152298 475814 152854
rect 475194 116854 475814 152298
rect 475194 116298 475226 116854
rect 475782 116298 475814 116854
rect 475194 80854 475814 116298
rect 475194 80298 475226 80854
rect 475782 80298 475814 80854
rect 475194 44854 475814 80298
rect 475194 44298 475226 44854
rect 475782 44298 475814 44854
rect 475194 8854 475814 44298
rect 475194 8298 475226 8854
rect 475782 8298 475814 8854
rect 475194 -5146 475814 8298
rect 475194 -5702 475226 -5146
rect 475782 -5702 475814 -5146
rect 475194 -7654 475814 -5702
rect 476434 226094 477054 261216
rect 476434 225538 476466 226094
rect 477022 225538 477054 226094
rect 476434 190094 477054 225538
rect 476434 189538 476466 190094
rect 477022 189538 477054 190094
rect 476434 154094 477054 189538
rect 476434 153538 476466 154094
rect 477022 153538 477054 154094
rect 476434 118094 477054 153538
rect 476434 117538 476466 118094
rect 477022 117538 477054 118094
rect 476434 82094 477054 117538
rect 476434 81538 476466 82094
rect 477022 81538 477054 82094
rect 476434 46094 477054 81538
rect 476434 45538 476466 46094
rect 477022 45538 477054 46094
rect 476434 10094 477054 45538
rect 476434 9538 476466 10094
rect 477022 9538 477054 10094
rect 476434 -6106 477054 9538
rect 476434 -6662 476466 -6106
rect 477022 -6662 477054 -6106
rect 476434 -7654 477054 -6662
rect 477674 227334 478294 261216
rect 477674 226778 477706 227334
rect 478262 226778 478294 227334
rect 477674 191334 478294 226778
rect 477674 190778 477706 191334
rect 478262 190778 478294 191334
rect 477674 155334 478294 190778
rect 477674 154778 477706 155334
rect 478262 154778 478294 155334
rect 477674 119334 478294 154778
rect 477674 118778 477706 119334
rect 478262 118778 478294 119334
rect 477674 83334 478294 118778
rect 477674 82778 477706 83334
rect 478262 82778 478294 83334
rect 477674 47334 478294 82778
rect 477674 46778 477706 47334
rect 478262 46778 478294 47334
rect 477674 11334 478294 46778
rect 477674 10778 477706 11334
rect 478262 10778 478294 11334
rect 477674 -7066 478294 10778
rect 477674 -7622 477706 -7066
rect 478262 -7622 478294 -7066
rect 477674 -7654 478294 -7622
rect 504994 254654 505614 290098
rect 504994 254098 505026 254654
rect 505582 254098 505614 254654
rect 504994 218654 505614 254098
rect 504994 218098 505026 218654
rect 505582 218098 505614 218654
rect 504994 182654 505614 218098
rect 504994 182098 505026 182654
rect 505582 182098 505614 182654
rect 504994 146654 505614 182098
rect 504994 146098 505026 146654
rect 505582 146098 505614 146654
rect 504994 110654 505614 146098
rect 504994 110098 505026 110654
rect 505582 110098 505614 110654
rect 504994 74654 505614 110098
rect 504994 74098 505026 74654
rect 505582 74098 505614 74654
rect 504994 38654 505614 74098
rect 504994 38098 505026 38654
rect 505582 38098 505614 38654
rect 504994 2654 505614 38098
rect 504994 2098 505026 2654
rect 505582 2098 505614 2654
rect 504994 -346 505614 2098
rect 504994 -902 505026 -346
rect 505582 -902 505614 -346
rect 504994 -7654 505614 -902
rect 506234 705798 506854 711590
rect 506234 705242 506266 705798
rect 506822 705242 506854 705798
rect 506234 687894 506854 705242
rect 506234 687338 506266 687894
rect 506822 687338 506854 687894
rect 506234 651894 506854 687338
rect 506234 651338 506266 651894
rect 506822 651338 506854 651894
rect 506234 615894 506854 651338
rect 506234 615338 506266 615894
rect 506822 615338 506854 615894
rect 506234 579894 506854 615338
rect 506234 579338 506266 579894
rect 506822 579338 506854 579894
rect 506234 543894 506854 579338
rect 506234 543338 506266 543894
rect 506822 543338 506854 543894
rect 506234 507894 506854 543338
rect 506234 507338 506266 507894
rect 506822 507338 506854 507894
rect 506234 471894 506854 507338
rect 506234 471338 506266 471894
rect 506822 471338 506854 471894
rect 506234 435894 506854 471338
rect 506234 435338 506266 435894
rect 506822 435338 506854 435894
rect 506234 399894 506854 435338
rect 506234 399338 506266 399894
rect 506822 399338 506854 399894
rect 506234 363894 506854 399338
rect 506234 363338 506266 363894
rect 506822 363338 506854 363894
rect 506234 327894 506854 363338
rect 506234 327338 506266 327894
rect 506822 327338 506854 327894
rect 506234 291894 506854 327338
rect 506234 291338 506266 291894
rect 506822 291338 506854 291894
rect 506234 255894 506854 291338
rect 506234 255338 506266 255894
rect 506822 255338 506854 255894
rect 506234 219894 506854 255338
rect 506234 219338 506266 219894
rect 506822 219338 506854 219894
rect 506234 183894 506854 219338
rect 506234 183338 506266 183894
rect 506822 183338 506854 183894
rect 506234 147894 506854 183338
rect 506234 147338 506266 147894
rect 506822 147338 506854 147894
rect 506234 111894 506854 147338
rect 506234 111338 506266 111894
rect 506822 111338 506854 111894
rect 506234 75894 506854 111338
rect 506234 75338 506266 75894
rect 506822 75338 506854 75894
rect 506234 39894 506854 75338
rect 506234 39338 506266 39894
rect 506822 39338 506854 39894
rect 506234 3894 506854 39338
rect 506234 3338 506266 3894
rect 506822 3338 506854 3894
rect 506234 -1306 506854 3338
rect 506234 -1862 506266 -1306
rect 506822 -1862 506854 -1306
rect 506234 -7654 506854 -1862
rect 507474 706758 508094 711590
rect 507474 706202 507506 706758
rect 508062 706202 508094 706758
rect 507474 689134 508094 706202
rect 507474 688578 507506 689134
rect 508062 688578 508094 689134
rect 507474 653134 508094 688578
rect 507474 652578 507506 653134
rect 508062 652578 508094 653134
rect 507474 617134 508094 652578
rect 507474 616578 507506 617134
rect 508062 616578 508094 617134
rect 507474 581134 508094 616578
rect 507474 580578 507506 581134
rect 508062 580578 508094 581134
rect 507474 545134 508094 580578
rect 507474 544578 507506 545134
rect 508062 544578 508094 545134
rect 507474 509134 508094 544578
rect 507474 508578 507506 509134
rect 508062 508578 508094 509134
rect 507474 473134 508094 508578
rect 507474 472578 507506 473134
rect 508062 472578 508094 473134
rect 507474 437134 508094 472578
rect 507474 436578 507506 437134
rect 508062 436578 508094 437134
rect 507474 401134 508094 436578
rect 507474 400578 507506 401134
rect 508062 400578 508094 401134
rect 507474 365134 508094 400578
rect 507474 364578 507506 365134
rect 508062 364578 508094 365134
rect 507474 329134 508094 364578
rect 507474 328578 507506 329134
rect 508062 328578 508094 329134
rect 507474 293134 508094 328578
rect 507474 292578 507506 293134
rect 508062 292578 508094 293134
rect 507474 257134 508094 292578
rect 507474 256578 507506 257134
rect 508062 256578 508094 257134
rect 507474 221134 508094 256578
rect 507474 220578 507506 221134
rect 508062 220578 508094 221134
rect 507474 185134 508094 220578
rect 507474 184578 507506 185134
rect 508062 184578 508094 185134
rect 507474 149134 508094 184578
rect 507474 148578 507506 149134
rect 508062 148578 508094 149134
rect 507474 113134 508094 148578
rect 507474 112578 507506 113134
rect 508062 112578 508094 113134
rect 507474 77134 508094 112578
rect 507474 76578 507506 77134
rect 508062 76578 508094 77134
rect 507474 41134 508094 76578
rect 507474 40578 507506 41134
rect 508062 40578 508094 41134
rect 507474 5134 508094 40578
rect 507474 4578 507506 5134
rect 508062 4578 508094 5134
rect 507474 -2266 508094 4578
rect 507474 -2822 507506 -2266
rect 508062 -2822 508094 -2266
rect 507474 -7654 508094 -2822
rect 508714 707718 509334 711590
rect 508714 707162 508746 707718
rect 509302 707162 509334 707718
rect 508714 690374 509334 707162
rect 508714 689818 508746 690374
rect 509302 689818 509334 690374
rect 508714 654374 509334 689818
rect 508714 653818 508746 654374
rect 509302 653818 509334 654374
rect 508714 618374 509334 653818
rect 508714 617818 508746 618374
rect 509302 617818 509334 618374
rect 508714 582374 509334 617818
rect 508714 581818 508746 582374
rect 509302 581818 509334 582374
rect 508714 546374 509334 581818
rect 508714 545818 508746 546374
rect 509302 545818 509334 546374
rect 508714 510374 509334 545818
rect 508714 509818 508746 510374
rect 509302 509818 509334 510374
rect 508714 474374 509334 509818
rect 508714 473818 508746 474374
rect 509302 473818 509334 474374
rect 508714 438374 509334 473818
rect 508714 437818 508746 438374
rect 509302 437818 509334 438374
rect 508714 402374 509334 437818
rect 508714 401818 508746 402374
rect 509302 401818 509334 402374
rect 508714 366374 509334 401818
rect 508714 365818 508746 366374
rect 509302 365818 509334 366374
rect 508714 330374 509334 365818
rect 508714 329818 508746 330374
rect 509302 329818 509334 330374
rect 508714 294374 509334 329818
rect 508714 293818 508746 294374
rect 509302 293818 509334 294374
rect 508714 258374 509334 293818
rect 508714 257818 508746 258374
rect 509302 257818 509334 258374
rect 508714 222374 509334 257818
rect 508714 221818 508746 222374
rect 509302 221818 509334 222374
rect 508714 186374 509334 221818
rect 508714 185818 508746 186374
rect 509302 185818 509334 186374
rect 508714 150374 509334 185818
rect 508714 149818 508746 150374
rect 509302 149818 509334 150374
rect 508714 114374 509334 149818
rect 508714 113818 508746 114374
rect 509302 113818 509334 114374
rect 508714 78374 509334 113818
rect 508714 77818 508746 78374
rect 509302 77818 509334 78374
rect 508714 42374 509334 77818
rect 508714 41818 508746 42374
rect 509302 41818 509334 42374
rect 508714 6374 509334 41818
rect 508714 5818 508746 6374
rect 509302 5818 509334 6374
rect 508714 -3226 509334 5818
rect 508714 -3782 508746 -3226
rect 509302 -3782 509334 -3226
rect 508714 -7654 509334 -3782
rect 509954 708678 510574 711590
rect 509954 708122 509986 708678
rect 510542 708122 510574 708678
rect 509954 691614 510574 708122
rect 509954 691058 509986 691614
rect 510542 691058 510574 691614
rect 509954 655614 510574 691058
rect 509954 655058 509986 655614
rect 510542 655058 510574 655614
rect 509954 619614 510574 655058
rect 509954 619058 509986 619614
rect 510542 619058 510574 619614
rect 509954 583614 510574 619058
rect 509954 583058 509986 583614
rect 510542 583058 510574 583614
rect 509954 547614 510574 583058
rect 509954 547058 509986 547614
rect 510542 547058 510574 547614
rect 509954 511614 510574 547058
rect 509954 511058 509986 511614
rect 510542 511058 510574 511614
rect 509954 475614 510574 511058
rect 509954 475058 509986 475614
rect 510542 475058 510574 475614
rect 509954 439614 510574 475058
rect 509954 439058 509986 439614
rect 510542 439058 510574 439614
rect 509954 403614 510574 439058
rect 509954 403058 509986 403614
rect 510542 403058 510574 403614
rect 509954 367614 510574 403058
rect 509954 367058 509986 367614
rect 510542 367058 510574 367614
rect 509954 331614 510574 367058
rect 509954 331058 509986 331614
rect 510542 331058 510574 331614
rect 509954 295614 510574 331058
rect 509954 295058 509986 295614
rect 510542 295058 510574 295614
rect 509954 259614 510574 295058
rect 509954 259058 509986 259614
rect 510542 259058 510574 259614
rect 509954 223614 510574 259058
rect 509954 223058 509986 223614
rect 510542 223058 510574 223614
rect 509954 187614 510574 223058
rect 509954 187058 509986 187614
rect 510542 187058 510574 187614
rect 509954 151614 510574 187058
rect 509954 151058 509986 151614
rect 510542 151058 510574 151614
rect 509954 115614 510574 151058
rect 509954 115058 509986 115614
rect 510542 115058 510574 115614
rect 509954 79614 510574 115058
rect 509954 79058 509986 79614
rect 510542 79058 510574 79614
rect 509954 43614 510574 79058
rect 509954 43058 509986 43614
rect 510542 43058 510574 43614
rect 509954 7614 510574 43058
rect 509954 7058 509986 7614
rect 510542 7058 510574 7614
rect 509954 -4186 510574 7058
rect 509954 -4742 509986 -4186
rect 510542 -4742 510574 -4186
rect 509954 -7654 510574 -4742
rect 511194 709638 511814 711590
rect 511194 709082 511226 709638
rect 511782 709082 511814 709638
rect 511194 692854 511814 709082
rect 511194 692298 511226 692854
rect 511782 692298 511814 692854
rect 511194 656854 511814 692298
rect 511194 656298 511226 656854
rect 511782 656298 511814 656854
rect 511194 620854 511814 656298
rect 511194 620298 511226 620854
rect 511782 620298 511814 620854
rect 511194 584854 511814 620298
rect 511194 584298 511226 584854
rect 511782 584298 511814 584854
rect 511194 548854 511814 584298
rect 511194 548298 511226 548854
rect 511782 548298 511814 548854
rect 511194 512854 511814 548298
rect 511194 512298 511226 512854
rect 511782 512298 511814 512854
rect 511194 476854 511814 512298
rect 511194 476298 511226 476854
rect 511782 476298 511814 476854
rect 511194 440854 511814 476298
rect 511194 440298 511226 440854
rect 511782 440298 511814 440854
rect 511194 404854 511814 440298
rect 511194 404298 511226 404854
rect 511782 404298 511814 404854
rect 511194 368854 511814 404298
rect 511194 368298 511226 368854
rect 511782 368298 511814 368854
rect 511194 332854 511814 368298
rect 511194 332298 511226 332854
rect 511782 332298 511814 332854
rect 511194 296854 511814 332298
rect 511194 296298 511226 296854
rect 511782 296298 511814 296854
rect 511194 260854 511814 296298
rect 511194 260298 511226 260854
rect 511782 260298 511814 260854
rect 511194 224854 511814 260298
rect 511194 224298 511226 224854
rect 511782 224298 511814 224854
rect 511194 188854 511814 224298
rect 511194 188298 511226 188854
rect 511782 188298 511814 188854
rect 511194 152854 511814 188298
rect 511194 152298 511226 152854
rect 511782 152298 511814 152854
rect 511194 116854 511814 152298
rect 511194 116298 511226 116854
rect 511782 116298 511814 116854
rect 511194 80854 511814 116298
rect 511194 80298 511226 80854
rect 511782 80298 511814 80854
rect 511194 44854 511814 80298
rect 511194 44298 511226 44854
rect 511782 44298 511814 44854
rect 511194 8854 511814 44298
rect 511194 8298 511226 8854
rect 511782 8298 511814 8854
rect 511194 -5146 511814 8298
rect 511194 -5702 511226 -5146
rect 511782 -5702 511814 -5146
rect 511194 -7654 511814 -5702
rect 512434 710598 513054 711590
rect 512434 710042 512466 710598
rect 513022 710042 513054 710598
rect 512434 694094 513054 710042
rect 512434 693538 512466 694094
rect 513022 693538 513054 694094
rect 512434 658094 513054 693538
rect 512434 657538 512466 658094
rect 513022 657538 513054 658094
rect 512434 622094 513054 657538
rect 512434 621538 512466 622094
rect 513022 621538 513054 622094
rect 512434 586094 513054 621538
rect 512434 585538 512466 586094
rect 513022 585538 513054 586094
rect 512434 550094 513054 585538
rect 512434 549538 512466 550094
rect 513022 549538 513054 550094
rect 512434 514094 513054 549538
rect 512434 513538 512466 514094
rect 513022 513538 513054 514094
rect 512434 478094 513054 513538
rect 512434 477538 512466 478094
rect 513022 477538 513054 478094
rect 512434 442094 513054 477538
rect 512434 441538 512466 442094
rect 513022 441538 513054 442094
rect 512434 406094 513054 441538
rect 512434 405538 512466 406094
rect 513022 405538 513054 406094
rect 512434 370094 513054 405538
rect 512434 369538 512466 370094
rect 513022 369538 513054 370094
rect 512434 334094 513054 369538
rect 512434 333538 512466 334094
rect 513022 333538 513054 334094
rect 512434 298094 513054 333538
rect 512434 297538 512466 298094
rect 513022 297538 513054 298094
rect 512434 262094 513054 297538
rect 512434 261538 512466 262094
rect 513022 261538 513054 262094
rect 512434 226094 513054 261538
rect 512434 225538 512466 226094
rect 513022 225538 513054 226094
rect 512434 190094 513054 225538
rect 512434 189538 512466 190094
rect 513022 189538 513054 190094
rect 512434 154094 513054 189538
rect 512434 153538 512466 154094
rect 513022 153538 513054 154094
rect 512434 118094 513054 153538
rect 512434 117538 512466 118094
rect 513022 117538 513054 118094
rect 512434 82094 513054 117538
rect 512434 81538 512466 82094
rect 513022 81538 513054 82094
rect 512434 46094 513054 81538
rect 512434 45538 512466 46094
rect 513022 45538 513054 46094
rect 512434 10094 513054 45538
rect 512434 9538 512466 10094
rect 513022 9538 513054 10094
rect 512434 -6106 513054 9538
rect 512434 -6662 512466 -6106
rect 513022 -6662 513054 -6106
rect 512434 -7654 513054 -6662
rect 513674 711558 514294 711590
rect 513674 711002 513706 711558
rect 514262 711002 514294 711558
rect 513674 695334 514294 711002
rect 513674 694778 513706 695334
rect 514262 694778 514294 695334
rect 513674 659334 514294 694778
rect 513674 658778 513706 659334
rect 514262 658778 514294 659334
rect 513674 623334 514294 658778
rect 513674 622778 513706 623334
rect 514262 622778 514294 623334
rect 513674 587334 514294 622778
rect 513674 586778 513706 587334
rect 514262 586778 514294 587334
rect 513674 551334 514294 586778
rect 513674 550778 513706 551334
rect 514262 550778 514294 551334
rect 513674 515334 514294 550778
rect 513674 514778 513706 515334
rect 514262 514778 514294 515334
rect 513674 479334 514294 514778
rect 513674 478778 513706 479334
rect 514262 478778 514294 479334
rect 513674 443334 514294 478778
rect 540994 704838 541614 711590
rect 540994 704282 541026 704838
rect 541582 704282 541614 704838
rect 540994 686654 541614 704282
rect 540994 686098 541026 686654
rect 541582 686098 541614 686654
rect 540994 650654 541614 686098
rect 540994 650098 541026 650654
rect 541582 650098 541614 650654
rect 540994 614654 541614 650098
rect 540994 614098 541026 614654
rect 541582 614098 541614 614654
rect 540994 578654 541614 614098
rect 540994 578098 541026 578654
rect 541582 578098 541614 578654
rect 540994 542654 541614 578098
rect 540994 542098 541026 542654
rect 541582 542098 541614 542654
rect 540994 506654 541614 542098
rect 540994 506098 541026 506654
rect 541582 506098 541614 506654
rect 540994 470654 541614 506098
rect 540994 470098 541026 470654
rect 541582 470098 541614 470654
rect 540994 445572 541614 470098
rect 542234 705798 542854 711590
rect 542234 705242 542266 705798
rect 542822 705242 542854 705798
rect 542234 687894 542854 705242
rect 542234 687338 542266 687894
rect 542822 687338 542854 687894
rect 542234 651894 542854 687338
rect 542234 651338 542266 651894
rect 542822 651338 542854 651894
rect 542234 615894 542854 651338
rect 542234 615338 542266 615894
rect 542822 615338 542854 615894
rect 542234 579894 542854 615338
rect 542234 579338 542266 579894
rect 542822 579338 542854 579894
rect 542234 543894 542854 579338
rect 542234 543338 542266 543894
rect 542822 543338 542854 543894
rect 542234 507894 542854 543338
rect 542234 507338 542266 507894
rect 542822 507338 542854 507894
rect 542234 471894 542854 507338
rect 542234 471338 542266 471894
rect 542822 471338 542854 471894
rect 542234 445572 542854 471338
rect 543474 706758 544094 711590
rect 543474 706202 543506 706758
rect 544062 706202 544094 706758
rect 543474 689134 544094 706202
rect 543474 688578 543506 689134
rect 544062 688578 544094 689134
rect 543474 653134 544094 688578
rect 543474 652578 543506 653134
rect 544062 652578 544094 653134
rect 543474 617134 544094 652578
rect 543474 616578 543506 617134
rect 544062 616578 544094 617134
rect 543474 581134 544094 616578
rect 543474 580578 543506 581134
rect 544062 580578 544094 581134
rect 543474 545134 544094 580578
rect 543474 544578 543506 545134
rect 544062 544578 544094 545134
rect 543474 509134 544094 544578
rect 543474 508578 543506 509134
rect 544062 508578 544094 509134
rect 543474 473134 544094 508578
rect 543474 472578 543506 473134
rect 544062 472578 544094 473134
rect 543474 445572 544094 472578
rect 544714 707718 545334 711590
rect 544714 707162 544746 707718
rect 545302 707162 545334 707718
rect 544714 690374 545334 707162
rect 544714 689818 544746 690374
rect 545302 689818 545334 690374
rect 544714 654374 545334 689818
rect 544714 653818 544746 654374
rect 545302 653818 545334 654374
rect 544714 618374 545334 653818
rect 544714 617818 544746 618374
rect 545302 617818 545334 618374
rect 544714 582374 545334 617818
rect 544714 581818 544746 582374
rect 545302 581818 545334 582374
rect 544714 546374 545334 581818
rect 544714 545818 544746 546374
rect 545302 545818 545334 546374
rect 544714 510374 545334 545818
rect 544714 509818 544746 510374
rect 545302 509818 545334 510374
rect 544714 474374 545334 509818
rect 544714 473818 544746 474374
rect 545302 473818 545334 474374
rect 544714 445572 545334 473818
rect 545954 708678 546574 711590
rect 545954 708122 545986 708678
rect 546542 708122 546574 708678
rect 545954 691614 546574 708122
rect 545954 691058 545986 691614
rect 546542 691058 546574 691614
rect 545954 655614 546574 691058
rect 545954 655058 545986 655614
rect 546542 655058 546574 655614
rect 545954 619614 546574 655058
rect 545954 619058 545986 619614
rect 546542 619058 546574 619614
rect 545954 583614 546574 619058
rect 545954 583058 545986 583614
rect 546542 583058 546574 583614
rect 545954 547614 546574 583058
rect 545954 547058 545986 547614
rect 546542 547058 546574 547614
rect 545954 511614 546574 547058
rect 545954 511058 545986 511614
rect 546542 511058 546574 511614
rect 545954 475614 546574 511058
rect 545954 475058 545986 475614
rect 546542 475058 546574 475614
rect 545954 445572 546574 475058
rect 547194 709638 547814 711590
rect 547194 709082 547226 709638
rect 547782 709082 547814 709638
rect 547194 692854 547814 709082
rect 547194 692298 547226 692854
rect 547782 692298 547814 692854
rect 547194 656854 547814 692298
rect 547194 656298 547226 656854
rect 547782 656298 547814 656854
rect 547194 620854 547814 656298
rect 547194 620298 547226 620854
rect 547782 620298 547814 620854
rect 547194 584854 547814 620298
rect 547194 584298 547226 584854
rect 547782 584298 547814 584854
rect 547194 548854 547814 584298
rect 547194 548298 547226 548854
rect 547782 548298 547814 548854
rect 547194 512854 547814 548298
rect 547194 512298 547226 512854
rect 547782 512298 547814 512854
rect 547194 476854 547814 512298
rect 547194 476298 547226 476854
rect 547782 476298 547814 476854
rect 513674 442778 513706 443334
rect 514262 442778 514294 443334
rect 513674 407334 514294 442778
rect 547194 440854 547814 476298
rect 547194 440298 547226 440854
rect 547782 440298 547814 440854
rect 540876 435894 541196 435926
rect 540876 435658 540918 435894
rect 541154 435658 541196 435894
rect 540876 435574 541196 435658
rect 540876 435338 540918 435574
rect 541154 435338 541196 435574
rect 540876 435306 541196 435338
rect 542808 435894 543128 435926
rect 542808 435658 542850 435894
rect 543086 435658 543128 435894
rect 542808 435574 543128 435658
rect 542808 435338 542850 435574
rect 543086 435338 543128 435574
rect 542808 435306 543128 435338
rect 544740 435894 545060 435926
rect 544740 435658 544782 435894
rect 545018 435658 545060 435894
rect 544740 435574 545060 435658
rect 544740 435338 544782 435574
rect 545018 435338 545060 435574
rect 544740 435306 545060 435338
rect 546672 435894 546992 435926
rect 546672 435658 546714 435894
rect 546950 435658 546992 435894
rect 546672 435574 546992 435658
rect 546672 435338 546714 435574
rect 546950 435338 546992 435574
rect 546672 435306 546992 435338
rect 539910 434654 540230 434686
rect 539910 434418 539952 434654
rect 540188 434418 540230 434654
rect 539910 434334 540230 434418
rect 539910 434098 539952 434334
rect 540188 434098 540230 434334
rect 539910 434066 540230 434098
rect 541842 434654 542162 434686
rect 541842 434418 541884 434654
rect 542120 434418 542162 434654
rect 541842 434334 542162 434418
rect 541842 434098 541884 434334
rect 542120 434098 542162 434334
rect 541842 434066 542162 434098
rect 543774 434654 544094 434686
rect 543774 434418 543816 434654
rect 544052 434418 544094 434654
rect 543774 434334 544094 434418
rect 543774 434098 543816 434334
rect 544052 434098 544094 434334
rect 543774 434066 544094 434098
rect 545706 434654 546026 434686
rect 545706 434418 545748 434654
rect 545984 434418 546026 434654
rect 545706 434334 546026 434418
rect 545706 434098 545748 434334
rect 545984 434098 546026 434334
rect 545706 434066 546026 434098
rect 513674 406778 513706 407334
rect 514262 406778 514294 407334
rect 513674 371334 514294 406778
rect 547194 404854 547814 440298
rect 547194 404298 547226 404854
rect 547782 404298 547814 404854
rect 540876 399894 541196 399926
rect 540876 399658 540918 399894
rect 541154 399658 541196 399894
rect 540876 399574 541196 399658
rect 540876 399338 540918 399574
rect 541154 399338 541196 399574
rect 540876 399306 541196 399338
rect 542808 399894 543128 399926
rect 542808 399658 542850 399894
rect 543086 399658 543128 399894
rect 542808 399574 543128 399658
rect 542808 399338 542850 399574
rect 543086 399338 543128 399574
rect 542808 399306 543128 399338
rect 544740 399894 545060 399926
rect 544740 399658 544782 399894
rect 545018 399658 545060 399894
rect 544740 399574 545060 399658
rect 544740 399338 544782 399574
rect 545018 399338 545060 399574
rect 544740 399306 545060 399338
rect 546672 399894 546992 399926
rect 546672 399658 546714 399894
rect 546950 399658 546992 399894
rect 546672 399574 546992 399658
rect 546672 399338 546714 399574
rect 546950 399338 546992 399574
rect 546672 399306 546992 399338
rect 539910 398654 540230 398686
rect 539910 398418 539952 398654
rect 540188 398418 540230 398654
rect 539910 398334 540230 398418
rect 539910 398098 539952 398334
rect 540188 398098 540230 398334
rect 539910 398066 540230 398098
rect 541842 398654 542162 398686
rect 541842 398418 541884 398654
rect 542120 398418 542162 398654
rect 541842 398334 542162 398418
rect 541842 398098 541884 398334
rect 542120 398098 542162 398334
rect 541842 398066 542162 398098
rect 543774 398654 544094 398686
rect 543774 398418 543816 398654
rect 544052 398418 544094 398654
rect 543774 398334 544094 398418
rect 543774 398098 543816 398334
rect 544052 398098 544094 398334
rect 543774 398066 544094 398098
rect 545706 398654 546026 398686
rect 545706 398418 545748 398654
rect 545984 398418 546026 398654
rect 545706 398334 546026 398418
rect 545706 398098 545748 398334
rect 545984 398098 546026 398334
rect 545706 398066 546026 398098
rect 513674 370778 513706 371334
rect 514262 370778 514294 371334
rect 513674 335334 514294 370778
rect 547194 368854 547814 404298
rect 547194 368298 547226 368854
rect 547782 368298 547814 368854
rect 540876 363894 541196 363926
rect 540876 363658 540918 363894
rect 541154 363658 541196 363894
rect 540876 363574 541196 363658
rect 540876 363338 540918 363574
rect 541154 363338 541196 363574
rect 540876 363306 541196 363338
rect 542808 363894 543128 363926
rect 542808 363658 542850 363894
rect 543086 363658 543128 363894
rect 542808 363574 543128 363658
rect 542808 363338 542850 363574
rect 543086 363338 543128 363574
rect 542808 363306 543128 363338
rect 544740 363894 545060 363926
rect 544740 363658 544782 363894
rect 545018 363658 545060 363894
rect 544740 363574 545060 363658
rect 544740 363338 544782 363574
rect 545018 363338 545060 363574
rect 544740 363306 545060 363338
rect 546672 363894 546992 363926
rect 546672 363658 546714 363894
rect 546950 363658 546992 363894
rect 546672 363574 546992 363658
rect 546672 363338 546714 363574
rect 546950 363338 546992 363574
rect 546672 363306 546992 363338
rect 539910 362654 540230 362686
rect 539910 362418 539952 362654
rect 540188 362418 540230 362654
rect 539910 362334 540230 362418
rect 539910 362098 539952 362334
rect 540188 362098 540230 362334
rect 539910 362066 540230 362098
rect 541842 362654 542162 362686
rect 541842 362418 541884 362654
rect 542120 362418 542162 362654
rect 541842 362334 542162 362418
rect 541842 362098 541884 362334
rect 542120 362098 542162 362334
rect 541842 362066 542162 362098
rect 543774 362654 544094 362686
rect 543774 362418 543816 362654
rect 544052 362418 544094 362654
rect 543774 362334 544094 362418
rect 543774 362098 543816 362334
rect 544052 362098 544094 362334
rect 543774 362066 544094 362098
rect 545706 362654 546026 362686
rect 545706 362418 545748 362654
rect 545984 362418 546026 362654
rect 545706 362334 546026 362418
rect 545706 362098 545748 362334
rect 545984 362098 546026 362334
rect 545706 362066 546026 362098
rect 513674 334778 513706 335334
rect 514262 334778 514294 335334
rect 513674 299334 514294 334778
rect 547194 332854 547814 368298
rect 547194 332298 547226 332854
rect 547782 332298 547814 332854
rect 540876 327894 541196 327926
rect 540876 327658 540918 327894
rect 541154 327658 541196 327894
rect 540876 327574 541196 327658
rect 540876 327338 540918 327574
rect 541154 327338 541196 327574
rect 540876 327306 541196 327338
rect 542808 327894 543128 327926
rect 542808 327658 542850 327894
rect 543086 327658 543128 327894
rect 542808 327574 543128 327658
rect 542808 327338 542850 327574
rect 543086 327338 543128 327574
rect 542808 327306 543128 327338
rect 544740 327894 545060 327926
rect 544740 327658 544782 327894
rect 545018 327658 545060 327894
rect 544740 327574 545060 327658
rect 544740 327338 544782 327574
rect 545018 327338 545060 327574
rect 544740 327306 545060 327338
rect 546672 327894 546992 327926
rect 546672 327658 546714 327894
rect 546950 327658 546992 327894
rect 546672 327574 546992 327658
rect 546672 327338 546714 327574
rect 546950 327338 546992 327574
rect 546672 327306 546992 327338
rect 539910 326654 540230 326686
rect 539910 326418 539952 326654
rect 540188 326418 540230 326654
rect 539910 326334 540230 326418
rect 539910 326098 539952 326334
rect 540188 326098 540230 326334
rect 539910 326066 540230 326098
rect 541842 326654 542162 326686
rect 541842 326418 541884 326654
rect 542120 326418 542162 326654
rect 541842 326334 542162 326418
rect 541842 326098 541884 326334
rect 542120 326098 542162 326334
rect 541842 326066 542162 326098
rect 543774 326654 544094 326686
rect 543774 326418 543816 326654
rect 544052 326418 544094 326654
rect 543774 326334 544094 326418
rect 543774 326098 543816 326334
rect 544052 326098 544094 326334
rect 543774 326066 544094 326098
rect 545706 326654 546026 326686
rect 545706 326418 545748 326654
rect 545984 326418 546026 326654
rect 545706 326334 546026 326418
rect 545706 326098 545748 326334
rect 545984 326098 546026 326334
rect 545706 326066 546026 326098
rect 513674 298778 513706 299334
rect 514262 298778 514294 299334
rect 513674 263334 514294 298778
rect 547194 296854 547814 332298
rect 547194 296298 547226 296854
rect 547782 296298 547814 296854
rect 540876 291894 541196 291926
rect 540876 291658 540918 291894
rect 541154 291658 541196 291894
rect 540876 291574 541196 291658
rect 540876 291338 540918 291574
rect 541154 291338 541196 291574
rect 540876 291306 541196 291338
rect 542808 291894 543128 291926
rect 542808 291658 542850 291894
rect 543086 291658 543128 291894
rect 542808 291574 543128 291658
rect 542808 291338 542850 291574
rect 543086 291338 543128 291574
rect 542808 291306 543128 291338
rect 544740 291894 545060 291926
rect 544740 291658 544782 291894
rect 545018 291658 545060 291894
rect 544740 291574 545060 291658
rect 544740 291338 544782 291574
rect 545018 291338 545060 291574
rect 544740 291306 545060 291338
rect 546672 291894 546992 291926
rect 546672 291658 546714 291894
rect 546950 291658 546992 291894
rect 546672 291574 546992 291658
rect 546672 291338 546714 291574
rect 546950 291338 546992 291574
rect 546672 291306 546992 291338
rect 539910 290654 540230 290686
rect 539910 290418 539952 290654
rect 540188 290418 540230 290654
rect 539910 290334 540230 290418
rect 539910 290098 539952 290334
rect 540188 290098 540230 290334
rect 539910 290066 540230 290098
rect 541842 290654 542162 290686
rect 541842 290418 541884 290654
rect 542120 290418 542162 290654
rect 541842 290334 542162 290418
rect 541842 290098 541884 290334
rect 542120 290098 542162 290334
rect 541842 290066 542162 290098
rect 543774 290654 544094 290686
rect 543774 290418 543816 290654
rect 544052 290418 544094 290654
rect 543774 290334 544094 290418
rect 543774 290098 543816 290334
rect 544052 290098 544094 290334
rect 543774 290066 544094 290098
rect 545706 290654 546026 290686
rect 545706 290418 545748 290654
rect 545984 290418 546026 290654
rect 545706 290334 546026 290418
rect 545706 290098 545748 290334
rect 545984 290098 546026 290334
rect 545706 290066 546026 290098
rect 513674 262778 513706 263334
rect 514262 262778 514294 263334
rect 513674 227334 514294 262778
rect 513674 226778 513706 227334
rect 514262 226778 514294 227334
rect 513674 191334 514294 226778
rect 513674 190778 513706 191334
rect 514262 190778 514294 191334
rect 513674 155334 514294 190778
rect 513674 154778 513706 155334
rect 514262 154778 514294 155334
rect 513674 119334 514294 154778
rect 513674 118778 513706 119334
rect 514262 118778 514294 119334
rect 513674 83334 514294 118778
rect 513674 82778 513706 83334
rect 514262 82778 514294 83334
rect 513674 47334 514294 82778
rect 513674 46778 513706 47334
rect 514262 46778 514294 47334
rect 513674 11334 514294 46778
rect 513674 10778 513706 11334
rect 514262 10778 514294 11334
rect 513674 -7066 514294 10778
rect 513674 -7622 513706 -7066
rect 514262 -7622 514294 -7066
rect 513674 -7654 514294 -7622
rect 540994 254654 541614 279788
rect 540994 254098 541026 254654
rect 541582 254098 541614 254654
rect 540994 218654 541614 254098
rect 540994 218098 541026 218654
rect 541582 218098 541614 218654
rect 540994 182654 541614 218098
rect 540994 182098 541026 182654
rect 541582 182098 541614 182654
rect 540994 146654 541614 182098
rect 540994 146098 541026 146654
rect 541582 146098 541614 146654
rect 540994 110654 541614 146098
rect 540994 110098 541026 110654
rect 541582 110098 541614 110654
rect 540994 74654 541614 110098
rect 540994 74098 541026 74654
rect 541582 74098 541614 74654
rect 540994 38654 541614 74098
rect 540994 38098 541026 38654
rect 541582 38098 541614 38654
rect 540994 2654 541614 38098
rect 540994 2098 541026 2654
rect 541582 2098 541614 2654
rect 540994 -346 541614 2098
rect 540994 -902 541026 -346
rect 541582 -902 541614 -346
rect 540994 -7654 541614 -902
rect 542234 255894 542854 279788
rect 542234 255338 542266 255894
rect 542822 255338 542854 255894
rect 542234 219894 542854 255338
rect 542234 219338 542266 219894
rect 542822 219338 542854 219894
rect 542234 183894 542854 219338
rect 542234 183338 542266 183894
rect 542822 183338 542854 183894
rect 542234 147894 542854 183338
rect 542234 147338 542266 147894
rect 542822 147338 542854 147894
rect 542234 111894 542854 147338
rect 542234 111338 542266 111894
rect 542822 111338 542854 111894
rect 542234 75894 542854 111338
rect 542234 75338 542266 75894
rect 542822 75338 542854 75894
rect 542234 39894 542854 75338
rect 542234 39338 542266 39894
rect 542822 39338 542854 39894
rect 542234 3894 542854 39338
rect 542234 3338 542266 3894
rect 542822 3338 542854 3894
rect 542234 -1306 542854 3338
rect 542234 -1862 542266 -1306
rect 542822 -1862 542854 -1306
rect 542234 -7654 542854 -1862
rect 543474 257134 544094 279788
rect 543474 256578 543506 257134
rect 544062 256578 544094 257134
rect 543474 221134 544094 256578
rect 543474 220578 543506 221134
rect 544062 220578 544094 221134
rect 543474 185134 544094 220578
rect 543474 184578 543506 185134
rect 544062 184578 544094 185134
rect 543474 149134 544094 184578
rect 543474 148578 543506 149134
rect 544062 148578 544094 149134
rect 543474 113134 544094 148578
rect 543474 112578 543506 113134
rect 544062 112578 544094 113134
rect 543474 77134 544094 112578
rect 543474 76578 543506 77134
rect 544062 76578 544094 77134
rect 543474 41134 544094 76578
rect 543474 40578 543506 41134
rect 544062 40578 544094 41134
rect 543474 5134 544094 40578
rect 543474 4578 543506 5134
rect 544062 4578 544094 5134
rect 543474 -2266 544094 4578
rect 543474 -2822 543506 -2266
rect 544062 -2822 544094 -2266
rect 543474 -7654 544094 -2822
rect 544714 258374 545334 279788
rect 544714 257818 544746 258374
rect 545302 257818 545334 258374
rect 544714 222374 545334 257818
rect 544714 221818 544746 222374
rect 545302 221818 545334 222374
rect 544714 186374 545334 221818
rect 544714 185818 544746 186374
rect 545302 185818 545334 186374
rect 544714 150374 545334 185818
rect 544714 149818 544746 150374
rect 545302 149818 545334 150374
rect 544714 114374 545334 149818
rect 544714 113818 544746 114374
rect 545302 113818 545334 114374
rect 544714 78374 545334 113818
rect 544714 77818 544746 78374
rect 545302 77818 545334 78374
rect 544714 42374 545334 77818
rect 544714 41818 544746 42374
rect 545302 41818 545334 42374
rect 544714 6374 545334 41818
rect 544714 5818 544746 6374
rect 545302 5818 545334 6374
rect 544714 -3226 545334 5818
rect 544714 -3782 544746 -3226
rect 545302 -3782 545334 -3226
rect 544714 -7654 545334 -3782
rect 545954 259614 546574 279788
rect 545954 259058 545986 259614
rect 546542 259058 546574 259614
rect 545954 223614 546574 259058
rect 545954 223058 545986 223614
rect 546542 223058 546574 223614
rect 545954 187614 546574 223058
rect 545954 187058 545986 187614
rect 546542 187058 546574 187614
rect 545954 151614 546574 187058
rect 545954 151058 545986 151614
rect 546542 151058 546574 151614
rect 545954 115614 546574 151058
rect 545954 115058 545986 115614
rect 546542 115058 546574 115614
rect 545954 79614 546574 115058
rect 545954 79058 545986 79614
rect 546542 79058 546574 79614
rect 545954 43614 546574 79058
rect 545954 43058 545986 43614
rect 546542 43058 546574 43614
rect 545954 7614 546574 43058
rect 545954 7058 545986 7614
rect 546542 7058 546574 7614
rect 545954 -4186 546574 7058
rect 545954 -4742 545986 -4186
rect 546542 -4742 546574 -4186
rect 545954 -7654 546574 -4742
rect 547194 260854 547814 296298
rect 547194 260298 547226 260854
rect 547782 260298 547814 260854
rect 547194 224854 547814 260298
rect 547194 224298 547226 224854
rect 547782 224298 547814 224854
rect 547194 188854 547814 224298
rect 547194 188298 547226 188854
rect 547782 188298 547814 188854
rect 547194 152854 547814 188298
rect 547194 152298 547226 152854
rect 547782 152298 547814 152854
rect 547194 116854 547814 152298
rect 547194 116298 547226 116854
rect 547782 116298 547814 116854
rect 547194 80854 547814 116298
rect 547194 80298 547226 80854
rect 547782 80298 547814 80854
rect 547194 44854 547814 80298
rect 547194 44298 547226 44854
rect 547782 44298 547814 44854
rect 547194 8854 547814 44298
rect 547194 8298 547226 8854
rect 547782 8298 547814 8854
rect 547194 -5146 547814 8298
rect 547194 -5702 547226 -5146
rect 547782 -5702 547814 -5146
rect 547194 -7654 547814 -5702
rect 548434 710598 549054 711590
rect 548434 710042 548466 710598
rect 549022 710042 549054 710598
rect 548434 694094 549054 710042
rect 548434 693538 548466 694094
rect 549022 693538 549054 694094
rect 548434 658094 549054 693538
rect 548434 657538 548466 658094
rect 549022 657538 549054 658094
rect 548434 622094 549054 657538
rect 548434 621538 548466 622094
rect 549022 621538 549054 622094
rect 548434 586094 549054 621538
rect 548434 585538 548466 586094
rect 549022 585538 549054 586094
rect 548434 550094 549054 585538
rect 548434 549538 548466 550094
rect 549022 549538 549054 550094
rect 548434 514094 549054 549538
rect 548434 513538 548466 514094
rect 549022 513538 549054 514094
rect 548434 478094 549054 513538
rect 548434 477538 548466 478094
rect 549022 477538 549054 478094
rect 548434 442094 549054 477538
rect 548434 441538 548466 442094
rect 549022 441538 549054 442094
rect 548434 406094 549054 441538
rect 548434 405538 548466 406094
rect 549022 405538 549054 406094
rect 548434 370094 549054 405538
rect 548434 369538 548466 370094
rect 549022 369538 549054 370094
rect 548434 334094 549054 369538
rect 548434 333538 548466 334094
rect 549022 333538 549054 334094
rect 548434 298094 549054 333538
rect 548434 297538 548466 298094
rect 549022 297538 549054 298094
rect 548434 262094 549054 297538
rect 548434 261538 548466 262094
rect 549022 261538 549054 262094
rect 548434 226094 549054 261538
rect 548434 225538 548466 226094
rect 549022 225538 549054 226094
rect 548434 190094 549054 225538
rect 548434 189538 548466 190094
rect 549022 189538 549054 190094
rect 548434 154094 549054 189538
rect 548434 153538 548466 154094
rect 549022 153538 549054 154094
rect 548434 118094 549054 153538
rect 548434 117538 548466 118094
rect 549022 117538 549054 118094
rect 548434 82094 549054 117538
rect 548434 81538 548466 82094
rect 549022 81538 549054 82094
rect 548434 46094 549054 81538
rect 548434 45538 548466 46094
rect 549022 45538 549054 46094
rect 548434 10094 549054 45538
rect 548434 9538 548466 10094
rect 549022 9538 549054 10094
rect 548434 -6106 549054 9538
rect 548434 -6662 548466 -6106
rect 549022 -6662 549054 -6106
rect 548434 -7654 549054 -6662
rect 549674 711558 550294 711590
rect 549674 711002 549706 711558
rect 550262 711002 550294 711558
rect 549674 695334 550294 711002
rect 549674 694778 549706 695334
rect 550262 694778 550294 695334
rect 549674 659334 550294 694778
rect 549674 658778 549706 659334
rect 550262 658778 550294 659334
rect 549674 623334 550294 658778
rect 549674 622778 549706 623334
rect 550262 622778 550294 623334
rect 549674 587334 550294 622778
rect 549674 586778 549706 587334
rect 550262 586778 550294 587334
rect 549674 551334 550294 586778
rect 549674 550778 549706 551334
rect 550262 550778 550294 551334
rect 549674 515334 550294 550778
rect 549674 514778 549706 515334
rect 550262 514778 550294 515334
rect 549674 479334 550294 514778
rect 549674 478778 549706 479334
rect 550262 478778 550294 479334
rect 549674 443334 550294 478778
rect 549674 442778 549706 443334
rect 550262 442778 550294 443334
rect 549674 407334 550294 442778
rect 549674 406778 549706 407334
rect 550262 406778 550294 407334
rect 549674 371334 550294 406778
rect 549674 370778 549706 371334
rect 550262 370778 550294 371334
rect 549674 335334 550294 370778
rect 549674 334778 549706 335334
rect 550262 334778 550294 335334
rect 549674 299334 550294 334778
rect 549674 298778 549706 299334
rect 550262 298778 550294 299334
rect 549674 263334 550294 298778
rect 549674 262778 549706 263334
rect 550262 262778 550294 263334
rect 549674 227334 550294 262778
rect 549674 226778 549706 227334
rect 550262 226778 550294 227334
rect 549674 191334 550294 226778
rect 549674 190778 549706 191334
rect 550262 190778 550294 191334
rect 549674 155334 550294 190778
rect 549674 154778 549706 155334
rect 550262 154778 550294 155334
rect 549674 119334 550294 154778
rect 549674 118778 549706 119334
rect 550262 118778 550294 119334
rect 549674 83334 550294 118778
rect 549674 82778 549706 83334
rect 550262 82778 550294 83334
rect 549674 47334 550294 82778
rect 549674 46778 549706 47334
rect 550262 46778 550294 47334
rect 549674 11334 550294 46778
rect 549674 10778 549706 11334
rect 550262 10778 550294 11334
rect 549674 -7066 550294 10778
rect 549674 -7622 549706 -7066
rect 550262 -7622 550294 -7066
rect 549674 -7654 550294 -7622
rect 576994 704838 577614 711590
rect 576994 704282 577026 704838
rect 577582 704282 577614 704838
rect 576994 686654 577614 704282
rect 576994 686098 577026 686654
rect 577582 686098 577614 686654
rect 576994 650654 577614 686098
rect 576994 650098 577026 650654
rect 577582 650098 577614 650654
rect 576994 614654 577614 650098
rect 576994 614098 577026 614654
rect 577582 614098 577614 614654
rect 576994 578654 577614 614098
rect 576994 578098 577026 578654
rect 577582 578098 577614 578654
rect 576994 542654 577614 578098
rect 576994 542098 577026 542654
rect 577582 542098 577614 542654
rect 576994 506654 577614 542098
rect 576994 506098 577026 506654
rect 577582 506098 577614 506654
rect 576994 470654 577614 506098
rect 576994 470098 577026 470654
rect 577582 470098 577614 470654
rect 576994 434654 577614 470098
rect 576994 434098 577026 434654
rect 577582 434098 577614 434654
rect 576994 398654 577614 434098
rect 576994 398098 577026 398654
rect 577582 398098 577614 398654
rect 576994 362654 577614 398098
rect 576994 362098 577026 362654
rect 577582 362098 577614 362654
rect 576994 326654 577614 362098
rect 576994 326098 577026 326654
rect 577582 326098 577614 326654
rect 576994 290654 577614 326098
rect 576994 290098 577026 290654
rect 577582 290098 577614 290654
rect 576994 254654 577614 290098
rect 576994 254098 577026 254654
rect 577582 254098 577614 254654
rect 576994 218654 577614 254098
rect 576994 218098 577026 218654
rect 577582 218098 577614 218654
rect 576994 182654 577614 218098
rect 576994 182098 577026 182654
rect 577582 182098 577614 182654
rect 576994 146654 577614 182098
rect 576994 146098 577026 146654
rect 577582 146098 577614 146654
rect 576994 110654 577614 146098
rect 576994 110098 577026 110654
rect 577582 110098 577614 110654
rect 576994 74654 577614 110098
rect 576994 74098 577026 74654
rect 577582 74098 577614 74654
rect 576994 38654 577614 74098
rect 576994 38098 577026 38654
rect 577582 38098 577614 38654
rect 576994 2654 577614 38098
rect 576994 2098 577026 2654
rect 577582 2098 577614 2654
rect 576994 -346 577614 2098
rect 576994 -902 577026 -346
rect 577582 -902 577614 -346
rect 576994 -7654 577614 -902
rect 578234 705798 578854 711590
rect 578234 705242 578266 705798
rect 578822 705242 578854 705798
rect 578234 687894 578854 705242
rect 578234 687338 578266 687894
rect 578822 687338 578854 687894
rect 578234 651894 578854 687338
rect 578234 651338 578266 651894
rect 578822 651338 578854 651894
rect 578234 615894 578854 651338
rect 578234 615338 578266 615894
rect 578822 615338 578854 615894
rect 578234 579894 578854 615338
rect 578234 579338 578266 579894
rect 578822 579338 578854 579894
rect 578234 543894 578854 579338
rect 578234 543338 578266 543894
rect 578822 543338 578854 543894
rect 578234 507894 578854 543338
rect 578234 507338 578266 507894
rect 578822 507338 578854 507894
rect 578234 471894 578854 507338
rect 578234 471338 578266 471894
rect 578822 471338 578854 471894
rect 578234 435894 578854 471338
rect 578234 435338 578266 435894
rect 578822 435338 578854 435894
rect 578234 399894 578854 435338
rect 578234 399338 578266 399894
rect 578822 399338 578854 399894
rect 578234 363894 578854 399338
rect 578234 363338 578266 363894
rect 578822 363338 578854 363894
rect 578234 327894 578854 363338
rect 578234 327338 578266 327894
rect 578822 327338 578854 327894
rect 578234 291894 578854 327338
rect 578234 291338 578266 291894
rect 578822 291338 578854 291894
rect 578234 255894 578854 291338
rect 578234 255338 578266 255894
rect 578822 255338 578854 255894
rect 578234 219894 578854 255338
rect 578234 219338 578266 219894
rect 578822 219338 578854 219894
rect 578234 183894 578854 219338
rect 578234 183338 578266 183894
rect 578822 183338 578854 183894
rect 578234 147894 578854 183338
rect 578234 147338 578266 147894
rect 578822 147338 578854 147894
rect 578234 111894 578854 147338
rect 578234 111338 578266 111894
rect 578822 111338 578854 111894
rect 578234 75894 578854 111338
rect 578234 75338 578266 75894
rect 578822 75338 578854 75894
rect 578234 39894 578854 75338
rect 578234 39338 578266 39894
rect 578822 39338 578854 39894
rect 578234 3894 578854 39338
rect 578234 3338 578266 3894
rect 578822 3338 578854 3894
rect 578234 -1306 578854 3338
rect 578234 -1862 578266 -1306
rect 578822 -1862 578854 -1306
rect 578234 -7654 578854 -1862
rect 579474 706758 580094 711590
rect 579474 706202 579506 706758
rect 580062 706202 580094 706758
rect 579474 689134 580094 706202
rect 579474 688578 579506 689134
rect 580062 688578 580094 689134
rect 579474 653134 580094 688578
rect 579474 652578 579506 653134
rect 580062 652578 580094 653134
rect 579474 617134 580094 652578
rect 579474 616578 579506 617134
rect 580062 616578 580094 617134
rect 579474 581134 580094 616578
rect 579474 580578 579506 581134
rect 580062 580578 580094 581134
rect 579474 545134 580094 580578
rect 579474 544578 579506 545134
rect 580062 544578 580094 545134
rect 579474 509134 580094 544578
rect 579474 508578 579506 509134
rect 580062 508578 580094 509134
rect 579474 473134 580094 508578
rect 579474 472578 579506 473134
rect 580062 472578 580094 473134
rect 579474 437134 580094 472578
rect 579474 436578 579506 437134
rect 580062 436578 580094 437134
rect 579474 401134 580094 436578
rect 579474 400578 579506 401134
rect 580062 400578 580094 401134
rect 579474 365134 580094 400578
rect 579474 364578 579506 365134
rect 580062 364578 580094 365134
rect 579474 329134 580094 364578
rect 579474 328578 579506 329134
rect 580062 328578 580094 329134
rect 579474 293134 580094 328578
rect 579474 292578 579506 293134
rect 580062 292578 580094 293134
rect 579474 257134 580094 292578
rect 579474 256578 579506 257134
rect 580062 256578 580094 257134
rect 579474 221134 580094 256578
rect 579474 220578 579506 221134
rect 580062 220578 580094 221134
rect 579474 185134 580094 220578
rect 579474 184578 579506 185134
rect 580062 184578 580094 185134
rect 579474 149134 580094 184578
rect 579474 148578 579506 149134
rect 580062 148578 580094 149134
rect 579474 113134 580094 148578
rect 579474 112578 579506 113134
rect 580062 112578 580094 113134
rect 579474 77134 580094 112578
rect 579474 76578 579506 77134
rect 580062 76578 580094 77134
rect 579474 41134 580094 76578
rect 579474 40578 579506 41134
rect 580062 40578 580094 41134
rect 579474 5134 580094 40578
rect 579474 4578 579506 5134
rect 580062 4578 580094 5134
rect 579474 -2266 580094 4578
rect 579474 -2822 579506 -2266
rect 580062 -2822 580094 -2266
rect 579474 -7654 580094 -2822
rect 580714 707718 581334 711590
rect 580714 707162 580746 707718
rect 581302 707162 581334 707718
rect 580714 690374 581334 707162
rect 580714 689818 580746 690374
rect 581302 689818 581334 690374
rect 580714 654374 581334 689818
rect 580714 653818 580746 654374
rect 581302 653818 581334 654374
rect 580714 618374 581334 653818
rect 580714 617818 580746 618374
rect 581302 617818 581334 618374
rect 580714 582374 581334 617818
rect 580714 581818 580746 582374
rect 581302 581818 581334 582374
rect 580714 546374 581334 581818
rect 580714 545818 580746 546374
rect 581302 545818 581334 546374
rect 580714 510374 581334 545818
rect 580714 509818 580746 510374
rect 581302 509818 581334 510374
rect 580714 474374 581334 509818
rect 580714 473818 580746 474374
rect 581302 473818 581334 474374
rect 580714 438374 581334 473818
rect 580714 437818 580746 438374
rect 581302 437818 581334 438374
rect 580714 402374 581334 437818
rect 580714 401818 580746 402374
rect 581302 401818 581334 402374
rect 580714 366374 581334 401818
rect 580714 365818 580746 366374
rect 581302 365818 581334 366374
rect 580714 330374 581334 365818
rect 580714 329818 580746 330374
rect 581302 329818 581334 330374
rect 580714 294374 581334 329818
rect 580714 293818 580746 294374
rect 581302 293818 581334 294374
rect 580714 258374 581334 293818
rect 580714 257818 580746 258374
rect 581302 257818 581334 258374
rect 580714 222374 581334 257818
rect 580714 221818 580746 222374
rect 581302 221818 581334 222374
rect 580714 186374 581334 221818
rect 580714 185818 580746 186374
rect 581302 185818 581334 186374
rect 580714 150374 581334 185818
rect 580714 149818 580746 150374
rect 581302 149818 581334 150374
rect 580714 114374 581334 149818
rect 580714 113818 580746 114374
rect 581302 113818 581334 114374
rect 580714 78374 581334 113818
rect 580714 77818 580746 78374
rect 581302 77818 581334 78374
rect 580714 42374 581334 77818
rect 580714 41818 580746 42374
rect 581302 41818 581334 42374
rect 580714 6374 581334 41818
rect 580714 5818 580746 6374
rect 581302 5818 581334 6374
rect 580714 -3226 581334 5818
rect 580714 -3782 580746 -3226
rect 581302 -3782 581334 -3226
rect 580714 -7654 581334 -3782
rect 581954 708678 582574 711590
rect 592030 711558 592650 711590
rect 592030 711002 592062 711558
rect 592618 711002 592650 711558
rect 591070 710598 591690 710630
rect 591070 710042 591102 710598
rect 591658 710042 591690 710598
rect 590110 709638 590730 709670
rect 590110 709082 590142 709638
rect 590698 709082 590730 709638
rect 581954 708122 581986 708678
rect 582542 708122 582574 708678
rect 581954 691614 582574 708122
rect 589150 708678 589770 708710
rect 589150 708122 589182 708678
rect 589738 708122 589770 708678
rect 588190 707718 588810 707750
rect 588190 707162 588222 707718
rect 588778 707162 588810 707718
rect 587230 706758 587850 706790
rect 587230 706202 587262 706758
rect 587818 706202 587850 706758
rect 586270 705798 586890 705830
rect 586270 705242 586302 705798
rect 586858 705242 586890 705798
rect 581954 691058 581986 691614
rect 582542 691058 582574 691614
rect 581954 655614 582574 691058
rect 581954 655058 581986 655614
rect 582542 655058 582574 655614
rect 581954 619614 582574 655058
rect 581954 619058 581986 619614
rect 582542 619058 582574 619614
rect 581954 583614 582574 619058
rect 581954 583058 581986 583614
rect 582542 583058 582574 583614
rect 581954 547614 582574 583058
rect 581954 547058 581986 547614
rect 582542 547058 582574 547614
rect 581954 511614 582574 547058
rect 581954 511058 581986 511614
rect 582542 511058 582574 511614
rect 581954 475614 582574 511058
rect 581954 475058 581986 475614
rect 582542 475058 582574 475614
rect 581954 439614 582574 475058
rect 581954 439058 581986 439614
rect 582542 439058 582574 439614
rect 581954 403614 582574 439058
rect 581954 403058 581986 403614
rect 582542 403058 582574 403614
rect 581954 367614 582574 403058
rect 581954 367058 581986 367614
rect 582542 367058 582574 367614
rect 581954 331614 582574 367058
rect 581954 331058 581986 331614
rect 582542 331058 582574 331614
rect 581954 295614 582574 331058
rect 581954 295058 581986 295614
rect 582542 295058 582574 295614
rect 581954 259614 582574 295058
rect 581954 259058 581986 259614
rect 582542 259058 582574 259614
rect 581954 223614 582574 259058
rect 581954 223058 581986 223614
rect 582542 223058 582574 223614
rect 581954 187614 582574 223058
rect 581954 187058 581986 187614
rect 582542 187058 582574 187614
rect 581954 151614 582574 187058
rect 581954 151058 581986 151614
rect 582542 151058 582574 151614
rect 581954 115614 582574 151058
rect 581954 115058 581986 115614
rect 582542 115058 582574 115614
rect 581954 79614 582574 115058
rect 581954 79058 581986 79614
rect 582542 79058 582574 79614
rect 581954 43614 582574 79058
rect 581954 43058 581986 43614
rect 582542 43058 582574 43614
rect 581954 7614 582574 43058
rect 581954 7058 581986 7614
rect 582542 7058 582574 7614
rect 581954 -4186 582574 7058
rect 585310 704838 585930 704870
rect 585310 704282 585342 704838
rect 585898 704282 585930 704838
rect 585310 686654 585930 704282
rect 585310 686098 585342 686654
rect 585898 686098 585930 686654
rect 585310 650654 585930 686098
rect 585310 650098 585342 650654
rect 585898 650098 585930 650654
rect 585310 614654 585930 650098
rect 585310 614098 585342 614654
rect 585898 614098 585930 614654
rect 585310 578654 585930 614098
rect 585310 578098 585342 578654
rect 585898 578098 585930 578654
rect 585310 542654 585930 578098
rect 585310 542098 585342 542654
rect 585898 542098 585930 542654
rect 585310 506654 585930 542098
rect 585310 506098 585342 506654
rect 585898 506098 585930 506654
rect 585310 470654 585930 506098
rect 585310 470098 585342 470654
rect 585898 470098 585930 470654
rect 585310 434654 585930 470098
rect 585310 434098 585342 434654
rect 585898 434098 585930 434654
rect 585310 398654 585930 434098
rect 585310 398098 585342 398654
rect 585898 398098 585930 398654
rect 585310 362654 585930 398098
rect 585310 362098 585342 362654
rect 585898 362098 585930 362654
rect 585310 326654 585930 362098
rect 585310 326098 585342 326654
rect 585898 326098 585930 326654
rect 585310 290654 585930 326098
rect 585310 290098 585342 290654
rect 585898 290098 585930 290654
rect 585310 254654 585930 290098
rect 585310 254098 585342 254654
rect 585898 254098 585930 254654
rect 585310 218654 585930 254098
rect 585310 218098 585342 218654
rect 585898 218098 585930 218654
rect 585310 182654 585930 218098
rect 585310 182098 585342 182654
rect 585898 182098 585930 182654
rect 585310 146654 585930 182098
rect 585310 146098 585342 146654
rect 585898 146098 585930 146654
rect 585310 110654 585930 146098
rect 585310 110098 585342 110654
rect 585898 110098 585930 110654
rect 585310 74654 585930 110098
rect 585310 74098 585342 74654
rect 585898 74098 585930 74654
rect 585310 38654 585930 74098
rect 585310 38098 585342 38654
rect 585898 38098 585930 38654
rect 585310 2654 585930 38098
rect 585310 2098 585342 2654
rect 585898 2098 585930 2654
rect 585310 -346 585930 2098
rect 585310 -902 585342 -346
rect 585898 -902 585930 -346
rect 585310 -934 585930 -902
rect 586270 687894 586890 705242
rect 586270 687338 586302 687894
rect 586858 687338 586890 687894
rect 586270 651894 586890 687338
rect 586270 651338 586302 651894
rect 586858 651338 586890 651894
rect 586270 615894 586890 651338
rect 586270 615338 586302 615894
rect 586858 615338 586890 615894
rect 586270 579894 586890 615338
rect 586270 579338 586302 579894
rect 586858 579338 586890 579894
rect 586270 543894 586890 579338
rect 586270 543338 586302 543894
rect 586858 543338 586890 543894
rect 586270 507894 586890 543338
rect 586270 507338 586302 507894
rect 586858 507338 586890 507894
rect 586270 471894 586890 507338
rect 586270 471338 586302 471894
rect 586858 471338 586890 471894
rect 586270 435894 586890 471338
rect 586270 435338 586302 435894
rect 586858 435338 586890 435894
rect 586270 399894 586890 435338
rect 586270 399338 586302 399894
rect 586858 399338 586890 399894
rect 586270 363894 586890 399338
rect 586270 363338 586302 363894
rect 586858 363338 586890 363894
rect 586270 327894 586890 363338
rect 586270 327338 586302 327894
rect 586858 327338 586890 327894
rect 586270 291894 586890 327338
rect 586270 291338 586302 291894
rect 586858 291338 586890 291894
rect 586270 255894 586890 291338
rect 586270 255338 586302 255894
rect 586858 255338 586890 255894
rect 586270 219894 586890 255338
rect 586270 219338 586302 219894
rect 586858 219338 586890 219894
rect 586270 183894 586890 219338
rect 586270 183338 586302 183894
rect 586858 183338 586890 183894
rect 586270 147894 586890 183338
rect 586270 147338 586302 147894
rect 586858 147338 586890 147894
rect 586270 111894 586890 147338
rect 586270 111338 586302 111894
rect 586858 111338 586890 111894
rect 586270 75894 586890 111338
rect 586270 75338 586302 75894
rect 586858 75338 586890 75894
rect 586270 39894 586890 75338
rect 586270 39338 586302 39894
rect 586858 39338 586890 39894
rect 586270 3894 586890 39338
rect 586270 3338 586302 3894
rect 586858 3338 586890 3894
rect 586270 -1306 586890 3338
rect 586270 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect 586270 -1894 586890 -1862
rect 587230 689134 587850 706202
rect 587230 688578 587262 689134
rect 587818 688578 587850 689134
rect 587230 653134 587850 688578
rect 587230 652578 587262 653134
rect 587818 652578 587850 653134
rect 587230 617134 587850 652578
rect 587230 616578 587262 617134
rect 587818 616578 587850 617134
rect 587230 581134 587850 616578
rect 587230 580578 587262 581134
rect 587818 580578 587850 581134
rect 587230 545134 587850 580578
rect 587230 544578 587262 545134
rect 587818 544578 587850 545134
rect 587230 509134 587850 544578
rect 587230 508578 587262 509134
rect 587818 508578 587850 509134
rect 587230 473134 587850 508578
rect 587230 472578 587262 473134
rect 587818 472578 587850 473134
rect 587230 437134 587850 472578
rect 587230 436578 587262 437134
rect 587818 436578 587850 437134
rect 587230 401134 587850 436578
rect 587230 400578 587262 401134
rect 587818 400578 587850 401134
rect 587230 365134 587850 400578
rect 587230 364578 587262 365134
rect 587818 364578 587850 365134
rect 587230 329134 587850 364578
rect 587230 328578 587262 329134
rect 587818 328578 587850 329134
rect 587230 293134 587850 328578
rect 587230 292578 587262 293134
rect 587818 292578 587850 293134
rect 587230 257134 587850 292578
rect 587230 256578 587262 257134
rect 587818 256578 587850 257134
rect 587230 221134 587850 256578
rect 587230 220578 587262 221134
rect 587818 220578 587850 221134
rect 587230 185134 587850 220578
rect 587230 184578 587262 185134
rect 587818 184578 587850 185134
rect 587230 149134 587850 184578
rect 587230 148578 587262 149134
rect 587818 148578 587850 149134
rect 587230 113134 587850 148578
rect 587230 112578 587262 113134
rect 587818 112578 587850 113134
rect 587230 77134 587850 112578
rect 587230 76578 587262 77134
rect 587818 76578 587850 77134
rect 587230 41134 587850 76578
rect 587230 40578 587262 41134
rect 587818 40578 587850 41134
rect 587230 5134 587850 40578
rect 587230 4578 587262 5134
rect 587818 4578 587850 5134
rect 587230 -2266 587850 4578
rect 587230 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect 587230 -2854 587850 -2822
rect 588190 690374 588810 707162
rect 588190 689818 588222 690374
rect 588778 689818 588810 690374
rect 588190 654374 588810 689818
rect 588190 653818 588222 654374
rect 588778 653818 588810 654374
rect 588190 618374 588810 653818
rect 588190 617818 588222 618374
rect 588778 617818 588810 618374
rect 588190 582374 588810 617818
rect 588190 581818 588222 582374
rect 588778 581818 588810 582374
rect 588190 546374 588810 581818
rect 588190 545818 588222 546374
rect 588778 545818 588810 546374
rect 588190 510374 588810 545818
rect 588190 509818 588222 510374
rect 588778 509818 588810 510374
rect 588190 474374 588810 509818
rect 588190 473818 588222 474374
rect 588778 473818 588810 474374
rect 588190 438374 588810 473818
rect 588190 437818 588222 438374
rect 588778 437818 588810 438374
rect 588190 402374 588810 437818
rect 588190 401818 588222 402374
rect 588778 401818 588810 402374
rect 588190 366374 588810 401818
rect 588190 365818 588222 366374
rect 588778 365818 588810 366374
rect 588190 330374 588810 365818
rect 588190 329818 588222 330374
rect 588778 329818 588810 330374
rect 588190 294374 588810 329818
rect 588190 293818 588222 294374
rect 588778 293818 588810 294374
rect 588190 258374 588810 293818
rect 588190 257818 588222 258374
rect 588778 257818 588810 258374
rect 588190 222374 588810 257818
rect 588190 221818 588222 222374
rect 588778 221818 588810 222374
rect 588190 186374 588810 221818
rect 588190 185818 588222 186374
rect 588778 185818 588810 186374
rect 588190 150374 588810 185818
rect 588190 149818 588222 150374
rect 588778 149818 588810 150374
rect 588190 114374 588810 149818
rect 588190 113818 588222 114374
rect 588778 113818 588810 114374
rect 588190 78374 588810 113818
rect 588190 77818 588222 78374
rect 588778 77818 588810 78374
rect 588190 42374 588810 77818
rect 588190 41818 588222 42374
rect 588778 41818 588810 42374
rect 588190 6374 588810 41818
rect 588190 5818 588222 6374
rect 588778 5818 588810 6374
rect 588190 -3226 588810 5818
rect 588190 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect 588190 -3814 588810 -3782
rect 589150 691614 589770 708122
rect 589150 691058 589182 691614
rect 589738 691058 589770 691614
rect 589150 655614 589770 691058
rect 589150 655058 589182 655614
rect 589738 655058 589770 655614
rect 589150 619614 589770 655058
rect 589150 619058 589182 619614
rect 589738 619058 589770 619614
rect 589150 583614 589770 619058
rect 589150 583058 589182 583614
rect 589738 583058 589770 583614
rect 589150 547614 589770 583058
rect 589150 547058 589182 547614
rect 589738 547058 589770 547614
rect 589150 511614 589770 547058
rect 589150 511058 589182 511614
rect 589738 511058 589770 511614
rect 589150 475614 589770 511058
rect 589150 475058 589182 475614
rect 589738 475058 589770 475614
rect 589150 439614 589770 475058
rect 589150 439058 589182 439614
rect 589738 439058 589770 439614
rect 589150 403614 589770 439058
rect 589150 403058 589182 403614
rect 589738 403058 589770 403614
rect 589150 367614 589770 403058
rect 589150 367058 589182 367614
rect 589738 367058 589770 367614
rect 589150 331614 589770 367058
rect 589150 331058 589182 331614
rect 589738 331058 589770 331614
rect 589150 295614 589770 331058
rect 589150 295058 589182 295614
rect 589738 295058 589770 295614
rect 589150 259614 589770 295058
rect 589150 259058 589182 259614
rect 589738 259058 589770 259614
rect 589150 223614 589770 259058
rect 589150 223058 589182 223614
rect 589738 223058 589770 223614
rect 589150 187614 589770 223058
rect 589150 187058 589182 187614
rect 589738 187058 589770 187614
rect 589150 151614 589770 187058
rect 589150 151058 589182 151614
rect 589738 151058 589770 151614
rect 589150 115614 589770 151058
rect 589150 115058 589182 115614
rect 589738 115058 589770 115614
rect 589150 79614 589770 115058
rect 589150 79058 589182 79614
rect 589738 79058 589770 79614
rect 589150 43614 589770 79058
rect 589150 43058 589182 43614
rect 589738 43058 589770 43614
rect 589150 7614 589770 43058
rect 589150 7058 589182 7614
rect 589738 7058 589770 7614
rect 581954 -4742 581986 -4186
rect 582542 -4742 582574 -4186
rect 581954 -7654 582574 -4742
rect 589150 -4186 589770 7058
rect 589150 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect 589150 -4774 589770 -4742
rect 590110 692854 590730 709082
rect 590110 692298 590142 692854
rect 590698 692298 590730 692854
rect 590110 656854 590730 692298
rect 590110 656298 590142 656854
rect 590698 656298 590730 656854
rect 590110 620854 590730 656298
rect 590110 620298 590142 620854
rect 590698 620298 590730 620854
rect 590110 584854 590730 620298
rect 590110 584298 590142 584854
rect 590698 584298 590730 584854
rect 590110 548854 590730 584298
rect 590110 548298 590142 548854
rect 590698 548298 590730 548854
rect 590110 512854 590730 548298
rect 590110 512298 590142 512854
rect 590698 512298 590730 512854
rect 590110 476854 590730 512298
rect 590110 476298 590142 476854
rect 590698 476298 590730 476854
rect 590110 440854 590730 476298
rect 590110 440298 590142 440854
rect 590698 440298 590730 440854
rect 590110 404854 590730 440298
rect 590110 404298 590142 404854
rect 590698 404298 590730 404854
rect 590110 368854 590730 404298
rect 590110 368298 590142 368854
rect 590698 368298 590730 368854
rect 590110 332854 590730 368298
rect 590110 332298 590142 332854
rect 590698 332298 590730 332854
rect 590110 296854 590730 332298
rect 590110 296298 590142 296854
rect 590698 296298 590730 296854
rect 590110 260854 590730 296298
rect 590110 260298 590142 260854
rect 590698 260298 590730 260854
rect 590110 224854 590730 260298
rect 590110 224298 590142 224854
rect 590698 224298 590730 224854
rect 590110 188854 590730 224298
rect 590110 188298 590142 188854
rect 590698 188298 590730 188854
rect 590110 152854 590730 188298
rect 590110 152298 590142 152854
rect 590698 152298 590730 152854
rect 590110 116854 590730 152298
rect 590110 116298 590142 116854
rect 590698 116298 590730 116854
rect 590110 80854 590730 116298
rect 590110 80298 590142 80854
rect 590698 80298 590730 80854
rect 590110 44854 590730 80298
rect 590110 44298 590142 44854
rect 590698 44298 590730 44854
rect 590110 8854 590730 44298
rect 590110 8298 590142 8854
rect 590698 8298 590730 8854
rect 590110 -5146 590730 8298
rect 590110 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect 590110 -5734 590730 -5702
rect 591070 694094 591690 710042
rect 591070 693538 591102 694094
rect 591658 693538 591690 694094
rect 591070 658094 591690 693538
rect 591070 657538 591102 658094
rect 591658 657538 591690 658094
rect 591070 622094 591690 657538
rect 591070 621538 591102 622094
rect 591658 621538 591690 622094
rect 591070 586094 591690 621538
rect 591070 585538 591102 586094
rect 591658 585538 591690 586094
rect 591070 550094 591690 585538
rect 591070 549538 591102 550094
rect 591658 549538 591690 550094
rect 591070 514094 591690 549538
rect 591070 513538 591102 514094
rect 591658 513538 591690 514094
rect 591070 478094 591690 513538
rect 591070 477538 591102 478094
rect 591658 477538 591690 478094
rect 591070 442094 591690 477538
rect 591070 441538 591102 442094
rect 591658 441538 591690 442094
rect 591070 406094 591690 441538
rect 591070 405538 591102 406094
rect 591658 405538 591690 406094
rect 591070 370094 591690 405538
rect 591070 369538 591102 370094
rect 591658 369538 591690 370094
rect 591070 334094 591690 369538
rect 591070 333538 591102 334094
rect 591658 333538 591690 334094
rect 591070 298094 591690 333538
rect 591070 297538 591102 298094
rect 591658 297538 591690 298094
rect 591070 262094 591690 297538
rect 591070 261538 591102 262094
rect 591658 261538 591690 262094
rect 591070 226094 591690 261538
rect 591070 225538 591102 226094
rect 591658 225538 591690 226094
rect 591070 190094 591690 225538
rect 591070 189538 591102 190094
rect 591658 189538 591690 190094
rect 591070 154094 591690 189538
rect 591070 153538 591102 154094
rect 591658 153538 591690 154094
rect 591070 118094 591690 153538
rect 591070 117538 591102 118094
rect 591658 117538 591690 118094
rect 591070 82094 591690 117538
rect 591070 81538 591102 82094
rect 591658 81538 591690 82094
rect 591070 46094 591690 81538
rect 591070 45538 591102 46094
rect 591658 45538 591690 46094
rect 591070 10094 591690 45538
rect 591070 9538 591102 10094
rect 591658 9538 591690 10094
rect 591070 -6106 591690 9538
rect 591070 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect 591070 -6694 591690 -6662
rect 592030 695334 592650 711002
rect 592030 694778 592062 695334
rect 592618 694778 592650 695334
rect 592030 659334 592650 694778
rect 592030 658778 592062 659334
rect 592618 658778 592650 659334
rect 592030 623334 592650 658778
rect 592030 622778 592062 623334
rect 592618 622778 592650 623334
rect 592030 587334 592650 622778
rect 592030 586778 592062 587334
rect 592618 586778 592650 587334
rect 592030 551334 592650 586778
rect 592030 550778 592062 551334
rect 592618 550778 592650 551334
rect 592030 515334 592650 550778
rect 592030 514778 592062 515334
rect 592618 514778 592650 515334
rect 592030 479334 592650 514778
rect 592030 478778 592062 479334
rect 592618 478778 592650 479334
rect 592030 443334 592650 478778
rect 592030 442778 592062 443334
rect 592618 442778 592650 443334
rect 592030 407334 592650 442778
rect 592030 406778 592062 407334
rect 592618 406778 592650 407334
rect 592030 371334 592650 406778
rect 592030 370778 592062 371334
rect 592618 370778 592650 371334
rect 592030 335334 592650 370778
rect 592030 334778 592062 335334
rect 592618 334778 592650 335334
rect 592030 299334 592650 334778
rect 592030 298778 592062 299334
rect 592618 298778 592650 299334
rect 592030 263334 592650 298778
rect 592030 262778 592062 263334
rect 592618 262778 592650 263334
rect 592030 227334 592650 262778
rect 592030 226778 592062 227334
rect 592618 226778 592650 227334
rect 592030 191334 592650 226778
rect 592030 190778 592062 191334
rect 592618 190778 592650 191334
rect 592030 155334 592650 190778
rect 592030 154778 592062 155334
rect 592618 154778 592650 155334
rect 592030 119334 592650 154778
rect 592030 118778 592062 119334
rect 592618 118778 592650 119334
rect 592030 83334 592650 118778
rect 592030 82778 592062 83334
rect 592618 82778 592650 83334
rect 592030 47334 592650 82778
rect 592030 46778 592062 47334
rect 592618 46778 592650 47334
rect 592030 11334 592650 46778
rect 592030 10778 592062 11334
rect 592618 10778 592650 11334
rect 592030 -7066 592650 10778
rect 592030 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711002 -8138 711558
rect -8694 694778 -8138 695334
rect -8694 658778 -8138 659334
rect -8694 622778 -8138 623334
rect -8694 586778 -8138 587334
rect -8694 550778 -8138 551334
rect -8694 514778 -8138 515334
rect -8694 478778 -8138 479334
rect -8694 442778 -8138 443334
rect -8694 406778 -8138 407334
rect -8694 370778 -8138 371334
rect -8694 334778 -8138 335334
rect -8694 298778 -8138 299334
rect -8694 262778 -8138 263334
rect -8694 226778 -8138 227334
rect -8694 190778 -8138 191334
rect -8694 154778 -8138 155334
rect -8694 118778 -8138 119334
rect -8694 82778 -8138 83334
rect -8694 46778 -8138 47334
rect -8694 10778 -8138 11334
rect -7734 710042 -7178 710598
rect -7734 693538 -7178 694094
rect -7734 657538 -7178 658094
rect -7734 621538 -7178 622094
rect -7734 585538 -7178 586094
rect -7734 549538 -7178 550094
rect -7734 513538 -7178 514094
rect -7734 477538 -7178 478094
rect -7734 441538 -7178 442094
rect -7734 405538 -7178 406094
rect -7734 369538 -7178 370094
rect -7734 333538 -7178 334094
rect -7734 297538 -7178 298094
rect -7734 261538 -7178 262094
rect -7734 225538 -7178 226094
rect -7734 189538 -7178 190094
rect -7734 153538 -7178 154094
rect -7734 117538 -7178 118094
rect -7734 81538 -7178 82094
rect -7734 45538 -7178 46094
rect -7734 9538 -7178 10094
rect -6774 709082 -6218 709638
rect -6774 692298 -6218 692854
rect -6774 656298 -6218 656854
rect -6774 620298 -6218 620854
rect -6774 584298 -6218 584854
rect -6774 548298 -6218 548854
rect -6774 512298 -6218 512854
rect -6774 476298 -6218 476854
rect -6774 440298 -6218 440854
rect -6774 404298 -6218 404854
rect -6774 368298 -6218 368854
rect -6774 332298 -6218 332854
rect -6774 296298 -6218 296854
rect -6774 260298 -6218 260854
rect -6774 224298 -6218 224854
rect -6774 188298 -6218 188854
rect -6774 152298 -6218 152854
rect -6774 116298 -6218 116854
rect -6774 80298 -6218 80854
rect -6774 44298 -6218 44854
rect -6774 8298 -6218 8854
rect -5814 708122 -5258 708678
rect -5814 691058 -5258 691614
rect -5814 655058 -5258 655614
rect -5814 619058 -5258 619614
rect -5814 583058 -5258 583614
rect -5814 547058 -5258 547614
rect -5814 511058 -5258 511614
rect -5814 475058 -5258 475614
rect -5814 439058 -5258 439614
rect -5814 403058 -5258 403614
rect -5814 367058 -5258 367614
rect -5814 331058 -5258 331614
rect -5814 295058 -5258 295614
rect -5814 259058 -5258 259614
rect -5814 223058 -5258 223614
rect -5814 187058 -5258 187614
rect -5814 151058 -5258 151614
rect -5814 115058 -5258 115614
rect -5814 79058 -5258 79614
rect -5814 43058 -5258 43614
rect -5814 7058 -5258 7614
rect -4854 707162 -4298 707718
rect -4854 689818 -4298 690374
rect -4854 653818 -4298 654374
rect -4854 617818 -4298 618374
rect -4854 581818 -4298 582374
rect -4854 545818 -4298 546374
rect -4854 509818 -4298 510374
rect -4854 473818 -4298 474374
rect -4854 437818 -4298 438374
rect -4854 401818 -4298 402374
rect -4854 365818 -4298 366374
rect -4854 329818 -4298 330374
rect -4854 293818 -4298 294374
rect -4854 257818 -4298 258374
rect -4854 221818 -4298 222374
rect -4854 185818 -4298 186374
rect -4854 149818 -4298 150374
rect -4854 113818 -4298 114374
rect -4854 77818 -4298 78374
rect -4854 41818 -4298 42374
rect -4854 5818 -4298 6374
rect -3894 706202 -3338 706758
rect -3894 688578 -3338 689134
rect -3894 652578 -3338 653134
rect -3894 616578 -3338 617134
rect -3894 580578 -3338 581134
rect -3894 544578 -3338 545134
rect -3894 508578 -3338 509134
rect -3894 472578 -3338 473134
rect -3894 436578 -3338 437134
rect -3894 400578 -3338 401134
rect -3894 364578 -3338 365134
rect -3894 328578 -3338 329134
rect -3894 292578 -3338 293134
rect -3894 256578 -3338 257134
rect -3894 220578 -3338 221134
rect -3894 184578 -3338 185134
rect -3894 148578 -3338 149134
rect -3894 112578 -3338 113134
rect -3894 76578 -3338 77134
rect -3894 40578 -3338 41134
rect -3894 4578 -3338 5134
rect -2934 705242 -2378 705798
rect -2934 687338 -2378 687894
rect -2934 651338 -2378 651894
rect -2934 615338 -2378 615894
rect -2934 579338 -2378 579894
rect -2934 543338 -2378 543894
rect -2934 507338 -2378 507894
rect -2934 471338 -2378 471894
rect -2934 435338 -2378 435894
rect -2934 399338 -2378 399894
rect -2934 363338 -2378 363894
rect -2934 327338 -2378 327894
rect -2934 291338 -2378 291894
rect -2934 255338 -2378 255894
rect -2934 219338 -2378 219894
rect -2934 183338 -2378 183894
rect -2934 147338 -2378 147894
rect -2934 111338 -2378 111894
rect -2934 75338 -2378 75894
rect -2934 39338 -2378 39894
rect -2934 3338 -2378 3894
rect -1974 704282 -1418 704838
rect -1974 686098 -1418 686654
rect -1974 650098 -1418 650654
rect -1974 614098 -1418 614654
rect -1974 578098 -1418 578654
rect -1974 542098 -1418 542654
rect -1974 506098 -1418 506654
rect -1974 470098 -1418 470654
rect -1974 434098 -1418 434654
rect -1974 398098 -1418 398654
rect -1974 362098 -1418 362654
rect -1974 326098 -1418 326654
rect -1974 290098 -1418 290654
rect -1974 254098 -1418 254654
rect -1974 218098 -1418 218654
rect -1974 182098 -1418 182654
rect -1974 146098 -1418 146654
rect -1974 110098 -1418 110654
rect -1974 74098 -1418 74654
rect -1974 38098 -1418 38654
rect -1974 2098 -1418 2654
rect -1974 -902 -1418 -346
rect 1026 704282 1582 704838
rect 1026 686098 1582 686654
rect 1026 650098 1582 650654
rect 1026 614098 1582 614654
rect 1026 578098 1582 578654
rect 1026 542098 1582 542654
rect 1026 506098 1582 506654
rect 1026 470098 1582 470654
rect 1026 434098 1582 434654
rect 1026 398098 1582 398654
rect 1026 362098 1582 362654
rect 1026 326098 1582 326654
rect 1026 290098 1582 290654
rect 1026 254098 1582 254654
rect 1026 218098 1582 218654
rect 1026 182098 1582 182654
rect 1026 146098 1582 146654
rect 1026 110098 1582 110654
rect 1026 74098 1582 74654
rect 1026 38098 1582 38654
rect 1026 2098 1582 2654
rect 1026 -902 1582 -346
rect -2934 -1862 -2378 -1306
rect -3894 -2822 -3338 -2266
rect -4854 -3782 -4298 -3226
rect -5814 -4742 -5258 -4186
rect -6774 -5702 -6218 -5146
rect -7734 -6662 -7178 -6106
rect -8694 -7622 -8138 -7066
rect 2266 705242 2822 705798
rect 2266 687338 2822 687894
rect 2266 651338 2822 651894
rect 2266 615338 2822 615894
rect 2266 579338 2822 579894
rect 2266 543338 2822 543894
rect 2266 507338 2822 507894
rect 2266 471338 2822 471894
rect 2266 435338 2822 435894
rect 2266 399338 2822 399894
rect 2266 363338 2822 363894
rect 2266 327338 2822 327894
rect 2266 291338 2822 291894
rect 2266 255338 2822 255894
rect 2266 219338 2822 219894
rect 2266 183338 2822 183894
rect 2266 147338 2822 147894
rect 2266 111338 2822 111894
rect 2266 75338 2822 75894
rect 2266 39338 2822 39894
rect 2266 3338 2822 3894
rect 2266 -1862 2822 -1306
rect 3506 706202 4062 706758
rect 3506 688578 4062 689134
rect 3506 652578 4062 653134
rect 3506 616578 4062 617134
rect 3506 580578 4062 581134
rect 3506 544578 4062 545134
rect 3506 508578 4062 509134
rect 3506 472578 4062 473134
rect 3506 436578 4062 437134
rect 3506 400578 4062 401134
rect 3506 364578 4062 365134
rect 3506 328578 4062 329134
rect 3506 292578 4062 293134
rect 3506 256578 4062 257134
rect 3506 220578 4062 221134
rect 3506 184578 4062 185134
rect 3506 148578 4062 149134
rect 3506 112578 4062 113134
rect 3506 76578 4062 77134
rect 3506 40578 4062 41134
rect 3506 4578 4062 5134
rect 3506 -2822 4062 -2266
rect 4746 707162 5302 707718
rect 4746 689818 5302 690374
rect 4746 653818 5302 654374
rect 4746 617818 5302 618374
rect 4746 581818 5302 582374
rect 4746 545818 5302 546374
rect 4746 509818 5302 510374
rect 4746 473818 5302 474374
rect 4746 437818 5302 438374
rect 4746 401818 5302 402374
rect 4746 365818 5302 366374
rect 4746 329818 5302 330374
rect 4746 293818 5302 294374
rect 4746 257818 5302 258374
rect 4746 221818 5302 222374
rect 4746 185818 5302 186374
rect 4746 149818 5302 150374
rect 4746 113818 5302 114374
rect 4746 77818 5302 78374
rect 4746 41818 5302 42374
rect 4746 5818 5302 6374
rect 4746 -3782 5302 -3226
rect 5986 708122 6542 708678
rect 5986 691058 6542 691614
rect 5986 655058 6542 655614
rect 5986 619058 6542 619614
rect 5986 583058 6542 583614
rect 5986 547058 6542 547614
rect 5986 511058 6542 511614
rect 5986 475058 6542 475614
rect 5986 439058 6542 439614
rect 5986 403058 6542 403614
rect 5986 367058 6542 367614
rect 5986 331058 6542 331614
rect 5986 295058 6542 295614
rect 5986 259058 6542 259614
rect 5986 223058 6542 223614
rect 5986 187058 6542 187614
rect 5986 151058 6542 151614
rect 5986 115058 6542 115614
rect 5986 79058 6542 79614
rect 5986 43058 6542 43614
rect 5986 7058 6542 7614
rect 5986 -4742 6542 -4186
rect 7226 709082 7782 709638
rect 7226 692298 7782 692854
rect 7226 656298 7782 656854
rect 7226 620298 7782 620854
rect 7226 584298 7782 584854
rect 7226 548298 7782 548854
rect 7226 512298 7782 512854
rect 7226 476298 7782 476854
rect 7226 440298 7782 440854
rect 7226 404298 7782 404854
rect 7226 368298 7782 368854
rect 7226 332298 7782 332854
rect 7226 296298 7782 296854
rect 7226 260298 7782 260854
rect 7226 224298 7782 224854
rect 7226 188298 7782 188854
rect 7226 152298 7782 152854
rect 7226 116298 7782 116854
rect 7226 80298 7782 80854
rect 7226 44298 7782 44854
rect 7226 8298 7782 8854
rect 7226 -5702 7782 -5146
rect 8466 710042 9022 710598
rect 8466 693538 9022 694094
rect 8466 657538 9022 658094
rect 8466 621538 9022 622094
rect 8466 585538 9022 586094
rect 8466 549538 9022 550094
rect 8466 513538 9022 514094
rect 8466 477538 9022 478094
rect 8466 441538 9022 442094
rect 8466 405538 9022 406094
rect 8466 369538 9022 370094
rect 8466 333538 9022 334094
rect 8466 297538 9022 298094
rect 8466 261538 9022 262094
rect 8466 225538 9022 226094
rect 8466 189538 9022 190094
rect 8466 153538 9022 154094
rect 8466 117538 9022 118094
rect 8466 81538 9022 82094
rect 8466 45538 9022 46094
rect 8466 9538 9022 10094
rect 8466 -6662 9022 -6106
rect 9706 711002 10262 711558
rect 9706 694778 10262 695334
rect 9706 658778 10262 659334
rect 9706 622778 10262 623334
rect 9706 586778 10262 587334
rect 9706 550778 10262 551334
rect 9706 514778 10262 515334
rect 9706 478778 10262 479334
rect 9706 442778 10262 443334
rect 9706 406778 10262 407334
rect 9706 370778 10262 371334
rect 9706 334778 10262 335334
rect 9706 298778 10262 299334
rect 9706 262778 10262 263334
rect 9706 226778 10262 227334
rect 9706 190778 10262 191334
rect 9706 154778 10262 155334
rect 9706 118778 10262 119334
rect 9706 82778 10262 83334
rect 9706 46778 10262 47334
rect 9706 10778 10262 11334
rect 9706 -7622 10262 -7066
rect 37026 704282 37582 704838
rect 37026 686098 37582 686654
rect 37026 650098 37582 650654
rect 37026 614098 37582 614654
rect 37026 578098 37582 578654
rect 37026 542098 37582 542654
rect 37026 506098 37582 506654
rect 37026 470098 37582 470654
rect 37026 434098 37582 434654
rect 37026 398098 37582 398654
rect 37026 362098 37582 362654
rect 37026 326098 37582 326654
rect 37026 290098 37582 290654
rect 37026 254098 37582 254654
rect 37026 218098 37582 218654
rect 37026 182098 37582 182654
rect 37026 146098 37582 146654
rect 37026 110098 37582 110654
rect 37026 74098 37582 74654
rect 37026 38098 37582 38654
rect 37026 2098 37582 2654
rect 37026 -902 37582 -346
rect 38266 705242 38822 705798
rect 38266 687338 38822 687894
rect 38266 651338 38822 651894
rect 38266 615338 38822 615894
rect 38266 579338 38822 579894
rect 38266 543338 38822 543894
rect 38266 507338 38822 507894
rect 38266 471338 38822 471894
rect 38266 435338 38822 435894
rect 38266 399338 38822 399894
rect 38266 363338 38822 363894
rect 38266 327338 38822 327894
rect 38266 291338 38822 291894
rect 38266 255338 38822 255894
rect 38266 219338 38822 219894
rect 38266 183338 38822 183894
rect 38266 147338 38822 147894
rect 38266 111338 38822 111894
rect 38266 75338 38822 75894
rect 38266 39338 38822 39894
rect 38266 3338 38822 3894
rect 38266 -1862 38822 -1306
rect 39506 706202 40062 706758
rect 39506 688578 40062 689134
rect 39506 652578 40062 653134
rect 39506 616578 40062 617134
rect 39506 580578 40062 581134
rect 39506 544578 40062 545134
rect 39506 508578 40062 509134
rect 39506 472578 40062 473134
rect 39506 436578 40062 437134
rect 39506 400578 40062 401134
rect 39506 364578 40062 365134
rect 39506 328578 40062 329134
rect 39506 292578 40062 293134
rect 39506 256578 40062 257134
rect 39506 220578 40062 221134
rect 39506 184578 40062 185134
rect 39506 148578 40062 149134
rect 39506 112578 40062 113134
rect 39506 76578 40062 77134
rect 39506 40578 40062 41134
rect 39506 4578 40062 5134
rect 39506 -2822 40062 -2266
rect 40746 707162 41302 707718
rect 40746 689818 41302 690374
rect 40746 653818 41302 654374
rect 40746 617818 41302 618374
rect 40746 581818 41302 582374
rect 40746 545818 41302 546374
rect 40746 509818 41302 510374
rect 40746 473818 41302 474374
rect 40746 437818 41302 438374
rect 40746 401818 41302 402374
rect 40746 365818 41302 366374
rect 40746 329818 41302 330374
rect 40746 293818 41302 294374
rect 40746 257818 41302 258374
rect 40746 221818 41302 222374
rect 40746 185818 41302 186374
rect 40746 149818 41302 150374
rect 40746 113818 41302 114374
rect 40746 77818 41302 78374
rect 40746 41818 41302 42374
rect 40746 5818 41302 6374
rect 40746 -3782 41302 -3226
rect 41986 708122 42542 708678
rect 41986 691058 42542 691614
rect 41986 655058 42542 655614
rect 41986 619058 42542 619614
rect 41986 583058 42542 583614
rect 41986 547058 42542 547614
rect 41986 511058 42542 511614
rect 41986 475058 42542 475614
rect 41986 439058 42542 439614
rect 41986 403058 42542 403614
rect 41986 367058 42542 367614
rect 41986 331058 42542 331614
rect 41986 295058 42542 295614
rect 41986 259058 42542 259614
rect 41986 223058 42542 223614
rect 41986 187058 42542 187614
rect 41986 151058 42542 151614
rect 41986 115058 42542 115614
rect 41986 79058 42542 79614
rect 41986 43058 42542 43614
rect 41986 7058 42542 7614
rect 41986 -4742 42542 -4186
rect 43226 709082 43782 709638
rect 43226 692298 43782 692854
rect 43226 656298 43782 656854
rect 43226 620298 43782 620854
rect 43226 584298 43782 584854
rect 43226 548298 43782 548854
rect 43226 512298 43782 512854
rect 43226 476298 43782 476854
rect 43226 440298 43782 440854
rect 43226 404298 43782 404854
rect 43226 368298 43782 368854
rect 43226 332298 43782 332854
rect 43226 296298 43782 296854
rect 43226 260298 43782 260854
rect 43226 224298 43782 224854
rect 43226 188298 43782 188854
rect 43226 152298 43782 152854
rect 43226 116298 43782 116854
rect 43226 80298 43782 80854
rect 43226 44298 43782 44854
rect 43226 8298 43782 8854
rect 43226 -5702 43782 -5146
rect 44466 710042 45022 710598
rect 44466 693538 45022 694094
rect 44466 657538 45022 658094
rect 44466 621538 45022 622094
rect 44466 585538 45022 586094
rect 44466 549538 45022 550094
rect 44466 513538 45022 514094
rect 44466 477538 45022 478094
rect 44466 441538 45022 442094
rect 44466 405538 45022 406094
rect 44466 369538 45022 370094
rect 44466 333538 45022 334094
rect 44466 297538 45022 298094
rect 44466 261538 45022 262094
rect 44466 225538 45022 226094
rect 44466 189538 45022 190094
rect 44466 153538 45022 154094
rect 44466 117538 45022 118094
rect 44466 81538 45022 82094
rect 44466 45538 45022 46094
rect 44466 9538 45022 10094
rect 44466 -6662 45022 -6106
rect 45706 711002 46262 711558
rect 45706 694778 46262 695334
rect 45706 658778 46262 659334
rect 45706 622778 46262 623334
rect 45706 586778 46262 587334
rect 45706 550778 46262 551334
rect 45706 514778 46262 515334
rect 45706 478778 46262 479334
rect 45706 442778 46262 443334
rect 45706 406778 46262 407334
rect 45706 370778 46262 371334
rect 45706 334778 46262 335334
rect 45706 298778 46262 299334
rect 45706 262778 46262 263334
rect 45706 226778 46262 227334
rect 45706 190778 46262 191334
rect 45706 154778 46262 155334
rect 45706 118778 46262 119334
rect 45706 82778 46262 83334
rect 45706 46778 46262 47334
rect 45706 10778 46262 11334
rect 45706 -7622 46262 -7066
rect 73026 704282 73582 704838
rect 73026 686098 73582 686654
rect 73026 650098 73582 650654
rect 73026 614098 73582 614654
rect 73026 578098 73582 578654
rect 73026 542098 73582 542654
rect 73026 506098 73582 506654
rect 73026 470098 73582 470654
rect 73026 434098 73582 434654
rect 73026 398098 73582 398654
rect 73026 362098 73582 362654
rect 73026 326098 73582 326654
rect 73026 290098 73582 290654
rect 73026 254098 73582 254654
rect 73026 218098 73582 218654
rect 73026 182098 73582 182654
rect 73026 146098 73582 146654
rect 73026 110098 73582 110654
rect 73026 74098 73582 74654
rect 73026 38098 73582 38654
rect 73026 2098 73582 2654
rect 73026 -902 73582 -346
rect 74266 705242 74822 705798
rect 74266 687338 74822 687894
rect 74266 651338 74822 651894
rect 74266 615338 74822 615894
rect 74266 579338 74822 579894
rect 74266 543338 74822 543894
rect 74266 507338 74822 507894
rect 74266 471338 74822 471894
rect 74266 435338 74822 435894
rect 74266 399338 74822 399894
rect 74266 363338 74822 363894
rect 74266 327338 74822 327894
rect 74266 291338 74822 291894
rect 74266 255338 74822 255894
rect 74266 219338 74822 219894
rect 74266 183338 74822 183894
rect 74266 147338 74822 147894
rect 74266 111338 74822 111894
rect 74266 75338 74822 75894
rect 74266 39338 74822 39894
rect 74266 3338 74822 3894
rect 74266 -1862 74822 -1306
rect 75506 706202 76062 706758
rect 75506 688578 76062 689134
rect 75506 652578 76062 653134
rect 75506 616578 76062 617134
rect 75506 580578 76062 581134
rect 75506 544578 76062 545134
rect 75506 508578 76062 509134
rect 75506 472578 76062 473134
rect 75506 436578 76062 437134
rect 75506 400578 76062 401134
rect 75506 364578 76062 365134
rect 75506 328578 76062 329134
rect 75506 292578 76062 293134
rect 75506 256578 76062 257134
rect 75506 220578 76062 221134
rect 75506 184578 76062 185134
rect 75506 148578 76062 149134
rect 75506 112578 76062 113134
rect 75506 76578 76062 77134
rect 75506 40578 76062 41134
rect 75506 4578 76062 5134
rect 75506 -2822 76062 -2266
rect 76746 707162 77302 707718
rect 76746 689818 77302 690374
rect 76746 653818 77302 654374
rect 76746 617818 77302 618374
rect 76746 581818 77302 582374
rect 76746 545818 77302 546374
rect 76746 509818 77302 510374
rect 76746 473818 77302 474374
rect 76746 437818 77302 438374
rect 76746 401818 77302 402374
rect 76746 365818 77302 366374
rect 76746 329818 77302 330374
rect 76746 293818 77302 294374
rect 76746 257818 77302 258374
rect 76746 221818 77302 222374
rect 76746 185818 77302 186374
rect 76746 149818 77302 150374
rect 76746 113818 77302 114374
rect 76746 77818 77302 78374
rect 76746 41818 77302 42374
rect 76746 5818 77302 6374
rect 76746 -3782 77302 -3226
rect 77986 708122 78542 708678
rect 77986 691058 78542 691614
rect 77986 655058 78542 655614
rect 77986 619058 78542 619614
rect 77986 583058 78542 583614
rect 77986 547058 78542 547614
rect 77986 511058 78542 511614
rect 77986 475058 78542 475614
rect 77986 439058 78542 439614
rect 77986 403058 78542 403614
rect 77986 367058 78542 367614
rect 77986 331058 78542 331614
rect 77986 295058 78542 295614
rect 77986 259058 78542 259614
rect 77986 223058 78542 223614
rect 77986 187058 78542 187614
rect 77986 151058 78542 151614
rect 77986 115058 78542 115614
rect 77986 79058 78542 79614
rect 77986 43058 78542 43614
rect 77986 7058 78542 7614
rect 77986 -4742 78542 -4186
rect 79226 709082 79782 709638
rect 79226 692298 79782 692854
rect 79226 656298 79782 656854
rect 79226 620298 79782 620854
rect 79226 584298 79782 584854
rect 79226 548298 79782 548854
rect 79226 512298 79782 512854
rect 79226 476298 79782 476854
rect 79226 440298 79782 440854
rect 79226 404298 79782 404854
rect 79226 368298 79782 368854
rect 79226 332298 79782 332854
rect 79226 296298 79782 296854
rect 79226 260298 79782 260854
rect 79226 224298 79782 224854
rect 79226 188298 79782 188854
rect 79226 152298 79782 152854
rect 79226 116298 79782 116854
rect 79226 80298 79782 80854
rect 79226 44298 79782 44854
rect 79226 8298 79782 8854
rect 79226 -5702 79782 -5146
rect 80466 710042 81022 710598
rect 80466 693538 81022 694094
rect 80466 657538 81022 658094
rect 80466 621538 81022 622094
rect 80466 585538 81022 586094
rect 80466 549538 81022 550094
rect 80466 513538 81022 514094
rect 80466 477538 81022 478094
rect 80466 441538 81022 442094
rect 80466 405538 81022 406094
rect 80466 369538 81022 370094
rect 80466 333538 81022 334094
rect 80466 297538 81022 298094
rect 80466 261538 81022 262094
rect 80466 225538 81022 226094
rect 80466 189538 81022 190094
rect 80466 153538 81022 154094
rect 80466 117538 81022 118094
rect 80466 81538 81022 82094
rect 80466 45538 81022 46094
rect 80466 9538 81022 10094
rect 80466 -6662 81022 -6106
rect 81706 711002 82262 711558
rect 81706 694778 82262 695334
rect 81706 658778 82262 659334
rect 81706 622778 82262 623334
rect 81706 586778 82262 587334
rect 81706 550778 82262 551334
rect 81706 514778 82262 515334
rect 81706 478778 82262 479334
rect 81706 442778 82262 443334
rect 81706 406778 82262 407334
rect 81706 370778 82262 371334
rect 81706 334778 82262 335334
rect 81706 298778 82262 299334
rect 81706 262778 82262 263334
rect 81706 226778 82262 227334
rect 81706 190778 82262 191334
rect 81706 154778 82262 155334
rect 81706 118778 82262 119334
rect 81706 82778 82262 83334
rect 81706 46778 82262 47334
rect 81706 10778 82262 11334
rect 81706 -7622 82262 -7066
rect 109026 704282 109582 704838
rect 109026 686098 109582 686654
rect 109026 650098 109582 650654
rect 109026 614098 109582 614654
rect 109026 578098 109582 578654
rect 109026 542098 109582 542654
rect 109026 506098 109582 506654
rect 109026 470098 109582 470654
rect 109026 434098 109582 434654
rect 109026 398098 109582 398654
rect 109026 362098 109582 362654
rect 109026 326098 109582 326654
rect 109026 290098 109582 290654
rect 109026 254098 109582 254654
rect 109026 218098 109582 218654
rect 109026 182098 109582 182654
rect 109026 146098 109582 146654
rect 109026 110098 109582 110654
rect 109026 74098 109582 74654
rect 109026 38098 109582 38654
rect 109026 2098 109582 2654
rect 109026 -902 109582 -346
rect 110266 705242 110822 705798
rect 110266 687338 110822 687894
rect 110266 651338 110822 651894
rect 110266 615338 110822 615894
rect 110266 579338 110822 579894
rect 110266 543338 110822 543894
rect 110266 507338 110822 507894
rect 110266 471338 110822 471894
rect 110266 435338 110822 435894
rect 110266 399338 110822 399894
rect 110266 363338 110822 363894
rect 110266 327338 110822 327894
rect 110266 291338 110822 291894
rect 110266 255338 110822 255894
rect 110266 219338 110822 219894
rect 110266 183338 110822 183894
rect 110266 147338 110822 147894
rect 110266 111338 110822 111894
rect 110266 75338 110822 75894
rect 110266 39338 110822 39894
rect 110266 3338 110822 3894
rect 110266 -1862 110822 -1306
rect 111506 706202 112062 706758
rect 111506 688578 112062 689134
rect 111506 652578 112062 653134
rect 111506 616578 112062 617134
rect 111506 580578 112062 581134
rect 111506 544578 112062 545134
rect 111506 508578 112062 509134
rect 111506 472578 112062 473134
rect 111506 436578 112062 437134
rect 111506 400578 112062 401134
rect 111506 364578 112062 365134
rect 111506 328578 112062 329134
rect 111506 292578 112062 293134
rect 111506 256578 112062 257134
rect 111506 220578 112062 221134
rect 111506 184578 112062 185134
rect 111506 148578 112062 149134
rect 111506 112578 112062 113134
rect 111506 76578 112062 77134
rect 111506 40578 112062 41134
rect 111506 4578 112062 5134
rect 111506 -2822 112062 -2266
rect 112746 707162 113302 707718
rect 112746 689818 113302 690374
rect 112746 653818 113302 654374
rect 112746 617818 113302 618374
rect 112746 581818 113302 582374
rect 112746 545818 113302 546374
rect 112746 509818 113302 510374
rect 112746 473818 113302 474374
rect 112746 437818 113302 438374
rect 112746 401818 113302 402374
rect 112746 365818 113302 366374
rect 112746 329818 113302 330374
rect 112746 293818 113302 294374
rect 112746 257818 113302 258374
rect 112746 221818 113302 222374
rect 112746 185818 113302 186374
rect 112746 149818 113302 150374
rect 112746 113818 113302 114374
rect 112746 77818 113302 78374
rect 112746 41818 113302 42374
rect 112746 5818 113302 6374
rect 112746 -3782 113302 -3226
rect 113986 708122 114542 708678
rect 113986 691058 114542 691614
rect 113986 655058 114542 655614
rect 113986 619058 114542 619614
rect 113986 583058 114542 583614
rect 113986 547058 114542 547614
rect 113986 511058 114542 511614
rect 113986 475058 114542 475614
rect 113986 439058 114542 439614
rect 113986 403058 114542 403614
rect 113986 367058 114542 367614
rect 113986 331058 114542 331614
rect 113986 295058 114542 295614
rect 113986 259058 114542 259614
rect 113986 223058 114542 223614
rect 113986 187058 114542 187614
rect 113986 151058 114542 151614
rect 113986 115058 114542 115614
rect 113986 79058 114542 79614
rect 113986 43058 114542 43614
rect 113986 7058 114542 7614
rect 113986 -4742 114542 -4186
rect 115226 709082 115782 709638
rect 115226 692298 115782 692854
rect 115226 656298 115782 656854
rect 115226 620298 115782 620854
rect 115226 584298 115782 584854
rect 115226 548298 115782 548854
rect 115226 512298 115782 512854
rect 115226 476298 115782 476854
rect 115226 440298 115782 440854
rect 115226 404298 115782 404854
rect 115226 368298 115782 368854
rect 115226 332298 115782 332854
rect 115226 296298 115782 296854
rect 115226 260298 115782 260854
rect 115226 224298 115782 224854
rect 115226 188298 115782 188854
rect 115226 152298 115782 152854
rect 115226 116298 115782 116854
rect 115226 80298 115782 80854
rect 115226 44298 115782 44854
rect 115226 8298 115782 8854
rect 115226 -5702 115782 -5146
rect 116466 710042 117022 710598
rect 116466 693538 117022 694094
rect 116466 657538 117022 658094
rect 116466 621538 117022 622094
rect 116466 585538 117022 586094
rect 116466 549538 117022 550094
rect 116466 513538 117022 514094
rect 116466 477538 117022 478094
rect 116466 441538 117022 442094
rect 116466 405538 117022 406094
rect 116466 369538 117022 370094
rect 116466 333538 117022 334094
rect 116466 297538 117022 298094
rect 116466 261538 117022 262094
rect 116466 225538 117022 226094
rect 116466 189538 117022 190094
rect 116466 153538 117022 154094
rect 116466 117538 117022 118094
rect 116466 81538 117022 82094
rect 116466 45538 117022 46094
rect 116466 9538 117022 10094
rect 116466 -6662 117022 -6106
rect 117706 711002 118262 711558
rect 117706 694778 118262 695334
rect 117706 658778 118262 659334
rect 117706 622778 118262 623334
rect 117706 586778 118262 587334
rect 117706 550778 118262 551334
rect 117706 514778 118262 515334
rect 117706 478778 118262 479334
rect 117706 442778 118262 443334
rect 117706 406778 118262 407334
rect 117706 370778 118262 371334
rect 117706 334778 118262 335334
rect 117706 298778 118262 299334
rect 117706 262778 118262 263334
rect 117706 226778 118262 227334
rect 117706 190778 118262 191334
rect 117706 154778 118262 155334
rect 117706 118778 118262 119334
rect 117706 82778 118262 83334
rect 117706 46778 118262 47334
rect 117706 10778 118262 11334
rect 117706 -7622 118262 -7066
rect 145026 704282 145582 704838
rect 145026 686098 145582 686654
rect 145026 650098 145582 650654
rect 145026 614098 145582 614654
rect 145026 578098 145582 578654
rect 145026 542098 145582 542654
rect 145026 506098 145582 506654
rect 145026 470098 145582 470654
rect 145026 434098 145582 434654
rect 145026 398098 145582 398654
rect 145026 362098 145582 362654
rect 145026 326098 145582 326654
rect 145026 290098 145582 290654
rect 145026 254098 145582 254654
rect 145026 218098 145582 218654
rect 145026 182098 145582 182654
rect 145026 146098 145582 146654
rect 145026 110098 145582 110654
rect 145026 74098 145582 74654
rect 145026 38098 145582 38654
rect 145026 2098 145582 2654
rect 145026 -902 145582 -346
rect 146266 705242 146822 705798
rect 146266 687338 146822 687894
rect 146266 651338 146822 651894
rect 146266 615338 146822 615894
rect 146266 579338 146822 579894
rect 146266 543338 146822 543894
rect 146266 507338 146822 507894
rect 146266 471338 146822 471894
rect 146266 435338 146822 435894
rect 146266 399338 146822 399894
rect 146266 363338 146822 363894
rect 146266 327338 146822 327894
rect 146266 291338 146822 291894
rect 146266 255338 146822 255894
rect 146266 219338 146822 219894
rect 146266 183338 146822 183894
rect 146266 147338 146822 147894
rect 146266 111338 146822 111894
rect 146266 75338 146822 75894
rect 146266 39338 146822 39894
rect 146266 3338 146822 3894
rect 146266 -1862 146822 -1306
rect 147506 706202 148062 706758
rect 147506 688578 148062 689134
rect 147506 652578 148062 653134
rect 147506 616578 148062 617134
rect 147506 580578 148062 581134
rect 147506 544578 148062 545134
rect 147506 508578 148062 509134
rect 147506 472578 148062 473134
rect 147506 436578 148062 437134
rect 147506 400578 148062 401134
rect 147506 364578 148062 365134
rect 147506 328578 148062 329134
rect 147506 292578 148062 293134
rect 147506 256578 148062 257134
rect 147506 220578 148062 221134
rect 147506 184578 148062 185134
rect 147506 148578 148062 149134
rect 147506 112578 148062 113134
rect 147506 76578 148062 77134
rect 147506 40578 148062 41134
rect 147506 4578 148062 5134
rect 147506 -2822 148062 -2266
rect 148746 707162 149302 707718
rect 148746 689818 149302 690374
rect 148746 653818 149302 654374
rect 148746 617818 149302 618374
rect 148746 581818 149302 582374
rect 148746 545818 149302 546374
rect 148746 509818 149302 510374
rect 148746 473818 149302 474374
rect 148746 437818 149302 438374
rect 148746 401818 149302 402374
rect 148746 365818 149302 366374
rect 148746 329818 149302 330374
rect 148746 293818 149302 294374
rect 148746 257818 149302 258374
rect 148746 221818 149302 222374
rect 148746 185818 149302 186374
rect 148746 149818 149302 150374
rect 148746 113818 149302 114374
rect 148746 77818 149302 78374
rect 148746 41818 149302 42374
rect 148746 5818 149302 6374
rect 148746 -3782 149302 -3226
rect 149986 708122 150542 708678
rect 149986 691058 150542 691614
rect 149986 655058 150542 655614
rect 149986 619058 150542 619614
rect 149986 583058 150542 583614
rect 149986 547058 150542 547614
rect 149986 511058 150542 511614
rect 149986 475058 150542 475614
rect 149986 439058 150542 439614
rect 149986 403058 150542 403614
rect 149986 367058 150542 367614
rect 149986 331058 150542 331614
rect 149986 295058 150542 295614
rect 149986 259058 150542 259614
rect 149986 223058 150542 223614
rect 149986 187058 150542 187614
rect 149986 151058 150542 151614
rect 149986 115058 150542 115614
rect 149986 79058 150542 79614
rect 149986 43058 150542 43614
rect 149986 7058 150542 7614
rect 149986 -4742 150542 -4186
rect 151226 709082 151782 709638
rect 151226 692298 151782 692854
rect 151226 656298 151782 656854
rect 151226 620298 151782 620854
rect 151226 584298 151782 584854
rect 151226 548298 151782 548854
rect 151226 512298 151782 512854
rect 151226 476298 151782 476854
rect 151226 440298 151782 440854
rect 151226 404298 151782 404854
rect 151226 368298 151782 368854
rect 151226 332298 151782 332854
rect 151226 296298 151782 296854
rect 151226 260298 151782 260854
rect 151226 224298 151782 224854
rect 151226 188298 151782 188854
rect 151226 152298 151782 152854
rect 151226 116298 151782 116854
rect 151226 80298 151782 80854
rect 151226 44298 151782 44854
rect 151226 8298 151782 8854
rect 151226 -5702 151782 -5146
rect 152466 710042 153022 710598
rect 152466 693538 153022 694094
rect 152466 657538 153022 658094
rect 152466 621538 153022 622094
rect 152466 585538 153022 586094
rect 152466 549538 153022 550094
rect 152466 513538 153022 514094
rect 152466 477538 153022 478094
rect 152466 441538 153022 442094
rect 152466 405538 153022 406094
rect 152466 369538 153022 370094
rect 152466 333538 153022 334094
rect 152466 297538 153022 298094
rect 152466 261538 153022 262094
rect 152466 225538 153022 226094
rect 152466 189538 153022 190094
rect 152466 153538 153022 154094
rect 152466 117538 153022 118094
rect 152466 81538 153022 82094
rect 152466 45538 153022 46094
rect 152466 9538 153022 10094
rect 152466 -6662 153022 -6106
rect 153706 711002 154262 711558
rect 153706 694778 154262 695334
rect 153706 658778 154262 659334
rect 153706 622778 154262 623334
rect 153706 586778 154262 587334
rect 153706 550778 154262 551334
rect 153706 514778 154262 515334
rect 153706 478778 154262 479334
rect 153706 442778 154262 443334
rect 153706 406778 154262 407334
rect 153706 370778 154262 371334
rect 153706 334778 154262 335334
rect 153706 298778 154262 299334
rect 153706 262778 154262 263334
rect 153706 226778 154262 227334
rect 153706 190778 154262 191334
rect 153706 154778 154262 155334
rect 153706 118778 154262 119334
rect 153706 82778 154262 83334
rect 153706 46778 154262 47334
rect 153706 10778 154262 11334
rect 153706 -7622 154262 -7066
rect 181026 704282 181582 704838
rect 181026 686098 181582 686654
rect 181026 650098 181582 650654
rect 181026 614098 181582 614654
rect 181026 578098 181582 578654
rect 181026 542098 181582 542654
rect 181026 506098 181582 506654
rect 181026 470098 181582 470654
rect 181026 434098 181582 434654
rect 181026 398098 181582 398654
rect 181026 362098 181582 362654
rect 181026 326098 181582 326654
rect 181026 290098 181582 290654
rect 181026 254098 181582 254654
rect 181026 218098 181582 218654
rect 181026 182098 181582 182654
rect 181026 146098 181582 146654
rect 181026 110098 181582 110654
rect 181026 74098 181582 74654
rect 181026 38098 181582 38654
rect 181026 2098 181582 2654
rect 181026 -902 181582 -346
rect 182266 705242 182822 705798
rect 182266 687338 182822 687894
rect 182266 651338 182822 651894
rect 182266 615338 182822 615894
rect 182266 579338 182822 579894
rect 182266 543338 182822 543894
rect 182266 507338 182822 507894
rect 182266 471338 182822 471894
rect 182266 435338 182822 435894
rect 182266 399338 182822 399894
rect 182266 363338 182822 363894
rect 182266 327338 182822 327894
rect 182266 291338 182822 291894
rect 182266 255338 182822 255894
rect 182266 219338 182822 219894
rect 182266 183338 182822 183894
rect 182266 147338 182822 147894
rect 182266 111338 182822 111894
rect 182266 75338 182822 75894
rect 182266 39338 182822 39894
rect 182266 3338 182822 3894
rect 182266 -1862 182822 -1306
rect 183506 706202 184062 706758
rect 183506 688578 184062 689134
rect 183506 652578 184062 653134
rect 183506 616578 184062 617134
rect 183506 580578 184062 581134
rect 183506 544578 184062 545134
rect 183506 508578 184062 509134
rect 183506 472578 184062 473134
rect 183506 436578 184062 437134
rect 183506 400578 184062 401134
rect 183506 364578 184062 365134
rect 183506 328578 184062 329134
rect 183506 292578 184062 293134
rect 183506 256578 184062 257134
rect 183506 220578 184062 221134
rect 183506 184578 184062 185134
rect 183506 148578 184062 149134
rect 183506 112578 184062 113134
rect 183506 76578 184062 77134
rect 183506 40578 184062 41134
rect 183506 4578 184062 5134
rect 183506 -2822 184062 -2266
rect 184746 707162 185302 707718
rect 184746 689818 185302 690374
rect 184746 653818 185302 654374
rect 184746 617818 185302 618374
rect 184746 581818 185302 582374
rect 184746 545818 185302 546374
rect 184746 509818 185302 510374
rect 184746 473818 185302 474374
rect 184746 437818 185302 438374
rect 184746 401818 185302 402374
rect 184746 365818 185302 366374
rect 184746 329818 185302 330374
rect 184746 293818 185302 294374
rect 184746 257818 185302 258374
rect 184746 221818 185302 222374
rect 184746 185818 185302 186374
rect 184746 149818 185302 150374
rect 184746 113818 185302 114374
rect 184746 77818 185302 78374
rect 184746 41818 185302 42374
rect 184746 5818 185302 6374
rect 184746 -3782 185302 -3226
rect 185986 708122 186542 708678
rect 185986 691058 186542 691614
rect 185986 655058 186542 655614
rect 185986 619058 186542 619614
rect 185986 583058 186542 583614
rect 185986 547058 186542 547614
rect 185986 511058 186542 511614
rect 185986 475058 186542 475614
rect 185986 439058 186542 439614
rect 185986 403058 186542 403614
rect 185986 367058 186542 367614
rect 185986 331058 186542 331614
rect 185986 295058 186542 295614
rect 185986 259058 186542 259614
rect 185986 223058 186542 223614
rect 185986 187058 186542 187614
rect 185986 151058 186542 151614
rect 185986 115058 186542 115614
rect 185986 79058 186542 79614
rect 185986 43058 186542 43614
rect 185986 7058 186542 7614
rect 185986 -4742 186542 -4186
rect 187226 709082 187782 709638
rect 187226 692298 187782 692854
rect 187226 656298 187782 656854
rect 187226 620298 187782 620854
rect 187226 584298 187782 584854
rect 187226 548298 187782 548854
rect 187226 512298 187782 512854
rect 187226 476298 187782 476854
rect 187226 440298 187782 440854
rect 187226 404298 187782 404854
rect 187226 368298 187782 368854
rect 187226 332298 187782 332854
rect 187226 296298 187782 296854
rect 187226 260298 187782 260854
rect 187226 224298 187782 224854
rect 187226 188298 187782 188854
rect 187226 152298 187782 152854
rect 187226 116298 187782 116854
rect 187226 80298 187782 80854
rect 187226 44298 187782 44854
rect 187226 8298 187782 8854
rect 187226 -5702 187782 -5146
rect 188466 710042 189022 710598
rect 188466 693538 189022 694094
rect 188466 657538 189022 658094
rect 188466 621538 189022 622094
rect 188466 585538 189022 586094
rect 188466 549538 189022 550094
rect 188466 513538 189022 514094
rect 188466 477538 189022 478094
rect 188466 441538 189022 442094
rect 188466 405538 189022 406094
rect 188466 369538 189022 370094
rect 188466 333538 189022 334094
rect 188466 297538 189022 298094
rect 188466 261538 189022 262094
rect 188466 225538 189022 226094
rect 188466 189538 189022 190094
rect 188466 153538 189022 154094
rect 188466 117538 189022 118094
rect 188466 81538 189022 82094
rect 188466 45538 189022 46094
rect 188466 9538 189022 10094
rect 188466 -6662 189022 -6106
rect 189706 711002 190262 711558
rect 189706 694778 190262 695334
rect 189706 658778 190262 659334
rect 189706 622778 190262 623334
rect 189706 586778 190262 587334
rect 189706 550778 190262 551334
rect 189706 514778 190262 515334
rect 189706 478778 190262 479334
rect 189706 442778 190262 443334
rect 189706 406778 190262 407334
rect 189706 370778 190262 371334
rect 189706 334778 190262 335334
rect 189706 298778 190262 299334
rect 189706 262778 190262 263334
rect 189706 226778 190262 227334
rect 189706 190778 190262 191334
rect 189706 154778 190262 155334
rect 189706 118778 190262 119334
rect 189706 82778 190262 83334
rect 189706 46778 190262 47334
rect 189706 10778 190262 11334
rect 189706 -7622 190262 -7066
rect 217026 704282 217582 704838
rect 217026 686098 217582 686654
rect 217026 650098 217582 650654
rect 217026 614098 217582 614654
rect 217026 578098 217582 578654
rect 217026 542098 217582 542654
rect 217026 506098 217582 506654
rect 217026 470098 217582 470654
rect 217026 434098 217582 434654
rect 217026 398098 217582 398654
rect 217026 362098 217582 362654
rect 217026 326098 217582 326654
rect 217026 290098 217582 290654
rect 217026 254098 217582 254654
rect 217026 218098 217582 218654
rect 217026 182098 217582 182654
rect 217026 146098 217582 146654
rect 217026 110098 217582 110654
rect 217026 74098 217582 74654
rect 217026 38098 217582 38654
rect 217026 2098 217582 2654
rect 217026 -902 217582 -346
rect 218266 705242 218822 705798
rect 218266 687338 218822 687894
rect 218266 651338 218822 651894
rect 218266 615338 218822 615894
rect 218266 579338 218822 579894
rect 218266 543338 218822 543894
rect 218266 507338 218822 507894
rect 218266 471338 218822 471894
rect 218266 435338 218822 435894
rect 218266 399338 218822 399894
rect 218266 363338 218822 363894
rect 218266 327338 218822 327894
rect 218266 291338 218822 291894
rect 218266 255338 218822 255894
rect 218266 219338 218822 219894
rect 218266 183338 218822 183894
rect 218266 147338 218822 147894
rect 218266 111338 218822 111894
rect 218266 75338 218822 75894
rect 218266 39338 218822 39894
rect 218266 3338 218822 3894
rect 218266 -1862 218822 -1306
rect 219506 706202 220062 706758
rect 219506 688578 220062 689134
rect 219506 652578 220062 653134
rect 219506 616578 220062 617134
rect 219506 580578 220062 581134
rect 219506 544578 220062 545134
rect 219506 508578 220062 509134
rect 219506 472578 220062 473134
rect 219506 436578 220062 437134
rect 219506 400578 220062 401134
rect 219506 364578 220062 365134
rect 219506 328578 220062 329134
rect 219506 292578 220062 293134
rect 219506 256578 220062 257134
rect 219506 220578 220062 221134
rect 219506 184578 220062 185134
rect 219506 148578 220062 149134
rect 219506 112578 220062 113134
rect 219506 76578 220062 77134
rect 219506 40578 220062 41134
rect 219506 4578 220062 5134
rect 219506 -2822 220062 -2266
rect 220746 707162 221302 707718
rect 220746 689818 221302 690374
rect 220746 653818 221302 654374
rect 220746 617818 221302 618374
rect 220746 581818 221302 582374
rect 220746 545818 221302 546374
rect 220746 509818 221302 510374
rect 220746 473818 221302 474374
rect 220746 437818 221302 438374
rect 220746 401818 221302 402374
rect 220746 365818 221302 366374
rect 220746 329818 221302 330374
rect 220746 293818 221302 294374
rect 220746 257818 221302 258374
rect 220746 221818 221302 222374
rect 220746 185818 221302 186374
rect 220746 149818 221302 150374
rect 220746 113818 221302 114374
rect 220746 77818 221302 78374
rect 220746 41818 221302 42374
rect 220746 5818 221302 6374
rect 220746 -3782 221302 -3226
rect 221986 708122 222542 708678
rect 221986 691058 222542 691614
rect 221986 655058 222542 655614
rect 221986 619058 222542 619614
rect 221986 583058 222542 583614
rect 221986 547058 222542 547614
rect 221986 511058 222542 511614
rect 221986 475058 222542 475614
rect 221986 439058 222542 439614
rect 221986 403058 222542 403614
rect 221986 367058 222542 367614
rect 221986 331058 222542 331614
rect 221986 295058 222542 295614
rect 221986 259058 222542 259614
rect 221986 223058 222542 223614
rect 221986 187058 222542 187614
rect 221986 151058 222542 151614
rect 221986 115058 222542 115614
rect 221986 79058 222542 79614
rect 221986 43058 222542 43614
rect 221986 7058 222542 7614
rect 221986 -4742 222542 -4186
rect 223226 709082 223782 709638
rect 223226 692298 223782 692854
rect 223226 656298 223782 656854
rect 223226 620298 223782 620854
rect 223226 584298 223782 584854
rect 223226 548298 223782 548854
rect 223226 512298 223782 512854
rect 223226 476298 223782 476854
rect 223226 440298 223782 440854
rect 223226 404298 223782 404854
rect 223226 368298 223782 368854
rect 223226 332298 223782 332854
rect 223226 296298 223782 296854
rect 223226 260298 223782 260854
rect 223226 224298 223782 224854
rect 223226 188298 223782 188854
rect 223226 152298 223782 152854
rect 223226 116298 223782 116854
rect 223226 80298 223782 80854
rect 223226 44298 223782 44854
rect 223226 8298 223782 8854
rect 223226 -5702 223782 -5146
rect 224466 710042 225022 710598
rect 224466 693538 225022 694094
rect 224466 657538 225022 658094
rect 224466 621538 225022 622094
rect 224466 585538 225022 586094
rect 224466 549538 225022 550094
rect 224466 513538 225022 514094
rect 224466 477538 225022 478094
rect 224466 441538 225022 442094
rect 224466 405538 225022 406094
rect 224466 369538 225022 370094
rect 224466 333538 225022 334094
rect 224466 297538 225022 298094
rect 224466 261538 225022 262094
rect 224466 225538 225022 226094
rect 224466 189538 225022 190094
rect 224466 153538 225022 154094
rect 224466 117538 225022 118094
rect 224466 81538 225022 82094
rect 224466 45538 225022 46094
rect 224466 9538 225022 10094
rect 224466 -6662 225022 -6106
rect 225706 711002 226262 711558
rect 225706 694778 226262 695334
rect 225706 658778 226262 659334
rect 225706 622778 226262 623334
rect 225706 586778 226262 587334
rect 225706 550778 226262 551334
rect 225706 514778 226262 515334
rect 225706 478778 226262 479334
rect 225706 442778 226262 443334
rect 225706 406778 226262 407334
rect 225706 370778 226262 371334
rect 225706 334778 226262 335334
rect 225706 298778 226262 299334
rect 225706 262778 226262 263334
rect 225706 226778 226262 227334
rect 225706 190778 226262 191334
rect 225706 154778 226262 155334
rect 225706 118778 226262 119334
rect 225706 82778 226262 83334
rect 225706 46778 226262 47334
rect 225706 10778 226262 11334
rect 225706 -7622 226262 -7066
rect 253026 704282 253582 704838
rect 253026 686098 253582 686654
rect 253026 650098 253582 650654
rect 253026 614098 253582 614654
rect 253026 578098 253582 578654
rect 253026 542098 253582 542654
rect 253026 506098 253582 506654
rect 253026 470098 253582 470654
rect 253026 434098 253582 434654
rect 253026 398098 253582 398654
rect 253026 362098 253582 362654
rect 253026 326098 253582 326654
rect 253026 290098 253582 290654
rect 253026 254098 253582 254654
rect 253026 218098 253582 218654
rect 253026 182098 253582 182654
rect 253026 146098 253582 146654
rect 253026 110098 253582 110654
rect 253026 74098 253582 74654
rect 253026 38098 253582 38654
rect 253026 2098 253582 2654
rect 253026 -902 253582 -346
rect 254266 705242 254822 705798
rect 254266 687338 254822 687894
rect 254266 651338 254822 651894
rect 254266 615338 254822 615894
rect 254266 579338 254822 579894
rect 254266 543338 254822 543894
rect 254266 507338 254822 507894
rect 254266 471338 254822 471894
rect 254266 435338 254822 435894
rect 254266 399338 254822 399894
rect 254266 363338 254822 363894
rect 254266 327338 254822 327894
rect 254266 291338 254822 291894
rect 254266 255338 254822 255894
rect 254266 219338 254822 219894
rect 254266 183338 254822 183894
rect 254266 147338 254822 147894
rect 254266 111338 254822 111894
rect 254266 75338 254822 75894
rect 254266 39338 254822 39894
rect 254266 3338 254822 3894
rect 254266 -1862 254822 -1306
rect 255506 706202 256062 706758
rect 255506 688578 256062 689134
rect 255506 652578 256062 653134
rect 255506 616578 256062 617134
rect 255506 580578 256062 581134
rect 255506 544578 256062 545134
rect 255506 508578 256062 509134
rect 255506 472578 256062 473134
rect 255506 436578 256062 437134
rect 255506 400578 256062 401134
rect 255506 364578 256062 365134
rect 255506 328578 256062 329134
rect 255506 292578 256062 293134
rect 255506 256578 256062 257134
rect 255506 220578 256062 221134
rect 255506 184578 256062 185134
rect 255506 148578 256062 149134
rect 255506 112578 256062 113134
rect 255506 76578 256062 77134
rect 255506 40578 256062 41134
rect 255506 4578 256062 5134
rect 255506 -2822 256062 -2266
rect 256746 707162 257302 707718
rect 256746 689818 257302 690374
rect 256746 653818 257302 654374
rect 256746 617818 257302 618374
rect 256746 581818 257302 582374
rect 256746 545818 257302 546374
rect 256746 509818 257302 510374
rect 256746 473818 257302 474374
rect 256746 437818 257302 438374
rect 256746 401818 257302 402374
rect 256746 365818 257302 366374
rect 256746 329818 257302 330374
rect 256746 293818 257302 294374
rect 256746 257818 257302 258374
rect 256746 221818 257302 222374
rect 256746 185818 257302 186374
rect 256746 149818 257302 150374
rect 256746 113818 257302 114374
rect 256746 77818 257302 78374
rect 256746 41818 257302 42374
rect 256746 5818 257302 6374
rect 256746 -3782 257302 -3226
rect 257986 708122 258542 708678
rect 257986 691058 258542 691614
rect 257986 655058 258542 655614
rect 257986 619058 258542 619614
rect 257986 583058 258542 583614
rect 257986 547058 258542 547614
rect 257986 511058 258542 511614
rect 257986 475058 258542 475614
rect 257986 439058 258542 439614
rect 257986 403058 258542 403614
rect 257986 367058 258542 367614
rect 257986 331058 258542 331614
rect 257986 295058 258542 295614
rect 257986 259058 258542 259614
rect 257986 223058 258542 223614
rect 257986 187058 258542 187614
rect 257986 151058 258542 151614
rect 257986 115058 258542 115614
rect 257986 79058 258542 79614
rect 257986 43058 258542 43614
rect 257986 7058 258542 7614
rect 257986 -4742 258542 -4186
rect 259226 709082 259782 709638
rect 259226 692298 259782 692854
rect 259226 656298 259782 656854
rect 259226 620298 259782 620854
rect 259226 584298 259782 584854
rect 259226 548298 259782 548854
rect 259226 512298 259782 512854
rect 259226 476298 259782 476854
rect 259226 440298 259782 440854
rect 259226 404298 259782 404854
rect 259226 368298 259782 368854
rect 259226 332298 259782 332854
rect 259226 296298 259782 296854
rect 259226 260298 259782 260854
rect 259226 224298 259782 224854
rect 259226 188298 259782 188854
rect 259226 152298 259782 152854
rect 259226 116298 259782 116854
rect 259226 80298 259782 80854
rect 259226 44298 259782 44854
rect 259226 8298 259782 8854
rect 259226 -5702 259782 -5146
rect 260466 710042 261022 710598
rect 260466 693538 261022 694094
rect 260466 657538 261022 658094
rect 260466 621538 261022 622094
rect 260466 585538 261022 586094
rect 260466 549538 261022 550094
rect 260466 513538 261022 514094
rect 260466 477538 261022 478094
rect 260466 441538 261022 442094
rect 260466 405538 261022 406094
rect 260466 369538 261022 370094
rect 260466 333538 261022 334094
rect 260466 297538 261022 298094
rect 260466 261538 261022 262094
rect 260466 225538 261022 226094
rect 260466 189538 261022 190094
rect 260466 153538 261022 154094
rect 260466 117538 261022 118094
rect 260466 81538 261022 82094
rect 260466 45538 261022 46094
rect 260466 9538 261022 10094
rect 260466 -6662 261022 -6106
rect 261706 711002 262262 711558
rect 261706 694778 262262 695334
rect 261706 658778 262262 659334
rect 261706 622778 262262 623334
rect 261706 586778 262262 587334
rect 261706 550778 262262 551334
rect 261706 514778 262262 515334
rect 261706 478778 262262 479334
rect 261706 442778 262262 443334
rect 261706 406778 262262 407334
rect 261706 370778 262262 371334
rect 261706 334778 262262 335334
rect 261706 298778 262262 299334
rect 261706 262778 262262 263334
rect 261706 226778 262262 227334
rect 261706 190778 262262 191334
rect 261706 154778 262262 155334
rect 261706 118778 262262 119334
rect 261706 82778 262262 83334
rect 261706 46778 262262 47334
rect 261706 10778 262262 11334
rect 261706 -7622 262262 -7066
rect 289026 704282 289582 704838
rect 289026 686098 289582 686654
rect 289026 650098 289582 650654
rect 289026 614098 289582 614654
rect 289026 578098 289582 578654
rect 289026 542098 289582 542654
rect 289026 506098 289582 506654
rect 289026 470098 289582 470654
rect 289026 434098 289582 434654
rect 289026 398098 289582 398654
rect 289026 362098 289582 362654
rect 289026 326098 289582 326654
rect 289026 290098 289582 290654
rect 289026 254098 289582 254654
rect 289026 218098 289582 218654
rect 289026 182098 289582 182654
rect 289026 146098 289582 146654
rect 289026 110098 289582 110654
rect 289026 74098 289582 74654
rect 289026 38098 289582 38654
rect 289026 2098 289582 2654
rect 289026 -902 289582 -346
rect 290266 705242 290822 705798
rect 290266 687338 290822 687894
rect 290266 651338 290822 651894
rect 290266 615338 290822 615894
rect 290266 579338 290822 579894
rect 290266 543338 290822 543894
rect 290266 507338 290822 507894
rect 290266 471338 290822 471894
rect 290266 435338 290822 435894
rect 290266 399338 290822 399894
rect 290266 363338 290822 363894
rect 290266 327338 290822 327894
rect 290266 291338 290822 291894
rect 290266 255338 290822 255894
rect 290266 219338 290822 219894
rect 290266 183338 290822 183894
rect 290266 147338 290822 147894
rect 290266 111338 290822 111894
rect 290266 75338 290822 75894
rect 290266 39338 290822 39894
rect 290266 3338 290822 3894
rect 290266 -1862 290822 -1306
rect 291506 706202 292062 706758
rect 291506 688578 292062 689134
rect 291506 652578 292062 653134
rect 291506 616578 292062 617134
rect 291506 580578 292062 581134
rect 291506 544578 292062 545134
rect 291506 508578 292062 509134
rect 291506 472578 292062 473134
rect 291506 436578 292062 437134
rect 291506 400578 292062 401134
rect 291506 364578 292062 365134
rect 291506 328578 292062 329134
rect 291506 292578 292062 293134
rect 291506 256578 292062 257134
rect 291506 220578 292062 221134
rect 291506 184578 292062 185134
rect 291506 148578 292062 149134
rect 291506 112578 292062 113134
rect 291506 76578 292062 77134
rect 291506 40578 292062 41134
rect 291506 4578 292062 5134
rect 291506 -2822 292062 -2266
rect 292746 707162 293302 707718
rect 292746 689818 293302 690374
rect 292746 653818 293302 654374
rect 292746 617818 293302 618374
rect 292746 581818 293302 582374
rect 292746 545818 293302 546374
rect 292746 509818 293302 510374
rect 292746 473818 293302 474374
rect 292746 437818 293302 438374
rect 292746 401818 293302 402374
rect 292746 365818 293302 366374
rect 292746 329818 293302 330374
rect 292746 293818 293302 294374
rect 292746 257818 293302 258374
rect 292746 221818 293302 222374
rect 292746 185818 293302 186374
rect 292746 149818 293302 150374
rect 292746 113818 293302 114374
rect 292746 77818 293302 78374
rect 292746 41818 293302 42374
rect 292746 5818 293302 6374
rect 292746 -3782 293302 -3226
rect 293986 708122 294542 708678
rect 293986 691058 294542 691614
rect 293986 655058 294542 655614
rect 293986 619058 294542 619614
rect 293986 583058 294542 583614
rect 293986 547058 294542 547614
rect 293986 511058 294542 511614
rect 293986 475058 294542 475614
rect 293986 439058 294542 439614
rect 293986 403058 294542 403614
rect 293986 367058 294542 367614
rect 293986 331058 294542 331614
rect 293986 295058 294542 295614
rect 293986 259058 294542 259614
rect 293986 223058 294542 223614
rect 293986 187058 294542 187614
rect 293986 151058 294542 151614
rect 293986 115058 294542 115614
rect 293986 79058 294542 79614
rect 293986 43058 294542 43614
rect 293986 7058 294542 7614
rect 293986 -4742 294542 -4186
rect 295226 709082 295782 709638
rect 295226 692298 295782 692854
rect 295226 656298 295782 656854
rect 295226 620298 295782 620854
rect 295226 584298 295782 584854
rect 295226 548298 295782 548854
rect 295226 512298 295782 512854
rect 295226 476298 295782 476854
rect 295226 440298 295782 440854
rect 295226 404298 295782 404854
rect 295226 368298 295782 368854
rect 295226 332298 295782 332854
rect 295226 296298 295782 296854
rect 295226 260298 295782 260854
rect 295226 224298 295782 224854
rect 295226 188298 295782 188854
rect 295226 152298 295782 152854
rect 295226 116298 295782 116854
rect 295226 80298 295782 80854
rect 295226 44298 295782 44854
rect 295226 8298 295782 8854
rect 295226 -5702 295782 -5146
rect 296466 710042 297022 710598
rect 296466 693538 297022 694094
rect 296466 657538 297022 658094
rect 296466 621538 297022 622094
rect 296466 585538 297022 586094
rect 296466 549538 297022 550094
rect 296466 513538 297022 514094
rect 296466 477538 297022 478094
rect 296466 441538 297022 442094
rect 296466 405538 297022 406094
rect 296466 369538 297022 370094
rect 296466 333538 297022 334094
rect 296466 297538 297022 298094
rect 296466 261538 297022 262094
rect 296466 225538 297022 226094
rect 296466 189538 297022 190094
rect 296466 153538 297022 154094
rect 296466 117538 297022 118094
rect 296466 81538 297022 82094
rect 296466 45538 297022 46094
rect 296466 9538 297022 10094
rect 296466 -6662 297022 -6106
rect 297706 711002 298262 711558
rect 297706 694778 298262 695334
rect 297706 658778 298262 659334
rect 297706 622778 298262 623334
rect 297706 586778 298262 587334
rect 297706 550778 298262 551334
rect 297706 514778 298262 515334
rect 297706 478778 298262 479334
rect 297706 442778 298262 443334
rect 297706 406778 298262 407334
rect 297706 370778 298262 371334
rect 297706 334778 298262 335334
rect 297706 298778 298262 299334
rect 297706 262778 298262 263334
rect 297706 226778 298262 227334
rect 297706 190778 298262 191334
rect 297706 154778 298262 155334
rect 297706 118778 298262 119334
rect 297706 82778 298262 83334
rect 297706 46778 298262 47334
rect 297706 10778 298262 11334
rect 297706 -7622 298262 -7066
rect 325026 704282 325582 704838
rect 325026 686098 325582 686654
rect 325026 650098 325582 650654
rect 325026 614098 325582 614654
rect 325026 578098 325582 578654
rect 325026 542098 325582 542654
rect 325026 506098 325582 506654
rect 325026 470098 325582 470654
rect 325026 434098 325582 434654
rect 325026 398098 325582 398654
rect 325026 362098 325582 362654
rect 325026 326098 325582 326654
rect 325026 290098 325582 290654
rect 325026 254098 325582 254654
rect 325026 218098 325582 218654
rect 325026 182098 325582 182654
rect 325026 146098 325582 146654
rect 325026 110098 325582 110654
rect 325026 74098 325582 74654
rect 325026 38098 325582 38654
rect 325026 2098 325582 2654
rect 325026 -902 325582 -346
rect 326266 705242 326822 705798
rect 326266 687338 326822 687894
rect 326266 651338 326822 651894
rect 326266 615338 326822 615894
rect 326266 579338 326822 579894
rect 326266 543338 326822 543894
rect 326266 507338 326822 507894
rect 326266 471338 326822 471894
rect 326266 435338 326822 435894
rect 326266 399338 326822 399894
rect 326266 363338 326822 363894
rect 326266 327338 326822 327894
rect 326266 291338 326822 291894
rect 326266 255338 326822 255894
rect 326266 219338 326822 219894
rect 326266 183338 326822 183894
rect 326266 147338 326822 147894
rect 326266 111338 326822 111894
rect 326266 75338 326822 75894
rect 326266 39338 326822 39894
rect 326266 3338 326822 3894
rect 326266 -1862 326822 -1306
rect 327506 706202 328062 706758
rect 327506 688578 328062 689134
rect 327506 652578 328062 653134
rect 327506 616578 328062 617134
rect 327506 580578 328062 581134
rect 327506 544578 328062 545134
rect 327506 508578 328062 509134
rect 327506 472578 328062 473134
rect 327506 436578 328062 437134
rect 327506 400578 328062 401134
rect 327506 364578 328062 365134
rect 327506 328578 328062 329134
rect 327506 292578 328062 293134
rect 327506 256578 328062 257134
rect 327506 220578 328062 221134
rect 327506 184578 328062 185134
rect 327506 148578 328062 149134
rect 327506 112578 328062 113134
rect 327506 76578 328062 77134
rect 327506 40578 328062 41134
rect 327506 4578 328062 5134
rect 327506 -2822 328062 -2266
rect 328746 707162 329302 707718
rect 328746 689818 329302 690374
rect 328746 653818 329302 654374
rect 328746 617818 329302 618374
rect 328746 581818 329302 582374
rect 328746 545818 329302 546374
rect 328746 509818 329302 510374
rect 328746 473818 329302 474374
rect 328746 437818 329302 438374
rect 328746 401818 329302 402374
rect 328746 365818 329302 366374
rect 328746 329818 329302 330374
rect 328746 293818 329302 294374
rect 328746 257818 329302 258374
rect 328746 221818 329302 222374
rect 328746 185818 329302 186374
rect 328746 149818 329302 150374
rect 328746 113818 329302 114374
rect 328746 77818 329302 78374
rect 328746 41818 329302 42374
rect 328746 5818 329302 6374
rect 328746 -3782 329302 -3226
rect 329986 708122 330542 708678
rect 329986 691058 330542 691614
rect 329986 655058 330542 655614
rect 329986 619058 330542 619614
rect 329986 583058 330542 583614
rect 329986 547058 330542 547614
rect 329986 511058 330542 511614
rect 329986 475058 330542 475614
rect 329986 439058 330542 439614
rect 329986 403058 330542 403614
rect 329986 367058 330542 367614
rect 329986 331058 330542 331614
rect 329986 295058 330542 295614
rect 329986 259058 330542 259614
rect 329986 223058 330542 223614
rect 329986 187058 330542 187614
rect 329986 151058 330542 151614
rect 329986 115058 330542 115614
rect 329986 79058 330542 79614
rect 329986 43058 330542 43614
rect 329986 7058 330542 7614
rect 329986 -4742 330542 -4186
rect 331226 709082 331782 709638
rect 331226 692298 331782 692854
rect 331226 656298 331782 656854
rect 331226 620298 331782 620854
rect 331226 584298 331782 584854
rect 331226 548298 331782 548854
rect 331226 512298 331782 512854
rect 331226 476298 331782 476854
rect 331226 440298 331782 440854
rect 331226 404298 331782 404854
rect 331226 368298 331782 368854
rect 331226 332298 331782 332854
rect 331226 296298 331782 296854
rect 331226 260298 331782 260854
rect 331226 224298 331782 224854
rect 331226 188298 331782 188854
rect 331226 152298 331782 152854
rect 331226 116298 331782 116854
rect 331226 80298 331782 80854
rect 331226 44298 331782 44854
rect 331226 8298 331782 8854
rect 331226 -5702 331782 -5146
rect 332466 710042 333022 710598
rect 332466 693538 333022 694094
rect 332466 657538 333022 658094
rect 332466 621538 333022 622094
rect 332466 585538 333022 586094
rect 332466 549538 333022 550094
rect 332466 513538 333022 514094
rect 332466 477538 333022 478094
rect 332466 441538 333022 442094
rect 332466 405538 333022 406094
rect 332466 369538 333022 370094
rect 332466 333538 333022 334094
rect 332466 297538 333022 298094
rect 332466 261538 333022 262094
rect 332466 225538 333022 226094
rect 332466 189538 333022 190094
rect 332466 153538 333022 154094
rect 332466 117538 333022 118094
rect 332466 81538 333022 82094
rect 332466 45538 333022 46094
rect 332466 9538 333022 10094
rect 332466 -6662 333022 -6106
rect 333706 711002 334262 711558
rect 333706 694778 334262 695334
rect 333706 658778 334262 659334
rect 333706 622778 334262 623334
rect 333706 586778 334262 587334
rect 333706 550778 334262 551334
rect 333706 514778 334262 515334
rect 333706 478778 334262 479334
rect 333706 442778 334262 443334
rect 333706 406778 334262 407334
rect 333706 370778 334262 371334
rect 333706 334778 334262 335334
rect 333706 298778 334262 299334
rect 333706 262778 334262 263334
rect 333706 226778 334262 227334
rect 333706 190778 334262 191334
rect 333706 154778 334262 155334
rect 333706 118778 334262 119334
rect 333706 82778 334262 83334
rect 333706 46778 334262 47334
rect 333706 10778 334262 11334
rect 333706 -7622 334262 -7066
rect 361026 704282 361582 704838
rect 361026 686098 361582 686654
rect 361026 650098 361582 650654
rect 361026 614098 361582 614654
rect 361026 578098 361582 578654
rect 361026 542098 361582 542654
rect 361026 506098 361582 506654
rect 361026 470098 361582 470654
rect 361026 434098 361582 434654
rect 361026 398098 361582 398654
rect 361026 362098 361582 362654
rect 361026 326098 361582 326654
rect 361026 290098 361582 290654
rect 361026 254098 361582 254654
rect 361026 218098 361582 218654
rect 361026 182098 361582 182654
rect 361026 146098 361582 146654
rect 361026 110098 361582 110654
rect 361026 74098 361582 74654
rect 361026 38098 361582 38654
rect 361026 2098 361582 2654
rect 361026 -902 361582 -346
rect 362266 705242 362822 705798
rect 362266 687338 362822 687894
rect 362266 651338 362822 651894
rect 362266 615338 362822 615894
rect 362266 579338 362822 579894
rect 362266 543338 362822 543894
rect 362266 507338 362822 507894
rect 362266 471338 362822 471894
rect 362266 435338 362822 435894
rect 362266 399338 362822 399894
rect 362266 363338 362822 363894
rect 362266 327338 362822 327894
rect 362266 291338 362822 291894
rect 362266 255338 362822 255894
rect 362266 219338 362822 219894
rect 362266 183338 362822 183894
rect 362266 147338 362822 147894
rect 362266 111338 362822 111894
rect 362266 75338 362822 75894
rect 362266 39338 362822 39894
rect 362266 3338 362822 3894
rect 362266 -1862 362822 -1306
rect 363506 706202 364062 706758
rect 363506 688578 364062 689134
rect 363506 652578 364062 653134
rect 363506 616578 364062 617134
rect 363506 580578 364062 581134
rect 363506 544578 364062 545134
rect 363506 508578 364062 509134
rect 363506 472578 364062 473134
rect 363506 436578 364062 437134
rect 363506 400578 364062 401134
rect 363506 364578 364062 365134
rect 363506 328578 364062 329134
rect 363506 292578 364062 293134
rect 363506 256578 364062 257134
rect 363506 220578 364062 221134
rect 363506 184578 364062 185134
rect 363506 148578 364062 149134
rect 363506 112578 364062 113134
rect 363506 76578 364062 77134
rect 363506 40578 364062 41134
rect 363506 4578 364062 5134
rect 363506 -2822 364062 -2266
rect 364746 707162 365302 707718
rect 364746 689818 365302 690374
rect 364746 653818 365302 654374
rect 364746 617818 365302 618374
rect 364746 581818 365302 582374
rect 364746 545818 365302 546374
rect 364746 509818 365302 510374
rect 364746 473818 365302 474374
rect 364746 437818 365302 438374
rect 364746 401818 365302 402374
rect 364746 365818 365302 366374
rect 364746 329818 365302 330374
rect 364746 293818 365302 294374
rect 364746 257818 365302 258374
rect 364746 221818 365302 222374
rect 364746 185818 365302 186374
rect 364746 149818 365302 150374
rect 364746 113818 365302 114374
rect 364746 77818 365302 78374
rect 364746 41818 365302 42374
rect 364746 5818 365302 6374
rect 364746 -3782 365302 -3226
rect 365986 708122 366542 708678
rect 365986 691058 366542 691614
rect 365986 655058 366542 655614
rect 365986 619058 366542 619614
rect 365986 583058 366542 583614
rect 365986 547058 366542 547614
rect 365986 511058 366542 511614
rect 365986 475058 366542 475614
rect 365986 439058 366542 439614
rect 365986 403058 366542 403614
rect 365986 367058 366542 367614
rect 365986 331058 366542 331614
rect 365986 295058 366542 295614
rect 365986 259058 366542 259614
rect 365986 223058 366542 223614
rect 365986 187058 366542 187614
rect 365986 151058 366542 151614
rect 365986 115058 366542 115614
rect 365986 79058 366542 79614
rect 365986 43058 366542 43614
rect 365986 7058 366542 7614
rect 365986 -4742 366542 -4186
rect 367226 709082 367782 709638
rect 367226 692298 367782 692854
rect 367226 656298 367782 656854
rect 367226 620298 367782 620854
rect 367226 584298 367782 584854
rect 367226 548298 367782 548854
rect 367226 512298 367782 512854
rect 367226 476298 367782 476854
rect 367226 440298 367782 440854
rect 367226 404298 367782 404854
rect 367226 368298 367782 368854
rect 367226 332298 367782 332854
rect 367226 296298 367782 296854
rect 367226 260298 367782 260854
rect 367226 224298 367782 224854
rect 367226 188298 367782 188854
rect 367226 152298 367782 152854
rect 367226 116298 367782 116854
rect 367226 80298 367782 80854
rect 367226 44298 367782 44854
rect 367226 8298 367782 8854
rect 367226 -5702 367782 -5146
rect 368466 710042 369022 710598
rect 368466 693538 369022 694094
rect 368466 657538 369022 658094
rect 368466 621538 369022 622094
rect 368466 585538 369022 586094
rect 368466 549538 369022 550094
rect 368466 513538 369022 514094
rect 368466 477538 369022 478094
rect 368466 441538 369022 442094
rect 368466 405538 369022 406094
rect 368466 369538 369022 370094
rect 368466 333538 369022 334094
rect 368466 297538 369022 298094
rect 368466 261538 369022 262094
rect 368466 225538 369022 226094
rect 368466 189538 369022 190094
rect 368466 153538 369022 154094
rect 368466 117538 369022 118094
rect 368466 81538 369022 82094
rect 368466 45538 369022 46094
rect 368466 9538 369022 10094
rect 368466 -6662 369022 -6106
rect 369706 711002 370262 711558
rect 369706 694778 370262 695334
rect 369706 658778 370262 659334
rect 369706 622778 370262 623334
rect 369706 586778 370262 587334
rect 369706 550778 370262 551334
rect 369706 514778 370262 515334
rect 369706 478778 370262 479334
rect 369706 442778 370262 443334
rect 369706 406778 370262 407334
rect 369706 370778 370262 371334
rect 369706 334778 370262 335334
rect 369706 298778 370262 299334
rect 369706 262778 370262 263334
rect 369706 226778 370262 227334
rect 369706 190778 370262 191334
rect 369706 154778 370262 155334
rect 369706 118778 370262 119334
rect 369706 82778 370262 83334
rect 369706 46778 370262 47334
rect 369706 10778 370262 11334
rect 369706 -7622 370262 -7066
rect 397026 704282 397582 704838
rect 397026 686098 397582 686654
rect 397026 650098 397582 650654
rect 397026 614098 397582 614654
rect 397026 578098 397582 578654
rect 397026 542098 397582 542654
rect 397026 506098 397582 506654
rect 397026 470098 397582 470654
rect 397026 434098 397582 434654
rect 397026 398098 397582 398654
rect 397026 362098 397582 362654
rect 397026 326098 397582 326654
rect 397026 290098 397582 290654
rect 397026 254098 397582 254654
rect 397026 218098 397582 218654
rect 397026 182098 397582 182654
rect 397026 146098 397582 146654
rect 397026 110098 397582 110654
rect 397026 74098 397582 74654
rect 397026 38098 397582 38654
rect 397026 2098 397582 2654
rect 397026 -902 397582 -346
rect 398266 705242 398822 705798
rect 398266 687338 398822 687894
rect 398266 651338 398822 651894
rect 398266 615338 398822 615894
rect 398266 579338 398822 579894
rect 398266 543338 398822 543894
rect 398266 507338 398822 507894
rect 398266 471338 398822 471894
rect 398266 435338 398822 435894
rect 398266 399338 398822 399894
rect 398266 363338 398822 363894
rect 398266 327338 398822 327894
rect 398266 291338 398822 291894
rect 398266 255338 398822 255894
rect 398266 219338 398822 219894
rect 398266 183338 398822 183894
rect 398266 147338 398822 147894
rect 398266 111338 398822 111894
rect 398266 75338 398822 75894
rect 398266 39338 398822 39894
rect 398266 3338 398822 3894
rect 398266 -1862 398822 -1306
rect 399506 706202 400062 706758
rect 399506 688578 400062 689134
rect 399506 652578 400062 653134
rect 399506 616578 400062 617134
rect 399506 580578 400062 581134
rect 399506 544578 400062 545134
rect 399506 508578 400062 509134
rect 399506 472578 400062 473134
rect 399506 436578 400062 437134
rect 399506 400578 400062 401134
rect 399506 364578 400062 365134
rect 399506 328578 400062 329134
rect 399506 292578 400062 293134
rect 399506 256578 400062 257134
rect 399506 220578 400062 221134
rect 399506 184578 400062 185134
rect 399506 148578 400062 149134
rect 399506 112578 400062 113134
rect 399506 76578 400062 77134
rect 399506 40578 400062 41134
rect 399506 4578 400062 5134
rect 399506 -2822 400062 -2266
rect 400746 707162 401302 707718
rect 400746 689818 401302 690374
rect 400746 653818 401302 654374
rect 400746 617818 401302 618374
rect 400746 581818 401302 582374
rect 400746 545818 401302 546374
rect 400746 509818 401302 510374
rect 400746 473818 401302 474374
rect 400746 437818 401302 438374
rect 400746 401818 401302 402374
rect 400746 365818 401302 366374
rect 400746 329818 401302 330374
rect 400746 293818 401302 294374
rect 400746 257818 401302 258374
rect 400746 221818 401302 222374
rect 400746 185818 401302 186374
rect 400746 149818 401302 150374
rect 400746 113818 401302 114374
rect 400746 77818 401302 78374
rect 400746 41818 401302 42374
rect 400746 5818 401302 6374
rect 400746 -3782 401302 -3226
rect 401986 708122 402542 708678
rect 401986 691058 402542 691614
rect 401986 655058 402542 655614
rect 401986 619058 402542 619614
rect 401986 583058 402542 583614
rect 401986 547058 402542 547614
rect 401986 511058 402542 511614
rect 401986 475058 402542 475614
rect 401986 439058 402542 439614
rect 401986 403058 402542 403614
rect 401986 367058 402542 367614
rect 401986 331058 402542 331614
rect 401986 295058 402542 295614
rect 401986 259058 402542 259614
rect 401986 223058 402542 223614
rect 401986 187058 402542 187614
rect 401986 151058 402542 151614
rect 401986 115058 402542 115614
rect 401986 79058 402542 79614
rect 401986 43058 402542 43614
rect 401986 7058 402542 7614
rect 401986 -4742 402542 -4186
rect 403226 709082 403782 709638
rect 403226 692298 403782 692854
rect 403226 656298 403782 656854
rect 403226 620298 403782 620854
rect 403226 584298 403782 584854
rect 403226 548298 403782 548854
rect 403226 512298 403782 512854
rect 403226 476298 403782 476854
rect 403226 440298 403782 440854
rect 403226 404298 403782 404854
rect 403226 368298 403782 368854
rect 403226 332298 403782 332854
rect 403226 296298 403782 296854
rect 403226 260298 403782 260854
rect 403226 224298 403782 224854
rect 403226 188298 403782 188854
rect 403226 152298 403782 152854
rect 403226 116298 403782 116854
rect 403226 80298 403782 80854
rect 403226 44298 403782 44854
rect 403226 8298 403782 8854
rect 403226 -5702 403782 -5146
rect 404466 710042 405022 710598
rect 404466 693538 405022 694094
rect 404466 657538 405022 658094
rect 404466 621538 405022 622094
rect 404466 585538 405022 586094
rect 404466 549538 405022 550094
rect 404466 513538 405022 514094
rect 404466 477538 405022 478094
rect 404466 441538 405022 442094
rect 404466 405538 405022 406094
rect 404466 369538 405022 370094
rect 404466 333538 405022 334094
rect 404466 297538 405022 298094
rect 404466 261538 405022 262094
rect 404466 225538 405022 226094
rect 404466 189538 405022 190094
rect 404466 153538 405022 154094
rect 404466 117538 405022 118094
rect 404466 81538 405022 82094
rect 404466 45538 405022 46094
rect 404466 9538 405022 10094
rect 404466 -6662 405022 -6106
rect 405706 711002 406262 711558
rect 405706 694778 406262 695334
rect 405706 658778 406262 659334
rect 405706 622778 406262 623334
rect 405706 586778 406262 587334
rect 405706 550778 406262 551334
rect 405706 514778 406262 515334
rect 405706 478778 406262 479334
rect 405706 442778 406262 443334
rect 405706 406778 406262 407334
rect 405706 370778 406262 371334
rect 405706 334778 406262 335334
rect 405706 298778 406262 299334
rect 405706 262778 406262 263334
rect 405706 226778 406262 227334
rect 405706 190778 406262 191334
rect 405706 154778 406262 155334
rect 405706 118778 406262 119334
rect 405706 82778 406262 83334
rect 405706 46778 406262 47334
rect 405706 10778 406262 11334
rect 405706 -7622 406262 -7066
rect 433026 704282 433582 704838
rect 433026 686098 433582 686654
rect 433026 650098 433582 650654
rect 433026 614098 433582 614654
rect 433026 578098 433582 578654
rect 433026 542098 433582 542654
rect 433026 506098 433582 506654
rect 433026 470098 433582 470654
rect 433026 434098 433582 434654
rect 433026 398098 433582 398654
rect 433026 362098 433582 362654
rect 433026 326098 433582 326654
rect 433026 290098 433582 290654
rect 433026 254098 433582 254654
rect 433026 218098 433582 218654
rect 433026 182098 433582 182654
rect 433026 146098 433582 146654
rect 433026 110098 433582 110654
rect 433026 74098 433582 74654
rect 433026 38098 433582 38654
rect 433026 2098 433582 2654
rect 433026 -902 433582 -346
rect 434266 705242 434822 705798
rect 434266 687338 434822 687894
rect 434266 651338 434822 651894
rect 434266 615338 434822 615894
rect 434266 579338 434822 579894
rect 434266 543338 434822 543894
rect 434266 507338 434822 507894
rect 434266 471338 434822 471894
rect 434266 435338 434822 435894
rect 434266 399338 434822 399894
rect 434266 363338 434822 363894
rect 434266 327338 434822 327894
rect 434266 291338 434822 291894
rect 434266 255338 434822 255894
rect 434266 219338 434822 219894
rect 434266 183338 434822 183894
rect 434266 147338 434822 147894
rect 434266 111338 434822 111894
rect 434266 75338 434822 75894
rect 434266 39338 434822 39894
rect 434266 3338 434822 3894
rect 434266 -1862 434822 -1306
rect 435506 706202 436062 706758
rect 435506 688578 436062 689134
rect 435506 652578 436062 653134
rect 435506 616578 436062 617134
rect 435506 580578 436062 581134
rect 435506 544578 436062 545134
rect 435506 508578 436062 509134
rect 435506 472578 436062 473134
rect 435506 436578 436062 437134
rect 435506 400578 436062 401134
rect 435506 364578 436062 365134
rect 435506 328578 436062 329134
rect 435506 292578 436062 293134
rect 435506 256578 436062 257134
rect 435506 220578 436062 221134
rect 435506 184578 436062 185134
rect 435506 148578 436062 149134
rect 435506 112578 436062 113134
rect 435506 76578 436062 77134
rect 435506 40578 436062 41134
rect 435506 4578 436062 5134
rect 435506 -2822 436062 -2266
rect 436746 707162 437302 707718
rect 436746 689818 437302 690374
rect 436746 653818 437302 654374
rect 436746 617818 437302 618374
rect 436746 581818 437302 582374
rect 436746 545818 437302 546374
rect 436746 509818 437302 510374
rect 436746 473818 437302 474374
rect 436746 437818 437302 438374
rect 436746 401818 437302 402374
rect 436746 365818 437302 366374
rect 436746 329818 437302 330374
rect 436746 293818 437302 294374
rect 436746 257818 437302 258374
rect 436746 221818 437302 222374
rect 436746 185818 437302 186374
rect 436746 149818 437302 150374
rect 436746 113818 437302 114374
rect 436746 77818 437302 78374
rect 436746 41818 437302 42374
rect 436746 5818 437302 6374
rect 436746 -3782 437302 -3226
rect 437986 708122 438542 708678
rect 437986 691058 438542 691614
rect 437986 655058 438542 655614
rect 437986 619058 438542 619614
rect 437986 583058 438542 583614
rect 437986 547058 438542 547614
rect 437986 511058 438542 511614
rect 437986 475058 438542 475614
rect 437986 439058 438542 439614
rect 437986 403058 438542 403614
rect 437986 367058 438542 367614
rect 437986 331058 438542 331614
rect 437986 295058 438542 295614
rect 437986 259058 438542 259614
rect 437986 223058 438542 223614
rect 437986 187058 438542 187614
rect 437986 151058 438542 151614
rect 437986 115058 438542 115614
rect 437986 79058 438542 79614
rect 437986 43058 438542 43614
rect 437986 7058 438542 7614
rect 437986 -4742 438542 -4186
rect 439226 709082 439782 709638
rect 439226 692298 439782 692854
rect 439226 656298 439782 656854
rect 439226 620298 439782 620854
rect 439226 584298 439782 584854
rect 439226 548298 439782 548854
rect 439226 512298 439782 512854
rect 439226 476298 439782 476854
rect 439226 440298 439782 440854
rect 439226 404298 439782 404854
rect 439226 368298 439782 368854
rect 439226 332298 439782 332854
rect 439226 296298 439782 296854
rect 439226 260298 439782 260854
rect 439226 224298 439782 224854
rect 439226 188298 439782 188854
rect 439226 152298 439782 152854
rect 439226 116298 439782 116854
rect 439226 80298 439782 80854
rect 439226 44298 439782 44854
rect 439226 8298 439782 8854
rect 439226 -5702 439782 -5146
rect 440466 710042 441022 710598
rect 440466 693538 441022 694094
rect 440466 657538 441022 658094
rect 440466 621538 441022 622094
rect 440466 585538 441022 586094
rect 440466 549538 441022 550094
rect 440466 513538 441022 514094
rect 440466 477538 441022 478094
rect 440466 441538 441022 442094
rect 440466 405538 441022 406094
rect 440466 369538 441022 370094
rect 440466 333538 441022 334094
rect 440466 297538 441022 298094
rect 440466 261538 441022 262094
rect 440466 225538 441022 226094
rect 440466 189538 441022 190094
rect 440466 153538 441022 154094
rect 440466 117538 441022 118094
rect 440466 81538 441022 82094
rect 440466 45538 441022 46094
rect 440466 9538 441022 10094
rect 440466 -6662 441022 -6106
rect 441706 711002 442262 711558
rect 441706 694778 442262 695334
rect 441706 658778 442262 659334
rect 441706 622778 442262 623334
rect 441706 586778 442262 587334
rect 441706 550778 442262 551334
rect 441706 514778 442262 515334
rect 441706 478778 442262 479334
rect 441706 442778 442262 443334
rect 441706 406778 442262 407334
rect 441706 370778 442262 371334
rect 441706 334778 442262 335334
rect 441706 298778 442262 299334
rect 441706 262778 442262 263334
rect 441706 226778 442262 227334
rect 441706 190778 442262 191334
rect 441706 154778 442262 155334
rect 441706 118778 442262 119334
rect 441706 82778 442262 83334
rect 441706 46778 442262 47334
rect 441706 10778 442262 11334
rect 441706 -7622 442262 -7066
rect 469026 704282 469582 704838
rect 469026 686098 469582 686654
rect 469026 650098 469582 650654
rect 469026 614098 469582 614654
rect 469026 578098 469582 578654
rect 469026 542098 469582 542654
rect 469026 506098 469582 506654
rect 469026 470098 469582 470654
rect 469026 434098 469582 434654
rect 469026 398098 469582 398654
rect 469026 362098 469582 362654
rect 469026 326098 469582 326654
rect 469026 290098 469582 290654
rect 469026 254098 469582 254654
rect 469026 218098 469582 218654
rect 469026 182098 469582 182654
rect 469026 146098 469582 146654
rect 469026 110098 469582 110654
rect 469026 74098 469582 74654
rect 469026 38098 469582 38654
rect 469026 2098 469582 2654
rect 469026 -902 469582 -346
rect 470266 705242 470822 705798
rect 470266 687338 470822 687894
rect 470266 651338 470822 651894
rect 470266 615338 470822 615894
rect 470266 579338 470822 579894
rect 470266 543338 470822 543894
rect 470266 507338 470822 507894
rect 470266 471338 470822 471894
rect 470266 435338 470822 435894
rect 470266 399338 470822 399894
rect 470266 363338 470822 363894
rect 470266 327780 470272 327894
rect 470272 327780 470816 327894
rect 470816 327780 470822 327894
rect 470266 327338 470822 327780
rect 470266 291338 470822 291894
rect 470266 255338 470822 255894
rect 470266 219338 470822 219894
rect 470266 183338 470822 183894
rect 470266 147338 470822 147894
rect 470266 111338 470822 111894
rect 470266 75338 470822 75894
rect 470266 39338 470822 39894
rect 470266 3338 470822 3894
rect 470266 -1862 470822 -1306
rect 471506 706202 472062 706758
rect 471506 688578 472062 689134
rect 471506 652578 472062 653134
rect 471506 616578 472062 617134
rect 471506 580578 472062 581134
rect 471506 544578 472062 545134
rect 471506 508578 472062 509134
rect 471506 472578 472062 473134
rect 471506 436578 472062 437134
rect 471506 400578 472062 401134
rect 472746 707162 473302 707718
rect 472746 689818 473302 690374
rect 472746 653818 473302 654374
rect 472746 617818 473302 618374
rect 472746 581818 473302 582374
rect 472746 545818 473302 546374
rect 472746 509818 473302 510374
rect 472746 473818 473302 474374
rect 472746 437818 473302 438374
rect 472746 401818 473302 402374
rect 473986 708122 474542 708678
rect 473986 691058 474542 691614
rect 473986 655058 474542 655614
rect 473986 619058 474542 619614
rect 473986 583058 474542 583614
rect 473986 547058 474542 547614
rect 473986 511058 474542 511614
rect 473986 475058 474542 475614
rect 473986 439058 474542 439614
rect 473986 403058 474542 403614
rect 475226 709082 475782 709638
rect 475226 692298 475782 692854
rect 475226 656298 475782 656854
rect 475226 620298 475782 620854
rect 475226 584298 475782 584854
rect 475226 548298 475782 548854
rect 475226 512298 475782 512854
rect 475226 476298 475782 476854
rect 475226 440298 475782 440854
rect 475226 404298 475782 404854
rect 476466 710042 477022 710598
rect 476466 693538 477022 694094
rect 476466 657538 477022 658094
rect 476466 621538 477022 622094
rect 476466 585538 477022 586094
rect 476466 549538 477022 550094
rect 476466 513538 477022 514094
rect 476466 477538 477022 478094
rect 476466 441538 477022 442094
rect 476466 405538 477022 406094
rect 477706 711002 478262 711558
rect 477706 694778 478262 695334
rect 477706 658778 478262 659334
rect 477706 622778 478262 623334
rect 477706 586778 478262 587334
rect 477706 550778 478262 551334
rect 477706 514778 478262 515334
rect 477706 478778 478262 479334
rect 477706 442778 478262 443334
rect 477706 406778 478262 407334
rect 477706 370778 478262 371334
rect 505026 704282 505582 704838
rect 505026 686098 505582 686654
rect 505026 650098 505582 650654
rect 505026 614098 505582 614654
rect 505026 578098 505582 578654
rect 505026 542098 505582 542654
rect 505026 506098 505582 506654
rect 505026 470098 505582 470654
rect 505026 434098 505582 434654
rect 505026 398098 505582 398654
rect 471506 364578 472062 365134
rect 471506 328578 472062 329134
rect 471506 292578 472062 293134
rect 472746 365883 472982 366119
rect 473066 365883 473302 366119
rect 472746 329818 473302 330374
rect 472746 293818 473302 294374
rect 473986 331058 474542 331614
rect 473986 295058 474542 295614
rect 475226 332298 475782 332854
rect 475226 296298 475782 296854
rect 476466 333538 477022 334094
rect 476466 297538 477022 298094
rect 477706 334778 478262 335334
rect 477706 298778 478262 299334
rect 505026 362098 505582 362654
rect 505026 326098 505582 326654
rect 505026 290098 505582 290654
rect 471506 256578 472062 257134
rect 471506 220578 472062 221134
rect 471506 184578 472062 185134
rect 471506 148578 472062 149134
rect 471506 112578 472062 113134
rect 471506 76578 472062 77134
rect 471506 40578 472062 41134
rect 471506 4578 472062 5134
rect 471506 -2822 472062 -2266
rect 472746 257818 473302 258374
rect 472746 221818 473302 222374
rect 472746 185818 473302 186374
rect 472746 149818 473302 150374
rect 472746 113818 473302 114374
rect 472746 77818 473302 78374
rect 472746 41818 473302 42374
rect 472746 5818 473302 6374
rect 472746 -3782 473302 -3226
rect 473986 259058 474542 259614
rect 473986 223058 474542 223614
rect 473986 187058 474542 187614
rect 473986 151058 474542 151614
rect 473986 115058 474542 115614
rect 473986 79058 474542 79614
rect 473986 43058 474542 43614
rect 473986 7058 474542 7614
rect 473986 -4742 474542 -4186
rect 475226 260298 475782 260854
rect 475226 224298 475782 224854
rect 475226 188298 475782 188854
rect 475226 152298 475782 152854
rect 475226 116298 475782 116854
rect 475226 80298 475782 80854
rect 475226 44298 475782 44854
rect 475226 8298 475782 8854
rect 475226 -5702 475782 -5146
rect 476466 225538 477022 226094
rect 476466 189538 477022 190094
rect 476466 153538 477022 154094
rect 476466 117538 477022 118094
rect 476466 81538 477022 82094
rect 476466 45538 477022 46094
rect 476466 9538 477022 10094
rect 476466 -6662 477022 -6106
rect 477706 226778 478262 227334
rect 477706 190778 478262 191334
rect 477706 154778 478262 155334
rect 477706 118778 478262 119334
rect 477706 82778 478262 83334
rect 477706 46778 478262 47334
rect 477706 10778 478262 11334
rect 477706 -7622 478262 -7066
rect 505026 254098 505582 254654
rect 505026 218098 505582 218654
rect 505026 182098 505582 182654
rect 505026 146098 505582 146654
rect 505026 110098 505582 110654
rect 505026 74098 505582 74654
rect 505026 38098 505582 38654
rect 505026 2098 505582 2654
rect 505026 -902 505582 -346
rect 506266 705242 506822 705798
rect 506266 687338 506822 687894
rect 506266 651338 506822 651894
rect 506266 615338 506822 615894
rect 506266 579338 506822 579894
rect 506266 543338 506822 543894
rect 506266 507338 506822 507894
rect 506266 471338 506822 471894
rect 506266 435338 506822 435894
rect 506266 399338 506822 399894
rect 506266 363338 506822 363894
rect 506266 327338 506822 327894
rect 506266 291338 506822 291894
rect 506266 255338 506822 255894
rect 506266 219338 506822 219894
rect 506266 183338 506822 183894
rect 506266 147338 506822 147894
rect 506266 111338 506822 111894
rect 506266 75338 506822 75894
rect 506266 39338 506822 39894
rect 506266 3338 506822 3894
rect 506266 -1862 506822 -1306
rect 507506 706202 508062 706758
rect 507506 688578 508062 689134
rect 507506 652578 508062 653134
rect 507506 616578 508062 617134
rect 507506 580578 508062 581134
rect 507506 544578 508062 545134
rect 507506 508578 508062 509134
rect 507506 472578 508062 473134
rect 507506 436578 508062 437134
rect 507506 400578 508062 401134
rect 507506 364578 508062 365134
rect 507506 328578 508062 329134
rect 507506 292578 508062 293134
rect 507506 256578 508062 257134
rect 507506 220578 508062 221134
rect 507506 184578 508062 185134
rect 507506 148578 508062 149134
rect 507506 112578 508062 113134
rect 507506 76578 508062 77134
rect 507506 40578 508062 41134
rect 507506 4578 508062 5134
rect 507506 -2822 508062 -2266
rect 508746 707162 509302 707718
rect 508746 689818 509302 690374
rect 508746 653818 509302 654374
rect 508746 617818 509302 618374
rect 508746 581818 509302 582374
rect 508746 545818 509302 546374
rect 508746 509818 509302 510374
rect 508746 473818 509302 474374
rect 508746 437818 509302 438374
rect 508746 401818 509302 402374
rect 508746 365818 509302 366374
rect 508746 329818 509302 330374
rect 508746 293818 509302 294374
rect 508746 257818 509302 258374
rect 508746 221818 509302 222374
rect 508746 185818 509302 186374
rect 508746 149818 509302 150374
rect 508746 113818 509302 114374
rect 508746 77818 509302 78374
rect 508746 41818 509302 42374
rect 508746 5818 509302 6374
rect 508746 -3782 509302 -3226
rect 509986 708122 510542 708678
rect 509986 691058 510542 691614
rect 509986 655058 510542 655614
rect 509986 619058 510542 619614
rect 509986 583058 510542 583614
rect 509986 547058 510542 547614
rect 509986 511058 510542 511614
rect 509986 475058 510542 475614
rect 509986 439058 510542 439614
rect 509986 403058 510542 403614
rect 509986 367058 510542 367614
rect 509986 331058 510542 331614
rect 509986 295058 510542 295614
rect 509986 259058 510542 259614
rect 509986 223058 510542 223614
rect 509986 187058 510542 187614
rect 509986 151058 510542 151614
rect 509986 115058 510542 115614
rect 509986 79058 510542 79614
rect 509986 43058 510542 43614
rect 509986 7058 510542 7614
rect 509986 -4742 510542 -4186
rect 511226 709082 511782 709638
rect 511226 692298 511782 692854
rect 511226 656298 511782 656854
rect 511226 620298 511782 620854
rect 511226 584298 511782 584854
rect 511226 548298 511782 548854
rect 511226 512298 511782 512854
rect 511226 476298 511782 476854
rect 511226 440298 511782 440854
rect 511226 404298 511782 404854
rect 511226 368298 511782 368854
rect 511226 332298 511782 332854
rect 511226 296298 511782 296854
rect 511226 260298 511782 260854
rect 511226 224298 511782 224854
rect 511226 188298 511782 188854
rect 511226 152298 511782 152854
rect 511226 116298 511782 116854
rect 511226 80298 511782 80854
rect 511226 44298 511782 44854
rect 511226 8298 511782 8854
rect 511226 -5702 511782 -5146
rect 512466 710042 513022 710598
rect 512466 693538 513022 694094
rect 512466 657538 513022 658094
rect 512466 621538 513022 622094
rect 512466 585538 513022 586094
rect 512466 549538 513022 550094
rect 512466 513538 513022 514094
rect 512466 477538 513022 478094
rect 512466 441538 513022 442094
rect 512466 405538 513022 406094
rect 512466 369538 513022 370094
rect 512466 333538 513022 334094
rect 512466 297538 513022 298094
rect 512466 261538 513022 262094
rect 512466 225538 513022 226094
rect 512466 189538 513022 190094
rect 512466 153538 513022 154094
rect 512466 117538 513022 118094
rect 512466 81538 513022 82094
rect 512466 45538 513022 46094
rect 512466 9538 513022 10094
rect 512466 -6662 513022 -6106
rect 513706 711002 514262 711558
rect 513706 694778 514262 695334
rect 513706 658778 514262 659334
rect 513706 622778 514262 623334
rect 513706 586778 514262 587334
rect 513706 550778 514262 551334
rect 513706 514778 514262 515334
rect 513706 478778 514262 479334
rect 541026 704282 541582 704838
rect 541026 686098 541582 686654
rect 541026 650098 541582 650654
rect 541026 614098 541582 614654
rect 541026 578098 541582 578654
rect 541026 542098 541582 542654
rect 541026 506098 541582 506654
rect 541026 470098 541582 470654
rect 542266 705242 542822 705798
rect 542266 687338 542822 687894
rect 542266 651338 542822 651894
rect 542266 615338 542822 615894
rect 542266 579338 542822 579894
rect 542266 543338 542822 543894
rect 542266 507338 542822 507894
rect 542266 471338 542822 471894
rect 543506 706202 544062 706758
rect 543506 688578 544062 689134
rect 543506 652578 544062 653134
rect 543506 616578 544062 617134
rect 543506 580578 544062 581134
rect 543506 544578 544062 545134
rect 543506 508578 544062 509134
rect 543506 472578 544062 473134
rect 544746 707162 545302 707718
rect 544746 689818 545302 690374
rect 544746 653818 545302 654374
rect 544746 617818 545302 618374
rect 544746 581818 545302 582374
rect 544746 545818 545302 546374
rect 544746 509818 545302 510374
rect 544746 473818 545302 474374
rect 545986 708122 546542 708678
rect 545986 691058 546542 691614
rect 545986 655058 546542 655614
rect 545986 619058 546542 619614
rect 545986 583058 546542 583614
rect 545986 547058 546542 547614
rect 545986 511058 546542 511614
rect 545986 475058 546542 475614
rect 547226 709082 547782 709638
rect 547226 692298 547782 692854
rect 547226 656298 547782 656854
rect 547226 620298 547782 620854
rect 547226 584298 547782 584854
rect 547226 548298 547782 548854
rect 547226 512298 547782 512854
rect 547226 476298 547782 476854
rect 513706 442778 514262 443334
rect 547226 440298 547782 440854
rect 540918 435658 541154 435894
rect 540918 435338 541154 435574
rect 542850 435658 543086 435894
rect 542850 435338 543086 435574
rect 544782 435658 545018 435894
rect 544782 435338 545018 435574
rect 546714 435658 546950 435894
rect 546714 435338 546950 435574
rect 539952 434418 540188 434654
rect 539952 434098 540188 434334
rect 541884 434418 542120 434654
rect 541884 434098 542120 434334
rect 543816 434418 544052 434654
rect 543816 434098 544052 434334
rect 545748 434418 545984 434654
rect 545748 434098 545984 434334
rect 513706 406778 514262 407334
rect 547226 404298 547782 404854
rect 540918 399658 541154 399894
rect 540918 399338 541154 399574
rect 542850 399658 543086 399894
rect 542850 399338 543086 399574
rect 544782 399658 545018 399894
rect 544782 399338 545018 399574
rect 546714 399658 546950 399894
rect 546714 399338 546950 399574
rect 539952 398418 540188 398654
rect 539952 398098 540188 398334
rect 541884 398418 542120 398654
rect 541884 398098 542120 398334
rect 543816 398418 544052 398654
rect 543816 398098 544052 398334
rect 545748 398418 545984 398654
rect 545748 398098 545984 398334
rect 513706 370778 514262 371334
rect 547226 368298 547782 368854
rect 540918 363658 541154 363894
rect 540918 363338 541154 363574
rect 542850 363658 543086 363894
rect 542850 363338 543086 363574
rect 544782 363658 545018 363894
rect 544782 363338 545018 363574
rect 546714 363658 546950 363894
rect 546714 363338 546950 363574
rect 539952 362418 540188 362654
rect 539952 362098 540188 362334
rect 541884 362418 542120 362654
rect 541884 362098 542120 362334
rect 543816 362418 544052 362654
rect 543816 362098 544052 362334
rect 545748 362418 545984 362654
rect 545748 362098 545984 362334
rect 513706 334778 514262 335334
rect 547226 332298 547782 332854
rect 540918 327658 541154 327894
rect 540918 327338 541154 327574
rect 542850 327658 543086 327894
rect 542850 327338 543086 327574
rect 544782 327658 545018 327894
rect 544782 327338 545018 327574
rect 546714 327658 546950 327894
rect 546714 327338 546950 327574
rect 539952 326418 540188 326654
rect 539952 326098 540188 326334
rect 541884 326418 542120 326654
rect 541884 326098 542120 326334
rect 543816 326418 544052 326654
rect 543816 326098 544052 326334
rect 545748 326418 545984 326654
rect 545748 326098 545984 326334
rect 513706 298778 514262 299334
rect 547226 296298 547782 296854
rect 540918 291658 541154 291894
rect 540918 291338 541154 291574
rect 542850 291658 543086 291894
rect 542850 291338 543086 291574
rect 544782 291658 545018 291894
rect 544782 291338 545018 291574
rect 546714 291658 546950 291894
rect 546714 291338 546950 291574
rect 539952 290418 540188 290654
rect 539952 290098 540188 290334
rect 541884 290418 542120 290654
rect 541884 290098 542120 290334
rect 543816 290418 544052 290654
rect 543816 290098 544052 290334
rect 545748 290418 545984 290654
rect 545748 290098 545984 290334
rect 513706 262778 514262 263334
rect 513706 226778 514262 227334
rect 513706 190778 514262 191334
rect 513706 154778 514262 155334
rect 513706 118778 514262 119334
rect 513706 82778 514262 83334
rect 513706 46778 514262 47334
rect 513706 10778 514262 11334
rect 513706 -7622 514262 -7066
rect 541026 254098 541582 254654
rect 541026 218098 541582 218654
rect 541026 182098 541582 182654
rect 541026 146098 541582 146654
rect 541026 110098 541582 110654
rect 541026 74098 541582 74654
rect 541026 38098 541582 38654
rect 541026 2098 541582 2654
rect 541026 -902 541582 -346
rect 542266 255338 542822 255894
rect 542266 219338 542822 219894
rect 542266 183338 542822 183894
rect 542266 147338 542822 147894
rect 542266 111338 542822 111894
rect 542266 75338 542822 75894
rect 542266 39338 542822 39894
rect 542266 3338 542822 3894
rect 542266 -1862 542822 -1306
rect 543506 256578 544062 257134
rect 543506 220578 544062 221134
rect 543506 184578 544062 185134
rect 543506 148578 544062 149134
rect 543506 112578 544062 113134
rect 543506 76578 544062 77134
rect 543506 40578 544062 41134
rect 543506 4578 544062 5134
rect 543506 -2822 544062 -2266
rect 544746 257818 545302 258374
rect 544746 221818 545302 222374
rect 544746 185818 545302 186374
rect 544746 149818 545302 150374
rect 544746 113818 545302 114374
rect 544746 77818 545302 78374
rect 544746 41818 545302 42374
rect 544746 5818 545302 6374
rect 544746 -3782 545302 -3226
rect 545986 259058 546542 259614
rect 545986 223058 546542 223614
rect 545986 187058 546542 187614
rect 545986 151058 546542 151614
rect 545986 115058 546542 115614
rect 545986 79058 546542 79614
rect 545986 43058 546542 43614
rect 545986 7058 546542 7614
rect 545986 -4742 546542 -4186
rect 547226 260298 547782 260854
rect 547226 224298 547782 224854
rect 547226 188298 547782 188854
rect 547226 152298 547782 152854
rect 547226 116298 547782 116854
rect 547226 80298 547782 80854
rect 547226 44298 547782 44854
rect 547226 8298 547782 8854
rect 547226 -5702 547782 -5146
rect 548466 710042 549022 710598
rect 548466 693538 549022 694094
rect 548466 657538 549022 658094
rect 548466 621538 549022 622094
rect 548466 585538 549022 586094
rect 548466 549538 549022 550094
rect 548466 513538 549022 514094
rect 548466 477538 549022 478094
rect 548466 441538 549022 442094
rect 548466 405538 549022 406094
rect 548466 369538 549022 370094
rect 548466 333538 549022 334094
rect 548466 297538 549022 298094
rect 548466 261538 549022 262094
rect 548466 225538 549022 226094
rect 548466 189538 549022 190094
rect 548466 153538 549022 154094
rect 548466 117538 549022 118094
rect 548466 81538 549022 82094
rect 548466 45538 549022 46094
rect 548466 9538 549022 10094
rect 548466 -6662 549022 -6106
rect 549706 711002 550262 711558
rect 549706 694778 550262 695334
rect 549706 658778 550262 659334
rect 549706 622778 550262 623334
rect 549706 586778 550262 587334
rect 549706 550778 550262 551334
rect 549706 514778 550262 515334
rect 549706 478778 550262 479334
rect 549706 442778 550262 443334
rect 549706 406778 550262 407334
rect 549706 370778 550262 371334
rect 549706 334778 550262 335334
rect 549706 298778 550262 299334
rect 549706 262778 550262 263334
rect 549706 226778 550262 227334
rect 549706 190778 550262 191334
rect 549706 154778 550262 155334
rect 549706 118778 550262 119334
rect 549706 82778 550262 83334
rect 549706 46778 550262 47334
rect 549706 10778 550262 11334
rect 549706 -7622 550262 -7066
rect 577026 704282 577582 704838
rect 577026 686098 577582 686654
rect 577026 650098 577582 650654
rect 577026 614098 577582 614654
rect 577026 578098 577582 578654
rect 577026 542098 577582 542654
rect 577026 506098 577582 506654
rect 577026 470098 577582 470654
rect 577026 434098 577582 434654
rect 577026 398098 577582 398654
rect 577026 362098 577582 362654
rect 577026 326098 577582 326654
rect 577026 290098 577582 290654
rect 577026 254098 577582 254654
rect 577026 218098 577582 218654
rect 577026 182098 577582 182654
rect 577026 146098 577582 146654
rect 577026 110098 577582 110654
rect 577026 74098 577582 74654
rect 577026 38098 577582 38654
rect 577026 2098 577582 2654
rect 577026 -902 577582 -346
rect 578266 705242 578822 705798
rect 578266 687338 578822 687894
rect 578266 651338 578822 651894
rect 578266 615338 578822 615894
rect 578266 579338 578822 579894
rect 578266 543338 578822 543894
rect 578266 507338 578822 507894
rect 578266 471338 578822 471894
rect 578266 435338 578822 435894
rect 578266 399338 578822 399894
rect 578266 363338 578822 363894
rect 578266 327338 578822 327894
rect 578266 291338 578822 291894
rect 578266 255338 578822 255894
rect 578266 219338 578822 219894
rect 578266 183338 578822 183894
rect 578266 147338 578822 147894
rect 578266 111338 578822 111894
rect 578266 75338 578822 75894
rect 578266 39338 578822 39894
rect 578266 3338 578822 3894
rect 578266 -1862 578822 -1306
rect 579506 706202 580062 706758
rect 579506 688578 580062 689134
rect 579506 652578 580062 653134
rect 579506 616578 580062 617134
rect 579506 580578 580062 581134
rect 579506 544578 580062 545134
rect 579506 508578 580062 509134
rect 579506 472578 580062 473134
rect 579506 436578 580062 437134
rect 579506 400578 580062 401134
rect 579506 364578 580062 365134
rect 579506 328578 580062 329134
rect 579506 292578 580062 293134
rect 579506 256578 580062 257134
rect 579506 220578 580062 221134
rect 579506 184578 580062 185134
rect 579506 148578 580062 149134
rect 579506 112578 580062 113134
rect 579506 76578 580062 77134
rect 579506 40578 580062 41134
rect 579506 4578 580062 5134
rect 579506 -2822 580062 -2266
rect 580746 707162 581302 707718
rect 580746 689818 581302 690374
rect 580746 653818 581302 654374
rect 580746 617818 581302 618374
rect 580746 581818 581302 582374
rect 580746 545818 581302 546374
rect 580746 509818 581302 510374
rect 580746 473818 581302 474374
rect 580746 437818 581302 438374
rect 580746 401818 581302 402374
rect 580746 365818 581302 366374
rect 580746 329818 581302 330374
rect 580746 293818 581302 294374
rect 580746 257818 581302 258374
rect 580746 221818 581302 222374
rect 580746 185818 581302 186374
rect 580746 149818 581302 150374
rect 580746 113818 581302 114374
rect 580746 77818 581302 78374
rect 580746 41818 581302 42374
rect 580746 5818 581302 6374
rect 580746 -3782 581302 -3226
rect 592062 711002 592618 711558
rect 591102 710042 591658 710598
rect 590142 709082 590698 709638
rect 581986 708122 582542 708678
rect 589182 708122 589738 708678
rect 588222 707162 588778 707718
rect 587262 706202 587818 706758
rect 586302 705242 586858 705798
rect 581986 691058 582542 691614
rect 581986 655058 582542 655614
rect 581986 619058 582542 619614
rect 581986 583058 582542 583614
rect 581986 547058 582542 547614
rect 581986 511058 582542 511614
rect 581986 475058 582542 475614
rect 581986 439058 582542 439614
rect 581986 403058 582542 403614
rect 581986 367058 582542 367614
rect 581986 331058 582542 331614
rect 581986 295058 582542 295614
rect 581986 259058 582542 259614
rect 581986 223058 582542 223614
rect 581986 187058 582542 187614
rect 581986 151058 582542 151614
rect 581986 115058 582542 115614
rect 581986 79058 582542 79614
rect 581986 43058 582542 43614
rect 581986 7058 582542 7614
rect 585342 704282 585898 704838
rect 585342 686098 585898 686654
rect 585342 650098 585898 650654
rect 585342 614098 585898 614654
rect 585342 578098 585898 578654
rect 585342 542098 585898 542654
rect 585342 506098 585898 506654
rect 585342 470098 585898 470654
rect 585342 434098 585898 434654
rect 585342 398098 585898 398654
rect 585342 362098 585898 362654
rect 585342 326098 585898 326654
rect 585342 290098 585898 290654
rect 585342 254098 585898 254654
rect 585342 218098 585898 218654
rect 585342 182098 585898 182654
rect 585342 146098 585898 146654
rect 585342 110098 585898 110654
rect 585342 74098 585898 74654
rect 585342 38098 585898 38654
rect 585342 2098 585898 2654
rect 585342 -902 585898 -346
rect 586302 687338 586858 687894
rect 586302 651338 586858 651894
rect 586302 615338 586858 615894
rect 586302 579338 586858 579894
rect 586302 543338 586858 543894
rect 586302 507338 586858 507894
rect 586302 471338 586858 471894
rect 586302 435338 586858 435894
rect 586302 399338 586858 399894
rect 586302 363338 586858 363894
rect 586302 327338 586858 327894
rect 586302 291338 586858 291894
rect 586302 255338 586858 255894
rect 586302 219338 586858 219894
rect 586302 183338 586858 183894
rect 586302 147338 586858 147894
rect 586302 111338 586858 111894
rect 586302 75338 586858 75894
rect 586302 39338 586858 39894
rect 586302 3338 586858 3894
rect 586302 -1862 586858 -1306
rect 587262 688578 587818 689134
rect 587262 652578 587818 653134
rect 587262 616578 587818 617134
rect 587262 580578 587818 581134
rect 587262 544578 587818 545134
rect 587262 508578 587818 509134
rect 587262 472578 587818 473134
rect 587262 436578 587818 437134
rect 587262 400578 587818 401134
rect 587262 364578 587818 365134
rect 587262 328578 587818 329134
rect 587262 292578 587818 293134
rect 587262 256578 587818 257134
rect 587262 220578 587818 221134
rect 587262 184578 587818 185134
rect 587262 148578 587818 149134
rect 587262 112578 587818 113134
rect 587262 76578 587818 77134
rect 587262 40578 587818 41134
rect 587262 4578 587818 5134
rect 587262 -2822 587818 -2266
rect 588222 689818 588778 690374
rect 588222 653818 588778 654374
rect 588222 617818 588778 618374
rect 588222 581818 588778 582374
rect 588222 545818 588778 546374
rect 588222 509818 588778 510374
rect 588222 473818 588778 474374
rect 588222 437818 588778 438374
rect 588222 401818 588778 402374
rect 588222 365818 588778 366374
rect 588222 329818 588778 330374
rect 588222 293818 588778 294374
rect 588222 257818 588778 258374
rect 588222 221818 588778 222374
rect 588222 185818 588778 186374
rect 588222 149818 588778 150374
rect 588222 113818 588778 114374
rect 588222 77818 588778 78374
rect 588222 41818 588778 42374
rect 588222 5818 588778 6374
rect 588222 -3782 588778 -3226
rect 589182 691058 589738 691614
rect 589182 655058 589738 655614
rect 589182 619058 589738 619614
rect 589182 583058 589738 583614
rect 589182 547058 589738 547614
rect 589182 511058 589738 511614
rect 589182 475058 589738 475614
rect 589182 439058 589738 439614
rect 589182 403058 589738 403614
rect 589182 367058 589738 367614
rect 589182 331058 589738 331614
rect 589182 295058 589738 295614
rect 589182 259058 589738 259614
rect 589182 223058 589738 223614
rect 589182 187058 589738 187614
rect 589182 151058 589738 151614
rect 589182 115058 589738 115614
rect 589182 79058 589738 79614
rect 589182 43058 589738 43614
rect 589182 7058 589738 7614
rect 581986 -4742 582542 -4186
rect 589182 -4742 589738 -4186
rect 590142 692298 590698 692854
rect 590142 656298 590698 656854
rect 590142 620298 590698 620854
rect 590142 584298 590698 584854
rect 590142 548298 590698 548854
rect 590142 512298 590698 512854
rect 590142 476298 590698 476854
rect 590142 440298 590698 440854
rect 590142 404298 590698 404854
rect 590142 368298 590698 368854
rect 590142 332298 590698 332854
rect 590142 296298 590698 296854
rect 590142 260298 590698 260854
rect 590142 224298 590698 224854
rect 590142 188298 590698 188854
rect 590142 152298 590698 152854
rect 590142 116298 590698 116854
rect 590142 80298 590698 80854
rect 590142 44298 590698 44854
rect 590142 8298 590698 8854
rect 590142 -5702 590698 -5146
rect 591102 693538 591658 694094
rect 591102 657538 591658 658094
rect 591102 621538 591658 622094
rect 591102 585538 591658 586094
rect 591102 549538 591658 550094
rect 591102 513538 591658 514094
rect 591102 477538 591658 478094
rect 591102 441538 591658 442094
rect 591102 405538 591658 406094
rect 591102 369538 591658 370094
rect 591102 333538 591658 334094
rect 591102 297538 591658 298094
rect 591102 261538 591658 262094
rect 591102 225538 591658 226094
rect 591102 189538 591658 190094
rect 591102 153538 591658 154094
rect 591102 117538 591658 118094
rect 591102 81538 591658 82094
rect 591102 45538 591658 46094
rect 591102 9538 591658 10094
rect 591102 -6662 591658 -6106
rect 592062 694778 592618 695334
rect 592062 658778 592618 659334
rect 592062 622778 592618 623334
rect 592062 586778 592618 587334
rect 592062 550778 592618 551334
rect 592062 514778 592618 515334
rect 592062 478778 592618 479334
rect 592062 442778 592618 443334
rect 592062 406778 592618 407334
rect 592062 370778 592618 371334
rect 592062 334778 592618 335334
rect 592062 298778 592618 299334
rect 592062 262778 592618 263334
rect 592062 226778 592618 227334
rect 592062 190778 592618 191334
rect 592062 154778 592618 155334
rect 592062 118778 592618 119334
rect 592062 82778 592618 83334
rect 592062 46778 592618 47334
rect 592062 10778 592618 11334
rect 592062 -7622 592618 -7066
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711002 -8694 711558
rect -8138 711002 9706 711558
rect 10262 711002 45706 711558
rect 46262 711002 81706 711558
rect 82262 711002 117706 711558
rect 118262 711002 153706 711558
rect 154262 711002 189706 711558
rect 190262 711002 225706 711558
rect 226262 711002 261706 711558
rect 262262 711002 297706 711558
rect 298262 711002 333706 711558
rect 334262 711002 369706 711558
rect 370262 711002 405706 711558
rect 406262 711002 441706 711558
rect 442262 711002 477706 711558
rect 478262 711002 513706 711558
rect 514262 711002 549706 711558
rect 550262 711002 592062 711558
rect 592618 711002 592650 711558
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710042 -7734 710598
rect -7178 710042 8466 710598
rect 9022 710042 44466 710598
rect 45022 710042 80466 710598
rect 81022 710042 116466 710598
rect 117022 710042 152466 710598
rect 153022 710042 188466 710598
rect 189022 710042 224466 710598
rect 225022 710042 260466 710598
rect 261022 710042 296466 710598
rect 297022 710042 332466 710598
rect 333022 710042 368466 710598
rect 369022 710042 404466 710598
rect 405022 710042 440466 710598
rect 441022 710042 476466 710598
rect 477022 710042 512466 710598
rect 513022 710042 548466 710598
rect 549022 710042 591102 710598
rect 591658 710042 591690 710598
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709082 -6774 709638
rect -6218 709082 7226 709638
rect 7782 709082 43226 709638
rect 43782 709082 79226 709638
rect 79782 709082 115226 709638
rect 115782 709082 151226 709638
rect 151782 709082 187226 709638
rect 187782 709082 223226 709638
rect 223782 709082 259226 709638
rect 259782 709082 295226 709638
rect 295782 709082 331226 709638
rect 331782 709082 367226 709638
rect 367782 709082 403226 709638
rect 403782 709082 439226 709638
rect 439782 709082 475226 709638
rect 475782 709082 511226 709638
rect 511782 709082 547226 709638
rect 547782 709082 590142 709638
rect 590698 709082 590730 709638
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708122 -5814 708678
rect -5258 708122 5986 708678
rect 6542 708122 41986 708678
rect 42542 708122 77986 708678
rect 78542 708122 113986 708678
rect 114542 708122 149986 708678
rect 150542 708122 185986 708678
rect 186542 708122 221986 708678
rect 222542 708122 257986 708678
rect 258542 708122 293986 708678
rect 294542 708122 329986 708678
rect 330542 708122 365986 708678
rect 366542 708122 401986 708678
rect 402542 708122 437986 708678
rect 438542 708122 473986 708678
rect 474542 708122 509986 708678
rect 510542 708122 545986 708678
rect 546542 708122 581986 708678
rect 582542 708122 589182 708678
rect 589738 708122 589770 708678
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707162 -4854 707718
rect -4298 707162 4746 707718
rect 5302 707162 40746 707718
rect 41302 707162 76746 707718
rect 77302 707162 112746 707718
rect 113302 707162 148746 707718
rect 149302 707162 184746 707718
rect 185302 707162 220746 707718
rect 221302 707162 256746 707718
rect 257302 707162 292746 707718
rect 293302 707162 328746 707718
rect 329302 707162 364746 707718
rect 365302 707162 400746 707718
rect 401302 707162 436746 707718
rect 437302 707162 472746 707718
rect 473302 707162 508746 707718
rect 509302 707162 544746 707718
rect 545302 707162 580746 707718
rect 581302 707162 588222 707718
rect 588778 707162 588810 707718
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706202 -3894 706758
rect -3338 706202 3506 706758
rect 4062 706202 39506 706758
rect 40062 706202 75506 706758
rect 76062 706202 111506 706758
rect 112062 706202 147506 706758
rect 148062 706202 183506 706758
rect 184062 706202 219506 706758
rect 220062 706202 255506 706758
rect 256062 706202 291506 706758
rect 292062 706202 327506 706758
rect 328062 706202 363506 706758
rect 364062 706202 399506 706758
rect 400062 706202 435506 706758
rect 436062 706202 471506 706758
rect 472062 706202 507506 706758
rect 508062 706202 543506 706758
rect 544062 706202 579506 706758
rect 580062 706202 587262 706758
rect 587818 706202 587850 706758
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705242 -2934 705798
rect -2378 705242 2266 705798
rect 2822 705242 38266 705798
rect 38822 705242 74266 705798
rect 74822 705242 110266 705798
rect 110822 705242 146266 705798
rect 146822 705242 182266 705798
rect 182822 705242 218266 705798
rect 218822 705242 254266 705798
rect 254822 705242 290266 705798
rect 290822 705242 326266 705798
rect 326822 705242 362266 705798
rect 362822 705242 398266 705798
rect 398822 705242 434266 705798
rect 434822 705242 470266 705798
rect 470822 705242 506266 705798
rect 506822 705242 542266 705798
rect 542822 705242 578266 705798
rect 578822 705242 586302 705798
rect 586858 705242 586890 705798
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704282 -1974 704838
rect -1418 704282 1026 704838
rect 1582 704282 37026 704838
rect 37582 704282 73026 704838
rect 73582 704282 109026 704838
rect 109582 704282 145026 704838
rect 145582 704282 181026 704838
rect 181582 704282 217026 704838
rect 217582 704282 253026 704838
rect 253582 704282 289026 704838
rect 289582 704282 325026 704838
rect 325582 704282 361026 704838
rect 361582 704282 397026 704838
rect 397582 704282 433026 704838
rect 433582 704282 469026 704838
rect 469582 704282 505026 704838
rect 505582 704282 541026 704838
rect 541582 704282 577026 704838
rect 577582 704282 585342 704838
rect 585898 704282 585930 704838
rect -2006 704250 585930 704282
rect -8726 695334 592650 695366
rect -8726 694778 -8694 695334
rect -8138 694778 9706 695334
rect 10262 694778 45706 695334
rect 46262 694778 81706 695334
rect 82262 694778 117706 695334
rect 118262 694778 153706 695334
rect 154262 694778 189706 695334
rect 190262 694778 225706 695334
rect 226262 694778 261706 695334
rect 262262 694778 297706 695334
rect 298262 694778 333706 695334
rect 334262 694778 369706 695334
rect 370262 694778 405706 695334
rect 406262 694778 441706 695334
rect 442262 694778 477706 695334
rect 478262 694778 513706 695334
rect 514262 694778 549706 695334
rect 550262 694778 592062 695334
rect 592618 694778 592650 695334
rect -8726 694746 592650 694778
rect -8726 694094 592650 694126
rect -8726 693538 -7734 694094
rect -7178 693538 8466 694094
rect 9022 693538 44466 694094
rect 45022 693538 80466 694094
rect 81022 693538 116466 694094
rect 117022 693538 152466 694094
rect 153022 693538 188466 694094
rect 189022 693538 224466 694094
rect 225022 693538 260466 694094
rect 261022 693538 296466 694094
rect 297022 693538 332466 694094
rect 333022 693538 368466 694094
rect 369022 693538 404466 694094
rect 405022 693538 440466 694094
rect 441022 693538 476466 694094
rect 477022 693538 512466 694094
rect 513022 693538 548466 694094
rect 549022 693538 591102 694094
rect 591658 693538 592650 694094
rect -8726 693506 592650 693538
rect -8726 692854 592650 692886
rect -8726 692298 -6774 692854
rect -6218 692298 7226 692854
rect 7782 692298 43226 692854
rect 43782 692298 79226 692854
rect 79782 692298 115226 692854
rect 115782 692298 151226 692854
rect 151782 692298 187226 692854
rect 187782 692298 223226 692854
rect 223782 692298 259226 692854
rect 259782 692298 295226 692854
rect 295782 692298 331226 692854
rect 331782 692298 367226 692854
rect 367782 692298 403226 692854
rect 403782 692298 439226 692854
rect 439782 692298 475226 692854
rect 475782 692298 511226 692854
rect 511782 692298 547226 692854
rect 547782 692298 590142 692854
rect 590698 692298 592650 692854
rect -8726 692266 592650 692298
rect -8726 691614 592650 691646
rect -8726 691058 -5814 691614
rect -5258 691058 5986 691614
rect 6542 691058 41986 691614
rect 42542 691058 77986 691614
rect 78542 691058 113986 691614
rect 114542 691058 149986 691614
rect 150542 691058 185986 691614
rect 186542 691058 221986 691614
rect 222542 691058 257986 691614
rect 258542 691058 293986 691614
rect 294542 691058 329986 691614
rect 330542 691058 365986 691614
rect 366542 691058 401986 691614
rect 402542 691058 437986 691614
rect 438542 691058 473986 691614
rect 474542 691058 509986 691614
rect 510542 691058 545986 691614
rect 546542 691058 581986 691614
rect 582542 691058 589182 691614
rect 589738 691058 592650 691614
rect -8726 691026 592650 691058
rect -8726 690374 592650 690406
rect -8726 689818 -4854 690374
rect -4298 689818 4746 690374
rect 5302 689818 40746 690374
rect 41302 689818 76746 690374
rect 77302 689818 112746 690374
rect 113302 689818 148746 690374
rect 149302 689818 184746 690374
rect 185302 689818 220746 690374
rect 221302 689818 256746 690374
rect 257302 689818 292746 690374
rect 293302 689818 328746 690374
rect 329302 689818 364746 690374
rect 365302 689818 400746 690374
rect 401302 689818 436746 690374
rect 437302 689818 472746 690374
rect 473302 689818 508746 690374
rect 509302 689818 544746 690374
rect 545302 689818 580746 690374
rect 581302 689818 588222 690374
rect 588778 689818 592650 690374
rect -8726 689786 592650 689818
rect -8726 689134 592650 689166
rect -8726 688578 -3894 689134
rect -3338 688578 3506 689134
rect 4062 688578 39506 689134
rect 40062 688578 75506 689134
rect 76062 688578 111506 689134
rect 112062 688578 147506 689134
rect 148062 688578 183506 689134
rect 184062 688578 219506 689134
rect 220062 688578 255506 689134
rect 256062 688578 291506 689134
rect 292062 688578 327506 689134
rect 328062 688578 363506 689134
rect 364062 688578 399506 689134
rect 400062 688578 435506 689134
rect 436062 688578 471506 689134
rect 472062 688578 507506 689134
rect 508062 688578 543506 689134
rect 544062 688578 579506 689134
rect 580062 688578 587262 689134
rect 587818 688578 592650 689134
rect -8726 688546 592650 688578
rect -8726 687894 592650 687926
rect -8726 687338 -2934 687894
rect -2378 687338 2266 687894
rect 2822 687338 38266 687894
rect 38822 687338 74266 687894
rect 74822 687338 110266 687894
rect 110822 687338 146266 687894
rect 146822 687338 182266 687894
rect 182822 687338 218266 687894
rect 218822 687338 254266 687894
rect 254822 687338 290266 687894
rect 290822 687338 326266 687894
rect 326822 687338 362266 687894
rect 362822 687338 398266 687894
rect 398822 687338 434266 687894
rect 434822 687338 470266 687894
rect 470822 687338 506266 687894
rect 506822 687338 542266 687894
rect 542822 687338 578266 687894
rect 578822 687338 586302 687894
rect 586858 687338 592650 687894
rect -8726 687306 592650 687338
rect -8726 686654 592650 686686
rect -8726 686098 -1974 686654
rect -1418 686098 1026 686654
rect 1582 686098 37026 686654
rect 37582 686098 73026 686654
rect 73582 686098 109026 686654
rect 109582 686098 145026 686654
rect 145582 686098 181026 686654
rect 181582 686098 217026 686654
rect 217582 686098 253026 686654
rect 253582 686098 289026 686654
rect 289582 686098 325026 686654
rect 325582 686098 361026 686654
rect 361582 686098 397026 686654
rect 397582 686098 433026 686654
rect 433582 686098 469026 686654
rect 469582 686098 505026 686654
rect 505582 686098 541026 686654
rect 541582 686098 577026 686654
rect 577582 686098 585342 686654
rect 585898 686098 592650 686654
rect -8726 686066 592650 686098
rect -8726 659334 592650 659366
rect -8726 658778 -8694 659334
rect -8138 658778 9706 659334
rect 10262 658778 45706 659334
rect 46262 658778 81706 659334
rect 82262 658778 117706 659334
rect 118262 658778 153706 659334
rect 154262 658778 189706 659334
rect 190262 658778 225706 659334
rect 226262 658778 261706 659334
rect 262262 658778 297706 659334
rect 298262 658778 333706 659334
rect 334262 658778 369706 659334
rect 370262 658778 405706 659334
rect 406262 658778 441706 659334
rect 442262 658778 477706 659334
rect 478262 658778 513706 659334
rect 514262 658778 549706 659334
rect 550262 658778 592062 659334
rect 592618 658778 592650 659334
rect -8726 658746 592650 658778
rect -8726 658094 592650 658126
rect -8726 657538 -7734 658094
rect -7178 657538 8466 658094
rect 9022 657538 44466 658094
rect 45022 657538 80466 658094
rect 81022 657538 116466 658094
rect 117022 657538 152466 658094
rect 153022 657538 188466 658094
rect 189022 657538 224466 658094
rect 225022 657538 260466 658094
rect 261022 657538 296466 658094
rect 297022 657538 332466 658094
rect 333022 657538 368466 658094
rect 369022 657538 404466 658094
rect 405022 657538 440466 658094
rect 441022 657538 476466 658094
rect 477022 657538 512466 658094
rect 513022 657538 548466 658094
rect 549022 657538 591102 658094
rect 591658 657538 592650 658094
rect -8726 657506 592650 657538
rect -8726 656854 592650 656886
rect -8726 656298 -6774 656854
rect -6218 656298 7226 656854
rect 7782 656298 43226 656854
rect 43782 656298 79226 656854
rect 79782 656298 115226 656854
rect 115782 656298 151226 656854
rect 151782 656298 187226 656854
rect 187782 656298 223226 656854
rect 223782 656298 259226 656854
rect 259782 656298 295226 656854
rect 295782 656298 331226 656854
rect 331782 656298 367226 656854
rect 367782 656298 403226 656854
rect 403782 656298 439226 656854
rect 439782 656298 475226 656854
rect 475782 656298 511226 656854
rect 511782 656298 547226 656854
rect 547782 656298 590142 656854
rect 590698 656298 592650 656854
rect -8726 656266 592650 656298
rect -8726 655614 592650 655646
rect -8726 655058 -5814 655614
rect -5258 655058 5986 655614
rect 6542 655058 41986 655614
rect 42542 655058 77986 655614
rect 78542 655058 113986 655614
rect 114542 655058 149986 655614
rect 150542 655058 185986 655614
rect 186542 655058 221986 655614
rect 222542 655058 257986 655614
rect 258542 655058 293986 655614
rect 294542 655058 329986 655614
rect 330542 655058 365986 655614
rect 366542 655058 401986 655614
rect 402542 655058 437986 655614
rect 438542 655058 473986 655614
rect 474542 655058 509986 655614
rect 510542 655058 545986 655614
rect 546542 655058 581986 655614
rect 582542 655058 589182 655614
rect 589738 655058 592650 655614
rect -8726 655026 592650 655058
rect -8726 654374 592650 654406
rect -8726 653818 -4854 654374
rect -4298 653818 4746 654374
rect 5302 653818 40746 654374
rect 41302 653818 76746 654374
rect 77302 653818 112746 654374
rect 113302 653818 148746 654374
rect 149302 653818 184746 654374
rect 185302 653818 220746 654374
rect 221302 653818 256746 654374
rect 257302 653818 292746 654374
rect 293302 653818 328746 654374
rect 329302 653818 364746 654374
rect 365302 653818 400746 654374
rect 401302 653818 436746 654374
rect 437302 653818 472746 654374
rect 473302 653818 508746 654374
rect 509302 653818 544746 654374
rect 545302 653818 580746 654374
rect 581302 653818 588222 654374
rect 588778 653818 592650 654374
rect -8726 653786 592650 653818
rect -8726 653134 592650 653166
rect -8726 652578 -3894 653134
rect -3338 652578 3506 653134
rect 4062 652578 39506 653134
rect 40062 652578 75506 653134
rect 76062 652578 111506 653134
rect 112062 652578 147506 653134
rect 148062 652578 183506 653134
rect 184062 652578 219506 653134
rect 220062 652578 255506 653134
rect 256062 652578 291506 653134
rect 292062 652578 327506 653134
rect 328062 652578 363506 653134
rect 364062 652578 399506 653134
rect 400062 652578 435506 653134
rect 436062 652578 471506 653134
rect 472062 652578 507506 653134
rect 508062 652578 543506 653134
rect 544062 652578 579506 653134
rect 580062 652578 587262 653134
rect 587818 652578 592650 653134
rect -8726 652546 592650 652578
rect -8726 651894 592650 651926
rect -8726 651338 -2934 651894
rect -2378 651338 2266 651894
rect 2822 651338 38266 651894
rect 38822 651338 74266 651894
rect 74822 651338 110266 651894
rect 110822 651338 146266 651894
rect 146822 651338 182266 651894
rect 182822 651338 218266 651894
rect 218822 651338 254266 651894
rect 254822 651338 290266 651894
rect 290822 651338 326266 651894
rect 326822 651338 362266 651894
rect 362822 651338 398266 651894
rect 398822 651338 434266 651894
rect 434822 651338 470266 651894
rect 470822 651338 506266 651894
rect 506822 651338 542266 651894
rect 542822 651338 578266 651894
rect 578822 651338 586302 651894
rect 586858 651338 592650 651894
rect -8726 651306 592650 651338
rect -8726 650654 592650 650686
rect -8726 650098 -1974 650654
rect -1418 650098 1026 650654
rect 1582 650098 37026 650654
rect 37582 650098 73026 650654
rect 73582 650098 109026 650654
rect 109582 650098 145026 650654
rect 145582 650098 181026 650654
rect 181582 650098 217026 650654
rect 217582 650098 253026 650654
rect 253582 650098 289026 650654
rect 289582 650098 325026 650654
rect 325582 650098 361026 650654
rect 361582 650098 397026 650654
rect 397582 650098 433026 650654
rect 433582 650098 469026 650654
rect 469582 650098 505026 650654
rect 505582 650098 541026 650654
rect 541582 650098 577026 650654
rect 577582 650098 585342 650654
rect 585898 650098 592650 650654
rect -8726 650066 592650 650098
rect -8726 623334 592650 623366
rect -8726 622778 -8694 623334
rect -8138 622778 9706 623334
rect 10262 622778 45706 623334
rect 46262 622778 81706 623334
rect 82262 622778 117706 623334
rect 118262 622778 153706 623334
rect 154262 622778 189706 623334
rect 190262 622778 225706 623334
rect 226262 622778 261706 623334
rect 262262 622778 297706 623334
rect 298262 622778 333706 623334
rect 334262 622778 369706 623334
rect 370262 622778 405706 623334
rect 406262 622778 441706 623334
rect 442262 622778 477706 623334
rect 478262 622778 513706 623334
rect 514262 622778 549706 623334
rect 550262 622778 592062 623334
rect 592618 622778 592650 623334
rect -8726 622746 592650 622778
rect -8726 622094 592650 622126
rect -8726 621538 -7734 622094
rect -7178 621538 8466 622094
rect 9022 621538 44466 622094
rect 45022 621538 80466 622094
rect 81022 621538 116466 622094
rect 117022 621538 152466 622094
rect 153022 621538 188466 622094
rect 189022 621538 224466 622094
rect 225022 621538 260466 622094
rect 261022 621538 296466 622094
rect 297022 621538 332466 622094
rect 333022 621538 368466 622094
rect 369022 621538 404466 622094
rect 405022 621538 440466 622094
rect 441022 621538 476466 622094
rect 477022 621538 512466 622094
rect 513022 621538 548466 622094
rect 549022 621538 591102 622094
rect 591658 621538 592650 622094
rect -8726 621506 592650 621538
rect -8726 620854 592650 620886
rect -8726 620298 -6774 620854
rect -6218 620298 7226 620854
rect 7782 620298 43226 620854
rect 43782 620298 79226 620854
rect 79782 620298 115226 620854
rect 115782 620298 151226 620854
rect 151782 620298 187226 620854
rect 187782 620298 223226 620854
rect 223782 620298 259226 620854
rect 259782 620298 295226 620854
rect 295782 620298 331226 620854
rect 331782 620298 367226 620854
rect 367782 620298 403226 620854
rect 403782 620298 439226 620854
rect 439782 620298 475226 620854
rect 475782 620298 511226 620854
rect 511782 620298 547226 620854
rect 547782 620298 590142 620854
rect 590698 620298 592650 620854
rect -8726 620266 592650 620298
rect -8726 619614 592650 619646
rect -8726 619058 -5814 619614
rect -5258 619058 5986 619614
rect 6542 619058 41986 619614
rect 42542 619058 77986 619614
rect 78542 619058 113986 619614
rect 114542 619058 149986 619614
rect 150542 619058 185986 619614
rect 186542 619058 221986 619614
rect 222542 619058 257986 619614
rect 258542 619058 293986 619614
rect 294542 619058 329986 619614
rect 330542 619058 365986 619614
rect 366542 619058 401986 619614
rect 402542 619058 437986 619614
rect 438542 619058 473986 619614
rect 474542 619058 509986 619614
rect 510542 619058 545986 619614
rect 546542 619058 581986 619614
rect 582542 619058 589182 619614
rect 589738 619058 592650 619614
rect -8726 619026 592650 619058
rect -8726 618374 592650 618406
rect -8726 617818 -4854 618374
rect -4298 617818 4746 618374
rect 5302 617818 40746 618374
rect 41302 617818 76746 618374
rect 77302 617818 112746 618374
rect 113302 617818 148746 618374
rect 149302 617818 184746 618374
rect 185302 617818 220746 618374
rect 221302 617818 256746 618374
rect 257302 617818 292746 618374
rect 293302 617818 328746 618374
rect 329302 617818 364746 618374
rect 365302 617818 400746 618374
rect 401302 617818 436746 618374
rect 437302 617818 472746 618374
rect 473302 617818 508746 618374
rect 509302 617818 544746 618374
rect 545302 617818 580746 618374
rect 581302 617818 588222 618374
rect 588778 617818 592650 618374
rect -8726 617786 592650 617818
rect -8726 617134 592650 617166
rect -8726 616578 -3894 617134
rect -3338 616578 3506 617134
rect 4062 616578 39506 617134
rect 40062 616578 75506 617134
rect 76062 616578 111506 617134
rect 112062 616578 147506 617134
rect 148062 616578 183506 617134
rect 184062 616578 219506 617134
rect 220062 616578 255506 617134
rect 256062 616578 291506 617134
rect 292062 616578 327506 617134
rect 328062 616578 363506 617134
rect 364062 616578 399506 617134
rect 400062 616578 435506 617134
rect 436062 616578 471506 617134
rect 472062 616578 507506 617134
rect 508062 616578 543506 617134
rect 544062 616578 579506 617134
rect 580062 616578 587262 617134
rect 587818 616578 592650 617134
rect -8726 616546 592650 616578
rect -8726 615894 592650 615926
rect -8726 615338 -2934 615894
rect -2378 615338 2266 615894
rect 2822 615338 38266 615894
rect 38822 615338 74266 615894
rect 74822 615338 110266 615894
rect 110822 615338 146266 615894
rect 146822 615338 182266 615894
rect 182822 615338 218266 615894
rect 218822 615338 254266 615894
rect 254822 615338 290266 615894
rect 290822 615338 326266 615894
rect 326822 615338 362266 615894
rect 362822 615338 398266 615894
rect 398822 615338 434266 615894
rect 434822 615338 470266 615894
rect 470822 615338 506266 615894
rect 506822 615338 542266 615894
rect 542822 615338 578266 615894
rect 578822 615338 586302 615894
rect 586858 615338 592650 615894
rect -8726 615306 592650 615338
rect -8726 614654 592650 614686
rect -8726 614098 -1974 614654
rect -1418 614098 1026 614654
rect 1582 614098 37026 614654
rect 37582 614098 73026 614654
rect 73582 614098 109026 614654
rect 109582 614098 145026 614654
rect 145582 614098 181026 614654
rect 181582 614098 217026 614654
rect 217582 614098 253026 614654
rect 253582 614098 289026 614654
rect 289582 614098 325026 614654
rect 325582 614098 361026 614654
rect 361582 614098 397026 614654
rect 397582 614098 433026 614654
rect 433582 614098 469026 614654
rect 469582 614098 505026 614654
rect 505582 614098 541026 614654
rect 541582 614098 577026 614654
rect 577582 614098 585342 614654
rect 585898 614098 592650 614654
rect -8726 614066 592650 614098
rect -8726 587334 592650 587366
rect -8726 586778 -8694 587334
rect -8138 586778 9706 587334
rect 10262 586778 45706 587334
rect 46262 586778 81706 587334
rect 82262 586778 117706 587334
rect 118262 586778 153706 587334
rect 154262 586778 189706 587334
rect 190262 586778 225706 587334
rect 226262 586778 261706 587334
rect 262262 586778 297706 587334
rect 298262 586778 333706 587334
rect 334262 586778 369706 587334
rect 370262 586778 405706 587334
rect 406262 586778 441706 587334
rect 442262 586778 477706 587334
rect 478262 586778 513706 587334
rect 514262 586778 549706 587334
rect 550262 586778 592062 587334
rect 592618 586778 592650 587334
rect -8726 586746 592650 586778
rect -8726 586094 592650 586126
rect -8726 585538 -7734 586094
rect -7178 585538 8466 586094
rect 9022 585538 44466 586094
rect 45022 585538 80466 586094
rect 81022 585538 116466 586094
rect 117022 585538 152466 586094
rect 153022 585538 188466 586094
rect 189022 585538 224466 586094
rect 225022 585538 260466 586094
rect 261022 585538 296466 586094
rect 297022 585538 332466 586094
rect 333022 585538 368466 586094
rect 369022 585538 404466 586094
rect 405022 585538 440466 586094
rect 441022 585538 476466 586094
rect 477022 585538 512466 586094
rect 513022 585538 548466 586094
rect 549022 585538 591102 586094
rect 591658 585538 592650 586094
rect -8726 585506 592650 585538
rect -8726 584854 592650 584886
rect -8726 584298 -6774 584854
rect -6218 584298 7226 584854
rect 7782 584298 43226 584854
rect 43782 584298 79226 584854
rect 79782 584298 115226 584854
rect 115782 584298 151226 584854
rect 151782 584298 187226 584854
rect 187782 584298 223226 584854
rect 223782 584298 259226 584854
rect 259782 584298 295226 584854
rect 295782 584298 331226 584854
rect 331782 584298 367226 584854
rect 367782 584298 403226 584854
rect 403782 584298 439226 584854
rect 439782 584298 475226 584854
rect 475782 584298 511226 584854
rect 511782 584298 547226 584854
rect 547782 584298 590142 584854
rect 590698 584298 592650 584854
rect -8726 584266 592650 584298
rect -8726 583614 592650 583646
rect -8726 583058 -5814 583614
rect -5258 583058 5986 583614
rect 6542 583058 41986 583614
rect 42542 583058 77986 583614
rect 78542 583058 113986 583614
rect 114542 583058 149986 583614
rect 150542 583058 185986 583614
rect 186542 583058 221986 583614
rect 222542 583058 257986 583614
rect 258542 583058 293986 583614
rect 294542 583058 329986 583614
rect 330542 583058 365986 583614
rect 366542 583058 401986 583614
rect 402542 583058 437986 583614
rect 438542 583058 473986 583614
rect 474542 583058 509986 583614
rect 510542 583058 545986 583614
rect 546542 583058 581986 583614
rect 582542 583058 589182 583614
rect 589738 583058 592650 583614
rect -8726 583026 592650 583058
rect -8726 582374 592650 582406
rect -8726 581818 -4854 582374
rect -4298 581818 4746 582374
rect 5302 581818 40746 582374
rect 41302 581818 76746 582374
rect 77302 581818 112746 582374
rect 113302 581818 148746 582374
rect 149302 581818 184746 582374
rect 185302 581818 220746 582374
rect 221302 581818 256746 582374
rect 257302 581818 292746 582374
rect 293302 581818 328746 582374
rect 329302 581818 364746 582374
rect 365302 581818 400746 582374
rect 401302 581818 436746 582374
rect 437302 581818 472746 582374
rect 473302 581818 508746 582374
rect 509302 581818 544746 582374
rect 545302 581818 580746 582374
rect 581302 581818 588222 582374
rect 588778 581818 592650 582374
rect -8726 581786 592650 581818
rect -8726 581134 592650 581166
rect -8726 580578 -3894 581134
rect -3338 580578 3506 581134
rect 4062 580578 39506 581134
rect 40062 580578 75506 581134
rect 76062 580578 111506 581134
rect 112062 580578 147506 581134
rect 148062 580578 183506 581134
rect 184062 580578 219506 581134
rect 220062 580578 255506 581134
rect 256062 580578 291506 581134
rect 292062 580578 327506 581134
rect 328062 580578 363506 581134
rect 364062 580578 399506 581134
rect 400062 580578 435506 581134
rect 436062 580578 471506 581134
rect 472062 580578 507506 581134
rect 508062 580578 543506 581134
rect 544062 580578 579506 581134
rect 580062 580578 587262 581134
rect 587818 580578 592650 581134
rect -8726 580546 592650 580578
rect -8726 579894 592650 579926
rect -8726 579338 -2934 579894
rect -2378 579338 2266 579894
rect 2822 579338 38266 579894
rect 38822 579338 74266 579894
rect 74822 579338 110266 579894
rect 110822 579338 146266 579894
rect 146822 579338 182266 579894
rect 182822 579338 218266 579894
rect 218822 579338 254266 579894
rect 254822 579338 290266 579894
rect 290822 579338 326266 579894
rect 326822 579338 362266 579894
rect 362822 579338 398266 579894
rect 398822 579338 434266 579894
rect 434822 579338 470266 579894
rect 470822 579338 506266 579894
rect 506822 579338 542266 579894
rect 542822 579338 578266 579894
rect 578822 579338 586302 579894
rect 586858 579338 592650 579894
rect -8726 579306 592650 579338
rect -8726 578654 592650 578686
rect -8726 578098 -1974 578654
rect -1418 578098 1026 578654
rect 1582 578098 37026 578654
rect 37582 578098 73026 578654
rect 73582 578098 109026 578654
rect 109582 578098 145026 578654
rect 145582 578098 181026 578654
rect 181582 578098 217026 578654
rect 217582 578098 253026 578654
rect 253582 578098 289026 578654
rect 289582 578098 325026 578654
rect 325582 578098 361026 578654
rect 361582 578098 397026 578654
rect 397582 578098 433026 578654
rect 433582 578098 469026 578654
rect 469582 578098 505026 578654
rect 505582 578098 541026 578654
rect 541582 578098 577026 578654
rect 577582 578098 585342 578654
rect 585898 578098 592650 578654
rect -8726 578066 592650 578098
rect -8726 551334 592650 551366
rect -8726 550778 -8694 551334
rect -8138 550778 9706 551334
rect 10262 550778 45706 551334
rect 46262 550778 81706 551334
rect 82262 550778 117706 551334
rect 118262 550778 153706 551334
rect 154262 550778 189706 551334
rect 190262 550778 225706 551334
rect 226262 550778 261706 551334
rect 262262 550778 297706 551334
rect 298262 550778 333706 551334
rect 334262 550778 369706 551334
rect 370262 550778 405706 551334
rect 406262 550778 441706 551334
rect 442262 550778 477706 551334
rect 478262 550778 513706 551334
rect 514262 550778 549706 551334
rect 550262 550778 592062 551334
rect 592618 550778 592650 551334
rect -8726 550746 592650 550778
rect -8726 550094 592650 550126
rect -8726 549538 -7734 550094
rect -7178 549538 8466 550094
rect 9022 549538 44466 550094
rect 45022 549538 80466 550094
rect 81022 549538 116466 550094
rect 117022 549538 152466 550094
rect 153022 549538 188466 550094
rect 189022 549538 224466 550094
rect 225022 549538 260466 550094
rect 261022 549538 296466 550094
rect 297022 549538 332466 550094
rect 333022 549538 368466 550094
rect 369022 549538 404466 550094
rect 405022 549538 440466 550094
rect 441022 549538 476466 550094
rect 477022 549538 512466 550094
rect 513022 549538 548466 550094
rect 549022 549538 591102 550094
rect 591658 549538 592650 550094
rect -8726 549506 592650 549538
rect -8726 548854 592650 548886
rect -8726 548298 -6774 548854
rect -6218 548298 7226 548854
rect 7782 548298 43226 548854
rect 43782 548298 79226 548854
rect 79782 548298 115226 548854
rect 115782 548298 151226 548854
rect 151782 548298 187226 548854
rect 187782 548298 223226 548854
rect 223782 548298 259226 548854
rect 259782 548298 295226 548854
rect 295782 548298 331226 548854
rect 331782 548298 367226 548854
rect 367782 548298 403226 548854
rect 403782 548298 439226 548854
rect 439782 548298 475226 548854
rect 475782 548298 511226 548854
rect 511782 548298 547226 548854
rect 547782 548298 590142 548854
rect 590698 548298 592650 548854
rect -8726 548266 592650 548298
rect -8726 547614 592650 547646
rect -8726 547058 -5814 547614
rect -5258 547058 5986 547614
rect 6542 547058 41986 547614
rect 42542 547058 77986 547614
rect 78542 547058 113986 547614
rect 114542 547058 149986 547614
rect 150542 547058 185986 547614
rect 186542 547058 221986 547614
rect 222542 547058 257986 547614
rect 258542 547058 293986 547614
rect 294542 547058 329986 547614
rect 330542 547058 365986 547614
rect 366542 547058 401986 547614
rect 402542 547058 437986 547614
rect 438542 547058 473986 547614
rect 474542 547058 509986 547614
rect 510542 547058 545986 547614
rect 546542 547058 581986 547614
rect 582542 547058 589182 547614
rect 589738 547058 592650 547614
rect -8726 547026 592650 547058
rect -8726 546374 592650 546406
rect -8726 545818 -4854 546374
rect -4298 545818 4746 546374
rect 5302 545818 40746 546374
rect 41302 545818 76746 546374
rect 77302 545818 112746 546374
rect 113302 545818 148746 546374
rect 149302 545818 184746 546374
rect 185302 545818 220746 546374
rect 221302 545818 256746 546374
rect 257302 545818 292746 546374
rect 293302 545818 328746 546374
rect 329302 545818 364746 546374
rect 365302 545818 400746 546374
rect 401302 545818 436746 546374
rect 437302 545818 472746 546374
rect 473302 545818 508746 546374
rect 509302 545818 544746 546374
rect 545302 545818 580746 546374
rect 581302 545818 588222 546374
rect 588778 545818 592650 546374
rect -8726 545786 592650 545818
rect -8726 545134 592650 545166
rect -8726 544578 -3894 545134
rect -3338 544578 3506 545134
rect 4062 544578 39506 545134
rect 40062 544578 75506 545134
rect 76062 544578 111506 545134
rect 112062 544578 147506 545134
rect 148062 544578 183506 545134
rect 184062 544578 219506 545134
rect 220062 544578 255506 545134
rect 256062 544578 291506 545134
rect 292062 544578 327506 545134
rect 328062 544578 363506 545134
rect 364062 544578 399506 545134
rect 400062 544578 435506 545134
rect 436062 544578 471506 545134
rect 472062 544578 507506 545134
rect 508062 544578 543506 545134
rect 544062 544578 579506 545134
rect 580062 544578 587262 545134
rect 587818 544578 592650 545134
rect -8726 544546 592650 544578
rect -8726 543894 592650 543926
rect -8726 543338 -2934 543894
rect -2378 543338 2266 543894
rect 2822 543338 38266 543894
rect 38822 543338 74266 543894
rect 74822 543338 110266 543894
rect 110822 543338 146266 543894
rect 146822 543338 182266 543894
rect 182822 543338 218266 543894
rect 218822 543338 254266 543894
rect 254822 543338 290266 543894
rect 290822 543338 326266 543894
rect 326822 543338 362266 543894
rect 362822 543338 398266 543894
rect 398822 543338 434266 543894
rect 434822 543338 470266 543894
rect 470822 543338 506266 543894
rect 506822 543338 542266 543894
rect 542822 543338 578266 543894
rect 578822 543338 586302 543894
rect 586858 543338 592650 543894
rect -8726 543306 592650 543338
rect -8726 542654 592650 542686
rect -8726 542098 -1974 542654
rect -1418 542098 1026 542654
rect 1582 542098 37026 542654
rect 37582 542098 73026 542654
rect 73582 542098 109026 542654
rect 109582 542098 145026 542654
rect 145582 542098 181026 542654
rect 181582 542098 217026 542654
rect 217582 542098 253026 542654
rect 253582 542098 289026 542654
rect 289582 542098 325026 542654
rect 325582 542098 361026 542654
rect 361582 542098 397026 542654
rect 397582 542098 433026 542654
rect 433582 542098 469026 542654
rect 469582 542098 505026 542654
rect 505582 542098 541026 542654
rect 541582 542098 577026 542654
rect 577582 542098 585342 542654
rect 585898 542098 592650 542654
rect -8726 542066 592650 542098
rect -8726 515334 592650 515366
rect -8726 514778 -8694 515334
rect -8138 514778 9706 515334
rect 10262 514778 45706 515334
rect 46262 514778 81706 515334
rect 82262 514778 117706 515334
rect 118262 514778 153706 515334
rect 154262 514778 189706 515334
rect 190262 514778 225706 515334
rect 226262 514778 261706 515334
rect 262262 514778 297706 515334
rect 298262 514778 333706 515334
rect 334262 514778 369706 515334
rect 370262 514778 405706 515334
rect 406262 514778 441706 515334
rect 442262 514778 477706 515334
rect 478262 514778 513706 515334
rect 514262 514778 549706 515334
rect 550262 514778 592062 515334
rect 592618 514778 592650 515334
rect -8726 514746 592650 514778
rect -8726 514094 592650 514126
rect -8726 513538 -7734 514094
rect -7178 513538 8466 514094
rect 9022 513538 44466 514094
rect 45022 513538 80466 514094
rect 81022 513538 116466 514094
rect 117022 513538 152466 514094
rect 153022 513538 188466 514094
rect 189022 513538 224466 514094
rect 225022 513538 260466 514094
rect 261022 513538 296466 514094
rect 297022 513538 332466 514094
rect 333022 513538 368466 514094
rect 369022 513538 404466 514094
rect 405022 513538 440466 514094
rect 441022 513538 476466 514094
rect 477022 513538 512466 514094
rect 513022 513538 548466 514094
rect 549022 513538 591102 514094
rect 591658 513538 592650 514094
rect -8726 513506 592650 513538
rect -8726 512854 592650 512886
rect -8726 512298 -6774 512854
rect -6218 512298 7226 512854
rect 7782 512298 43226 512854
rect 43782 512298 79226 512854
rect 79782 512298 115226 512854
rect 115782 512298 151226 512854
rect 151782 512298 187226 512854
rect 187782 512298 223226 512854
rect 223782 512298 259226 512854
rect 259782 512298 295226 512854
rect 295782 512298 331226 512854
rect 331782 512298 367226 512854
rect 367782 512298 403226 512854
rect 403782 512298 439226 512854
rect 439782 512298 475226 512854
rect 475782 512298 511226 512854
rect 511782 512298 547226 512854
rect 547782 512298 590142 512854
rect 590698 512298 592650 512854
rect -8726 512266 592650 512298
rect -8726 511614 592650 511646
rect -8726 511058 -5814 511614
rect -5258 511058 5986 511614
rect 6542 511058 41986 511614
rect 42542 511058 77986 511614
rect 78542 511058 113986 511614
rect 114542 511058 149986 511614
rect 150542 511058 185986 511614
rect 186542 511058 221986 511614
rect 222542 511058 257986 511614
rect 258542 511058 293986 511614
rect 294542 511058 329986 511614
rect 330542 511058 365986 511614
rect 366542 511058 401986 511614
rect 402542 511058 437986 511614
rect 438542 511058 473986 511614
rect 474542 511058 509986 511614
rect 510542 511058 545986 511614
rect 546542 511058 581986 511614
rect 582542 511058 589182 511614
rect 589738 511058 592650 511614
rect -8726 511026 592650 511058
rect -8726 510374 592650 510406
rect -8726 509818 -4854 510374
rect -4298 509818 4746 510374
rect 5302 509818 40746 510374
rect 41302 509818 76746 510374
rect 77302 509818 112746 510374
rect 113302 509818 148746 510374
rect 149302 509818 184746 510374
rect 185302 509818 220746 510374
rect 221302 509818 256746 510374
rect 257302 509818 292746 510374
rect 293302 509818 328746 510374
rect 329302 509818 364746 510374
rect 365302 509818 400746 510374
rect 401302 509818 436746 510374
rect 437302 509818 472746 510374
rect 473302 509818 508746 510374
rect 509302 509818 544746 510374
rect 545302 509818 580746 510374
rect 581302 509818 588222 510374
rect 588778 509818 592650 510374
rect -8726 509786 592650 509818
rect -8726 509134 592650 509166
rect -8726 508578 -3894 509134
rect -3338 508578 3506 509134
rect 4062 508578 39506 509134
rect 40062 508578 75506 509134
rect 76062 508578 111506 509134
rect 112062 508578 147506 509134
rect 148062 508578 183506 509134
rect 184062 508578 219506 509134
rect 220062 508578 255506 509134
rect 256062 508578 291506 509134
rect 292062 508578 327506 509134
rect 328062 508578 363506 509134
rect 364062 508578 399506 509134
rect 400062 508578 435506 509134
rect 436062 508578 471506 509134
rect 472062 508578 507506 509134
rect 508062 508578 543506 509134
rect 544062 508578 579506 509134
rect 580062 508578 587262 509134
rect 587818 508578 592650 509134
rect -8726 508546 592650 508578
rect -8726 507894 592650 507926
rect -8726 507338 -2934 507894
rect -2378 507338 2266 507894
rect 2822 507338 38266 507894
rect 38822 507338 74266 507894
rect 74822 507338 110266 507894
rect 110822 507338 146266 507894
rect 146822 507338 182266 507894
rect 182822 507338 218266 507894
rect 218822 507338 254266 507894
rect 254822 507338 290266 507894
rect 290822 507338 326266 507894
rect 326822 507338 362266 507894
rect 362822 507338 398266 507894
rect 398822 507338 434266 507894
rect 434822 507338 470266 507894
rect 470822 507338 506266 507894
rect 506822 507338 542266 507894
rect 542822 507338 578266 507894
rect 578822 507338 586302 507894
rect 586858 507338 592650 507894
rect -8726 507306 592650 507338
rect -8726 506654 592650 506686
rect -8726 506098 -1974 506654
rect -1418 506098 1026 506654
rect 1582 506098 37026 506654
rect 37582 506098 73026 506654
rect 73582 506098 109026 506654
rect 109582 506098 145026 506654
rect 145582 506098 181026 506654
rect 181582 506098 217026 506654
rect 217582 506098 253026 506654
rect 253582 506098 289026 506654
rect 289582 506098 325026 506654
rect 325582 506098 361026 506654
rect 361582 506098 397026 506654
rect 397582 506098 433026 506654
rect 433582 506098 469026 506654
rect 469582 506098 505026 506654
rect 505582 506098 541026 506654
rect 541582 506098 577026 506654
rect 577582 506098 585342 506654
rect 585898 506098 592650 506654
rect -8726 506066 592650 506098
rect -8726 479334 592650 479366
rect -8726 478778 -8694 479334
rect -8138 478778 9706 479334
rect 10262 478778 45706 479334
rect 46262 478778 81706 479334
rect 82262 478778 117706 479334
rect 118262 478778 153706 479334
rect 154262 478778 189706 479334
rect 190262 478778 225706 479334
rect 226262 478778 261706 479334
rect 262262 478778 297706 479334
rect 298262 478778 333706 479334
rect 334262 478778 369706 479334
rect 370262 478778 405706 479334
rect 406262 478778 441706 479334
rect 442262 478778 477706 479334
rect 478262 478778 513706 479334
rect 514262 478778 549706 479334
rect 550262 478778 592062 479334
rect 592618 478778 592650 479334
rect -8726 478746 592650 478778
rect -8726 478094 592650 478126
rect -8726 477538 -7734 478094
rect -7178 477538 8466 478094
rect 9022 477538 44466 478094
rect 45022 477538 80466 478094
rect 81022 477538 116466 478094
rect 117022 477538 152466 478094
rect 153022 477538 188466 478094
rect 189022 477538 224466 478094
rect 225022 477538 260466 478094
rect 261022 477538 296466 478094
rect 297022 477538 332466 478094
rect 333022 477538 368466 478094
rect 369022 477538 404466 478094
rect 405022 477538 440466 478094
rect 441022 477538 476466 478094
rect 477022 477538 512466 478094
rect 513022 477538 548466 478094
rect 549022 477538 591102 478094
rect 591658 477538 592650 478094
rect -8726 477506 592650 477538
rect -8726 476854 592650 476886
rect -8726 476298 -6774 476854
rect -6218 476298 7226 476854
rect 7782 476298 43226 476854
rect 43782 476298 79226 476854
rect 79782 476298 115226 476854
rect 115782 476298 151226 476854
rect 151782 476298 187226 476854
rect 187782 476298 223226 476854
rect 223782 476298 259226 476854
rect 259782 476298 295226 476854
rect 295782 476298 331226 476854
rect 331782 476298 367226 476854
rect 367782 476298 403226 476854
rect 403782 476298 439226 476854
rect 439782 476298 475226 476854
rect 475782 476298 511226 476854
rect 511782 476298 547226 476854
rect 547782 476298 590142 476854
rect 590698 476298 592650 476854
rect -8726 476266 592650 476298
rect -8726 475614 592650 475646
rect -8726 475058 -5814 475614
rect -5258 475058 5986 475614
rect 6542 475058 41986 475614
rect 42542 475058 77986 475614
rect 78542 475058 113986 475614
rect 114542 475058 149986 475614
rect 150542 475058 185986 475614
rect 186542 475058 221986 475614
rect 222542 475058 257986 475614
rect 258542 475058 293986 475614
rect 294542 475058 329986 475614
rect 330542 475058 365986 475614
rect 366542 475058 401986 475614
rect 402542 475058 437986 475614
rect 438542 475058 473986 475614
rect 474542 475058 509986 475614
rect 510542 475058 545986 475614
rect 546542 475058 581986 475614
rect 582542 475058 589182 475614
rect 589738 475058 592650 475614
rect -8726 475026 592650 475058
rect -8726 474374 592650 474406
rect -8726 473818 -4854 474374
rect -4298 473818 4746 474374
rect 5302 473818 40746 474374
rect 41302 473818 76746 474374
rect 77302 473818 112746 474374
rect 113302 473818 148746 474374
rect 149302 473818 184746 474374
rect 185302 473818 220746 474374
rect 221302 473818 256746 474374
rect 257302 473818 292746 474374
rect 293302 473818 328746 474374
rect 329302 473818 364746 474374
rect 365302 473818 400746 474374
rect 401302 473818 436746 474374
rect 437302 473818 472746 474374
rect 473302 473818 508746 474374
rect 509302 473818 544746 474374
rect 545302 473818 580746 474374
rect 581302 473818 588222 474374
rect 588778 473818 592650 474374
rect -8726 473786 592650 473818
rect -8726 473134 592650 473166
rect -8726 472578 -3894 473134
rect -3338 472578 3506 473134
rect 4062 472578 39506 473134
rect 40062 472578 75506 473134
rect 76062 472578 111506 473134
rect 112062 472578 147506 473134
rect 148062 472578 183506 473134
rect 184062 472578 219506 473134
rect 220062 472578 255506 473134
rect 256062 472578 291506 473134
rect 292062 472578 327506 473134
rect 328062 472578 363506 473134
rect 364062 472578 399506 473134
rect 400062 472578 435506 473134
rect 436062 472578 471506 473134
rect 472062 472578 507506 473134
rect 508062 472578 543506 473134
rect 544062 472578 579506 473134
rect 580062 472578 587262 473134
rect 587818 472578 592650 473134
rect -8726 472546 592650 472578
rect -8726 471894 592650 471926
rect -8726 471338 -2934 471894
rect -2378 471338 2266 471894
rect 2822 471338 38266 471894
rect 38822 471338 74266 471894
rect 74822 471338 110266 471894
rect 110822 471338 146266 471894
rect 146822 471338 182266 471894
rect 182822 471338 218266 471894
rect 218822 471338 254266 471894
rect 254822 471338 290266 471894
rect 290822 471338 326266 471894
rect 326822 471338 362266 471894
rect 362822 471338 398266 471894
rect 398822 471338 434266 471894
rect 434822 471338 470266 471894
rect 470822 471338 506266 471894
rect 506822 471338 542266 471894
rect 542822 471338 578266 471894
rect 578822 471338 586302 471894
rect 586858 471338 592650 471894
rect -8726 471306 592650 471338
rect -8726 470654 592650 470686
rect -8726 470098 -1974 470654
rect -1418 470098 1026 470654
rect 1582 470098 37026 470654
rect 37582 470098 73026 470654
rect 73582 470098 109026 470654
rect 109582 470098 145026 470654
rect 145582 470098 181026 470654
rect 181582 470098 217026 470654
rect 217582 470098 253026 470654
rect 253582 470098 289026 470654
rect 289582 470098 325026 470654
rect 325582 470098 361026 470654
rect 361582 470098 397026 470654
rect 397582 470098 433026 470654
rect 433582 470098 469026 470654
rect 469582 470098 505026 470654
rect 505582 470098 541026 470654
rect 541582 470098 577026 470654
rect 577582 470098 585342 470654
rect 585898 470098 592650 470654
rect -8726 470066 592650 470098
rect -8726 443334 592650 443366
rect -8726 442778 -8694 443334
rect -8138 442778 9706 443334
rect 10262 442778 45706 443334
rect 46262 442778 81706 443334
rect 82262 442778 117706 443334
rect 118262 442778 153706 443334
rect 154262 442778 189706 443334
rect 190262 442778 225706 443334
rect 226262 442778 261706 443334
rect 262262 442778 297706 443334
rect 298262 442778 333706 443334
rect 334262 442778 369706 443334
rect 370262 442778 405706 443334
rect 406262 442778 441706 443334
rect 442262 442778 477706 443334
rect 478262 442778 513706 443334
rect 514262 442778 549706 443334
rect 550262 442778 592062 443334
rect 592618 442778 592650 443334
rect -8726 442746 592650 442778
rect -8726 442094 592650 442126
rect -8726 441538 -7734 442094
rect -7178 441538 8466 442094
rect 9022 441538 44466 442094
rect 45022 441538 80466 442094
rect 81022 441538 116466 442094
rect 117022 441538 152466 442094
rect 153022 441538 188466 442094
rect 189022 441538 224466 442094
rect 225022 441538 260466 442094
rect 261022 441538 296466 442094
rect 297022 441538 332466 442094
rect 333022 441538 368466 442094
rect 369022 441538 404466 442094
rect 405022 441538 440466 442094
rect 441022 441538 476466 442094
rect 477022 441538 512466 442094
rect 513022 441538 548466 442094
rect 549022 441538 591102 442094
rect 591658 441538 592650 442094
rect -8726 441506 592650 441538
rect -8726 440854 592650 440886
rect -8726 440298 -6774 440854
rect -6218 440298 7226 440854
rect 7782 440298 43226 440854
rect 43782 440298 79226 440854
rect 79782 440298 115226 440854
rect 115782 440298 151226 440854
rect 151782 440298 187226 440854
rect 187782 440298 223226 440854
rect 223782 440298 259226 440854
rect 259782 440298 295226 440854
rect 295782 440298 331226 440854
rect 331782 440298 367226 440854
rect 367782 440298 403226 440854
rect 403782 440298 439226 440854
rect 439782 440298 475226 440854
rect 475782 440298 511226 440854
rect 511782 440298 547226 440854
rect 547782 440298 590142 440854
rect 590698 440298 592650 440854
rect -8726 440266 592650 440298
rect -8726 439614 592650 439646
rect -8726 439058 -5814 439614
rect -5258 439058 5986 439614
rect 6542 439058 41986 439614
rect 42542 439058 77986 439614
rect 78542 439058 113986 439614
rect 114542 439058 149986 439614
rect 150542 439058 185986 439614
rect 186542 439058 221986 439614
rect 222542 439058 257986 439614
rect 258542 439058 293986 439614
rect 294542 439058 329986 439614
rect 330542 439058 365986 439614
rect 366542 439058 401986 439614
rect 402542 439058 437986 439614
rect 438542 439058 473986 439614
rect 474542 439058 509986 439614
rect 510542 439058 581986 439614
rect 582542 439058 589182 439614
rect 589738 439058 592650 439614
rect -8726 439026 592650 439058
rect -8726 438374 592650 438406
rect -8726 437818 -4854 438374
rect -4298 437818 4746 438374
rect 5302 437818 40746 438374
rect 41302 437818 76746 438374
rect 77302 437818 112746 438374
rect 113302 437818 148746 438374
rect 149302 437818 184746 438374
rect 185302 437818 220746 438374
rect 221302 437818 256746 438374
rect 257302 437818 292746 438374
rect 293302 437818 328746 438374
rect 329302 437818 364746 438374
rect 365302 437818 400746 438374
rect 401302 437818 436746 438374
rect 437302 437818 472746 438374
rect 473302 437818 508746 438374
rect 509302 437818 580746 438374
rect 581302 437818 588222 438374
rect 588778 437818 592650 438374
rect -8726 437786 592650 437818
rect -8726 437134 592650 437166
rect -8726 436578 -3894 437134
rect -3338 436578 3506 437134
rect 4062 436578 39506 437134
rect 40062 436578 75506 437134
rect 76062 436578 111506 437134
rect 112062 436578 147506 437134
rect 148062 436578 183506 437134
rect 184062 436578 219506 437134
rect 220062 436578 255506 437134
rect 256062 436578 291506 437134
rect 292062 436578 327506 437134
rect 328062 436578 363506 437134
rect 364062 436578 399506 437134
rect 400062 436578 435506 437134
rect 436062 436578 471506 437134
rect 472062 436578 507506 437134
rect 508062 436578 579506 437134
rect 580062 436578 587262 437134
rect 587818 436578 592650 437134
rect -8726 436546 592650 436578
rect -8726 435894 592650 435926
rect -8726 435338 -2934 435894
rect -2378 435338 2266 435894
rect 2822 435338 38266 435894
rect 38822 435338 74266 435894
rect 74822 435338 110266 435894
rect 110822 435338 146266 435894
rect 146822 435338 182266 435894
rect 182822 435338 218266 435894
rect 218822 435338 254266 435894
rect 254822 435338 290266 435894
rect 290822 435338 326266 435894
rect 326822 435338 362266 435894
rect 362822 435338 398266 435894
rect 398822 435338 434266 435894
rect 434822 435338 470266 435894
rect 470822 435338 506266 435894
rect 506822 435658 540918 435894
rect 541154 435658 542850 435894
rect 543086 435658 544782 435894
rect 545018 435658 546714 435894
rect 546950 435658 578266 435894
rect 506822 435574 578266 435658
rect 506822 435338 540918 435574
rect 541154 435338 542850 435574
rect 543086 435338 544782 435574
rect 545018 435338 546714 435574
rect 546950 435338 578266 435574
rect 578822 435338 586302 435894
rect 586858 435338 592650 435894
rect -8726 435306 592650 435338
rect -8726 434654 592650 434686
rect -8726 434098 -1974 434654
rect -1418 434098 1026 434654
rect 1582 434098 37026 434654
rect 37582 434098 73026 434654
rect 73582 434098 109026 434654
rect 109582 434098 145026 434654
rect 145582 434098 181026 434654
rect 181582 434098 217026 434654
rect 217582 434098 253026 434654
rect 253582 434098 289026 434654
rect 289582 434098 325026 434654
rect 325582 434098 361026 434654
rect 361582 434098 397026 434654
rect 397582 434098 433026 434654
rect 433582 434098 469026 434654
rect 469582 434098 505026 434654
rect 505582 434418 539952 434654
rect 540188 434418 541884 434654
rect 542120 434418 543816 434654
rect 544052 434418 545748 434654
rect 545984 434418 577026 434654
rect 505582 434334 577026 434418
rect 505582 434098 539952 434334
rect 540188 434098 541884 434334
rect 542120 434098 543816 434334
rect 544052 434098 545748 434334
rect 545984 434098 577026 434334
rect 577582 434098 585342 434654
rect 585898 434098 592650 434654
rect -8726 434066 592650 434098
rect -8726 407334 592650 407366
rect -8726 406778 -8694 407334
rect -8138 406778 9706 407334
rect 10262 406778 45706 407334
rect 46262 406778 81706 407334
rect 82262 406778 117706 407334
rect 118262 406778 153706 407334
rect 154262 406778 189706 407334
rect 190262 406778 225706 407334
rect 226262 406778 261706 407334
rect 262262 406778 297706 407334
rect 298262 406778 333706 407334
rect 334262 406778 369706 407334
rect 370262 406778 405706 407334
rect 406262 406778 441706 407334
rect 442262 406778 477706 407334
rect 478262 406778 513706 407334
rect 514262 406778 549706 407334
rect 550262 406778 592062 407334
rect 592618 406778 592650 407334
rect -8726 406746 592650 406778
rect -8726 406094 592650 406126
rect -8726 405538 -7734 406094
rect -7178 405538 8466 406094
rect 9022 405538 44466 406094
rect 45022 405538 80466 406094
rect 81022 405538 116466 406094
rect 117022 405538 152466 406094
rect 153022 405538 188466 406094
rect 189022 405538 224466 406094
rect 225022 405538 260466 406094
rect 261022 405538 296466 406094
rect 297022 405538 332466 406094
rect 333022 405538 368466 406094
rect 369022 405538 404466 406094
rect 405022 405538 440466 406094
rect 441022 405538 476466 406094
rect 477022 405538 512466 406094
rect 513022 405538 548466 406094
rect 549022 405538 591102 406094
rect 591658 405538 592650 406094
rect -8726 405506 592650 405538
rect -8726 404854 592650 404886
rect -8726 404298 -6774 404854
rect -6218 404298 7226 404854
rect 7782 404298 43226 404854
rect 43782 404298 79226 404854
rect 79782 404298 115226 404854
rect 115782 404298 151226 404854
rect 151782 404298 187226 404854
rect 187782 404298 223226 404854
rect 223782 404298 259226 404854
rect 259782 404298 295226 404854
rect 295782 404298 331226 404854
rect 331782 404298 367226 404854
rect 367782 404298 403226 404854
rect 403782 404298 439226 404854
rect 439782 404298 475226 404854
rect 475782 404298 511226 404854
rect 511782 404298 547226 404854
rect 547782 404298 590142 404854
rect 590698 404298 592650 404854
rect -8726 404266 592650 404298
rect -8726 403614 592650 403646
rect -8726 403058 -5814 403614
rect -5258 403058 5986 403614
rect 6542 403058 41986 403614
rect 42542 403058 77986 403614
rect 78542 403058 113986 403614
rect 114542 403058 149986 403614
rect 150542 403058 185986 403614
rect 186542 403058 221986 403614
rect 222542 403058 257986 403614
rect 258542 403058 293986 403614
rect 294542 403058 329986 403614
rect 330542 403058 365986 403614
rect 366542 403058 401986 403614
rect 402542 403058 437986 403614
rect 438542 403058 473986 403614
rect 474542 403058 509986 403614
rect 510542 403058 581986 403614
rect 582542 403058 589182 403614
rect 589738 403058 592650 403614
rect -8726 403026 592650 403058
rect -8726 402374 592650 402406
rect -8726 401818 -4854 402374
rect -4298 401818 4746 402374
rect 5302 401818 40746 402374
rect 41302 401818 76746 402374
rect 77302 401818 112746 402374
rect 113302 401818 148746 402374
rect 149302 401818 184746 402374
rect 185302 401818 220746 402374
rect 221302 401818 256746 402374
rect 257302 401818 292746 402374
rect 293302 401818 328746 402374
rect 329302 401818 364746 402374
rect 365302 401818 400746 402374
rect 401302 401818 436746 402374
rect 437302 401818 472746 402374
rect 473302 401818 508746 402374
rect 509302 401818 580746 402374
rect 581302 401818 588222 402374
rect 588778 401818 592650 402374
rect -8726 401786 592650 401818
rect -8726 401134 592650 401166
rect -8726 400578 -3894 401134
rect -3338 400578 3506 401134
rect 4062 400578 39506 401134
rect 40062 400578 75506 401134
rect 76062 400578 111506 401134
rect 112062 400578 147506 401134
rect 148062 400578 183506 401134
rect 184062 400578 219506 401134
rect 220062 400578 255506 401134
rect 256062 400578 291506 401134
rect 292062 400578 327506 401134
rect 328062 400578 363506 401134
rect 364062 400578 399506 401134
rect 400062 400578 435506 401134
rect 436062 400578 471506 401134
rect 472062 400578 507506 401134
rect 508062 400578 579506 401134
rect 580062 400578 587262 401134
rect 587818 400578 592650 401134
rect -8726 400546 592650 400578
rect -8726 399894 592650 399926
rect -8726 399338 -2934 399894
rect -2378 399338 2266 399894
rect 2822 399338 38266 399894
rect 38822 399338 74266 399894
rect 74822 399338 110266 399894
rect 110822 399338 146266 399894
rect 146822 399338 182266 399894
rect 182822 399338 218266 399894
rect 218822 399338 254266 399894
rect 254822 399338 290266 399894
rect 290822 399338 326266 399894
rect 326822 399338 362266 399894
rect 362822 399338 398266 399894
rect 398822 399338 434266 399894
rect 434822 399338 470266 399894
rect 470822 399338 506266 399894
rect 506822 399658 540918 399894
rect 541154 399658 542850 399894
rect 543086 399658 544782 399894
rect 545018 399658 546714 399894
rect 546950 399658 578266 399894
rect 506822 399574 578266 399658
rect 506822 399338 540918 399574
rect 541154 399338 542850 399574
rect 543086 399338 544782 399574
rect 545018 399338 546714 399574
rect 546950 399338 578266 399574
rect 578822 399338 586302 399894
rect 586858 399338 592650 399894
rect -8726 399306 592650 399338
rect -8726 398654 592650 398686
rect -8726 398098 -1974 398654
rect -1418 398098 1026 398654
rect 1582 398098 37026 398654
rect 37582 398098 73026 398654
rect 73582 398098 109026 398654
rect 109582 398098 145026 398654
rect 145582 398098 181026 398654
rect 181582 398098 217026 398654
rect 217582 398098 253026 398654
rect 253582 398098 289026 398654
rect 289582 398098 325026 398654
rect 325582 398098 361026 398654
rect 361582 398098 397026 398654
rect 397582 398098 433026 398654
rect 433582 398098 469026 398654
rect 469582 398098 505026 398654
rect 505582 398418 539952 398654
rect 540188 398418 541884 398654
rect 542120 398418 543816 398654
rect 544052 398418 545748 398654
rect 545984 398418 577026 398654
rect 505582 398334 577026 398418
rect 505582 398098 539952 398334
rect 540188 398098 541884 398334
rect 542120 398098 543816 398334
rect 544052 398098 545748 398334
rect 545984 398098 577026 398334
rect 577582 398098 585342 398654
rect 585898 398098 592650 398654
rect -8726 398066 592650 398098
rect -8726 371334 592650 371366
rect -8726 370778 -8694 371334
rect -8138 370778 9706 371334
rect 10262 370778 45706 371334
rect 46262 370778 81706 371334
rect 82262 370778 117706 371334
rect 118262 370778 153706 371334
rect 154262 370778 189706 371334
rect 190262 370778 225706 371334
rect 226262 370778 261706 371334
rect 262262 370778 297706 371334
rect 298262 370778 333706 371334
rect 334262 370778 369706 371334
rect 370262 370778 405706 371334
rect 406262 370778 441706 371334
rect 442262 370778 477706 371334
rect 478262 370778 513706 371334
rect 514262 370778 549706 371334
rect 550262 370778 592062 371334
rect 592618 370778 592650 371334
rect -8726 370746 592650 370778
rect -8726 370094 592650 370126
rect -8726 369538 -7734 370094
rect -7178 369538 8466 370094
rect 9022 369538 44466 370094
rect 45022 369538 80466 370094
rect 81022 369538 116466 370094
rect 117022 369538 152466 370094
rect 153022 369538 188466 370094
rect 189022 369538 224466 370094
rect 225022 369538 260466 370094
rect 261022 369538 296466 370094
rect 297022 369538 332466 370094
rect 333022 369538 368466 370094
rect 369022 369538 404466 370094
rect 405022 369538 440466 370094
rect 441022 369538 512466 370094
rect 513022 369538 548466 370094
rect 549022 369538 591102 370094
rect 591658 369538 592650 370094
rect -8726 369506 592650 369538
rect -8726 368854 592650 368886
rect -8726 368298 -6774 368854
rect -6218 368298 7226 368854
rect 7782 368298 43226 368854
rect 43782 368298 79226 368854
rect 79782 368298 115226 368854
rect 115782 368298 151226 368854
rect 151782 368298 187226 368854
rect 187782 368298 223226 368854
rect 223782 368298 259226 368854
rect 259782 368298 295226 368854
rect 295782 368298 331226 368854
rect 331782 368298 367226 368854
rect 367782 368298 403226 368854
rect 403782 368298 439226 368854
rect 439782 368298 511226 368854
rect 511782 368298 547226 368854
rect 547782 368298 590142 368854
rect 590698 368298 592650 368854
rect -8726 368266 592650 368298
rect -8726 367614 592650 367646
rect -8726 367058 -5814 367614
rect -5258 367058 5986 367614
rect 6542 367058 41986 367614
rect 42542 367058 77986 367614
rect 78542 367058 113986 367614
rect 114542 367058 149986 367614
rect 150542 367058 185986 367614
rect 186542 367058 221986 367614
rect 222542 367058 257986 367614
rect 258542 367058 293986 367614
rect 294542 367058 329986 367614
rect 330542 367058 365986 367614
rect 366542 367058 401986 367614
rect 402542 367058 437986 367614
rect 438542 367058 509986 367614
rect 510542 367058 581986 367614
rect 582542 367058 589182 367614
rect 589738 367058 592650 367614
rect -8726 367026 592650 367058
rect -8726 366374 592650 366406
rect -8726 365818 -4854 366374
rect -4298 365818 4746 366374
rect 5302 365818 40746 366374
rect 41302 365818 76746 366374
rect 77302 365818 112746 366374
rect 113302 365818 148746 366374
rect 149302 365818 184746 366374
rect 185302 365818 220746 366374
rect 221302 365818 256746 366374
rect 257302 365818 292746 366374
rect 293302 365818 328746 366374
rect 329302 365818 364746 366374
rect 365302 365818 400746 366374
rect 401302 365818 436746 366374
rect 437302 366119 508746 366374
rect 437302 365883 472746 366119
rect 472982 365883 473066 366119
rect 473302 365883 508746 366119
rect 437302 365818 508746 365883
rect 509302 365818 580746 366374
rect 581302 365818 588222 366374
rect 588778 365818 592650 366374
rect -8726 365786 592650 365818
rect -8726 365134 592650 365166
rect -8726 364578 -3894 365134
rect -3338 364578 3506 365134
rect 4062 364578 39506 365134
rect 40062 364578 75506 365134
rect 76062 364578 111506 365134
rect 112062 364578 147506 365134
rect 148062 364578 183506 365134
rect 184062 364578 219506 365134
rect 220062 364578 255506 365134
rect 256062 364578 291506 365134
rect 292062 364578 327506 365134
rect 328062 364578 363506 365134
rect 364062 364578 399506 365134
rect 400062 364578 435506 365134
rect 436062 364578 471506 365134
rect 472062 364578 507506 365134
rect 508062 364578 579506 365134
rect 580062 364578 587262 365134
rect 587818 364578 592650 365134
rect -8726 364546 592650 364578
rect -8726 363894 592650 363926
rect -8726 363338 -2934 363894
rect -2378 363338 2266 363894
rect 2822 363338 38266 363894
rect 38822 363338 74266 363894
rect 74822 363338 110266 363894
rect 110822 363338 146266 363894
rect 146822 363338 182266 363894
rect 182822 363338 218266 363894
rect 218822 363338 254266 363894
rect 254822 363338 290266 363894
rect 290822 363338 326266 363894
rect 326822 363338 362266 363894
rect 362822 363338 398266 363894
rect 398822 363338 434266 363894
rect 434822 363338 470266 363894
rect 470822 363338 506266 363894
rect 506822 363658 540918 363894
rect 541154 363658 542850 363894
rect 543086 363658 544782 363894
rect 545018 363658 546714 363894
rect 546950 363658 578266 363894
rect 506822 363574 578266 363658
rect 506822 363338 540918 363574
rect 541154 363338 542850 363574
rect 543086 363338 544782 363574
rect 545018 363338 546714 363574
rect 546950 363338 578266 363574
rect 578822 363338 586302 363894
rect 586858 363338 592650 363894
rect -8726 363306 592650 363338
rect -8726 362654 592650 362686
rect -8726 362098 -1974 362654
rect -1418 362098 1026 362654
rect 1582 362098 37026 362654
rect 37582 362098 73026 362654
rect 73582 362098 109026 362654
rect 109582 362098 145026 362654
rect 145582 362098 181026 362654
rect 181582 362098 217026 362654
rect 217582 362098 253026 362654
rect 253582 362098 289026 362654
rect 289582 362098 325026 362654
rect 325582 362098 361026 362654
rect 361582 362098 397026 362654
rect 397582 362098 433026 362654
rect 433582 362098 469026 362654
rect 469582 362098 505026 362654
rect 505582 362418 539952 362654
rect 540188 362418 541884 362654
rect 542120 362418 543816 362654
rect 544052 362418 545748 362654
rect 545984 362418 577026 362654
rect 505582 362334 577026 362418
rect 505582 362098 539952 362334
rect 540188 362098 541884 362334
rect 542120 362098 543816 362334
rect 544052 362098 545748 362334
rect 545984 362098 577026 362334
rect 577582 362098 585342 362654
rect 585898 362098 592650 362654
rect -8726 362066 592650 362098
rect -8726 335334 592650 335366
rect -8726 334778 -8694 335334
rect -8138 334778 9706 335334
rect 10262 334778 45706 335334
rect 46262 334778 81706 335334
rect 82262 334778 117706 335334
rect 118262 334778 153706 335334
rect 154262 334778 189706 335334
rect 190262 334778 225706 335334
rect 226262 334778 261706 335334
rect 262262 334778 297706 335334
rect 298262 334778 333706 335334
rect 334262 334778 369706 335334
rect 370262 334778 405706 335334
rect 406262 334778 441706 335334
rect 442262 334778 477706 335334
rect 478262 334778 513706 335334
rect 514262 334778 549706 335334
rect 550262 334778 592062 335334
rect 592618 334778 592650 335334
rect -8726 334746 592650 334778
rect -8726 334094 592650 334126
rect -8726 333538 -7734 334094
rect -7178 333538 8466 334094
rect 9022 333538 44466 334094
rect 45022 333538 80466 334094
rect 81022 333538 116466 334094
rect 117022 333538 152466 334094
rect 153022 333538 188466 334094
rect 189022 333538 224466 334094
rect 225022 333538 260466 334094
rect 261022 333538 296466 334094
rect 297022 333538 332466 334094
rect 333022 333538 368466 334094
rect 369022 333538 404466 334094
rect 405022 333538 440466 334094
rect 441022 333538 476466 334094
rect 477022 333538 512466 334094
rect 513022 333538 548466 334094
rect 549022 333538 591102 334094
rect 591658 333538 592650 334094
rect -8726 333506 592650 333538
rect -8726 332854 592650 332886
rect -8726 332298 -6774 332854
rect -6218 332298 7226 332854
rect 7782 332298 43226 332854
rect 43782 332298 79226 332854
rect 79782 332298 115226 332854
rect 115782 332298 151226 332854
rect 151782 332298 187226 332854
rect 187782 332298 223226 332854
rect 223782 332298 259226 332854
rect 259782 332298 295226 332854
rect 295782 332298 331226 332854
rect 331782 332298 367226 332854
rect 367782 332298 403226 332854
rect 403782 332298 439226 332854
rect 439782 332298 475226 332854
rect 475782 332298 511226 332854
rect 511782 332298 547226 332854
rect 547782 332298 590142 332854
rect 590698 332298 592650 332854
rect -8726 332266 592650 332298
rect -8726 331614 592650 331646
rect -8726 331058 -5814 331614
rect -5258 331058 5986 331614
rect 6542 331058 41986 331614
rect 42542 331058 77986 331614
rect 78542 331058 113986 331614
rect 114542 331058 149986 331614
rect 150542 331058 185986 331614
rect 186542 331058 221986 331614
rect 222542 331058 257986 331614
rect 258542 331058 293986 331614
rect 294542 331058 329986 331614
rect 330542 331058 365986 331614
rect 366542 331058 401986 331614
rect 402542 331058 437986 331614
rect 438542 331058 473986 331614
rect 474542 331058 509986 331614
rect 510542 331058 581986 331614
rect 582542 331058 589182 331614
rect 589738 331058 592650 331614
rect -8726 331026 592650 331058
rect -8726 330374 592650 330406
rect -8726 329818 -4854 330374
rect -4298 329818 4746 330374
rect 5302 329818 40746 330374
rect 41302 329818 76746 330374
rect 77302 329818 112746 330374
rect 113302 329818 148746 330374
rect 149302 329818 184746 330374
rect 185302 329818 220746 330374
rect 221302 329818 256746 330374
rect 257302 329818 292746 330374
rect 293302 329818 328746 330374
rect 329302 329818 364746 330374
rect 365302 329818 400746 330374
rect 401302 329818 436746 330374
rect 437302 329818 472746 330374
rect 473302 329818 508746 330374
rect 509302 329818 580746 330374
rect 581302 329818 588222 330374
rect 588778 329818 592650 330374
rect -8726 329786 592650 329818
rect -8726 329134 592650 329166
rect -8726 328578 -3894 329134
rect -3338 328578 3506 329134
rect 4062 328578 39506 329134
rect 40062 328578 75506 329134
rect 76062 328578 111506 329134
rect 112062 328578 147506 329134
rect 148062 328578 183506 329134
rect 184062 328578 219506 329134
rect 220062 328578 255506 329134
rect 256062 328578 291506 329134
rect 292062 328578 327506 329134
rect 328062 328578 363506 329134
rect 364062 328578 399506 329134
rect 400062 328578 435506 329134
rect 436062 328578 471506 329134
rect 472062 328578 507506 329134
rect 508062 328578 579506 329134
rect 580062 328578 587262 329134
rect 587818 328578 592650 329134
rect -8726 328546 592650 328578
rect -8726 327894 592650 327926
rect -8726 327338 -2934 327894
rect -2378 327338 2266 327894
rect 2822 327338 38266 327894
rect 38822 327338 74266 327894
rect 74822 327338 110266 327894
rect 110822 327338 146266 327894
rect 146822 327338 182266 327894
rect 182822 327338 218266 327894
rect 218822 327338 254266 327894
rect 254822 327338 290266 327894
rect 290822 327338 326266 327894
rect 326822 327338 362266 327894
rect 362822 327338 398266 327894
rect 398822 327338 434266 327894
rect 434822 327338 470266 327894
rect 470822 327338 506266 327894
rect 506822 327658 540918 327894
rect 541154 327658 542850 327894
rect 543086 327658 544782 327894
rect 545018 327658 546714 327894
rect 546950 327658 578266 327894
rect 506822 327574 578266 327658
rect 506822 327338 540918 327574
rect 541154 327338 542850 327574
rect 543086 327338 544782 327574
rect 545018 327338 546714 327574
rect 546950 327338 578266 327574
rect 578822 327338 586302 327894
rect 586858 327338 592650 327894
rect -8726 327306 592650 327338
rect -8726 326654 592650 326686
rect -8726 326098 -1974 326654
rect -1418 326098 1026 326654
rect 1582 326098 37026 326654
rect 37582 326098 73026 326654
rect 73582 326098 109026 326654
rect 109582 326098 145026 326654
rect 145582 326098 181026 326654
rect 181582 326098 217026 326654
rect 217582 326098 253026 326654
rect 253582 326098 289026 326654
rect 289582 326098 325026 326654
rect 325582 326098 361026 326654
rect 361582 326098 397026 326654
rect 397582 326098 433026 326654
rect 433582 326098 469026 326654
rect 469582 326098 505026 326654
rect 505582 326418 539952 326654
rect 540188 326418 541884 326654
rect 542120 326418 543816 326654
rect 544052 326418 545748 326654
rect 545984 326418 577026 326654
rect 505582 326334 577026 326418
rect 505582 326098 539952 326334
rect 540188 326098 541884 326334
rect 542120 326098 543816 326334
rect 544052 326098 545748 326334
rect 545984 326098 577026 326334
rect 577582 326098 585342 326654
rect 585898 326098 592650 326654
rect -8726 326066 592650 326098
rect -8726 299334 592650 299366
rect -8726 298778 -8694 299334
rect -8138 298778 9706 299334
rect 10262 298778 45706 299334
rect 46262 298778 81706 299334
rect 82262 298778 117706 299334
rect 118262 298778 153706 299334
rect 154262 298778 189706 299334
rect 190262 298778 225706 299334
rect 226262 298778 261706 299334
rect 262262 298778 297706 299334
rect 298262 298778 333706 299334
rect 334262 298778 369706 299334
rect 370262 298778 405706 299334
rect 406262 298778 441706 299334
rect 442262 298778 477706 299334
rect 478262 298778 513706 299334
rect 514262 298778 549706 299334
rect 550262 298778 592062 299334
rect 592618 298778 592650 299334
rect -8726 298746 592650 298778
rect -8726 298094 592650 298126
rect -8726 297538 -7734 298094
rect -7178 297538 8466 298094
rect 9022 297538 44466 298094
rect 45022 297538 80466 298094
rect 81022 297538 116466 298094
rect 117022 297538 152466 298094
rect 153022 297538 188466 298094
rect 189022 297538 224466 298094
rect 225022 297538 260466 298094
rect 261022 297538 296466 298094
rect 297022 297538 332466 298094
rect 333022 297538 368466 298094
rect 369022 297538 404466 298094
rect 405022 297538 440466 298094
rect 441022 297538 476466 298094
rect 477022 297538 512466 298094
rect 513022 297538 548466 298094
rect 549022 297538 591102 298094
rect 591658 297538 592650 298094
rect -8726 297506 592650 297538
rect -8726 296854 592650 296886
rect -8726 296298 -6774 296854
rect -6218 296298 7226 296854
rect 7782 296298 43226 296854
rect 43782 296298 79226 296854
rect 79782 296298 115226 296854
rect 115782 296298 151226 296854
rect 151782 296298 187226 296854
rect 187782 296298 223226 296854
rect 223782 296298 259226 296854
rect 259782 296298 295226 296854
rect 295782 296298 331226 296854
rect 331782 296298 367226 296854
rect 367782 296298 403226 296854
rect 403782 296298 439226 296854
rect 439782 296298 475226 296854
rect 475782 296298 511226 296854
rect 511782 296298 547226 296854
rect 547782 296298 590142 296854
rect 590698 296298 592650 296854
rect -8726 296266 592650 296298
rect -8726 295614 592650 295646
rect -8726 295058 -5814 295614
rect -5258 295058 5986 295614
rect 6542 295058 41986 295614
rect 42542 295058 77986 295614
rect 78542 295058 113986 295614
rect 114542 295058 149986 295614
rect 150542 295058 185986 295614
rect 186542 295058 221986 295614
rect 222542 295058 257986 295614
rect 258542 295058 293986 295614
rect 294542 295058 329986 295614
rect 330542 295058 365986 295614
rect 366542 295058 401986 295614
rect 402542 295058 437986 295614
rect 438542 295058 473986 295614
rect 474542 295058 509986 295614
rect 510542 295058 581986 295614
rect 582542 295058 589182 295614
rect 589738 295058 592650 295614
rect -8726 295026 592650 295058
rect -8726 294374 592650 294406
rect -8726 293818 -4854 294374
rect -4298 293818 4746 294374
rect 5302 293818 40746 294374
rect 41302 293818 76746 294374
rect 77302 293818 112746 294374
rect 113302 293818 148746 294374
rect 149302 293818 184746 294374
rect 185302 293818 220746 294374
rect 221302 293818 256746 294374
rect 257302 293818 292746 294374
rect 293302 293818 328746 294374
rect 329302 293818 364746 294374
rect 365302 293818 400746 294374
rect 401302 293818 436746 294374
rect 437302 293818 472746 294374
rect 473302 293818 508746 294374
rect 509302 293818 580746 294374
rect 581302 293818 588222 294374
rect 588778 293818 592650 294374
rect -8726 293786 592650 293818
rect -8726 293134 592650 293166
rect -8726 292578 -3894 293134
rect -3338 292578 3506 293134
rect 4062 292578 39506 293134
rect 40062 292578 75506 293134
rect 76062 292578 111506 293134
rect 112062 292578 147506 293134
rect 148062 292578 183506 293134
rect 184062 292578 219506 293134
rect 220062 292578 255506 293134
rect 256062 292578 291506 293134
rect 292062 292578 327506 293134
rect 328062 292578 363506 293134
rect 364062 292578 399506 293134
rect 400062 292578 435506 293134
rect 436062 292578 471506 293134
rect 472062 292578 507506 293134
rect 508062 292578 579506 293134
rect 580062 292578 587262 293134
rect 587818 292578 592650 293134
rect -8726 292546 592650 292578
rect -8726 291894 592650 291926
rect -8726 291338 -2934 291894
rect -2378 291338 2266 291894
rect 2822 291338 38266 291894
rect 38822 291338 74266 291894
rect 74822 291338 110266 291894
rect 110822 291338 146266 291894
rect 146822 291338 182266 291894
rect 182822 291338 218266 291894
rect 218822 291338 254266 291894
rect 254822 291338 290266 291894
rect 290822 291338 326266 291894
rect 326822 291338 362266 291894
rect 362822 291338 398266 291894
rect 398822 291338 434266 291894
rect 434822 291338 470266 291894
rect 470822 291338 506266 291894
rect 506822 291658 540918 291894
rect 541154 291658 542850 291894
rect 543086 291658 544782 291894
rect 545018 291658 546714 291894
rect 546950 291658 578266 291894
rect 506822 291574 578266 291658
rect 506822 291338 540918 291574
rect 541154 291338 542850 291574
rect 543086 291338 544782 291574
rect 545018 291338 546714 291574
rect 546950 291338 578266 291574
rect 578822 291338 586302 291894
rect 586858 291338 592650 291894
rect -8726 291306 592650 291338
rect -8726 290654 592650 290686
rect -8726 290098 -1974 290654
rect -1418 290098 1026 290654
rect 1582 290098 37026 290654
rect 37582 290098 73026 290654
rect 73582 290098 109026 290654
rect 109582 290098 145026 290654
rect 145582 290098 181026 290654
rect 181582 290098 217026 290654
rect 217582 290098 253026 290654
rect 253582 290098 289026 290654
rect 289582 290098 325026 290654
rect 325582 290098 361026 290654
rect 361582 290098 397026 290654
rect 397582 290098 433026 290654
rect 433582 290098 469026 290654
rect 469582 290098 505026 290654
rect 505582 290418 539952 290654
rect 540188 290418 541884 290654
rect 542120 290418 543816 290654
rect 544052 290418 545748 290654
rect 545984 290418 577026 290654
rect 505582 290334 577026 290418
rect 505582 290098 539952 290334
rect 540188 290098 541884 290334
rect 542120 290098 543816 290334
rect 544052 290098 545748 290334
rect 545984 290098 577026 290334
rect 577582 290098 585342 290654
rect 585898 290098 592650 290654
rect -8726 290066 592650 290098
rect -8726 263334 592650 263366
rect -8726 262778 -8694 263334
rect -8138 262778 9706 263334
rect 10262 262778 45706 263334
rect 46262 262778 81706 263334
rect 82262 262778 117706 263334
rect 118262 262778 153706 263334
rect 154262 262778 189706 263334
rect 190262 262778 225706 263334
rect 226262 262778 261706 263334
rect 262262 262778 297706 263334
rect 298262 262778 333706 263334
rect 334262 262778 369706 263334
rect 370262 262778 405706 263334
rect 406262 262778 441706 263334
rect 442262 262778 513706 263334
rect 514262 262778 549706 263334
rect 550262 262778 592062 263334
rect 592618 262778 592650 263334
rect -8726 262746 592650 262778
rect -8726 262094 592650 262126
rect -8726 261538 -7734 262094
rect -7178 261538 8466 262094
rect 9022 261538 44466 262094
rect 45022 261538 80466 262094
rect 81022 261538 116466 262094
rect 117022 261538 152466 262094
rect 153022 261538 188466 262094
rect 189022 261538 224466 262094
rect 225022 261538 260466 262094
rect 261022 261538 296466 262094
rect 297022 261538 332466 262094
rect 333022 261538 368466 262094
rect 369022 261538 404466 262094
rect 405022 261538 440466 262094
rect 441022 261538 512466 262094
rect 513022 261538 548466 262094
rect 549022 261538 591102 262094
rect 591658 261538 592650 262094
rect -8726 261506 592650 261538
rect -8726 260854 592650 260886
rect -8726 260298 -6774 260854
rect -6218 260298 7226 260854
rect 7782 260298 43226 260854
rect 43782 260298 79226 260854
rect 79782 260298 115226 260854
rect 115782 260298 151226 260854
rect 151782 260298 187226 260854
rect 187782 260298 223226 260854
rect 223782 260298 259226 260854
rect 259782 260298 295226 260854
rect 295782 260298 331226 260854
rect 331782 260298 367226 260854
rect 367782 260298 403226 260854
rect 403782 260298 439226 260854
rect 439782 260298 475226 260854
rect 475782 260298 511226 260854
rect 511782 260298 547226 260854
rect 547782 260298 590142 260854
rect 590698 260298 592650 260854
rect -8726 260266 592650 260298
rect -8726 259614 592650 259646
rect -8726 259058 -5814 259614
rect -5258 259058 5986 259614
rect 6542 259058 41986 259614
rect 42542 259058 77986 259614
rect 78542 259058 113986 259614
rect 114542 259058 149986 259614
rect 150542 259058 185986 259614
rect 186542 259058 221986 259614
rect 222542 259058 257986 259614
rect 258542 259058 293986 259614
rect 294542 259058 329986 259614
rect 330542 259058 365986 259614
rect 366542 259058 401986 259614
rect 402542 259058 437986 259614
rect 438542 259058 473986 259614
rect 474542 259058 509986 259614
rect 510542 259058 545986 259614
rect 546542 259058 581986 259614
rect 582542 259058 589182 259614
rect 589738 259058 592650 259614
rect -8726 259026 592650 259058
rect -8726 258374 592650 258406
rect -8726 257818 -4854 258374
rect -4298 257818 4746 258374
rect 5302 257818 40746 258374
rect 41302 257818 76746 258374
rect 77302 257818 112746 258374
rect 113302 257818 148746 258374
rect 149302 257818 184746 258374
rect 185302 257818 220746 258374
rect 221302 257818 256746 258374
rect 257302 257818 292746 258374
rect 293302 257818 328746 258374
rect 329302 257818 364746 258374
rect 365302 257818 400746 258374
rect 401302 257818 436746 258374
rect 437302 257818 472746 258374
rect 473302 257818 508746 258374
rect 509302 257818 544746 258374
rect 545302 257818 580746 258374
rect 581302 257818 588222 258374
rect 588778 257818 592650 258374
rect -8726 257786 592650 257818
rect -8726 257134 592650 257166
rect -8726 256578 -3894 257134
rect -3338 256578 3506 257134
rect 4062 256578 39506 257134
rect 40062 256578 75506 257134
rect 76062 256578 111506 257134
rect 112062 256578 147506 257134
rect 148062 256578 183506 257134
rect 184062 256578 219506 257134
rect 220062 256578 255506 257134
rect 256062 256578 291506 257134
rect 292062 256578 327506 257134
rect 328062 256578 363506 257134
rect 364062 256578 399506 257134
rect 400062 256578 435506 257134
rect 436062 256578 471506 257134
rect 472062 256578 507506 257134
rect 508062 256578 543506 257134
rect 544062 256578 579506 257134
rect 580062 256578 587262 257134
rect 587818 256578 592650 257134
rect -8726 256546 592650 256578
rect -8726 255894 592650 255926
rect -8726 255338 -2934 255894
rect -2378 255338 2266 255894
rect 2822 255338 38266 255894
rect 38822 255338 74266 255894
rect 74822 255338 110266 255894
rect 110822 255338 146266 255894
rect 146822 255338 182266 255894
rect 182822 255338 218266 255894
rect 218822 255338 254266 255894
rect 254822 255338 290266 255894
rect 290822 255338 326266 255894
rect 326822 255338 362266 255894
rect 362822 255338 398266 255894
rect 398822 255338 434266 255894
rect 434822 255338 470266 255894
rect 470822 255338 506266 255894
rect 506822 255338 542266 255894
rect 542822 255338 578266 255894
rect 578822 255338 586302 255894
rect 586858 255338 592650 255894
rect -8726 255306 592650 255338
rect -8726 254654 592650 254686
rect -8726 254098 -1974 254654
rect -1418 254098 1026 254654
rect 1582 254098 37026 254654
rect 37582 254098 73026 254654
rect 73582 254098 109026 254654
rect 109582 254098 145026 254654
rect 145582 254098 181026 254654
rect 181582 254098 217026 254654
rect 217582 254098 253026 254654
rect 253582 254098 289026 254654
rect 289582 254098 325026 254654
rect 325582 254098 361026 254654
rect 361582 254098 397026 254654
rect 397582 254098 433026 254654
rect 433582 254098 469026 254654
rect 469582 254098 505026 254654
rect 505582 254098 541026 254654
rect 541582 254098 577026 254654
rect 577582 254098 585342 254654
rect 585898 254098 592650 254654
rect -8726 254066 592650 254098
rect -8726 227334 592650 227366
rect -8726 226778 -8694 227334
rect -8138 226778 9706 227334
rect 10262 226778 45706 227334
rect 46262 226778 81706 227334
rect 82262 226778 117706 227334
rect 118262 226778 153706 227334
rect 154262 226778 189706 227334
rect 190262 226778 225706 227334
rect 226262 226778 261706 227334
rect 262262 226778 297706 227334
rect 298262 226778 333706 227334
rect 334262 226778 369706 227334
rect 370262 226778 405706 227334
rect 406262 226778 441706 227334
rect 442262 226778 477706 227334
rect 478262 226778 513706 227334
rect 514262 226778 549706 227334
rect 550262 226778 592062 227334
rect 592618 226778 592650 227334
rect -8726 226746 592650 226778
rect -8726 226094 592650 226126
rect -8726 225538 -7734 226094
rect -7178 225538 8466 226094
rect 9022 225538 44466 226094
rect 45022 225538 80466 226094
rect 81022 225538 116466 226094
rect 117022 225538 152466 226094
rect 153022 225538 188466 226094
rect 189022 225538 224466 226094
rect 225022 225538 260466 226094
rect 261022 225538 296466 226094
rect 297022 225538 332466 226094
rect 333022 225538 368466 226094
rect 369022 225538 404466 226094
rect 405022 225538 440466 226094
rect 441022 225538 476466 226094
rect 477022 225538 512466 226094
rect 513022 225538 548466 226094
rect 549022 225538 591102 226094
rect 591658 225538 592650 226094
rect -8726 225506 592650 225538
rect -8726 224854 592650 224886
rect -8726 224298 -6774 224854
rect -6218 224298 7226 224854
rect 7782 224298 43226 224854
rect 43782 224298 79226 224854
rect 79782 224298 115226 224854
rect 115782 224298 151226 224854
rect 151782 224298 187226 224854
rect 187782 224298 223226 224854
rect 223782 224298 259226 224854
rect 259782 224298 295226 224854
rect 295782 224298 331226 224854
rect 331782 224298 367226 224854
rect 367782 224298 403226 224854
rect 403782 224298 439226 224854
rect 439782 224298 475226 224854
rect 475782 224298 511226 224854
rect 511782 224298 547226 224854
rect 547782 224298 590142 224854
rect 590698 224298 592650 224854
rect -8726 224266 592650 224298
rect -8726 223614 592650 223646
rect -8726 223058 -5814 223614
rect -5258 223058 5986 223614
rect 6542 223058 41986 223614
rect 42542 223058 77986 223614
rect 78542 223058 113986 223614
rect 114542 223058 149986 223614
rect 150542 223058 185986 223614
rect 186542 223058 221986 223614
rect 222542 223058 257986 223614
rect 258542 223058 293986 223614
rect 294542 223058 329986 223614
rect 330542 223058 365986 223614
rect 366542 223058 401986 223614
rect 402542 223058 437986 223614
rect 438542 223058 473986 223614
rect 474542 223058 509986 223614
rect 510542 223058 545986 223614
rect 546542 223058 581986 223614
rect 582542 223058 589182 223614
rect 589738 223058 592650 223614
rect -8726 223026 592650 223058
rect -8726 222374 592650 222406
rect -8726 221818 -4854 222374
rect -4298 221818 4746 222374
rect 5302 221818 40746 222374
rect 41302 221818 76746 222374
rect 77302 221818 112746 222374
rect 113302 221818 148746 222374
rect 149302 221818 184746 222374
rect 185302 221818 220746 222374
rect 221302 221818 256746 222374
rect 257302 221818 292746 222374
rect 293302 221818 328746 222374
rect 329302 221818 364746 222374
rect 365302 221818 400746 222374
rect 401302 221818 436746 222374
rect 437302 221818 472746 222374
rect 473302 221818 508746 222374
rect 509302 221818 544746 222374
rect 545302 221818 580746 222374
rect 581302 221818 588222 222374
rect 588778 221818 592650 222374
rect -8726 221786 592650 221818
rect -8726 221134 592650 221166
rect -8726 220578 -3894 221134
rect -3338 220578 3506 221134
rect 4062 220578 39506 221134
rect 40062 220578 75506 221134
rect 76062 220578 111506 221134
rect 112062 220578 147506 221134
rect 148062 220578 183506 221134
rect 184062 220578 219506 221134
rect 220062 220578 255506 221134
rect 256062 220578 291506 221134
rect 292062 220578 327506 221134
rect 328062 220578 363506 221134
rect 364062 220578 399506 221134
rect 400062 220578 435506 221134
rect 436062 220578 471506 221134
rect 472062 220578 507506 221134
rect 508062 220578 543506 221134
rect 544062 220578 579506 221134
rect 580062 220578 587262 221134
rect 587818 220578 592650 221134
rect -8726 220546 592650 220578
rect -8726 219894 592650 219926
rect -8726 219338 -2934 219894
rect -2378 219338 2266 219894
rect 2822 219338 38266 219894
rect 38822 219338 74266 219894
rect 74822 219338 110266 219894
rect 110822 219338 146266 219894
rect 146822 219338 182266 219894
rect 182822 219338 218266 219894
rect 218822 219338 254266 219894
rect 254822 219338 290266 219894
rect 290822 219338 326266 219894
rect 326822 219338 362266 219894
rect 362822 219338 398266 219894
rect 398822 219338 434266 219894
rect 434822 219338 470266 219894
rect 470822 219338 506266 219894
rect 506822 219338 542266 219894
rect 542822 219338 578266 219894
rect 578822 219338 586302 219894
rect 586858 219338 592650 219894
rect -8726 219306 592650 219338
rect -8726 218654 592650 218686
rect -8726 218098 -1974 218654
rect -1418 218098 1026 218654
rect 1582 218098 37026 218654
rect 37582 218098 73026 218654
rect 73582 218098 109026 218654
rect 109582 218098 145026 218654
rect 145582 218098 181026 218654
rect 181582 218098 217026 218654
rect 217582 218098 253026 218654
rect 253582 218098 289026 218654
rect 289582 218098 325026 218654
rect 325582 218098 361026 218654
rect 361582 218098 397026 218654
rect 397582 218098 433026 218654
rect 433582 218098 469026 218654
rect 469582 218098 505026 218654
rect 505582 218098 541026 218654
rect 541582 218098 577026 218654
rect 577582 218098 585342 218654
rect 585898 218098 592650 218654
rect -8726 218066 592650 218098
rect -8726 191334 592650 191366
rect -8726 190778 -8694 191334
rect -8138 190778 9706 191334
rect 10262 190778 45706 191334
rect 46262 190778 81706 191334
rect 82262 190778 117706 191334
rect 118262 190778 153706 191334
rect 154262 190778 189706 191334
rect 190262 190778 225706 191334
rect 226262 190778 261706 191334
rect 262262 190778 297706 191334
rect 298262 190778 333706 191334
rect 334262 190778 369706 191334
rect 370262 190778 405706 191334
rect 406262 190778 441706 191334
rect 442262 190778 477706 191334
rect 478262 190778 513706 191334
rect 514262 190778 549706 191334
rect 550262 190778 592062 191334
rect 592618 190778 592650 191334
rect -8726 190746 592650 190778
rect -8726 190094 592650 190126
rect -8726 189538 -7734 190094
rect -7178 189538 8466 190094
rect 9022 189538 44466 190094
rect 45022 189538 80466 190094
rect 81022 189538 116466 190094
rect 117022 189538 152466 190094
rect 153022 189538 188466 190094
rect 189022 189538 224466 190094
rect 225022 189538 260466 190094
rect 261022 189538 296466 190094
rect 297022 189538 332466 190094
rect 333022 189538 368466 190094
rect 369022 189538 404466 190094
rect 405022 189538 440466 190094
rect 441022 189538 476466 190094
rect 477022 189538 512466 190094
rect 513022 189538 548466 190094
rect 549022 189538 591102 190094
rect 591658 189538 592650 190094
rect -8726 189506 592650 189538
rect -8726 188854 592650 188886
rect -8726 188298 -6774 188854
rect -6218 188298 7226 188854
rect 7782 188298 43226 188854
rect 43782 188298 79226 188854
rect 79782 188298 115226 188854
rect 115782 188298 151226 188854
rect 151782 188298 187226 188854
rect 187782 188298 223226 188854
rect 223782 188298 259226 188854
rect 259782 188298 295226 188854
rect 295782 188298 331226 188854
rect 331782 188298 367226 188854
rect 367782 188298 403226 188854
rect 403782 188298 439226 188854
rect 439782 188298 475226 188854
rect 475782 188298 511226 188854
rect 511782 188298 547226 188854
rect 547782 188298 590142 188854
rect 590698 188298 592650 188854
rect -8726 188266 592650 188298
rect -8726 187614 592650 187646
rect -8726 187058 -5814 187614
rect -5258 187058 5986 187614
rect 6542 187058 41986 187614
rect 42542 187058 77986 187614
rect 78542 187058 113986 187614
rect 114542 187058 149986 187614
rect 150542 187058 185986 187614
rect 186542 187058 221986 187614
rect 222542 187058 257986 187614
rect 258542 187058 293986 187614
rect 294542 187058 329986 187614
rect 330542 187058 365986 187614
rect 366542 187058 401986 187614
rect 402542 187058 437986 187614
rect 438542 187058 473986 187614
rect 474542 187058 509986 187614
rect 510542 187058 545986 187614
rect 546542 187058 581986 187614
rect 582542 187058 589182 187614
rect 589738 187058 592650 187614
rect -8726 187026 592650 187058
rect -8726 186374 592650 186406
rect -8726 185818 -4854 186374
rect -4298 185818 4746 186374
rect 5302 185818 40746 186374
rect 41302 185818 76746 186374
rect 77302 185818 112746 186374
rect 113302 185818 148746 186374
rect 149302 185818 184746 186374
rect 185302 185818 220746 186374
rect 221302 185818 256746 186374
rect 257302 185818 292746 186374
rect 293302 185818 328746 186374
rect 329302 185818 364746 186374
rect 365302 185818 400746 186374
rect 401302 185818 436746 186374
rect 437302 185818 472746 186374
rect 473302 185818 508746 186374
rect 509302 185818 544746 186374
rect 545302 185818 580746 186374
rect 581302 185818 588222 186374
rect 588778 185818 592650 186374
rect -8726 185786 592650 185818
rect -8726 185134 592650 185166
rect -8726 184578 -3894 185134
rect -3338 184578 3506 185134
rect 4062 184578 39506 185134
rect 40062 184578 75506 185134
rect 76062 184578 111506 185134
rect 112062 184578 147506 185134
rect 148062 184578 183506 185134
rect 184062 184578 219506 185134
rect 220062 184578 255506 185134
rect 256062 184578 291506 185134
rect 292062 184578 327506 185134
rect 328062 184578 363506 185134
rect 364062 184578 399506 185134
rect 400062 184578 435506 185134
rect 436062 184578 471506 185134
rect 472062 184578 507506 185134
rect 508062 184578 543506 185134
rect 544062 184578 579506 185134
rect 580062 184578 587262 185134
rect 587818 184578 592650 185134
rect -8726 184546 592650 184578
rect -8726 183894 592650 183926
rect -8726 183338 -2934 183894
rect -2378 183338 2266 183894
rect 2822 183338 38266 183894
rect 38822 183338 74266 183894
rect 74822 183338 110266 183894
rect 110822 183338 146266 183894
rect 146822 183338 182266 183894
rect 182822 183338 218266 183894
rect 218822 183338 254266 183894
rect 254822 183338 290266 183894
rect 290822 183338 326266 183894
rect 326822 183338 362266 183894
rect 362822 183338 398266 183894
rect 398822 183338 434266 183894
rect 434822 183338 470266 183894
rect 470822 183338 506266 183894
rect 506822 183338 542266 183894
rect 542822 183338 578266 183894
rect 578822 183338 586302 183894
rect 586858 183338 592650 183894
rect -8726 183306 592650 183338
rect -8726 182654 592650 182686
rect -8726 182098 -1974 182654
rect -1418 182098 1026 182654
rect 1582 182098 37026 182654
rect 37582 182098 73026 182654
rect 73582 182098 109026 182654
rect 109582 182098 145026 182654
rect 145582 182098 181026 182654
rect 181582 182098 217026 182654
rect 217582 182098 253026 182654
rect 253582 182098 289026 182654
rect 289582 182098 325026 182654
rect 325582 182098 361026 182654
rect 361582 182098 397026 182654
rect 397582 182098 433026 182654
rect 433582 182098 469026 182654
rect 469582 182098 505026 182654
rect 505582 182098 541026 182654
rect 541582 182098 577026 182654
rect 577582 182098 585342 182654
rect 585898 182098 592650 182654
rect -8726 182066 592650 182098
rect -8726 155334 592650 155366
rect -8726 154778 -8694 155334
rect -8138 154778 9706 155334
rect 10262 154778 45706 155334
rect 46262 154778 81706 155334
rect 82262 154778 117706 155334
rect 118262 154778 153706 155334
rect 154262 154778 189706 155334
rect 190262 154778 225706 155334
rect 226262 154778 261706 155334
rect 262262 154778 297706 155334
rect 298262 154778 333706 155334
rect 334262 154778 369706 155334
rect 370262 154778 405706 155334
rect 406262 154778 441706 155334
rect 442262 154778 477706 155334
rect 478262 154778 513706 155334
rect 514262 154778 549706 155334
rect 550262 154778 592062 155334
rect 592618 154778 592650 155334
rect -8726 154746 592650 154778
rect -8726 154094 592650 154126
rect -8726 153538 -7734 154094
rect -7178 153538 8466 154094
rect 9022 153538 44466 154094
rect 45022 153538 80466 154094
rect 81022 153538 116466 154094
rect 117022 153538 152466 154094
rect 153022 153538 188466 154094
rect 189022 153538 224466 154094
rect 225022 153538 260466 154094
rect 261022 153538 296466 154094
rect 297022 153538 332466 154094
rect 333022 153538 368466 154094
rect 369022 153538 404466 154094
rect 405022 153538 440466 154094
rect 441022 153538 476466 154094
rect 477022 153538 512466 154094
rect 513022 153538 548466 154094
rect 549022 153538 591102 154094
rect 591658 153538 592650 154094
rect -8726 153506 592650 153538
rect -8726 152854 592650 152886
rect -8726 152298 -6774 152854
rect -6218 152298 7226 152854
rect 7782 152298 43226 152854
rect 43782 152298 79226 152854
rect 79782 152298 115226 152854
rect 115782 152298 151226 152854
rect 151782 152298 187226 152854
rect 187782 152298 223226 152854
rect 223782 152298 259226 152854
rect 259782 152298 295226 152854
rect 295782 152298 331226 152854
rect 331782 152298 367226 152854
rect 367782 152298 403226 152854
rect 403782 152298 439226 152854
rect 439782 152298 475226 152854
rect 475782 152298 511226 152854
rect 511782 152298 547226 152854
rect 547782 152298 590142 152854
rect 590698 152298 592650 152854
rect -8726 152266 592650 152298
rect -8726 151614 592650 151646
rect -8726 151058 -5814 151614
rect -5258 151058 5986 151614
rect 6542 151058 41986 151614
rect 42542 151058 77986 151614
rect 78542 151058 113986 151614
rect 114542 151058 149986 151614
rect 150542 151058 185986 151614
rect 186542 151058 221986 151614
rect 222542 151058 257986 151614
rect 258542 151058 293986 151614
rect 294542 151058 329986 151614
rect 330542 151058 365986 151614
rect 366542 151058 401986 151614
rect 402542 151058 437986 151614
rect 438542 151058 473986 151614
rect 474542 151058 509986 151614
rect 510542 151058 545986 151614
rect 546542 151058 581986 151614
rect 582542 151058 589182 151614
rect 589738 151058 592650 151614
rect -8726 151026 592650 151058
rect -8726 150374 592650 150406
rect -8726 149818 -4854 150374
rect -4298 149818 4746 150374
rect 5302 149818 40746 150374
rect 41302 149818 76746 150374
rect 77302 149818 112746 150374
rect 113302 149818 148746 150374
rect 149302 149818 184746 150374
rect 185302 149818 220746 150374
rect 221302 149818 256746 150374
rect 257302 149818 292746 150374
rect 293302 149818 328746 150374
rect 329302 149818 364746 150374
rect 365302 149818 400746 150374
rect 401302 149818 436746 150374
rect 437302 149818 472746 150374
rect 473302 149818 508746 150374
rect 509302 149818 544746 150374
rect 545302 149818 580746 150374
rect 581302 149818 588222 150374
rect 588778 149818 592650 150374
rect -8726 149786 592650 149818
rect -8726 149134 592650 149166
rect -8726 148578 -3894 149134
rect -3338 148578 3506 149134
rect 4062 148578 39506 149134
rect 40062 148578 75506 149134
rect 76062 148578 111506 149134
rect 112062 148578 147506 149134
rect 148062 148578 183506 149134
rect 184062 148578 219506 149134
rect 220062 148578 255506 149134
rect 256062 148578 291506 149134
rect 292062 148578 327506 149134
rect 328062 148578 363506 149134
rect 364062 148578 399506 149134
rect 400062 148578 435506 149134
rect 436062 148578 471506 149134
rect 472062 148578 507506 149134
rect 508062 148578 543506 149134
rect 544062 148578 579506 149134
rect 580062 148578 587262 149134
rect 587818 148578 592650 149134
rect -8726 148546 592650 148578
rect -8726 147894 592650 147926
rect -8726 147338 -2934 147894
rect -2378 147338 2266 147894
rect 2822 147338 38266 147894
rect 38822 147338 74266 147894
rect 74822 147338 110266 147894
rect 110822 147338 146266 147894
rect 146822 147338 182266 147894
rect 182822 147338 218266 147894
rect 218822 147338 254266 147894
rect 254822 147338 290266 147894
rect 290822 147338 326266 147894
rect 326822 147338 362266 147894
rect 362822 147338 398266 147894
rect 398822 147338 434266 147894
rect 434822 147338 470266 147894
rect 470822 147338 506266 147894
rect 506822 147338 542266 147894
rect 542822 147338 578266 147894
rect 578822 147338 586302 147894
rect 586858 147338 592650 147894
rect -8726 147306 592650 147338
rect -8726 146654 592650 146686
rect -8726 146098 -1974 146654
rect -1418 146098 1026 146654
rect 1582 146098 37026 146654
rect 37582 146098 73026 146654
rect 73582 146098 109026 146654
rect 109582 146098 145026 146654
rect 145582 146098 181026 146654
rect 181582 146098 217026 146654
rect 217582 146098 253026 146654
rect 253582 146098 289026 146654
rect 289582 146098 325026 146654
rect 325582 146098 361026 146654
rect 361582 146098 397026 146654
rect 397582 146098 433026 146654
rect 433582 146098 469026 146654
rect 469582 146098 505026 146654
rect 505582 146098 541026 146654
rect 541582 146098 577026 146654
rect 577582 146098 585342 146654
rect 585898 146098 592650 146654
rect -8726 146066 592650 146098
rect -8726 119334 592650 119366
rect -8726 118778 -8694 119334
rect -8138 118778 9706 119334
rect 10262 118778 45706 119334
rect 46262 118778 81706 119334
rect 82262 118778 117706 119334
rect 118262 118778 153706 119334
rect 154262 118778 189706 119334
rect 190262 118778 225706 119334
rect 226262 118778 261706 119334
rect 262262 118778 297706 119334
rect 298262 118778 333706 119334
rect 334262 118778 369706 119334
rect 370262 118778 405706 119334
rect 406262 118778 441706 119334
rect 442262 118778 477706 119334
rect 478262 118778 513706 119334
rect 514262 118778 549706 119334
rect 550262 118778 592062 119334
rect 592618 118778 592650 119334
rect -8726 118746 592650 118778
rect -8726 118094 592650 118126
rect -8726 117538 -7734 118094
rect -7178 117538 8466 118094
rect 9022 117538 44466 118094
rect 45022 117538 80466 118094
rect 81022 117538 116466 118094
rect 117022 117538 152466 118094
rect 153022 117538 188466 118094
rect 189022 117538 224466 118094
rect 225022 117538 260466 118094
rect 261022 117538 296466 118094
rect 297022 117538 332466 118094
rect 333022 117538 368466 118094
rect 369022 117538 404466 118094
rect 405022 117538 440466 118094
rect 441022 117538 476466 118094
rect 477022 117538 512466 118094
rect 513022 117538 548466 118094
rect 549022 117538 591102 118094
rect 591658 117538 592650 118094
rect -8726 117506 592650 117538
rect -8726 116854 592650 116886
rect -8726 116298 -6774 116854
rect -6218 116298 7226 116854
rect 7782 116298 43226 116854
rect 43782 116298 79226 116854
rect 79782 116298 115226 116854
rect 115782 116298 151226 116854
rect 151782 116298 187226 116854
rect 187782 116298 223226 116854
rect 223782 116298 259226 116854
rect 259782 116298 295226 116854
rect 295782 116298 331226 116854
rect 331782 116298 367226 116854
rect 367782 116298 403226 116854
rect 403782 116298 439226 116854
rect 439782 116298 475226 116854
rect 475782 116298 511226 116854
rect 511782 116298 547226 116854
rect 547782 116298 590142 116854
rect 590698 116298 592650 116854
rect -8726 116266 592650 116298
rect -8726 115614 592650 115646
rect -8726 115058 -5814 115614
rect -5258 115058 5986 115614
rect 6542 115058 41986 115614
rect 42542 115058 77986 115614
rect 78542 115058 113986 115614
rect 114542 115058 149986 115614
rect 150542 115058 185986 115614
rect 186542 115058 221986 115614
rect 222542 115058 257986 115614
rect 258542 115058 293986 115614
rect 294542 115058 329986 115614
rect 330542 115058 365986 115614
rect 366542 115058 401986 115614
rect 402542 115058 437986 115614
rect 438542 115058 473986 115614
rect 474542 115058 509986 115614
rect 510542 115058 545986 115614
rect 546542 115058 581986 115614
rect 582542 115058 589182 115614
rect 589738 115058 592650 115614
rect -8726 115026 592650 115058
rect -8726 114374 592650 114406
rect -8726 113818 -4854 114374
rect -4298 113818 4746 114374
rect 5302 113818 40746 114374
rect 41302 113818 76746 114374
rect 77302 113818 112746 114374
rect 113302 113818 148746 114374
rect 149302 113818 184746 114374
rect 185302 113818 220746 114374
rect 221302 113818 256746 114374
rect 257302 113818 292746 114374
rect 293302 113818 328746 114374
rect 329302 113818 364746 114374
rect 365302 113818 400746 114374
rect 401302 113818 436746 114374
rect 437302 113818 472746 114374
rect 473302 113818 508746 114374
rect 509302 113818 544746 114374
rect 545302 113818 580746 114374
rect 581302 113818 588222 114374
rect 588778 113818 592650 114374
rect -8726 113786 592650 113818
rect -8726 113134 592650 113166
rect -8726 112578 -3894 113134
rect -3338 112578 3506 113134
rect 4062 112578 39506 113134
rect 40062 112578 75506 113134
rect 76062 112578 111506 113134
rect 112062 112578 147506 113134
rect 148062 112578 183506 113134
rect 184062 112578 219506 113134
rect 220062 112578 255506 113134
rect 256062 112578 291506 113134
rect 292062 112578 327506 113134
rect 328062 112578 363506 113134
rect 364062 112578 399506 113134
rect 400062 112578 435506 113134
rect 436062 112578 471506 113134
rect 472062 112578 507506 113134
rect 508062 112578 543506 113134
rect 544062 112578 579506 113134
rect 580062 112578 587262 113134
rect 587818 112578 592650 113134
rect -8726 112546 592650 112578
rect -8726 111894 592650 111926
rect -8726 111338 -2934 111894
rect -2378 111338 2266 111894
rect 2822 111338 38266 111894
rect 38822 111338 74266 111894
rect 74822 111338 110266 111894
rect 110822 111338 146266 111894
rect 146822 111338 182266 111894
rect 182822 111338 218266 111894
rect 218822 111338 254266 111894
rect 254822 111338 290266 111894
rect 290822 111338 326266 111894
rect 326822 111338 362266 111894
rect 362822 111338 398266 111894
rect 398822 111338 434266 111894
rect 434822 111338 470266 111894
rect 470822 111338 506266 111894
rect 506822 111338 542266 111894
rect 542822 111338 578266 111894
rect 578822 111338 586302 111894
rect 586858 111338 592650 111894
rect -8726 111306 592650 111338
rect -8726 110654 592650 110686
rect -8726 110098 -1974 110654
rect -1418 110098 1026 110654
rect 1582 110098 37026 110654
rect 37582 110098 73026 110654
rect 73582 110098 109026 110654
rect 109582 110098 145026 110654
rect 145582 110098 181026 110654
rect 181582 110098 217026 110654
rect 217582 110098 253026 110654
rect 253582 110098 289026 110654
rect 289582 110098 325026 110654
rect 325582 110098 361026 110654
rect 361582 110098 397026 110654
rect 397582 110098 433026 110654
rect 433582 110098 469026 110654
rect 469582 110098 505026 110654
rect 505582 110098 541026 110654
rect 541582 110098 577026 110654
rect 577582 110098 585342 110654
rect 585898 110098 592650 110654
rect -8726 110066 592650 110098
rect -8726 83334 592650 83366
rect -8726 82778 -8694 83334
rect -8138 82778 9706 83334
rect 10262 82778 45706 83334
rect 46262 82778 81706 83334
rect 82262 82778 117706 83334
rect 118262 82778 153706 83334
rect 154262 82778 189706 83334
rect 190262 82778 225706 83334
rect 226262 82778 261706 83334
rect 262262 82778 297706 83334
rect 298262 82778 333706 83334
rect 334262 82778 369706 83334
rect 370262 82778 405706 83334
rect 406262 82778 441706 83334
rect 442262 82778 477706 83334
rect 478262 82778 513706 83334
rect 514262 82778 549706 83334
rect 550262 82778 592062 83334
rect 592618 82778 592650 83334
rect -8726 82746 592650 82778
rect -8726 82094 592650 82126
rect -8726 81538 -7734 82094
rect -7178 81538 8466 82094
rect 9022 81538 44466 82094
rect 45022 81538 80466 82094
rect 81022 81538 116466 82094
rect 117022 81538 152466 82094
rect 153022 81538 188466 82094
rect 189022 81538 224466 82094
rect 225022 81538 260466 82094
rect 261022 81538 296466 82094
rect 297022 81538 332466 82094
rect 333022 81538 368466 82094
rect 369022 81538 404466 82094
rect 405022 81538 440466 82094
rect 441022 81538 476466 82094
rect 477022 81538 512466 82094
rect 513022 81538 548466 82094
rect 549022 81538 591102 82094
rect 591658 81538 592650 82094
rect -8726 81506 592650 81538
rect -8726 80854 592650 80886
rect -8726 80298 -6774 80854
rect -6218 80298 7226 80854
rect 7782 80298 43226 80854
rect 43782 80298 79226 80854
rect 79782 80298 115226 80854
rect 115782 80298 151226 80854
rect 151782 80298 187226 80854
rect 187782 80298 223226 80854
rect 223782 80298 259226 80854
rect 259782 80298 295226 80854
rect 295782 80298 331226 80854
rect 331782 80298 367226 80854
rect 367782 80298 403226 80854
rect 403782 80298 439226 80854
rect 439782 80298 475226 80854
rect 475782 80298 511226 80854
rect 511782 80298 547226 80854
rect 547782 80298 590142 80854
rect 590698 80298 592650 80854
rect -8726 80266 592650 80298
rect -8726 79614 592650 79646
rect -8726 79058 -5814 79614
rect -5258 79058 5986 79614
rect 6542 79058 41986 79614
rect 42542 79058 77986 79614
rect 78542 79058 113986 79614
rect 114542 79058 149986 79614
rect 150542 79058 185986 79614
rect 186542 79058 221986 79614
rect 222542 79058 257986 79614
rect 258542 79058 293986 79614
rect 294542 79058 329986 79614
rect 330542 79058 365986 79614
rect 366542 79058 401986 79614
rect 402542 79058 437986 79614
rect 438542 79058 473986 79614
rect 474542 79058 509986 79614
rect 510542 79058 545986 79614
rect 546542 79058 581986 79614
rect 582542 79058 589182 79614
rect 589738 79058 592650 79614
rect -8726 79026 592650 79058
rect -8726 78374 592650 78406
rect -8726 77818 -4854 78374
rect -4298 77818 4746 78374
rect 5302 77818 40746 78374
rect 41302 77818 76746 78374
rect 77302 77818 112746 78374
rect 113302 77818 148746 78374
rect 149302 77818 184746 78374
rect 185302 77818 220746 78374
rect 221302 77818 256746 78374
rect 257302 77818 292746 78374
rect 293302 77818 328746 78374
rect 329302 77818 364746 78374
rect 365302 77818 400746 78374
rect 401302 77818 436746 78374
rect 437302 77818 472746 78374
rect 473302 77818 508746 78374
rect 509302 77818 544746 78374
rect 545302 77818 580746 78374
rect 581302 77818 588222 78374
rect 588778 77818 592650 78374
rect -8726 77786 592650 77818
rect -8726 77134 592650 77166
rect -8726 76578 -3894 77134
rect -3338 76578 3506 77134
rect 4062 76578 39506 77134
rect 40062 76578 75506 77134
rect 76062 76578 111506 77134
rect 112062 76578 147506 77134
rect 148062 76578 183506 77134
rect 184062 76578 219506 77134
rect 220062 76578 255506 77134
rect 256062 76578 291506 77134
rect 292062 76578 327506 77134
rect 328062 76578 363506 77134
rect 364062 76578 399506 77134
rect 400062 76578 435506 77134
rect 436062 76578 471506 77134
rect 472062 76578 507506 77134
rect 508062 76578 543506 77134
rect 544062 76578 579506 77134
rect 580062 76578 587262 77134
rect 587818 76578 592650 77134
rect -8726 76546 592650 76578
rect -8726 75894 592650 75926
rect -8726 75338 -2934 75894
rect -2378 75338 2266 75894
rect 2822 75338 38266 75894
rect 38822 75338 74266 75894
rect 74822 75338 110266 75894
rect 110822 75338 146266 75894
rect 146822 75338 182266 75894
rect 182822 75338 218266 75894
rect 218822 75338 254266 75894
rect 254822 75338 290266 75894
rect 290822 75338 326266 75894
rect 326822 75338 362266 75894
rect 362822 75338 398266 75894
rect 398822 75338 434266 75894
rect 434822 75338 470266 75894
rect 470822 75338 506266 75894
rect 506822 75338 542266 75894
rect 542822 75338 578266 75894
rect 578822 75338 586302 75894
rect 586858 75338 592650 75894
rect -8726 75306 592650 75338
rect -8726 74654 592650 74686
rect -8726 74098 -1974 74654
rect -1418 74098 1026 74654
rect 1582 74098 37026 74654
rect 37582 74098 73026 74654
rect 73582 74098 109026 74654
rect 109582 74098 145026 74654
rect 145582 74098 181026 74654
rect 181582 74098 217026 74654
rect 217582 74098 253026 74654
rect 253582 74098 289026 74654
rect 289582 74098 325026 74654
rect 325582 74098 361026 74654
rect 361582 74098 397026 74654
rect 397582 74098 433026 74654
rect 433582 74098 469026 74654
rect 469582 74098 505026 74654
rect 505582 74098 541026 74654
rect 541582 74098 577026 74654
rect 577582 74098 585342 74654
rect 585898 74098 592650 74654
rect -8726 74066 592650 74098
rect -8726 47334 592650 47366
rect -8726 46778 -8694 47334
rect -8138 46778 9706 47334
rect 10262 46778 45706 47334
rect 46262 46778 81706 47334
rect 82262 46778 117706 47334
rect 118262 46778 153706 47334
rect 154262 46778 189706 47334
rect 190262 46778 225706 47334
rect 226262 46778 261706 47334
rect 262262 46778 297706 47334
rect 298262 46778 333706 47334
rect 334262 46778 369706 47334
rect 370262 46778 405706 47334
rect 406262 46778 441706 47334
rect 442262 46778 477706 47334
rect 478262 46778 513706 47334
rect 514262 46778 549706 47334
rect 550262 46778 592062 47334
rect 592618 46778 592650 47334
rect -8726 46746 592650 46778
rect -8726 46094 592650 46126
rect -8726 45538 -7734 46094
rect -7178 45538 8466 46094
rect 9022 45538 44466 46094
rect 45022 45538 80466 46094
rect 81022 45538 116466 46094
rect 117022 45538 152466 46094
rect 153022 45538 188466 46094
rect 189022 45538 224466 46094
rect 225022 45538 260466 46094
rect 261022 45538 296466 46094
rect 297022 45538 332466 46094
rect 333022 45538 368466 46094
rect 369022 45538 404466 46094
rect 405022 45538 440466 46094
rect 441022 45538 476466 46094
rect 477022 45538 512466 46094
rect 513022 45538 548466 46094
rect 549022 45538 591102 46094
rect 591658 45538 592650 46094
rect -8726 45506 592650 45538
rect -8726 44854 592650 44886
rect -8726 44298 -6774 44854
rect -6218 44298 7226 44854
rect 7782 44298 43226 44854
rect 43782 44298 79226 44854
rect 79782 44298 115226 44854
rect 115782 44298 151226 44854
rect 151782 44298 187226 44854
rect 187782 44298 223226 44854
rect 223782 44298 259226 44854
rect 259782 44298 295226 44854
rect 295782 44298 331226 44854
rect 331782 44298 367226 44854
rect 367782 44298 403226 44854
rect 403782 44298 439226 44854
rect 439782 44298 475226 44854
rect 475782 44298 511226 44854
rect 511782 44298 547226 44854
rect 547782 44298 590142 44854
rect 590698 44298 592650 44854
rect -8726 44266 592650 44298
rect -8726 43614 592650 43646
rect -8726 43058 -5814 43614
rect -5258 43058 5986 43614
rect 6542 43058 41986 43614
rect 42542 43058 77986 43614
rect 78542 43058 113986 43614
rect 114542 43058 149986 43614
rect 150542 43058 185986 43614
rect 186542 43058 221986 43614
rect 222542 43058 257986 43614
rect 258542 43058 293986 43614
rect 294542 43058 329986 43614
rect 330542 43058 365986 43614
rect 366542 43058 401986 43614
rect 402542 43058 437986 43614
rect 438542 43058 473986 43614
rect 474542 43058 509986 43614
rect 510542 43058 545986 43614
rect 546542 43058 581986 43614
rect 582542 43058 589182 43614
rect 589738 43058 592650 43614
rect -8726 43026 592650 43058
rect -8726 42374 592650 42406
rect -8726 41818 -4854 42374
rect -4298 41818 4746 42374
rect 5302 41818 40746 42374
rect 41302 41818 76746 42374
rect 77302 41818 112746 42374
rect 113302 41818 148746 42374
rect 149302 41818 184746 42374
rect 185302 41818 220746 42374
rect 221302 41818 256746 42374
rect 257302 41818 292746 42374
rect 293302 41818 328746 42374
rect 329302 41818 364746 42374
rect 365302 41818 400746 42374
rect 401302 41818 436746 42374
rect 437302 41818 472746 42374
rect 473302 41818 508746 42374
rect 509302 41818 544746 42374
rect 545302 41818 580746 42374
rect 581302 41818 588222 42374
rect 588778 41818 592650 42374
rect -8726 41786 592650 41818
rect -8726 41134 592650 41166
rect -8726 40578 -3894 41134
rect -3338 40578 3506 41134
rect 4062 40578 39506 41134
rect 40062 40578 75506 41134
rect 76062 40578 111506 41134
rect 112062 40578 147506 41134
rect 148062 40578 183506 41134
rect 184062 40578 219506 41134
rect 220062 40578 255506 41134
rect 256062 40578 291506 41134
rect 292062 40578 327506 41134
rect 328062 40578 363506 41134
rect 364062 40578 399506 41134
rect 400062 40578 435506 41134
rect 436062 40578 471506 41134
rect 472062 40578 507506 41134
rect 508062 40578 543506 41134
rect 544062 40578 579506 41134
rect 580062 40578 587262 41134
rect 587818 40578 592650 41134
rect -8726 40546 592650 40578
rect -8726 39894 592650 39926
rect -8726 39338 -2934 39894
rect -2378 39338 2266 39894
rect 2822 39338 38266 39894
rect 38822 39338 74266 39894
rect 74822 39338 110266 39894
rect 110822 39338 146266 39894
rect 146822 39338 182266 39894
rect 182822 39338 218266 39894
rect 218822 39338 254266 39894
rect 254822 39338 290266 39894
rect 290822 39338 326266 39894
rect 326822 39338 362266 39894
rect 362822 39338 398266 39894
rect 398822 39338 434266 39894
rect 434822 39338 470266 39894
rect 470822 39338 506266 39894
rect 506822 39338 542266 39894
rect 542822 39338 578266 39894
rect 578822 39338 586302 39894
rect 586858 39338 592650 39894
rect -8726 39306 592650 39338
rect -8726 38654 592650 38686
rect -8726 38098 -1974 38654
rect -1418 38098 1026 38654
rect 1582 38098 37026 38654
rect 37582 38098 73026 38654
rect 73582 38098 109026 38654
rect 109582 38098 145026 38654
rect 145582 38098 181026 38654
rect 181582 38098 217026 38654
rect 217582 38098 253026 38654
rect 253582 38098 289026 38654
rect 289582 38098 325026 38654
rect 325582 38098 361026 38654
rect 361582 38098 397026 38654
rect 397582 38098 433026 38654
rect 433582 38098 469026 38654
rect 469582 38098 505026 38654
rect 505582 38098 541026 38654
rect 541582 38098 577026 38654
rect 577582 38098 585342 38654
rect 585898 38098 592650 38654
rect -8726 38066 592650 38098
rect -8726 11334 592650 11366
rect -8726 10778 -8694 11334
rect -8138 10778 9706 11334
rect 10262 10778 45706 11334
rect 46262 10778 81706 11334
rect 82262 10778 117706 11334
rect 118262 10778 153706 11334
rect 154262 10778 189706 11334
rect 190262 10778 225706 11334
rect 226262 10778 261706 11334
rect 262262 10778 297706 11334
rect 298262 10778 333706 11334
rect 334262 10778 369706 11334
rect 370262 10778 405706 11334
rect 406262 10778 441706 11334
rect 442262 10778 477706 11334
rect 478262 10778 513706 11334
rect 514262 10778 549706 11334
rect 550262 10778 592062 11334
rect 592618 10778 592650 11334
rect -8726 10746 592650 10778
rect -8726 10094 592650 10126
rect -8726 9538 -7734 10094
rect -7178 9538 8466 10094
rect 9022 9538 44466 10094
rect 45022 9538 80466 10094
rect 81022 9538 116466 10094
rect 117022 9538 152466 10094
rect 153022 9538 188466 10094
rect 189022 9538 224466 10094
rect 225022 9538 260466 10094
rect 261022 9538 296466 10094
rect 297022 9538 332466 10094
rect 333022 9538 368466 10094
rect 369022 9538 404466 10094
rect 405022 9538 440466 10094
rect 441022 9538 476466 10094
rect 477022 9538 512466 10094
rect 513022 9538 548466 10094
rect 549022 9538 591102 10094
rect 591658 9538 592650 10094
rect -8726 9506 592650 9538
rect -8726 8854 592650 8886
rect -8726 8298 -6774 8854
rect -6218 8298 7226 8854
rect 7782 8298 43226 8854
rect 43782 8298 79226 8854
rect 79782 8298 115226 8854
rect 115782 8298 151226 8854
rect 151782 8298 187226 8854
rect 187782 8298 223226 8854
rect 223782 8298 259226 8854
rect 259782 8298 295226 8854
rect 295782 8298 331226 8854
rect 331782 8298 367226 8854
rect 367782 8298 403226 8854
rect 403782 8298 439226 8854
rect 439782 8298 475226 8854
rect 475782 8298 511226 8854
rect 511782 8298 547226 8854
rect 547782 8298 590142 8854
rect 590698 8298 592650 8854
rect -8726 8266 592650 8298
rect -8726 7614 592650 7646
rect -8726 7058 -5814 7614
rect -5258 7058 5986 7614
rect 6542 7058 41986 7614
rect 42542 7058 77986 7614
rect 78542 7058 113986 7614
rect 114542 7058 149986 7614
rect 150542 7058 185986 7614
rect 186542 7058 221986 7614
rect 222542 7058 257986 7614
rect 258542 7058 293986 7614
rect 294542 7058 329986 7614
rect 330542 7058 365986 7614
rect 366542 7058 401986 7614
rect 402542 7058 437986 7614
rect 438542 7058 473986 7614
rect 474542 7058 509986 7614
rect 510542 7058 545986 7614
rect 546542 7058 581986 7614
rect 582542 7058 589182 7614
rect 589738 7058 592650 7614
rect -8726 7026 592650 7058
rect -8726 6374 592650 6406
rect -8726 5818 -4854 6374
rect -4298 5818 4746 6374
rect 5302 5818 40746 6374
rect 41302 5818 76746 6374
rect 77302 5818 112746 6374
rect 113302 5818 148746 6374
rect 149302 5818 184746 6374
rect 185302 5818 220746 6374
rect 221302 5818 256746 6374
rect 257302 5818 292746 6374
rect 293302 5818 328746 6374
rect 329302 5818 364746 6374
rect 365302 5818 400746 6374
rect 401302 5818 436746 6374
rect 437302 5818 472746 6374
rect 473302 5818 508746 6374
rect 509302 5818 544746 6374
rect 545302 5818 580746 6374
rect 581302 5818 588222 6374
rect 588778 5818 592650 6374
rect -8726 5786 592650 5818
rect -8726 5134 592650 5166
rect -8726 4578 -3894 5134
rect -3338 4578 3506 5134
rect 4062 4578 39506 5134
rect 40062 4578 75506 5134
rect 76062 4578 111506 5134
rect 112062 4578 147506 5134
rect 148062 4578 183506 5134
rect 184062 4578 219506 5134
rect 220062 4578 255506 5134
rect 256062 4578 291506 5134
rect 292062 4578 327506 5134
rect 328062 4578 363506 5134
rect 364062 4578 399506 5134
rect 400062 4578 435506 5134
rect 436062 4578 471506 5134
rect 472062 4578 507506 5134
rect 508062 4578 543506 5134
rect 544062 4578 579506 5134
rect 580062 4578 587262 5134
rect 587818 4578 592650 5134
rect -8726 4546 592650 4578
rect -8726 3894 592650 3926
rect -8726 3338 -2934 3894
rect -2378 3338 2266 3894
rect 2822 3338 38266 3894
rect 38822 3338 74266 3894
rect 74822 3338 110266 3894
rect 110822 3338 146266 3894
rect 146822 3338 182266 3894
rect 182822 3338 218266 3894
rect 218822 3338 254266 3894
rect 254822 3338 290266 3894
rect 290822 3338 326266 3894
rect 326822 3338 362266 3894
rect 362822 3338 398266 3894
rect 398822 3338 434266 3894
rect 434822 3338 470266 3894
rect 470822 3338 506266 3894
rect 506822 3338 542266 3894
rect 542822 3338 578266 3894
rect 578822 3338 586302 3894
rect 586858 3338 592650 3894
rect -8726 3306 592650 3338
rect -8726 2654 592650 2686
rect -8726 2098 -1974 2654
rect -1418 2098 1026 2654
rect 1582 2098 37026 2654
rect 37582 2098 73026 2654
rect 73582 2098 109026 2654
rect 109582 2098 145026 2654
rect 145582 2098 181026 2654
rect 181582 2098 217026 2654
rect 217582 2098 253026 2654
rect 253582 2098 289026 2654
rect 289582 2098 325026 2654
rect 325582 2098 361026 2654
rect 361582 2098 397026 2654
rect 397582 2098 433026 2654
rect 433582 2098 469026 2654
rect 469582 2098 505026 2654
rect 505582 2098 541026 2654
rect 541582 2098 577026 2654
rect 577582 2098 585342 2654
rect 585898 2098 592650 2654
rect -8726 2066 592650 2098
rect -2006 -346 585930 -314
rect -2006 -902 -1974 -346
rect -1418 -902 1026 -346
rect 1582 -902 37026 -346
rect 37582 -902 73026 -346
rect 73582 -902 109026 -346
rect 109582 -902 145026 -346
rect 145582 -902 181026 -346
rect 181582 -902 217026 -346
rect 217582 -902 253026 -346
rect 253582 -902 289026 -346
rect 289582 -902 325026 -346
rect 325582 -902 361026 -346
rect 361582 -902 397026 -346
rect 397582 -902 433026 -346
rect 433582 -902 469026 -346
rect 469582 -902 505026 -346
rect 505582 -902 541026 -346
rect 541582 -902 577026 -346
rect 577582 -902 585342 -346
rect 585898 -902 585930 -346
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1862 -2934 -1306
rect -2378 -1862 2266 -1306
rect 2822 -1862 38266 -1306
rect 38822 -1862 74266 -1306
rect 74822 -1862 110266 -1306
rect 110822 -1862 146266 -1306
rect 146822 -1862 182266 -1306
rect 182822 -1862 218266 -1306
rect 218822 -1862 254266 -1306
rect 254822 -1862 290266 -1306
rect 290822 -1862 326266 -1306
rect 326822 -1862 362266 -1306
rect 362822 -1862 398266 -1306
rect 398822 -1862 434266 -1306
rect 434822 -1862 470266 -1306
rect 470822 -1862 506266 -1306
rect 506822 -1862 542266 -1306
rect 542822 -1862 578266 -1306
rect 578822 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2822 -3894 -2266
rect -3338 -2822 3506 -2266
rect 4062 -2822 39506 -2266
rect 40062 -2822 75506 -2266
rect 76062 -2822 111506 -2266
rect 112062 -2822 147506 -2266
rect 148062 -2822 183506 -2266
rect 184062 -2822 219506 -2266
rect 220062 -2822 255506 -2266
rect 256062 -2822 291506 -2266
rect 292062 -2822 327506 -2266
rect 328062 -2822 363506 -2266
rect 364062 -2822 399506 -2266
rect 400062 -2822 435506 -2266
rect 436062 -2822 471506 -2266
rect 472062 -2822 507506 -2266
rect 508062 -2822 543506 -2266
rect 544062 -2822 579506 -2266
rect 580062 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3782 -4854 -3226
rect -4298 -3782 4746 -3226
rect 5302 -3782 40746 -3226
rect 41302 -3782 76746 -3226
rect 77302 -3782 112746 -3226
rect 113302 -3782 148746 -3226
rect 149302 -3782 184746 -3226
rect 185302 -3782 220746 -3226
rect 221302 -3782 256746 -3226
rect 257302 -3782 292746 -3226
rect 293302 -3782 328746 -3226
rect 329302 -3782 364746 -3226
rect 365302 -3782 400746 -3226
rect 401302 -3782 436746 -3226
rect 437302 -3782 472746 -3226
rect 473302 -3782 508746 -3226
rect 509302 -3782 544746 -3226
rect 545302 -3782 580746 -3226
rect 581302 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4742 -5814 -4186
rect -5258 -4742 5986 -4186
rect 6542 -4742 41986 -4186
rect 42542 -4742 77986 -4186
rect 78542 -4742 113986 -4186
rect 114542 -4742 149986 -4186
rect 150542 -4742 185986 -4186
rect 186542 -4742 221986 -4186
rect 222542 -4742 257986 -4186
rect 258542 -4742 293986 -4186
rect 294542 -4742 329986 -4186
rect 330542 -4742 365986 -4186
rect 366542 -4742 401986 -4186
rect 402542 -4742 437986 -4186
rect 438542 -4742 473986 -4186
rect 474542 -4742 509986 -4186
rect 510542 -4742 545986 -4186
rect 546542 -4742 581986 -4186
rect 582542 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5702 -6774 -5146
rect -6218 -5702 7226 -5146
rect 7782 -5702 43226 -5146
rect 43782 -5702 79226 -5146
rect 79782 -5702 115226 -5146
rect 115782 -5702 151226 -5146
rect 151782 -5702 187226 -5146
rect 187782 -5702 223226 -5146
rect 223782 -5702 259226 -5146
rect 259782 -5702 295226 -5146
rect 295782 -5702 331226 -5146
rect 331782 -5702 367226 -5146
rect 367782 -5702 403226 -5146
rect 403782 -5702 439226 -5146
rect 439782 -5702 475226 -5146
rect 475782 -5702 511226 -5146
rect 511782 -5702 547226 -5146
rect 547782 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6662 -7734 -6106
rect -7178 -6662 8466 -6106
rect 9022 -6662 44466 -6106
rect 45022 -6662 80466 -6106
rect 81022 -6662 116466 -6106
rect 117022 -6662 152466 -6106
rect 153022 -6662 188466 -6106
rect 189022 -6662 224466 -6106
rect 225022 -6662 260466 -6106
rect 261022 -6662 296466 -6106
rect 297022 -6662 332466 -6106
rect 333022 -6662 368466 -6106
rect 369022 -6662 404466 -6106
rect 405022 -6662 440466 -6106
rect 441022 -6662 476466 -6106
rect 477022 -6662 512466 -6106
rect 513022 -6662 548466 -6106
rect 549022 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7622 -8694 -7066
rect -8138 -7622 9706 -7066
rect 10262 -7622 45706 -7066
rect 46262 -7622 81706 -7066
rect 82262 -7622 117706 -7066
rect 118262 -7622 153706 -7066
rect 154262 -7622 189706 -7066
rect 190262 -7622 225706 -7066
rect 226262 -7622 261706 -7066
rect 262262 -7622 297706 -7066
rect 298262 -7622 333706 -7066
rect 334262 -7622 369706 -7066
rect 370262 -7622 405706 -7066
rect 406262 -7622 441706 -7066
rect 442262 -7622 477706 -7066
rect 478262 -7622 513706 -7066
rect 514262 -7622 549706 -7066
rect 550262 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect -8726 -7654 592650 -7622
use mux16x1_project  mprj1
timestamp 0
transform 1 0 538000 0 1 423800
box 0 552 10000 22000
use mux16x1_project  mprj2
timestamp 0
transform 1 0 538000 0 1 387800
box 0 552 10000 22000
use mux16x1_project  mprj3
timestamp 0
transform 1 0 538000 0 1 351800
box 0 552 10000 22000
use mux16x1_project  mprj4
timestamp 0
transform 1 0 538000 0 1 315800
box 0 552 10000 22000
use mux16x1_project  mprj5
timestamp 0
transform 1 0 538000 0 1 279800
box 0 552 10000 22000
use sky130_osu_ring_oscillator_mpr2ca_8_b0r1  ro1
timestamp 0
transform 1 0 468600 0 1 449000
box 0 0 20145 2491
use sky130_osu_ring_oscillator_mpr2ct_8_b0r1  ro2
timestamp 0
transform 1 0 468600 0 1 430600
box 0 0 20785 2492
use sky130_osu_ring_oscillator_mpr2ea_8_b0r1  ro3
timestamp 0
transform 1 0 468600 0 1 409600
box 0 0 19886 2492
use sky130_osu_ring_oscillator_mpr2et_8_b0r1  ro4
timestamp 0
transform 1 0 468600 0 1 388600
box 0 0 22123 2493
use sky130_osu_ring_oscillator_mpr2xa_8_b0r1  ro5
timestamp 0
transform 1 0 468600 0 1 367600
box 0 0 20809 2493
use sky130_osu_ring_oscillator_mpr2ca_8_b0r2  ro6
timestamp 0
transform 1 0 468600 0 1 346600
box 0 0 20217 2494
use sky130_osu_ring_oscillator_mpr2ct_8_b0r2  ro7
timestamp 0
transform 1 0 468600 0 1 325600
box 0 0 20783 2493
use sky130_osu_ring_oscillator_mpr2ea_8_b0r2  ro8
timestamp 0
transform 1 0 468600 0 1 304600
box 0 0 19885 2492
use sky130_osu_ring_oscillator_mpr2et_8_b0r2  ro9
timestamp 0
transform 1 0 468600 0 1 283600
box 0 0 22120 2493
use sky130_osu_ring_oscillator_mpr2xa_8_b0r2  ro10
timestamp 0
transform 1 0 468600 0 1 262600
box 0 0 20819 2493
use sky130_fd_sc_hd__conb_1  TIE_ZERO_zero_
timestamp 0
transform -1 0 544364 0 -1 213248
box -38 -48 314 592
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 1200 0 0 0 analog_io[0]
port 1 nsew
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 560 90 0 0 analog_io[10]
port 2 nsew
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 560 90 0 0 analog_io[11]
port 3 nsew
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 560 90 0 0 analog_io[12]
port 4 nsew
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 560 90 0 0 analog_io[13]
port 5 nsew
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 560 90 0 0 analog_io[14]
port 6 nsew
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 560 90 0 0 analog_io[15]
port 7 nsew
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 560 90 0 0 analog_io[16]
port 8 nsew
flabel metal3 s -960 697220 480 697460 0 FreeSans 1200 0 0 0 analog_io[17]
port 9 nsew
flabel metal3 s -960 644996 480 645236 0 FreeSans 1200 0 0 0 analog_io[18]
port 10 nsew
flabel metal3 s -960 592908 480 593148 0 FreeSans 1200 0 0 0 analog_io[19]
port 11 nsew
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 1200 0 0 0 analog_io[1]
port 12 nsew
flabel metal3 s -960 540684 480 540924 0 FreeSans 1200 0 0 0 analog_io[20]
port 13 nsew
flabel metal3 s -960 488596 480 488836 0 FreeSans 1200 0 0 0 analog_io[21]
port 14 nsew
flabel metal3 s -960 436508 480 436748 0 FreeSans 1200 0 0 0 analog_io[22]
port 15 nsew
flabel metal3 s -960 384284 480 384524 0 FreeSans 1200 0 0 0 analog_io[23]
port 16 nsew
flabel metal3 s -960 332196 480 332436 0 FreeSans 1200 0 0 0 analog_io[24]
port 17 nsew
flabel metal3 s -960 279972 480 280212 0 FreeSans 1200 0 0 0 analog_io[25]
port 18 nsew
flabel metal3 s -960 227884 480 228124 0 FreeSans 1200 0 0 0 analog_io[26]
port 19 nsew
flabel metal3 s -960 175796 480 176036 0 FreeSans 1200 0 0 0 analog_io[27]
port 20 nsew
flabel metal3 s -960 123572 480 123812 0 FreeSans 1200 0 0 0 analog_io[28]
port 21 nsew
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 1200 0 0 0 analog_io[2]
port 22 nsew
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 1200 0 0 0 analog_io[3]
port 23 nsew
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 1200 0 0 0 analog_io[4]
port 24 nsew
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 1200 0 0 0 analog_io[5]
port 25 nsew
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 1200 0 0 0 analog_io[6]
port 26 nsew
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 1200 0 0 0 analog_io[7]
port 27 nsew
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 560 90 0 0 analog_io[8]
port 28 nsew
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 560 90 0 0 analog_io[9]
port 29 nsew
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 1200 0 0 0 io_in[0]
port 30 nsew
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 1200 0 0 0 io_in[10]
port 31 nsew
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 1200 0 0 0 io_in[11]
port 32 nsew
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 1200 0 0 0 io_in[12]
port 33 nsew
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 1200 0 0 0 io_in[13]
port 34 nsew
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 1200 0 0 0 io_in[14]
port 35 nsew
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 560 90 0 0 io_in[15]
port 36 nsew
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 560 90 0 0 io_in[16]
port 37 nsew
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 560 90 0 0 io_in[17]
port 38 nsew
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 560 90 0 0 io_in[18]
port 39 nsew
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 560 90 0 0 io_in[19]
port 40 nsew
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 1200 0 0 0 io_in[1]
port 41 nsew
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 560 90 0 0 io_in[20]
port 42 nsew
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 560 90 0 0 io_in[21]
port 43 nsew
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 560 90 0 0 io_in[22]
port 44 nsew
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 560 90 0 0 io_in[23]
port 45 nsew
flabel metal3 s -960 684164 480 684404 0 FreeSans 1200 0 0 0 io_in[24]
port 46 nsew
flabel metal3 s -960 631940 480 632180 0 FreeSans 1200 0 0 0 io_in[25]
port 47 nsew
flabel metal3 s -960 579852 480 580092 0 FreeSans 1200 0 0 0 io_in[26]
port 48 nsew
flabel metal3 s -960 527764 480 528004 0 FreeSans 1200 0 0 0 io_in[27]
port 49 nsew
flabel metal3 s -960 475540 480 475780 0 FreeSans 1200 0 0 0 io_in[28]
port 50 nsew
flabel metal3 s -960 423452 480 423692 0 FreeSans 1200 0 0 0 io_in[29]
port 51 nsew
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 1200 0 0 0 io_in[2]
port 52 nsew
flabel metal3 s -960 371228 480 371468 0 FreeSans 1200 0 0 0 io_in[30]
port 53 nsew
flabel metal3 s -960 319140 480 319380 0 FreeSans 1200 0 0 0 io_in[31]
port 54 nsew
flabel metal3 s -960 267052 480 267292 0 FreeSans 1200 0 0 0 io_in[32]
port 55 nsew
flabel metal3 s -960 214828 480 215068 0 FreeSans 1200 0 0 0 io_in[33]
port 56 nsew
flabel metal3 s -960 162740 480 162980 0 FreeSans 1200 0 0 0 io_in[34]
port 57 nsew
flabel metal3 s -960 110516 480 110756 0 FreeSans 1200 0 0 0 io_in[35]
port 58 nsew
flabel metal3 s -960 71484 480 71724 0 FreeSans 1200 0 0 0 io_in[36]
port 59 nsew
flabel metal3 s -960 32316 480 32556 0 FreeSans 1200 0 0 0 io_in[37]
port 60 nsew
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 1200 0 0 0 io_in[3]
port 61 nsew
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 1200 0 0 0 io_in[4]
port 62 nsew
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 1200 0 0 0 io_in[5]
port 63 nsew
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 1200 0 0 0 io_in[6]
port 64 nsew
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 1200 0 0 0 io_in[7]
port 65 nsew
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 1200 0 0 0 io_in[8]
port 66 nsew
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 1200 0 0 0 io_in[9]
port 67 nsew
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 1200 0 0 0 io_oeb[0]
port 68 nsew
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 1200 0 0 0 io_oeb[10]
port 69 nsew
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 1200 0 0 0 io_oeb[11]
port 70 nsew
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 1200 0 0 0 io_oeb[12]
port 71 nsew
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 1200 0 0 0 io_oeb[13]
port 72 nsew
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 1200 0 0 0 io_oeb[14]
port 73 nsew
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 560 90 0 0 io_oeb[15]
port 74 nsew
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 560 90 0 0 io_oeb[16]
port 75 nsew
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 560 90 0 0 io_oeb[17]
port 76 nsew
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 560 90 0 0 io_oeb[18]
port 77 nsew
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 560 90 0 0 io_oeb[19]
port 78 nsew
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 1200 0 0 0 io_oeb[1]
port 79 nsew
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 560 90 0 0 io_oeb[20]
port 80 nsew
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 560 90 0 0 io_oeb[21]
port 81 nsew
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 560 90 0 0 io_oeb[22]
port 82 nsew
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 560 90 0 0 io_oeb[23]
port 83 nsew
flabel metal3 s -960 658052 480 658292 0 FreeSans 1200 0 0 0 io_oeb[24]
port 84 nsew
flabel metal3 s -960 605964 480 606204 0 FreeSans 1200 0 0 0 io_oeb[25]
port 85 nsew
flabel metal3 s -960 553740 480 553980 0 FreeSans 1200 0 0 0 io_oeb[26]
port 86 nsew
flabel metal3 s -960 501652 480 501892 0 FreeSans 1200 0 0 0 io_oeb[27]
port 87 nsew
flabel metal3 s -960 449428 480 449668 0 FreeSans 1200 0 0 0 io_oeb[28]
port 88 nsew
flabel metal3 s -960 397340 480 397580 0 FreeSans 1200 0 0 0 io_oeb[29]
port 89 nsew
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 1200 0 0 0 io_oeb[2]
port 90 nsew
flabel metal3 s -960 345252 480 345492 0 FreeSans 1200 0 0 0 io_oeb[30]
port 91 nsew
flabel metal3 s -960 293028 480 293268 0 FreeSans 1200 0 0 0 io_oeb[31]
port 92 nsew
flabel metal3 s -960 240940 480 241180 0 FreeSans 1200 0 0 0 io_oeb[32]
port 93 nsew
flabel metal3 s -960 188716 480 188956 0 FreeSans 1200 0 0 0 io_oeb[33]
port 94 nsew
flabel metal3 s -960 136628 480 136868 0 FreeSans 1200 0 0 0 io_oeb[34]
port 95 nsew
flabel metal3 s -960 84540 480 84780 0 FreeSans 1200 0 0 0 io_oeb[35]
port 96 nsew
flabel metal3 s -960 45372 480 45612 0 FreeSans 1200 0 0 0 io_oeb[36]
port 97 nsew
flabel metal3 s -960 6340 480 6580 0 FreeSans 1200 0 0 0 io_oeb[37]
port 98 nsew
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 1200 0 0 0 io_oeb[3]
port 99 nsew
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 1200 0 0 0 io_oeb[4]
port 100 nsew
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 1200 0 0 0 io_oeb[5]
port 101 nsew
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 1200 0 0 0 io_oeb[6]
port 102 nsew
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 1200 0 0 0 io_oeb[7]
port 103 nsew
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 1200 0 0 0 io_oeb[8]
port 104 nsew
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 1200 0 0 0 io_oeb[9]
port 105 nsew
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 1200 0 0 0 io_out[0]
port 106 nsew
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 1200 0 0 0 io_out[10]
port 107 nsew
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 1200 0 0 0 io_out[11]
port 108 nsew
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 1200 0 0 0 io_out[12]
port 109 nsew
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 1200 0 0 0 io_out[13]
port 110 nsew
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 1200 0 0 0 io_out[14]
port 111 nsew
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 560 90 0 0 io_out[15]
port 112 nsew
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 560 90 0 0 io_out[16]
port 113 nsew
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 560 90 0 0 io_out[17]
port 114 nsew
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 560 90 0 0 io_out[18]
port 115 nsew
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 560 90 0 0 io_out[19]
port 116 nsew
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 1200 0 0 0 io_out[1]
port 117 nsew
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 560 90 0 0 io_out[20]
port 118 nsew
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 560 90 0 0 io_out[21]
port 119 nsew
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 560 90 0 0 io_out[22]
port 120 nsew
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 560 90 0 0 io_out[23]
port 121 nsew
flabel metal3 s -960 671108 480 671348 0 FreeSans 1200 0 0 0 io_out[24]
port 122 nsew
flabel metal3 s -960 619020 480 619260 0 FreeSans 1200 0 0 0 io_out[25]
port 123 nsew
flabel metal3 s -960 566796 480 567036 0 FreeSans 1200 0 0 0 io_out[26]
port 124 nsew
flabel metal3 s -960 514708 480 514948 0 FreeSans 1200 0 0 0 io_out[27]
port 125 nsew
flabel metal3 s -960 462484 480 462724 0 FreeSans 1200 0 0 0 io_out[28]
port 126 nsew
flabel metal3 s -960 410396 480 410636 0 FreeSans 1200 0 0 0 io_out[29]
port 127 nsew
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 1200 0 0 0 io_out[2]
port 128 nsew
flabel metal3 s -960 358308 480 358548 0 FreeSans 1200 0 0 0 io_out[30]
port 129 nsew
flabel metal3 s -960 306084 480 306324 0 FreeSans 1200 0 0 0 io_out[31]
port 130 nsew
flabel metal3 s -960 253996 480 254236 0 FreeSans 1200 0 0 0 io_out[32]
port 131 nsew
flabel metal3 s -960 201772 480 202012 0 FreeSans 1200 0 0 0 io_out[33]
port 132 nsew
flabel metal3 s -960 149684 480 149924 0 FreeSans 1200 0 0 0 io_out[34]
port 133 nsew
flabel metal3 s -960 97460 480 97700 0 FreeSans 1200 0 0 0 io_out[35]
port 134 nsew
flabel metal3 s -960 58428 480 58668 0 FreeSans 1200 0 0 0 io_out[36]
port 135 nsew
flabel metal3 s -960 19260 480 19500 0 FreeSans 1200 0 0 0 io_out[37]
port 136 nsew
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 1200 0 0 0 io_out[3]
port 137 nsew
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 1200 0 0 0 io_out[4]
port 138 nsew
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 1200 0 0 0 io_out[5]
port 139 nsew
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 1200 0 0 0 io_out[6]
port 140 nsew
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 1200 0 0 0 io_out[7]
port 141 nsew
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 1200 0 0 0 io_out[8]
port 142 nsew
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 1200 0 0 0 io_out[9]
port 143 nsew
flabel metal2 s 125846 -960 125958 480 0 FreeSans 560 90 0 0 la_data_in[0]
port 144 nsew
flabel metal2 s 480506 -960 480618 480 0 FreeSans 560 90 0 0 la_data_in[100]
port 145 nsew
flabel metal2 s 484002 -960 484114 480 0 FreeSans 560 90 0 0 la_data_in[101]
port 146 nsew
flabel metal2 s 487590 -960 487702 480 0 FreeSans 560 90 0 0 la_data_in[102]
port 147 nsew
flabel metal2 s 491086 -960 491198 480 0 FreeSans 560 90 0 0 la_data_in[103]
port 148 nsew
flabel metal2 s 494674 -960 494786 480 0 FreeSans 560 90 0 0 la_data_in[104]
port 149 nsew
flabel metal2 s 498170 -960 498282 480 0 FreeSans 560 90 0 0 la_data_in[105]
port 150 nsew
flabel metal2 s 501758 -960 501870 480 0 FreeSans 560 90 0 0 la_data_in[106]
port 151 nsew
flabel metal2 s 505346 -960 505458 480 0 FreeSans 560 90 0 0 la_data_in[107]
port 152 nsew
flabel metal2 s 508842 -960 508954 480 0 FreeSans 560 90 0 0 la_data_in[108]
port 153 nsew
flabel metal2 s 512430 -960 512542 480 0 FreeSans 560 90 0 0 la_data_in[109]
port 154 nsew
flabel metal2 s 161266 -960 161378 480 0 FreeSans 560 90 0 0 la_data_in[10]
port 155 nsew
flabel metal2 s 515926 -960 516038 480 0 FreeSans 560 90 0 0 la_data_in[110]
port 156 nsew
flabel metal2 s 519514 -960 519626 480 0 FreeSans 560 90 0 0 la_data_in[111]
port 157 nsew
flabel metal2 s 523010 -960 523122 480 0 FreeSans 560 90 0 0 la_data_in[112]
port 158 nsew
flabel metal2 s 526598 -960 526710 480 0 FreeSans 560 90 0 0 la_data_in[113]
port 159 nsew
flabel metal2 s 530094 -960 530206 480 0 FreeSans 560 90 0 0 la_data_in[114]
port 160 nsew
flabel metal2 s 533682 -960 533794 480 0 FreeSans 560 90 0 0 la_data_in[115]
port 161 nsew
flabel metal2 s 537178 -960 537290 480 0 FreeSans 560 90 0 0 la_data_in[116]
port 162 nsew
flabel metal2 s 540766 -960 540878 480 0 FreeSans 560 90 0 0 la_data_in[117]
port 163 nsew
flabel metal2 s 544354 -960 544466 480 0 FreeSans 560 90 0 0 la_data_in[118]
port 164 nsew
flabel metal2 s 547850 -960 547962 480 0 FreeSans 560 90 0 0 la_data_in[119]
port 165 nsew
flabel metal2 s 164854 -960 164966 480 0 FreeSans 560 90 0 0 la_data_in[11]
port 166 nsew
flabel metal2 s 551438 -960 551550 480 0 FreeSans 560 90 0 0 la_data_in[120]
port 167 nsew
flabel metal2 s 554934 -960 555046 480 0 FreeSans 560 90 0 0 la_data_in[121]
port 168 nsew
flabel metal2 s 558522 -960 558634 480 0 FreeSans 560 90 0 0 la_data_in[122]
port 169 nsew
flabel metal2 s 562018 -960 562130 480 0 FreeSans 560 90 0 0 la_data_in[123]
port 170 nsew
flabel metal2 s 565606 -960 565718 480 0 FreeSans 560 90 0 0 la_data_in[124]
port 171 nsew
flabel metal2 s 569102 -960 569214 480 0 FreeSans 560 90 0 0 la_data_in[125]
port 172 nsew
flabel metal2 s 572690 -960 572802 480 0 FreeSans 560 90 0 0 la_data_in[126]
port 173 nsew
flabel metal2 s 576278 -960 576390 480 0 FreeSans 560 90 0 0 la_data_in[127]
port 174 nsew
flabel metal2 s 168350 -960 168462 480 0 FreeSans 560 90 0 0 la_data_in[12]
port 175 nsew
flabel metal2 s 171938 -960 172050 480 0 FreeSans 560 90 0 0 la_data_in[13]
port 176 nsew
flabel metal2 s 175434 -960 175546 480 0 FreeSans 560 90 0 0 la_data_in[14]
port 177 nsew
flabel metal2 s 179022 -960 179134 480 0 FreeSans 560 90 0 0 la_data_in[15]
port 178 nsew
flabel metal2 s 182518 -960 182630 480 0 FreeSans 560 90 0 0 la_data_in[16]
port 179 nsew
flabel metal2 s 186106 -960 186218 480 0 FreeSans 560 90 0 0 la_data_in[17]
port 180 nsew
flabel metal2 s 189694 -960 189806 480 0 FreeSans 560 90 0 0 la_data_in[18]
port 181 nsew
flabel metal2 s 193190 -960 193302 480 0 FreeSans 560 90 0 0 la_data_in[19]
port 182 nsew
flabel metal2 s 129342 -960 129454 480 0 FreeSans 560 90 0 0 la_data_in[1]
port 183 nsew
flabel metal2 s 196778 -960 196890 480 0 FreeSans 560 90 0 0 la_data_in[20]
port 184 nsew
flabel metal2 s 200274 -960 200386 480 0 FreeSans 560 90 0 0 la_data_in[21]
port 185 nsew
flabel metal2 s 203862 -960 203974 480 0 FreeSans 560 90 0 0 la_data_in[22]
port 186 nsew
flabel metal2 s 207358 -960 207470 480 0 FreeSans 560 90 0 0 la_data_in[23]
port 187 nsew
flabel metal2 s 210946 -960 211058 480 0 FreeSans 560 90 0 0 la_data_in[24]
port 188 nsew
flabel metal2 s 214442 -960 214554 480 0 FreeSans 560 90 0 0 la_data_in[25]
port 189 nsew
flabel metal2 s 218030 -960 218142 480 0 FreeSans 560 90 0 0 la_data_in[26]
port 190 nsew
flabel metal2 s 221526 -960 221638 480 0 FreeSans 560 90 0 0 la_data_in[27]
port 191 nsew
flabel metal2 s 225114 -960 225226 480 0 FreeSans 560 90 0 0 la_data_in[28]
port 192 nsew
flabel metal2 s 228702 -960 228814 480 0 FreeSans 560 90 0 0 la_data_in[29]
port 193 nsew
flabel metal2 s 132930 -960 133042 480 0 FreeSans 560 90 0 0 la_data_in[2]
port 194 nsew
flabel metal2 s 232198 -960 232310 480 0 FreeSans 560 90 0 0 la_data_in[30]
port 195 nsew
flabel metal2 s 235786 -960 235898 480 0 FreeSans 560 90 0 0 la_data_in[31]
port 196 nsew
flabel metal2 s 239282 -960 239394 480 0 FreeSans 560 90 0 0 la_data_in[32]
port 197 nsew
flabel metal2 s 242870 -960 242982 480 0 FreeSans 560 90 0 0 la_data_in[33]
port 198 nsew
flabel metal2 s 246366 -960 246478 480 0 FreeSans 560 90 0 0 la_data_in[34]
port 199 nsew
flabel metal2 s 249954 -960 250066 480 0 FreeSans 560 90 0 0 la_data_in[35]
port 200 nsew
flabel metal2 s 253450 -960 253562 480 0 FreeSans 560 90 0 0 la_data_in[36]
port 201 nsew
flabel metal2 s 257038 -960 257150 480 0 FreeSans 560 90 0 0 la_data_in[37]
port 202 nsew
flabel metal2 s 260626 -960 260738 480 0 FreeSans 560 90 0 0 la_data_in[38]
port 203 nsew
flabel metal2 s 264122 -960 264234 480 0 FreeSans 560 90 0 0 la_data_in[39]
port 204 nsew
flabel metal2 s 136426 -960 136538 480 0 FreeSans 560 90 0 0 la_data_in[3]
port 205 nsew
flabel metal2 s 267710 -960 267822 480 0 FreeSans 560 90 0 0 la_data_in[40]
port 206 nsew
flabel metal2 s 271206 -960 271318 480 0 FreeSans 560 90 0 0 la_data_in[41]
port 207 nsew
flabel metal2 s 274794 -960 274906 480 0 FreeSans 560 90 0 0 la_data_in[42]
port 208 nsew
flabel metal2 s 278290 -960 278402 480 0 FreeSans 560 90 0 0 la_data_in[43]
port 209 nsew
flabel metal2 s 281878 -960 281990 480 0 FreeSans 560 90 0 0 la_data_in[44]
port 210 nsew
flabel metal2 s 285374 -960 285486 480 0 FreeSans 560 90 0 0 la_data_in[45]
port 211 nsew
flabel metal2 s 288962 -960 289074 480 0 FreeSans 560 90 0 0 la_data_in[46]
port 212 nsew
flabel metal2 s 292550 -960 292662 480 0 FreeSans 560 90 0 0 la_data_in[47]
port 213 nsew
flabel metal2 s 296046 -960 296158 480 0 FreeSans 560 90 0 0 la_data_in[48]
port 214 nsew
flabel metal2 s 299634 -960 299746 480 0 FreeSans 560 90 0 0 la_data_in[49]
port 215 nsew
flabel metal2 s 140014 -960 140126 480 0 FreeSans 560 90 0 0 la_data_in[4]
port 216 nsew
flabel metal2 s 303130 -960 303242 480 0 FreeSans 560 90 0 0 la_data_in[50]
port 217 nsew
flabel metal2 s 306718 -960 306830 480 0 FreeSans 560 90 0 0 la_data_in[51]
port 218 nsew
flabel metal2 s 310214 -960 310326 480 0 FreeSans 560 90 0 0 la_data_in[52]
port 219 nsew
flabel metal2 s 313802 -960 313914 480 0 FreeSans 560 90 0 0 la_data_in[53]
port 220 nsew
flabel metal2 s 317298 -960 317410 480 0 FreeSans 560 90 0 0 la_data_in[54]
port 221 nsew
flabel metal2 s 320886 -960 320998 480 0 FreeSans 560 90 0 0 la_data_in[55]
port 222 nsew
flabel metal2 s 324382 -960 324494 480 0 FreeSans 560 90 0 0 la_data_in[56]
port 223 nsew
flabel metal2 s 327970 -960 328082 480 0 FreeSans 560 90 0 0 la_data_in[57]
port 224 nsew
flabel metal2 s 331558 -960 331670 480 0 FreeSans 560 90 0 0 la_data_in[58]
port 225 nsew
flabel metal2 s 335054 -960 335166 480 0 FreeSans 560 90 0 0 la_data_in[59]
port 226 nsew
flabel metal2 s 143510 -960 143622 480 0 FreeSans 560 90 0 0 la_data_in[5]
port 227 nsew
flabel metal2 s 338642 -960 338754 480 0 FreeSans 560 90 0 0 la_data_in[60]
port 228 nsew
flabel metal2 s 342138 -960 342250 480 0 FreeSans 560 90 0 0 la_data_in[61]
port 229 nsew
flabel metal2 s 345726 -960 345838 480 0 FreeSans 560 90 0 0 la_data_in[62]
port 230 nsew
flabel metal2 s 349222 -960 349334 480 0 FreeSans 560 90 0 0 la_data_in[63]
port 231 nsew
flabel metal2 s 352810 -960 352922 480 0 FreeSans 560 90 0 0 la_data_in[64]
port 232 nsew
flabel metal2 s 356306 -960 356418 480 0 FreeSans 560 90 0 0 la_data_in[65]
port 233 nsew
flabel metal2 s 359894 -960 360006 480 0 FreeSans 560 90 0 0 la_data_in[66]
port 234 nsew
flabel metal2 s 363482 -960 363594 480 0 FreeSans 560 90 0 0 la_data_in[67]
port 235 nsew
flabel metal2 s 366978 -960 367090 480 0 FreeSans 560 90 0 0 la_data_in[68]
port 236 nsew
flabel metal2 s 370566 -960 370678 480 0 FreeSans 560 90 0 0 la_data_in[69]
port 237 nsew
flabel metal2 s 147098 -960 147210 480 0 FreeSans 560 90 0 0 la_data_in[6]
port 238 nsew
flabel metal2 s 374062 -960 374174 480 0 FreeSans 560 90 0 0 la_data_in[70]
port 239 nsew
flabel metal2 s 377650 -960 377762 480 0 FreeSans 560 90 0 0 la_data_in[71]
port 240 nsew
flabel metal2 s 381146 -960 381258 480 0 FreeSans 560 90 0 0 la_data_in[72]
port 241 nsew
flabel metal2 s 384734 -960 384846 480 0 FreeSans 560 90 0 0 la_data_in[73]
port 242 nsew
flabel metal2 s 388230 -960 388342 480 0 FreeSans 560 90 0 0 la_data_in[74]
port 243 nsew
flabel metal2 s 391818 -960 391930 480 0 FreeSans 560 90 0 0 la_data_in[75]
port 244 nsew
flabel metal2 s 395314 -960 395426 480 0 FreeSans 560 90 0 0 la_data_in[76]
port 245 nsew
flabel metal2 s 398902 -960 399014 480 0 FreeSans 560 90 0 0 la_data_in[77]
port 246 nsew
flabel metal2 s 402490 -960 402602 480 0 FreeSans 560 90 0 0 la_data_in[78]
port 247 nsew
flabel metal2 s 405986 -960 406098 480 0 FreeSans 560 90 0 0 la_data_in[79]
port 248 nsew
flabel metal2 s 150594 -960 150706 480 0 FreeSans 560 90 0 0 la_data_in[7]
port 249 nsew
flabel metal2 s 409574 -960 409686 480 0 FreeSans 560 90 0 0 la_data_in[80]
port 250 nsew
flabel metal2 s 413070 -960 413182 480 0 FreeSans 560 90 0 0 la_data_in[81]
port 251 nsew
flabel metal2 s 416658 -960 416770 480 0 FreeSans 560 90 0 0 la_data_in[82]
port 252 nsew
flabel metal2 s 420154 -960 420266 480 0 FreeSans 560 90 0 0 la_data_in[83]
port 253 nsew
flabel metal2 s 423742 -960 423854 480 0 FreeSans 560 90 0 0 la_data_in[84]
port 254 nsew
flabel metal2 s 427238 -960 427350 480 0 FreeSans 560 90 0 0 la_data_in[85]
port 255 nsew
flabel metal2 s 430826 -960 430938 480 0 FreeSans 560 90 0 0 la_data_in[86]
port 256 nsew
flabel metal2 s 434414 -960 434526 480 0 FreeSans 560 90 0 0 la_data_in[87]
port 257 nsew
flabel metal2 s 437910 -960 438022 480 0 FreeSans 560 90 0 0 la_data_in[88]
port 258 nsew
flabel metal2 s 441498 -960 441610 480 0 FreeSans 560 90 0 0 la_data_in[89]
port 259 nsew
flabel metal2 s 154182 -960 154294 480 0 FreeSans 560 90 0 0 la_data_in[8]
port 260 nsew
flabel metal2 s 444994 -960 445106 480 0 FreeSans 560 90 0 0 la_data_in[90]
port 261 nsew
flabel metal2 s 448582 -960 448694 480 0 FreeSans 560 90 0 0 la_data_in[91]
port 262 nsew
flabel metal2 s 452078 -960 452190 480 0 FreeSans 560 90 0 0 la_data_in[92]
port 263 nsew
flabel metal2 s 455666 -960 455778 480 0 FreeSans 560 90 0 0 la_data_in[93]
port 264 nsew
flabel metal2 s 459162 -960 459274 480 0 FreeSans 560 90 0 0 la_data_in[94]
port 265 nsew
flabel metal2 s 462750 -960 462862 480 0 FreeSans 560 90 0 0 la_data_in[95]
port 266 nsew
flabel metal2 s 466246 -960 466358 480 0 FreeSans 560 90 0 0 la_data_in[96]
port 267 nsew
flabel metal2 s 469834 -960 469946 480 0 FreeSans 560 90 0 0 la_data_in[97]
port 268 nsew
flabel metal2 s 473422 -960 473534 480 0 FreeSans 560 90 0 0 la_data_in[98]
port 269 nsew
flabel metal2 s 476918 -960 477030 480 0 FreeSans 560 90 0 0 la_data_in[99]
port 270 nsew
flabel metal2 s 157770 -960 157882 480 0 FreeSans 560 90 0 0 la_data_in[9]
port 271 nsew
flabel metal2 s 126950 -960 127062 480 0 FreeSans 560 90 0 0 la_data_out[0]
port 272 nsew
flabel metal2 s 481702 -960 481814 480 0 FreeSans 560 90 0 0 la_data_out[100]
port 273 nsew
flabel metal2 s 485198 -960 485310 480 0 FreeSans 560 90 0 0 la_data_out[101]
port 274 nsew
flabel metal2 s 488786 -960 488898 480 0 FreeSans 560 90 0 0 la_data_out[102]
port 275 nsew
flabel metal2 s 492282 -960 492394 480 0 FreeSans 560 90 0 0 la_data_out[103]
port 276 nsew
flabel metal2 s 495870 -960 495982 480 0 FreeSans 560 90 0 0 la_data_out[104]
port 277 nsew
flabel metal2 s 499366 -960 499478 480 0 FreeSans 560 90 0 0 la_data_out[105]
port 278 nsew
flabel metal2 s 502954 -960 503066 480 0 FreeSans 560 90 0 0 la_data_out[106]
port 279 nsew
flabel metal2 s 506450 -960 506562 480 0 FreeSans 560 90 0 0 la_data_out[107]
port 280 nsew
flabel metal2 s 510038 -960 510150 480 0 FreeSans 560 90 0 0 la_data_out[108]
port 281 nsew
flabel metal2 s 513534 -960 513646 480 0 FreeSans 560 90 0 0 la_data_out[109]
port 282 nsew
flabel metal2 s 162462 -960 162574 480 0 FreeSans 560 90 0 0 la_data_out[10]
port 283 nsew
flabel metal2 s 517122 -960 517234 480 0 FreeSans 560 90 0 0 la_data_out[110]
port 284 nsew
flabel metal2 s 520710 -960 520822 480 0 FreeSans 560 90 0 0 la_data_out[111]
port 285 nsew
flabel metal2 s 524206 -960 524318 480 0 FreeSans 560 90 0 0 la_data_out[112]
port 286 nsew
flabel metal2 s 527794 -960 527906 480 0 FreeSans 560 90 0 0 la_data_out[113]
port 287 nsew
flabel metal2 s 531290 -960 531402 480 0 FreeSans 560 90 0 0 la_data_out[114]
port 288 nsew
flabel metal2 s 534878 -960 534990 480 0 FreeSans 560 90 0 0 la_data_out[115]
port 289 nsew
flabel metal2 s 538374 -960 538486 480 0 FreeSans 560 90 0 0 la_data_out[116]
port 290 nsew
flabel metal2 s 541962 -960 542074 480 0 FreeSans 560 90 0 0 la_data_out[117]
port 291 nsew
flabel metal2 s 545458 -960 545570 480 0 FreeSans 560 90 0 0 la_data_out[118]
port 292 nsew
flabel metal2 s 549046 -960 549158 480 0 FreeSans 560 90 0 0 la_data_out[119]
port 293 nsew
flabel metal2 s 166050 -960 166162 480 0 FreeSans 560 90 0 0 la_data_out[11]
port 294 nsew
flabel metal2 s 552634 -960 552746 480 0 FreeSans 560 90 0 0 la_data_out[120]
port 295 nsew
flabel metal2 s 556130 -960 556242 480 0 FreeSans 560 90 0 0 la_data_out[121]
port 296 nsew
flabel metal2 s 559718 -960 559830 480 0 FreeSans 560 90 0 0 la_data_out[122]
port 297 nsew
flabel metal2 s 563214 -960 563326 480 0 FreeSans 560 90 0 0 la_data_out[123]
port 298 nsew
flabel metal2 s 566802 -960 566914 480 0 FreeSans 560 90 0 0 la_data_out[124]
port 299 nsew
flabel metal2 s 570298 -960 570410 480 0 FreeSans 560 90 0 0 la_data_out[125]
port 300 nsew
flabel metal2 s 573886 -960 573998 480 0 FreeSans 560 90 0 0 la_data_out[126]
port 301 nsew
flabel metal2 s 577382 -960 577494 480 0 FreeSans 560 90 0 0 la_data_out[127]
port 302 nsew
flabel metal2 s 169546 -960 169658 480 0 FreeSans 560 90 0 0 la_data_out[12]
port 303 nsew
flabel metal2 s 173134 -960 173246 480 0 FreeSans 560 90 0 0 la_data_out[13]
port 304 nsew
flabel metal2 s 176630 -960 176742 480 0 FreeSans 560 90 0 0 la_data_out[14]
port 305 nsew
flabel metal2 s 180218 -960 180330 480 0 FreeSans 560 90 0 0 la_data_out[15]
port 306 nsew
flabel metal2 s 183714 -960 183826 480 0 FreeSans 560 90 0 0 la_data_out[16]
port 307 nsew
flabel metal2 s 187302 -960 187414 480 0 FreeSans 560 90 0 0 la_data_out[17]
port 308 nsew
flabel metal2 s 190798 -960 190910 480 0 FreeSans 560 90 0 0 la_data_out[18]
port 309 nsew
flabel metal2 s 194386 -960 194498 480 0 FreeSans 560 90 0 0 la_data_out[19]
port 310 nsew
flabel metal2 s 130538 -960 130650 480 0 FreeSans 560 90 0 0 la_data_out[1]
port 311 nsew
flabel metal2 s 197882 -960 197994 480 0 FreeSans 560 90 0 0 la_data_out[20]
port 312 nsew
flabel metal2 s 201470 -960 201582 480 0 FreeSans 560 90 0 0 la_data_out[21]
port 313 nsew
flabel metal2 s 205058 -960 205170 480 0 FreeSans 560 90 0 0 la_data_out[22]
port 314 nsew
flabel metal2 s 208554 -960 208666 480 0 FreeSans 560 90 0 0 la_data_out[23]
port 315 nsew
flabel metal2 s 212142 -960 212254 480 0 FreeSans 560 90 0 0 la_data_out[24]
port 316 nsew
flabel metal2 s 215638 -960 215750 480 0 FreeSans 560 90 0 0 la_data_out[25]
port 317 nsew
flabel metal2 s 219226 -960 219338 480 0 FreeSans 560 90 0 0 la_data_out[26]
port 318 nsew
flabel metal2 s 222722 -960 222834 480 0 FreeSans 560 90 0 0 la_data_out[27]
port 319 nsew
flabel metal2 s 226310 -960 226422 480 0 FreeSans 560 90 0 0 la_data_out[28]
port 320 nsew
flabel metal2 s 229806 -960 229918 480 0 FreeSans 560 90 0 0 la_data_out[29]
port 321 nsew
flabel metal2 s 134126 -960 134238 480 0 FreeSans 560 90 0 0 la_data_out[2]
port 322 nsew
flabel metal2 s 233394 -960 233506 480 0 FreeSans 560 90 0 0 la_data_out[30]
port 323 nsew
flabel metal2 s 236982 -960 237094 480 0 FreeSans 560 90 0 0 la_data_out[31]
port 324 nsew
flabel metal2 s 240478 -960 240590 480 0 FreeSans 560 90 0 0 la_data_out[32]
port 325 nsew
flabel metal2 s 244066 -960 244178 480 0 FreeSans 560 90 0 0 la_data_out[33]
port 326 nsew
flabel metal2 s 247562 -960 247674 480 0 FreeSans 560 90 0 0 la_data_out[34]
port 327 nsew
flabel metal2 s 251150 -960 251262 480 0 FreeSans 560 90 0 0 la_data_out[35]
port 328 nsew
flabel metal2 s 254646 -960 254758 480 0 FreeSans 560 90 0 0 la_data_out[36]
port 329 nsew
flabel metal2 s 258234 -960 258346 480 0 FreeSans 560 90 0 0 la_data_out[37]
port 330 nsew
flabel metal2 s 261730 -960 261842 480 0 FreeSans 560 90 0 0 la_data_out[38]
port 331 nsew
flabel metal2 s 265318 -960 265430 480 0 FreeSans 560 90 0 0 la_data_out[39]
port 332 nsew
flabel metal2 s 137622 -960 137734 480 0 FreeSans 560 90 0 0 la_data_out[3]
port 333 nsew
flabel metal2 s 268814 -960 268926 480 0 FreeSans 560 90 0 0 la_data_out[40]
port 334 nsew
flabel metal2 s 272402 -960 272514 480 0 FreeSans 560 90 0 0 la_data_out[41]
port 335 nsew
flabel metal2 s 275990 -960 276102 480 0 FreeSans 560 90 0 0 la_data_out[42]
port 336 nsew
flabel metal2 s 279486 -960 279598 480 0 FreeSans 560 90 0 0 la_data_out[43]
port 337 nsew
flabel metal2 s 283074 -960 283186 480 0 FreeSans 560 90 0 0 la_data_out[44]
port 338 nsew
flabel metal2 s 286570 -960 286682 480 0 FreeSans 560 90 0 0 la_data_out[45]
port 339 nsew
flabel metal2 s 290158 -960 290270 480 0 FreeSans 560 90 0 0 la_data_out[46]
port 340 nsew
flabel metal2 s 293654 -960 293766 480 0 FreeSans 560 90 0 0 la_data_out[47]
port 341 nsew
flabel metal2 s 297242 -960 297354 480 0 FreeSans 560 90 0 0 la_data_out[48]
port 342 nsew
flabel metal2 s 300738 -960 300850 480 0 FreeSans 560 90 0 0 la_data_out[49]
port 343 nsew
flabel metal2 s 141210 -960 141322 480 0 FreeSans 560 90 0 0 la_data_out[4]
port 344 nsew
flabel metal2 s 304326 -960 304438 480 0 FreeSans 560 90 0 0 la_data_out[50]
port 345 nsew
flabel metal2 s 307914 -960 308026 480 0 FreeSans 560 90 0 0 la_data_out[51]
port 346 nsew
flabel metal2 s 311410 -960 311522 480 0 FreeSans 560 90 0 0 la_data_out[52]
port 347 nsew
flabel metal2 s 314998 -960 315110 480 0 FreeSans 560 90 0 0 la_data_out[53]
port 348 nsew
flabel metal2 s 318494 -960 318606 480 0 FreeSans 560 90 0 0 la_data_out[54]
port 349 nsew
flabel metal2 s 322082 -960 322194 480 0 FreeSans 560 90 0 0 la_data_out[55]
port 350 nsew
flabel metal2 s 325578 -960 325690 480 0 FreeSans 560 90 0 0 la_data_out[56]
port 351 nsew
flabel metal2 s 329166 -960 329278 480 0 FreeSans 560 90 0 0 la_data_out[57]
port 352 nsew
flabel metal2 s 332662 -960 332774 480 0 FreeSans 560 90 0 0 la_data_out[58]
port 353 nsew
flabel metal2 s 336250 -960 336362 480 0 FreeSans 560 90 0 0 la_data_out[59]
port 354 nsew
flabel metal2 s 144706 -960 144818 480 0 FreeSans 560 90 0 0 la_data_out[5]
port 355 nsew
flabel metal2 s 339838 -960 339950 480 0 FreeSans 560 90 0 0 la_data_out[60]
port 356 nsew
flabel metal2 s 343334 -960 343446 480 0 FreeSans 560 90 0 0 la_data_out[61]
port 357 nsew
flabel metal2 s 346922 -960 347034 480 0 FreeSans 560 90 0 0 la_data_out[62]
port 358 nsew
flabel metal2 s 350418 -960 350530 480 0 FreeSans 560 90 0 0 la_data_out[63]
port 359 nsew
flabel metal2 s 354006 -960 354118 480 0 FreeSans 560 90 0 0 la_data_out[64]
port 360 nsew
flabel metal2 s 357502 -960 357614 480 0 FreeSans 560 90 0 0 la_data_out[65]
port 361 nsew
flabel metal2 s 361090 -960 361202 480 0 FreeSans 560 90 0 0 la_data_out[66]
port 362 nsew
flabel metal2 s 364586 -960 364698 480 0 FreeSans 560 90 0 0 la_data_out[67]
port 363 nsew
flabel metal2 s 368174 -960 368286 480 0 FreeSans 560 90 0 0 la_data_out[68]
port 364 nsew
flabel metal2 s 371670 -960 371782 480 0 FreeSans 560 90 0 0 la_data_out[69]
port 365 nsew
flabel metal2 s 148294 -960 148406 480 0 FreeSans 560 90 0 0 la_data_out[6]
port 366 nsew
flabel metal2 s 375258 -960 375370 480 0 FreeSans 560 90 0 0 la_data_out[70]
port 367 nsew
flabel metal2 s 378846 -960 378958 480 0 FreeSans 560 90 0 0 la_data_out[71]
port 368 nsew
flabel metal2 s 382342 -960 382454 480 0 FreeSans 560 90 0 0 la_data_out[72]
port 369 nsew
flabel metal2 s 385930 -960 386042 480 0 FreeSans 560 90 0 0 la_data_out[73]
port 370 nsew
flabel metal2 s 389426 -960 389538 480 0 FreeSans 560 90 0 0 la_data_out[74]
port 371 nsew
flabel metal2 s 393014 -960 393126 480 0 FreeSans 560 90 0 0 la_data_out[75]
port 372 nsew
flabel metal2 s 396510 -960 396622 480 0 FreeSans 560 90 0 0 la_data_out[76]
port 373 nsew
flabel metal2 s 400098 -960 400210 480 0 FreeSans 560 90 0 0 la_data_out[77]
port 374 nsew
flabel metal2 s 403594 -960 403706 480 0 FreeSans 560 90 0 0 la_data_out[78]
port 375 nsew
flabel metal2 s 407182 -960 407294 480 0 FreeSans 560 90 0 0 la_data_out[79]
port 376 nsew
flabel metal2 s 151790 -960 151902 480 0 FreeSans 560 90 0 0 la_data_out[7]
port 377 nsew
flabel metal2 s 410770 -960 410882 480 0 FreeSans 560 90 0 0 la_data_out[80]
port 378 nsew
flabel metal2 s 414266 -960 414378 480 0 FreeSans 560 90 0 0 la_data_out[81]
port 379 nsew
flabel metal2 s 417854 -960 417966 480 0 FreeSans 560 90 0 0 la_data_out[82]
port 380 nsew
flabel metal2 s 421350 -960 421462 480 0 FreeSans 560 90 0 0 la_data_out[83]
port 381 nsew
flabel metal2 s 424938 -960 425050 480 0 FreeSans 560 90 0 0 la_data_out[84]
port 382 nsew
flabel metal2 s 428434 -960 428546 480 0 FreeSans 560 90 0 0 la_data_out[85]
port 383 nsew
flabel metal2 s 432022 -960 432134 480 0 FreeSans 560 90 0 0 la_data_out[86]
port 384 nsew
flabel metal2 s 435518 -960 435630 480 0 FreeSans 560 90 0 0 la_data_out[87]
port 385 nsew
flabel metal2 s 439106 -960 439218 480 0 FreeSans 560 90 0 0 la_data_out[88]
port 386 nsew
flabel metal2 s 442602 -960 442714 480 0 FreeSans 560 90 0 0 la_data_out[89]
port 387 nsew
flabel metal2 s 155378 -960 155490 480 0 FreeSans 560 90 0 0 la_data_out[8]
port 388 nsew
flabel metal2 s 446190 -960 446302 480 0 FreeSans 560 90 0 0 la_data_out[90]
port 389 nsew
flabel metal2 s 449778 -960 449890 480 0 FreeSans 560 90 0 0 la_data_out[91]
port 390 nsew
flabel metal2 s 453274 -960 453386 480 0 FreeSans 560 90 0 0 la_data_out[92]
port 391 nsew
flabel metal2 s 456862 -960 456974 480 0 FreeSans 560 90 0 0 la_data_out[93]
port 392 nsew
flabel metal2 s 460358 -960 460470 480 0 FreeSans 560 90 0 0 la_data_out[94]
port 393 nsew
flabel metal2 s 463946 -960 464058 480 0 FreeSans 560 90 0 0 la_data_out[95]
port 394 nsew
flabel metal2 s 467442 -960 467554 480 0 FreeSans 560 90 0 0 la_data_out[96]
port 395 nsew
flabel metal2 s 471030 -960 471142 480 0 FreeSans 560 90 0 0 la_data_out[97]
port 396 nsew
flabel metal2 s 474526 -960 474638 480 0 FreeSans 560 90 0 0 la_data_out[98]
port 397 nsew
flabel metal2 s 478114 -960 478226 480 0 FreeSans 560 90 0 0 la_data_out[99]
port 398 nsew
flabel metal2 s 158874 -960 158986 480 0 FreeSans 560 90 0 0 la_data_out[9]
port 399 nsew
flabel metal2 s 128146 -960 128258 480 0 FreeSans 560 90 0 0 la_oenb[0]
port 400 nsew
flabel metal2 s 482806 -960 482918 480 0 FreeSans 560 90 0 0 la_oenb[100]
port 401 nsew
flabel metal2 s 486394 -960 486506 480 0 FreeSans 560 90 0 0 la_oenb[101]
port 402 nsew
flabel metal2 s 489890 -960 490002 480 0 FreeSans 560 90 0 0 la_oenb[102]
port 403 nsew
flabel metal2 s 493478 -960 493590 480 0 FreeSans 560 90 0 0 la_oenb[103]
port 404 nsew
flabel metal2 s 497066 -960 497178 480 0 FreeSans 560 90 0 0 la_oenb[104]
port 405 nsew
flabel metal2 s 500562 -960 500674 480 0 FreeSans 560 90 0 0 la_oenb[105]
port 406 nsew
flabel metal2 s 504150 -960 504262 480 0 FreeSans 560 90 0 0 la_oenb[106]
port 407 nsew
flabel metal2 s 507646 -960 507758 480 0 FreeSans 560 90 0 0 la_oenb[107]
port 408 nsew
flabel metal2 s 511234 -960 511346 480 0 FreeSans 560 90 0 0 la_oenb[108]
port 409 nsew
flabel metal2 s 514730 -960 514842 480 0 FreeSans 560 90 0 0 la_oenb[109]
port 410 nsew
flabel metal2 s 163658 -960 163770 480 0 FreeSans 560 90 0 0 la_oenb[10]
port 411 nsew
flabel metal2 s 518318 -960 518430 480 0 FreeSans 560 90 0 0 la_oenb[110]
port 412 nsew
flabel metal2 s 521814 -960 521926 480 0 FreeSans 560 90 0 0 la_oenb[111]
port 413 nsew
flabel metal2 s 525402 -960 525514 480 0 FreeSans 560 90 0 0 la_oenb[112]
port 414 nsew
flabel metal2 s 528990 -960 529102 480 0 FreeSans 560 90 0 0 la_oenb[113]
port 415 nsew
flabel metal2 s 532486 -960 532598 480 0 FreeSans 560 90 0 0 la_oenb[114]
port 416 nsew
flabel metal2 s 536074 -960 536186 480 0 FreeSans 560 90 0 0 la_oenb[115]
port 417 nsew
flabel metal2 s 539570 -960 539682 480 0 FreeSans 560 90 0 0 la_oenb[116]
port 418 nsew
flabel metal2 s 543158 -960 543270 480 0 FreeSans 560 90 0 0 la_oenb[117]
port 419 nsew
flabel metal2 s 546654 -960 546766 480 0 FreeSans 560 90 0 0 la_oenb[118]
port 420 nsew
flabel metal2 s 550242 -960 550354 480 0 FreeSans 560 90 0 0 la_oenb[119]
port 421 nsew
flabel metal2 s 167154 -960 167266 480 0 FreeSans 560 90 0 0 la_oenb[11]
port 422 nsew
flabel metal2 s 553738 -960 553850 480 0 FreeSans 560 90 0 0 la_oenb[120]
port 423 nsew
flabel metal2 s 557326 -960 557438 480 0 FreeSans 560 90 0 0 la_oenb[121]
port 424 nsew
flabel metal2 s 560822 -960 560934 480 0 FreeSans 560 90 0 0 la_oenb[122]
port 425 nsew
flabel metal2 s 564410 -960 564522 480 0 FreeSans 560 90 0 0 la_oenb[123]
port 426 nsew
flabel metal2 s 567998 -960 568110 480 0 FreeSans 560 90 0 0 la_oenb[124]
port 427 nsew
flabel metal2 s 571494 -960 571606 480 0 FreeSans 560 90 0 0 la_oenb[125]
port 428 nsew
flabel metal2 s 575082 -960 575194 480 0 FreeSans 560 90 0 0 la_oenb[126]
port 429 nsew
flabel metal2 s 578578 -960 578690 480 0 FreeSans 560 90 0 0 la_oenb[127]
port 430 nsew
flabel metal2 s 170742 -960 170854 480 0 FreeSans 560 90 0 0 la_oenb[12]
port 431 nsew
flabel metal2 s 174238 -960 174350 480 0 FreeSans 560 90 0 0 la_oenb[13]
port 432 nsew
flabel metal2 s 177826 -960 177938 480 0 FreeSans 560 90 0 0 la_oenb[14]
port 433 nsew
flabel metal2 s 181414 -960 181526 480 0 FreeSans 560 90 0 0 la_oenb[15]
port 434 nsew
flabel metal2 s 184910 -960 185022 480 0 FreeSans 560 90 0 0 la_oenb[16]
port 435 nsew
flabel metal2 s 188498 -960 188610 480 0 FreeSans 560 90 0 0 la_oenb[17]
port 436 nsew
flabel metal2 s 191994 -960 192106 480 0 FreeSans 560 90 0 0 la_oenb[18]
port 437 nsew
flabel metal2 s 195582 -960 195694 480 0 FreeSans 560 90 0 0 la_oenb[19]
port 438 nsew
flabel metal2 s 131734 -960 131846 480 0 FreeSans 560 90 0 0 la_oenb[1]
port 439 nsew
flabel metal2 s 199078 -960 199190 480 0 FreeSans 560 90 0 0 la_oenb[20]
port 440 nsew
flabel metal2 s 202666 -960 202778 480 0 FreeSans 560 90 0 0 la_oenb[21]
port 441 nsew
flabel metal2 s 206162 -960 206274 480 0 FreeSans 560 90 0 0 la_oenb[22]
port 442 nsew
flabel metal2 s 209750 -960 209862 480 0 FreeSans 560 90 0 0 la_oenb[23]
port 443 nsew
flabel metal2 s 213338 -960 213450 480 0 FreeSans 560 90 0 0 la_oenb[24]
port 444 nsew
flabel metal2 s 216834 -960 216946 480 0 FreeSans 560 90 0 0 la_oenb[25]
port 445 nsew
flabel metal2 s 220422 -960 220534 480 0 FreeSans 560 90 0 0 la_oenb[26]
port 446 nsew
flabel metal2 s 223918 -960 224030 480 0 FreeSans 560 90 0 0 la_oenb[27]
port 447 nsew
flabel metal2 s 227506 -960 227618 480 0 FreeSans 560 90 0 0 la_oenb[28]
port 448 nsew
flabel metal2 s 231002 -960 231114 480 0 FreeSans 560 90 0 0 la_oenb[29]
port 449 nsew
flabel metal2 s 135230 -960 135342 480 0 FreeSans 560 90 0 0 la_oenb[2]
port 450 nsew
flabel metal2 s 234590 -960 234702 480 0 FreeSans 560 90 0 0 la_oenb[30]
port 451 nsew
flabel metal2 s 238086 -960 238198 480 0 FreeSans 560 90 0 0 la_oenb[31]
port 452 nsew
flabel metal2 s 241674 -960 241786 480 0 FreeSans 560 90 0 0 la_oenb[32]
port 453 nsew
flabel metal2 s 245170 -960 245282 480 0 FreeSans 560 90 0 0 la_oenb[33]
port 454 nsew
flabel metal2 s 248758 -960 248870 480 0 FreeSans 560 90 0 0 la_oenb[34]
port 455 nsew
flabel metal2 s 252346 -960 252458 480 0 FreeSans 560 90 0 0 la_oenb[35]
port 456 nsew
flabel metal2 s 255842 -960 255954 480 0 FreeSans 560 90 0 0 la_oenb[36]
port 457 nsew
flabel metal2 s 259430 -960 259542 480 0 FreeSans 560 90 0 0 la_oenb[37]
port 458 nsew
flabel metal2 s 262926 -960 263038 480 0 FreeSans 560 90 0 0 la_oenb[38]
port 459 nsew
flabel metal2 s 266514 -960 266626 480 0 FreeSans 560 90 0 0 la_oenb[39]
port 460 nsew
flabel metal2 s 138818 -960 138930 480 0 FreeSans 560 90 0 0 la_oenb[3]
port 461 nsew
flabel metal2 s 270010 -960 270122 480 0 FreeSans 560 90 0 0 la_oenb[40]
port 462 nsew
flabel metal2 s 273598 -960 273710 480 0 FreeSans 560 90 0 0 la_oenb[41]
port 463 nsew
flabel metal2 s 277094 -960 277206 480 0 FreeSans 560 90 0 0 la_oenb[42]
port 464 nsew
flabel metal2 s 280682 -960 280794 480 0 FreeSans 560 90 0 0 la_oenb[43]
port 465 nsew
flabel metal2 s 284270 -960 284382 480 0 FreeSans 560 90 0 0 la_oenb[44]
port 466 nsew
flabel metal2 s 287766 -960 287878 480 0 FreeSans 560 90 0 0 la_oenb[45]
port 467 nsew
flabel metal2 s 291354 -960 291466 480 0 FreeSans 560 90 0 0 la_oenb[46]
port 468 nsew
flabel metal2 s 294850 -960 294962 480 0 FreeSans 560 90 0 0 la_oenb[47]
port 469 nsew
flabel metal2 s 298438 -960 298550 480 0 FreeSans 560 90 0 0 la_oenb[48]
port 470 nsew
flabel metal2 s 301934 -960 302046 480 0 FreeSans 560 90 0 0 la_oenb[49]
port 471 nsew
flabel metal2 s 142406 -960 142518 480 0 FreeSans 560 90 0 0 la_oenb[4]
port 472 nsew
flabel metal2 s 305522 -960 305634 480 0 FreeSans 560 90 0 0 la_oenb[50]
port 473 nsew
flabel metal2 s 309018 -960 309130 480 0 FreeSans 560 90 0 0 la_oenb[51]
port 474 nsew
flabel metal2 s 312606 -960 312718 480 0 FreeSans 560 90 0 0 la_oenb[52]
port 475 nsew
flabel metal2 s 316194 -960 316306 480 0 FreeSans 560 90 0 0 la_oenb[53]
port 476 nsew
flabel metal2 s 319690 -960 319802 480 0 FreeSans 560 90 0 0 la_oenb[54]
port 477 nsew
flabel metal2 s 323278 -960 323390 480 0 FreeSans 560 90 0 0 la_oenb[55]
port 478 nsew
flabel metal2 s 326774 -960 326886 480 0 FreeSans 560 90 0 0 la_oenb[56]
port 479 nsew
flabel metal2 s 330362 -960 330474 480 0 FreeSans 560 90 0 0 la_oenb[57]
port 480 nsew
flabel metal2 s 333858 -960 333970 480 0 FreeSans 560 90 0 0 la_oenb[58]
port 481 nsew
flabel metal2 s 337446 -960 337558 480 0 FreeSans 560 90 0 0 la_oenb[59]
port 482 nsew
flabel metal2 s 145902 -960 146014 480 0 FreeSans 560 90 0 0 la_oenb[5]
port 483 nsew
flabel metal2 s 340942 -960 341054 480 0 FreeSans 560 90 0 0 la_oenb[60]
port 484 nsew
flabel metal2 s 344530 -960 344642 480 0 FreeSans 560 90 0 0 la_oenb[61]
port 485 nsew
flabel metal2 s 348026 -960 348138 480 0 FreeSans 560 90 0 0 la_oenb[62]
port 486 nsew
flabel metal2 s 351614 -960 351726 480 0 FreeSans 560 90 0 0 la_oenb[63]
port 487 nsew
flabel metal2 s 355202 -960 355314 480 0 FreeSans 560 90 0 0 la_oenb[64]
port 488 nsew
flabel metal2 s 358698 -960 358810 480 0 FreeSans 560 90 0 0 la_oenb[65]
port 489 nsew
flabel metal2 s 362286 -960 362398 480 0 FreeSans 560 90 0 0 la_oenb[66]
port 490 nsew
flabel metal2 s 365782 -960 365894 480 0 FreeSans 560 90 0 0 la_oenb[67]
port 491 nsew
flabel metal2 s 369370 -960 369482 480 0 FreeSans 560 90 0 0 la_oenb[68]
port 492 nsew
flabel metal2 s 372866 -960 372978 480 0 FreeSans 560 90 0 0 la_oenb[69]
port 493 nsew
flabel metal2 s 149490 -960 149602 480 0 FreeSans 560 90 0 0 la_oenb[6]
port 494 nsew
flabel metal2 s 376454 -960 376566 480 0 FreeSans 560 90 0 0 la_oenb[70]
port 495 nsew
flabel metal2 s 379950 -960 380062 480 0 FreeSans 560 90 0 0 la_oenb[71]
port 496 nsew
flabel metal2 s 383538 -960 383650 480 0 FreeSans 560 90 0 0 la_oenb[72]
port 497 nsew
flabel metal2 s 387126 -960 387238 480 0 FreeSans 560 90 0 0 la_oenb[73]
port 498 nsew
flabel metal2 s 390622 -960 390734 480 0 FreeSans 560 90 0 0 la_oenb[74]
port 499 nsew
flabel metal2 s 394210 -960 394322 480 0 FreeSans 560 90 0 0 la_oenb[75]
port 500 nsew
flabel metal2 s 397706 -960 397818 480 0 FreeSans 560 90 0 0 la_oenb[76]
port 501 nsew
flabel metal2 s 401294 -960 401406 480 0 FreeSans 560 90 0 0 la_oenb[77]
port 502 nsew
flabel metal2 s 404790 -960 404902 480 0 FreeSans 560 90 0 0 la_oenb[78]
port 503 nsew
flabel metal2 s 408378 -960 408490 480 0 FreeSans 560 90 0 0 la_oenb[79]
port 504 nsew
flabel metal2 s 152986 -960 153098 480 0 FreeSans 560 90 0 0 la_oenb[7]
port 505 nsew
flabel metal2 s 411874 -960 411986 480 0 FreeSans 560 90 0 0 la_oenb[80]
port 506 nsew
flabel metal2 s 415462 -960 415574 480 0 FreeSans 560 90 0 0 la_oenb[81]
port 507 nsew
flabel metal2 s 418958 -960 419070 480 0 FreeSans 560 90 0 0 la_oenb[82]
port 508 nsew
flabel metal2 s 422546 -960 422658 480 0 FreeSans 560 90 0 0 la_oenb[83]
port 509 nsew
flabel metal2 s 426134 -960 426246 480 0 FreeSans 560 90 0 0 la_oenb[84]
port 510 nsew
flabel metal2 s 429630 -960 429742 480 0 FreeSans 560 90 0 0 la_oenb[85]
port 511 nsew
flabel metal2 s 433218 -960 433330 480 0 FreeSans 560 90 0 0 la_oenb[86]
port 512 nsew
flabel metal2 s 436714 -960 436826 480 0 FreeSans 560 90 0 0 la_oenb[87]
port 513 nsew
flabel metal2 s 440302 -960 440414 480 0 FreeSans 560 90 0 0 la_oenb[88]
port 514 nsew
flabel metal2 s 443798 -960 443910 480 0 FreeSans 560 90 0 0 la_oenb[89]
port 515 nsew
flabel metal2 s 156574 -960 156686 480 0 FreeSans 560 90 0 0 la_oenb[8]
port 516 nsew
flabel metal2 s 447386 -960 447498 480 0 FreeSans 560 90 0 0 la_oenb[90]
port 517 nsew
flabel metal2 s 450882 -960 450994 480 0 FreeSans 560 90 0 0 la_oenb[91]
port 518 nsew
flabel metal2 s 454470 -960 454582 480 0 FreeSans 560 90 0 0 la_oenb[92]
port 519 nsew
flabel metal2 s 458058 -960 458170 480 0 FreeSans 560 90 0 0 la_oenb[93]
port 520 nsew
flabel metal2 s 461554 -960 461666 480 0 FreeSans 560 90 0 0 la_oenb[94]
port 521 nsew
flabel metal2 s 465142 -960 465254 480 0 FreeSans 560 90 0 0 la_oenb[95]
port 522 nsew
flabel metal2 s 468638 -960 468750 480 0 FreeSans 560 90 0 0 la_oenb[96]
port 523 nsew
flabel metal2 s 472226 -960 472338 480 0 FreeSans 560 90 0 0 la_oenb[97]
port 524 nsew
flabel metal2 s 475722 -960 475834 480 0 FreeSans 560 90 0 0 la_oenb[98]
port 525 nsew
flabel metal2 s 479310 -960 479422 480 0 FreeSans 560 90 0 0 la_oenb[99]
port 526 nsew
flabel metal2 s 160070 -960 160182 480 0 FreeSans 560 90 0 0 la_oenb[9]
port 527 nsew
flabel metal2 s 579774 -960 579886 480 0 FreeSans 560 90 0 0 user_clock2
port 528 nsew
flabel metal2 s 580970 -960 581082 480 0 FreeSans 560 90 0 0 user_irq[0]
port 529 nsew
flabel metal2 s 582166 -960 582278 480 0 FreeSans 560 90 0 0 user_irq[1]
port 530 nsew
flabel metal2 s 583362 -960 583474 480 0 FreeSans 560 90 0 0 user_irq[2]
port 531 nsew
flabel metal5 s -8726 686066 592650 686686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 650066 592650 650686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 614066 592650 614686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 578066 592650 578686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 542066 592650 542686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 506066 592650 506686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 470066 592650 470686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 434066 592650 434686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 398066 592650 398686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 362066 592650 362686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 326066 592650 326686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 290066 592650 290686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 254066 592650 254686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 218066 592650 218686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 182066 592650 182686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 146066 592650 146686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 110066 592650 110686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 74066 592650 74686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 38066 592650 38686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 2066 592650 2686 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal4 s 576994 -7654 577614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 540994 445572 541614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 540994 -7654 541614 279788 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 504994 -7654 505614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 468994 -7654 469614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 432994 -7654 433614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 396994 -7654 397614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 360994 -7654 361614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 324994 -7654 325614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 288994 -7654 289614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 252994 -7654 253614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 216994 -7654 217614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 180994 -7654 181614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 144994 -7654 145614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 108994 -7654 109614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 72994 -7654 73614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 36994 -7654 37614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 994 -7654 1614 711590 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 3200 0 0 0 vccd1
port 532 nsew
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 4800 90 0 0 vccd1
port 532 nsew
flabel metal5 s -8726 688546 592650 689166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 652546 592650 653166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 616546 592650 617166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 580546 592650 581166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 544546 592650 545166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 508546 592650 509166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 472546 592650 473166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 436546 592650 437166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 400546 592650 401166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 364546 592650 365166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 328546 592650 329166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 292546 592650 293166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 256546 592650 257166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 220546 592650 221166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 184546 592650 185166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 148546 592650 149166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 112546 592650 113166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 76546 592650 77166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 40546 592650 41166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 4546 592650 5166 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal4 s 579474 -7654 580094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 543474 445572 544094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 543474 -7654 544094 279788 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 507474 -7654 508094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 471474 -7654 472094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 435474 -7654 436094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 399474 -7654 400094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 363474 -7654 364094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 327474 -7654 328094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 291474 -7654 292094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 255474 -7654 256094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 219474 -7654 220094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 183474 -7654 184094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 147474 -7654 148094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 111474 -7654 112094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 75474 -7654 76094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 39474 -7654 40094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 3474 -7654 4094 711590 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 3200 0 0 0 vccd2
port 533 nsew
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 4800 90 0 0 vccd2
port 533 nsew
flabel metal5 s -8726 691026 592650 691646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 655026 592650 655646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 619026 592650 619646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 583026 592650 583646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 547026 592650 547646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 511026 592650 511646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 475026 592650 475646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 439026 592650 439646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 403026 592650 403646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 367026 592650 367646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 331026 592650 331646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 295026 592650 295646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 259026 592650 259646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 223026 592650 223646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 187026 592650 187646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 151026 592650 151646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 115026 592650 115646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 79026 592650 79646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 43026 592650 43646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 7026 592650 7646 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal4 s 581954 -7654 582574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 545954 445572 546574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 545954 -7654 546574 279788 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 509954 -7654 510574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 473954 370660 474574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 473954 265660 474574 366216 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 473954 -7654 474574 261216 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 437954 -7654 438574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 401954 -7654 402574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 365954 -7654 366574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 329954 -7654 330574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 293954 -7654 294574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 257954 -7654 258574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 221954 -7654 222574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 185954 -7654 186574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 149954 -7654 150574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 113954 -7654 114574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 77954 -7654 78574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 41954 -7654 42574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 5954 -7654 6574 711590 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 3200 0 0 0 vdda1
port 534 nsew
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 4800 90 0 0 vdda1
port 534 nsew
flabel metal5 s -8726 693506 592650 694126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 657506 592650 658126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 621506 592650 622126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 585506 592650 586126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 549506 592650 550126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 513506 592650 514126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 477506 592650 478126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 441506 592650 442126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 405506 592650 406126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 369506 592650 370126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 333506 592650 334126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 297506 592650 298126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 261506 592650 262126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 225506 592650 226126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 189506 592650 190126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 153506 592650 154126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 117506 592650 118126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 81506 592650 82126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 45506 592650 46126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 9506 592650 10126 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal4 s 548434 -7654 549054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 512434 -7654 513054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 476434 370660 477054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 476434 265660 477054 366216 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 476434 -7654 477054 261216 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 440434 -7654 441054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 404434 -7654 405054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 368434 -7654 369054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 332434 -7654 333054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 296434 -7654 297054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 260434 -7654 261054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 224434 -7654 225054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 188434 -7654 189054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 152434 -7654 153054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 116434 -7654 117054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 80434 -7654 81054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 44434 -7654 45054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 8434 -7654 9054 711590 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 3200 0 0 0 vdda2
port 535 nsew
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 4800 90 0 0 vdda2
port 535 nsew
flabel metal5 s -8726 692266 592650 692886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 656266 592650 656886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 620266 592650 620886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 584266 592650 584886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 548266 592650 548886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 512266 592650 512886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 476266 592650 476886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 440266 592650 440886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 404266 592650 404886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 368266 592650 368886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 332266 592650 332886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 296266 592650 296886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 260266 592650 260886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 224266 592650 224886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 188266 592650 188886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 152266 592650 152886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 116266 592650 116886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 80266 592650 80886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 44266 592650 44886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 8266 592650 8886 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal4 s 547194 -7654 547814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 511194 -7654 511814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 475194 370660 475814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 475194 265660 475814 366216 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 475194 -7654 475814 261216 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 439194 -7654 439814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 403194 -7654 403814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 367194 -7654 367814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 331194 -7654 331814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 295194 -7654 295814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 259194 -7654 259814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 223194 -7654 223814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 187194 -7654 187814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 151194 -7654 151814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 115194 -7654 115814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 79194 -7654 79814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 43194 -7654 43814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 7194 -7654 7814 711590 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 3200 0 0 0 vssa1
port 536 nsew
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 4800 90 0 0 vssa1
port 536 nsew
flabel metal5 s -8726 694746 592650 695366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 658746 592650 659366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 622746 592650 623366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 586746 592650 587366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 550746 592650 551366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 514746 592650 515366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 478746 592650 479366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 442746 592650 443366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 406746 592650 407366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 370746 592650 371366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 334746 592650 335366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 298746 592650 299366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 262746 592650 263366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 226746 592650 227366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 190746 592650 191366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 154746 592650 155366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 118746 592650 119366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 82746 592650 83366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 46746 592650 47366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 10746 592650 11366 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal4 s 549674 -7654 550294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 513674 -7654 514294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 477674 370660 478294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 477674 265660 478294 366216 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 477674 -7654 478294 261216 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 441674 -7654 442294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 405674 -7654 406294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 369674 -7654 370294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 333674 -7654 334294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 297674 -7654 298294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 261674 -7654 262294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 225674 -7654 226294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 189674 -7654 190294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 153674 -7654 154294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 117674 -7654 118294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 81674 -7654 82294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 45674 -7654 46294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 9674 -7654 10294 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 3200 0 0 0 vssa2
port 537 nsew
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 4800 90 0 0 vssa2
port 537 nsew
flabel metal5 s -8726 687306 592650 687926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 651306 592650 651926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 615306 592650 615926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 579306 592650 579926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 543306 592650 543926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 507306 592650 507926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 471306 592650 471926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 435306 592650 435926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 399306 592650 399926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 363306 592650 363926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 327306 592650 327926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 291306 592650 291926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 255306 592650 255926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 219306 592650 219926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 183306 592650 183926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 147306 592650 147926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 111306 592650 111926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 75306 592650 75926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 39306 592650 39926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 3306 592650 3926 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal4 s 578234 -7654 578854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 542234 445572 542854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 542234 -7654 542854 279788 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 506234 -7654 506854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 470234 -7654 470854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 434234 -7654 434854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 398234 -7654 398854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 362234 -7654 362854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 326234 -7654 326854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 290234 -7654 290854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 254234 -7654 254854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 218234 -7654 218854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 182234 -7654 182854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 146234 -7654 146854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 110234 -7654 110854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 74234 -7654 74854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 38234 -7654 38854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 2234 -7654 2854 711590 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 3200 0 0 0 vssd1
port 538 nsew
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 4800 90 0 0 vssd1
port 538 nsew
flabel metal5 s -8726 689786 592650 690406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 653786 592650 654406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 617786 592650 618406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 581786 592650 582406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 545786 592650 546406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 509786 592650 510406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 473786 592650 474406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 437786 592650 438406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 401786 592650 402406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 365786 592650 366406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 329786 592650 330406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 293786 592650 294406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 257786 592650 258406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 221786 592650 222406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 185786 592650 186406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 149786 592650 150406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 113786 592650 114406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 77786 592650 78406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 41786 592650 42406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -8726 5786 592650 6406 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal4 s 580714 -7654 581334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 544714 445572 545334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 544714 -7654 545334 279788 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 508714 -7654 509334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 472714 370660 473334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 472714 265660 473334 366216 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 472714 -7654 473334 261216 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 436714 -7654 437334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 400714 -7654 401334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 364714 -7654 365334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 328714 -7654 329334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 292714 -7654 293334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 256714 -7654 257334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 220714 -7654 221334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 184714 -7654 185334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 148714 -7654 149334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 112714 -7654 113334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 76714 -7654 77334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 40714 -7654 41334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 4714 -7654 5334 711590 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 3200 0 0 0 vssd2
port 539 nsew
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 4800 90 0 0 vssd2
port 539 nsew
flabel metal2 s 542 -960 654 480 0 FreeSans 560 90 0 0 wb_clk_i
port 540 nsew
flabel metal2 s 1646 -960 1758 480 0 FreeSans 560 90 0 0 wb_rst_i
port 541 nsew
flabel metal2 s 2842 -960 2954 480 0 FreeSans 560 90 0 0 wbs_ack_o
port 542 nsew
flabel metal2 s 7626 -960 7738 480 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 543 nsew
flabel metal2 s 47830 -960 47942 480 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 544 nsew
flabel metal2 s 51326 -960 51438 480 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 545 nsew
flabel metal2 s 54914 -960 55026 480 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 546 nsew
flabel metal2 s 58410 -960 58522 480 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 547 nsew
flabel metal2 s 61998 -960 62110 480 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 548 nsew
flabel metal2 s 65494 -960 65606 480 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 549 nsew
flabel metal2 s 69082 -960 69194 480 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 550 nsew
flabel metal2 s 72578 -960 72690 480 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 551 nsew
flabel metal2 s 76166 -960 76278 480 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 552 nsew
flabel metal2 s 79662 -960 79774 480 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 553 nsew
flabel metal2 s 12318 -960 12430 480 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 554 nsew
flabel metal2 s 83250 -960 83362 480 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 555 nsew
flabel metal2 s 86838 -960 86950 480 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 556 nsew
flabel metal2 s 90334 -960 90446 480 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 557 nsew
flabel metal2 s 93922 -960 94034 480 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 558 nsew
flabel metal2 s 97418 -960 97530 480 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 559 nsew
flabel metal2 s 101006 -960 101118 480 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 560 nsew
flabel metal2 s 104502 -960 104614 480 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 561 nsew
flabel metal2 s 108090 -960 108202 480 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 562 nsew
flabel metal2 s 111586 -960 111698 480 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 563 nsew
flabel metal2 s 115174 -960 115286 480 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 564 nsew
flabel metal2 s 17010 -960 17122 480 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 565 nsew
flabel metal2 s 118762 -960 118874 480 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 566 nsew
flabel metal2 s 122258 -960 122370 480 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 567 nsew
flabel metal2 s 21794 -960 21906 480 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 568 nsew
flabel metal2 s 26486 -960 26598 480 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 569 nsew
flabel metal2 s 30074 -960 30186 480 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 570 nsew
flabel metal2 s 33570 -960 33682 480 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 571 nsew
flabel metal2 s 37158 -960 37270 480 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 572 nsew
flabel metal2 s 40654 -960 40766 480 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 573 nsew
flabel metal2 s 44242 -960 44354 480 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 574 nsew
flabel metal2 s 4038 -960 4150 480 0 FreeSans 560 90 0 0 wbs_cyc_i
port 575 nsew
flabel metal2 s 8730 -960 8842 480 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 576 nsew
flabel metal2 s 48934 -960 49046 480 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 577 nsew
flabel metal2 s 52522 -960 52634 480 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 578 nsew
flabel metal2 s 56018 -960 56130 480 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 579 nsew
flabel metal2 s 59606 -960 59718 480 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 580 nsew
flabel metal2 s 63194 -960 63306 480 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 581 nsew
flabel metal2 s 66690 -960 66802 480 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 582 nsew
flabel metal2 s 70278 -960 70390 480 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 583 nsew
flabel metal2 s 73774 -960 73886 480 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 584 nsew
flabel metal2 s 77362 -960 77474 480 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 585 nsew
flabel metal2 s 80858 -960 80970 480 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 586 nsew
flabel metal2 s 13514 -960 13626 480 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 587 nsew
flabel metal2 s 84446 -960 84558 480 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 588 nsew
flabel metal2 s 87942 -960 88054 480 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 589 nsew
flabel metal2 s 91530 -960 91642 480 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 590 nsew
flabel metal2 s 95118 -960 95230 480 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 591 nsew
flabel metal2 s 98614 -960 98726 480 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 592 nsew
flabel metal2 s 102202 -960 102314 480 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 593 nsew
flabel metal2 s 105698 -960 105810 480 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 594 nsew
flabel metal2 s 109286 -960 109398 480 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 595 nsew
flabel metal2 s 112782 -960 112894 480 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 596 nsew
flabel metal2 s 116370 -960 116482 480 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 597 nsew
flabel metal2 s 18206 -960 18318 480 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 598 nsew
flabel metal2 s 119866 -960 119978 480 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 599 nsew
flabel metal2 s 123454 -960 123566 480 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 600 nsew
flabel metal2 s 22990 -960 23102 480 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 601 nsew
flabel metal2 s 27682 -960 27794 480 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 602 nsew
flabel metal2 s 31270 -960 31382 480 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 603 nsew
flabel metal2 s 34766 -960 34878 480 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 604 nsew
flabel metal2 s 38354 -960 38466 480 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 605 nsew
flabel metal2 s 41850 -960 41962 480 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 606 nsew
flabel metal2 s 45438 -960 45550 480 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 607 nsew
flabel metal2 s 9926 -960 10038 480 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 608 nsew
flabel metal2 s 50130 -960 50242 480 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 609 nsew
flabel metal2 s 53718 -960 53830 480 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 610 nsew
flabel metal2 s 57214 -960 57326 480 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 611 nsew
flabel metal2 s 60802 -960 60914 480 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 612 nsew
flabel metal2 s 64298 -960 64410 480 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 613 nsew
flabel metal2 s 67886 -960 67998 480 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 614 nsew
flabel metal2 s 71474 -960 71586 480 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 615 nsew
flabel metal2 s 74970 -960 75082 480 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 616 nsew
flabel metal2 s 78558 -960 78670 480 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 617 nsew
flabel metal2 s 82054 -960 82166 480 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 618 nsew
flabel metal2 s 14710 -960 14822 480 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 619 nsew
flabel metal2 s 85642 -960 85754 480 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 620 nsew
flabel metal2 s 89138 -960 89250 480 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 621 nsew
flabel metal2 s 92726 -960 92838 480 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 622 nsew
flabel metal2 s 96222 -960 96334 480 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 623 nsew
flabel metal2 s 99810 -960 99922 480 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 624 nsew
flabel metal2 s 103306 -960 103418 480 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 625 nsew
flabel metal2 s 106894 -960 107006 480 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 626 nsew
flabel metal2 s 110482 -960 110594 480 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 627 nsew
flabel metal2 s 113978 -960 114090 480 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 628 nsew
flabel metal2 s 117566 -960 117678 480 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 629 nsew
flabel metal2 s 19402 -960 19514 480 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 630 nsew
flabel metal2 s 121062 -960 121174 480 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 631 nsew
flabel metal2 s 124650 -960 124762 480 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 632 nsew
flabel metal2 s 24186 -960 24298 480 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 633 nsew
flabel metal2 s 28878 -960 28990 480 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 634 nsew
flabel metal2 s 32374 -960 32486 480 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 635 nsew
flabel metal2 s 35962 -960 36074 480 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 636 nsew
flabel metal2 s 39550 -960 39662 480 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 637 nsew
flabel metal2 s 43046 -960 43158 480 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 638 nsew
flabel metal2 s 46634 -960 46746 480 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 639 nsew
flabel metal2 s 11122 -960 11234 480 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 640 nsew
flabel metal2 s 15906 -960 16018 480 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 641 nsew
flabel metal2 s 20598 -960 20710 480 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 642 nsew
flabel metal2 s 25290 -960 25402 480 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 643 nsew
flabel metal2 s 5234 -960 5346 480 0 FreeSans 560 90 0 0 wbs_stb_i
port 644 nsew
flabel metal2 s 6430 -960 6542 480 0 FreeSans 560 90 0 0 wbs_we_i
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
